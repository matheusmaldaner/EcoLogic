library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(10239 downto 0);
    signal layer1_outputs: std_logic_vector(10239 downto 0);
    signal layer2_outputs: std_logic_vector(10239 downto 0);
    signal layer3_outputs: std_logic_vector(10239 downto 0);
    signal layer4_outputs: std_logic_vector(10239 downto 0);

begin
    layer0_outputs(0) <= not b or a;
    layer0_outputs(1) <= a and b;
    layer0_outputs(2) <= 1'b0;
    layer0_outputs(3) <= a and b;
    layer0_outputs(4) <= not b;
    layer0_outputs(5) <= not (a or b);
    layer0_outputs(6) <= not a or b;
    layer0_outputs(7) <= not a;
    layer0_outputs(8) <= not a;
    layer0_outputs(9) <= not (a and b);
    layer0_outputs(10) <= a and not b;
    layer0_outputs(11) <= not a or b;
    layer0_outputs(12) <= not b or a;
    layer0_outputs(13) <= a xor b;
    layer0_outputs(14) <= not a or b;
    layer0_outputs(15) <= a;
    layer0_outputs(16) <= b;
    layer0_outputs(17) <= not b;
    layer0_outputs(18) <= a xor b;
    layer0_outputs(19) <= b;
    layer0_outputs(20) <= a and not b;
    layer0_outputs(21) <= a;
    layer0_outputs(22) <= a or b;
    layer0_outputs(23) <= not a;
    layer0_outputs(24) <= a and not b;
    layer0_outputs(25) <= a xor b;
    layer0_outputs(26) <= not b;
    layer0_outputs(27) <= not a or b;
    layer0_outputs(28) <= not a or b;
    layer0_outputs(29) <= a or b;
    layer0_outputs(30) <= b;
    layer0_outputs(31) <= 1'b0;
    layer0_outputs(32) <= not b;
    layer0_outputs(33) <= not (a or b);
    layer0_outputs(34) <= a xor b;
    layer0_outputs(35) <= not (a xor b);
    layer0_outputs(36) <= not (a xor b);
    layer0_outputs(37) <= not b or a;
    layer0_outputs(38) <= not (a or b);
    layer0_outputs(39) <= a;
    layer0_outputs(40) <= not a;
    layer0_outputs(41) <= not (a and b);
    layer0_outputs(42) <= a or b;
    layer0_outputs(43) <= not (a xor b);
    layer0_outputs(44) <= not (a and b);
    layer0_outputs(45) <= not a;
    layer0_outputs(46) <= a xor b;
    layer0_outputs(47) <= not (a and b);
    layer0_outputs(48) <= not b;
    layer0_outputs(49) <= 1'b1;
    layer0_outputs(50) <= not a;
    layer0_outputs(51) <= not b;
    layer0_outputs(52) <= b;
    layer0_outputs(53) <= not a;
    layer0_outputs(54) <= a or b;
    layer0_outputs(55) <= a and b;
    layer0_outputs(56) <= a and b;
    layer0_outputs(57) <= a or b;
    layer0_outputs(58) <= a or b;
    layer0_outputs(59) <= not (a xor b);
    layer0_outputs(60) <= not a;
    layer0_outputs(61) <= not (a xor b);
    layer0_outputs(62) <= b;
    layer0_outputs(63) <= b and not a;
    layer0_outputs(64) <= not b;
    layer0_outputs(65) <= b;
    layer0_outputs(66) <= not (a or b);
    layer0_outputs(67) <= a and not b;
    layer0_outputs(68) <= b;
    layer0_outputs(69) <= not (a xor b);
    layer0_outputs(70) <= not b or a;
    layer0_outputs(71) <= a xor b;
    layer0_outputs(72) <= a and not b;
    layer0_outputs(73) <= not (a xor b);
    layer0_outputs(74) <= not b;
    layer0_outputs(75) <= not (a or b);
    layer0_outputs(76) <= not a;
    layer0_outputs(77) <= not a;
    layer0_outputs(78) <= 1'b0;
    layer0_outputs(79) <= not (a xor b);
    layer0_outputs(80) <= a or b;
    layer0_outputs(81) <= a and b;
    layer0_outputs(82) <= not b;
    layer0_outputs(83) <= not (a xor b);
    layer0_outputs(84) <= not (a and b);
    layer0_outputs(85) <= b;
    layer0_outputs(86) <= 1'b1;
    layer0_outputs(87) <= not (a xor b);
    layer0_outputs(88) <= not a;
    layer0_outputs(89) <= not b;
    layer0_outputs(90) <= a xor b;
    layer0_outputs(91) <= not a or b;
    layer0_outputs(92) <= a or b;
    layer0_outputs(93) <= a and b;
    layer0_outputs(94) <= not a or b;
    layer0_outputs(95) <= not b;
    layer0_outputs(96) <= b and not a;
    layer0_outputs(97) <= not a or b;
    layer0_outputs(98) <= a or b;
    layer0_outputs(99) <= a xor b;
    layer0_outputs(100) <= 1'b1;
    layer0_outputs(101) <= not (a or b);
    layer0_outputs(102) <= 1'b1;
    layer0_outputs(103) <= a and b;
    layer0_outputs(104) <= not (a xor b);
    layer0_outputs(105) <= not b or a;
    layer0_outputs(106) <= not (a xor b);
    layer0_outputs(107) <= not (a xor b);
    layer0_outputs(108) <= a;
    layer0_outputs(109) <= not (a or b);
    layer0_outputs(110) <= a and b;
    layer0_outputs(111) <= not a or b;
    layer0_outputs(112) <= not b;
    layer0_outputs(113) <= not (a or b);
    layer0_outputs(114) <= b and not a;
    layer0_outputs(115) <= not a or b;
    layer0_outputs(116) <= not (a xor b);
    layer0_outputs(117) <= not (a or b);
    layer0_outputs(118) <= a xor b;
    layer0_outputs(119) <= not b;
    layer0_outputs(120) <= not (a xor b);
    layer0_outputs(121) <= a;
    layer0_outputs(122) <= b and not a;
    layer0_outputs(123) <= b and not a;
    layer0_outputs(124) <= not a;
    layer0_outputs(125) <= a or b;
    layer0_outputs(126) <= not (a or b);
    layer0_outputs(127) <= a xor b;
    layer0_outputs(128) <= not (a and b);
    layer0_outputs(129) <= not (a or b);
    layer0_outputs(130) <= b and not a;
    layer0_outputs(131) <= not (a xor b);
    layer0_outputs(132) <= not a;
    layer0_outputs(133) <= a;
    layer0_outputs(134) <= not (a or b);
    layer0_outputs(135) <= not a or b;
    layer0_outputs(136) <= not b;
    layer0_outputs(137) <= a or b;
    layer0_outputs(138) <= a and b;
    layer0_outputs(139) <= 1'b0;
    layer0_outputs(140) <= not a;
    layer0_outputs(141) <= b;
    layer0_outputs(142) <= not a or b;
    layer0_outputs(143) <= a;
    layer0_outputs(144) <= a and not b;
    layer0_outputs(145) <= a and b;
    layer0_outputs(146) <= 1'b0;
    layer0_outputs(147) <= not a or b;
    layer0_outputs(148) <= 1'b0;
    layer0_outputs(149) <= b and not a;
    layer0_outputs(150) <= a and b;
    layer0_outputs(151) <= not b;
    layer0_outputs(152) <= 1'b1;
    layer0_outputs(153) <= 1'b1;
    layer0_outputs(154) <= not a;
    layer0_outputs(155) <= not (a or b);
    layer0_outputs(156) <= a or b;
    layer0_outputs(157) <= not (a xor b);
    layer0_outputs(158) <= not (a or b);
    layer0_outputs(159) <= not a;
    layer0_outputs(160) <= a or b;
    layer0_outputs(161) <= 1'b0;
    layer0_outputs(162) <= not (a and b);
    layer0_outputs(163) <= not (a or b);
    layer0_outputs(164) <= a xor b;
    layer0_outputs(165) <= a;
    layer0_outputs(166) <= not b or a;
    layer0_outputs(167) <= not (a xor b);
    layer0_outputs(168) <= not b or a;
    layer0_outputs(169) <= not b or a;
    layer0_outputs(170) <= not b or a;
    layer0_outputs(171) <= not a;
    layer0_outputs(172) <= not (a or b);
    layer0_outputs(173) <= not a or b;
    layer0_outputs(174) <= not b or a;
    layer0_outputs(175) <= not a;
    layer0_outputs(176) <= b and not a;
    layer0_outputs(177) <= not b;
    layer0_outputs(178) <= not (a or b);
    layer0_outputs(179) <= a or b;
    layer0_outputs(180) <= b and not a;
    layer0_outputs(181) <= a or b;
    layer0_outputs(182) <= a xor b;
    layer0_outputs(183) <= not a or b;
    layer0_outputs(184) <= a or b;
    layer0_outputs(185) <= not b or a;
    layer0_outputs(186) <= a or b;
    layer0_outputs(187) <= not a or b;
    layer0_outputs(188) <= b;
    layer0_outputs(189) <= not (a xor b);
    layer0_outputs(190) <= not b;
    layer0_outputs(191) <= not a;
    layer0_outputs(192) <= a or b;
    layer0_outputs(193) <= a xor b;
    layer0_outputs(194) <= not (a xor b);
    layer0_outputs(195) <= not (a xor b);
    layer0_outputs(196) <= a and b;
    layer0_outputs(197) <= a and b;
    layer0_outputs(198) <= not (a or b);
    layer0_outputs(199) <= not (a and b);
    layer0_outputs(200) <= not (a and b);
    layer0_outputs(201) <= not b or a;
    layer0_outputs(202) <= a xor b;
    layer0_outputs(203) <= not a;
    layer0_outputs(204) <= not a;
    layer0_outputs(205) <= not (a xor b);
    layer0_outputs(206) <= a xor b;
    layer0_outputs(207) <= b and not a;
    layer0_outputs(208) <= not a;
    layer0_outputs(209) <= not a;
    layer0_outputs(210) <= not b;
    layer0_outputs(211) <= not b or a;
    layer0_outputs(212) <= not (a or b);
    layer0_outputs(213) <= not b;
    layer0_outputs(214) <= a or b;
    layer0_outputs(215) <= not (a xor b);
    layer0_outputs(216) <= not (a and b);
    layer0_outputs(217) <= not b;
    layer0_outputs(218) <= a and not b;
    layer0_outputs(219) <= not (a xor b);
    layer0_outputs(220) <= a;
    layer0_outputs(221) <= not (a or b);
    layer0_outputs(222) <= a and not b;
    layer0_outputs(223) <= not b or a;
    layer0_outputs(224) <= not b;
    layer0_outputs(225) <= b;
    layer0_outputs(226) <= not a or b;
    layer0_outputs(227) <= not (a or b);
    layer0_outputs(228) <= not (a or b);
    layer0_outputs(229) <= a and not b;
    layer0_outputs(230) <= not b or a;
    layer0_outputs(231) <= not (a or b);
    layer0_outputs(232) <= not b or a;
    layer0_outputs(233) <= not (a xor b);
    layer0_outputs(234) <= b;
    layer0_outputs(235) <= not (a and b);
    layer0_outputs(236) <= not b;
    layer0_outputs(237) <= a xor b;
    layer0_outputs(238) <= a xor b;
    layer0_outputs(239) <= a and not b;
    layer0_outputs(240) <= not a;
    layer0_outputs(241) <= not (a or b);
    layer0_outputs(242) <= 1'b0;
    layer0_outputs(243) <= not b or a;
    layer0_outputs(244) <= not b;
    layer0_outputs(245) <= b and not a;
    layer0_outputs(246) <= 1'b0;
    layer0_outputs(247) <= b and not a;
    layer0_outputs(248) <= not (a or b);
    layer0_outputs(249) <= not a or b;
    layer0_outputs(250) <= not a;
    layer0_outputs(251) <= a or b;
    layer0_outputs(252) <= a;
    layer0_outputs(253) <= a and not b;
    layer0_outputs(254) <= b;
    layer0_outputs(255) <= a xor b;
    layer0_outputs(256) <= a and not b;
    layer0_outputs(257) <= a xor b;
    layer0_outputs(258) <= b and not a;
    layer0_outputs(259) <= not b;
    layer0_outputs(260) <= not b or a;
    layer0_outputs(261) <= b;
    layer0_outputs(262) <= b and not a;
    layer0_outputs(263) <= 1'b0;
    layer0_outputs(264) <= 1'b1;
    layer0_outputs(265) <= 1'b0;
    layer0_outputs(266) <= not (a xor b);
    layer0_outputs(267) <= b and not a;
    layer0_outputs(268) <= not (a xor b);
    layer0_outputs(269) <= not (a or b);
    layer0_outputs(270) <= not (a and b);
    layer0_outputs(271) <= not b;
    layer0_outputs(272) <= not (a or b);
    layer0_outputs(273) <= a xor b;
    layer0_outputs(274) <= not b or a;
    layer0_outputs(275) <= not b;
    layer0_outputs(276) <= 1'b1;
    layer0_outputs(277) <= not (a or b);
    layer0_outputs(278) <= a;
    layer0_outputs(279) <= b;
    layer0_outputs(280) <= not a;
    layer0_outputs(281) <= a or b;
    layer0_outputs(282) <= a or b;
    layer0_outputs(283) <= not (a or b);
    layer0_outputs(284) <= 1'b1;
    layer0_outputs(285) <= a or b;
    layer0_outputs(286) <= not (a xor b);
    layer0_outputs(287) <= not b or a;
    layer0_outputs(288) <= a xor b;
    layer0_outputs(289) <= not a or b;
    layer0_outputs(290) <= not (a xor b);
    layer0_outputs(291) <= a;
    layer0_outputs(292) <= a or b;
    layer0_outputs(293) <= not a;
    layer0_outputs(294) <= not a;
    layer0_outputs(295) <= a xor b;
    layer0_outputs(296) <= a;
    layer0_outputs(297) <= b;
    layer0_outputs(298) <= not (a and b);
    layer0_outputs(299) <= not (a or b);
    layer0_outputs(300) <= a xor b;
    layer0_outputs(301) <= b;
    layer0_outputs(302) <= b;
    layer0_outputs(303) <= a xor b;
    layer0_outputs(304) <= not a;
    layer0_outputs(305) <= b and not a;
    layer0_outputs(306) <= a and not b;
    layer0_outputs(307) <= a or b;
    layer0_outputs(308) <= 1'b0;
    layer0_outputs(309) <= a or b;
    layer0_outputs(310) <= not b or a;
    layer0_outputs(311) <= 1'b0;
    layer0_outputs(312) <= b;
    layer0_outputs(313) <= a and not b;
    layer0_outputs(314) <= a or b;
    layer0_outputs(315) <= not b;
    layer0_outputs(316) <= a and b;
    layer0_outputs(317) <= a xor b;
    layer0_outputs(318) <= b;
    layer0_outputs(319) <= a and not b;
    layer0_outputs(320) <= not b;
    layer0_outputs(321) <= a and not b;
    layer0_outputs(322) <= not b;
    layer0_outputs(323) <= not a;
    layer0_outputs(324) <= not (a or b);
    layer0_outputs(325) <= 1'b0;
    layer0_outputs(326) <= a or b;
    layer0_outputs(327) <= not (a or b);
    layer0_outputs(328) <= b;
    layer0_outputs(329) <= a xor b;
    layer0_outputs(330) <= a or b;
    layer0_outputs(331) <= a and not b;
    layer0_outputs(332) <= b;
    layer0_outputs(333) <= not a;
    layer0_outputs(334) <= not b;
    layer0_outputs(335) <= not (a xor b);
    layer0_outputs(336) <= not b;
    layer0_outputs(337) <= a and not b;
    layer0_outputs(338) <= not a;
    layer0_outputs(339) <= not b;
    layer0_outputs(340) <= not b or a;
    layer0_outputs(341) <= not b or a;
    layer0_outputs(342) <= not (a or b);
    layer0_outputs(343) <= a and not b;
    layer0_outputs(344) <= b and not a;
    layer0_outputs(345) <= not a;
    layer0_outputs(346) <= not b;
    layer0_outputs(347) <= b and not a;
    layer0_outputs(348) <= not a or b;
    layer0_outputs(349) <= b;
    layer0_outputs(350) <= 1'b0;
    layer0_outputs(351) <= not b or a;
    layer0_outputs(352) <= a xor b;
    layer0_outputs(353) <= b and not a;
    layer0_outputs(354) <= a;
    layer0_outputs(355) <= b and not a;
    layer0_outputs(356) <= a or b;
    layer0_outputs(357) <= b;
    layer0_outputs(358) <= a or b;
    layer0_outputs(359) <= not (a or b);
    layer0_outputs(360) <= a xor b;
    layer0_outputs(361) <= a or b;
    layer0_outputs(362) <= not a or b;
    layer0_outputs(363) <= not (a or b);
    layer0_outputs(364) <= b;
    layer0_outputs(365) <= not a;
    layer0_outputs(366) <= not b;
    layer0_outputs(367) <= not a;
    layer0_outputs(368) <= a and b;
    layer0_outputs(369) <= a and not b;
    layer0_outputs(370) <= a xor b;
    layer0_outputs(371) <= a or b;
    layer0_outputs(372) <= not (a xor b);
    layer0_outputs(373) <= a or b;
    layer0_outputs(374) <= not a or b;
    layer0_outputs(375) <= not b;
    layer0_outputs(376) <= b and not a;
    layer0_outputs(377) <= not a;
    layer0_outputs(378) <= not (a and b);
    layer0_outputs(379) <= a and b;
    layer0_outputs(380) <= a xor b;
    layer0_outputs(381) <= b and not a;
    layer0_outputs(382) <= 1'b0;
    layer0_outputs(383) <= not b or a;
    layer0_outputs(384) <= not a;
    layer0_outputs(385) <= b;
    layer0_outputs(386) <= a and b;
    layer0_outputs(387) <= not b or a;
    layer0_outputs(388) <= not b;
    layer0_outputs(389) <= not (a or b);
    layer0_outputs(390) <= a and b;
    layer0_outputs(391) <= not a or b;
    layer0_outputs(392) <= not (a or b);
    layer0_outputs(393) <= a and not b;
    layer0_outputs(394) <= not a;
    layer0_outputs(395) <= a or b;
    layer0_outputs(396) <= a and not b;
    layer0_outputs(397) <= not a or b;
    layer0_outputs(398) <= not b;
    layer0_outputs(399) <= not b or a;
    layer0_outputs(400) <= a xor b;
    layer0_outputs(401) <= not a;
    layer0_outputs(402) <= not b;
    layer0_outputs(403) <= not (a or b);
    layer0_outputs(404) <= a or b;
    layer0_outputs(405) <= a and b;
    layer0_outputs(406) <= not b or a;
    layer0_outputs(407) <= not (a xor b);
    layer0_outputs(408) <= a or b;
    layer0_outputs(409) <= a;
    layer0_outputs(410) <= not a;
    layer0_outputs(411) <= not (a or b);
    layer0_outputs(412) <= b and not a;
    layer0_outputs(413) <= not b;
    layer0_outputs(414) <= b and not a;
    layer0_outputs(415) <= not (a or b);
    layer0_outputs(416) <= not (a xor b);
    layer0_outputs(417) <= 1'b0;
    layer0_outputs(418) <= a;
    layer0_outputs(419) <= not (a or b);
    layer0_outputs(420) <= not a;
    layer0_outputs(421) <= b;
    layer0_outputs(422) <= a or b;
    layer0_outputs(423) <= not a or b;
    layer0_outputs(424) <= a;
    layer0_outputs(425) <= b and not a;
    layer0_outputs(426) <= a and b;
    layer0_outputs(427) <= not (a xor b);
    layer0_outputs(428) <= a or b;
    layer0_outputs(429) <= not a or b;
    layer0_outputs(430) <= not b;
    layer0_outputs(431) <= 1'b1;
    layer0_outputs(432) <= not a or b;
    layer0_outputs(433) <= not (a or b);
    layer0_outputs(434) <= 1'b0;
    layer0_outputs(435) <= not (a or b);
    layer0_outputs(436) <= not (a or b);
    layer0_outputs(437) <= not (a or b);
    layer0_outputs(438) <= not (a or b);
    layer0_outputs(439) <= b and not a;
    layer0_outputs(440) <= a or b;
    layer0_outputs(441) <= not b or a;
    layer0_outputs(442) <= b;
    layer0_outputs(443) <= a or b;
    layer0_outputs(444) <= not b;
    layer0_outputs(445) <= not (a or b);
    layer0_outputs(446) <= not (a or b);
    layer0_outputs(447) <= a and b;
    layer0_outputs(448) <= not (a or b);
    layer0_outputs(449) <= a xor b;
    layer0_outputs(450) <= a and b;
    layer0_outputs(451) <= b and not a;
    layer0_outputs(452) <= a;
    layer0_outputs(453) <= not (a and b);
    layer0_outputs(454) <= a or b;
    layer0_outputs(455) <= a;
    layer0_outputs(456) <= a and b;
    layer0_outputs(457) <= 1'b1;
    layer0_outputs(458) <= b and not a;
    layer0_outputs(459) <= not (a or b);
    layer0_outputs(460) <= not (a xor b);
    layer0_outputs(461) <= not (a or b);
    layer0_outputs(462) <= a;
    layer0_outputs(463) <= b;
    layer0_outputs(464) <= 1'b1;
    layer0_outputs(465) <= a and not b;
    layer0_outputs(466) <= a xor b;
    layer0_outputs(467) <= b;
    layer0_outputs(468) <= a xor b;
    layer0_outputs(469) <= a or b;
    layer0_outputs(470) <= not (a xor b);
    layer0_outputs(471) <= b;
    layer0_outputs(472) <= not b or a;
    layer0_outputs(473) <= a or b;
    layer0_outputs(474) <= b and not a;
    layer0_outputs(475) <= not b;
    layer0_outputs(476) <= not b;
    layer0_outputs(477) <= not (a xor b);
    layer0_outputs(478) <= a or b;
    layer0_outputs(479) <= not a;
    layer0_outputs(480) <= b and not a;
    layer0_outputs(481) <= a xor b;
    layer0_outputs(482) <= b;
    layer0_outputs(483) <= a or b;
    layer0_outputs(484) <= a and b;
    layer0_outputs(485) <= not a or b;
    layer0_outputs(486) <= not a or b;
    layer0_outputs(487) <= 1'b1;
    layer0_outputs(488) <= not (a xor b);
    layer0_outputs(489) <= b and not a;
    layer0_outputs(490) <= not a or b;
    layer0_outputs(491) <= not (a or b);
    layer0_outputs(492) <= not b;
    layer0_outputs(493) <= not a or b;
    layer0_outputs(494) <= not b;
    layer0_outputs(495) <= a or b;
    layer0_outputs(496) <= not b;
    layer0_outputs(497) <= b;
    layer0_outputs(498) <= b;
    layer0_outputs(499) <= b and not a;
    layer0_outputs(500) <= not b or a;
    layer0_outputs(501) <= a or b;
    layer0_outputs(502) <= 1'b1;
    layer0_outputs(503) <= 1'b0;
    layer0_outputs(504) <= not (a xor b);
    layer0_outputs(505) <= b;
    layer0_outputs(506) <= a or b;
    layer0_outputs(507) <= a;
    layer0_outputs(508) <= not b;
    layer0_outputs(509) <= b;
    layer0_outputs(510) <= a xor b;
    layer0_outputs(511) <= not b or a;
    layer0_outputs(512) <= a or b;
    layer0_outputs(513) <= a or b;
    layer0_outputs(514) <= not (a and b);
    layer0_outputs(515) <= not (a or b);
    layer0_outputs(516) <= not b or a;
    layer0_outputs(517) <= not b;
    layer0_outputs(518) <= not b;
    layer0_outputs(519) <= not a;
    layer0_outputs(520) <= not b or a;
    layer0_outputs(521) <= b;
    layer0_outputs(522) <= a;
    layer0_outputs(523) <= not b or a;
    layer0_outputs(524) <= not a or b;
    layer0_outputs(525) <= not (a xor b);
    layer0_outputs(526) <= a xor b;
    layer0_outputs(527) <= not b or a;
    layer0_outputs(528) <= a and not b;
    layer0_outputs(529) <= b;
    layer0_outputs(530) <= a and not b;
    layer0_outputs(531) <= a xor b;
    layer0_outputs(532) <= not a or b;
    layer0_outputs(533) <= a;
    layer0_outputs(534) <= b;
    layer0_outputs(535) <= not (a and b);
    layer0_outputs(536) <= b and not a;
    layer0_outputs(537) <= a;
    layer0_outputs(538) <= 1'b1;
    layer0_outputs(539) <= a xor b;
    layer0_outputs(540) <= not a;
    layer0_outputs(541) <= a or b;
    layer0_outputs(542) <= not (a or b);
    layer0_outputs(543) <= not a or b;
    layer0_outputs(544) <= a;
    layer0_outputs(545) <= a and not b;
    layer0_outputs(546) <= 1'b1;
    layer0_outputs(547) <= not b;
    layer0_outputs(548) <= b;
    layer0_outputs(549) <= b;
    layer0_outputs(550) <= b;
    layer0_outputs(551) <= not a or b;
    layer0_outputs(552) <= a xor b;
    layer0_outputs(553) <= not a;
    layer0_outputs(554) <= a or b;
    layer0_outputs(555) <= b and not a;
    layer0_outputs(556) <= a xor b;
    layer0_outputs(557) <= a xor b;
    layer0_outputs(558) <= b;
    layer0_outputs(559) <= a or b;
    layer0_outputs(560) <= not a or b;
    layer0_outputs(561) <= not b or a;
    layer0_outputs(562) <= not b or a;
    layer0_outputs(563) <= not (a or b);
    layer0_outputs(564) <= not b;
    layer0_outputs(565) <= a xor b;
    layer0_outputs(566) <= not (a or b);
    layer0_outputs(567) <= not b;
    layer0_outputs(568) <= not b;
    layer0_outputs(569) <= a or b;
    layer0_outputs(570) <= not (a xor b);
    layer0_outputs(571) <= not (a or b);
    layer0_outputs(572) <= not (a or b);
    layer0_outputs(573) <= not a;
    layer0_outputs(574) <= not (a xor b);
    layer0_outputs(575) <= a and not b;
    layer0_outputs(576) <= 1'b1;
    layer0_outputs(577) <= not (a xor b);
    layer0_outputs(578) <= b;
    layer0_outputs(579) <= a and not b;
    layer0_outputs(580) <= a and not b;
    layer0_outputs(581) <= not a;
    layer0_outputs(582) <= a or b;
    layer0_outputs(583) <= not b;
    layer0_outputs(584) <= not (a or b);
    layer0_outputs(585) <= b;
    layer0_outputs(586) <= a;
    layer0_outputs(587) <= not b;
    layer0_outputs(588) <= not (a or b);
    layer0_outputs(589) <= b;
    layer0_outputs(590) <= a;
    layer0_outputs(591) <= a or b;
    layer0_outputs(592) <= not b or a;
    layer0_outputs(593) <= b;
    layer0_outputs(594) <= not (a or b);
    layer0_outputs(595) <= not b or a;
    layer0_outputs(596) <= not a;
    layer0_outputs(597) <= not a;
    layer0_outputs(598) <= a xor b;
    layer0_outputs(599) <= not (a xor b);
    layer0_outputs(600) <= not b or a;
    layer0_outputs(601) <= a;
    layer0_outputs(602) <= not (a and b);
    layer0_outputs(603) <= not b;
    layer0_outputs(604) <= not b or a;
    layer0_outputs(605) <= not (a or b);
    layer0_outputs(606) <= a xor b;
    layer0_outputs(607) <= not (a or b);
    layer0_outputs(608) <= a xor b;
    layer0_outputs(609) <= a;
    layer0_outputs(610) <= a;
    layer0_outputs(611) <= not a;
    layer0_outputs(612) <= a or b;
    layer0_outputs(613) <= not (a or b);
    layer0_outputs(614) <= not (a or b);
    layer0_outputs(615) <= a and not b;
    layer0_outputs(616) <= not b or a;
    layer0_outputs(617) <= a or b;
    layer0_outputs(618) <= a;
    layer0_outputs(619) <= a and b;
    layer0_outputs(620) <= not (a and b);
    layer0_outputs(621) <= not a or b;
    layer0_outputs(622) <= a and not b;
    layer0_outputs(623) <= 1'b0;
    layer0_outputs(624) <= not a or b;
    layer0_outputs(625) <= b;
    layer0_outputs(626) <= a;
    layer0_outputs(627) <= not b;
    layer0_outputs(628) <= b;
    layer0_outputs(629) <= not (a or b);
    layer0_outputs(630) <= not (a and b);
    layer0_outputs(631) <= not b;
    layer0_outputs(632) <= b;
    layer0_outputs(633) <= b;
    layer0_outputs(634) <= a xor b;
    layer0_outputs(635) <= a xor b;
    layer0_outputs(636) <= a and not b;
    layer0_outputs(637) <= a xor b;
    layer0_outputs(638) <= a and b;
    layer0_outputs(639) <= not a or b;
    layer0_outputs(640) <= a or b;
    layer0_outputs(641) <= a xor b;
    layer0_outputs(642) <= 1'b1;
    layer0_outputs(643) <= a or b;
    layer0_outputs(644) <= a or b;
    layer0_outputs(645) <= a;
    layer0_outputs(646) <= not b;
    layer0_outputs(647) <= not (a or b);
    layer0_outputs(648) <= a;
    layer0_outputs(649) <= not (a xor b);
    layer0_outputs(650) <= 1'b1;
    layer0_outputs(651) <= 1'b1;
    layer0_outputs(652) <= not b;
    layer0_outputs(653) <= a;
    layer0_outputs(654) <= a;
    layer0_outputs(655) <= a;
    layer0_outputs(656) <= not a or b;
    layer0_outputs(657) <= a or b;
    layer0_outputs(658) <= not (a xor b);
    layer0_outputs(659) <= not a or b;
    layer0_outputs(660) <= not a or b;
    layer0_outputs(661) <= b and not a;
    layer0_outputs(662) <= not b or a;
    layer0_outputs(663) <= not a or b;
    layer0_outputs(664) <= a or b;
    layer0_outputs(665) <= a;
    layer0_outputs(666) <= not (a or b);
    layer0_outputs(667) <= not (a and b);
    layer0_outputs(668) <= a or b;
    layer0_outputs(669) <= 1'b0;
    layer0_outputs(670) <= a xor b;
    layer0_outputs(671) <= a;
    layer0_outputs(672) <= a xor b;
    layer0_outputs(673) <= 1'b1;
    layer0_outputs(674) <= not a or b;
    layer0_outputs(675) <= not a or b;
    layer0_outputs(676) <= not a or b;
    layer0_outputs(677) <= a xor b;
    layer0_outputs(678) <= b and not a;
    layer0_outputs(679) <= a or b;
    layer0_outputs(680) <= not b;
    layer0_outputs(681) <= a and b;
    layer0_outputs(682) <= 1'b1;
    layer0_outputs(683) <= not (a xor b);
    layer0_outputs(684) <= not a or b;
    layer0_outputs(685) <= a or b;
    layer0_outputs(686) <= a xor b;
    layer0_outputs(687) <= a xor b;
    layer0_outputs(688) <= not (a and b);
    layer0_outputs(689) <= not (a or b);
    layer0_outputs(690) <= not b or a;
    layer0_outputs(691) <= not a or b;
    layer0_outputs(692) <= not b or a;
    layer0_outputs(693) <= not (a or b);
    layer0_outputs(694) <= a or b;
    layer0_outputs(695) <= not b or a;
    layer0_outputs(696) <= b;
    layer0_outputs(697) <= b;
    layer0_outputs(698) <= a or b;
    layer0_outputs(699) <= a or b;
    layer0_outputs(700) <= a and b;
    layer0_outputs(701) <= 1'b0;
    layer0_outputs(702) <= a xor b;
    layer0_outputs(703) <= not a;
    layer0_outputs(704) <= not (a and b);
    layer0_outputs(705) <= not (a or b);
    layer0_outputs(706) <= not a;
    layer0_outputs(707) <= not a;
    layer0_outputs(708) <= a or b;
    layer0_outputs(709) <= a xor b;
    layer0_outputs(710) <= not (a xor b);
    layer0_outputs(711) <= b and not a;
    layer0_outputs(712) <= not (a or b);
    layer0_outputs(713) <= not a or b;
    layer0_outputs(714) <= not a;
    layer0_outputs(715) <= not a;
    layer0_outputs(716) <= not (a xor b);
    layer0_outputs(717) <= not b or a;
    layer0_outputs(718) <= not (a xor b);
    layer0_outputs(719) <= a or b;
    layer0_outputs(720) <= a;
    layer0_outputs(721) <= not (a or b);
    layer0_outputs(722) <= b and not a;
    layer0_outputs(723) <= not b or a;
    layer0_outputs(724) <= not a or b;
    layer0_outputs(725) <= a and not b;
    layer0_outputs(726) <= not a or b;
    layer0_outputs(727) <= 1'b0;
    layer0_outputs(728) <= a xor b;
    layer0_outputs(729) <= a and b;
    layer0_outputs(730) <= not a;
    layer0_outputs(731) <= 1'b0;
    layer0_outputs(732) <= not a;
    layer0_outputs(733) <= a or b;
    layer0_outputs(734) <= b and not a;
    layer0_outputs(735) <= b and not a;
    layer0_outputs(736) <= not b;
    layer0_outputs(737) <= not a;
    layer0_outputs(738) <= not (a xor b);
    layer0_outputs(739) <= not a or b;
    layer0_outputs(740) <= not (a xor b);
    layer0_outputs(741) <= b and not a;
    layer0_outputs(742) <= not (a and b);
    layer0_outputs(743) <= not b or a;
    layer0_outputs(744) <= a or b;
    layer0_outputs(745) <= b;
    layer0_outputs(746) <= a and not b;
    layer0_outputs(747) <= a or b;
    layer0_outputs(748) <= not (a or b);
    layer0_outputs(749) <= a;
    layer0_outputs(750) <= not (a and b);
    layer0_outputs(751) <= not a;
    layer0_outputs(752) <= a;
    layer0_outputs(753) <= not (a xor b);
    layer0_outputs(754) <= not b or a;
    layer0_outputs(755) <= not a or b;
    layer0_outputs(756) <= b;
    layer0_outputs(757) <= not a or b;
    layer0_outputs(758) <= a and not b;
    layer0_outputs(759) <= a xor b;
    layer0_outputs(760) <= a or b;
    layer0_outputs(761) <= a or b;
    layer0_outputs(762) <= a xor b;
    layer0_outputs(763) <= a and not b;
    layer0_outputs(764) <= not (a or b);
    layer0_outputs(765) <= not b or a;
    layer0_outputs(766) <= a or b;
    layer0_outputs(767) <= a or b;
    layer0_outputs(768) <= not b or a;
    layer0_outputs(769) <= 1'b1;
    layer0_outputs(770) <= b and not a;
    layer0_outputs(771) <= b;
    layer0_outputs(772) <= b;
    layer0_outputs(773) <= a;
    layer0_outputs(774) <= a;
    layer0_outputs(775) <= not b or a;
    layer0_outputs(776) <= not (a or b);
    layer0_outputs(777) <= not (a or b);
    layer0_outputs(778) <= not a or b;
    layer0_outputs(779) <= b;
    layer0_outputs(780) <= not (a xor b);
    layer0_outputs(781) <= a;
    layer0_outputs(782) <= not (a or b);
    layer0_outputs(783) <= not a;
    layer0_outputs(784) <= not a;
    layer0_outputs(785) <= 1'b1;
    layer0_outputs(786) <= not b or a;
    layer0_outputs(787) <= a and b;
    layer0_outputs(788) <= not b;
    layer0_outputs(789) <= not (a and b);
    layer0_outputs(790) <= a and not b;
    layer0_outputs(791) <= not (a or b);
    layer0_outputs(792) <= not a;
    layer0_outputs(793) <= a and b;
    layer0_outputs(794) <= not b or a;
    layer0_outputs(795) <= not a or b;
    layer0_outputs(796) <= a xor b;
    layer0_outputs(797) <= 1'b1;
    layer0_outputs(798) <= a or b;
    layer0_outputs(799) <= not (a or b);
    layer0_outputs(800) <= a or b;
    layer0_outputs(801) <= b;
    layer0_outputs(802) <= not b or a;
    layer0_outputs(803) <= a xor b;
    layer0_outputs(804) <= a or b;
    layer0_outputs(805) <= not (a xor b);
    layer0_outputs(806) <= 1'b1;
    layer0_outputs(807) <= not (a or b);
    layer0_outputs(808) <= not a;
    layer0_outputs(809) <= a or b;
    layer0_outputs(810) <= a xor b;
    layer0_outputs(811) <= b and not a;
    layer0_outputs(812) <= not a;
    layer0_outputs(813) <= not b or a;
    layer0_outputs(814) <= 1'b0;
    layer0_outputs(815) <= not b or a;
    layer0_outputs(816) <= not b;
    layer0_outputs(817) <= b;
    layer0_outputs(818) <= 1'b0;
    layer0_outputs(819) <= 1'b0;
    layer0_outputs(820) <= a or b;
    layer0_outputs(821) <= not a or b;
    layer0_outputs(822) <= b;
    layer0_outputs(823) <= not b or a;
    layer0_outputs(824) <= a or b;
    layer0_outputs(825) <= not (a and b);
    layer0_outputs(826) <= not (a xor b);
    layer0_outputs(827) <= not (a or b);
    layer0_outputs(828) <= not b or a;
    layer0_outputs(829) <= 1'b1;
    layer0_outputs(830) <= b;
    layer0_outputs(831) <= a and not b;
    layer0_outputs(832) <= b;
    layer0_outputs(833) <= not b;
    layer0_outputs(834) <= b;
    layer0_outputs(835) <= b;
    layer0_outputs(836) <= a and not b;
    layer0_outputs(837) <= not b or a;
    layer0_outputs(838) <= a xor b;
    layer0_outputs(839) <= not (a or b);
    layer0_outputs(840) <= a;
    layer0_outputs(841) <= b;
    layer0_outputs(842) <= a and not b;
    layer0_outputs(843) <= a or b;
    layer0_outputs(844) <= a;
    layer0_outputs(845) <= a xor b;
    layer0_outputs(846) <= b and not a;
    layer0_outputs(847) <= not a;
    layer0_outputs(848) <= a and not b;
    layer0_outputs(849) <= a and not b;
    layer0_outputs(850) <= not (a or b);
    layer0_outputs(851) <= not b;
    layer0_outputs(852) <= a and b;
    layer0_outputs(853) <= not b;
    layer0_outputs(854) <= not a or b;
    layer0_outputs(855) <= 1'b0;
    layer0_outputs(856) <= not (a xor b);
    layer0_outputs(857) <= not (a and b);
    layer0_outputs(858) <= not (a or b);
    layer0_outputs(859) <= a and not b;
    layer0_outputs(860) <= 1'b0;
    layer0_outputs(861) <= a or b;
    layer0_outputs(862) <= not b;
    layer0_outputs(863) <= a or b;
    layer0_outputs(864) <= not (a xor b);
    layer0_outputs(865) <= not a;
    layer0_outputs(866) <= not a or b;
    layer0_outputs(867) <= a xor b;
    layer0_outputs(868) <= a xor b;
    layer0_outputs(869) <= 1'b0;
    layer0_outputs(870) <= not (a or b);
    layer0_outputs(871) <= not (a or b);
    layer0_outputs(872) <= 1'b1;
    layer0_outputs(873) <= a and not b;
    layer0_outputs(874) <= a or b;
    layer0_outputs(875) <= not (a and b);
    layer0_outputs(876) <= not a or b;
    layer0_outputs(877) <= not a;
    layer0_outputs(878) <= a and not b;
    layer0_outputs(879) <= a;
    layer0_outputs(880) <= a;
    layer0_outputs(881) <= not b or a;
    layer0_outputs(882) <= b;
    layer0_outputs(883) <= a;
    layer0_outputs(884) <= a and b;
    layer0_outputs(885) <= a and not b;
    layer0_outputs(886) <= a and b;
    layer0_outputs(887) <= not (a xor b);
    layer0_outputs(888) <= not b or a;
    layer0_outputs(889) <= b and not a;
    layer0_outputs(890) <= a xor b;
    layer0_outputs(891) <= b;
    layer0_outputs(892) <= not (a or b);
    layer0_outputs(893) <= a and not b;
    layer0_outputs(894) <= not a or b;
    layer0_outputs(895) <= not (a xor b);
    layer0_outputs(896) <= not a;
    layer0_outputs(897) <= not a;
    layer0_outputs(898) <= b;
    layer0_outputs(899) <= a or b;
    layer0_outputs(900) <= a and not b;
    layer0_outputs(901) <= not a;
    layer0_outputs(902) <= not a or b;
    layer0_outputs(903) <= not a or b;
    layer0_outputs(904) <= not a or b;
    layer0_outputs(905) <= not (a or b);
    layer0_outputs(906) <= not b or a;
    layer0_outputs(907) <= a and b;
    layer0_outputs(908) <= not b or a;
    layer0_outputs(909) <= a or b;
    layer0_outputs(910) <= not b;
    layer0_outputs(911) <= not a or b;
    layer0_outputs(912) <= a;
    layer0_outputs(913) <= a;
    layer0_outputs(914) <= a xor b;
    layer0_outputs(915) <= not b;
    layer0_outputs(916) <= b;
    layer0_outputs(917) <= a;
    layer0_outputs(918) <= b;
    layer0_outputs(919) <= a and not b;
    layer0_outputs(920) <= b and not a;
    layer0_outputs(921) <= a;
    layer0_outputs(922) <= not (a xor b);
    layer0_outputs(923) <= not b or a;
    layer0_outputs(924) <= 1'b0;
    layer0_outputs(925) <= b;
    layer0_outputs(926) <= a;
    layer0_outputs(927) <= not a;
    layer0_outputs(928) <= a or b;
    layer0_outputs(929) <= not a;
    layer0_outputs(930) <= not (a and b);
    layer0_outputs(931) <= not (a xor b);
    layer0_outputs(932) <= a;
    layer0_outputs(933) <= a xor b;
    layer0_outputs(934) <= not (a or b);
    layer0_outputs(935) <= not a or b;
    layer0_outputs(936) <= not b;
    layer0_outputs(937) <= not a;
    layer0_outputs(938) <= not (a xor b);
    layer0_outputs(939) <= not b;
    layer0_outputs(940) <= not (a and b);
    layer0_outputs(941) <= b and not a;
    layer0_outputs(942) <= not (a or b);
    layer0_outputs(943) <= not a;
    layer0_outputs(944) <= not (a xor b);
    layer0_outputs(945) <= a xor b;
    layer0_outputs(946) <= not (a xor b);
    layer0_outputs(947) <= a or b;
    layer0_outputs(948) <= b;
    layer0_outputs(949) <= not (a or b);
    layer0_outputs(950) <= not (a or b);
    layer0_outputs(951) <= not a;
    layer0_outputs(952) <= a or b;
    layer0_outputs(953) <= a and not b;
    layer0_outputs(954) <= not a;
    layer0_outputs(955) <= b;
    layer0_outputs(956) <= a or b;
    layer0_outputs(957) <= 1'b1;
    layer0_outputs(958) <= a xor b;
    layer0_outputs(959) <= 1'b0;
    layer0_outputs(960) <= not (a xor b);
    layer0_outputs(961) <= not (a xor b);
    layer0_outputs(962) <= not (a xor b);
    layer0_outputs(963) <= a or b;
    layer0_outputs(964) <= not (a xor b);
    layer0_outputs(965) <= a and b;
    layer0_outputs(966) <= a xor b;
    layer0_outputs(967) <= b and not a;
    layer0_outputs(968) <= a xor b;
    layer0_outputs(969) <= a and not b;
    layer0_outputs(970) <= not (a xor b);
    layer0_outputs(971) <= a xor b;
    layer0_outputs(972) <= not (a or b);
    layer0_outputs(973) <= not b;
    layer0_outputs(974) <= a;
    layer0_outputs(975) <= a;
    layer0_outputs(976) <= not b or a;
    layer0_outputs(977) <= b and not a;
    layer0_outputs(978) <= not b;
    layer0_outputs(979) <= not a or b;
    layer0_outputs(980) <= b and not a;
    layer0_outputs(981) <= a or b;
    layer0_outputs(982) <= not b or a;
    layer0_outputs(983) <= not a or b;
    layer0_outputs(984) <= 1'b0;
    layer0_outputs(985) <= b and not a;
    layer0_outputs(986) <= a;
    layer0_outputs(987) <= a or b;
    layer0_outputs(988) <= a xor b;
    layer0_outputs(989) <= a xor b;
    layer0_outputs(990) <= a;
    layer0_outputs(991) <= not b or a;
    layer0_outputs(992) <= not (a or b);
    layer0_outputs(993) <= 1'b0;
    layer0_outputs(994) <= a;
    layer0_outputs(995) <= a and b;
    layer0_outputs(996) <= a or b;
    layer0_outputs(997) <= a;
    layer0_outputs(998) <= not (a and b);
    layer0_outputs(999) <= a;
    layer0_outputs(1000) <= 1'b1;
    layer0_outputs(1001) <= a or b;
    layer0_outputs(1002) <= b;
    layer0_outputs(1003) <= not a or b;
    layer0_outputs(1004) <= not b;
    layer0_outputs(1005) <= not (a xor b);
    layer0_outputs(1006) <= not (a xor b);
    layer0_outputs(1007) <= a;
    layer0_outputs(1008) <= b and not a;
    layer0_outputs(1009) <= a and not b;
    layer0_outputs(1010) <= not b or a;
    layer0_outputs(1011) <= not (a xor b);
    layer0_outputs(1012) <= a or b;
    layer0_outputs(1013) <= a;
    layer0_outputs(1014) <= not b or a;
    layer0_outputs(1015) <= not (a and b);
    layer0_outputs(1016) <= not a or b;
    layer0_outputs(1017) <= b and not a;
    layer0_outputs(1018) <= not b;
    layer0_outputs(1019) <= a;
    layer0_outputs(1020) <= a xor b;
    layer0_outputs(1021) <= not b;
    layer0_outputs(1022) <= not a;
    layer0_outputs(1023) <= not b or a;
    layer0_outputs(1024) <= a xor b;
    layer0_outputs(1025) <= a xor b;
    layer0_outputs(1026) <= a;
    layer0_outputs(1027) <= a;
    layer0_outputs(1028) <= a xor b;
    layer0_outputs(1029) <= b and not a;
    layer0_outputs(1030) <= b and not a;
    layer0_outputs(1031) <= not a;
    layer0_outputs(1032) <= a;
    layer0_outputs(1033) <= a;
    layer0_outputs(1034) <= not (a or b);
    layer0_outputs(1035) <= a or b;
    layer0_outputs(1036) <= not (a xor b);
    layer0_outputs(1037) <= a or b;
    layer0_outputs(1038) <= a xor b;
    layer0_outputs(1039) <= b and not a;
    layer0_outputs(1040) <= b and not a;
    layer0_outputs(1041) <= not b;
    layer0_outputs(1042) <= a and b;
    layer0_outputs(1043) <= not (a or b);
    layer0_outputs(1044) <= b and not a;
    layer0_outputs(1045) <= not (a or b);
    layer0_outputs(1046) <= not (a or b);
    layer0_outputs(1047) <= not a;
    layer0_outputs(1048) <= not a;
    layer0_outputs(1049) <= a and not b;
    layer0_outputs(1050) <= b and not a;
    layer0_outputs(1051) <= not (a or b);
    layer0_outputs(1052) <= b and not a;
    layer0_outputs(1053) <= a;
    layer0_outputs(1054) <= not a or b;
    layer0_outputs(1055) <= b;
    layer0_outputs(1056) <= a or b;
    layer0_outputs(1057) <= not (a and b);
    layer0_outputs(1058) <= a or b;
    layer0_outputs(1059) <= not (a or b);
    layer0_outputs(1060) <= a;
    layer0_outputs(1061) <= a or b;
    layer0_outputs(1062) <= not a or b;
    layer0_outputs(1063) <= a and not b;
    layer0_outputs(1064) <= not b or a;
    layer0_outputs(1065) <= not a;
    layer0_outputs(1066) <= a or b;
    layer0_outputs(1067) <= not a or b;
    layer0_outputs(1068) <= not b;
    layer0_outputs(1069) <= not b or a;
    layer0_outputs(1070) <= not b or a;
    layer0_outputs(1071) <= not (a xor b);
    layer0_outputs(1072) <= a xor b;
    layer0_outputs(1073) <= 1'b1;
    layer0_outputs(1074) <= not a or b;
    layer0_outputs(1075) <= a and b;
    layer0_outputs(1076) <= not a;
    layer0_outputs(1077) <= a or b;
    layer0_outputs(1078) <= not (a or b);
    layer0_outputs(1079) <= not (a or b);
    layer0_outputs(1080) <= 1'b0;
    layer0_outputs(1081) <= a and not b;
    layer0_outputs(1082) <= not b;
    layer0_outputs(1083) <= not (a or b);
    layer0_outputs(1084) <= not b or a;
    layer0_outputs(1085) <= not b;
    layer0_outputs(1086) <= a or b;
    layer0_outputs(1087) <= b;
    layer0_outputs(1088) <= b;
    layer0_outputs(1089) <= b;
    layer0_outputs(1090) <= a xor b;
    layer0_outputs(1091) <= 1'b0;
    layer0_outputs(1092) <= a;
    layer0_outputs(1093) <= b;
    layer0_outputs(1094) <= a and b;
    layer0_outputs(1095) <= b and not a;
    layer0_outputs(1096) <= not a;
    layer0_outputs(1097) <= not a or b;
    layer0_outputs(1098) <= not (a or b);
    layer0_outputs(1099) <= not (a or b);
    layer0_outputs(1100) <= not a;
    layer0_outputs(1101) <= 1'b0;
    layer0_outputs(1102) <= not (a and b);
    layer0_outputs(1103) <= not b;
    layer0_outputs(1104) <= not (a or b);
    layer0_outputs(1105) <= not b;
    layer0_outputs(1106) <= a xor b;
    layer0_outputs(1107) <= not a;
    layer0_outputs(1108) <= a;
    layer0_outputs(1109) <= not (a xor b);
    layer0_outputs(1110) <= 1'b0;
    layer0_outputs(1111) <= not (a or b);
    layer0_outputs(1112) <= not a;
    layer0_outputs(1113) <= not (a xor b);
    layer0_outputs(1114) <= not b;
    layer0_outputs(1115) <= not b;
    layer0_outputs(1116) <= a or b;
    layer0_outputs(1117) <= not b;
    layer0_outputs(1118) <= a or b;
    layer0_outputs(1119) <= not a or b;
    layer0_outputs(1120) <= not (a xor b);
    layer0_outputs(1121) <= a or b;
    layer0_outputs(1122) <= a;
    layer0_outputs(1123) <= not b or a;
    layer0_outputs(1124) <= a or b;
    layer0_outputs(1125) <= not a;
    layer0_outputs(1126) <= not (a and b);
    layer0_outputs(1127) <= a;
    layer0_outputs(1128) <= a or b;
    layer0_outputs(1129) <= not (a and b);
    layer0_outputs(1130) <= b;
    layer0_outputs(1131) <= a xor b;
    layer0_outputs(1132) <= b;
    layer0_outputs(1133) <= not b or a;
    layer0_outputs(1134) <= not (a xor b);
    layer0_outputs(1135) <= not (a or b);
    layer0_outputs(1136) <= not (a or b);
    layer0_outputs(1137) <= not b;
    layer0_outputs(1138) <= a xor b;
    layer0_outputs(1139) <= a xor b;
    layer0_outputs(1140) <= a and not b;
    layer0_outputs(1141) <= 1'b0;
    layer0_outputs(1142) <= 1'b1;
    layer0_outputs(1143) <= not b or a;
    layer0_outputs(1144) <= 1'b1;
    layer0_outputs(1145) <= not b;
    layer0_outputs(1146) <= not (a xor b);
    layer0_outputs(1147) <= not a or b;
    layer0_outputs(1148) <= a and b;
    layer0_outputs(1149) <= 1'b1;
    layer0_outputs(1150) <= a and not b;
    layer0_outputs(1151) <= not (a or b);
    layer0_outputs(1152) <= a or b;
    layer0_outputs(1153) <= a and not b;
    layer0_outputs(1154) <= a and not b;
    layer0_outputs(1155) <= not b;
    layer0_outputs(1156) <= not a or b;
    layer0_outputs(1157) <= b and not a;
    layer0_outputs(1158) <= b;
    layer0_outputs(1159) <= a;
    layer0_outputs(1160) <= b;
    layer0_outputs(1161) <= b and not a;
    layer0_outputs(1162) <= not b;
    layer0_outputs(1163) <= a xor b;
    layer0_outputs(1164) <= not a;
    layer0_outputs(1165) <= not a or b;
    layer0_outputs(1166) <= a;
    layer0_outputs(1167) <= not a or b;
    layer0_outputs(1168) <= b;
    layer0_outputs(1169) <= not (a and b);
    layer0_outputs(1170) <= not (a or b);
    layer0_outputs(1171) <= 1'b0;
    layer0_outputs(1172) <= a or b;
    layer0_outputs(1173) <= not (a xor b);
    layer0_outputs(1174) <= a or b;
    layer0_outputs(1175) <= a xor b;
    layer0_outputs(1176) <= b;
    layer0_outputs(1177) <= not (a xor b);
    layer0_outputs(1178) <= not b or a;
    layer0_outputs(1179) <= a and b;
    layer0_outputs(1180) <= not (a or b);
    layer0_outputs(1181) <= not b or a;
    layer0_outputs(1182) <= not a or b;
    layer0_outputs(1183) <= not b;
    layer0_outputs(1184) <= not a or b;
    layer0_outputs(1185) <= b;
    layer0_outputs(1186) <= a or b;
    layer0_outputs(1187) <= b;
    layer0_outputs(1188) <= not a;
    layer0_outputs(1189) <= a or b;
    layer0_outputs(1190) <= a and not b;
    layer0_outputs(1191) <= b;
    layer0_outputs(1192) <= not (a or b);
    layer0_outputs(1193) <= not b or a;
    layer0_outputs(1194) <= a and b;
    layer0_outputs(1195) <= a xor b;
    layer0_outputs(1196) <= b;
    layer0_outputs(1197) <= a xor b;
    layer0_outputs(1198) <= b;
    layer0_outputs(1199) <= not b;
    layer0_outputs(1200) <= a or b;
    layer0_outputs(1201) <= not b;
    layer0_outputs(1202) <= not b;
    layer0_outputs(1203) <= not a;
    layer0_outputs(1204) <= b;
    layer0_outputs(1205) <= not a;
    layer0_outputs(1206) <= b;
    layer0_outputs(1207) <= not (a and b);
    layer0_outputs(1208) <= a and not b;
    layer0_outputs(1209) <= not (a and b);
    layer0_outputs(1210) <= a;
    layer0_outputs(1211) <= not (a and b);
    layer0_outputs(1212) <= a;
    layer0_outputs(1213) <= b and not a;
    layer0_outputs(1214) <= a and not b;
    layer0_outputs(1215) <= a xor b;
    layer0_outputs(1216) <= 1'b0;
    layer0_outputs(1217) <= not b;
    layer0_outputs(1218) <= not a;
    layer0_outputs(1219) <= not b or a;
    layer0_outputs(1220) <= not b;
    layer0_outputs(1221) <= a or b;
    layer0_outputs(1222) <= not (a xor b);
    layer0_outputs(1223) <= a and b;
    layer0_outputs(1224) <= b and not a;
    layer0_outputs(1225) <= not a or b;
    layer0_outputs(1226) <= 1'b1;
    layer0_outputs(1227) <= b;
    layer0_outputs(1228) <= b;
    layer0_outputs(1229) <= not b or a;
    layer0_outputs(1230) <= 1'b0;
    layer0_outputs(1231) <= not a;
    layer0_outputs(1232) <= a or b;
    layer0_outputs(1233) <= a and b;
    layer0_outputs(1234) <= 1'b0;
    layer0_outputs(1235) <= not (a xor b);
    layer0_outputs(1236) <= b and not a;
    layer0_outputs(1237) <= not (a or b);
    layer0_outputs(1238) <= not (a and b);
    layer0_outputs(1239) <= not (a or b);
    layer0_outputs(1240) <= a and not b;
    layer0_outputs(1241) <= a or b;
    layer0_outputs(1242) <= a;
    layer0_outputs(1243) <= not (a or b);
    layer0_outputs(1244) <= not b;
    layer0_outputs(1245) <= a xor b;
    layer0_outputs(1246) <= a and not b;
    layer0_outputs(1247) <= not a;
    layer0_outputs(1248) <= b;
    layer0_outputs(1249) <= not (a or b);
    layer0_outputs(1250) <= not b or a;
    layer0_outputs(1251) <= a and not b;
    layer0_outputs(1252) <= a xor b;
    layer0_outputs(1253) <= not (a xor b);
    layer0_outputs(1254) <= a and not b;
    layer0_outputs(1255) <= a;
    layer0_outputs(1256) <= a;
    layer0_outputs(1257) <= not b;
    layer0_outputs(1258) <= not (a or b);
    layer0_outputs(1259) <= b;
    layer0_outputs(1260) <= 1'b0;
    layer0_outputs(1261) <= not a or b;
    layer0_outputs(1262) <= a xor b;
    layer0_outputs(1263) <= not (a and b);
    layer0_outputs(1264) <= not (a or b);
    layer0_outputs(1265) <= not (a or b);
    layer0_outputs(1266) <= 1'b0;
    layer0_outputs(1267) <= b;
    layer0_outputs(1268) <= not a;
    layer0_outputs(1269) <= not (a xor b);
    layer0_outputs(1270) <= b and not a;
    layer0_outputs(1271) <= a xor b;
    layer0_outputs(1272) <= b;
    layer0_outputs(1273) <= not a;
    layer0_outputs(1274) <= not (a or b);
    layer0_outputs(1275) <= a and not b;
    layer0_outputs(1276) <= not (a xor b);
    layer0_outputs(1277) <= 1'b0;
    layer0_outputs(1278) <= b and not a;
    layer0_outputs(1279) <= b;
    layer0_outputs(1280) <= a and not b;
    layer0_outputs(1281) <= a and not b;
    layer0_outputs(1282) <= not a;
    layer0_outputs(1283) <= not a;
    layer0_outputs(1284) <= a and b;
    layer0_outputs(1285) <= b;
    layer0_outputs(1286) <= not a or b;
    layer0_outputs(1287) <= not (a and b);
    layer0_outputs(1288) <= not (a or b);
    layer0_outputs(1289) <= not b or a;
    layer0_outputs(1290) <= not b;
    layer0_outputs(1291) <= a xor b;
    layer0_outputs(1292) <= 1'b1;
    layer0_outputs(1293) <= not b;
    layer0_outputs(1294) <= a;
    layer0_outputs(1295) <= a;
    layer0_outputs(1296) <= not a;
    layer0_outputs(1297) <= a xor b;
    layer0_outputs(1298) <= not b or a;
    layer0_outputs(1299) <= not b;
    layer0_outputs(1300) <= a xor b;
    layer0_outputs(1301) <= a and not b;
    layer0_outputs(1302) <= a or b;
    layer0_outputs(1303) <= a xor b;
    layer0_outputs(1304) <= a and not b;
    layer0_outputs(1305) <= not (a xor b);
    layer0_outputs(1306) <= a;
    layer0_outputs(1307) <= a or b;
    layer0_outputs(1308) <= a xor b;
    layer0_outputs(1309) <= b and not a;
    layer0_outputs(1310) <= not b;
    layer0_outputs(1311) <= a and not b;
    layer0_outputs(1312) <= a or b;
    layer0_outputs(1313) <= a or b;
    layer0_outputs(1314) <= not (a or b);
    layer0_outputs(1315) <= a and not b;
    layer0_outputs(1316) <= not (a or b);
    layer0_outputs(1317) <= a or b;
    layer0_outputs(1318) <= a and not b;
    layer0_outputs(1319) <= not (a or b);
    layer0_outputs(1320) <= not b or a;
    layer0_outputs(1321) <= not (a or b);
    layer0_outputs(1322) <= a or b;
    layer0_outputs(1323) <= not b or a;
    layer0_outputs(1324) <= a or b;
    layer0_outputs(1325) <= 1'b1;
    layer0_outputs(1326) <= not (a or b);
    layer0_outputs(1327) <= not (a xor b);
    layer0_outputs(1328) <= a and b;
    layer0_outputs(1329) <= not a or b;
    layer0_outputs(1330) <= not a or b;
    layer0_outputs(1331) <= b;
    layer0_outputs(1332) <= not (a or b);
    layer0_outputs(1333) <= not a;
    layer0_outputs(1334) <= not (a or b);
    layer0_outputs(1335) <= a;
    layer0_outputs(1336) <= 1'b0;
    layer0_outputs(1337) <= 1'b1;
    layer0_outputs(1338) <= not (a xor b);
    layer0_outputs(1339) <= b;
    layer0_outputs(1340) <= b;
    layer0_outputs(1341) <= b;
    layer0_outputs(1342) <= a and not b;
    layer0_outputs(1343) <= not (a xor b);
    layer0_outputs(1344) <= 1'b1;
    layer0_outputs(1345) <= a xor b;
    layer0_outputs(1346) <= not (a xor b);
    layer0_outputs(1347) <= b and not a;
    layer0_outputs(1348) <= 1'b1;
    layer0_outputs(1349) <= a and not b;
    layer0_outputs(1350) <= not (a or b);
    layer0_outputs(1351) <= a or b;
    layer0_outputs(1352) <= 1'b0;
    layer0_outputs(1353) <= not a;
    layer0_outputs(1354) <= not (a xor b);
    layer0_outputs(1355) <= not b;
    layer0_outputs(1356) <= a;
    layer0_outputs(1357) <= a and not b;
    layer0_outputs(1358) <= not (a or b);
    layer0_outputs(1359) <= 1'b0;
    layer0_outputs(1360) <= a or b;
    layer0_outputs(1361) <= not (a or b);
    layer0_outputs(1362) <= a and b;
    layer0_outputs(1363) <= a;
    layer0_outputs(1364) <= b and not a;
    layer0_outputs(1365) <= a xor b;
    layer0_outputs(1366) <= a and b;
    layer0_outputs(1367) <= a and not b;
    layer0_outputs(1368) <= not a or b;
    layer0_outputs(1369) <= not (a or b);
    layer0_outputs(1370) <= b;
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= b and not a;
    layer0_outputs(1373) <= a and b;
    layer0_outputs(1374) <= b and not a;
    layer0_outputs(1375) <= not (a xor b);
    layer0_outputs(1376) <= 1'b0;
    layer0_outputs(1377) <= a xor b;
    layer0_outputs(1378) <= not (a or b);
    layer0_outputs(1379) <= b;
    layer0_outputs(1380) <= b and not a;
    layer0_outputs(1381) <= not b;
    layer0_outputs(1382) <= a;
    layer0_outputs(1383) <= b and not a;
    layer0_outputs(1384) <= a;
    layer0_outputs(1385) <= a or b;
    layer0_outputs(1386) <= not (a or b);
    layer0_outputs(1387) <= a and not b;
    layer0_outputs(1388) <= 1'b0;
    layer0_outputs(1389) <= a and b;
    layer0_outputs(1390) <= not (a xor b);
    layer0_outputs(1391) <= a xor b;
    layer0_outputs(1392) <= a or b;
    layer0_outputs(1393) <= not (a xor b);
    layer0_outputs(1394) <= a and not b;
    layer0_outputs(1395) <= a or b;
    layer0_outputs(1396) <= b and not a;
    layer0_outputs(1397) <= a;
    layer0_outputs(1398) <= a xor b;
    layer0_outputs(1399) <= a;
    layer0_outputs(1400) <= not (a or b);
    layer0_outputs(1401) <= b and not a;
    layer0_outputs(1402) <= not a or b;
    layer0_outputs(1403) <= not (a and b);
    layer0_outputs(1404) <= b and not a;
    layer0_outputs(1405) <= not (a or b);
    layer0_outputs(1406) <= not a;
    layer0_outputs(1407) <= not a or b;
    layer0_outputs(1408) <= a or b;
    layer0_outputs(1409) <= a or b;
    layer0_outputs(1410) <= not a;
    layer0_outputs(1411) <= not a;
    layer0_outputs(1412) <= not a or b;
    layer0_outputs(1413) <= not a;
    layer0_outputs(1414) <= not (a xor b);
    layer0_outputs(1415) <= a and not b;
    layer0_outputs(1416) <= not a;
    layer0_outputs(1417) <= not a;
    layer0_outputs(1418) <= 1'b1;
    layer0_outputs(1419) <= a xor b;
    layer0_outputs(1420) <= 1'b1;
    layer0_outputs(1421) <= not b;
    layer0_outputs(1422) <= a;
    layer0_outputs(1423) <= not b or a;
    layer0_outputs(1424) <= not a;
    layer0_outputs(1425) <= not (a xor b);
    layer0_outputs(1426) <= not (a or b);
    layer0_outputs(1427) <= a xor b;
    layer0_outputs(1428) <= b and not a;
    layer0_outputs(1429) <= not (a or b);
    layer0_outputs(1430) <= 1'b1;
    layer0_outputs(1431) <= not (a xor b);
    layer0_outputs(1432) <= a and not b;
    layer0_outputs(1433) <= a and not b;
    layer0_outputs(1434) <= a and not b;
    layer0_outputs(1435) <= a and b;
    layer0_outputs(1436) <= b;
    layer0_outputs(1437) <= a and b;
    layer0_outputs(1438) <= 1'b0;
    layer0_outputs(1439) <= not b;
    layer0_outputs(1440) <= not a or b;
    layer0_outputs(1441) <= not a or b;
    layer0_outputs(1442) <= not b;
    layer0_outputs(1443) <= 1'b0;
    layer0_outputs(1444) <= not b;
    layer0_outputs(1445) <= not (a or b);
    layer0_outputs(1446) <= a and b;
    layer0_outputs(1447) <= not (a xor b);
    layer0_outputs(1448) <= a xor b;
    layer0_outputs(1449) <= not (a or b);
    layer0_outputs(1450) <= not a;
    layer0_outputs(1451) <= not b;
    layer0_outputs(1452) <= a or b;
    layer0_outputs(1453) <= not b or a;
    layer0_outputs(1454) <= b;
    layer0_outputs(1455) <= b;
    layer0_outputs(1456) <= a or b;
    layer0_outputs(1457) <= a and not b;
    layer0_outputs(1458) <= not (a xor b);
    layer0_outputs(1459) <= a or b;
    layer0_outputs(1460) <= a and not b;
    layer0_outputs(1461) <= not (a xor b);
    layer0_outputs(1462) <= 1'b0;
    layer0_outputs(1463) <= a and not b;
    layer0_outputs(1464) <= not a or b;
    layer0_outputs(1465) <= b and not a;
    layer0_outputs(1466) <= a or b;
    layer0_outputs(1467) <= a and not b;
    layer0_outputs(1468) <= a xor b;
    layer0_outputs(1469) <= b and not a;
    layer0_outputs(1470) <= not (a or b);
    layer0_outputs(1471) <= b and not a;
    layer0_outputs(1472) <= not (a xor b);
    layer0_outputs(1473) <= not (a or b);
    layer0_outputs(1474) <= not (a and b);
    layer0_outputs(1475) <= 1'b1;
    layer0_outputs(1476) <= a;
    layer0_outputs(1477) <= a;
    layer0_outputs(1478) <= not (a or b);
    layer0_outputs(1479) <= a and not b;
    layer0_outputs(1480) <= not b;
    layer0_outputs(1481) <= not b;
    layer0_outputs(1482) <= a;
    layer0_outputs(1483) <= not a;
    layer0_outputs(1484) <= 1'b0;
    layer0_outputs(1485) <= not (a or b);
    layer0_outputs(1486) <= a or b;
    layer0_outputs(1487) <= not (a or b);
    layer0_outputs(1488) <= a or b;
    layer0_outputs(1489) <= 1'b1;
    layer0_outputs(1490) <= b and not a;
    layer0_outputs(1491) <= a;
    layer0_outputs(1492) <= a or b;
    layer0_outputs(1493) <= a or b;
    layer0_outputs(1494) <= not b or a;
    layer0_outputs(1495) <= 1'b1;
    layer0_outputs(1496) <= a and b;
    layer0_outputs(1497) <= not b;
    layer0_outputs(1498) <= not a;
    layer0_outputs(1499) <= not (a or b);
    layer0_outputs(1500) <= 1'b1;
    layer0_outputs(1501) <= not (a or b);
    layer0_outputs(1502) <= not a;
    layer0_outputs(1503) <= b and not a;
    layer0_outputs(1504) <= a and not b;
    layer0_outputs(1505) <= b and not a;
    layer0_outputs(1506) <= b and not a;
    layer0_outputs(1507) <= 1'b0;
    layer0_outputs(1508) <= a and not b;
    layer0_outputs(1509) <= not a or b;
    layer0_outputs(1510) <= not (a and b);
    layer0_outputs(1511) <= not (a or b);
    layer0_outputs(1512) <= 1'b0;
    layer0_outputs(1513) <= a or b;
    layer0_outputs(1514) <= b;
    layer0_outputs(1515) <= a or b;
    layer0_outputs(1516) <= not b or a;
    layer0_outputs(1517) <= a and b;
    layer0_outputs(1518) <= a or b;
    layer0_outputs(1519) <= not (a and b);
    layer0_outputs(1520) <= a xor b;
    layer0_outputs(1521) <= a xor b;
    layer0_outputs(1522) <= 1'b1;
    layer0_outputs(1523) <= not a;
    layer0_outputs(1524) <= a xor b;
    layer0_outputs(1525) <= not (a xor b);
    layer0_outputs(1526) <= not b or a;
    layer0_outputs(1527) <= not a or b;
    layer0_outputs(1528) <= not (a xor b);
    layer0_outputs(1529) <= not b;
    layer0_outputs(1530) <= not b;
    layer0_outputs(1531) <= not (a or b);
    layer0_outputs(1532) <= not b;
    layer0_outputs(1533) <= a;
    layer0_outputs(1534) <= a;
    layer0_outputs(1535) <= b;
    layer0_outputs(1536) <= not (a xor b);
    layer0_outputs(1537) <= not b;
    layer0_outputs(1538) <= a xor b;
    layer0_outputs(1539) <= b and not a;
    layer0_outputs(1540) <= a or b;
    layer0_outputs(1541) <= not a or b;
    layer0_outputs(1542) <= not b or a;
    layer0_outputs(1543) <= b and not a;
    layer0_outputs(1544) <= not (a or b);
    layer0_outputs(1545) <= not (a xor b);
    layer0_outputs(1546) <= not b;
    layer0_outputs(1547) <= a xor b;
    layer0_outputs(1548) <= a and not b;
    layer0_outputs(1549) <= a or b;
    layer0_outputs(1550) <= not a or b;
    layer0_outputs(1551) <= 1'b0;
    layer0_outputs(1552) <= not (a or b);
    layer0_outputs(1553) <= not a or b;
    layer0_outputs(1554) <= b and not a;
    layer0_outputs(1555) <= a and not b;
    layer0_outputs(1556) <= not a or b;
    layer0_outputs(1557) <= a xor b;
    layer0_outputs(1558) <= a and not b;
    layer0_outputs(1559) <= b;
    layer0_outputs(1560) <= a or b;
    layer0_outputs(1561) <= not (a or b);
    layer0_outputs(1562) <= 1'b0;
    layer0_outputs(1563) <= not (a or b);
    layer0_outputs(1564) <= not a;
    layer0_outputs(1565) <= b;
    layer0_outputs(1566) <= not b or a;
    layer0_outputs(1567) <= a xor b;
    layer0_outputs(1568) <= a;
    layer0_outputs(1569) <= 1'b0;
    layer0_outputs(1570) <= a and b;
    layer0_outputs(1571) <= 1'b1;
    layer0_outputs(1572) <= not (a or b);
    layer0_outputs(1573) <= a or b;
    layer0_outputs(1574) <= not b or a;
    layer0_outputs(1575) <= b and not a;
    layer0_outputs(1576) <= not b;
    layer0_outputs(1577) <= b;
    layer0_outputs(1578) <= not (a or b);
    layer0_outputs(1579) <= not a or b;
    layer0_outputs(1580) <= b;
    layer0_outputs(1581) <= a or b;
    layer0_outputs(1582) <= a;
    layer0_outputs(1583) <= not a;
    layer0_outputs(1584) <= a;
    layer0_outputs(1585) <= a xor b;
    layer0_outputs(1586) <= a;
    layer0_outputs(1587) <= a or b;
    layer0_outputs(1588) <= not a or b;
    layer0_outputs(1589) <= 1'b0;
    layer0_outputs(1590) <= not b;
    layer0_outputs(1591) <= not a;
    layer0_outputs(1592) <= a xor b;
    layer0_outputs(1593) <= a xor b;
    layer0_outputs(1594) <= not (a or b);
    layer0_outputs(1595) <= b and not a;
    layer0_outputs(1596) <= not b or a;
    layer0_outputs(1597) <= not b or a;
    layer0_outputs(1598) <= 1'b1;
    layer0_outputs(1599) <= a xor b;
    layer0_outputs(1600) <= not (a or b);
    layer0_outputs(1601) <= a or b;
    layer0_outputs(1602) <= not (a or b);
    layer0_outputs(1603) <= not (a or b);
    layer0_outputs(1604) <= not (a xor b);
    layer0_outputs(1605) <= a xor b;
    layer0_outputs(1606) <= a xor b;
    layer0_outputs(1607) <= a or b;
    layer0_outputs(1608) <= a and b;
    layer0_outputs(1609) <= a and not b;
    layer0_outputs(1610) <= not b;
    layer0_outputs(1611) <= not b;
    layer0_outputs(1612) <= not (a or b);
    layer0_outputs(1613) <= a;
    layer0_outputs(1614) <= not (a or b);
    layer0_outputs(1615) <= not (a or b);
    layer0_outputs(1616) <= not b;
    layer0_outputs(1617) <= a and b;
    layer0_outputs(1618) <= 1'b1;
    layer0_outputs(1619) <= not a;
    layer0_outputs(1620) <= 1'b1;
    layer0_outputs(1621) <= not b;
    layer0_outputs(1622) <= not a;
    layer0_outputs(1623) <= a xor b;
    layer0_outputs(1624) <= not (a xor b);
    layer0_outputs(1625) <= 1'b0;
    layer0_outputs(1626) <= b and not a;
    layer0_outputs(1627) <= not (a and b);
    layer0_outputs(1628) <= a xor b;
    layer0_outputs(1629) <= b and not a;
    layer0_outputs(1630) <= b;
    layer0_outputs(1631) <= not a;
    layer0_outputs(1632) <= b;
    layer0_outputs(1633) <= not a or b;
    layer0_outputs(1634) <= not a or b;
    layer0_outputs(1635) <= not a or b;
    layer0_outputs(1636) <= 1'b1;
    layer0_outputs(1637) <= not a or b;
    layer0_outputs(1638) <= not a;
    layer0_outputs(1639) <= not (a and b);
    layer0_outputs(1640) <= not (a and b);
    layer0_outputs(1641) <= a xor b;
    layer0_outputs(1642) <= not a;
    layer0_outputs(1643) <= not b or a;
    layer0_outputs(1644) <= a or b;
    layer0_outputs(1645) <= b;
    layer0_outputs(1646) <= a or b;
    layer0_outputs(1647) <= b;
    layer0_outputs(1648) <= not (a or b);
    layer0_outputs(1649) <= b;
    layer0_outputs(1650) <= a or b;
    layer0_outputs(1651) <= not (a xor b);
    layer0_outputs(1652) <= not b or a;
    layer0_outputs(1653) <= a and not b;
    layer0_outputs(1654) <= a and b;
    layer0_outputs(1655) <= a xor b;
    layer0_outputs(1656) <= not b;
    layer0_outputs(1657) <= a xor b;
    layer0_outputs(1658) <= not b or a;
    layer0_outputs(1659) <= not (a xor b);
    layer0_outputs(1660) <= not a;
    layer0_outputs(1661) <= a;
    layer0_outputs(1662) <= 1'b0;
    layer0_outputs(1663) <= a and not b;
    layer0_outputs(1664) <= not (a and b);
    layer0_outputs(1665) <= not a;
    layer0_outputs(1666) <= not a or b;
    layer0_outputs(1667) <= a;
    layer0_outputs(1668) <= b;
    layer0_outputs(1669) <= not a;
    layer0_outputs(1670) <= not b or a;
    layer0_outputs(1671) <= not b;
    layer0_outputs(1672) <= a and not b;
    layer0_outputs(1673) <= a;
    layer0_outputs(1674) <= a and b;
    layer0_outputs(1675) <= not b or a;
    layer0_outputs(1676) <= not (a xor b);
    layer0_outputs(1677) <= b;
    layer0_outputs(1678) <= not b or a;
    layer0_outputs(1679) <= a or b;
    layer0_outputs(1680) <= a and b;
    layer0_outputs(1681) <= a;
    layer0_outputs(1682) <= a;
    layer0_outputs(1683) <= a and b;
    layer0_outputs(1684) <= not a or b;
    layer0_outputs(1685) <= a and b;
    layer0_outputs(1686) <= a and b;
    layer0_outputs(1687) <= not b;
    layer0_outputs(1688) <= a or b;
    layer0_outputs(1689) <= b;
    layer0_outputs(1690) <= not (a or b);
    layer0_outputs(1691) <= a or b;
    layer0_outputs(1692) <= not a;
    layer0_outputs(1693) <= not (a xor b);
    layer0_outputs(1694) <= not b or a;
    layer0_outputs(1695) <= not b;
    layer0_outputs(1696) <= a;
    layer0_outputs(1697) <= not a;
    layer0_outputs(1698) <= a and not b;
    layer0_outputs(1699) <= not (a xor b);
    layer0_outputs(1700) <= a or b;
    layer0_outputs(1701) <= a xor b;
    layer0_outputs(1702) <= b;
    layer0_outputs(1703) <= not b;
    layer0_outputs(1704) <= a and not b;
    layer0_outputs(1705) <= b;
    layer0_outputs(1706) <= b;
    layer0_outputs(1707) <= a and b;
    layer0_outputs(1708) <= b;
    layer0_outputs(1709) <= 1'b1;
    layer0_outputs(1710) <= b;
    layer0_outputs(1711) <= b and not a;
    layer0_outputs(1712) <= 1'b1;
    layer0_outputs(1713) <= a and b;
    layer0_outputs(1714) <= 1'b0;
    layer0_outputs(1715) <= not (a or b);
    layer0_outputs(1716) <= a or b;
    layer0_outputs(1717) <= a;
    layer0_outputs(1718) <= a xor b;
    layer0_outputs(1719) <= a or b;
    layer0_outputs(1720) <= not a;
    layer0_outputs(1721) <= not (a or b);
    layer0_outputs(1722) <= not (a and b);
    layer0_outputs(1723) <= b and not a;
    layer0_outputs(1724) <= a or b;
    layer0_outputs(1725) <= a and not b;
    layer0_outputs(1726) <= not a;
    layer0_outputs(1727) <= not a or b;
    layer0_outputs(1728) <= a xor b;
    layer0_outputs(1729) <= not (a or b);
    layer0_outputs(1730) <= a;
    layer0_outputs(1731) <= not (a xor b);
    layer0_outputs(1732) <= b;
    layer0_outputs(1733) <= a or b;
    layer0_outputs(1734) <= 1'b1;
    layer0_outputs(1735) <= 1'b1;
    layer0_outputs(1736) <= a and b;
    layer0_outputs(1737) <= not a;
    layer0_outputs(1738) <= not a or b;
    layer0_outputs(1739) <= a xor b;
    layer0_outputs(1740) <= not (a xor b);
    layer0_outputs(1741) <= a;
    layer0_outputs(1742) <= b;
    layer0_outputs(1743) <= not b or a;
    layer0_outputs(1744) <= b;
    layer0_outputs(1745) <= not b or a;
    layer0_outputs(1746) <= not b or a;
    layer0_outputs(1747) <= b and not a;
    layer0_outputs(1748) <= not a or b;
    layer0_outputs(1749) <= not (a and b);
    layer0_outputs(1750) <= a or b;
    layer0_outputs(1751) <= not (a xor b);
    layer0_outputs(1752) <= not (a xor b);
    layer0_outputs(1753) <= 1'b0;
    layer0_outputs(1754) <= 1'b0;
    layer0_outputs(1755) <= b and not a;
    layer0_outputs(1756) <= not (a or b);
    layer0_outputs(1757) <= not a or b;
    layer0_outputs(1758) <= not (a xor b);
    layer0_outputs(1759) <= b and not a;
    layer0_outputs(1760) <= a and not b;
    layer0_outputs(1761) <= not b or a;
    layer0_outputs(1762) <= not b or a;
    layer0_outputs(1763) <= not (a and b);
    layer0_outputs(1764) <= not a;
    layer0_outputs(1765) <= b;
    layer0_outputs(1766) <= not b;
    layer0_outputs(1767) <= not (a or b);
    layer0_outputs(1768) <= not a or b;
    layer0_outputs(1769) <= a or b;
    layer0_outputs(1770) <= a and not b;
    layer0_outputs(1771) <= b;
    layer0_outputs(1772) <= b and not a;
    layer0_outputs(1773) <= a;
    layer0_outputs(1774) <= not (a or b);
    layer0_outputs(1775) <= 1'b0;
    layer0_outputs(1776) <= not (a xor b);
    layer0_outputs(1777) <= a;
    layer0_outputs(1778) <= a;
    layer0_outputs(1779) <= not a or b;
    layer0_outputs(1780) <= not b;
    layer0_outputs(1781) <= b and not a;
    layer0_outputs(1782) <= not (a or b);
    layer0_outputs(1783) <= not (a xor b);
    layer0_outputs(1784) <= a;
    layer0_outputs(1785) <= a xor b;
    layer0_outputs(1786) <= not (a and b);
    layer0_outputs(1787) <= not b;
    layer0_outputs(1788) <= not a;
    layer0_outputs(1789) <= not (a or b);
    layer0_outputs(1790) <= a or b;
    layer0_outputs(1791) <= not (a or b);
    layer0_outputs(1792) <= not a;
    layer0_outputs(1793) <= not b or a;
    layer0_outputs(1794) <= not (a xor b);
    layer0_outputs(1795) <= not b;
    layer0_outputs(1796) <= 1'b0;
    layer0_outputs(1797) <= not a or b;
    layer0_outputs(1798) <= not b;
    layer0_outputs(1799) <= not (a and b);
    layer0_outputs(1800) <= not (a and b);
    layer0_outputs(1801) <= not a;
    layer0_outputs(1802) <= 1'b1;
    layer0_outputs(1803) <= not a or b;
    layer0_outputs(1804) <= not (a xor b);
    layer0_outputs(1805) <= b;
    layer0_outputs(1806) <= not (a or b);
    layer0_outputs(1807) <= not b or a;
    layer0_outputs(1808) <= b and not a;
    layer0_outputs(1809) <= a and not b;
    layer0_outputs(1810) <= not (a or b);
    layer0_outputs(1811) <= 1'b1;
    layer0_outputs(1812) <= not (a or b);
    layer0_outputs(1813) <= not (a or b);
    layer0_outputs(1814) <= not a;
    layer0_outputs(1815) <= not (a xor b);
    layer0_outputs(1816) <= a xor b;
    layer0_outputs(1817) <= a or b;
    layer0_outputs(1818) <= not (a xor b);
    layer0_outputs(1819) <= not (a or b);
    layer0_outputs(1820) <= b;
    layer0_outputs(1821) <= not a;
    layer0_outputs(1822) <= b;
    layer0_outputs(1823) <= not (a and b);
    layer0_outputs(1824) <= b;
    layer0_outputs(1825) <= b;
    layer0_outputs(1826) <= a and b;
    layer0_outputs(1827) <= b;
    layer0_outputs(1828) <= not b;
    layer0_outputs(1829) <= b;
    layer0_outputs(1830) <= 1'b0;
    layer0_outputs(1831) <= 1'b0;
    layer0_outputs(1832) <= not (a and b);
    layer0_outputs(1833) <= b and not a;
    layer0_outputs(1834) <= a or b;
    layer0_outputs(1835) <= a and not b;
    layer0_outputs(1836) <= not a;
    layer0_outputs(1837) <= 1'b0;
    layer0_outputs(1838) <= 1'b0;
    layer0_outputs(1839) <= not (a or b);
    layer0_outputs(1840) <= b and not a;
    layer0_outputs(1841) <= b;
    layer0_outputs(1842) <= a xor b;
    layer0_outputs(1843) <= not (a and b);
    layer0_outputs(1844) <= not (a and b);
    layer0_outputs(1845) <= a xor b;
    layer0_outputs(1846) <= not (a xor b);
    layer0_outputs(1847) <= not a or b;
    layer0_outputs(1848) <= a or b;
    layer0_outputs(1849) <= b and not a;
    layer0_outputs(1850) <= b and not a;
    layer0_outputs(1851) <= a and b;
    layer0_outputs(1852) <= 1'b0;
    layer0_outputs(1853) <= a;
    layer0_outputs(1854) <= a or b;
    layer0_outputs(1855) <= not a;
    layer0_outputs(1856) <= not (a and b);
    layer0_outputs(1857) <= not (a or b);
    layer0_outputs(1858) <= a and not b;
    layer0_outputs(1859) <= not b;
    layer0_outputs(1860) <= a xor b;
    layer0_outputs(1861) <= b and not a;
    layer0_outputs(1862) <= not b;
    layer0_outputs(1863) <= b;
    layer0_outputs(1864) <= not b;
    layer0_outputs(1865) <= not b;
    layer0_outputs(1866) <= not b or a;
    layer0_outputs(1867) <= not b;
    layer0_outputs(1868) <= 1'b1;
    layer0_outputs(1869) <= a;
    layer0_outputs(1870) <= b;
    layer0_outputs(1871) <= a or b;
    layer0_outputs(1872) <= a and b;
    layer0_outputs(1873) <= 1'b1;
    layer0_outputs(1874) <= a;
    layer0_outputs(1875) <= a xor b;
    layer0_outputs(1876) <= b and not a;
    layer0_outputs(1877) <= a and b;
    layer0_outputs(1878) <= a or b;
    layer0_outputs(1879) <= a xor b;
    layer0_outputs(1880) <= not a or b;
    layer0_outputs(1881) <= b;
    layer0_outputs(1882) <= a or b;
    layer0_outputs(1883) <= a or b;
    layer0_outputs(1884) <= not (a or b);
    layer0_outputs(1885) <= a or b;
    layer0_outputs(1886) <= not b;
    layer0_outputs(1887) <= a and not b;
    layer0_outputs(1888) <= b and not a;
    layer0_outputs(1889) <= not b;
    layer0_outputs(1890) <= a or b;
    layer0_outputs(1891) <= 1'b0;
    layer0_outputs(1892) <= b;
    layer0_outputs(1893) <= b and not a;
    layer0_outputs(1894) <= a or b;
    layer0_outputs(1895) <= b;
    layer0_outputs(1896) <= not a;
    layer0_outputs(1897) <= not a;
    layer0_outputs(1898) <= not (a xor b);
    layer0_outputs(1899) <= a or b;
    layer0_outputs(1900) <= not (a or b);
    layer0_outputs(1901) <= not (a xor b);
    layer0_outputs(1902) <= not b or a;
    layer0_outputs(1903) <= b;
    layer0_outputs(1904) <= not (a or b);
    layer0_outputs(1905) <= not (a or b);
    layer0_outputs(1906) <= not (a or b);
    layer0_outputs(1907) <= b;
    layer0_outputs(1908) <= not a;
    layer0_outputs(1909) <= not b or a;
    layer0_outputs(1910) <= a and not b;
    layer0_outputs(1911) <= b and not a;
    layer0_outputs(1912) <= not (a or b);
    layer0_outputs(1913) <= b and not a;
    layer0_outputs(1914) <= not a or b;
    layer0_outputs(1915) <= a or b;
    layer0_outputs(1916) <= not b or a;
    layer0_outputs(1917) <= a or b;
    layer0_outputs(1918) <= b;
    layer0_outputs(1919) <= not b or a;
    layer0_outputs(1920) <= a or b;
    layer0_outputs(1921) <= not a;
    layer0_outputs(1922) <= a and not b;
    layer0_outputs(1923) <= 1'b1;
    layer0_outputs(1924) <= not b or a;
    layer0_outputs(1925) <= not b;
    layer0_outputs(1926) <= not a;
    layer0_outputs(1927) <= not (a and b);
    layer0_outputs(1928) <= a;
    layer0_outputs(1929) <= a or b;
    layer0_outputs(1930) <= not a or b;
    layer0_outputs(1931) <= 1'b0;
    layer0_outputs(1932) <= a xor b;
    layer0_outputs(1933) <= not a;
    layer0_outputs(1934) <= not a;
    layer0_outputs(1935) <= not (a or b);
    layer0_outputs(1936) <= not (a xor b);
    layer0_outputs(1937) <= not (a and b);
    layer0_outputs(1938) <= b;
    layer0_outputs(1939) <= not (a or b);
    layer0_outputs(1940) <= b and not a;
    layer0_outputs(1941) <= not (a or b);
    layer0_outputs(1942) <= a or b;
    layer0_outputs(1943) <= not b;
    layer0_outputs(1944) <= not b;
    layer0_outputs(1945) <= not b or a;
    layer0_outputs(1946) <= a;
    layer0_outputs(1947) <= a;
    layer0_outputs(1948) <= 1'b1;
    layer0_outputs(1949) <= a;
    layer0_outputs(1950) <= 1'b1;
    layer0_outputs(1951) <= not b or a;
    layer0_outputs(1952) <= not b;
    layer0_outputs(1953) <= not (a or b);
    layer0_outputs(1954) <= 1'b0;
    layer0_outputs(1955) <= not a;
    layer0_outputs(1956) <= not b;
    layer0_outputs(1957) <= not (a xor b);
    layer0_outputs(1958) <= a and not b;
    layer0_outputs(1959) <= 1'b1;
    layer0_outputs(1960) <= not a or b;
    layer0_outputs(1961) <= a or b;
    layer0_outputs(1962) <= not b;
    layer0_outputs(1963) <= a xor b;
    layer0_outputs(1964) <= not (a and b);
    layer0_outputs(1965) <= a and b;
    layer0_outputs(1966) <= not a;
    layer0_outputs(1967) <= not (a and b);
    layer0_outputs(1968) <= a and b;
    layer0_outputs(1969) <= b and not a;
    layer0_outputs(1970) <= a or b;
    layer0_outputs(1971) <= a and b;
    layer0_outputs(1972) <= not (a or b);
    layer0_outputs(1973) <= a and b;
    layer0_outputs(1974) <= a or b;
    layer0_outputs(1975) <= a and not b;
    layer0_outputs(1976) <= a xor b;
    layer0_outputs(1977) <= b;
    layer0_outputs(1978) <= a and not b;
    layer0_outputs(1979) <= not b or a;
    layer0_outputs(1980) <= not (a or b);
    layer0_outputs(1981) <= b and not a;
    layer0_outputs(1982) <= not b;
    layer0_outputs(1983) <= a or b;
    layer0_outputs(1984) <= a and b;
    layer0_outputs(1985) <= 1'b0;
    layer0_outputs(1986) <= a;
    layer0_outputs(1987) <= not b or a;
    layer0_outputs(1988) <= not a;
    layer0_outputs(1989) <= not (a xor b);
    layer0_outputs(1990) <= b;
    layer0_outputs(1991) <= a or b;
    layer0_outputs(1992) <= 1'b0;
    layer0_outputs(1993) <= a xor b;
    layer0_outputs(1994) <= a and b;
    layer0_outputs(1995) <= not (a and b);
    layer0_outputs(1996) <= not a or b;
    layer0_outputs(1997) <= 1'b0;
    layer0_outputs(1998) <= a and not b;
    layer0_outputs(1999) <= not (a or b);
    layer0_outputs(2000) <= not b;
    layer0_outputs(2001) <= 1'b0;
    layer0_outputs(2002) <= a;
    layer0_outputs(2003) <= a or b;
    layer0_outputs(2004) <= not a;
    layer0_outputs(2005) <= not a or b;
    layer0_outputs(2006) <= not b;
    layer0_outputs(2007) <= 1'b0;
    layer0_outputs(2008) <= b and not a;
    layer0_outputs(2009) <= not (a or b);
    layer0_outputs(2010) <= a and b;
    layer0_outputs(2011) <= 1'b0;
    layer0_outputs(2012) <= b;
    layer0_outputs(2013) <= 1'b1;
    layer0_outputs(2014) <= not (a xor b);
    layer0_outputs(2015) <= not (a or b);
    layer0_outputs(2016) <= a and not b;
    layer0_outputs(2017) <= a and not b;
    layer0_outputs(2018) <= b and not a;
    layer0_outputs(2019) <= a and b;
    layer0_outputs(2020) <= a or b;
    layer0_outputs(2021) <= not (a or b);
    layer0_outputs(2022) <= not b or a;
    layer0_outputs(2023) <= not (a or b);
    layer0_outputs(2024) <= b;
    layer0_outputs(2025) <= not (a and b);
    layer0_outputs(2026) <= not (a or b);
    layer0_outputs(2027) <= not b;
    layer0_outputs(2028) <= a and b;
    layer0_outputs(2029) <= a;
    layer0_outputs(2030) <= a or b;
    layer0_outputs(2031) <= not (a or b);
    layer0_outputs(2032) <= not (a or b);
    layer0_outputs(2033) <= a;
    layer0_outputs(2034) <= b and not a;
    layer0_outputs(2035) <= b and not a;
    layer0_outputs(2036) <= not a or b;
    layer0_outputs(2037) <= not b;
    layer0_outputs(2038) <= not b;
    layer0_outputs(2039) <= a or b;
    layer0_outputs(2040) <= not (a and b);
    layer0_outputs(2041) <= a and not b;
    layer0_outputs(2042) <= a;
    layer0_outputs(2043) <= b and not a;
    layer0_outputs(2044) <= b;
    layer0_outputs(2045) <= a or b;
    layer0_outputs(2046) <= not (a xor b);
    layer0_outputs(2047) <= not (a xor b);
    layer0_outputs(2048) <= not (a or b);
    layer0_outputs(2049) <= not a or b;
    layer0_outputs(2050) <= not (a xor b);
    layer0_outputs(2051) <= a xor b;
    layer0_outputs(2052) <= not (a xor b);
    layer0_outputs(2053) <= not (a or b);
    layer0_outputs(2054) <= not a;
    layer0_outputs(2055) <= a or b;
    layer0_outputs(2056) <= not a or b;
    layer0_outputs(2057) <= not (a or b);
    layer0_outputs(2058) <= not a or b;
    layer0_outputs(2059) <= a and not b;
    layer0_outputs(2060) <= not b or a;
    layer0_outputs(2061) <= not (a or b);
    layer0_outputs(2062) <= not a or b;
    layer0_outputs(2063) <= not b;
    layer0_outputs(2064) <= not a or b;
    layer0_outputs(2065) <= not b;
    layer0_outputs(2066) <= b;
    layer0_outputs(2067) <= not (a xor b);
    layer0_outputs(2068) <= a or b;
    layer0_outputs(2069) <= a or b;
    layer0_outputs(2070) <= a or b;
    layer0_outputs(2071) <= a and not b;
    layer0_outputs(2072) <= not a or b;
    layer0_outputs(2073) <= b and not a;
    layer0_outputs(2074) <= a and not b;
    layer0_outputs(2075) <= a xor b;
    layer0_outputs(2076) <= a or b;
    layer0_outputs(2077) <= a;
    layer0_outputs(2078) <= not (a or b);
    layer0_outputs(2079) <= not (a xor b);
    layer0_outputs(2080) <= a;
    layer0_outputs(2081) <= not a;
    layer0_outputs(2082) <= not b or a;
    layer0_outputs(2083) <= b and not a;
    layer0_outputs(2084) <= a and b;
    layer0_outputs(2085) <= a;
    layer0_outputs(2086) <= not a or b;
    layer0_outputs(2087) <= a;
    layer0_outputs(2088) <= not a or b;
    layer0_outputs(2089) <= not (a or b);
    layer0_outputs(2090) <= not (a or b);
    layer0_outputs(2091) <= a;
    layer0_outputs(2092) <= a xor b;
    layer0_outputs(2093) <= not a or b;
    layer0_outputs(2094) <= a xor b;
    layer0_outputs(2095) <= not (a xor b);
    layer0_outputs(2096) <= b;
    layer0_outputs(2097) <= b;
    layer0_outputs(2098) <= not a or b;
    layer0_outputs(2099) <= a and b;
    layer0_outputs(2100) <= not b;
    layer0_outputs(2101) <= a and b;
    layer0_outputs(2102) <= b;
    layer0_outputs(2103) <= a or b;
    layer0_outputs(2104) <= not (a xor b);
    layer0_outputs(2105) <= not b;
    layer0_outputs(2106) <= a and b;
    layer0_outputs(2107) <= a and not b;
    layer0_outputs(2108) <= a and b;
    layer0_outputs(2109) <= not a;
    layer0_outputs(2110) <= a or b;
    layer0_outputs(2111) <= a and b;
    layer0_outputs(2112) <= a;
    layer0_outputs(2113) <= not (a and b);
    layer0_outputs(2114) <= b and not a;
    layer0_outputs(2115) <= not (a xor b);
    layer0_outputs(2116) <= b;
    layer0_outputs(2117) <= not b;
    layer0_outputs(2118) <= a or b;
    layer0_outputs(2119) <= not (a xor b);
    layer0_outputs(2120) <= b;
    layer0_outputs(2121) <= 1'b1;
    layer0_outputs(2122) <= not b;
    layer0_outputs(2123) <= not b;
    layer0_outputs(2124) <= not (a and b);
    layer0_outputs(2125) <= b and not a;
    layer0_outputs(2126) <= a and b;
    layer0_outputs(2127) <= b;
    layer0_outputs(2128) <= not b or a;
    layer0_outputs(2129) <= a xor b;
    layer0_outputs(2130) <= not b or a;
    layer0_outputs(2131) <= b;
    layer0_outputs(2132) <= b;
    layer0_outputs(2133) <= a or b;
    layer0_outputs(2134) <= not (a and b);
    layer0_outputs(2135) <= a or b;
    layer0_outputs(2136) <= not b or a;
    layer0_outputs(2137) <= a or b;
    layer0_outputs(2138) <= a and not b;
    layer0_outputs(2139) <= a or b;
    layer0_outputs(2140) <= b;
    layer0_outputs(2141) <= b and not a;
    layer0_outputs(2142) <= not (a xor b);
    layer0_outputs(2143) <= 1'b0;
    layer0_outputs(2144) <= a or b;
    layer0_outputs(2145) <= not a or b;
    layer0_outputs(2146) <= not a;
    layer0_outputs(2147) <= a and not b;
    layer0_outputs(2148) <= a or b;
    layer0_outputs(2149) <= not a;
    layer0_outputs(2150) <= not b or a;
    layer0_outputs(2151) <= not b;
    layer0_outputs(2152) <= not a;
    layer0_outputs(2153) <= a or b;
    layer0_outputs(2154) <= a xor b;
    layer0_outputs(2155) <= a or b;
    layer0_outputs(2156) <= not b or a;
    layer0_outputs(2157) <= not a or b;
    layer0_outputs(2158) <= b;
    layer0_outputs(2159) <= not (a and b);
    layer0_outputs(2160) <= a and b;
    layer0_outputs(2161) <= not a or b;
    layer0_outputs(2162) <= a or b;
    layer0_outputs(2163) <= not a;
    layer0_outputs(2164) <= not a or b;
    layer0_outputs(2165) <= not (a xor b);
    layer0_outputs(2166) <= a xor b;
    layer0_outputs(2167) <= a and not b;
    layer0_outputs(2168) <= not a;
    layer0_outputs(2169) <= 1'b0;
    layer0_outputs(2170) <= a xor b;
    layer0_outputs(2171) <= not (a or b);
    layer0_outputs(2172) <= a;
    layer0_outputs(2173) <= not (a xor b);
    layer0_outputs(2174) <= a or b;
    layer0_outputs(2175) <= 1'b0;
    layer0_outputs(2176) <= not (a or b);
    layer0_outputs(2177) <= a;
    layer0_outputs(2178) <= 1'b1;
    layer0_outputs(2179) <= a or b;
    layer0_outputs(2180) <= b and not a;
    layer0_outputs(2181) <= not b;
    layer0_outputs(2182) <= a;
    layer0_outputs(2183) <= not (a or b);
    layer0_outputs(2184) <= 1'b0;
    layer0_outputs(2185) <= not (a or b);
    layer0_outputs(2186) <= b;
    layer0_outputs(2187) <= b;
    layer0_outputs(2188) <= not a;
    layer0_outputs(2189) <= b;
    layer0_outputs(2190) <= a and not b;
    layer0_outputs(2191) <= b;
    layer0_outputs(2192) <= b;
    layer0_outputs(2193) <= b and not a;
    layer0_outputs(2194) <= 1'b0;
    layer0_outputs(2195) <= not (a or b);
    layer0_outputs(2196) <= not a;
    layer0_outputs(2197) <= a and not b;
    layer0_outputs(2198) <= not (a or b);
    layer0_outputs(2199) <= a and b;
    layer0_outputs(2200) <= not b or a;
    layer0_outputs(2201) <= not b or a;
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= a;
    layer0_outputs(2204) <= a and not b;
    layer0_outputs(2205) <= not (a or b);
    layer0_outputs(2206) <= not a or b;
    layer0_outputs(2207) <= not (a or b);
    layer0_outputs(2208) <= a or b;
    layer0_outputs(2209) <= a and not b;
    layer0_outputs(2210) <= a or b;
    layer0_outputs(2211) <= a;
    layer0_outputs(2212) <= b;
    layer0_outputs(2213) <= a xor b;
    layer0_outputs(2214) <= 1'b0;
    layer0_outputs(2215) <= a xor b;
    layer0_outputs(2216) <= a or b;
    layer0_outputs(2217) <= a or b;
    layer0_outputs(2218) <= not b;
    layer0_outputs(2219) <= not b;
    layer0_outputs(2220) <= 1'b0;
    layer0_outputs(2221) <= b and not a;
    layer0_outputs(2222) <= a xor b;
    layer0_outputs(2223) <= not a or b;
    layer0_outputs(2224) <= b and not a;
    layer0_outputs(2225) <= a and not b;
    layer0_outputs(2226) <= not a or b;
    layer0_outputs(2227) <= a and b;
    layer0_outputs(2228) <= 1'b0;
    layer0_outputs(2229) <= not b;
    layer0_outputs(2230) <= a;
    layer0_outputs(2231) <= not a;
    layer0_outputs(2232) <= not b;
    layer0_outputs(2233) <= a or b;
    layer0_outputs(2234) <= a and b;
    layer0_outputs(2235) <= a and not b;
    layer0_outputs(2236) <= b;
    layer0_outputs(2237) <= a xor b;
    layer0_outputs(2238) <= a and b;
    layer0_outputs(2239) <= not (a xor b);
    layer0_outputs(2240) <= a and b;
    layer0_outputs(2241) <= 1'b0;
    layer0_outputs(2242) <= a or b;
    layer0_outputs(2243) <= not (a or b);
    layer0_outputs(2244) <= a and not b;
    layer0_outputs(2245) <= not b or a;
    layer0_outputs(2246) <= 1'b1;
    layer0_outputs(2247) <= not a or b;
    layer0_outputs(2248) <= a or b;
    layer0_outputs(2249) <= a or b;
    layer0_outputs(2250) <= not (a or b);
    layer0_outputs(2251) <= not b or a;
    layer0_outputs(2252) <= not a;
    layer0_outputs(2253) <= not (a and b);
    layer0_outputs(2254) <= not (a or b);
    layer0_outputs(2255) <= b and not a;
    layer0_outputs(2256) <= a and b;
    layer0_outputs(2257) <= a or b;
    layer0_outputs(2258) <= not b or a;
    layer0_outputs(2259) <= b;
    layer0_outputs(2260) <= not (a or b);
    layer0_outputs(2261) <= not (a xor b);
    layer0_outputs(2262) <= a and not b;
    layer0_outputs(2263) <= b;
    layer0_outputs(2264) <= not (a and b);
    layer0_outputs(2265) <= a or b;
    layer0_outputs(2266) <= not a;
    layer0_outputs(2267) <= not b;
    layer0_outputs(2268) <= not a;
    layer0_outputs(2269) <= a and not b;
    layer0_outputs(2270) <= 1'b1;
    layer0_outputs(2271) <= a and not b;
    layer0_outputs(2272) <= a xor b;
    layer0_outputs(2273) <= not (a xor b);
    layer0_outputs(2274) <= b;
    layer0_outputs(2275) <= b;
    layer0_outputs(2276) <= not a;
    layer0_outputs(2277) <= a;
    layer0_outputs(2278) <= a;
    layer0_outputs(2279) <= a or b;
    layer0_outputs(2280) <= not a or b;
    layer0_outputs(2281) <= not b or a;
    layer0_outputs(2282) <= not b;
    layer0_outputs(2283) <= a;
    layer0_outputs(2284) <= not a;
    layer0_outputs(2285) <= a and not b;
    layer0_outputs(2286) <= a;
    layer0_outputs(2287) <= 1'b1;
    layer0_outputs(2288) <= a or b;
    layer0_outputs(2289) <= a xor b;
    layer0_outputs(2290) <= not (a or b);
    layer0_outputs(2291) <= not a;
    layer0_outputs(2292) <= a or b;
    layer0_outputs(2293) <= not b;
    layer0_outputs(2294) <= not (a or b);
    layer0_outputs(2295) <= b;
    layer0_outputs(2296) <= not (a or b);
    layer0_outputs(2297) <= not b or a;
    layer0_outputs(2298) <= a or b;
    layer0_outputs(2299) <= not a;
    layer0_outputs(2300) <= not b or a;
    layer0_outputs(2301) <= 1'b1;
    layer0_outputs(2302) <= a or b;
    layer0_outputs(2303) <= not b or a;
    layer0_outputs(2304) <= a;
    layer0_outputs(2305) <= 1'b1;
    layer0_outputs(2306) <= not b or a;
    layer0_outputs(2307) <= a;
    layer0_outputs(2308) <= not a;
    layer0_outputs(2309) <= not a;
    layer0_outputs(2310) <= a and b;
    layer0_outputs(2311) <= b;
    layer0_outputs(2312) <= a or b;
    layer0_outputs(2313) <= a xor b;
    layer0_outputs(2314) <= a and not b;
    layer0_outputs(2315) <= not (a or b);
    layer0_outputs(2316) <= a;
    layer0_outputs(2317) <= a and not b;
    layer0_outputs(2318) <= b;
    layer0_outputs(2319) <= 1'b0;
    layer0_outputs(2320) <= a or b;
    layer0_outputs(2321) <= not (a or b);
    layer0_outputs(2322) <= b and not a;
    layer0_outputs(2323) <= a and b;
    layer0_outputs(2324) <= a xor b;
    layer0_outputs(2325) <= a or b;
    layer0_outputs(2326) <= not b or a;
    layer0_outputs(2327) <= a or b;
    layer0_outputs(2328) <= not b;
    layer0_outputs(2329) <= not (a xor b);
    layer0_outputs(2330) <= not (a and b);
    layer0_outputs(2331) <= a and not b;
    layer0_outputs(2332) <= not (a or b);
    layer0_outputs(2333) <= a;
    layer0_outputs(2334) <= a and b;
    layer0_outputs(2335) <= not (a and b);
    layer0_outputs(2336) <= b and not a;
    layer0_outputs(2337) <= not a;
    layer0_outputs(2338) <= 1'b0;
    layer0_outputs(2339) <= not b or a;
    layer0_outputs(2340) <= not (a xor b);
    layer0_outputs(2341) <= b and not a;
    layer0_outputs(2342) <= a;
    layer0_outputs(2343) <= not b or a;
    layer0_outputs(2344) <= a and not b;
    layer0_outputs(2345) <= not (a xor b);
    layer0_outputs(2346) <= not b;
    layer0_outputs(2347) <= not (a or b);
    layer0_outputs(2348) <= a or b;
    layer0_outputs(2349) <= not (a xor b);
    layer0_outputs(2350) <= b and not a;
    layer0_outputs(2351) <= not (a or b);
    layer0_outputs(2352) <= a;
    layer0_outputs(2353) <= a;
    layer0_outputs(2354) <= not b or a;
    layer0_outputs(2355) <= a and not b;
    layer0_outputs(2356) <= a xor b;
    layer0_outputs(2357) <= b;
    layer0_outputs(2358) <= not b;
    layer0_outputs(2359) <= not b or a;
    layer0_outputs(2360) <= 1'b0;
    layer0_outputs(2361) <= not (a xor b);
    layer0_outputs(2362) <= b;
    layer0_outputs(2363) <= a and b;
    layer0_outputs(2364) <= a;
    layer0_outputs(2365) <= a or b;
    layer0_outputs(2366) <= a xor b;
    layer0_outputs(2367) <= a;
    layer0_outputs(2368) <= not (a and b);
    layer0_outputs(2369) <= not (a xor b);
    layer0_outputs(2370) <= a or b;
    layer0_outputs(2371) <= not (a or b);
    layer0_outputs(2372) <= not b;
    layer0_outputs(2373) <= 1'b1;
    layer0_outputs(2374) <= b;
    layer0_outputs(2375) <= a and b;
    layer0_outputs(2376) <= not b;
    layer0_outputs(2377) <= 1'b0;
    layer0_outputs(2378) <= not a;
    layer0_outputs(2379) <= a xor b;
    layer0_outputs(2380) <= not (a or b);
    layer0_outputs(2381) <= not b or a;
    layer0_outputs(2382) <= not b or a;
    layer0_outputs(2383) <= a;
    layer0_outputs(2384) <= not (a and b);
    layer0_outputs(2385) <= not a;
    layer0_outputs(2386) <= a and not b;
    layer0_outputs(2387) <= a xor b;
    layer0_outputs(2388) <= not b;
    layer0_outputs(2389) <= 1'b1;
    layer0_outputs(2390) <= a xor b;
    layer0_outputs(2391) <= a;
    layer0_outputs(2392) <= b;
    layer0_outputs(2393) <= b;
    layer0_outputs(2394) <= not b;
    layer0_outputs(2395) <= a;
    layer0_outputs(2396) <= not (a xor b);
    layer0_outputs(2397) <= b;
    layer0_outputs(2398) <= a xor b;
    layer0_outputs(2399) <= a xor b;
    layer0_outputs(2400) <= a and not b;
    layer0_outputs(2401) <= 1'b0;
    layer0_outputs(2402) <= b;
    layer0_outputs(2403) <= a or b;
    layer0_outputs(2404) <= b and not a;
    layer0_outputs(2405) <= not a or b;
    layer0_outputs(2406) <= not (a xor b);
    layer0_outputs(2407) <= not b or a;
    layer0_outputs(2408) <= 1'b1;
    layer0_outputs(2409) <= not (a and b);
    layer0_outputs(2410) <= a or b;
    layer0_outputs(2411) <= not (a and b);
    layer0_outputs(2412) <= a;
    layer0_outputs(2413) <= not a or b;
    layer0_outputs(2414) <= a xor b;
    layer0_outputs(2415) <= not (a or b);
    layer0_outputs(2416) <= not (a or b);
    layer0_outputs(2417) <= 1'b1;
    layer0_outputs(2418) <= not b;
    layer0_outputs(2419) <= a and not b;
    layer0_outputs(2420) <= b and not a;
    layer0_outputs(2421) <= not a;
    layer0_outputs(2422) <= not b;
    layer0_outputs(2423) <= a or b;
    layer0_outputs(2424) <= not a or b;
    layer0_outputs(2425) <= 1'b0;
    layer0_outputs(2426) <= not b;
    layer0_outputs(2427) <= a and not b;
    layer0_outputs(2428) <= not b or a;
    layer0_outputs(2429) <= not b;
    layer0_outputs(2430) <= not a;
    layer0_outputs(2431) <= a xor b;
    layer0_outputs(2432) <= b;
    layer0_outputs(2433) <= not a or b;
    layer0_outputs(2434) <= not a;
    layer0_outputs(2435) <= not b;
    layer0_outputs(2436) <= a and b;
    layer0_outputs(2437) <= not b;
    layer0_outputs(2438) <= a and b;
    layer0_outputs(2439) <= 1'b0;
    layer0_outputs(2440) <= not b or a;
    layer0_outputs(2441) <= not (a xor b);
    layer0_outputs(2442) <= not (a and b);
    layer0_outputs(2443) <= not b or a;
    layer0_outputs(2444) <= not b or a;
    layer0_outputs(2445) <= a xor b;
    layer0_outputs(2446) <= not (a or b);
    layer0_outputs(2447) <= a xor b;
    layer0_outputs(2448) <= not b or a;
    layer0_outputs(2449) <= 1'b1;
    layer0_outputs(2450) <= a and not b;
    layer0_outputs(2451) <= 1'b1;
    layer0_outputs(2452) <= not (a or b);
    layer0_outputs(2453) <= a and b;
    layer0_outputs(2454) <= a or b;
    layer0_outputs(2455) <= a and not b;
    layer0_outputs(2456) <= a or b;
    layer0_outputs(2457) <= 1'b0;
    layer0_outputs(2458) <= a and not b;
    layer0_outputs(2459) <= 1'b1;
    layer0_outputs(2460) <= b;
    layer0_outputs(2461) <= 1'b0;
    layer0_outputs(2462) <= a xor b;
    layer0_outputs(2463) <= not a or b;
    layer0_outputs(2464) <= not b;
    layer0_outputs(2465) <= not a;
    layer0_outputs(2466) <= not a or b;
    layer0_outputs(2467) <= not a or b;
    layer0_outputs(2468) <= not (a or b);
    layer0_outputs(2469) <= not (a or b);
    layer0_outputs(2470) <= b;
    layer0_outputs(2471) <= not (a xor b);
    layer0_outputs(2472) <= a;
    layer0_outputs(2473) <= not (a or b);
    layer0_outputs(2474) <= b;
    layer0_outputs(2475) <= a and not b;
    layer0_outputs(2476) <= b;
    layer0_outputs(2477) <= not b;
    layer0_outputs(2478) <= a xor b;
    layer0_outputs(2479) <= a xor b;
    layer0_outputs(2480) <= b and not a;
    layer0_outputs(2481) <= not a;
    layer0_outputs(2482) <= not (a or b);
    layer0_outputs(2483) <= not b or a;
    layer0_outputs(2484) <= a and b;
    layer0_outputs(2485) <= not b or a;
    layer0_outputs(2486) <= not (a or b);
    layer0_outputs(2487) <= not b;
    layer0_outputs(2488) <= 1'b0;
    layer0_outputs(2489) <= a xor b;
    layer0_outputs(2490) <= a and not b;
    layer0_outputs(2491) <= not b or a;
    layer0_outputs(2492) <= 1'b1;
    layer0_outputs(2493) <= a or b;
    layer0_outputs(2494) <= b and not a;
    layer0_outputs(2495) <= not b;
    layer0_outputs(2496) <= not a;
    layer0_outputs(2497) <= a or b;
    layer0_outputs(2498) <= a or b;
    layer0_outputs(2499) <= a or b;
    layer0_outputs(2500) <= 1'b1;
    layer0_outputs(2501) <= a and not b;
    layer0_outputs(2502) <= not b or a;
    layer0_outputs(2503) <= not (a or b);
    layer0_outputs(2504) <= not b;
    layer0_outputs(2505) <= 1'b0;
    layer0_outputs(2506) <= a or b;
    layer0_outputs(2507) <= not (a or b);
    layer0_outputs(2508) <= a and b;
    layer0_outputs(2509) <= a;
    layer0_outputs(2510) <= a or b;
    layer0_outputs(2511) <= b and not a;
    layer0_outputs(2512) <= a xor b;
    layer0_outputs(2513) <= not a;
    layer0_outputs(2514) <= b and not a;
    layer0_outputs(2515) <= not a;
    layer0_outputs(2516) <= not (a xor b);
    layer0_outputs(2517) <= not b;
    layer0_outputs(2518) <= not (a or b);
    layer0_outputs(2519) <= a;
    layer0_outputs(2520) <= not (a xor b);
    layer0_outputs(2521) <= a and not b;
    layer0_outputs(2522) <= not (a and b);
    layer0_outputs(2523) <= a and not b;
    layer0_outputs(2524) <= b and not a;
    layer0_outputs(2525) <= not b;
    layer0_outputs(2526) <= a xor b;
    layer0_outputs(2527) <= a or b;
    layer0_outputs(2528) <= b and not a;
    layer0_outputs(2529) <= not (a or b);
    layer0_outputs(2530) <= 1'b1;
    layer0_outputs(2531) <= not a or b;
    layer0_outputs(2532) <= a or b;
    layer0_outputs(2533) <= a and not b;
    layer0_outputs(2534) <= b;
    layer0_outputs(2535) <= not a;
    layer0_outputs(2536) <= not b or a;
    layer0_outputs(2537) <= a xor b;
    layer0_outputs(2538) <= a and b;
    layer0_outputs(2539) <= not a;
    layer0_outputs(2540) <= b and not a;
    layer0_outputs(2541) <= 1'b0;
    layer0_outputs(2542) <= a or b;
    layer0_outputs(2543) <= not a or b;
    layer0_outputs(2544) <= a and not b;
    layer0_outputs(2545) <= a and b;
    layer0_outputs(2546) <= not b or a;
    layer0_outputs(2547) <= not (a or b);
    layer0_outputs(2548) <= a or b;
    layer0_outputs(2549) <= not (a xor b);
    layer0_outputs(2550) <= a xor b;
    layer0_outputs(2551) <= not (a and b);
    layer0_outputs(2552) <= not (a or b);
    layer0_outputs(2553) <= a;
    layer0_outputs(2554) <= not b or a;
    layer0_outputs(2555) <= a and not b;
    layer0_outputs(2556) <= not (a or b);
    layer0_outputs(2557) <= not b or a;
    layer0_outputs(2558) <= not a or b;
    layer0_outputs(2559) <= not b or a;
    layer0_outputs(2560) <= a or b;
    layer0_outputs(2561) <= not b;
    layer0_outputs(2562) <= a;
    layer0_outputs(2563) <= not (a or b);
    layer0_outputs(2564) <= not b or a;
    layer0_outputs(2565) <= not (a or b);
    layer0_outputs(2566) <= not (a xor b);
    layer0_outputs(2567) <= a and not b;
    layer0_outputs(2568) <= b and not a;
    layer0_outputs(2569) <= not (a xor b);
    layer0_outputs(2570) <= a and b;
    layer0_outputs(2571) <= not (a or b);
    layer0_outputs(2572) <= a and not b;
    layer0_outputs(2573) <= 1'b0;
    layer0_outputs(2574) <= b and not a;
    layer0_outputs(2575) <= not (a or b);
    layer0_outputs(2576) <= a;
    layer0_outputs(2577) <= 1'b0;
    layer0_outputs(2578) <= a and not b;
    layer0_outputs(2579) <= a or b;
    layer0_outputs(2580) <= not b;
    layer0_outputs(2581) <= a;
    layer0_outputs(2582) <= not (a xor b);
    layer0_outputs(2583) <= a xor b;
    layer0_outputs(2584) <= not b;
    layer0_outputs(2585) <= 1'b0;
    layer0_outputs(2586) <= b and not a;
    layer0_outputs(2587) <= not (a or b);
    layer0_outputs(2588) <= a;
    layer0_outputs(2589) <= a xor b;
    layer0_outputs(2590) <= not b or a;
    layer0_outputs(2591) <= 1'b1;
    layer0_outputs(2592) <= a and not b;
    layer0_outputs(2593) <= a;
    layer0_outputs(2594) <= a or b;
    layer0_outputs(2595) <= b and not a;
    layer0_outputs(2596) <= not a;
    layer0_outputs(2597) <= not (a or b);
    layer0_outputs(2598) <= not a;
    layer0_outputs(2599) <= 1'b0;
    layer0_outputs(2600) <= a xor b;
    layer0_outputs(2601) <= a or b;
    layer0_outputs(2602) <= a xor b;
    layer0_outputs(2603) <= b;
    layer0_outputs(2604) <= not b;
    layer0_outputs(2605) <= not a or b;
    layer0_outputs(2606) <= not (a xor b);
    layer0_outputs(2607) <= not a;
    layer0_outputs(2608) <= not (a xor b);
    layer0_outputs(2609) <= a;
    layer0_outputs(2610) <= not b;
    layer0_outputs(2611) <= b and not a;
    layer0_outputs(2612) <= a;
    layer0_outputs(2613) <= 1'b0;
    layer0_outputs(2614) <= a;
    layer0_outputs(2615) <= a and b;
    layer0_outputs(2616) <= not a;
    layer0_outputs(2617) <= a and not b;
    layer0_outputs(2618) <= a and not b;
    layer0_outputs(2619) <= a or b;
    layer0_outputs(2620) <= b;
    layer0_outputs(2621) <= a or b;
    layer0_outputs(2622) <= not b or a;
    layer0_outputs(2623) <= not b;
    layer0_outputs(2624) <= not (a xor b);
    layer0_outputs(2625) <= not a;
    layer0_outputs(2626) <= not a or b;
    layer0_outputs(2627) <= not b or a;
    layer0_outputs(2628) <= a or b;
    layer0_outputs(2629) <= not a or b;
    layer0_outputs(2630) <= b and not a;
    layer0_outputs(2631) <= 1'b1;
    layer0_outputs(2632) <= not a or b;
    layer0_outputs(2633) <= 1'b1;
    layer0_outputs(2634) <= a and not b;
    layer0_outputs(2635) <= not (a and b);
    layer0_outputs(2636) <= a and b;
    layer0_outputs(2637) <= not (a or b);
    layer0_outputs(2638) <= not b;
    layer0_outputs(2639) <= b and not a;
    layer0_outputs(2640) <= not (a and b);
    layer0_outputs(2641) <= a and not b;
    layer0_outputs(2642) <= not a;
    layer0_outputs(2643) <= a or b;
    layer0_outputs(2644) <= not a or b;
    layer0_outputs(2645) <= not a;
    layer0_outputs(2646) <= b and not a;
    layer0_outputs(2647) <= b and not a;
    layer0_outputs(2648) <= not a;
    layer0_outputs(2649) <= not b;
    layer0_outputs(2650) <= not a;
    layer0_outputs(2651) <= 1'b0;
    layer0_outputs(2652) <= a and b;
    layer0_outputs(2653) <= not (a or b);
    layer0_outputs(2654) <= b and not a;
    layer0_outputs(2655) <= not a or b;
    layer0_outputs(2656) <= a and not b;
    layer0_outputs(2657) <= b;
    layer0_outputs(2658) <= 1'b0;
    layer0_outputs(2659) <= not b or a;
    layer0_outputs(2660) <= a and b;
    layer0_outputs(2661) <= not (a and b);
    layer0_outputs(2662) <= a or b;
    layer0_outputs(2663) <= b and not a;
    layer0_outputs(2664) <= not b;
    layer0_outputs(2665) <= not b or a;
    layer0_outputs(2666) <= b;
    layer0_outputs(2667) <= 1'b0;
    layer0_outputs(2668) <= a xor b;
    layer0_outputs(2669) <= not a or b;
    layer0_outputs(2670) <= not b;
    layer0_outputs(2671) <= b;
    layer0_outputs(2672) <= b;
    layer0_outputs(2673) <= not b or a;
    layer0_outputs(2674) <= not b;
    layer0_outputs(2675) <= not (a or b);
    layer0_outputs(2676) <= not b;
    layer0_outputs(2677) <= a or b;
    layer0_outputs(2678) <= 1'b1;
    layer0_outputs(2679) <= a xor b;
    layer0_outputs(2680) <= not a or b;
    layer0_outputs(2681) <= b and not a;
    layer0_outputs(2682) <= not (a and b);
    layer0_outputs(2683) <= a or b;
    layer0_outputs(2684) <= b and not a;
    layer0_outputs(2685) <= not (a or b);
    layer0_outputs(2686) <= not b or a;
    layer0_outputs(2687) <= not (a or b);
    layer0_outputs(2688) <= not b;
    layer0_outputs(2689) <= a or b;
    layer0_outputs(2690) <= not b;
    layer0_outputs(2691) <= not a or b;
    layer0_outputs(2692) <= not (a or b);
    layer0_outputs(2693) <= not b;
    layer0_outputs(2694) <= not (a xor b);
    layer0_outputs(2695) <= not (a or b);
    layer0_outputs(2696) <= not a or b;
    layer0_outputs(2697) <= not (a or b);
    layer0_outputs(2698) <= not a or b;
    layer0_outputs(2699) <= b and not a;
    layer0_outputs(2700) <= a and b;
    layer0_outputs(2701) <= not (a or b);
    layer0_outputs(2702) <= b and not a;
    layer0_outputs(2703) <= not (a xor b);
    layer0_outputs(2704) <= not b;
    layer0_outputs(2705) <= not (a xor b);
    layer0_outputs(2706) <= not (a and b);
    layer0_outputs(2707) <= not b;
    layer0_outputs(2708) <= not a;
    layer0_outputs(2709) <= b;
    layer0_outputs(2710) <= a xor b;
    layer0_outputs(2711) <= not (a or b);
    layer0_outputs(2712) <= not a or b;
    layer0_outputs(2713) <= not (a xor b);
    layer0_outputs(2714) <= a or b;
    layer0_outputs(2715) <= not a;
    layer0_outputs(2716) <= not (a or b);
    layer0_outputs(2717) <= not b or a;
    layer0_outputs(2718) <= not b or a;
    layer0_outputs(2719) <= not (a and b);
    layer0_outputs(2720) <= not a or b;
    layer0_outputs(2721) <= not b;
    layer0_outputs(2722) <= a;
    layer0_outputs(2723) <= not (a or b);
    layer0_outputs(2724) <= b and not a;
    layer0_outputs(2725) <= not (a and b);
    layer0_outputs(2726) <= not b or a;
    layer0_outputs(2727) <= not b;
    layer0_outputs(2728) <= not (a xor b);
    layer0_outputs(2729) <= not b or a;
    layer0_outputs(2730) <= 1'b1;
    layer0_outputs(2731) <= a or b;
    layer0_outputs(2732) <= a xor b;
    layer0_outputs(2733) <= not (a or b);
    layer0_outputs(2734) <= b;
    layer0_outputs(2735) <= not b or a;
    layer0_outputs(2736) <= not (a or b);
    layer0_outputs(2737) <= a or b;
    layer0_outputs(2738) <= b;
    layer0_outputs(2739) <= b;
    layer0_outputs(2740) <= not b or a;
    layer0_outputs(2741) <= not b or a;
    layer0_outputs(2742) <= a or b;
    layer0_outputs(2743) <= b;
    layer0_outputs(2744) <= b;
    layer0_outputs(2745) <= a;
    layer0_outputs(2746) <= not (a or b);
    layer0_outputs(2747) <= not (a or b);
    layer0_outputs(2748) <= not (a xor b);
    layer0_outputs(2749) <= a and b;
    layer0_outputs(2750) <= a and b;
    layer0_outputs(2751) <= b and not a;
    layer0_outputs(2752) <= not (a or b);
    layer0_outputs(2753) <= not (a or b);
    layer0_outputs(2754) <= not b;
    layer0_outputs(2755) <= a and not b;
    layer0_outputs(2756) <= not a;
    layer0_outputs(2757) <= not (a or b);
    layer0_outputs(2758) <= not a;
    layer0_outputs(2759) <= not b or a;
    layer0_outputs(2760) <= not b or a;
    layer0_outputs(2761) <= not b;
    layer0_outputs(2762) <= not a;
    layer0_outputs(2763) <= b;
    layer0_outputs(2764) <= a xor b;
    layer0_outputs(2765) <= a;
    layer0_outputs(2766) <= not a or b;
    layer0_outputs(2767) <= not (a or b);
    layer0_outputs(2768) <= a and not b;
    layer0_outputs(2769) <= a;
    layer0_outputs(2770) <= a xor b;
    layer0_outputs(2771) <= 1'b1;
    layer0_outputs(2772) <= not a or b;
    layer0_outputs(2773) <= not (a xor b);
    layer0_outputs(2774) <= not a or b;
    layer0_outputs(2775) <= a xor b;
    layer0_outputs(2776) <= not a or b;
    layer0_outputs(2777) <= a and not b;
    layer0_outputs(2778) <= a;
    layer0_outputs(2779) <= a;
    layer0_outputs(2780) <= a xor b;
    layer0_outputs(2781) <= a xor b;
    layer0_outputs(2782) <= not (a xor b);
    layer0_outputs(2783) <= not (a or b);
    layer0_outputs(2784) <= a and b;
    layer0_outputs(2785) <= not b or a;
    layer0_outputs(2786) <= a and not b;
    layer0_outputs(2787) <= not b or a;
    layer0_outputs(2788) <= not a;
    layer0_outputs(2789) <= not a;
    layer0_outputs(2790) <= not (a or b);
    layer0_outputs(2791) <= 1'b0;
    layer0_outputs(2792) <= 1'b0;
    layer0_outputs(2793) <= not a;
    layer0_outputs(2794) <= not b;
    layer0_outputs(2795) <= not (a or b);
    layer0_outputs(2796) <= a or b;
    layer0_outputs(2797) <= b and not a;
    layer0_outputs(2798) <= not a or b;
    layer0_outputs(2799) <= b and not a;
    layer0_outputs(2800) <= b and not a;
    layer0_outputs(2801) <= a;
    layer0_outputs(2802) <= not b;
    layer0_outputs(2803) <= not a;
    layer0_outputs(2804) <= not (a or b);
    layer0_outputs(2805) <= not (a xor b);
    layer0_outputs(2806) <= not (a or b);
    layer0_outputs(2807) <= a xor b;
    layer0_outputs(2808) <= not (a xor b);
    layer0_outputs(2809) <= not (a and b);
    layer0_outputs(2810) <= a or b;
    layer0_outputs(2811) <= a and b;
    layer0_outputs(2812) <= 1'b1;
    layer0_outputs(2813) <= a xor b;
    layer0_outputs(2814) <= a or b;
    layer0_outputs(2815) <= b;
    layer0_outputs(2816) <= a and not b;
    layer0_outputs(2817) <= not b or a;
    layer0_outputs(2818) <= 1'b1;
    layer0_outputs(2819) <= not (a xor b);
    layer0_outputs(2820) <= a xor b;
    layer0_outputs(2821) <= a xor b;
    layer0_outputs(2822) <= not a;
    layer0_outputs(2823) <= not (a xor b);
    layer0_outputs(2824) <= not (a and b);
    layer0_outputs(2825) <= b and not a;
    layer0_outputs(2826) <= not a;
    layer0_outputs(2827) <= b;
    layer0_outputs(2828) <= 1'b1;
    layer0_outputs(2829) <= not a or b;
    layer0_outputs(2830) <= a and not b;
    layer0_outputs(2831) <= b;
    layer0_outputs(2832) <= b;
    layer0_outputs(2833) <= not b;
    layer0_outputs(2834) <= a and not b;
    layer0_outputs(2835) <= b and not a;
    layer0_outputs(2836) <= a xor b;
    layer0_outputs(2837) <= not b;
    layer0_outputs(2838) <= b;
    layer0_outputs(2839) <= not b or a;
    layer0_outputs(2840) <= a or b;
    layer0_outputs(2841) <= a and b;
    layer0_outputs(2842) <= not (a or b);
    layer0_outputs(2843) <= not (a xor b);
    layer0_outputs(2844) <= a;
    layer0_outputs(2845) <= a and b;
    layer0_outputs(2846) <= not (a xor b);
    layer0_outputs(2847) <= not (a xor b);
    layer0_outputs(2848) <= not (a and b);
    layer0_outputs(2849) <= not (a or b);
    layer0_outputs(2850) <= a;
    layer0_outputs(2851) <= a;
    layer0_outputs(2852) <= not b;
    layer0_outputs(2853) <= 1'b0;
    layer0_outputs(2854) <= a and b;
    layer0_outputs(2855) <= 1'b1;
    layer0_outputs(2856) <= a;
    layer0_outputs(2857) <= a or b;
    layer0_outputs(2858) <= not a;
    layer0_outputs(2859) <= not b;
    layer0_outputs(2860) <= 1'b0;
    layer0_outputs(2861) <= b;
    layer0_outputs(2862) <= not a or b;
    layer0_outputs(2863) <= a;
    layer0_outputs(2864) <= a xor b;
    layer0_outputs(2865) <= not (a or b);
    layer0_outputs(2866) <= b;
    layer0_outputs(2867) <= not (a xor b);
    layer0_outputs(2868) <= not b;
    layer0_outputs(2869) <= not a;
    layer0_outputs(2870) <= a or b;
    layer0_outputs(2871) <= not b;
    layer0_outputs(2872) <= a or b;
    layer0_outputs(2873) <= a and b;
    layer0_outputs(2874) <= b;
    layer0_outputs(2875) <= a and not b;
    layer0_outputs(2876) <= not (a or b);
    layer0_outputs(2877) <= a or b;
    layer0_outputs(2878) <= not (a xor b);
    layer0_outputs(2879) <= a;
    layer0_outputs(2880) <= b;
    layer0_outputs(2881) <= not (a xor b);
    layer0_outputs(2882) <= not a;
    layer0_outputs(2883) <= not (a or b);
    layer0_outputs(2884) <= a or b;
    layer0_outputs(2885) <= not (a or b);
    layer0_outputs(2886) <= 1'b1;
    layer0_outputs(2887) <= not (a or b);
    layer0_outputs(2888) <= a and not b;
    layer0_outputs(2889) <= b;
    layer0_outputs(2890) <= 1'b0;
    layer0_outputs(2891) <= not b or a;
    layer0_outputs(2892) <= b and not a;
    layer0_outputs(2893) <= 1'b1;
    layer0_outputs(2894) <= a and b;
    layer0_outputs(2895) <= not a or b;
    layer0_outputs(2896) <= not a or b;
    layer0_outputs(2897) <= not (a xor b);
    layer0_outputs(2898) <= not b or a;
    layer0_outputs(2899) <= a or b;
    layer0_outputs(2900) <= b;
    layer0_outputs(2901) <= not b or a;
    layer0_outputs(2902) <= b and not a;
    layer0_outputs(2903) <= a or b;
    layer0_outputs(2904) <= a or b;
    layer0_outputs(2905) <= a xor b;
    layer0_outputs(2906) <= b and not a;
    layer0_outputs(2907) <= b and not a;
    layer0_outputs(2908) <= not (a and b);
    layer0_outputs(2909) <= not b or a;
    layer0_outputs(2910) <= not (a or b);
    layer0_outputs(2911) <= 1'b1;
    layer0_outputs(2912) <= not b or a;
    layer0_outputs(2913) <= not (a xor b);
    layer0_outputs(2914) <= not a or b;
    layer0_outputs(2915) <= a;
    layer0_outputs(2916) <= not b;
    layer0_outputs(2917) <= b and not a;
    layer0_outputs(2918) <= not (a or b);
    layer0_outputs(2919) <= not a;
    layer0_outputs(2920) <= b and not a;
    layer0_outputs(2921) <= a or b;
    layer0_outputs(2922) <= not b;
    layer0_outputs(2923) <= not b;
    layer0_outputs(2924) <= a;
    layer0_outputs(2925) <= 1'b1;
    layer0_outputs(2926) <= not (a xor b);
    layer0_outputs(2927) <= not b;
    layer0_outputs(2928) <= b and not a;
    layer0_outputs(2929) <= 1'b1;
    layer0_outputs(2930) <= not a;
    layer0_outputs(2931) <= not b or a;
    layer0_outputs(2932) <= not b or a;
    layer0_outputs(2933) <= b and not a;
    layer0_outputs(2934) <= not (a or b);
    layer0_outputs(2935) <= not b or a;
    layer0_outputs(2936) <= a;
    layer0_outputs(2937) <= b and not a;
    layer0_outputs(2938) <= 1'b0;
    layer0_outputs(2939) <= not b;
    layer0_outputs(2940) <= a xor b;
    layer0_outputs(2941) <= 1'b0;
    layer0_outputs(2942) <= not (a xor b);
    layer0_outputs(2943) <= not a;
    layer0_outputs(2944) <= not a;
    layer0_outputs(2945) <= not a;
    layer0_outputs(2946) <= not (a or b);
    layer0_outputs(2947) <= not b;
    layer0_outputs(2948) <= a and not b;
    layer0_outputs(2949) <= a and not b;
    layer0_outputs(2950) <= b;
    layer0_outputs(2951) <= not b;
    layer0_outputs(2952) <= not b or a;
    layer0_outputs(2953) <= not (a or b);
    layer0_outputs(2954) <= 1'b0;
    layer0_outputs(2955) <= not a;
    layer0_outputs(2956) <= not a or b;
    layer0_outputs(2957) <= not (a xor b);
    layer0_outputs(2958) <= not a or b;
    layer0_outputs(2959) <= not a;
    layer0_outputs(2960) <= not (a xor b);
    layer0_outputs(2961) <= not (a xor b);
    layer0_outputs(2962) <= not b;
    layer0_outputs(2963) <= b;
    layer0_outputs(2964) <= a xor b;
    layer0_outputs(2965) <= not (a or b);
    layer0_outputs(2966) <= b and not a;
    layer0_outputs(2967) <= a xor b;
    layer0_outputs(2968) <= not b or a;
    layer0_outputs(2969) <= not (a xor b);
    layer0_outputs(2970) <= a;
    layer0_outputs(2971) <= b;
    layer0_outputs(2972) <= 1'b1;
    layer0_outputs(2973) <= a xor b;
    layer0_outputs(2974) <= not (a and b);
    layer0_outputs(2975) <= not b;
    layer0_outputs(2976) <= not b or a;
    layer0_outputs(2977) <= not a;
    layer0_outputs(2978) <= not (a or b);
    layer0_outputs(2979) <= b and not a;
    layer0_outputs(2980) <= a;
    layer0_outputs(2981) <= not (a xor b);
    layer0_outputs(2982) <= 1'b1;
    layer0_outputs(2983) <= not b;
    layer0_outputs(2984) <= b;
    layer0_outputs(2985) <= a or b;
    layer0_outputs(2986) <= a;
    layer0_outputs(2987) <= not b;
    layer0_outputs(2988) <= 1'b0;
    layer0_outputs(2989) <= 1'b0;
    layer0_outputs(2990) <= a xor b;
    layer0_outputs(2991) <= a or b;
    layer0_outputs(2992) <= not a or b;
    layer0_outputs(2993) <= b;
    layer0_outputs(2994) <= a;
    layer0_outputs(2995) <= b and not a;
    layer0_outputs(2996) <= not (a xor b);
    layer0_outputs(2997) <= b;
    layer0_outputs(2998) <= not b or a;
    layer0_outputs(2999) <= b and not a;
    layer0_outputs(3000) <= a;
    layer0_outputs(3001) <= not (a and b);
    layer0_outputs(3002) <= a and b;
    layer0_outputs(3003) <= a or b;
    layer0_outputs(3004) <= not (a or b);
    layer0_outputs(3005) <= a and not b;
    layer0_outputs(3006) <= not (a xor b);
    layer0_outputs(3007) <= a or b;
    layer0_outputs(3008) <= not b;
    layer0_outputs(3009) <= a xor b;
    layer0_outputs(3010) <= b and not a;
    layer0_outputs(3011) <= a and not b;
    layer0_outputs(3012) <= not (a or b);
    layer0_outputs(3013) <= not b or a;
    layer0_outputs(3014) <= b and not a;
    layer0_outputs(3015) <= not (a xor b);
    layer0_outputs(3016) <= a or b;
    layer0_outputs(3017) <= not b or a;
    layer0_outputs(3018) <= b and not a;
    layer0_outputs(3019) <= a and not b;
    layer0_outputs(3020) <= 1'b0;
    layer0_outputs(3021) <= 1'b1;
    layer0_outputs(3022) <= a xor b;
    layer0_outputs(3023) <= b and not a;
    layer0_outputs(3024) <= a or b;
    layer0_outputs(3025) <= a;
    layer0_outputs(3026) <= not b or a;
    layer0_outputs(3027) <= a xor b;
    layer0_outputs(3028) <= a and b;
    layer0_outputs(3029) <= b and not a;
    layer0_outputs(3030) <= not (a xor b);
    layer0_outputs(3031) <= a and b;
    layer0_outputs(3032) <= a and b;
    layer0_outputs(3033) <= not b or a;
    layer0_outputs(3034) <= not a or b;
    layer0_outputs(3035) <= 1'b1;
    layer0_outputs(3036) <= not (a or b);
    layer0_outputs(3037) <= a and not b;
    layer0_outputs(3038) <= not (a or b);
    layer0_outputs(3039) <= not a;
    layer0_outputs(3040) <= a and b;
    layer0_outputs(3041) <= a;
    layer0_outputs(3042) <= a;
    layer0_outputs(3043) <= not a;
    layer0_outputs(3044) <= a and b;
    layer0_outputs(3045) <= a xor b;
    layer0_outputs(3046) <= not b;
    layer0_outputs(3047) <= not (a or b);
    layer0_outputs(3048) <= 1'b1;
    layer0_outputs(3049) <= not (a xor b);
    layer0_outputs(3050) <= b;
    layer0_outputs(3051) <= a and not b;
    layer0_outputs(3052) <= a or b;
    layer0_outputs(3053) <= not (a or b);
    layer0_outputs(3054) <= a or b;
    layer0_outputs(3055) <= a xor b;
    layer0_outputs(3056) <= a or b;
    layer0_outputs(3057) <= not b;
    layer0_outputs(3058) <= b;
    layer0_outputs(3059) <= not b;
    layer0_outputs(3060) <= not (a or b);
    layer0_outputs(3061) <= not (a xor b);
    layer0_outputs(3062) <= a and not b;
    layer0_outputs(3063) <= b and not a;
    layer0_outputs(3064) <= a and not b;
    layer0_outputs(3065) <= a or b;
    layer0_outputs(3066) <= not a;
    layer0_outputs(3067) <= a and not b;
    layer0_outputs(3068) <= a and not b;
    layer0_outputs(3069) <= not b;
    layer0_outputs(3070) <= not (a or b);
    layer0_outputs(3071) <= not a or b;
    layer0_outputs(3072) <= a and b;
    layer0_outputs(3073) <= not (a xor b);
    layer0_outputs(3074) <= not b or a;
    layer0_outputs(3075) <= not (a xor b);
    layer0_outputs(3076) <= not a or b;
    layer0_outputs(3077) <= a;
    layer0_outputs(3078) <= not (a or b);
    layer0_outputs(3079) <= a;
    layer0_outputs(3080) <= not b;
    layer0_outputs(3081) <= a and not b;
    layer0_outputs(3082) <= b and not a;
    layer0_outputs(3083) <= not a;
    layer0_outputs(3084) <= b;
    layer0_outputs(3085) <= a;
    layer0_outputs(3086) <= not b or a;
    layer0_outputs(3087) <= a or b;
    layer0_outputs(3088) <= a;
    layer0_outputs(3089) <= 1'b0;
    layer0_outputs(3090) <= 1'b1;
    layer0_outputs(3091) <= not a or b;
    layer0_outputs(3092) <= 1'b0;
    layer0_outputs(3093) <= a and not b;
    layer0_outputs(3094) <= a;
    layer0_outputs(3095) <= not a;
    layer0_outputs(3096) <= not b;
    layer0_outputs(3097) <= 1'b0;
    layer0_outputs(3098) <= a;
    layer0_outputs(3099) <= not (a and b);
    layer0_outputs(3100) <= not (a or b);
    layer0_outputs(3101) <= b and not a;
    layer0_outputs(3102) <= 1'b0;
    layer0_outputs(3103) <= a xor b;
    layer0_outputs(3104) <= not (a xor b);
    layer0_outputs(3105) <= a xor b;
    layer0_outputs(3106) <= not (a xor b);
    layer0_outputs(3107) <= a or b;
    layer0_outputs(3108) <= a xor b;
    layer0_outputs(3109) <= not a;
    layer0_outputs(3110) <= a or b;
    layer0_outputs(3111) <= a;
    layer0_outputs(3112) <= a;
    layer0_outputs(3113) <= a and b;
    layer0_outputs(3114) <= not a;
    layer0_outputs(3115) <= b;
    layer0_outputs(3116) <= not b;
    layer0_outputs(3117) <= a or b;
    layer0_outputs(3118) <= not b;
    layer0_outputs(3119) <= a and not b;
    layer0_outputs(3120) <= not a or b;
    layer0_outputs(3121) <= not (a xor b);
    layer0_outputs(3122) <= a or b;
    layer0_outputs(3123) <= not b or a;
    layer0_outputs(3124) <= b;
    layer0_outputs(3125) <= a;
    layer0_outputs(3126) <= a or b;
    layer0_outputs(3127) <= b;
    layer0_outputs(3128) <= not b or a;
    layer0_outputs(3129) <= b;
    layer0_outputs(3130) <= not b;
    layer0_outputs(3131) <= a and not b;
    layer0_outputs(3132) <= a or b;
    layer0_outputs(3133) <= a or b;
    layer0_outputs(3134) <= a and not b;
    layer0_outputs(3135) <= a or b;
    layer0_outputs(3136) <= not (a or b);
    layer0_outputs(3137) <= not b;
    layer0_outputs(3138) <= a or b;
    layer0_outputs(3139) <= a;
    layer0_outputs(3140) <= a or b;
    layer0_outputs(3141) <= b and not a;
    layer0_outputs(3142) <= not (a or b);
    layer0_outputs(3143) <= a;
    layer0_outputs(3144) <= a;
    layer0_outputs(3145) <= b;
    layer0_outputs(3146) <= a and b;
    layer0_outputs(3147) <= b and not a;
    layer0_outputs(3148) <= not a or b;
    layer0_outputs(3149) <= not b;
    layer0_outputs(3150) <= a;
    layer0_outputs(3151) <= b and not a;
    layer0_outputs(3152) <= not b or a;
    layer0_outputs(3153) <= a and not b;
    layer0_outputs(3154) <= a xor b;
    layer0_outputs(3155) <= not b;
    layer0_outputs(3156) <= not a;
    layer0_outputs(3157) <= a or b;
    layer0_outputs(3158) <= a xor b;
    layer0_outputs(3159) <= 1'b1;
    layer0_outputs(3160) <= not a or b;
    layer0_outputs(3161) <= not (a or b);
    layer0_outputs(3162) <= b and not a;
    layer0_outputs(3163) <= not (a and b);
    layer0_outputs(3164) <= b and not a;
    layer0_outputs(3165) <= a and not b;
    layer0_outputs(3166) <= not a or b;
    layer0_outputs(3167) <= a or b;
    layer0_outputs(3168) <= not (a or b);
    layer0_outputs(3169) <= not (a or b);
    layer0_outputs(3170) <= not b;
    layer0_outputs(3171) <= not b;
    layer0_outputs(3172) <= not b;
    layer0_outputs(3173) <= not b or a;
    layer0_outputs(3174) <= not a;
    layer0_outputs(3175) <= a or b;
    layer0_outputs(3176) <= not (a or b);
    layer0_outputs(3177) <= not a;
    layer0_outputs(3178) <= a xor b;
    layer0_outputs(3179) <= b and not a;
    layer0_outputs(3180) <= a and b;
    layer0_outputs(3181) <= not (a xor b);
    layer0_outputs(3182) <= a xor b;
    layer0_outputs(3183) <= a or b;
    layer0_outputs(3184) <= b;
    layer0_outputs(3185) <= not (a or b);
    layer0_outputs(3186) <= b and not a;
    layer0_outputs(3187) <= not (a or b);
    layer0_outputs(3188) <= a and not b;
    layer0_outputs(3189) <= not a or b;
    layer0_outputs(3190) <= 1'b0;
    layer0_outputs(3191) <= 1'b0;
    layer0_outputs(3192) <= b;
    layer0_outputs(3193) <= not (a xor b);
    layer0_outputs(3194) <= b;
    layer0_outputs(3195) <= a and not b;
    layer0_outputs(3196) <= a and not b;
    layer0_outputs(3197) <= not (a xor b);
    layer0_outputs(3198) <= a xor b;
    layer0_outputs(3199) <= a and b;
    layer0_outputs(3200) <= not b or a;
    layer0_outputs(3201) <= not (a or b);
    layer0_outputs(3202) <= b and not a;
    layer0_outputs(3203) <= not (a and b);
    layer0_outputs(3204) <= a;
    layer0_outputs(3205) <= not (a or b);
    layer0_outputs(3206) <= not b;
    layer0_outputs(3207) <= not (a or b);
    layer0_outputs(3208) <= a or b;
    layer0_outputs(3209) <= not b;
    layer0_outputs(3210) <= a or b;
    layer0_outputs(3211) <= a and b;
    layer0_outputs(3212) <= not a;
    layer0_outputs(3213) <= 1'b1;
    layer0_outputs(3214) <= b and not a;
    layer0_outputs(3215) <= not b;
    layer0_outputs(3216) <= a and not b;
    layer0_outputs(3217) <= not (a or b);
    layer0_outputs(3218) <= a xor b;
    layer0_outputs(3219) <= a or b;
    layer0_outputs(3220) <= not a or b;
    layer0_outputs(3221) <= a xor b;
    layer0_outputs(3222) <= not a or b;
    layer0_outputs(3223) <= b;
    layer0_outputs(3224) <= not b or a;
    layer0_outputs(3225) <= b;
    layer0_outputs(3226) <= not b;
    layer0_outputs(3227) <= a xor b;
    layer0_outputs(3228) <= a xor b;
    layer0_outputs(3229) <= a or b;
    layer0_outputs(3230) <= a or b;
    layer0_outputs(3231) <= a;
    layer0_outputs(3232) <= a or b;
    layer0_outputs(3233) <= not (a and b);
    layer0_outputs(3234) <= a or b;
    layer0_outputs(3235) <= a and not b;
    layer0_outputs(3236) <= a xor b;
    layer0_outputs(3237) <= a xor b;
    layer0_outputs(3238) <= a;
    layer0_outputs(3239) <= b;
    layer0_outputs(3240) <= not a or b;
    layer0_outputs(3241) <= not (a and b);
    layer0_outputs(3242) <= a;
    layer0_outputs(3243) <= not b;
    layer0_outputs(3244) <= not b;
    layer0_outputs(3245) <= a or b;
    layer0_outputs(3246) <= a and not b;
    layer0_outputs(3247) <= a xor b;
    layer0_outputs(3248) <= not b or a;
    layer0_outputs(3249) <= b and not a;
    layer0_outputs(3250) <= a or b;
    layer0_outputs(3251) <= not (a or b);
    layer0_outputs(3252) <= a xor b;
    layer0_outputs(3253) <= a or b;
    layer0_outputs(3254) <= a;
    layer0_outputs(3255) <= a xor b;
    layer0_outputs(3256) <= not a or b;
    layer0_outputs(3257) <= b and not a;
    layer0_outputs(3258) <= 1'b0;
    layer0_outputs(3259) <= not a or b;
    layer0_outputs(3260) <= a or b;
    layer0_outputs(3261) <= a;
    layer0_outputs(3262) <= a or b;
    layer0_outputs(3263) <= a xor b;
    layer0_outputs(3264) <= a and b;
    layer0_outputs(3265) <= not b;
    layer0_outputs(3266) <= not (a xor b);
    layer0_outputs(3267) <= not b or a;
    layer0_outputs(3268) <= a and not b;
    layer0_outputs(3269) <= not b;
    layer0_outputs(3270) <= not a;
    layer0_outputs(3271) <= not b or a;
    layer0_outputs(3272) <= 1'b0;
    layer0_outputs(3273) <= not (a xor b);
    layer0_outputs(3274) <= a and not b;
    layer0_outputs(3275) <= b;
    layer0_outputs(3276) <= not b or a;
    layer0_outputs(3277) <= a;
    layer0_outputs(3278) <= b and not a;
    layer0_outputs(3279) <= not b;
    layer0_outputs(3280) <= a and not b;
    layer0_outputs(3281) <= a and not b;
    layer0_outputs(3282) <= not (a xor b);
    layer0_outputs(3283) <= 1'b0;
    layer0_outputs(3284) <= not a;
    layer0_outputs(3285) <= a;
    layer0_outputs(3286) <= a or b;
    layer0_outputs(3287) <= b;
    layer0_outputs(3288) <= a or b;
    layer0_outputs(3289) <= a or b;
    layer0_outputs(3290) <= not a or b;
    layer0_outputs(3291) <= a and not b;
    layer0_outputs(3292) <= a;
    layer0_outputs(3293) <= not (a and b);
    layer0_outputs(3294) <= not (a xor b);
    layer0_outputs(3295) <= not (a or b);
    layer0_outputs(3296) <= not (a xor b);
    layer0_outputs(3297) <= a and not b;
    layer0_outputs(3298) <= a or b;
    layer0_outputs(3299) <= a and not b;
    layer0_outputs(3300) <= a and not b;
    layer0_outputs(3301) <= not (a or b);
    layer0_outputs(3302) <= not a;
    layer0_outputs(3303) <= not (a or b);
    layer0_outputs(3304) <= a xor b;
    layer0_outputs(3305) <= not (a or b);
    layer0_outputs(3306) <= b;
    layer0_outputs(3307) <= not b;
    layer0_outputs(3308) <= b;
    layer0_outputs(3309) <= not a;
    layer0_outputs(3310) <= a or b;
    layer0_outputs(3311) <= b;
    layer0_outputs(3312) <= a and not b;
    layer0_outputs(3313) <= not b;
    layer0_outputs(3314) <= not a;
    layer0_outputs(3315) <= a xor b;
    layer0_outputs(3316) <= a xor b;
    layer0_outputs(3317) <= not (a and b);
    layer0_outputs(3318) <= not b;
    layer0_outputs(3319) <= not b;
    layer0_outputs(3320) <= 1'b1;
    layer0_outputs(3321) <= not (a xor b);
    layer0_outputs(3322) <= not (a xor b);
    layer0_outputs(3323) <= not a;
    layer0_outputs(3324) <= a and not b;
    layer0_outputs(3325) <= not a or b;
    layer0_outputs(3326) <= a;
    layer0_outputs(3327) <= a;
    layer0_outputs(3328) <= a or b;
    layer0_outputs(3329) <= not (a or b);
    layer0_outputs(3330) <= not (a or b);
    layer0_outputs(3331) <= b;
    layer0_outputs(3332) <= not a or b;
    layer0_outputs(3333) <= not b or a;
    layer0_outputs(3334) <= a and b;
    layer0_outputs(3335) <= 1'b1;
    layer0_outputs(3336) <= not a or b;
    layer0_outputs(3337) <= a;
    layer0_outputs(3338) <= not (a or b);
    layer0_outputs(3339) <= a and b;
    layer0_outputs(3340) <= b;
    layer0_outputs(3341) <= not a;
    layer0_outputs(3342) <= not a;
    layer0_outputs(3343) <= b and not a;
    layer0_outputs(3344) <= a or b;
    layer0_outputs(3345) <= not b;
    layer0_outputs(3346) <= a or b;
    layer0_outputs(3347) <= a xor b;
    layer0_outputs(3348) <= not b;
    layer0_outputs(3349) <= 1'b1;
    layer0_outputs(3350) <= a or b;
    layer0_outputs(3351) <= not b;
    layer0_outputs(3352) <= b;
    layer0_outputs(3353) <= not b or a;
    layer0_outputs(3354) <= not (a xor b);
    layer0_outputs(3355) <= a;
    layer0_outputs(3356) <= not (a and b);
    layer0_outputs(3357) <= not a;
    layer0_outputs(3358) <= 1'b1;
    layer0_outputs(3359) <= a and b;
    layer0_outputs(3360) <= not a;
    layer0_outputs(3361) <= not (a xor b);
    layer0_outputs(3362) <= not b;
    layer0_outputs(3363) <= not a;
    layer0_outputs(3364) <= 1'b1;
    layer0_outputs(3365) <= a;
    layer0_outputs(3366) <= a or b;
    layer0_outputs(3367) <= not (a or b);
    layer0_outputs(3368) <= not (a xor b);
    layer0_outputs(3369) <= not b;
    layer0_outputs(3370) <= b and not a;
    layer0_outputs(3371) <= not b or a;
    layer0_outputs(3372) <= b and not a;
    layer0_outputs(3373) <= not b;
    layer0_outputs(3374) <= not b or a;
    layer0_outputs(3375) <= not a;
    layer0_outputs(3376) <= a xor b;
    layer0_outputs(3377) <= b;
    layer0_outputs(3378) <= not (a and b);
    layer0_outputs(3379) <= a;
    layer0_outputs(3380) <= a and not b;
    layer0_outputs(3381) <= a and b;
    layer0_outputs(3382) <= a;
    layer0_outputs(3383) <= not b or a;
    layer0_outputs(3384) <= not (a xor b);
    layer0_outputs(3385) <= 1'b1;
    layer0_outputs(3386) <= not (a or b);
    layer0_outputs(3387) <= a;
    layer0_outputs(3388) <= b and not a;
    layer0_outputs(3389) <= a or b;
    layer0_outputs(3390) <= b and not a;
    layer0_outputs(3391) <= b;
    layer0_outputs(3392) <= not (a or b);
    layer0_outputs(3393) <= not (a xor b);
    layer0_outputs(3394) <= a xor b;
    layer0_outputs(3395) <= a or b;
    layer0_outputs(3396) <= not a or b;
    layer0_outputs(3397) <= a or b;
    layer0_outputs(3398) <= b and not a;
    layer0_outputs(3399) <= 1'b0;
    layer0_outputs(3400) <= 1'b1;
    layer0_outputs(3401) <= a and not b;
    layer0_outputs(3402) <= a or b;
    layer0_outputs(3403) <= b;
    layer0_outputs(3404) <= 1'b1;
    layer0_outputs(3405) <= not (a or b);
    layer0_outputs(3406) <= a;
    layer0_outputs(3407) <= not (a xor b);
    layer0_outputs(3408) <= not (a and b);
    layer0_outputs(3409) <= not b;
    layer0_outputs(3410) <= not a or b;
    layer0_outputs(3411) <= not (a xor b);
    layer0_outputs(3412) <= not (a or b);
    layer0_outputs(3413) <= a;
    layer0_outputs(3414) <= a and not b;
    layer0_outputs(3415) <= a or b;
    layer0_outputs(3416) <= a or b;
    layer0_outputs(3417) <= not a or b;
    layer0_outputs(3418) <= 1'b1;
    layer0_outputs(3419) <= not a or b;
    layer0_outputs(3420) <= not (a xor b);
    layer0_outputs(3421) <= not a;
    layer0_outputs(3422) <= b and not a;
    layer0_outputs(3423) <= b;
    layer0_outputs(3424) <= not a;
    layer0_outputs(3425) <= not b;
    layer0_outputs(3426) <= not (a and b);
    layer0_outputs(3427) <= not a or b;
    layer0_outputs(3428) <= a xor b;
    layer0_outputs(3429) <= not b;
    layer0_outputs(3430) <= not b or a;
    layer0_outputs(3431) <= not a or b;
    layer0_outputs(3432) <= a or b;
    layer0_outputs(3433) <= not a;
    layer0_outputs(3434) <= a;
    layer0_outputs(3435) <= not b;
    layer0_outputs(3436) <= a xor b;
    layer0_outputs(3437) <= a;
    layer0_outputs(3438) <= 1'b0;
    layer0_outputs(3439) <= not a;
    layer0_outputs(3440) <= not a;
    layer0_outputs(3441) <= a and not b;
    layer0_outputs(3442) <= b and not a;
    layer0_outputs(3443) <= b and not a;
    layer0_outputs(3444) <= a and not b;
    layer0_outputs(3445) <= not a or b;
    layer0_outputs(3446) <= not b;
    layer0_outputs(3447) <= b;
    layer0_outputs(3448) <= not a;
    layer0_outputs(3449) <= not a;
    layer0_outputs(3450) <= b;
    layer0_outputs(3451) <= not a;
    layer0_outputs(3452) <= not b;
    layer0_outputs(3453) <= not (a xor b);
    layer0_outputs(3454) <= a or b;
    layer0_outputs(3455) <= a and b;
    layer0_outputs(3456) <= not b;
    layer0_outputs(3457) <= b;
    layer0_outputs(3458) <= not a or b;
    layer0_outputs(3459) <= b and not a;
    layer0_outputs(3460) <= a or b;
    layer0_outputs(3461) <= 1'b1;
    layer0_outputs(3462) <= not (a and b);
    layer0_outputs(3463) <= b;
    layer0_outputs(3464) <= b;
    layer0_outputs(3465) <= b;
    layer0_outputs(3466) <= not b;
    layer0_outputs(3467) <= a xor b;
    layer0_outputs(3468) <= a;
    layer0_outputs(3469) <= a or b;
    layer0_outputs(3470) <= not b;
    layer0_outputs(3471) <= a or b;
    layer0_outputs(3472) <= a;
    layer0_outputs(3473) <= a xor b;
    layer0_outputs(3474) <= a xor b;
    layer0_outputs(3475) <= not b;
    layer0_outputs(3476) <= not (a xor b);
    layer0_outputs(3477) <= not b;
    layer0_outputs(3478) <= a xor b;
    layer0_outputs(3479) <= 1'b1;
    layer0_outputs(3480) <= not (a and b);
    layer0_outputs(3481) <= b;
    layer0_outputs(3482) <= not a;
    layer0_outputs(3483) <= a and not b;
    layer0_outputs(3484) <= not b;
    layer0_outputs(3485) <= not a;
    layer0_outputs(3486) <= a;
    layer0_outputs(3487) <= a xor b;
    layer0_outputs(3488) <= not b or a;
    layer0_outputs(3489) <= not a;
    layer0_outputs(3490) <= a or b;
    layer0_outputs(3491) <= 1'b1;
    layer0_outputs(3492) <= not a;
    layer0_outputs(3493) <= not b or a;
    layer0_outputs(3494) <= not (a and b);
    layer0_outputs(3495) <= 1'b0;
    layer0_outputs(3496) <= not b or a;
    layer0_outputs(3497) <= a or b;
    layer0_outputs(3498) <= not b or a;
    layer0_outputs(3499) <= not a;
    layer0_outputs(3500) <= a or b;
    layer0_outputs(3501) <= 1'b1;
    layer0_outputs(3502) <= not b or a;
    layer0_outputs(3503) <= not b or a;
    layer0_outputs(3504) <= not (a and b);
    layer0_outputs(3505) <= not a;
    layer0_outputs(3506) <= b;
    layer0_outputs(3507) <= not b;
    layer0_outputs(3508) <= a and b;
    layer0_outputs(3509) <= b and not a;
    layer0_outputs(3510) <= a and not b;
    layer0_outputs(3511) <= a and not b;
    layer0_outputs(3512) <= a or b;
    layer0_outputs(3513) <= not b;
    layer0_outputs(3514) <= a;
    layer0_outputs(3515) <= not b or a;
    layer0_outputs(3516) <= not b;
    layer0_outputs(3517) <= not a;
    layer0_outputs(3518) <= a;
    layer0_outputs(3519) <= not b or a;
    layer0_outputs(3520) <= not (a or b);
    layer0_outputs(3521) <= 1'b1;
    layer0_outputs(3522) <= not (a or b);
    layer0_outputs(3523) <= a and not b;
    layer0_outputs(3524) <= 1'b0;
    layer0_outputs(3525) <= 1'b0;
    layer0_outputs(3526) <= not a or b;
    layer0_outputs(3527) <= a or b;
    layer0_outputs(3528) <= a or b;
    layer0_outputs(3529) <= not (a or b);
    layer0_outputs(3530) <= not (a and b);
    layer0_outputs(3531) <= a or b;
    layer0_outputs(3532) <= not b;
    layer0_outputs(3533) <= a and b;
    layer0_outputs(3534) <= a xor b;
    layer0_outputs(3535) <= b;
    layer0_outputs(3536) <= a xor b;
    layer0_outputs(3537) <= a and b;
    layer0_outputs(3538) <= not (a xor b);
    layer0_outputs(3539) <= a and b;
    layer0_outputs(3540) <= a;
    layer0_outputs(3541) <= not (a or b);
    layer0_outputs(3542) <= not a;
    layer0_outputs(3543) <= not (a or b);
    layer0_outputs(3544) <= a xor b;
    layer0_outputs(3545) <= 1'b0;
    layer0_outputs(3546) <= not b;
    layer0_outputs(3547) <= not (a or b);
    layer0_outputs(3548) <= not (a or b);
    layer0_outputs(3549) <= not a;
    layer0_outputs(3550) <= a xor b;
    layer0_outputs(3551) <= not (a or b);
    layer0_outputs(3552) <= a xor b;
    layer0_outputs(3553) <= not (a or b);
    layer0_outputs(3554) <= not a or b;
    layer0_outputs(3555) <= not b;
    layer0_outputs(3556) <= 1'b0;
    layer0_outputs(3557) <= b and not a;
    layer0_outputs(3558) <= not b or a;
    layer0_outputs(3559) <= not (a xor b);
    layer0_outputs(3560) <= not (a xor b);
    layer0_outputs(3561) <= not (a or b);
    layer0_outputs(3562) <= a;
    layer0_outputs(3563) <= not b;
    layer0_outputs(3564) <= 1'b1;
    layer0_outputs(3565) <= a and not b;
    layer0_outputs(3566) <= 1'b1;
    layer0_outputs(3567) <= not b;
    layer0_outputs(3568) <= 1'b0;
    layer0_outputs(3569) <= a or b;
    layer0_outputs(3570) <= not (a xor b);
    layer0_outputs(3571) <= not b;
    layer0_outputs(3572) <= not (a or b);
    layer0_outputs(3573) <= not b or a;
    layer0_outputs(3574) <= b and not a;
    layer0_outputs(3575) <= not (a or b);
    layer0_outputs(3576) <= not a;
    layer0_outputs(3577) <= not b or a;
    layer0_outputs(3578) <= a or b;
    layer0_outputs(3579) <= not (a and b);
    layer0_outputs(3580) <= b and not a;
    layer0_outputs(3581) <= a and not b;
    layer0_outputs(3582) <= b and not a;
    layer0_outputs(3583) <= not (a or b);
    layer0_outputs(3584) <= not a or b;
    layer0_outputs(3585) <= a xor b;
    layer0_outputs(3586) <= not b;
    layer0_outputs(3587) <= a or b;
    layer0_outputs(3588) <= not a;
    layer0_outputs(3589) <= not (a or b);
    layer0_outputs(3590) <= a and not b;
    layer0_outputs(3591) <= b and not a;
    layer0_outputs(3592) <= a or b;
    layer0_outputs(3593) <= a xor b;
    layer0_outputs(3594) <= not (a xor b);
    layer0_outputs(3595) <= not (a and b);
    layer0_outputs(3596) <= not b or a;
    layer0_outputs(3597) <= b and not a;
    layer0_outputs(3598) <= 1'b1;
    layer0_outputs(3599) <= not (a and b);
    layer0_outputs(3600) <= b and not a;
    layer0_outputs(3601) <= not (a or b);
    layer0_outputs(3602) <= not b;
    layer0_outputs(3603) <= a and not b;
    layer0_outputs(3604) <= not (a or b);
    layer0_outputs(3605) <= b and not a;
    layer0_outputs(3606) <= a xor b;
    layer0_outputs(3607) <= a or b;
    layer0_outputs(3608) <= 1'b0;
    layer0_outputs(3609) <= not a;
    layer0_outputs(3610) <= a xor b;
    layer0_outputs(3611) <= a xor b;
    layer0_outputs(3612) <= b and not a;
    layer0_outputs(3613) <= a or b;
    layer0_outputs(3614) <= a or b;
    layer0_outputs(3615) <= a xor b;
    layer0_outputs(3616) <= not b;
    layer0_outputs(3617) <= a or b;
    layer0_outputs(3618) <= a and b;
    layer0_outputs(3619) <= not b;
    layer0_outputs(3620) <= not (a or b);
    layer0_outputs(3621) <= b;
    layer0_outputs(3622) <= not (a xor b);
    layer0_outputs(3623) <= not (a or b);
    layer0_outputs(3624) <= b;
    layer0_outputs(3625) <= not b or a;
    layer0_outputs(3626) <= a;
    layer0_outputs(3627) <= not b;
    layer0_outputs(3628) <= a;
    layer0_outputs(3629) <= a and not b;
    layer0_outputs(3630) <= b and not a;
    layer0_outputs(3631) <= a xor b;
    layer0_outputs(3632) <= not (a xor b);
    layer0_outputs(3633) <= a or b;
    layer0_outputs(3634) <= b;
    layer0_outputs(3635) <= 1'b1;
    layer0_outputs(3636) <= b and not a;
    layer0_outputs(3637) <= not b or a;
    layer0_outputs(3638) <= not b or a;
    layer0_outputs(3639) <= a or b;
    layer0_outputs(3640) <= b;
    layer0_outputs(3641) <= 1'b0;
    layer0_outputs(3642) <= not b or a;
    layer0_outputs(3643) <= a or b;
    layer0_outputs(3644) <= not a;
    layer0_outputs(3645) <= a xor b;
    layer0_outputs(3646) <= a;
    layer0_outputs(3647) <= a;
    layer0_outputs(3648) <= a and b;
    layer0_outputs(3649) <= 1'b0;
    layer0_outputs(3650) <= a or b;
    layer0_outputs(3651) <= a and b;
    layer0_outputs(3652) <= not a;
    layer0_outputs(3653) <= a xor b;
    layer0_outputs(3654) <= a xor b;
    layer0_outputs(3655) <= a xor b;
    layer0_outputs(3656) <= a;
    layer0_outputs(3657) <= not a or b;
    layer0_outputs(3658) <= a xor b;
    layer0_outputs(3659) <= not (a xor b);
    layer0_outputs(3660) <= not (a xor b);
    layer0_outputs(3661) <= b and not a;
    layer0_outputs(3662) <= not a;
    layer0_outputs(3663) <= not b;
    layer0_outputs(3664) <= 1'b1;
    layer0_outputs(3665) <= not a or b;
    layer0_outputs(3666) <= a or b;
    layer0_outputs(3667) <= not (a xor b);
    layer0_outputs(3668) <= not b or a;
    layer0_outputs(3669) <= b;
    layer0_outputs(3670) <= not a;
    layer0_outputs(3671) <= b;
    layer0_outputs(3672) <= b and not a;
    layer0_outputs(3673) <= a and b;
    layer0_outputs(3674) <= not b;
    layer0_outputs(3675) <= not (a or b);
    layer0_outputs(3676) <= not a;
    layer0_outputs(3677) <= not b;
    layer0_outputs(3678) <= b and not a;
    layer0_outputs(3679) <= 1'b0;
    layer0_outputs(3680) <= b;
    layer0_outputs(3681) <= 1'b1;
    layer0_outputs(3682) <= b and not a;
    layer0_outputs(3683) <= not b;
    layer0_outputs(3684) <= b;
    layer0_outputs(3685) <= not (a and b);
    layer0_outputs(3686) <= not (a or b);
    layer0_outputs(3687) <= a;
    layer0_outputs(3688) <= a;
    layer0_outputs(3689) <= not b;
    layer0_outputs(3690) <= a;
    layer0_outputs(3691) <= not b or a;
    layer0_outputs(3692) <= not b;
    layer0_outputs(3693) <= not a;
    layer0_outputs(3694) <= not a;
    layer0_outputs(3695) <= a or b;
    layer0_outputs(3696) <= not (a or b);
    layer0_outputs(3697) <= 1'b0;
    layer0_outputs(3698) <= not (a or b);
    layer0_outputs(3699) <= not (a xor b);
    layer0_outputs(3700) <= 1'b0;
    layer0_outputs(3701) <= not b or a;
    layer0_outputs(3702) <= not a or b;
    layer0_outputs(3703) <= a xor b;
    layer0_outputs(3704) <= not (a xor b);
    layer0_outputs(3705) <= not (a xor b);
    layer0_outputs(3706) <= a or b;
    layer0_outputs(3707) <= b and not a;
    layer0_outputs(3708) <= a and b;
    layer0_outputs(3709) <= not b;
    layer0_outputs(3710) <= not a;
    layer0_outputs(3711) <= 1'b0;
    layer0_outputs(3712) <= not (a or b);
    layer0_outputs(3713) <= 1'b1;
    layer0_outputs(3714) <= a;
    layer0_outputs(3715) <= not (a or b);
    layer0_outputs(3716) <= not (a and b);
    layer0_outputs(3717) <= a;
    layer0_outputs(3718) <= not a;
    layer0_outputs(3719) <= not b;
    layer0_outputs(3720) <= a or b;
    layer0_outputs(3721) <= b;
    layer0_outputs(3722) <= a xor b;
    layer0_outputs(3723) <= b;
    layer0_outputs(3724) <= b and not a;
    layer0_outputs(3725) <= a;
    layer0_outputs(3726) <= not b;
    layer0_outputs(3727) <= not (a xor b);
    layer0_outputs(3728) <= not b;
    layer0_outputs(3729) <= 1'b1;
    layer0_outputs(3730) <= a xor b;
    layer0_outputs(3731) <= not (a xor b);
    layer0_outputs(3732) <= a;
    layer0_outputs(3733) <= b;
    layer0_outputs(3734) <= not b;
    layer0_outputs(3735) <= not b or a;
    layer0_outputs(3736) <= not b or a;
    layer0_outputs(3737) <= a and not b;
    layer0_outputs(3738) <= a xor b;
    layer0_outputs(3739) <= a xor b;
    layer0_outputs(3740) <= not a or b;
    layer0_outputs(3741) <= a and not b;
    layer0_outputs(3742) <= a or b;
    layer0_outputs(3743) <= not b;
    layer0_outputs(3744) <= a;
    layer0_outputs(3745) <= not a;
    layer0_outputs(3746) <= a or b;
    layer0_outputs(3747) <= a or b;
    layer0_outputs(3748) <= not (a or b);
    layer0_outputs(3749) <= not a or b;
    layer0_outputs(3750) <= b;
    layer0_outputs(3751) <= a or b;
    layer0_outputs(3752) <= b;
    layer0_outputs(3753) <= 1'b0;
    layer0_outputs(3754) <= a;
    layer0_outputs(3755) <= b;
    layer0_outputs(3756) <= not a or b;
    layer0_outputs(3757) <= 1'b0;
    layer0_outputs(3758) <= a;
    layer0_outputs(3759) <= a and b;
    layer0_outputs(3760) <= not (a or b);
    layer0_outputs(3761) <= not (a or b);
    layer0_outputs(3762) <= not b or a;
    layer0_outputs(3763) <= a and not b;
    layer0_outputs(3764) <= not (a xor b);
    layer0_outputs(3765) <= not (a and b);
    layer0_outputs(3766) <= b;
    layer0_outputs(3767) <= a;
    layer0_outputs(3768) <= not (a or b);
    layer0_outputs(3769) <= b and not a;
    layer0_outputs(3770) <= not (a or b);
    layer0_outputs(3771) <= a xor b;
    layer0_outputs(3772) <= not (a xor b);
    layer0_outputs(3773) <= b and not a;
    layer0_outputs(3774) <= a;
    layer0_outputs(3775) <= not a or b;
    layer0_outputs(3776) <= not b;
    layer0_outputs(3777) <= 1'b1;
    layer0_outputs(3778) <= not b or a;
    layer0_outputs(3779) <= b;
    layer0_outputs(3780) <= a xor b;
    layer0_outputs(3781) <= not a;
    layer0_outputs(3782) <= not a or b;
    layer0_outputs(3783) <= a;
    layer0_outputs(3784) <= not b;
    layer0_outputs(3785) <= a and not b;
    layer0_outputs(3786) <= b and not a;
    layer0_outputs(3787) <= not (a xor b);
    layer0_outputs(3788) <= not b or a;
    layer0_outputs(3789) <= a xor b;
    layer0_outputs(3790) <= not b or a;
    layer0_outputs(3791) <= a xor b;
    layer0_outputs(3792) <= not (a xor b);
    layer0_outputs(3793) <= not a or b;
    layer0_outputs(3794) <= not a or b;
    layer0_outputs(3795) <= not a or b;
    layer0_outputs(3796) <= b;
    layer0_outputs(3797) <= 1'b0;
    layer0_outputs(3798) <= a xor b;
    layer0_outputs(3799) <= a or b;
    layer0_outputs(3800) <= not b;
    layer0_outputs(3801) <= a or b;
    layer0_outputs(3802) <= not b;
    layer0_outputs(3803) <= b;
    layer0_outputs(3804) <= 1'b0;
    layer0_outputs(3805) <= not a or b;
    layer0_outputs(3806) <= a and not b;
    layer0_outputs(3807) <= 1'b0;
    layer0_outputs(3808) <= not (a xor b);
    layer0_outputs(3809) <= a or b;
    layer0_outputs(3810) <= not (a xor b);
    layer0_outputs(3811) <= a or b;
    layer0_outputs(3812) <= not a or b;
    layer0_outputs(3813) <= not (a xor b);
    layer0_outputs(3814) <= not (a or b);
    layer0_outputs(3815) <= not (a xor b);
    layer0_outputs(3816) <= b and not a;
    layer0_outputs(3817) <= not b or a;
    layer0_outputs(3818) <= not a or b;
    layer0_outputs(3819) <= b;
    layer0_outputs(3820) <= not b;
    layer0_outputs(3821) <= a or b;
    layer0_outputs(3822) <= b;
    layer0_outputs(3823) <= b and not a;
    layer0_outputs(3824) <= a xor b;
    layer0_outputs(3825) <= not a;
    layer0_outputs(3826) <= b and not a;
    layer0_outputs(3827) <= 1'b1;
    layer0_outputs(3828) <= b;
    layer0_outputs(3829) <= not a;
    layer0_outputs(3830) <= not a or b;
    layer0_outputs(3831) <= not b;
    layer0_outputs(3832) <= not (a xor b);
    layer0_outputs(3833) <= not b;
    layer0_outputs(3834) <= not (a or b);
    layer0_outputs(3835) <= not (a xor b);
    layer0_outputs(3836) <= not a;
    layer0_outputs(3837) <= b and not a;
    layer0_outputs(3838) <= not (a or b);
    layer0_outputs(3839) <= not (a or b);
    layer0_outputs(3840) <= a xor b;
    layer0_outputs(3841) <= not a or b;
    layer0_outputs(3842) <= a or b;
    layer0_outputs(3843) <= a;
    layer0_outputs(3844) <= 1'b1;
    layer0_outputs(3845) <= not (a or b);
    layer0_outputs(3846) <= b;
    layer0_outputs(3847) <= not (a xor b);
    layer0_outputs(3848) <= b and not a;
    layer0_outputs(3849) <= not (a xor b);
    layer0_outputs(3850) <= a xor b;
    layer0_outputs(3851) <= a xor b;
    layer0_outputs(3852) <= not b;
    layer0_outputs(3853) <= not a or b;
    layer0_outputs(3854) <= a;
    layer0_outputs(3855) <= not a;
    layer0_outputs(3856) <= b and not a;
    layer0_outputs(3857) <= not a or b;
    layer0_outputs(3858) <= not a or b;
    layer0_outputs(3859) <= 1'b1;
    layer0_outputs(3860) <= not b or a;
    layer0_outputs(3861) <= b;
    layer0_outputs(3862) <= a xor b;
    layer0_outputs(3863) <= a or b;
    layer0_outputs(3864) <= not a or b;
    layer0_outputs(3865) <= b and not a;
    layer0_outputs(3866) <= 1'b0;
    layer0_outputs(3867) <= a or b;
    layer0_outputs(3868) <= a;
    layer0_outputs(3869) <= not (a xor b);
    layer0_outputs(3870) <= not a;
    layer0_outputs(3871) <= not (a xor b);
    layer0_outputs(3872) <= not b;
    layer0_outputs(3873) <= a or b;
    layer0_outputs(3874) <= 1'b1;
    layer0_outputs(3875) <= a or b;
    layer0_outputs(3876) <= not a;
    layer0_outputs(3877) <= 1'b1;
    layer0_outputs(3878) <= not (a or b);
    layer0_outputs(3879) <= b and not a;
    layer0_outputs(3880) <= a;
    layer0_outputs(3881) <= a;
    layer0_outputs(3882) <= not (a xor b);
    layer0_outputs(3883) <= not a;
    layer0_outputs(3884) <= a or b;
    layer0_outputs(3885) <= b;
    layer0_outputs(3886) <= a xor b;
    layer0_outputs(3887) <= 1'b0;
    layer0_outputs(3888) <= not b;
    layer0_outputs(3889) <= not (a xor b);
    layer0_outputs(3890) <= a xor b;
    layer0_outputs(3891) <= 1'b1;
    layer0_outputs(3892) <= not a;
    layer0_outputs(3893) <= a and b;
    layer0_outputs(3894) <= b;
    layer0_outputs(3895) <= a and not b;
    layer0_outputs(3896) <= not (a and b);
    layer0_outputs(3897) <= a;
    layer0_outputs(3898) <= a xor b;
    layer0_outputs(3899) <= a or b;
    layer0_outputs(3900) <= not (a or b);
    layer0_outputs(3901) <= b;
    layer0_outputs(3902) <= b and not a;
    layer0_outputs(3903) <= not b;
    layer0_outputs(3904) <= a and b;
    layer0_outputs(3905) <= not b or a;
    layer0_outputs(3906) <= a or b;
    layer0_outputs(3907) <= not (a xor b);
    layer0_outputs(3908) <= b;
    layer0_outputs(3909) <= a and b;
    layer0_outputs(3910) <= not a;
    layer0_outputs(3911) <= a and not b;
    layer0_outputs(3912) <= not a or b;
    layer0_outputs(3913) <= not a;
    layer0_outputs(3914) <= a xor b;
    layer0_outputs(3915) <= 1'b0;
    layer0_outputs(3916) <= not a;
    layer0_outputs(3917) <= not (a xor b);
    layer0_outputs(3918) <= b;
    layer0_outputs(3919) <= b and not a;
    layer0_outputs(3920) <= not (a and b);
    layer0_outputs(3921) <= a;
    layer0_outputs(3922) <= a or b;
    layer0_outputs(3923) <= 1'b1;
    layer0_outputs(3924) <= not a;
    layer0_outputs(3925) <= b and not a;
    layer0_outputs(3926) <= not (a xor b);
    layer0_outputs(3927) <= a;
    layer0_outputs(3928) <= not b;
    layer0_outputs(3929) <= not b or a;
    layer0_outputs(3930) <= a and not b;
    layer0_outputs(3931) <= not a or b;
    layer0_outputs(3932) <= a and not b;
    layer0_outputs(3933) <= not b;
    layer0_outputs(3934) <= not a;
    layer0_outputs(3935) <= not a;
    layer0_outputs(3936) <= not (a or b);
    layer0_outputs(3937) <= not (a xor b);
    layer0_outputs(3938) <= 1'b0;
    layer0_outputs(3939) <= not b or a;
    layer0_outputs(3940) <= not b or a;
    layer0_outputs(3941) <= a or b;
    layer0_outputs(3942) <= not b;
    layer0_outputs(3943) <= a;
    layer0_outputs(3944) <= not (a or b);
    layer0_outputs(3945) <= not a or b;
    layer0_outputs(3946) <= a and b;
    layer0_outputs(3947) <= a or b;
    layer0_outputs(3948) <= not b;
    layer0_outputs(3949) <= a or b;
    layer0_outputs(3950) <= not b;
    layer0_outputs(3951) <= b;
    layer0_outputs(3952) <= not (a or b);
    layer0_outputs(3953) <= not (a xor b);
    layer0_outputs(3954) <= not b or a;
    layer0_outputs(3955) <= a and not b;
    layer0_outputs(3956) <= not b or a;
    layer0_outputs(3957) <= b;
    layer0_outputs(3958) <= b;
    layer0_outputs(3959) <= not b or a;
    layer0_outputs(3960) <= b;
    layer0_outputs(3961) <= b and not a;
    layer0_outputs(3962) <= not (a or b);
    layer0_outputs(3963) <= 1'b1;
    layer0_outputs(3964) <= a or b;
    layer0_outputs(3965) <= not (a xor b);
    layer0_outputs(3966) <= b;
    layer0_outputs(3967) <= not (a or b);
    layer0_outputs(3968) <= b and not a;
    layer0_outputs(3969) <= b;
    layer0_outputs(3970) <= a xor b;
    layer0_outputs(3971) <= not b;
    layer0_outputs(3972) <= not (a or b);
    layer0_outputs(3973) <= a and b;
    layer0_outputs(3974) <= not b or a;
    layer0_outputs(3975) <= a and not b;
    layer0_outputs(3976) <= a xor b;
    layer0_outputs(3977) <= a and not b;
    layer0_outputs(3978) <= a or b;
    layer0_outputs(3979) <= not a or b;
    layer0_outputs(3980) <= not (a xor b);
    layer0_outputs(3981) <= not a or b;
    layer0_outputs(3982) <= b;
    layer0_outputs(3983) <= a or b;
    layer0_outputs(3984) <= not a;
    layer0_outputs(3985) <= a and b;
    layer0_outputs(3986) <= not b;
    layer0_outputs(3987) <= not (a or b);
    layer0_outputs(3988) <= 1'b0;
    layer0_outputs(3989) <= b;
    layer0_outputs(3990) <= b;
    layer0_outputs(3991) <= a;
    layer0_outputs(3992) <= a;
    layer0_outputs(3993) <= not a or b;
    layer0_outputs(3994) <= a and not b;
    layer0_outputs(3995) <= 1'b1;
    layer0_outputs(3996) <= not a or b;
    layer0_outputs(3997) <= a or b;
    layer0_outputs(3998) <= not b or a;
    layer0_outputs(3999) <= a xor b;
    layer0_outputs(4000) <= b;
    layer0_outputs(4001) <= not (a xor b);
    layer0_outputs(4002) <= a and b;
    layer0_outputs(4003) <= a or b;
    layer0_outputs(4004) <= not (a or b);
    layer0_outputs(4005) <= b;
    layer0_outputs(4006) <= not (a or b);
    layer0_outputs(4007) <= 1'b0;
    layer0_outputs(4008) <= not a;
    layer0_outputs(4009) <= b and not a;
    layer0_outputs(4010) <= not a or b;
    layer0_outputs(4011) <= not b;
    layer0_outputs(4012) <= not (a or b);
    layer0_outputs(4013) <= a;
    layer0_outputs(4014) <= 1'b1;
    layer0_outputs(4015) <= b and not a;
    layer0_outputs(4016) <= b and not a;
    layer0_outputs(4017) <= a;
    layer0_outputs(4018) <= not (a and b);
    layer0_outputs(4019) <= a;
    layer0_outputs(4020) <= 1'b1;
    layer0_outputs(4021) <= b;
    layer0_outputs(4022) <= a and not b;
    layer0_outputs(4023) <= not a;
    layer0_outputs(4024) <= a xor b;
    layer0_outputs(4025) <= b and not a;
    layer0_outputs(4026) <= a or b;
    layer0_outputs(4027) <= not a or b;
    layer0_outputs(4028) <= not (a or b);
    layer0_outputs(4029) <= not (a or b);
    layer0_outputs(4030) <= not b or a;
    layer0_outputs(4031) <= not (a xor b);
    layer0_outputs(4032) <= a and not b;
    layer0_outputs(4033) <= b and not a;
    layer0_outputs(4034) <= not (a or b);
    layer0_outputs(4035) <= a and b;
    layer0_outputs(4036) <= not a;
    layer0_outputs(4037) <= a or b;
    layer0_outputs(4038) <= not b;
    layer0_outputs(4039) <= not b or a;
    layer0_outputs(4040) <= not (a and b);
    layer0_outputs(4041) <= not b or a;
    layer0_outputs(4042) <= 1'b1;
    layer0_outputs(4043) <= b;
    layer0_outputs(4044) <= a;
    layer0_outputs(4045) <= not b or a;
    layer0_outputs(4046) <= not a;
    layer0_outputs(4047) <= not b;
    layer0_outputs(4048) <= a;
    layer0_outputs(4049) <= not a;
    layer0_outputs(4050) <= not b or a;
    layer0_outputs(4051) <= a;
    layer0_outputs(4052) <= 1'b1;
    layer0_outputs(4053) <= not (a xor b);
    layer0_outputs(4054) <= not (a xor b);
    layer0_outputs(4055) <= a and b;
    layer0_outputs(4056) <= a or b;
    layer0_outputs(4057) <= a or b;
    layer0_outputs(4058) <= b and not a;
    layer0_outputs(4059) <= not b;
    layer0_outputs(4060) <= 1'b1;
    layer0_outputs(4061) <= b and not a;
    layer0_outputs(4062) <= b and not a;
    layer0_outputs(4063) <= a and not b;
    layer0_outputs(4064) <= not b or a;
    layer0_outputs(4065) <= not (a xor b);
    layer0_outputs(4066) <= a xor b;
    layer0_outputs(4067) <= 1'b1;
    layer0_outputs(4068) <= a or b;
    layer0_outputs(4069) <= a and b;
    layer0_outputs(4070) <= not b or a;
    layer0_outputs(4071) <= a;
    layer0_outputs(4072) <= not a;
    layer0_outputs(4073) <= 1'b0;
    layer0_outputs(4074) <= not (a xor b);
    layer0_outputs(4075) <= not (a or b);
    layer0_outputs(4076) <= a;
    layer0_outputs(4077) <= not (a or b);
    layer0_outputs(4078) <= not (a xor b);
    layer0_outputs(4079) <= not (a or b);
    layer0_outputs(4080) <= a or b;
    layer0_outputs(4081) <= not b;
    layer0_outputs(4082) <= not (a xor b);
    layer0_outputs(4083) <= 1'b0;
    layer0_outputs(4084) <= 1'b1;
    layer0_outputs(4085) <= a xor b;
    layer0_outputs(4086) <= not (a or b);
    layer0_outputs(4087) <= 1'b1;
    layer0_outputs(4088) <= not (a or b);
    layer0_outputs(4089) <= b;
    layer0_outputs(4090) <= not a or b;
    layer0_outputs(4091) <= b and not a;
    layer0_outputs(4092) <= b;
    layer0_outputs(4093) <= not (a xor b);
    layer0_outputs(4094) <= not a;
    layer0_outputs(4095) <= not a or b;
    layer0_outputs(4096) <= b;
    layer0_outputs(4097) <= b and not a;
    layer0_outputs(4098) <= not (a xor b);
    layer0_outputs(4099) <= a;
    layer0_outputs(4100) <= not (a and b);
    layer0_outputs(4101) <= not (a or b);
    layer0_outputs(4102) <= not a or b;
    layer0_outputs(4103) <= not (a xor b);
    layer0_outputs(4104) <= not b;
    layer0_outputs(4105) <= a;
    layer0_outputs(4106) <= b;
    layer0_outputs(4107) <= b and not a;
    layer0_outputs(4108) <= not a;
    layer0_outputs(4109) <= not (a and b);
    layer0_outputs(4110) <= a and b;
    layer0_outputs(4111) <= not (a and b);
    layer0_outputs(4112) <= b and not a;
    layer0_outputs(4113) <= a;
    layer0_outputs(4114) <= not a;
    layer0_outputs(4115) <= b;
    layer0_outputs(4116) <= not (a and b);
    layer0_outputs(4117) <= not (a xor b);
    layer0_outputs(4118) <= not a;
    layer0_outputs(4119) <= a xor b;
    layer0_outputs(4120) <= b and not a;
    layer0_outputs(4121) <= not (a or b);
    layer0_outputs(4122) <= not a;
    layer0_outputs(4123) <= not (a and b);
    layer0_outputs(4124) <= a or b;
    layer0_outputs(4125) <= not a;
    layer0_outputs(4126) <= a or b;
    layer0_outputs(4127) <= not b;
    layer0_outputs(4128) <= 1'b0;
    layer0_outputs(4129) <= not b;
    layer0_outputs(4130) <= a and not b;
    layer0_outputs(4131) <= a or b;
    layer0_outputs(4132) <= a or b;
    layer0_outputs(4133) <= not a;
    layer0_outputs(4134) <= not (a xor b);
    layer0_outputs(4135) <= a or b;
    layer0_outputs(4136) <= not b or a;
    layer0_outputs(4137) <= not (a or b);
    layer0_outputs(4138) <= a or b;
    layer0_outputs(4139) <= 1'b0;
    layer0_outputs(4140) <= not (a or b);
    layer0_outputs(4141) <= not b;
    layer0_outputs(4142) <= not (a xor b);
    layer0_outputs(4143) <= a and not b;
    layer0_outputs(4144) <= not b;
    layer0_outputs(4145) <= not (a or b);
    layer0_outputs(4146) <= 1'b1;
    layer0_outputs(4147) <= a xor b;
    layer0_outputs(4148) <= not (a or b);
    layer0_outputs(4149) <= not (a xor b);
    layer0_outputs(4150) <= a and b;
    layer0_outputs(4151) <= not (a and b);
    layer0_outputs(4152) <= not (a or b);
    layer0_outputs(4153) <= a;
    layer0_outputs(4154) <= not (a or b);
    layer0_outputs(4155) <= a xor b;
    layer0_outputs(4156) <= a;
    layer0_outputs(4157) <= a or b;
    layer0_outputs(4158) <= not (a or b);
    layer0_outputs(4159) <= not a;
    layer0_outputs(4160) <= b and not a;
    layer0_outputs(4161) <= not (a or b);
    layer0_outputs(4162) <= not a or b;
    layer0_outputs(4163) <= a or b;
    layer0_outputs(4164) <= b and not a;
    layer0_outputs(4165) <= not (a xor b);
    layer0_outputs(4166) <= not (a xor b);
    layer0_outputs(4167) <= a and b;
    layer0_outputs(4168) <= not a or b;
    layer0_outputs(4169) <= not (a or b);
    layer0_outputs(4170) <= not b;
    layer0_outputs(4171) <= a and not b;
    layer0_outputs(4172) <= 1'b0;
    layer0_outputs(4173) <= a and not b;
    layer0_outputs(4174) <= not a or b;
    layer0_outputs(4175) <= a and not b;
    layer0_outputs(4176) <= a and b;
    layer0_outputs(4177) <= not a or b;
    layer0_outputs(4178) <= not a;
    layer0_outputs(4179) <= not (a xor b);
    layer0_outputs(4180) <= not a;
    layer0_outputs(4181) <= b;
    layer0_outputs(4182) <= 1'b1;
    layer0_outputs(4183) <= not (a or b);
    layer0_outputs(4184) <= a or b;
    layer0_outputs(4185) <= a and b;
    layer0_outputs(4186) <= not a or b;
    layer0_outputs(4187) <= not b;
    layer0_outputs(4188) <= b and not a;
    layer0_outputs(4189) <= not a or b;
    layer0_outputs(4190) <= not (a xor b);
    layer0_outputs(4191) <= not b;
    layer0_outputs(4192) <= not a;
    layer0_outputs(4193) <= not (a xor b);
    layer0_outputs(4194) <= a;
    layer0_outputs(4195) <= 1'b0;
    layer0_outputs(4196) <= not b or a;
    layer0_outputs(4197) <= not b or a;
    layer0_outputs(4198) <= a and not b;
    layer0_outputs(4199) <= a xor b;
    layer0_outputs(4200) <= a or b;
    layer0_outputs(4201) <= not a;
    layer0_outputs(4202) <= not b or a;
    layer0_outputs(4203) <= 1'b1;
    layer0_outputs(4204) <= 1'b1;
    layer0_outputs(4205) <= not b or a;
    layer0_outputs(4206) <= not b or a;
    layer0_outputs(4207) <= a;
    layer0_outputs(4208) <= a or b;
    layer0_outputs(4209) <= 1'b0;
    layer0_outputs(4210) <= a xor b;
    layer0_outputs(4211) <= not b;
    layer0_outputs(4212) <= a;
    layer0_outputs(4213) <= a and not b;
    layer0_outputs(4214) <= a and not b;
    layer0_outputs(4215) <= a or b;
    layer0_outputs(4216) <= not (a or b);
    layer0_outputs(4217) <= not (a or b);
    layer0_outputs(4218) <= not b or a;
    layer0_outputs(4219) <= not b;
    layer0_outputs(4220) <= 1'b1;
    layer0_outputs(4221) <= not b or a;
    layer0_outputs(4222) <= b;
    layer0_outputs(4223) <= a;
    layer0_outputs(4224) <= 1'b0;
    layer0_outputs(4225) <= not (a or b);
    layer0_outputs(4226) <= not a or b;
    layer0_outputs(4227) <= not b or a;
    layer0_outputs(4228) <= 1'b1;
    layer0_outputs(4229) <= b and not a;
    layer0_outputs(4230) <= not b;
    layer0_outputs(4231) <= not a;
    layer0_outputs(4232) <= not a;
    layer0_outputs(4233) <= not (a xor b);
    layer0_outputs(4234) <= a;
    layer0_outputs(4235) <= not a;
    layer0_outputs(4236) <= not a or b;
    layer0_outputs(4237) <= not (a and b);
    layer0_outputs(4238) <= a or b;
    layer0_outputs(4239) <= 1'b1;
    layer0_outputs(4240) <= not b;
    layer0_outputs(4241) <= a;
    layer0_outputs(4242) <= not a;
    layer0_outputs(4243) <= not (a xor b);
    layer0_outputs(4244) <= b;
    layer0_outputs(4245) <= not (a and b);
    layer0_outputs(4246) <= not (a and b);
    layer0_outputs(4247) <= a xor b;
    layer0_outputs(4248) <= not a or b;
    layer0_outputs(4249) <= not b or a;
    layer0_outputs(4250) <= not a;
    layer0_outputs(4251) <= not b;
    layer0_outputs(4252) <= a and b;
    layer0_outputs(4253) <= a and not b;
    layer0_outputs(4254) <= not a or b;
    layer0_outputs(4255) <= a;
    layer0_outputs(4256) <= not b;
    layer0_outputs(4257) <= b;
    layer0_outputs(4258) <= not a;
    layer0_outputs(4259) <= not a;
    layer0_outputs(4260) <= not b or a;
    layer0_outputs(4261) <= not (a or b);
    layer0_outputs(4262) <= a;
    layer0_outputs(4263) <= not a or b;
    layer0_outputs(4264) <= a xor b;
    layer0_outputs(4265) <= a or b;
    layer0_outputs(4266) <= a;
    layer0_outputs(4267) <= a or b;
    layer0_outputs(4268) <= a and not b;
    layer0_outputs(4269) <= not (a or b);
    layer0_outputs(4270) <= not (a or b);
    layer0_outputs(4271) <= not (a or b);
    layer0_outputs(4272) <= not b;
    layer0_outputs(4273) <= a and b;
    layer0_outputs(4274) <= not a or b;
    layer0_outputs(4275) <= not a or b;
    layer0_outputs(4276) <= a and not b;
    layer0_outputs(4277) <= a xor b;
    layer0_outputs(4278) <= a xor b;
    layer0_outputs(4279) <= not b;
    layer0_outputs(4280) <= a and not b;
    layer0_outputs(4281) <= not (a or b);
    layer0_outputs(4282) <= a xor b;
    layer0_outputs(4283) <= not (a or b);
    layer0_outputs(4284) <= a;
    layer0_outputs(4285) <= a and not b;
    layer0_outputs(4286) <= not b or a;
    layer0_outputs(4287) <= a and b;
    layer0_outputs(4288) <= b;
    layer0_outputs(4289) <= not b;
    layer0_outputs(4290) <= a or b;
    layer0_outputs(4291) <= not a;
    layer0_outputs(4292) <= b;
    layer0_outputs(4293) <= not (a or b);
    layer0_outputs(4294) <= not b;
    layer0_outputs(4295) <= not a or b;
    layer0_outputs(4296) <= a;
    layer0_outputs(4297) <= not b;
    layer0_outputs(4298) <= not b;
    layer0_outputs(4299) <= a xor b;
    layer0_outputs(4300) <= a or b;
    layer0_outputs(4301) <= a and not b;
    layer0_outputs(4302) <= not a;
    layer0_outputs(4303) <= b and not a;
    layer0_outputs(4304) <= 1'b1;
    layer0_outputs(4305) <= a and not b;
    layer0_outputs(4306) <= not a;
    layer0_outputs(4307) <= not b;
    layer0_outputs(4308) <= not (a xor b);
    layer0_outputs(4309) <= not a or b;
    layer0_outputs(4310) <= not (a xor b);
    layer0_outputs(4311) <= 1'b1;
    layer0_outputs(4312) <= 1'b1;
    layer0_outputs(4313) <= b and not a;
    layer0_outputs(4314) <= b;
    layer0_outputs(4315) <= 1'b1;
    layer0_outputs(4316) <= a;
    layer0_outputs(4317) <= not b or a;
    layer0_outputs(4318) <= b;
    layer0_outputs(4319) <= a xor b;
    layer0_outputs(4320) <= a or b;
    layer0_outputs(4321) <= not (a or b);
    layer0_outputs(4322) <= not (a xor b);
    layer0_outputs(4323) <= not (a or b);
    layer0_outputs(4324) <= not a;
    layer0_outputs(4325) <= a or b;
    layer0_outputs(4326) <= not (a or b);
    layer0_outputs(4327) <= not b or a;
    layer0_outputs(4328) <= not a;
    layer0_outputs(4329) <= a;
    layer0_outputs(4330) <= not (a or b);
    layer0_outputs(4331) <= not a or b;
    layer0_outputs(4332) <= not a;
    layer0_outputs(4333) <= not (a and b);
    layer0_outputs(4334) <= a and b;
    layer0_outputs(4335) <= b and not a;
    layer0_outputs(4336) <= 1'b0;
    layer0_outputs(4337) <= not a;
    layer0_outputs(4338) <= a;
    layer0_outputs(4339) <= not b or a;
    layer0_outputs(4340) <= 1'b1;
    layer0_outputs(4341) <= b;
    layer0_outputs(4342) <= not (a or b);
    layer0_outputs(4343) <= not (a or b);
    layer0_outputs(4344) <= a xor b;
    layer0_outputs(4345) <= not b or a;
    layer0_outputs(4346) <= a and not b;
    layer0_outputs(4347) <= not a or b;
    layer0_outputs(4348) <= a and b;
    layer0_outputs(4349) <= a xor b;
    layer0_outputs(4350) <= not a or b;
    layer0_outputs(4351) <= a and b;
    layer0_outputs(4352) <= a xor b;
    layer0_outputs(4353) <= a xor b;
    layer0_outputs(4354) <= not (a or b);
    layer0_outputs(4355) <= not a;
    layer0_outputs(4356) <= not (a or b);
    layer0_outputs(4357) <= not (a or b);
    layer0_outputs(4358) <= a;
    layer0_outputs(4359) <= not (a or b);
    layer0_outputs(4360) <= b and not a;
    layer0_outputs(4361) <= a and not b;
    layer0_outputs(4362) <= not a or b;
    layer0_outputs(4363) <= a or b;
    layer0_outputs(4364) <= 1'b0;
    layer0_outputs(4365) <= not a;
    layer0_outputs(4366) <= a or b;
    layer0_outputs(4367) <= not a or b;
    layer0_outputs(4368) <= a or b;
    layer0_outputs(4369) <= 1'b0;
    layer0_outputs(4370) <= b and not a;
    layer0_outputs(4371) <= b;
    layer0_outputs(4372) <= a xor b;
    layer0_outputs(4373) <= not a;
    layer0_outputs(4374) <= a or b;
    layer0_outputs(4375) <= a or b;
    layer0_outputs(4376) <= 1'b1;
    layer0_outputs(4377) <= a or b;
    layer0_outputs(4378) <= a and not b;
    layer0_outputs(4379) <= a and b;
    layer0_outputs(4380) <= 1'b0;
    layer0_outputs(4381) <= a or b;
    layer0_outputs(4382) <= a and b;
    layer0_outputs(4383) <= a and not b;
    layer0_outputs(4384) <= not (a or b);
    layer0_outputs(4385) <= a xor b;
    layer0_outputs(4386) <= a or b;
    layer0_outputs(4387) <= not a;
    layer0_outputs(4388) <= not a;
    layer0_outputs(4389) <= not (a or b);
    layer0_outputs(4390) <= not b;
    layer0_outputs(4391) <= b and not a;
    layer0_outputs(4392) <= a or b;
    layer0_outputs(4393) <= a and not b;
    layer0_outputs(4394) <= a xor b;
    layer0_outputs(4395) <= a;
    layer0_outputs(4396) <= not b;
    layer0_outputs(4397) <= not (a and b);
    layer0_outputs(4398) <= b;
    layer0_outputs(4399) <= a or b;
    layer0_outputs(4400) <= a;
    layer0_outputs(4401) <= not a or b;
    layer0_outputs(4402) <= 1'b0;
    layer0_outputs(4403) <= a or b;
    layer0_outputs(4404) <= not (a or b);
    layer0_outputs(4405) <= a or b;
    layer0_outputs(4406) <= a and not b;
    layer0_outputs(4407) <= not (a or b);
    layer0_outputs(4408) <= not b or a;
    layer0_outputs(4409) <= not a;
    layer0_outputs(4410) <= 1'b1;
    layer0_outputs(4411) <= b;
    layer0_outputs(4412) <= not (a or b);
    layer0_outputs(4413) <= 1'b1;
    layer0_outputs(4414) <= b and not a;
    layer0_outputs(4415) <= not b;
    layer0_outputs(4416) <= not b;
    layer0_outputs(4417) <= a and b;
    layer0_outputs(4418) <= a and not b;
    layer0_outputs(4419) <= a or b;
    layer0_outputs(4420) <= a and not b;
    layer0_outputs(4421) <= b;
    layer0_outputs(4422) <= a and not b;
    layer0_outputs(4423) <= not b or a;
    layer0_outputs(4424) <= b;
    layer0_outputs(4425) <= a;
    layer0_outputs(4426) <= a xor b;
    layer0_outputs(4427) <= not b;
    layer0_outputs(4428) <= a and not b;
    layer0_outputs(4429) <= not (a xor b);
    layer0_outputs(4430) <= not (a or b);
    layer0_outputs(4431) <= not b or a;
    layer0_outputs(4432) <= a and not b;
    layer0_outputs(4433) <= not a;
    layer0_outputs(4434) <= a and not b;
    layer0_outputs(4435) <= b;
    layer0_outputs(4436) <= not b or a;
    layer0_outputs(4437) <= not b;
    layer0_outputs(4438) <= b and not a;
    layer0_outputs(4439) <= not a or b;
    layer0_outputs(4440) <= a or b;
    layer0_outputs(4441) <= not a;
    layer0_outputs(4442) <= 1'b0;
    layer0_outputs(4443) <= a xor b;
    layer0_outputs(4444) <= not a or b;
    layer0_outputs(4445) <= not a or b;
    layer0_outputs(4446) <= not (a xor b);
    layer0_outputs(4447) <= a and not b;
    layer0_outputs(4448) <= not a;
    layer0_outputs(4449) <= a;
    layer0_outputs(4450) <= 1'b0;
    layer0_outputs(4451) <= not (a xor b);
    layer0_outputs(4452) <= not (a or b);
    layer0_outputs(4453) <= a and not b;
    layer0_outputs(4454) <= a xor b;
    layer0_outputs(4455) <= a xor b;
    layer0_outputs(4456) <= a and not b;
    layer0_outputs(4457) <= not (a or b);
    layer0_outputs(4458) <= a and not b;
    layer0_outputs(4459) <= a xor b;
    layer0_outputs(4460) <= a;
    layer0_outputs(4461) <= a xor b;
    layer0_outputs(4462) <= not (a xor b);
    layer0_outputs(4463) <= not (a and b);
    layer0_outputs(4464) <= a or b;
    layer0_outputs(4465) <= not (a or b);
    layer0_outputs(4466) <= not (a or b);
    layer0_outputs(4467) <= a xor b;
    layer0_outputs(4468) <= not (a and b);
    layer0_outputs(4469) <= a and b;
    layer0_outputs(4470) <= a xor b;
    layer0_outputs(4471) <= not b or a;
    layer0_outputs(4472) <= 1'b0;
    layer0_outputs(4473) <= b;
    layer0_outputs(4474) <= not (a or b);
    layer0_outputs(4475) <= not a or b;
    layer0_outputs(4476) <= not (a xor b);
    layer0_outputs(4477) <= a;
    layer0_outputs(4478) <= a xor b;
    layer0_outputs(4479) <= a xor b;
    layer0_outputs(4480) <= not b or a;
    layer0_outputs(4481) <= b;
    layer0_outputs(4482) <= not a;
    layer0_outputs(4483) <= a and not b;
    layer0_outputs(4484) <= a;
    layer0_outputs(4485) <= not (a and b);
    layer0_outputs(4486) <= a and not b;
    layer0_outputs(4487) <= 1'b1;
    layer0_outputs(4488) <= not (a or b);
    layer0_outputs(4489) <= b;
    layer0_outputs(4490) <= a xor b;
    layer0_outputs(4491) <= a or b;
    layer0_outputs(4492) <= a;
    layer0_outputs(4493) <= not (a or b);
    layer0_outputs(4494) <= not (a xor b);
    layer0_outputs(4495) <= a and b;
    layer0_outputs(4496) <= a and b;
    layer0_outputs(4497) <= a or b;
    layer0_outputs(4498) <= not b or a;
    layer0_outputs(4499) <= not (a and b);
    layer0_outputs(4500) <= not (a or b);
    layer0_outputs(4501) <= b and not a;
    layer0_outputs(4502) <= not (a or b);
    layer0_outputs(4503) <= not b;
    layer0_outputs(4504) <= not (a or b);
    layer0_outputs(4505) <= not (a and b);
    layer0_outputs(4506) <= not (a or b);
    layer0_outputs(4507) <= not (a or b);
    layer0_outputs(4508) <= a and not b;
    layer0_outputs(4509) <= not a;
    layer0_outputs(4510) <= a;
    layer0_outputs(4511) <= not (a xor b);
    layer0_outputs(4512) <= not b;
    layer0_outputs(4513) <= b and not a;
    layer0_outputs(4514) <= 1'b0;
    layer0_outputs(4515) <= b and not a;
    layer0_outputs(4516) <= not a or b;
    layer0_outputs(4517) <= b and not a;
    layer0_outputs(4518) <= a xor b;
    layer0_outputs(4519) <= not (a xor b);
    layer0_outputs(4520) <= b;
    layer0_outputs(4521) <= a and b;
    layer0_outputs(4522) <= a xor b;
    layer0_outputs(4523) <= not (a or b);
    layer0_outputs(4524) <= a and not b;
    layer0_outputs(4525) <= b and not a;
    layer0_outputs(4526) <= b and not a;
    layer0_outputs(4527) <= a xor b;
    layer0_outputs(4528) <= not (a or b);
    layer0_outputs(4529) <= not a;
    layer0_outputs(4530) <= b and not a;
    layer0_outputs(4531) <= not (a or b);
    layer0_outputs(4532) <= a;
    layer0_outputs(4533) <= a;
    layer0_outputs(4534) <= not (a xor b);
    layer0_outputs(4535) <= not (a xor b);
    layer0_outputs(4536) <= 1'b1;
    layer0_outputs(4537) <= a;
    layer0_outputs(4538) <= a and b;
    layer0_outputs(4539) <= a and not b;
    layer0_outputs(4540) <= not (a xor b);
    layer0_outputs(4541) <= not (a and b);
    layer0_outputs(4542) <= not (a or b);
    layer0_outputs(4543) <= not (a or b);
    layer0_outputs(4544) <= a and not b;
    layer0_outputs(4545) <= a xor b;
    layer0_outputs(4546) <= not a or b;
    layer0_outputs(4547) <= b;
    layer0_outputs(4548) <= b;
    layer0_outputs(4549) <= a or b;
    layer0_outputs(4550) <= not (a and b);
    layer0_outputs(4551) <= not (a and b);
    layer0_outputs(4552) <= a xor b;
    layer0_outputs(4553) <= not (a xor b);
    layer0_outputs(4554) <= a or b;
    layer0_outputs(4555) <= not b or a;
    layer0_outputs(4556) <= a;
    layer0_outputs(4557) <= not (a and b);
    layer0_outputs(4558) <= not b;
    layer0_outputs(4559) <= a xor b;
    layer0_outputs(4560) <= not a or b;
    layer0_outputs(4561) <= a or b;
    layer0_outputs(4562) <= b and not a;
    layer0_outputs(4563) <= a or b;
    layer0_outputs(4564) <= not (a xor b);
    layer0_outputs(4565) <= not b or a;
    layer0_outputs(4566) <= not (a or b);
    layer0_outputs(4567) <= b;
    layer0_outputs(4568) <= b;
    layer0_outputs(4569) <= 1'b0;
    layer0_outputs(4570) <= 1'b0;
    layer0_outputs(4571) <= not (a or b);
    layer0_outputs(4572) <= not b or a;
    layer0_outputs(4573) <= not b;
    layer0_outputs(4574) <= a xor b;
    layer0_outputs(4575) <= 1'b0;
    layer0_outputs(4576) <= not (a or b);
    layer0_outputs(4577) <= a;
    layer0_outputs(4578) <= b and not a;
    layer0_outputs(4579) <= not (a xor b);
    layer0_outputs(4580) <= not (a or b);
    layer0_outputs(4581) <= a or b;
    layer0_outputs(4582) <= not (a and b);
    layer0_outputs(4583) <= a xor b;
    layer0_outputs(4584) <= not a or b;
    layer0_outputs(4585) <= b and not a;
    layer0_outputs(4586) <= not a or b;
    layer0_outputs(4587) <= not b;
    layer0_outputs(4588) <= a and not b;
    layer0_outputs(4589) <= a and not b;
    layer0_outputs(4590) <= b and not a;
    layer0_outputs(4591) <= not a;
    layer0_outputs(4592) <= not b or a;
    layer0_outputs(4593) <= a;
    layer0_outputs(4594) <= a;
    layer0_outputs(4595) <= a xor b;
    layer0_outputs(4596) <= not a or b;
    layer0_outputs(4597) <= not b;
    layer0_outputs(4598) <= 1'b0;
    layer0_outputs(4599) <= not a;
    layer0_outputs(4600) <= not b;
    layer0_outputs(4601) <= not (a xor b);
    layer0_outputs(4602) <= a or b;
    layer0_outputs(4603) <= not (a and b);
    layer0_outputs(4604) <= a;
    layer0_outputs(4605) <= b;
    layer0_outputs(4606) <= not (a and b);
    layer0_outputs(4607) <= not b or a;
    layer0_outputs(4608) <= not (a xor b);
    layer0_outputs(4609) <= 1'b1;
    layer0_outputs(4610) <= b;
    layer0_outputs(4611) <= 1'b0;
    layer0_outputs(4612) <= b and not a;
    layer0_outputs(4613) <= not (a or b);
    layer0_outputs(4614) <= not b;
    layer0_outputs(4615) <= not (a or b);
    layer0_outputs(4616) <= not b or a;
    layer0_outputs(4617) <= not (a or b);
    layer0_outputs(4618) <= a xor b;
    layer0_outputs(4619) <= a and b;
    layer0_outputs(4620) <= not a or b;
    layer0_outputs(4621) <= not (a or b);
    layer0_outputs(4622) <= a and b;
    layer0_outputs(4623) <= a;
    layer0_outputs(4624) <= not (a or b);
    layer0_outputs(4625) <= a or b;
    layer0_outputs(4626) <= 1'b1;
    layer0_outputs(4627) <= a xor b;
    layer0_outputs(4628) <= a and b;
    layer0_outputs(4629) <= not a or b;
    layer0_outputs(4630) <= a and b;
    layer0_outputs(4631) <= 1'b1;
    layer0_outputs(4632) <= a or b;
    layer0_outputs(4633) <= not b;
    layer0_outputs(4634) <= a xor b;
    layer0_outputs(4635) <= b and not a;
    layer0_outputs(4636) <= not b or a;
    layer0_outputs(4637) <= not (a xor b);
    layer0_outputs(4638) <= 1'b0;
    layer0_outputs(4639) <= a and b;
    layer0_outputs(4640) <= a;
    layer0_outputs(4641) <= 1'b0;
    layer0_outputs(4642) <= a;
    layer0_outputs(4643) <= not a;
    layer0_outputs(4644) <= not a;
    layer0_outputs(4645) <= not (a or b);
    layer0_outputs(4646) <= not b or a;
    layer0_outputs(4647) <= a and not b;
    layer0_outputs(4648) <= not a or b;
    layer0_outputs(4649) <= b and not a;
    layer0_outputs(4650) <= not a or b;
    layer0_outputs(4651) <= 1'b1;
    layer0_outputs(4652) <= not (a or b);
    layer0_outputs(4653) <= b;
    layer0_outputs(4654) <= b;
    layer0_outputs(4655) <= not b;
    layer0_outputs(4656) <= not a or b;
    layer0_outputs(4657) <= not a;
    layer0_outputs(4658) <= a xor b;
    layer0_outputs(4659) <= not (a or b);
    layer0_outputs(4660) <= a;
    layer0_outputs(4661) <= not (a and b);
    layer0_outputs(4662) <= 1'b0;
    layer0_outputs(4663) <= not a;
    layer0_outputs(4664) <= a;
    layer0_outputs(4665) <= not b;
    layer0_outputs(4666) <= a;
    layer0_outputs(4667) <= not b;
    layer0_outputs(4668) <= b and not a;
    layer0_outputs(4669) <= 1'b1;
    layer0_outputs(4670) <= not b;
    layer0_outputs(4671) <= not b or a;
    layer0_outputs(4672) <= not (a or b);
    layer0_outputs(4673) <= b;
    layer0_outputs(4674) <= not (a and b);
    layer0_outputs(4675) <= a or b;
    layer0_outputs(4676) <= not b;
    layer0_outputs(4677) <= not (a xor b);
    layer0_outputs(4678) <= b;
    layer0_outputs(4679) <= 1'b1;
    layer0_outputs(4680) <= a xor b;
    layer0_outputs(4681) <= not b or a;
    layer0_outputs(4682) <= a and b;
    layer0_outputs(4683) <= not (a or b);
    layer0_outputs(4684) <= b;
    layer0_outputs(4685) <= a or b;
    layer0_outputs(4686) <= a;
    layer0_outputs(4687) <= a xor b;
    layer0_outputs(4688) <= not a;
    layer0_outputs(4689) <= not a;
    layer0_outputs(4690) <= not (a and b);
    layer0_outputs(4691) <= not (a or b);
    layer0_outputs(4692) <= 1'b0;
    layer0_outputs(4693) <= b;
    layer0_outputs(4694) <= a or b;
    layer0_outputs(4695) <= a and not b;
    layer0_outputs(4696) <= not a;
    layer0_outputs(4697) <= a or b;
    layer0_outputs(4698) <= a xor b;
    layer0_outputs(4699) <= a or b;
    layer0_outputs(4700) <= a;
    layer0_outputs(4701) <= a;
    layer0_outputs(4702) <= a and b;
    layer0_outputs(4703) <= b and not a;
    layer0_outputs(4704) <= not (a or b);
    layer0_outputs(4705) <= not a or b;
    layer0_outputs(4706) <= not b or a;
    layer0_outputs(4707) <= not a;
    layer0_outputs(4708) <= not (a or b);
    layer0_outputs(4709) <= not (a xor b);
    layer0_outputs(4710) <= 1'b0;
    layer0_outputs(4711) <= b and not a;
    layer0_outputs(4712) <= a or b;
    layer0_outputs(4713) <= not b;
    layer0_outputs(4714) <= b and not a;
    layer0_outputs(4715) <= not b;
    layer0_outputs(4716) <= not b or a;
    layer0_outputs(4717) <= not (a xor b);
    layer0_outputs(4718) <= not (a or b);
    layer0_outputs(4719) <= a;
    layer0_outputs(4720) <= not (a and b);
    layer0_outputs(4721) <= a and b;
    layer0_outputs(4722) <= not b;
    layer0_outputs(4723) <= b;
    layer0_outputs(4724) <= a xor b;
    layer0_outputs(4725) <= b;
    layer0_outputs(4726) <= 1'b0;
    layer0_outputs(4727) <= a xor b;
    layer0_outputs(4728) <= a and not b;
    layer0_outputs(4729) <= b and not a;
    layer0_outputs(4730) <= not (a xor b);
    layer0_outputs(4731) <= not (a or b);
    layer0_outputs(4732) <= a or b;
    layer0_outputs(4733) <= not a or b;
    layer0_outputs(4734) <= not (a xor b);
    layer0_outputs(4735) <= not (a xor b);
    layer0_outputs(4736) <= b;
    layer0_outputs(4737) <= not (a or b);
    layer0_outputs(4738) <= a xor b;
    layer0_outputs(4739) <= not a or b;
    layer0_outputs(4740) <= a and not b;
    layer0_outputs(4741) <= not (a and b);
    layer0_outputs(4742) <= not a;
    layer0_outputs(4743) <= not (a and b);
    layer0_outputs(4744) <= a;
    layer0_outputs(4745) <= not b;
    layer0_outputs(4746) <= a or b;
    layer0_outputs(4747) <= not (a or b);
    layer0_outputs(4748) <= not a;
    layer0_outputs(4749) <= not b;
    layer0_outputs(4750) <= a xor b;
    layer0_outputs(4751) <= not a or b;
    layer0_outputs(4752) <= not a;
    layer0_outputs(4753) <= not a or b;
    layer0_outputs(4754) <= not a or b;
    layer0_outputs(4755) <= 1'b0;
    layer0_outputs(4756) <= not a;
    layer0_outputs(4757) <= not a;
    layer0_outputs(4758) <= a xor b;
    layer0_outputs(4759) <= not (a or b);
    layer0_outputs(4760) <= a xor b;
    layer0_outputs(4761) <= a xor b;
    layer0_outputs(4762) <= not (a xor b);
    layer0_outputs(4763) <= 1'b0;
    layer0_outputs(4764) <= b;
    layer0_outputs(4765) <= b;
    layer0_outputs(4766) <= not (a or b);
    layer0_outputs(4767) <= a;
    layer0_outputs(4768) <= a xor b;
    layer0_outputs(4769) <= not (a xor b);
    layer0_outputs(4770) <= not b or a;
    layer0_outputs(4771) <= not (a xor b);
    layer0_outputs(4772) <= not b;
    layer0_outputs(4773) <= a or b;
    layer0_outputs(4774) <= b and not a;
    layer0_outputs(4775) <= not (a or b);
    layer0_outputs(4776) <= a;
    layer0_outputs(4777) <= a and b;
    layer0_outputs(4778) <= not (a or b);
    layer0_outputs(4779) <= not b or a;
    layer0_outputs(4780) <= not b;
    layer0_outputs(4781) <= a and not b;
    layer0_outputs(4782) <= 1'b0;
    layer0_outputs(4783) <= not (a and b);
    layer0_outputs(4784) <= not b or a;
    layer0_outputs(4785) <= a or b;
    layer0_outputs(4786) <= not (a or b);
    layer0_outputs(4787) <= a;
    layer0_outputs(4788) <= a xor b;
    layer0_outputs(4789) <= not (a or b);
    layer0_outputs(4790) <= b and not a;
    layer0_outputs(4791) <= a or b;
    layer0_outputs(4792) <= not (a xor b);
    layer0_outputs(4793) <= not (a xor b);
    layer0_outputs(4794) <= not b;
    layer0_outputs(4795) <= b;
    layer0_outputs(4796) <= a or b;
    layer0_outputs(4797) <= a xor b;
    layer0_outputs(4798) <= b and not a;
    layer0_outputs(4799) <= not (a and b);
    layer0_outputs(4800) <= not (a or b);
    layer0_outputs(4801) <= a and b;
    layer0_outputs(4802) <= b;
    layer0_outputs(4803) <= not a or b;
    layer0_outputs(4804) <= 1'b1;
    layer0_outputs(4805) <= a or b;
    layer0_outputs(4806) <= not b or a;
    layer0_outputs(4807) <= not (a or b);
    layer0_outputs(4808) <= 1'b1;
    layer0_outputs(4809) <= not a or b;
    layer0_outputs(4810) <= not (a or b);
    layer0_outputs(4811) <= not b;
    layer0_outputs(4812) <= not b;
    layer0_outputs(4813) <= not b;
    layer0_outputs(4814) <= 1'b0;
    layer0_outputs(4815) <= not a;
    layer0_outputs(4816) <= a;
    layer0_outputs(4817) <= a and not b;
    layer0_outputs(4818) <= not (a xor b);
    layer0_outputs(4819) <= not b;
    layer0_outputs(4820) <= not (a or b);
    layer0_outputs(4821) <= a and not b;
    layer0_outputs(4822) <= not (a and b);
    layer0_outputs(4823) <= not (a or b);
    layer0_outputs(4824) <= not (a xor b);
    layer0_outputs(4825) <= a and b;
    layer0_outputs(4826) <= not b;
    layer0_outputs(4827) <= not (a or b);
    layer0_outputs(4828) <= a and not b;
    layer0_outputs(4829) <= not a;
    layer0_outputs(4830) <= a;
    layer0_outputs(4831) <= a xor b;
    layer0_outputs(4832) <= not (a xor b);
    layer0_outputs(4833) <= not (a xor b);
    layer0_outputs(4834) <= b and not a;
    layer0_outputs(4835) <= 1'b0;
    layer0_outputs(4836) <= a;
    layer0_outputs(4837) <= a or b;
    layer0_outputs(4838) <= not (a and b);
    layer0_outputs(4839) <= a xor b;
    layer0_outputs(4840) <= not (a or b);
    layer0_outputs(4841) <= not (a xor b);
    layer0_outputs(4842) <= not a or b;
    layer0_outputs(4843) <= not (a and b);
    layer0_outputs(4844) <= not (a and b);
    layer0_outputs(4845) <= a xor b;
    layer0_outputs(4846) <= not a or b;
    layer0_outputs(4847) <= a or b;
    layer0_outputs(4848) <= a and not b;
    layer0_outputs(4849) <= not a;
    layer0_outputs(4850) <= a or b;
    layer0_outputs(4851) <= a and not b;
    layer0_outputs(4852) <= not a;
    layer0_outputs(4853) <= b and not a;
    layer0_outputs(4854) <= b;
    layer0_outputs(4855) <= not b;
    layer0_outputs(4856) <= a or b;
    layer0_outputs(4857) <= not a;
    layer0_outputs(4858) <= a and b;
    layer0_outputs(4859) <= a and not b;
    layer0_outputs(4860) <= 1'b1;
    layer0_outputs(4861) <= not b;
    layer0_outputs(4862) <= not b;
    layer0_outputs(4863) <= a xor b;
    layer0_outputs(4864) <= not b or a;
    layer0_outputs(4865) <= a or b;
    layer0_outputs(4866) <= a and not b;
    layer0_outputs(4867) <= not b;
    layer0_outputs(4868) <= not (a and b);
    layer0_outputs(4869) <= not a or b;
    layer0_outputs(4870) <= not (a and b);
    layer0_outputs(4871) <= a xor b;
    layer0_outputs(4872) <= not b or a;
    layer0_outputs(4873) <= not a;
    layer0_outputs(4874) <= not b;
    layer0_outputs(4875) <= a xor b;
    layer0_outputs(4876) <= b;
    layer0_outputs(4877) <= not (a or b);
    layer0_outputs(4878) <= 1'b1;
    layer0_outputs(4879) <= a xor b;
    layer0_outputs(4880) <= a and not b;
    layer0_outputs(4881) <= not a or b;
    layer0_outputs(4882) <= b;
    layer0_outputs(4883) <= a xor b;
    layer0_outputs(4884) <= not (a or b);
    layer0_outputs(4885) <= not (a or b);
    layer0_outputs(4886) <= b;
    layer0_outputs(4887) <= not (a or b);
    layer0_outputs(4888) <= a xor b;
    layer0_outputs(4889) <= not (a xor b);
    layer0_outputs(4890) <= b;
    layer0_outputs(4891) <= a or b;
    layer0_outputs(4892) <= a xor b;
    layer0_outputs(4893) <= not a;
    layer0_outputs(4894) <= a xor b;
    layer0_outputs(4895) <= not a or b;
    layer0_outputs(4896) <= b;
    layer0_outputs(4897) <= a and not b;
    layer0_outputs(4898) <= not a or b;
    layer0_outputs(4899) <= not a or b;
    layer0_outputs(4900) <= a xor b;
    layer0_outputs(4901) <= a or b;
    layer0_outputs(4902) <= not a or b;
    layer0_outputs(4903) <= not a;
    layer0_outputs(4904) <= a;
    layer0_outputs(4905) <= a xor b;
    layer0_outputs(4906) <= b;
    layer0_outputs(4907) <= not (a and b);
    layer0_outputs(4908) <= not (a xor b);
    layer0_outputs(4909) <= not b or a;
    layer0_outputs(4910) <= a or b;
    layer0_outputs(4911) <= a and b;
    layer0_outputs(4912) <= b;
    layer0_outputs(4913) <= not (a and b);
    layer0_outputs(4914) <= not a;
    layer0_outputs(4915) <= not b;
    layer0_outputs(4916) <= a;
    layer0_outputs(4917) <= not a or b;
    layer0_outputs(4918) <= not a or b;
    layer0_outputs(4919) <= not b or a;
    layer0_outputs(4920) <= a and not b;
    layer0_outputs(4921) <= a;
    layer0_outputs(4922) <= a or b;
    layer0_outputs(4923) <= not (a xor b);
    layer0_outputs(4924) <= b;
    layer0_outputs(4925) <= b;
    layer0_outputs(4926) <= a or b;
    layer0_outputs(4927) <= not (a or b);
    layer0_outputs(4928) <= a or b;
    layer0_outputs(4929) <= not b;
    layer0_outputs(4930) <= a and b;
    layer0_outputs(4931) <= not (a or b);
    layer0_outputs(4932) <= a;
    layer0_outputs(4933) <= not (a or b);
    layer0_outputs(4934) <= a and not b;
    layer0_outputs(4935) <= a xor b;
    layer0_outputs(4936) <= not a;
    layer0_outputs(4937) <= not (a or b);
    layer0_outputs(4938) <= not b or a;
    layer0_outputs(4939) <= a or b;
    layer0_outputs(4940) <= 1'b1;
    layer0_outputs(4941) <= not (a xor b);
    layer0_outputs(4942) <= a xor b;
    layer0_outputs(4943) <= not (a or b);
    layer0_outputs(4944) <= not a;
    layer0_outputs(4945) <= b;
    layer0_outputs(4946) <= not (a xor b);
    layer0_outputs(4947) <= not (a xor b);
    layer0_outputs(4948) <= a;
    layer0_outputs(4949) <= 1'b0;
    layer0_outputs(4950) <= b and not a;
    layer0_outputs(4951) <= a;
    layer0_outputs(4952) <= not a;
    layer0_outputs(4953) <= not b;
    layer0_outputs(4954) <= not b or a;
    layer0_outputs(4955) <= b and not a;
    layer0_outputs(4956) <= b and not a;
    layer0_outputs(4957) <= not a;
    layer0_outputs(4958) <= a xor b;
    layer0_outputs(4959) <= not (a xor b);
    layer0_outputs(4960) <= not (a and b);
    layer0_outputs(4961) <= not a;
    layer0_outputs(4962) <= not (a xor b);
    layer0_outputs(4963) <= 1'b1;
    layer0_outputs(4964) <= not (a or b);
    layer0_outputs(4965) <= 1'b1;
    layer0_outputs(4966) <= not (a or b);
    layer0_outputs(4967) <= a xor b;
    layer0_outputs(4968) <= b and not a;
    layer0_outputs(4969) <= a or b;
    layer0_outputs(4970) <= not (a and b);
    layer0_outputs(4971) <= not a;
    layer0_outputs(4972) <= 1'b1;
    layer0_outputs(4973) <= not a or b;
    layer0_outputs(4974) <= not a or b;
    layer0_outputs(4975) <= b;
    layer0_outputs(4976) <= not b;
    layer0_outputs(4977) <= a xor b;
    layer0_outputs(4978) <= 1'b0;
    layer0_outputs(4979) <= b;
    layer0_outputs(4980) <= not (a xor b);
    layer0_outputs(4981) <= b;
    layer0_outputs(4982) <= 1'b1;
    layer0_outputs(4983) <= b and not a;
    layer0_outputs(4984) <= a;
    layer0_outputs(4985) <= not a;
    layer0_outputs(4986) <= not a;
    layer0_outputs(4987) <= not b;
    layer0_outputs(4988) <= a xor b;
    layer0_outputs(4989) <= b;
    layer0_outputs(4990) <= not (a or b);
    layer0_outputs(4991) <= a or b;
    layer0_outputs(4992) <= b;
    layer0_outputs(4993) <= not (a or b);
    layer0_outputs(4994) <= not b or a;
    layer0_outputs(4995) <= not (a or b);
    layer0_outputs(4996) <= 1'b1;
    layer0_outputs(4997) <= a and not b;
    layer0_outputs(4998) <= not a or b;
    layer0_outputs(4999) <= not b;
    layer0_outputs(5000) <= not b;
    layer0_outputs(5001) <= a;
    layer0_outputs(5002) <= b and not a;
    layer0_outputs(5003) <= not b;
    layer0_outputs(5004) <= not a or b;
    layer0_outputs(5005) <= a and not b;
    layer0_outputs(5006) <= a;
    layer0_outputs(5007) <= b;
    layer0_outputs(5008) <= a xor b;
    layer0_outputs(5009) <= not (a and b);
    layer0_outputs(5010) <= 1'b0;
    layer0_outputs(5011) <= not (a xor b);
    layer0_outputs(5012) <= b and not a;
    layer0_outputs(5013) <= b;
    layer0_outputs(5014) <= not a or b;
    layer0_outputs(5015) <= a and b;
    layer0_outputs(5016) <= 1'b1;
    layer0_outputs(5017) <= 1'b0;
    layer0_outputs(5018) <= not b or a;
    layer0_outputs(5019) <= a;
    layer0_outputs(5020) <= not (a or b);
    layer0_outputs(5021) <= not (a xor b);
    layer0_outputs(5022) <= not a;
    layer0_outputs(5023) <= b;
    layer0_outputs(5024) <= not (a or b);
    layer0_outputs(5025) <= not (a xor b);
    layer0_outputs(5026) <= a and not b;
    layer0_outputs(5027) <= b and not a;
    layer0_outputs(5028) <= not (a or b);
    layer0_outputs(5029) <= b;
    layer0_outputs(5030) <= not (a and b);
    layer0_outputs(5031) <= 1'b1;
    layer0_outputs(5032) <= a and not b;
    layer0_outputs(5033) <= not (a xor b);
    layer0_outputs(5034) <= not b;
    layer0_outputs(5035) <= b and not a;
    layer0_outputs(5036) <= a;
    layer0_outputs(5037) <= a or b;
    layer0_outputs(5038) <= a and b;
    layer0_outputs(5039) <= not b;
    layer0_outputs(5040) <= 1'b0;
    layer0_outputs(5041) <= b;
    layer0_outputs(5042) <= b and not a;
    layer0_outputs(5043) <= not (a xor b);
    layer0_outputs(5044) <= a xor b;
    layer0_outputs(5045) <= not b;
    layer0_outputs(5046) <= a or b;
    layer0_outputs(5047) <= not b;
    layer0_outputs(5048) <= a or b;
    layer0_outputs(5049) <= a or b;
    layer0_outputs(5050) <= not a;
    layer0_outputs(5051) <= not (a xor b);
    layer0_outputs(5052) <= not (a and b);
    layer0_outputs(5053) <= not b;
    layer0_outputs(5054) <= not a or b;
    layer0_outputs(5055) <= not (a or b);
    layer0_outputs(5056) <= a and not b;
    layer0_outputs(5057) <= not b or a;
    layer0_outputs(5058) <= b;
    layer0_outputs(5059) <= not b;
    layer0_outputs(5060) <= not (a or b);
    layer0_outputs(5061) <= not (a or b);
    layer0_outputs(5062) <= b and not a;
    layer0_outputs(5063) <= b;
    layer0_outputs(5064) <= not (a xor b);
    layer0_outputs(5065) <= 1'b0;
    layer0_outputs(5066) <= not (a xor b);
    layer0_outputs(5067) <= a xor b;
    layer0_outputs(5068) <= not (a or b);
    layer0_outputs(5069) <= a xor b;
    layer0_outputs(5070) <= b and not a;
    layer0_outputs(5071) <= b and not a;
    layer0_outputs(5072) <= not (a or b);
    layer0_outputs(5073) <= a xor b;
    layer0_outputs(5074) <= a and not b;
    layer0_outputs(5075) <= a and not b;
    layer0_outputs(5076) <= a and b;
    layer0_outputs(5077) <= not b;
    layer0_outputs(5078) <= not b or a;
    layer0_outputs(5079) <= not (a or b);
    layer0_outputs(5080) <= not (a xor b);
    layer0_outputs(5081) <= not (a or b);
    layer0_outputs(5082) <= not a;
    layer0_outputs(5083) <= not a;
    layer0_outputs(5084) <= not b or a;
    layer0_outputs(5085) <= a;
    layer0_outputs(5086) <= b;
    layer0_outputs(5087) <= not (a and b);
    layer0_outputs(5088) <= not b;
    layer0_outputs(5089) <= a or b;
    layer0_outputs(5090) <= a and not b;
    layer0_outputs(5091) <= not b;
    layer0_outputs(5092) <= not a or b;
    layer0_outputs(5093) <= not a or b;
    layer0_outputs(5094) <= b and not a;
    layer0_outputs(5095) <= a;
    layer0_outputs(5096) <= not a or b;
    layer0_outputs(5097) <= a or b;
    layer0_outputs(5098) <= a and not b;
    layer0_outputs(5099) <= not a;
    layer0_outputs(5100) <= b and not a;
    layer0_outputs(5101) <= a and not b;
    layer0_outputs(5102) <= not (a or b);
    layer0_outputs(5103) <= not a or b;
    layer0_outputs(5104) <= not (a or b);
    layer0_outputs(5105) <= b and not a;
    layer0_outputs(5106) <= a;
    layer0_outputs(5107) <= not a or b;
    layer0_outputs(5108) <= 1'b1;
    layer0_outputs(5109) <= not a or b;
    layer0_outputs(5110) <= a xor b;
    layer0_outputs(5111) <= not (a xor b);
    layer0_outputs(5112) <= 1'b1;
    layer0_outputs(5113) <= b and not a;
    layer0_outputs(5114) <= not a;
    layer0_outputs(5115) <= a and not b;
    layer0_outputs(5116) <= a xor b;
    layer0_outputs(5117) <= not (a and b);
    layer0_outputs(5118) <= a and not b;
    layer0_outputs(5119) <= b and not a;
    layer0_outputs(5120) <= a or b;
    layer0_outputs(5121) <= a xor b;
    layer0_outputs(5122) <= a or b;
    layer0_outputs(5123) <= not a or b;
    layer0_outputs(5124) <= b and not a;
    layer0_outputs(5125) <= not (a xor b);
    layer0_outputs(5126) <= not a;
    layer0_outputs(5127) <= a and not b;
    layer0_outputs(5128) <= b;
    layer0_outputs(5129) <= b;
    layer0_outputs(5130) <= a and b;
    layer0_outputs(5131) <= 1'b1;
    layer0_outputs(5132) <= not b or a;
    layer0_outputs(5133) <= a;
    layer0_outputs(5134) <= a;
    layer0_outputs(5135) <= b;
    layer0_outputs(5136) <= not (a xor b);
    layer0_outputs(5137) <= a and b;
    layer0_outputs(5138) <= b and not a;
    layer0_outputs(5139) <= not (a or b);
    layer0_outputs(5140) <= not b;
    layer0_outputs(5141) <= b;
    layer0_outputs(5142) <= a or b;
    layer0_outputs(5143) <= a or b;
    layer0_outputs(5144) <= a;
    layer0_outputs(5145) <= b;
    layer0_outputs(5146) <= not a;
    layer0_outputs(5147) <= not (a or b);
    layer0_outputs(5148) <= not a or b;
    layer0_outputs(5149) <= a xor b;
    layer0_outputs(5150) <= a;
    layer0_outputs(5151) <= not a;
    layer0_outputs(5152) <= not a;
    layer0_outputs(5153) <= not a or b;
    layer0_outputs(5154) <= not b or a;
    layer0_outputs(5155) <= not b or a;
    layer0_outputs(5156) <= a or b;
    layer0_outputs(5157) <= not (a xor b);
    layer0_outputs(5158) <= not (a xor b);
    layer0_outputs(5159) <= not (a xor b);
    layer0_outputs(5160) <= not (a or b);
    layer0_outputs(5161) <= a xor b;
    layer0_outputs(5162) <= not (a or b);
    layer0_outputs(5163) <= not b;
    layer0_outputs(5164) <= not (a xor b);
    layer0_outputs(5165) <= not (a or b);
    layer0_outputs(5166) <= a and not b;
    layer0_outputs(5167) <= a;
    layer0_outputs(5168) <= a;
    layer0_outputs(5169) <= not (a or b);
    layer0_outputs(5170) <= a or b;
    layer0_outputs(5171) <= not (a xor b);
    layer0_outputs(5172) <= not a;
    layer0_outputs(5173) <= a and b;
    layer0_outputs(5174) <= not b;
    layer0_outputs(5175) <= a and not b;
    layer0_outputs(5176) <= not (a and b);
    layer0_outputs(5177) <= b;
    layer0_outputs(5178) <= not a;
    layer0_outputs(5179) <= b and not a;
    layer0_outputs(5180) <= not (a or b);
    layer0_outputs(5181) <= 1'b0;
    layer0_outputs(5182) <= not b;
    layer0_outputs(5183) <= a and b;
    layer0_outputs(5184) <= not a or b;
    layer0_outputs(5185) <= a xor b;
    layer0_outputs(5186) <= 1'b0;
    layer0_outputs(5187) <= not a or b;
    layer0_outputs(5188) <= not (a or b);
    layer0_outputs(5189) <= a xor b;
    layer0_outputs(5190) <= b and not a;
    layer0_outputs(5191) <= not (a or b);
    layer0_outputs(5192) <= not b;
    layer0_outputs(5193) <= not b or a;
    layer0_outputs(5194) <= 1'b0;
    layer0_outputs(5195) <= 1'b1;
    layer0_outputs(5196) <= a or b;
    layer0_outputs(5197) <= a and not b;
    layer0_outputs(5198) <= b;
    layer0_outputs(5199) <= a;
    layer0_outputs(5200) <= not (a or b);
    layer0_outputs(5201) <= a or b;
    layer0_outputs(5202) <= a and not b;
    layer0_outputs(5203) <= not (a or b);
    layer0_outputs(5204) <= not b or a;
    layer0_outputs(5205) <= a or b;
    layer0_outputs(5206) <= not a;
    layer0_outputs(5207) <= a xor b;
    layer0_outputs(5208) <= not (a and b);
    layer0_outputs(5209) <= a xor b;
    layer0_outputs(5210) <= not (a and b);
    layer0_outputs(5211) <= not (a or b);
    layer0_outputs(5212) <= not (a or b);
    layer0_outputs(5213) <= a and b;
    layer0_outputs(5214) <= not b;
    layer0_outputs(5215) <= not (a or b);
    layer0_outputs(5216) <= not b or a;
    layer0_outputs(5217) <= a or b;
    layer0_outputs(5218) <= not a or b;
    layer0_outputs(5219) <= a or b;
    layer0_outputs(5220) <= a or b;
    layer0_outputs(5221) <= not a;
    layer0_outputs(5222) <= not a;
    layer0_outputs(5223) <= a;
    layer0_outputs(5224) <= not (a and b);
    layer0_outputs(5225) <= not b;
    layer0_outputs(5226) <= not (a xor b);
    layer0_outputs(5227) <= a and b;
    layer0_outputs(5228) <= b;
    layer0_outputs(5229) <= not (a or b);
    layer0_outputs(5230) <= b;
    layer0_outputs(5231) <= a or b;
    layer0_outputs(5232) <= a or b;
    layer0_outputs(5233) <= a or b;
    layer0_outputs(5234) <= not a;
    layer0_outputs(5235) <= not b;
    layer0_outputs(5236) <= b;
    layer0_outputs(5237) <= not (a or b);
    layer0_outputs(5238) <= not a or b;
    layer0_outputs(5239) <= not (a or b);
    layer0_outputs(5240) <= a or b;
    layer0_outputs(5241) <= 1'b0;
    layer0_outputs(5242) <= a or b;
    layer0_outputs(5243) <= not a or b;
    layer0_outputs(5244) <= not (a or b);
    layer0_outputs(5245) <= not (a xor b);
    layer0_outputs(5246) <= not b or a;
    layer0_outputs(5247) <= not (a or b);
    layer0_outputs(5248) <= 1'b0;
    layer0_outputs(5249) <= a;
    layer0_outputs(5250) <= 1'b1;
    layer0_outputs(5251) <= not b;
    layer0_outputs(5252) <= a or b;
    layer0_outputs(5253) <= not a;
    layer0_outputs(5254) <= not a;
    layer0_outputs(5255) <= a and b;
    layer0_outputs(5256) <= not a;
    layer0_outputs(5257) <= not a;
    layer0_outputs(5258) <= a or b;
    layer0_outputs(5259) <= a;
    layer0_outputs(5260) <= not b or a;
    layer0_outputs(5261) <= 1'b0;
    layer0_outputs(5262) <= not (a xor b);
    layer0_outputs(5263) <= a and b;
    layer0_outputs(5264) <= a xor b;
    layer0_outputs(5265) <= not a or b;
    layer0_outputs(5266) <= not (a xor b);
    layer0_outputs(5267) <= a and b;
    layer0_outputs(5268) <= not (a xor b);
    layer0_outputs(5269) <= not b;
    layer0_outputs(5270) <= not (a or b);
    layer0_outputs(5271) <= not (a or b);
    layer0_outputs(5272) <= not b;
    layer0_outputs(5273) <= not a;
    layer0_outputs(5274) <= not b or a;
    layer0_outputs(5275) <= a xor b;
    layer0_outputs(5276) <= not (a xor b);
    layer0_outputs(5277) <= b;
    layer0_outputs(5278) <= a or b;
    layer0_outputs(5279) <= a xor b;
    layer0_outputs(5280) <= not (a xor b);
    layer0_outputs(5281) <= a or b;
    layer0_outputs(5282) <= b;
    layer0_outputs(5283) <= 1'b0;
    layer0_outputs(5284) <= b and not a;
    layer0_outputs(5285) <= 1'b0;
    layer0_outputs(5286) <= 1'b0;
    layer0_outputs(5287) <= a;
    layer0_outputs(5288) <= not b;
    layer0_outputs(5289) <= not (a xor b);
    layer0_outputs(5290) <= not a;
    layer0_outputs(5291) <= not b;
    layer0_outputs(5292) <= not b;
    layer0_outputs(5293) <= not a or b;
    layer0_outputs(5294) <= not (a and b);
    layer0_outputs(5295) <= a or b;
    layer0_outputs(5296) <= a and not b;
    layer0_outputs(5297) <= not b;
    layer0_outputs(5298) <= a and not b;
    layer0_outputs(5299) <= a;
    layer0_outputs(5300) <= a;
    layer0_outputs(5301) <= not b;
    layer0_outputs(5302) <= not (a xor b);
    layer0_outputs(5303) <= not a;
    layer0_outputs(5304) <= not a or b;
    layer0_outputs(5305) <= a;
    layer0_outputs(5306) <= 1'b1;
    layer0_outputs(5307) <= a or b;
    layer0_outputs(5308) <= not b or a;
    layer0_outputs(5309) <= not (a and b);
    layer0_outputs(5310) <= a or b;
    layer0_outputs(5311) <= not (a xor b);
    layer0_outputs(5312) <= b and not a;
    layer0_outputs(5313) <= not (a xor b);
    layer0_outputs(5314) <= b and not a;
    layer0_outputs(5315) <= not b;
    layer0_outputs(5316) <= a and b;
    layer0_outputs(5317) <= a and not b;
    layer0_outputs(5318) <= not b or a;
    layer0_outputs(5319) <= b and not a;
    layer0_outputs(5320) <= b and not a;
    layer0_outputs(5321) <= a xor b;
    layer0_outputs(5322) <= 1'b1;
    layer0_outputs(5323) <= a xor b;
    layer0_outputs(5324) <= not a;
    layer0_outputs(5325) <= not (a or b);
    layer0_outputs(5326) <= a;
    layer0_outputs(5327) <= b;
    layer0_outputs(5328) <= not a or b;
    layer0_outputs(5329) <= a and b;
    layer0_outputs(5330) <= b;
    layer0_outputs(5331) <= a and b;
    layer0_outputs(5332) <= a and not b;
    layer0_outputs(5333) <= a xor b;
    layer0_outputs(5334) <= b;
    layer0_outputs(5335) <= a or b;
    layer0_outputs(5336) <= not a or b;
    layer0_outputs(5337) <= a xor b;
    layer0_outputs(5338) <= b;
    layer0_outputs(5339) <= b;
    layer0_outputs(5340) <= 1'b1;
    layer0_outputs(5341) <= not (a xor b);
    layer0_outputs(5342) <= not (a or b);
    layer0_outputs(5343) <= a xor b;
    layer0_outputs(5344) <= b;
    layer0_outputs(5345) <= not a or b;
    layer0_outputs(5346) <= 1'b0;
    layer0_outputs(5347) <= a and not b;
    layer0_outputs(5348) <= a xor b;
    layer0_outputs(5349) <= b and not a;
    layer0_outputs(5350) <= 1'b1;
    layer0_outputs(5351) <= 1'b1;
    layer0_outputs(5352) <= a or b;
    layer0_outputs(5353) <= not (a and b);
    layer0_outputs(5354) <= a xor b;
    layer0_outputs(5355) <= not a or b;
    layer0_outputs(5356) <= a xor b;
    layer0_outputs(5357) <= a;
    layer0_outputs(5358) <= b;
    layer0_outputs(5359) <= not b or a;
    layer0_outputs(5360) <= not a;
    layer0_outputs(5361) <= a;
    layer0_outputs(5362) <= not a or b;
    layer0_outputs(5363) <= not b or a;
    layer0_outputs(5364) <= b and not a;
    layer0_outputs(5365) <= a and b;
    layer0_outputs(5366) <= not b;
    layer0_outputs(5367) <= not (a xor b);
    layer0_outputs(5368) <= not (a xor b);
    layer0_outputs(5369) <= b and not a;
    layer0_outputs(5370) <= b;
    layer0_outputs(5371) <= b;
    layer0_outputs(5372) <= a and not b;
    layer0_outputs(5373) <= a and not b;
    layer0_outputs(5374) <= not (a or b);
    layer0_outputs(5375) <= a and not b;
    layer0_outputs(5376) <= not b or a;
    layer0_outputs(5377) <= not a or b;
    layer0_outputs(5378) <= a or b;
    layer0_outputs(5379) <= not (a xor b);
    layer0_outputs(5380) <= not (a xor b);
    layer0_outputs(5381) <= a xor b;
    layer0_outputs(5382) <= b;
    layer0_outputs(5383) <= not (a or b);
    layer0_outputs(5384) <= not b or a;
    layer0_outputs(5385) <= a and not b;
    layer0_outputs(5386) <= a or b;
    layer0_outputs(5387) <= not (a xor b);
    layer0_outputs(5388) <= not a or b;
    layer0_outputs(5389) <= not b;
    layer0_outputs(5390) <= not b;
    layer0_outputs(5391) <= a or b;
    layer0_outputs(5392) <= a xor b;
    layer0_outputs(5393) <= a;
    layer0_outputs(5394) <= not a;
    layer0_outputs(5395) <= not a or b;
    layer0_outputs(5396) <= not a or b;
    layer0_outputs(5397) <= b and not a;
    layer0_outputs(5398) <= a;
    layer0_outputs(5399) <= a and b;
    layer0_outputs(5400) <= a xor b;
    layer0_outputs(5401) <= not (a or b);
    layer0_outputs(5402) <= not (a xor b);
    layer0_outputs(5403) <= a or b;
    layer0_outputs(5404) <= not b or a;
    layer0_outputs(5405) <= a or b;
    layer0_outputs(5406) <= b and not a;
    layer0_outputs(5407) <= not b;
    layer0_outputs(5408) <= not (a and b);
    layer0_outputs(5409) <= a xor b;
    layer0_outputs(5410) <= not (a xor b);
    layer0_outputs(5411) <= not b;
    layer0_outputs(5412) <= not a or b;
    layer0_outputs(5413) <= b;
    layer0_outputs(5414) <= b;
    layer0_outputs(5415) <= a and b;
    layer0_outputs(5416) <= not (a or b);
    layer0_outputs(5417) <= a and not b;
    layer0_outputs(5418) <= not b or a;
    layer0_outputs(5419) <= a and b;
    layer0_outputs(5420) <= not (a xor b);
    layer0_outputs(5421) <= not (a or b);
    layer0_outputs(5422) <= not (a or b);
    layer0_outputs(5423) <= not b or a;
    layer0_outputs(5424) <= b;
    layer0_outputs(5425) <= not a;
    layer0_outputs(5426) <= a and not b;
    layer0_outputs(5427) <= b;
    layer0_outputs(5428) <= 1'b1;
    layer0_outputs(5429) <= b;
    layer0_outputs(5430) <= not a;
    layer0_outputs(5431) <= b;
    layer0_outputs(5432) <= not a or b;
    layer0_outputs(5433) <= a or b;
    layer0_outputs(5434) <= not (a xor b);
    layer0_outputs(5435) <= 1'b1;
    layer0_outputs(5436) <= not a or b;
    layer0_outputs(5437) <= not (a or b);
    layer0_outputs(5438) <= a and not b;
    layer0_outputs(5439) <= not b;
    layer0_outputs(5440) <= not a;
    layer0_outputs(5441) <= b;
    layer0_outputs(5442) <= 1'b0;
    layer0_outputs(5443) <= b and not a;
    layer0_outputs(5444) <= not a;
    layer0_outputs(5445) <= b and not a;
    layer0_outputs(5446) <= b;
    layer0_outputs(5447) <= not (a or b);
    layer0_outputs(5448) <= not (a xor b);
    layer0_outputs(5449) <= b;
    layer0_outputs(5450) <= b;
    layer0_outputs(5451) <= not b;
    layer0_outputs(5452) <= a xor b;
    layer0_outputs(5453) <= not a or b;
    layer0_outputs(5454) <= not a or b;
    layer0_outputs(5455) <= a or b;
    layer0_outputs(5456) <= a xor b;
    layer0_outputs(5457) <= not (a xor b);
    layer0_outputs(5458) <= a and b;
    layer0_outputs(5459) <= not b;
    layer0_outputs(5460) <= not a or b;
    layer0_outputs(5461) <= 1'b0;
    layer0_outputs(5462) <= not (a or b);
    layer0_outputs(5463) <= a or b;
    layer0_outputs(5464) <= not (a or b);
    layer0_outputs(5465) <= a xor b;
    layer0_outputs(5466) <= not (a or b);
    layer0_outputs(5467) <= not (a or b);
    layer0_outputs(5468) <= not a;
    layer0_outputs(5469) <= not (a or b);
    layer0_outputs(5470) <= a or b;
    layer0_outputs(5471) <= not a;
    layer0_outputs(5472) <= a and not b;
    layer0_outputs(5473) <= not a;
    layer0_outputs(5474) <= a or b;
    layer0_outputs(5475) <= a and b;
    layer0_outputs(5476) <= a;
    layer0_outputs(5477) <= not (a or b);
    layer0_outputs(5478) <= a and not b;
    layer0_outputs(5479) <= a or b;
    layer0_outputs(5480) <= a xor b;
    layer0_outputs(5481) <= not (a xor b);
    layer0_outputs(5482) <= not a;
    layer0_outputs(5483) <= a;
    layer0_outputs(5484) <= b and not a;
    layer0_outputs(5485) <= a;
    layer0_outputs(5486) <= not (a xor b);
    layer0_outputs(5487) <= not b;
    layer0_outputs(5488) <= not a;
    layer0_outputs(5489) <= not a or b;
    layer0_outputs(5490) <= not (a or b);
    layer0_outputs(5491) <= a;
    layer0_outputs(5492) <= 1'b1;
    layer0_outputs(5493) <= not (a or b);
    layer0_outputs(5494) <= a;
    layer0_outputs(5495) <= not a or b;
    layer0_outputs(5496) <= not b;
    layer0_outputs(5497) <= not (a or b);
    layer0_outputs(5498) <= a or b;
    layer0_outputs(5499) <= not (a or b);
    layer0_outputs(5500) <= a;
    layer0_outputs(5501) <= not a or b;
    layer0_outputs(5502) <= a xor b;
    layer0_outputs(5503) <= a xor b;
    layer0_outputs(5504) <= a and not b;
    layer0_outputs(5505) <= not a or b;
    layer0_outputs(5506) <= not a;
    layer0_outputs(5507) <= not (a xor b);
    layer0_outputs(5508) <= b and not a;
    layer0_outputs(5509) <= not b or a;
    layer0_outputs(5510) <= 1'b1;
    layer0_outputs(5511) <= a and b;
    layer0_outputs(5512) <= not b or a;
    layer0_outputs(5513) <= a;
    layer0_outputs(5514) <= a and not b;
    layer0_outputs(5515) <= not a;
    layer0_outputs(5516) <= b and not a;
    layer0_outputs(5517) <= a or b;
    layer0_outputs(5518) <= b and not a;
    layer0_outputs(5519) <= 1'b0;
    layer0_outputs(5520) <= not (a or b);
    layer0_outputs(5521) <= a or b;
    layer0_outputs(5522) <= a;
    layer0_outputs(5523) <= not (a and b);
    layer0_outputs(5524) <= 1'b0;
    layer0_outputs(5525) <= not a or b;
    layer0_outputs(5526) <= not a or b;
    layer0_outputs(5527) <= not (a or b);
    layer0_outputs(5528) <= a;
    layer0_outputs(5529) <= not b or a;
    layer0_outputs(5530) <= a xor b;
    layer0_outputs(5531) <= a or b;
    layer0_outputs(5532) <= a;
    layer0_outputs(5533) <= 1'b0;
    layer0_outputs(5534) <= a or b;
    layer0_outputs(5535) <= 1'b0;
    layer0_outputs(5536) <= not a;
    layer0_outputs(5537) <= b and not a;
    layer0_outputs(5538) <= not (a or b);
    layer0_outputs(5539) <= not b or a;
    layer0_outputs(5540) <= 1'b1;
    layer0_outputs(5541) <= a;
    layer0_outputs(5542) <= a or b;
    layer0_outputs(5543) <= not b or a;
    layer0_outputs(5544) <= not (a xor b);
    layer0_outputs(5545) <= not (a or b);
    layer0_outputs(5546) <= not b;
    layer0_outputs(5547) <= not (a or b);
    layer0_outputs(5548) <= b and not a;
    layer0_outputs(5549) <= a xor b;
    layer0_outputs(5550) <= not a;
    layer0_outputs(5551) <= b;
    layer0_outputs(5552) <= a and not b;
    layer0_outputs(5553) <= a xor b;
    layer0_outputs(5554) <= b;
    layer0_outputs(5555) <= a xor b;
    layer0_outputs(5556) <= a and not b;
    layer0_outputs(5557) <= a xor b;
    layer0_outputs(5558) <= b and not a;
    layer0_outputs(5559) <= not (a or b);
    layer0_outputs(5560) <= b and not a;
    layer0_outputs(5561) <= b;
    layer0_outputs(5562) <= b;
    layer0_outputs(5563) <= a xor b;
    layer0_outputs(5564) <= a;
    layer0_outputs(5565) <= a and b;
    layer0_outputs(5566) <= not (a xor b);
    layer0_outputs(5567) <= not (a xor b);
    layer0_outputs(5568) <= b;
    layer0_outputs(5569) <= a;
    layer0_outputs(5570) <= a and not b;
    layer0_outputs(5571) <= not b or a;
    layer0_outputs(5572) <= a or b;
    layer0_outputs(5573) <= a and b;
    layer0_outputs(5574) <= not b;
    layer0_outputs(5575) <= not a or b;
    layer0_outputs(5576) <= not (a xor b);
    layer0_outputs(5577) <= not a or b;
    layer0_outputs(5578) <= not (a and b);
    layer0_outputs(5579) <= a;
    layer0_outputs(5580) <= not (a and b);
    layer0_outputs(5581) <= not (a or b);
    layer0_outputs(5582) <= not a or b;
    layer0_outputs(5583) <= not b;
    layer0_outputs(5584) <= b;
    layer0_outputs(5585) <= not a;
    layer0_outputs(5586) <= a or b;
    layer0_outputs(5587) <= a and b;
    layer0_outputs(5588) <= not a;
    layer0_outputs(5589) <= a or b;
    layer0_outputs(5590) <= not (a or b);
    layer0_outputs(5591) <= not a;
    layer0_outputs(5592) <= a and not b;
    layer0_outputs(5593) <= not a;
    layer0_outputs(5594) <= a;
    layer0_outputs(5595) <= not a or b;
    layer0_outputs(5596) <= not (a or b);
    layer0_outputs(5597) <= not (a xor b);
    layer0_outputs(5598) <= b and not a;
    layer0_outputs(5599) <= a;
    layer0_outputs(5600) <= a and not b;
    layer0_outputs(5601) <= not b;
    layer0_outputs(5602) <= not b or a;
    layer0_outputs(5603) <= not a;
    layer0_outputs(5604) <= b;
    layer0_outputs(5605) <= 1'b1;
    layer0_outputs(5606) <= b;
    layer0_outputs(5607) <= 1'b1;
    layer0_outputs(5608) <= not b or a;
    layer0_outputs(5609) <= not (a xor b);
    layer0_outputs(5610) <= b;
    layer0_outputs(5611) <= not b;
    layer0_outputs(5612) <= not b;
    layer0_outputs(5613) <= not b or a;
    layer0_outputs(5614) <= 1'b1;
    layer0_outputs(5615) <= a or b;
    layer0_outputs(5616) <= not b;
    layer0_outputs(5617) <= a;
    layer0_outputs(5618) <= a;
    layer0_outputs(5619) <= not (a xor b);
    layer0_outputs(5620) <= b and not a;
    layer0_outputs(5621) <= not (a xor b);
    layer0_outputs(5622) <= a and not b;
    layer0_outputs(5623) <= not (a xor b);
    layer0_outputs(5624) <= not a;
    layer0_outputs(5625) <= not (a xor b);
    layer0_outputs(5626) <= not (a or b);
    layer0_outputs(5627) <= a and not b;
    layer0_outputs(5628) <= b and not a;
    layer0_outputs(5629) <= 1'b0;
    layer0_outputs(5630) <= a and not b;
    layer0_outputs(5631) <= a or b;
    layer0_outputs(5632) <= not (a or b);
    layer0_outputs(5633) <= 1'b1;
    layer0_outputs(5634) <= a xor b;
    layer0_outputs(5635) <= not b;
    layer0_outputs(5636) <= not a;
    layer0_outputs(5637) <= b;
    layer0_outputs(5638) <= not (a xor b);
    layer0_outputs(5639) <= b;
    layer0_outputs(5640) <= b;
    layer0_outputs(5641) <= not a or b;
    layer0_outputs(5642) <= a or b;
    layer0_outputs(5643) <= a xor b;
    layer0_outputs(5644) <= not b;
    layer0_outputs(5645) <= 1'b1;
    layer0_outputs(5646) <= b;
    layer0_outputs(5647) <= not b;
    layer0_outputs(5648) <= b;
    layer0_outputs(5649) <= a;
    layer0_outputs(5650) <= not a or b;
    layer0_outputs(5651) <= a or b;
    layer0_outputs(5652) <= a xor b;
    layer0_outputs(5653) <= not (a or b);
    layer0_outputs(5654) <= a;
    layer0_outputs(5655) <= not (a or b);
    layer0_outputs(5656) <= not b;
    layer0_outputs(5657) <= not (a xor b);
    layer0_outputs(5658) <= not (a or b);
    layer0_outputs(5659) <= not a;
    layer0_outputs(5660) <= b and not a;
    layer0_outputs(5661) <= a;
    layer0_outputs(5662) <= not (a or b);
    layer0_outputs(5663) <= not (a and b);
    layer0_outputs(5664) <= not a;
    layer0_outputs(5665) <= a and not b;
    layer0_outputs(5666) <= not b;
    layer0_outputs(5667) <= not b;
    layer0_outputs(5668) <= not (a and b);
    layer0_outputs(5669) <= not b;
    layer0_outputs(5670) <= not b or a;
    layer0_outputs(5671) <= not b;
    layer0_outputs(5672) <= 1'b1;
    layer0_outputs(5673) <= not (a and b);
    layer0_outputs(5674) <= a xor b;
    layer0_outputs(5675) <= a or b;
    layer0_outputs(5676) <= not (a or b);
    layer0_outputs(5677) <= not (a and b);
    layer0_outputs(5678) <= 1'b0;
    layer0_outputs(5679) <= not b or a;
    layer0_outputs(5680) <= b;
    layer0_outputs(5681) <= 1'b1;
    layer0_outputs(5682) <= b;
    layer0_outputs(5683) <= 1'b0;
    layer0_outputs(5684) <= a;
    layer0_outputs(5685) <= a or b;
    layer0_outputs(5686) <= not a;
    layer0_outputs(5687) <= not b or a;
    layer0_outputs(5688) <= not a or b;
    layer0_outputs(5689) <= a xor b;
    layer0_outputs(5690) <= a or b;
    layer0_outputs(5691) <= not b;
    layer0_outputs(5692) <= a or b;
    layer0_outputs(5693) <= a and b;
    layer0_outputs(5694) <= not (a xor b);
    layer0_outputs(5695) <= 1'b0;
    layer0_outputs(5696) <= not a;
    layer0_outputs(5697) <= a and b;
    layer0_outputs(5698) <= not a or b;
    layer0_outputs(5699) <= not a;
    layer0_outputs(5700) <= not (a xor b);
    layer0_outputs(5701) <= not b;
    layer0_outputs(5702) <= not (a or b);
    layer0_outputs(5703) <= a or b;
    layer0_outputs(5704) <= not (a or b);
    layer0_outputs(5705) <= a;
    layer0_outputs(5706) <= b;
    layer0_outputs(5707) <= not a or b;
    layer0_outputs(5708) <= not (a and b);
    layer0_outputs(5709) <= b and not a;
    layer0_outputs(5710) <= 1'b1;
    layer0_outputs(5711) <= a xor b;
    layer0_outputs(5712) <= not (a or b);
    layer0_outputs(5713) <= not a or b;
    layer0_outputs(5714) <= a or b;
    layer0_outputs(5715) <= b and not a;
    layer0_outputs(5716) <= not (a and b);
    layer0_outputs(5717) <= not b;
    layer0_outputs(5718) <= not (a xor b);
    layer0_outputs(5719) <= not (a or b);
    layer0_outputs(5720) <= not (a xor b);
    layer0_outputs(5721) <= not a or b;
    layer0_outputs(5722) <= 1'b0;
    layer0_outputs(5723) <= not (a xor b);
    layer0_outputs(5724) <= not (a and b);
    layer0_outputs(5725) <= not a;
    layer0_outputs(5726) <= a xor b;
    layer0_outputs(5727) <= 1'b0;
    layer0_outputs(5728) <= not a;
    layer0_outputs(5729) <= 1'b0;
    layer0_outputs(5730) <= a;
    layer0_outputs(5731) <= a or b;
    layer0_outputs(5732) <= not b;
    layer0_outputs(5733) <= a xor b;
    layer0_outputs(5734) <= b;
    layer0_outputs(5735) <= a or b;
    layer0_outputs(5736) <= not b;
    layer0_outputs(5737) <= not (a xor b);
    layer0_outputs(5738) <= not a or b;
    layer0_outputs(5739) <= not a;
    layer0_outputs(5740) <= not a or b;
    layer0_outputs(5741) <= 1'b0;
    layer0_outputs(5742) <= a or b;
    layer0_outputs(5743) <= b and not a;
    layer0_outputs(5744) <= not b or a;
    layer0_outputs(5745) <= a xor b;
    layer0_outputs(5746) <= a and b;
    layer0_outputs(5747) <= 1'b0;
    layer0_outputs(5748) <= a and not b;
    layer0_outputs(5749) <= a;
    layer0_outputs(5750) <= not b;
    layer0_outputs(5751) <= not (a or b);
    layer0_outputs(5752) <= not a or b;
    layer0_outputs(5753) <= a or b;
    layer0_outputs(5754) <= a xor b;
    layer0_outputs(5755) <= a;
    layer0_outputs(5756) <= not b;
    layer0_outputs(5757) <= not (a and b);
    layer0_outputs(5758) <= a;
    layer0_outputs(5759) <= not b;
    layer0_outputs(5760) <= not a or b;
    layer0_outputs(5761) <= not (a and b);
    layer0_outputs(5762) <= a;
    layer0_outputs(5763) <= not (a xor b);
    layer0_outputs(5764) <= a xor b;
    layer0_outputs(5765) <= not a;
    layer0_outputs(5766) <= a;
    layer0_outputs(5767) <= not a or b;
    layer0_outputs(5768) <= not (a and b);
    layer0_outputs(5769) <= not b;
    layer0_outputs(5770) <= not b;
    layer0_outputs(5771) <= a;
    layer0_outputs(5772) <= a;
    layer0_outputs(5773) <= not (a or b);
    layer0_outputs(5774) <= not b;
    layer0_outputs(5775) <= a and not b;
    layer0_outputs(5776) <= a xor b;
    layer0_outputs(5777) <= a xor b;
    layer0_outputs(5778) <= not b;
    layer0_outputs(5779) <= not (a or b);
    layer0_outputs(5780) <= a or b;
    layer0_outputs(5781) <= not b;
    layer0_outputs(5782) <= a;
    layer0_outputs(5783) <= b;
    layer0_outputs(5784) <= not (a or b);
    layer0_outputs(5785) <= not a or b;
    layer0_outputs(5786) <= a;
    layer0_outputs(5787) <= not (a xor b);
    layer0_outputs(5788) <= not b or a;
    layer0_outputs(5789) <= b;
    layer0_outputs(5790) <= not (a and b);
    layer0_outputs(5791) <= a and not b;
    layer0_outputs(5792) <= a;
    layer0_outputs(5793) <= a;
    layer0_outputs(5794) <= not (a or b);
    layer0_outputs(5795) <= not (a or b);
    layer0_outputs(5796) <= a xor b;
    layer0_outputs(5797) <= not (a or b);
    layer0_outputs(5798) <= a or b;
    layer0_outputs(5799) <= not a or b;
    layer0_outputs(5800) <= not a;
    layer0_outputs(5801) <= a or b;
    layer0_outputs(5802) <= a or b;
    layer0_outputs(5803) <= not (a and b);
    layer0_outputs(5804) <= not b;
    layer0_outputs(5805) <= b and not a;
    layer0_outputs(5806) <= a and not b;
    layer0_outputs(5807) <= not (a xor b);
    layer0_outputs(5808) <= not (a xor b);
    layer0_outputs(5809) <= a or b;
    layer0_outputs(5810) <= a;
    layer0_outputs(5811) <= not a or b;
    layer0_outputs(5812) <= b;
    layer0_outputs(5813) <= not b or a;
    layer0_outputs(5814) <= not (a and b);
    layer0_outputs(5815) <= a xor b;
    layer0_outputs(5816) <= a xor b;
    layer0_outputs(5817) <= not (a or b);
    layer0_outputs(5818) <= not b;
    layer0_outputs(5819) <= not (a or b);
    layer0_outputs(5820) <= not (a xor b);
    layer0_outputs(5821) <= 1'b0;
    layer0_outputs(5822) <= 1'b1;
    layer0_outputs(5823) <= not a or b;
    layer0_outputs(5824) <= b;
    layer0_outputs(5825) <= not (a or b);
    layer0_outputs(5826) <= a or b;
    layer0_outputs(5827) <= not b or a;
    layer0_outputs(5828) <= b;
    layer0_outputs(5829) <= a or b;
    layer0_outputs(5830) <= a xor b;
    layer0_outputs(5831) <= not a;
    layer0_outputs(5832) <= b and not a;
    layer0_outputs(5833) <= not b;
    layer0_outputs(5834) <= a or b;
    layer0_outputs(5835) <= a or b;
    layer0_outputs(5836) <= a and not b;
    layer0_outputs(5837) <= 1'b0;
    layer0_outputs(5838) <= a or b;
    layer0_outputs(5839) <= b and not a;
    layer0_outputs(5840) <= a or b;
    layer0_outputs(5841) <= a;
    layer0_outputs(5842) <= a or b;
    layer0_outputs(5843) <= b and not a;
    layer0_outputs(5844) <= a;
    layer0_outputs(5845) <= a;
    layer0_outputs(5846) <= b and not a;
    layer0_outputs(5847) <= not (a xor b);
    layer0_outputs(5848) <= b;
    layer0_outputs(5849) <= a or b;
    layer0_outputs(5850) <= not (a or b);
    layer0_outputs(5851) <= a;
    layer0_outputs(5852) <= 1'b1;
    layer0_outputs(5853) <= a xor b;
    layer0_outputs(5854) <= a or b;
    layer0_outputs(5855) <= not (a or b);
    layer0_outputs(5856) <= not (a or b);
    layer0_outputs(5857) <= not b or a;
    layer0_outputs(5858) <= not (a or b);
    layer0_outputs(5859) <= a and not b;
    layer0_outputs(5860) <= not a;
    layer0_outputs(5861) <= not (a xor b);
    layer0_outputs(5862) <= not a;
    layer0_outputs(5863) <= not b;
    layer0_outputs(5864) <= 1'b1;
    layer0_outputs(5865) <= not b;
    layer0_outputs(5866) <= not a or b;
    layer0_outputs(5867) <= not b or a;
    layer0_outputs(5868) <= not b;
    layer0_outputs(5869) <= not (a xor b);
    layer0_outputs(5870) <= a and not b;
    layer0_outputs(5871) <= not (a or b);
    layer0_outputs(5872) <= a and not b;
    layer0_outputs(5873) <= not b;
    layer0_outputs(5874) <= not a or b;
    layer0_outputs(5875) <= a;
    layer0_outputs(5876) <= not b;
    layer0_outputs(5877) <= b and not a;
    layer0_outputs(5878) <= not a;
    layer0_outputs(5879) <= not b or a;
    layer0_outputs(5880) <= a xor b;
    layer0_outputs(5881) <= not (a xor b);
    layer0_outputs(5882) <= not (a or b);
    layer0_outputs(5883) <= a and not b;
    layer0_outputs(5884) <= a and not b;
    layer0_outputs(5885) <= not (a xor b);
    layer0_outputs(5886) <= a;
    layer0_outputs(5887) <= a and b;
    layer0_outputs(5888) <= a or b;
    layer0_outputs(5889) <= not b;
    layer0_outputs(5890) <= not (a xor b);
    layer0_outputs(5891) <= a and not b;
    layer0_outputs(5892) <= 1'b1;
    layer0_outputs(5893) <= 1'b0;
    layer0_outputs(5894) <= not (a and b);
    layer0_outputs(5895) <= a and not b;
    layer0_outputs(5896) <= a or b;
    layer0_outputs(5897) <= a and not b;
    layer0_outputs(5898) <= a and b;
    layer0_outputs(5899) <= not (a or b);
    layer0_outputs(5900) <= a xor b;
    layer0_outputs(5901) <= a and not b;
    layer0_outputs(5902) <= not (a xor b);
    layer0_outputs(5903) <= a xor b;
    layer0_outputs(5904) <= not b;
    layer0_outputs(5905) <= not (a xor b);
    layer0_outputs(5906) <= a and not b;
    layer0_outputs(5907) <= a or b;
    layer0_outputs(5908) <= a xor b;
    layer0_outputs(5909) <= a and b;
    layer0_outputs(5910) <= a and not b;
    layer0_outputs(5911) <= a;
    layer0_outputs(5912) <= a;
    layer0_outputs(5913) <= b and not a;
    layer0_outputs(5914) <= a xor b;
    layer0_outputs(5915) <= not (a or b);
    layer0_outputs(5916) <= not a or b;
    layer0_outputs(5917) <= not b or a;
    layer0_outputs(5918) <= a xor b;
    layer0_outputs(5919) <= a or b;
    layer0_outputs(5920) <= a or b;
    layer0_outputs(5921) <= a or b;
    layer0_outputs(5922) <= not (a xor b);
    layer0_outputs(5923) <= b;
    layer0_outputs(5924) <= b;
    layer0_outputs(5925) <= a;
    layer0_outputs(5926) <= a and b;
    layer0_outputs(5927) <= a or b;
    layer0_outputs(5928) <= b;
    layer0_outputs(5929) <= a or b;
    layer0_outputs(5930) <= a and not b;
    layer0_outputs(5931) <= a and b;
    layer0_outputs(5932) <= not b or a;
    layer0_outputs(5933) <= not b;
    layer0_outputs(5934) <= not b;
    layer0_outputs(5935) <= not a;
    layer0_outputs(5936) <= a xor b;
    layer0_outputs(5937) <= not b;
    layer0_outputs(5938) <= not (a or b);
    layer0_outputs(5939) <= not (a xor b);
    layer0_outputs(5940) <= 1'b0;
    layer0_outputs(5941) <= not (a or b);
    layer0_outputs(5942) <= not a;
    layer0_outputs(5943) <= b;
    layer0_outputs(5944) <= b and not a;
    layer0_outputs(5945) <= not (a xor b);
    layer0_outputs(5946) <= 1'b1;
    layer0_outputs(5947) <= a;
    layer0_outputs(5948) <= a and not b;
    layer0_outputs(5949) <= 1'b1;
    layer0_outputs(5950) <= b;
    layer0_outputs(5951) <= a;
    layer0_outputs(5952) <= a;
    layer0_outputs(5953) <= b;
    layer0_outputs(5954) <= not a or b;
    layer0_outputs(5955) <= not b;
    layer0_outputs(5956) <= not (a or b);
    layer0_outputs(5957) <= not (a or b);
    layer0_outputs(5958) <= a xor b;
    layer0_outputs(5959) <= not a;
    layer0_outputs(5960) <= not a;
    layer0_outputs(5961) <= b and not a;
    layer0_outputs(5962) <= not (a or b);
    layer0_outputs(5963) <= not a or b;
    layer0_outputs(5964) <= 1'b1;
    layer0_outputs(5965) <= not a;
    layer0_outputs(5966) <= not a;
    layer0_outputs(5967) <= a and not b;
    layer0_outputs(5968) <= not a;
    layer0_outputs(5969) <= 1'b1;
    layer0_outputs(5970) <= not a;
    layer0_outputs(5971) <= not b or a;
    layer0_outputs(5972) <= a or b;
    layer0_outputs(5973) <= not (a or b);
    layer0_outputs(5974) <= not a or b;
    layer0_outputs(5975) <= a and b;
    layer0_outputs(5976) <= b;
    layer0_outputs(5977) <= not a;
    layer0_outputs(5978) <= not (a or b);
    layer0_outputs(5979) <= 1'b0;
    layer0_outputs(5980) <= not a;
    layer0_outputs(5981) <= a and not b;
    layer0_outputs(5982) <= a;
    layer0_outputs(5983) <= not a;
    layer0_outputs(5984) <= a and b;
    layer0_outputs(5985) <= not a or b;
    layer0_outputs(5986) <= 1'b1;
    layer0_outputs(5987) <= not b or a;
    layer0_outputs(5988) <= a or b;
    layer0_outputs(5989) <= not (a or b);
    layer0_outputs(5990) <= a xor b;
    layer0_outputs(5991) <= 1'b0;
    layer0_outputs(5992) <= 1'b0;
    layer0_outputs(5993) <= a and not b;
    layer0_outputs(5994) <= not a or b;
    layer0_outputs(5995) <= 1'b0;
    layer0_outputs(5996) <= not (a xor b);
    layer0_outputs(5997) <= not (a and b);
    layer0_outputs(5998) <= not (a xor b);
    layer0_outputs(5999) <= not a;
    layer0_outputs(6000) <= a or b;
    layer0_outputs(6001) <= a and not b;
    layer0_outputs(6002) <= not b or a;
    layer0_outputs(6003) <= not (a xor b);
    layer0_outputs(6004) <= 1'b1;
    layer0_outputs(6005) <= a and not b;
    layer0_outputs(6006) <= a or b;
    layer0_outputs(6007) <= a and b;
    layer0_outputs(6008) <= b;
    layer0_outputs(6009) <= not b;
    layer0_outputs(6010) <= not b;
    layer0_outputs(6011) <= not (a or b);
    layer0_outputs(6012) <= not (a xor b);
    layer0_outputs(6013) <= a and not b;
    layer0_outputs(6014) <= not (a or b);
    layer0_outputs(6015) <= not a or b;
    layer0_outputs(6016) <= not (a or b);
    layer0_outputs(6017) <= not b or a;
    layer0_outputs(6018) <= not (a or b);
    layer0_outputs(6019) <= a and not b;
    layer0_outputs(6020) <= a;
    layer0_outputs(6021) <= 1'b1;
    layer0_outputs(6022) <= 1'b1;
    layer0_outputs(6023) <= not b;
    layer0_outputs(6024) <= a and not b;
    layer0_outputs(6025) <= b and not a;
    layer0_outputs(6026) <= a or b;
    layer0_outputs(6027) <= a and not b;
    layer0_outputs(6028) <= a or b;
    layer0_outputs(6029) <= not (a xor b);
    layer0_outputs(6030) <= not b or a;
    layer0_outputs(6031) <= not (a or b);
    layer0_outputs(6032) <= not a or b;
    layer0_outputs(6033) <= not (a and b);
    layer0_outputs(6034) <= a or b;
    layer0_outputs(6035) <= not b or a;
    layer0_outputs(6036) <= not b;
    layer0_outputs(6037) <= not b;
    layer0_outputs(6038) <= not (a xor b);
    layer0_outputs(6039) <= a or b;
    layer0_outputs(6040) <= not (a or b);
    layer0_outputs(6041) <= a xor b;
    layer0_outputs(6042) <= a and not b;
    layer0_outputs(6043) <= a;
    layer0_outputs(6044) <= b and not a;
    layer0_outputs(6045) <= not a or b;
    layer0_outputs(6046) <= not a or b;
    layer0_outputs(6047) <= not a or b;
    layer0_outputs(6048) <= not a;
    layer0_outputs(6049) <= a or b;
    layer0_outputs(6050) <= 1'b1;
    layer0_outputs(6051) <= a xor b;
    layer0_outputs(6052) <= a or b;
    layer0_outputs(6053) <= a or b;
    layer0_outputs(6054) <= b;
    layer0_outputs(6055) <= a xor b;
    layer0_outputs(6056) <= not b;
    layer0_outputs(6057) <= not (a or b);
    layer0_outputs(6058) <= a;
    layer0_outputs(6059) <= not a or b;
    layer0_outputs(6060) <= not a;
    layer0_outputs(6061) <= not b or a;
    layer0_outputs(6062) <= a and b;
    layer0_outputs(6063) <= a;
    layer0_outputs(6064) <= a and b;
    layer0_outputs(6065) <= a;
    layer0_outputs(6066) <= not a or b;
    layer0_outputs(6067) <= a;
    layer0_outputs(6068) <= not (a xor b);
    layer0_outputs(6069) <= not a or b;
    layer0_outputs(6070) <= 1'b0;
    layer0_outputs(6071) <= 1'b1;
    layer0_outputs(6072) <= not a;
    layer0_outputs(6073) <= not a or b;
    layer0_outputs(6074) <= not a or b;
    layer0_outputs(6075) <= 1'b1;
    layer0_outputs(6076) <= not b or a;
    layer0_outputs(6077) <= a xor b;
    layer0_outputs(6078) <= a or b;
    layer0_outputs(6079) <= a xor b;
    layer0_outputs(6080) <= b;
    layer0_outputs(6081) <= a and not b;
    layer0_outputs(6082) <= a xor b;
    layer0_outputs(6083) <= not (a or b);
    layer0_outputs(6084) <= not (a xor b);
    layer0_outputs(6085) <= 1'b1;
    layer0_outputs(6086) <= not (a or b);
    layer0_outputs(6087) <= not b or a;
    layer0_outputs(6088) <= not a;
    layer0_outputs(6089) <= a and b;
    layer0_outputs(6090) <= a xor b;
    layer0_outputs(6091) <= not b or a;
    layer0_outputs(6092) <= b;
    layer0_outputs(6093) <= not a or b;
    layer0_outputs(6094) <= not (a or b);
    layer0_outputs(6095) <= not (a or b);
    layer0_outputs(6096) <= 1'b1;
    layer0_outputs(6097) <= not (a xor b);
    layer0_outputs(6098) <= not b;
    layer0_outputs(6099) <= a xor b;
    layer0_outputs(6100) <= not a or b;
    layer0_outputs(6101) <= not b or a;
    layer0_outputs(6102) <= not b or a;
    layer0_outputs(6103) <= b;
    layer0_outputs(6104) <= a;
    layer0_outputs(6105) <= not a or b;
    layer0_outputs(6106) <= b;
    layer0_outputs(6107) <= not b;
    layer0_outputs(6108) <= not a or b;
    layer0_outputs(6109) <= a;
    layer0_outputs(6110) <= not a;
    layer0_outputs(6111) <= not (a or b);
    layer0_outputs(6112) <= b;
    layer0_outputs(6113) <= not (a and b);
    layer0_outputs(6114) <= b;
    layer0_outputs(6115) <= a xor b;
    layer0_outputs(6116) <= not (a or b);
    layer0_outputs(6117) <= a xor b;
    layer0_outputs(6118) <= a;
    layer0_outputs(6119) <= a or b;
    layer0_outputs(6120) <= b;
    layer0_outputs(6121) <= not a;
    layer0_outputs(6122) <= a or b;
    layer0_outputs(6123) <= a xor b;
    layer0_outputs(6124) <= not b or a;
    layer0_outputs(6125) <= a and b;
    layer0_outputs(6126) <= b and not a;
    layer0_outputs(6127) <= b and not a;
    layer0_outputs(6128) <= not b or a;
    layer0_outputs(6129) <= not (a xor b);
    layer0_outputs(6130) <= not (a xor b);
    layer0_outputs(6131) <= a;
    layer0_outputs(6132) <= 1'b1;
    layer0_outputs(6133) <= b;
    layer0_outputs(6134) <= a xor b;
    layer0_outputs(6135) <= a and not b;
    layer0_outputs(6136) <= not b;
    layer0_outputs(6137) <= 1'b1;
    layer0_outputs(6138) <= a;
    layer0_outputs(6139) <= not (a and b);
    layer0_outputs(6140) <= not a or b;
    layer0_outputs(6141) <= a;
    layer0_outputs(6142) <= a or b;
    layer0_outputs(6143) <= a and not b;
    layer0_outputs(6144) <= a and not b;
    layer0_outputs(6145) <= not b;
    layer0_outputs(6146) <= b;
    layer0_outputs(6147) <= a or b;
    layer0_outputs(6148) <= not b;
    layer0_outputs(6149) <= not (a xor b);
    layer0_outputs(6150) <= not b;
    layer0_outputs(6151) <= not a or b;
    layer0_outputs(6152) <= not b;
    layer0_outputs(6153) <= a or b;
    layer0_outputs(6154) <= not (a and b);
    layer0_outputs(6155) <= a xor b;
    layer0_outputs(6156) <= a and not b;
    layer0_outputs(6157) <= a and not b;
    layer0_outputs(6158) <= not (a or b);
    layer0_outputs(6159) <= 1'b0;
    layer0_outputs(6160) <= 1'b0;
    layer0_outputs(6161) <= a and b;
    layer0_outputs(6162) <= not (a or b);
    layer0_outputs(6163) <= not b;
    layer0_outputs(6164) <= a xor b;
    layer0_outputs(6165) <= not b;
    layer0_outputs(6166) <= not a or b;
    layer0_outputs(6167) <= a and not b;
    layer0_outputs(6168) <= not (a or b);
    layer0_outputs(6169) <= not (a or b);
    layer0_outputs(6170) <= a or b;
    layer0_outputs(6171) <= a or b;
    layer0_outputs(6172) <= a and b;
    layer0_outputs(6173) <= not a;
    layer0_outputs(6174) <= a xor b;
    layer0_outputs(6175) <= not a;
    layer0_outputs(6176) <= a and not b;
    layer0_outputs(6177) <= a xor b;
    layer0_outputs(6178) <= not (a or b);
    layer0_outputs(6179) <= a and not b;
    layer0_outputs(6180) <= 1'b0;
    layer0_outputs(6181) <= a or b;
    layer0_outputs(6182) <= a or b;
    layer0_outputs(6183) <= a xor b;
    layer0_outputs(6184) <= a;
    layer0_outputs(6185) <= not a;
    layer0_outputs(6186) <= a xor b;
    layer0_outputs(6187) <= not a;
    layer0_outputs(6188) <= not a or b;
    layer0_outputs(6189) <= not a;
    layer0_outputs(6190) <= b;
    layer0_outputs(6191) <= a and b;
    layer0_outputs(6192) <= not a or b;
    layer0_outputs(6193) <= 1'b0;
    layer0_outputs(6194) <= not a or b;
    layer0_outputs(6195) <= a xor b;
    layer0_outputs(6196) <= not (a xor b);
    layer0_outputs(6197) <= not b or a;
    layer0_outputs(6198) <= not b or a;
    layer0_outputs(6199) <= not (a or b);
    layer0_outputs(6200) <= 1'b0;
    layer0_outputs(6201) <= not (a or b);
    layer0_outputs(6202) <= not (a xor b);
    layer0_outputs(6203) <= b;
    layer0_outputs(6204) <= b;
    layer0_outputs(6205) <= not a or b;
    layer0_outputs(6206) <= b;
    layer0_outputs(6207) <= not (a or b);
    layer0_outputs(6208) <= a;
    layer0_outputs(6209) <= not a;
    layer0_outputs(6210) <= not b;
    layer0_outputs(6211) <= 1'b1;
    layer0_outputs(6212) <= not b or a;
    layer0_outputs(6213) <= b and not a;
    layer0_outputs(6214) <= 1'b1;
    layer0_outputs(6215) <= a;
    layer0_outputs(6216) <= a and not b;
    layer0_outputs(6217) <= not (a or b);
    layer0_outputs(6218) <= 1'b0;
    layer0_outputs(6219) <= not b or a;
    layer0_outputs(6220) <= a or b;
    layer0_outputs(6221) <= 1'b1;
    layer0_outputs(6222) <= not (a or b);
    layer0_outputs(6223) <= not b;
    layer0_outputs(6224) <= not b;
    layer0_outputs(6225) <= not (a xor b);
    layer0_outputs(6226) <= not b;
    layer0_outputs(6227) <= not (a or b);
    layer0_outputs(6228) <= not (a xor b);
    layer0_outputs(6229) <= not (a and b);
    layer0_outputs(6230) <= not (a xor b);
    layer0_outputs(6231) <= a xor b;
    layer0_outputs(6232) <= a xor b;
    layer0_outputs(6233) <= a;
    layer0_outputs(6234) <= a;
    layer0_outputs(6235) <= not (a and b);
    layer0_outputs(6236) <= a;
    layer0_outputs(6237) <= a;
    layer0_outputs(6238) <= not (a or b);
    layer0_outputs(6239) <= a xor b;
    layer0_outputs(6240) <= a or b;
    layer0_outputs(6241) <= a xor b;
    layer0_outputs(6242) <= a and not b;
    layer0_outputs(6243) <= not a or b;
    layer0_outputs(6244) <= a xor b;
    layer0_outputs(6245) <= a;
    layer0_outputs(6246) <= a or b;
    layer0_outputs(6247) <= not (a or b);
    layer0_outputs(6248) <= a xor b;
    layer0_outputs(6249) <= not (a and b);
    layer0_outputs(6250) <= b and not a;
    layer0_outputs(6251) <= a or b;
    layer0_outputs(6252) <= b and not a;
    layer0_outputs(6253) <= a;
    layer0_outputs(6254) <= b and not a;
    layer0_outputs(6255) <= a and not b;
    layer0_outputs(6256) <= not a or b;
    layer0_outputs(6257) <= not a or b;
    layer0_outputs(6258) <= a or b;
    layer0_outputs(6259) <= not (a or b);
    layer0_outputs(6260) <= a and b;
    layer0_outputs(6261) <= a and not b;
    layer0_outputs(6262) <= b;
    layer0_outputs(6263) <= not a;
    layer0_outputs(6264) <= 1'b1;
    layer0_outputs(6265) <= a;
    layer0_outputs(6266) <= not (a or b);
    layer0_outputs(6267) <= a xor b;
    layer0_outputs(6268) <= not b;
    layer0_outputs(6269) <= not b;
    layer0_outputs(6270) <= not a;
    layer0_outputs(6271) <= not (a or b);
    layer0_outputs(6272) <= a xor b;
    layer0_outputs(6273) <= b;
    layer0_outputs(6274) <= not b or a;
    layer0_outputs(6275) <= a and not b;
    layer0_outputs(6276) <= not (a and b);
    layer0_outputs(6277) <= a;
    layer0_outputs(6278) <= not b or a;
    layer0_outputs(6279) <= a xor b;
    layer0_outputs(6280) <= not a or b;
    layer0_outputs(6281) <= a or b;
    layer0_outputs(6282) <= not a or b;
    layer0_outputs(6283) <= not (a or b);
    layer0_outputs(6284) <= not (a or b);
    layer0_outputs(6285) <= b;
    layer0_outputs(6286) <= not a;
    layer0_outputs(6287) <= 1'b0;
    layer0_outputs(6288) <= 1'b0;
    layer0_outputs(6289) <= not (a or b);
    layer0_outputs(6290) <= a and not b;
    layer0_outputs(6291) <= b;
    layer0_outputs(6292) <= not b;
    layer0_outputs(6293) <= a or b;
    layer0_outputs(6294) <= a or b;
    layer0_outputs(6295) <= not b;
    layer0_outputs(6296) <= a or b;
    layer0_outputs(6297) <= a;
    layer0_outputs(6298) <= not b or a;
    layer0_outputs(6299) <= not (a or b);
    layer0_outputs(6300) <= a and b;
    layer0_outputs(6301) <= a and not b;
    layer0_outputs(6302) <= not (a or b);
    layer0_outputs(6303) <= a xor b;
    layer0_outputs(6304) <= not (a or b);
    layer0_outputs(6305) <= not a or b;
    layer0_outputs(6306) <= 1'b0;
    layer0_outputs(6307) <= b and not a;
    layer0_outputs(6308) <= a and not b;
    layer0_outputs(6309) <= a xor b;
    layer0_outputs(6310) <= a and b;
    layer0_outputs(6311) <= a or b;
    layer0_outputs(6312) <= b;
    layer0_outputs(6313) <= a;
    layer0_outputs(6314) <= a or b;
    layer0_outputs(6315) <= a or b;
    layer0_outputs(6316) <= b;
    layer0_outputs(6317) <= not (a or b);
    layer0_outputs(6318) <= a and not b;
    layer0_outputs(6319) <= not (a xor b);
    layer0_outputs(6320) <= b and not a;
    layer0_outputs(6321) <= a or b;
    layer0_outputs(6322) <= b;
    layer0_outputs(6323) <= 1'b0;
    layer0_outputs(6324) <= a xor b;
    layer0_outputs(6325) <= not (a xor b);
    layer0_outputs(6326) <= not (a and b);
    layer0_outputs(6327) <= b and not a;
    layer0_outputs(6328) <= a;
    layer0_outputs(6329) <= a and not b;
    layer0_outputs(6330) <= b;
    layer0_outputs(6331) <= not b or a;
    layer0_outputs(6332) <= a or b;
    layer0_outputs(6333) <= b;
    layer0_outputs(6334) <= not (a and b);
    layer0_outputs(6335) <= not b;
    layer0_outputs(6336) <= not a;
    layer0_outputs(6337) <= b and not a;
    layer0_outputs(6338) <= a or b;
    layer0_outputs(6339) <= not a;
    layer0_outputs(6340) <= b;
    layer0_outputs(6341) <= a and b;
    layer0_outputs(6342) <= b;
    layer0_outputs(6343) <= a and b;
    layer0_outputs(6344) <= a or b;
    layer0_outputs(6345) <= 1'b1;
    layer0_outputs(6346) <= not b or a;
    layer0_outputs(6347) <= a;
    layer0_outputs(6348) <= a xor b;
    layer0_outputs(6349) <= a or b;
    layer0_outputs(6350) <= b and not a;
    layer0_outputs(6351) <= not (a and b);
    layer0_outputs(6352) <= not (a xor b);
    layer0_outputs(6353) <= a xor b;
    layer0_outputs(6354) <= a and b;
    layer0_outputs(6355) <= a or b;
    layer0_outputs(6356) <= a and not b;
    layer0_outputs(6357) <= b and not a;
    layer0_outputs(6358) <= a or b;
    layer0_outputs(6359) <= a and b;
    layer0_outputs(6360) <= a or b;
    layer0_outputs(6361) <= not b;
    layer0_outputs(6362) <= 1'b1;
    layer0_outputs(6363) <= not b or a;
    layer0_outputs(6364) <= a;
    layer0_outputs(6365) <= not (a xor b);
    layer0_outputs(6366) <= not a;
    layer0_outputs(6367) <= b and not a;
    layer0_outputs(6368) <= not (a xor b);
    layer0_outputs(6369) <= not b;
    layer0_outputs(6370) <= not b or a;
    layer0_outputs(6371) <= not b or a;
    layer0_outputs(6372) <= b;
    layer0_outputs(6373) <= b;
    layer0_outputs(6374) <= not (a xor b);
    layer0_outputs(6375) <= a and not b;
    layer0_outputs(6376) <= not b or a;
    layer0_outputs(6377) <= a;
    layer0_outputs(6378) <= not (a and b);
    layer0_outputs(6379) <= a;
    layer0_outputs(6380) <= not (a or b);
    layer0_outputs(6381) <= not a or b;
    layer0_outputs(6382) <= not b;
    layer0_outputs(6383) <= b;
    layer0_outputs(6384) <= a and not b;
    layer0_outputs(6385) <= not a or b;
    layer0_outputs(6386) <= a or b;
    layer0_outputs(6387) <= b;
    layer0_outputs(6388) <= a or b;
    layer0_outputs(6389) <= 1'b1;
    layer0_outputs(6390) <= a xor b;
    layer0_outputs(6391) <= a and b;
    layer0_outputs(6392) <= a xor b;
    layer0_outputs(6393) <= a and not b;
    layer0_outputs(6394) <= not a or b;
    layer0_outputs(6395) <= not b;
    layer0_outputs(6396) <= not b or a;
    layer0_outputs(6397) <= 1'b1;
    layer0_outputs(6398) <= a and not b;
    layer0_outputs(6399) <= not (a or b);
    layer0_outputs(6400) <= a and not b;
    layer0_outputs(6401) <= a or b;
    layer0_outputs(6402) <= a and b;
    layer0_outputs(6403) <= not (a or b);
    layer0_outputs(6404) <= not (a and b);
    layer0_outputs(6405) <= 1'b0;
    layer0_outputs(6406) <= not a;
    layer0_outputs(6407) <= not a or b;
    layer0_outputs(6408) <= b and not a;
    layer0_outputs(6409) <= not (a or b);
    layer0_outputs(6410) <= a and not b;
    layer0_outputs(6411) <= b and not a;
    layer0_outputs(6412) <= a xor b;
    layer0_outputs(6413) <= not b;
    layer0_outputs(6414) <= not a;
    layer0_outputs(6415) <= not a;
    layer0_outputs(6416) <= a or b;
    layer0_outputs(6417) <= a or b;
    layer0_outputs(6418) <= b;
    layer0_outputs(6419) <= not a;
    layer0_outputs(6420) <= a and not b;
    layer0_outputs(6421) <= not b or a;
    layer0_outputs(6422) <= a xor b;
    layer0_outputs(6423) <= not (a or b);
    layer0_outputs(6424) <= a or b;
    layer0_outputs(6425) <= not a;
    layer0_outputs(6426) <= 1'b1;
    layer0_outputs(6427) <= not (a and b);
    layer0_outputs(6428) <= a xor b;
    layer0_outputs(6429) <= b and not a;
    layer0_outputs(6430) <= a;
    layer0_outputs(6431) <= 1'b1;
    layer0_outputs(6432) <= a and not b;
    layer0_outputs(6433) <= a xor b;
    layer0_outputs(6434) <= not (a xor b);
    layer0_outputs(6435) <= not (a or b);
    layer0_outputs(6436) <= not a or b;
    layer0_outputs(6437) <= not a or b;
    layer0_outputs(6438) <= not (a xor b);
    layer0_outputs(6439) <= b and not a;
    layer0_outputs(6440) <= 1'b1;
    layer0_outputs(6441) <= not (a xor b);
    layer0_outputs(6442) <= b;
    layer0_outputs(6443) <= 1'b1;
    layer0_outputs(6444) <= 1'b1;
    layer0_outputs(6445) <= not (a xor b);
    layer0_outputs(6446) <= not (a and b);
    layer0_outputs(6447) <= b and not a;
    layer0_outputs(6448) <= a xor b;
    layer0_outputs(6449) <= not (a or b);
    layer0_outputs(6450) <= 1'b0;
    layer0_outputs(6451) <= not b or a;
    layer0_outputs(6452) <= a or b;
    layer0_outputs(6453) <= a and not b;
    layer0_outputs(6454) <= a xor b;
    layer0_outputs(6455) <= not (a xor b);
    layer0_outputs(6456) <= not (a or b);
    layer0_outputs(6457) <= not (a and b);
    layer0_outputs(6458) <= not a;
    layer0_outputs(6459) <= not a;
    layer0_outputs(6460) <= b and not a;
    layer0_outputs(6461) <= a or b;
    layer0_outputs(6462) <= not (a or b);
    layer0_outputs(6463) <= not a or b;
    layer0_outputs(6464) <= b;
    layer0_outputs(6465) <= a;
    layer0_outputs(6466) <= b;
    layer0_outputs(6467) <= a;
    layer0_outputs(6468) <= not (a or b);
    layer0_outputs(6469) <= not (a or b);
    layer0_outputs(6470) <= not (a or b);
    layer0_outputs(6471) <= not (a xor b);
    layer0_outputs(6472) <= not a;
    layer0_outputs(6473) <= not b;
    layer0_outputs(6474) <= not b;
    layer0_outputs(6475) <= a or b;
    layer0_outputs(6476) <= a and b;
    layer0_outputs(6477) <= not a;
    layer0_outputs(6478) <= b;
    layer0_outputs(6479) <= b;
    layer0_outputs(6480) <= a xor b;
    layer0_outputs(6481) <= a and b;
    layer0_outputs(6482) <= a and b;
    layer0_outputs(6483) <= not (a xor b);
    layer0_outputs(6484) <= not a;
    layer0_outputs(6485) <= a or b;
    layer0_outputs(6486) <= not b or a;
    layer0_outputs(6487) <= not (a xor b);
    layer0_outputs(6488) <= not (a and b);
    layer0_outputs(6489) <= a and not b;
    layer0_outputs(6490) <= not (a or b);
    layer0_outputs(6491) <= b;
    layer0_outputs(6492) <= not a or b;
    layer0_outputs(6493) <= a or b;
    layer0_outputs(6494) <= not (a xor b);
    layer0_outputs(6495) <= a;
    layer0_outputs(6496) <= a;
    layer0_outputs(6497) <= not (a or b);
    layer0_outputs(6498) <= not (a xor b);
    layer0_outputs(6499) <= not (a or b);
    layer0_outputs(6500) <= a;
    layer0_outputs(6501) <= not (a or b);
    layer0_outputs(6502) <= a and not b;
    layer0_outputs(6503) <= not b or a;
    layer0_outputs(6504) <= a or b;
    layer0_outputs(6505) <= a xor b;
    layer0_outputs(6506) <= not (a or b);
    layer0_outputs(6507) <= not (a xor b);
    layer0_outputs(6508) <= not (a or b);
    layer0_outputs(6509) <= not a;
    layer0_outputs(6510) <= a and not b;
    layer0_outputs(6511) <= a or b;
    layer0_outputs(6512) <= a and not b;
    layer0_outputs(6513) <= a or b;
    layer0_outputs(6514) <= a and not b;
    layer0_outputs(6515) <= a xor b;
    layer0_outputs(6516) <= 1'b0;
    layer0_outputs(6517) <= 1'b1;
    layer0_outputs(6518) <= not b or a;
    layer0_outputs(6519) <= 1'b1;
    layer0_outputs(6520) <= not (a xor b);
    layer0_outputs(6521) <= a;
    layer0_outputs(6522) <= b;
    layer0_outputs(6523) <= not (a or b);
    layer0_outputs(6524) <= 1'b0;
    layer0_outputs(6525) <= not a or b;
    layer0_outputs(6526) <= a and not b;
    layer0_outputs(6527) <= not (a and b);
    layer0_outputs(6528) <= not a or b;
    layer0_outputs(6529) <= a;
    layer0_outputs(6530) <= not a;
    layer0_outputs(6531) <= a or b;
    layer0_outputs(6532) <= a or b;
    layer0_outputs(6533) <= a xor b;
    layer0_outputs(6534) <= b and not a;
    layer0_outputs(6535) <= not b;
    layer0_outputs(6536) <= a xor b;
    layer0_outputs(6537) <= a;
    layer0_outputs(6538) <= a xor b;
    layer0_outputs(6539) <= not (a or b);
    layer0_outputs(6540) <= not b;
    layer0_outputs(6541) <= b and not a;
    layer0_outputs(6542) <= b;
    layer0_outputs(6543) <= not a or b;
    layer0_outputs(6544) <= a or b;
    layer0_outputs(6545) <= b;
    layer0_outputs(6546) <= b and not a;
    layer0_outputs(6547) <= not b or a;
    layer0_outputs(6548) <= a;
    layer0_outputs(6549) <= a or b;
    layer0_outputs(6550) <= not (a or b);
    layer0_outputs(6551) <= not (a or b);
    layer0_outputs(6552) <= not b or a;
    layer0_outputs(6553) <= not a;
    layer0_outputs(6554) <= b and not a;
    layer0_outputs(6555) <= a;
    layer0_outputs(6556) <= a xor b;
    layer0_outputs(6557) <= not a;
    layer0_outputs(6558) <= 1'b0;
    layer0_outputs(6559) <= not (a xor b);
    layer0_outputs(6560) <= 1'b1;
    layer0_outputs(6561) <= a;
    layer0_outputs(6562) <= not (a and b);
    layer0_outputs(6563) <= a and b;
    layer0_outputs(6564) <= a and not b;
    layer0_outputs(6565) <= a or b;
    layer0_outputs(6566) <= not a;
    layer0_outputs(6567) <= b and not a;
    layer0_outputs(6568) <= not (a xor b);
    layer0_outputs(6569) <= not b or a;
    layer0_outputs(6570) <= not b;
    layer0_outputs(6571) <= not (a or b);
    layer0_outputs(6572) <= b;
    layer0_outputs(6573) <= not (a or b);
    layer0_outputs(6574) <= a and not b;
    layer0_outputs(6575) <= not b;
    layer0_outputs(6576) <= not a;
    layer0_outputs(6577) <= not a;
    layer0_outputs(6578) <= not (a xor b);
    layer0_outputs(6579) <= not (a xor b);
    layer0_outputs(6580) <= 1'b0;
    layer0_outputs(6581) <= a and not b;
    layer0_outputs(6582) <= not (a or b);
    layer0_outputs(6583) <= 1'b1;
    layer0_outputs(6584) <= not a or b;
    layer0_outputs(6585) <= a;
    layer0_outputs(6586) <= a and b;
    layer0_outputs(6587) <= a and not b;
    layer0_outputs(6588) <= not a or b;
    layer0_outputs(6589) <= a and b;
    layer0_outputs(6590) <= not a;
    layer0_outputs(6591) <= not (a xor b);
    layer0_outputs(6592) <= not (a xor b);
    layer0_outputs(6593) <= a xor b;
    layer0_outputs(6594) <= not a;
    layer0_outputs(6595) <= a;
    layer0_outputs(6596) <= a or b;
    layer0_outputs(6597) <= a and b;
    layer0_outputs(6598) <= 1'b1;
    layer0_outputs(6599) <= not a;
    layer0_outputs(6600) <= a xor b;
    layer0_outputs(6601) <= not a;
    layer0_outputs(6602) <= a;
    layer0_outputs(6603) <= b and not a;
    layer0_outputs(6604) <= not b;
    layer0_outputs(6605) <= a or b;
    layer0_outputs(6606) <= b and not a;
    layer0_outputs(6607) <= a;
    layer0_outputs(6608) <= not b or a;
    layer0_outputs(6609) <= not (a and b);
    layer0_outputs(6610) <= a xor b;
    layer0_outputs(6611) <= b and not a;
    layer0_outputs(6612) <= a xor b;
    layer0_outputs(6613) <= not (a or b);
    layer0_outputs(6614) <= 1'b0;
    layer0_outputs(6615) <= b;
    layer0_outputs(6616) <= 1'b0;
    layer0_outputs(6617) <= a xor b;
    layer0_outputs(6618) <= a;
    layer0_outputs(6619) <= b and not a;
    layer0_outputs(6620) <= not a;
    layer0_outputs(6621) <= a or b;
    layer0_outputs(6622) <= b;
    layer0_outputs(6623) <= not (a xor b);
    layer0_outputs(6624) <= not (a or b);
    layer0_outputs(6625) <= a xor b;
    layer0_outputs(6626) <= a xor b;
    layer0_outputs(6627) <= a or b;
    layer0_outputs(6628) <= b;
    layer0_outputs(6629) <= not (a or b);
    layer0_outputs(6630) <= not (a xor b);
    layer0_outputs(6631) <= not (a or b);
    layer0_outputs(6632) <= a or b;
    layer0_outputs(6633) <= a or b;
    layer0_outputs(6634) <= not a or b;
    layer0_outputs(6635) <= not a;
    layer0_outputs(6636) <= a or b;
    layer0_outputs(6637) <= a xor b;
    layer0_outputs(6638) <= not (a xor b);
    layer0_outputs(6639) <= b;
    layer0_outputs(6640) <= not (a or b);
    layer0_outputs(6641) <= not b;
    layer0_outputs(6642) <= a or b;
    layer0_outputs(6643) <= b;
    layer0_outputs(6644) <= a and not b;
    layer0_outputs(6645) <= a;
    layer0_outputs(6646) <= not (a and b);
    layer0_outputs(6647) <= a xor b;
    layer0_outputs(6648) <= not a or b;
    layer0_outputs(6649) <= a;
    layer0_outputs(6650) <= not a or b;
    layer0_outputs(6651) <= b and not a;
    layer0_outputs(6652) <= not (a or b);
    layer0_outputs(6653) <= not a or b;
    layer0_outputs(6654) <= a;
    layer0_outputs(6655) <= b and not a;
    layer0_outputs(6656) <= a;
    layer0_outputs(6657) <= not (a xor b);
    layer0_outputs(6658) <= 1'b1;
    layer0_outputs(6659) <= b and not a;
    layer0_outputs(6660) <= not (a xor b);
    layer0_outputs(6661) <= not b;
    layer0_outputs(6662) <= b and not a;
    layer0_outputs(6663) <= not (a or b);
    layer0_outputs(6664) <= not b;
    layer0_outputs(6665) <= not a or b;
    layer0_outputs(6666) <= not a;
    layer0_outputs(6667) <= a or b;
    layer0_outputs(6668) <= not b;
    layer0_outputs(6669) <= not a;
    layer0_outputs(6670) <= not a;
    layer0_outputs(6671) <= not (a or b);
    layer0_outputs(6672) <= a xor b;
    layer0_outputs(6673) <= b;
    layer0_outputs(6674) <= a xor b;
    layer0_outputs(6675) <= not b;
    layer0_outputs(6676) <= not a;
    layer0_outputs(6677) <= not (a or b);
    layer0_outputs(6678) <= 1'b0;
    layer0_outputs(6679) <= 1'b0;
    layer0_outputs(6680) <= not (a and b);
    layer0_outputs(6681) <= not a or b;
    layer0_outputs(6682) <= a or b;
    layer0_outputs(6683) <= b;
    layer0_outputs(6684) <= not a;
    layer0_outputs(6685) <= not (a or b);
    layer0_outputs(6686) <= b;
    layer0_outputs(6687) <= b and not a;
    layer0_outputs(6688) <= b and not a;
    layer0_outputs(6689) <= not (a or b);
    layer0_outputs(6690) <= not (a or b);
    layer0_outputs(6691) <= not a;
    layer0_outputs(6692) <= not (a and b);
    layer0_outputs(6693) <= a and not b;
    layer0_outputs(6694) <= not a;
    layer0_outputs(6695) <= a and b;
    layer0_outputs(6696) <= a;
    layer0_outputs(6697) <= not (a or b);
    layer0_outputs(6698) <= not (a xor b);
    layer0_outputs(6699) <= a and b;
    layer0_outputs(6700) <= not (a or b);
    layer0_outputs(6701) <= not b;
    layer0_outputs(6702) <= not b;
    layer0_outputs(6703) <= a and b;
    layer0_outputs(6704) <= not (a and b);
    layer0_outputs(6705) <= 1'b1;
    layer0_outputs(6706) <= a or b;
    layer0_outputs(6707) <= b and not a;
    layer0_outputs(6708) <= not a;
    layer0_outputs(6709) <= a xor b;
    layer0_outputs(6710) <= not (a or b);
    layer0_outputs(6711) <= not b or a;
    layer0_outputs(6712) <= b;
    layer0_outputs(6713) <= not (a xor b);
    layer0_outputs(6714) <= not b or a;
    layer0_outputs(6715) <= a or b;
    layer0_outputs(6716) <= not a or b;
    layer0_outputs(6717) <= not a or b;
    layer0_outputs(6718) <= a or b;
    layer0_outputs(6719) <= a or b;
    layer0_outputs(6720) <= b;
    layer0_outputs(6721) <= not b;
    layer0_outputs(6722) <= a or b;
    layer0_outputs(6723) <= not (a and b);
    layer0_outputs(6724) <= not (a or b);
    layer0_outputs(6725) <= not a or b;
    layer0_outputs(6726) <= not a or b;
    layer0_outputs(6727) <= a;
    layer0_outputs(6728) <= not a;
    layer0_outputs(6729) <= a;
    layer0_outputs(6730) <= 1'b0;
    layer0_outputs(6731) <= not (a or b);
    layer0_outputs(6732) <= b;
    layer0_outputs(6733) <= a and b;
    layer0_outputs(6734) <= b and not a;
    layer0_outputs(6735) <= b;
    layer0_outputs(6736) <= not a or b;
    layer0_outputs(6737) <= 1'b1;
    layer0_outputs(6738) <= b and not a;
    layer0_outputs(6739) <= not (a and b);
    layer0_outputs(6740) <= a xor b;
    layer0_outputs(6741) <= 1'b0;
    layer0_outputs(6742) <= not (a or b);
    layer0_outputs(6743) <= a and b;
    layer0_outputs(6744) <= not (a and b);
    layer0_outputs(6745) <= 1'b1;
    layer0_outputs(6746) <= not (a or b);
    layer0_outputs(6747) <= not (a or b);
    layer0_outputs(6748) <= a or b;
    layer0_outputs(6749) <= a and not b;
    layer0_outputs(6750) <= not b or a;
    layer0_outputs(6751) <= b;
    layer0_outputs(6752) <= not (a or b);
    layer0_outputs(6753) <= a xor b;
    layer0_outputs(6754) <= not (a or b);
    layer0_outputs(6755) <= b and not a;
    layer0_outputs(6756) <= a and not b;
    layer0_outputs(6757) <= not (a or b);
    layer0_outputs(6758) <= not (a or b);
    layer0_outputs(6759) <= not a;
    layer0_outputs(6760) <= not (a xor b);
    layer0_outputs(6761) <= not b or a;
    layer0_outputs(6762) <= b;
    layer0_outputs(6763) <= not a;
    layer0_outputs(6764) <= b;
    layer0_outputs(6765) <= not (a and b);
    layer0_outputs(6766) <= not b or a;
    layer0_outputs(6767) <= not a or b;
    layer0_outputs(6768) <= not a or b;
    layer0_outputs(6769) <= not b;
    layer0_outputs(6770) <= b;
    layer0_outputs(6771) <= a or b;
    layer0_outputs(6772) <= a and not b;
    layer0_outputs(6773) <= 1'b1;
    layer0_outputs(6774) <= not b;
    layer0_outputs(6775) <= not (a or b);
    layer0_outputs(6776) <= not b or a;
    layer0_outputs(6777) <= 1'b0;
    layer0_outputs(6778) <= a;
    layer0_outputs(6779) <= a and b;
    layer0_outputs(6780) <= a;
    layer0_outputs(6781) <= a and not b;
    layer0_outputs(6782) <= 1'b0;
    layer0_outputs(6783) <= a xor b;
    layer0_outputs(6784) <= not b;
    layer0_outputs(6785) <= not (a or b);
    layer0_outputs(6786) <= not (a xor b);
    layer0_outputs(6787) <= a or b;
    layer0_outputs(6788) <= 1'b0;
    layer0_outputs(6789) <= b and not a;
    layer0_outputs(6790) <= a xor b;
    layer0_outputs(6791) <= not a;
    layer0_outputs(6792) <= a xor b;
    layer0_outputs(6793) <= not (a xor b);
    layer0_outputs(6794) <= b and not a;
    layer0_outputs(6795) <= a or b;
    layer0_outputs(6796) <= a xor b;
    layer0_outputs(6797) <= not b;
    layer0_outputs(6798) <= a and not b;
    layer0_outputs(6799) <= a or b;
    layer0_outputs(6800) <= not b or a;
    layer0_outputs(6801) <= a and not b;
    layer0_outputs(6802) <= b and not a;
    layer0_outputs(6803) <= not a or b;
    layer0_outputs(6804) <= not a;
    layer0_outputs(6805) <= not (a xor b);
    layer0_outputs(6806) <= b and not a;
    layer0_outputs(6807) <= a or b;
    layer0_outputs(6808) <= not (a or b);
    layer0_outputs(6809) <= a xor b;
    layer0_outputs(6810) <= a and not b;
    layer0_outputs(6811) <= 1'b0;
    layer0_outputs(6812) <= a xor b;
    layer0_outputs(6813) <= a or b;
    layer0_outputs(6814) <= 1'b0;
    layer0_outputs(6815) <= a or b;
    layer0_outputs(6816) <= b and not a;
    layer0_outputs(6817) <= not a or b;
    layer0_outputs(6818) <= not b or a;
    layer0_outputs(6819) <= not a;
    layer0_outputs(6820) <= a;
    layer0_outputs(6821) <= a and not b;
    layer0_outputs(6822) <= not b;
    layer0_outputs(6823) <= not a;
    layer0_outputs(6824) <= b and not a;
    layer0_outputs(6825) <= a or b;
    layer0_outputs(6826) <= not b or a;
    layer0_outputs(6827) <= a xor b;
    layer0_outputs(6828) <= not (a or b);
    layer0_outputs(6829) <= a and not b;
    layer0_outputs(6830) <= a;
    layer0_outputs(6831) <= not (a or b);
    layer0_outputs(6832) <= a or b;
    layer0_outputs(6833) <= a;
    layer0_outputs(6834) <= not a;
    layer0_outputs(6835) <= a;
    layer0_outputs(6836) <= a and b;
    layer0_outputs(6837) <= not (a or b);
    layer0_outputs(6838) <= not a;
    layer0_outputs(6839) <= a and b;
    layer0_outputs(6840) <= a xor b;
    layer0_outputs(6841) <= not (a xor b);
    layer0_outputs(6842) <= a xor b;
    layer0_outputs(6843) <= not b;
    layer0_outputs(6844) <= not (a or b);
    layer0_outputs(6845) <= not a or b;
    layer0_outputs(6846) <= not b or a;
    layer0_outputs(6847) <= a and not b;
    layer0_outputs(6848) <= not (a xor b);
    layer0_outputs(6849) <= a xor b;
    layer0_outputs(6850) <= not a or b;
    layer0_outputs(6851) <= b and not a;
    layer0_outputs(6852) <= b;
    layer0_outputs(6853) <= not a;
    layer0_outputs(6854) <= b;
    layer0_outputs(6855) <= a and b;
    layer0_outputs(6856) <= not a;
    layer0_outputs(6857) <= not (a xor b);
    layer0_outputs(6858) <= a;
    layer0_outputs(6859) <= b and not a;
    layer0_outputs(6860) <= not (a or b);
    layer0_outputs(6861) <= not a or b;
    layer0_outputs(6862) <= not b;
    layer0_outputs(6863) <= not (a xor b);
    layer0_outputs(6864) <= a or b;
    layer0_outputs(6865) <= a and not b;
    layer0_outputs(6866) <= b;
    layer0_outputs(6867) <= not (a and b);
    layer0_outputs(6868) <= not b or a;
    layer0_outputs(6869) <= not (a xor b);
    layer0_outputs(6870) <= not (a or b);
    layer0_outputs(6871) <= a;
    layer0_outputs(6872) <= not a;
    layer0_outputs(6873) <= not b or a;
    layer0_outputs(6874) <= b;
    layer0_outputs(6875) <= b and not a;
    layer0_outputs(6876) <= a and not b;
    layer0_outputs(6877) <= not a;
    layer0_outputs(6878) <= a or b;
    layer0_outputs(6879) <= not (a or b);
    layer0_outputs(6880) <= b and not a;
    layer0_outputs(6881) <= a xor b;
    layer0_outputs(6882) <= a and not b;
    layer0_outputs(6883) <= a or b;
    layer0_outputs(6884) <= a or b;
    layer0_outputs(6885) <= not b or a;
    layer0_outputs(6886) <= not (a and b);
    layer0_outputs(6887) <= a and not b;
    layer0_outputs(6888) <= not (a or b);
    layer0_outputs(6889) <= not (a and b);
    layer0_outputs(6890) <= not b;
    layer0_outputs(6891) <= not a;
    layer0_outputs(6892) <= b;
    layer0_outputs(6893) <= a;
    layer0_outputs(6894) <= 1'b0;
    layer0_outputs(6895) <= not a or b;
    layer0_outputs(6896) <= a and b;
    layer0_outputs(6897) <= 1'b0;
    layer0_outputs(6898) <= not (a or b);
    layer0_outputs(6899) <= not b;
    layer0_outputs(6900) <= a and b;
    layer0_outputs(6901) <= b;
    layer0_outputs(6902) <= not a or b;
    layer0_outputs(6903) <= not (a xor b);
    layer0_outputs(6904) <= not a;
    layer0_outputs(6905) <= not b or a;
    layer0_outputs(6906) <= not (a or b);
    layer0_outputs(6907) <= not (a xor b);
    layer0_outputs(6908) <= not (a xor b);
    layer0_outputs(6909) <= b;
    layer0_outputs(6910) <= not b or a;
    layer0_outputs(6911) <= not b;
    layer0_outputs(6912) <= a and not b;
    layer0_outputs(6913) <= not b;
    layer0_outputs(6914) <= not (a xor b);
    layer0_outputs(6915) <= not (a xor b);
    layer0_outputs(6916) <= not (a and b);
    layer0_outputs(6917) <= a and b;
    layer0_outputs(6918) <= b and not a;
    layer0_outputs(6919) <= not b;
    layer0_outputs(6920) <= b;
    layer0_outputs(6921) <= not (a xor b);
    layer0_outputs(6922) <= not (a and b);
    layer0_outputs(6923) <= not a;
    layer0_outputs(6924) <= not b or a;
    layer0_outputs(6925) <= b and not a;
    layer0_outputs(6926) <= not (a xor b);
    layer0_outputs(6927) <= a;
    layer0_outputs(6928) <= a or b;
    layer0_outputs(6929) <= not (a or b);
    layer0_outputs(6930) <= not a;
    layer0_outputs(6931) <= not b;
    layer0_outputs(6932) <= not b or a;
    layer0_outputs(6933) <= b and not a;
    layer0_outputs(6934) <= a;
    layer0_outputs(6935) <= a and b;
    layer0_outputs(6936) <= b;
    layer0_outputs(6937) <= a or b;
    layer0_outputs(6938) <= not b;
    layer0_outputs(6939) <= a and b;
    layer0_outputs(6940) <= not (a xor b);
    layer0_outputs(6941) <= not (a or b);
    layer0_outputs(6942) <= not b or a;
    layer0_outputs(6943) <= not b or a;
    layer0_outputs(6944) <= not (a or b);
    layer0_outputs(6945) <= 1'b1;
    layer0_outputs(6946) <= not b or a;
    layer0_outputs(6947) <= b;
    layer0_outputs(6948) <= not a;
    layer0_outputs(6949) <= not b;
    layer0_outputs(6950) <= not b;
    layer0_outputs(6951) <= not (a or b);
    layer0_outputs(6952) <= b and not a;
    layer0_outputs(6953) <= not (a and b);
    layer0_outputs(6954) <= not (a xor b);
    layer0_outputs(6955) <= b and not a;
    layer0_outputs(6956) <= not (a and b);
    layer0_outputs(6957) <= a;
    layer0_outputs(6958) <= b;
    layer0_outputs(6959) <= not a;
    layer0_outputs(6960) <= a or b;
    layer0_outputs(6961) <= 1'b0;
    layer0_outputs(6962) <= not a;
    layer0_outputs(6963) <= not (a xor b);
    layer0_outputs(6964) <= a or b;
    layer0_outputs(6965) <= 1'b1;
    layer0_outputs(6966) <= b and not a;
    layer0_outputs(6967) <= 1'b0;
    layer0_outputs(6968) <= b;
    layer0_outputs(6969) <= 1'b1;
    layer0_outputs(6970) <= not a or b;
    layer0_outputs(6971) <= 1'b0;
    layer0_outputs(6972) <= not b;
    layer0_outputs(6973) <= b;
    layer0_outputs(6974) <= b;
    layer0_outputs(6975) <= a;
    layer0_outputs(6976) <= not a or b;
    layer0_outputs(6977) <= a or b;
    layer0_outputs(6978) <= a or b;
    layer0_outputs(6979) <= not a or b;
    layer0_outputs(6980) <= not (a and b);
    layer0_outputs(6981) <= a or b;
    layer0_outputs(6982) <= not a;
    layer0_outputs(6983) <= 1'b0;
    layer0_outputs(6984) <= a xor b;
    layer0_outputs(6985) <= not (a xor b);
    layer0_outputs(6986) <= not b;
    layer0_outputs(6987) <= not (a or b);
    layer0_outputs(6988) <= not (a or b);
    layer0_outputs(6989) <= not (a or b);
    layer0_outputs(6990) <= not b;
    layer0_outputs(6991) <= not (a xor b);
    layer0_outputs(6992) <= not (a and b);
    layer0_outputs(6993) <= not (a xor b);
    layer0_outputs(6994) <= not b or a;
    layer0_outputs(6995) <= b and not a;
    layer0_outputs(6996) <= a or b;
    layer0_outputs(6997) <= not a;
    layer0_outputs(6998) <= a and not b;
    layer0_outputs(6999) <= not (a or b);
    layer0_outputs(7000) <= a or b;
    layer0_outputs(7001) <= b;
    layer0_outputs(7002) <= a and not b;
    layer0_outputs(7003) <= 1'b0;
    layer0_outputs(7004) <= not b or a;
    layer0_outputs(7005) <= b;
    layer0_outputs(7006) <= not a;
    layer0_outputs(7007) <= a or b;
    layer0_outputs(7008) <= b;
    layer0_outputs(7009) <= a xor b;
    layer0_outputs(7010) <= a xor b;
    layer0_outputs(7011) <= a xor b;
    layer0_outputs(7012) <= not a;
    layer0_outputs(7013) <= a;
    layer0_outputs(7014) <= b and not a;
    layer0_outputs(7015) <= a and b;
    layer0_outputs(7016) <= not (a xor b);
    layer0_outputs(7017) <= not b;
    layer0_outputs(7018) <= a and not b;
    layer0_outputs(7019) <= b;
    layer0_outputs(7020) <= not (a xor b);
    layer0_outputs(7021) <= not a;
    layer0_outputs(7022) <= a or b;
    layer0_outputs(7023) <= b and not a;
    layer0_outputs(7024) <= not (a or b);
    layer0_outputs(7025) <= not a;
    layer0_outputs(7026) <= a or b;
    layer0_outputs(7027) <= a and b;
    layer0_outputs(7028) <= 1'b0;
    layer0_outputs(7029) <= a xor b;
    layer0_outputs(7030) <= not b or a;
    layer0_outputs(7031) <= a xor b;
    layer0_outputs(7032) <= a xor b;
    layer0_outputs(7033) <= a;
    layer0_outputs(7034) <= a and b;
    layer0_outputs(7035) <= b and not a;
    layer0_outputs(7036) <= 1'b0;
    layer0_outputs(7037) <= b;
    layer0_outputs(7038) <= not (a xor b);
    layer0_outputs(7039) <= 1'b0;
    layer0_outputs(7040) <= a and b;
    layer0_outputs(7041) <= a;
    layer0_outputs(7042) <= not b or a;
    layer0_outputs(7043) <= a xor b;
    layer0_outputs(7044) <= a;
    layer0_outputs(7045) <= a and not b;
    layer0_outputs(7046) <= a or b;
    layer0_outputs(7047) <= not a;
    layer0_outputs(7048) <= not b;
    layer0_outputs(7049) <= a;
    layer0_outputs(7050) <= not b or a;
    layer0_outputs(7051) <= b and not a;
    layer0_outputs(7052) <= b;
    layer0_outputs(7053) <= not a;
    layer0_outputs(7054) <= not (a or b);
    layer0_outputs(7055) <= a or b;
    layer0_outputs(7056) <= a and b;
    layer0_outputs(7057) <= not (a or b);
    layer0_outputs(7058) <= b and not a;
    layer0_outputs(7059) <= not (a or b);
    layer0_outputs(7060) <= not (a xor b);
    layer0_outputs(7061) <= not (a or b);
    layer0_outputs(7062) <= not a;
    layer0_outputs(7063) <= not b;
    layer0_outputs(7064) <= not a;
    layer0_outputs(7065) <= not a or b;
    layer0_outputs(7066) <= not (a xor b);
    layer0_outputs(7067) <= a;
    layer0_outputs(7068) <= not (a and b);
    layer0_outputs(7069) <= a or b;
    layer0_outputs(7070) <= a or b;
    layer0_outputs(7071) <= b;
    layer0_outputs(7072) <= a;
    layer0_outputs(7073) <= not (a or b);
    layer0_outputs(7074) <= not b or a;
    layer0_outputs(7075) <= 1'b1;
    layer0_outputs(7076) <= a;
    layer0_outputs(7077) <= a and not b;
    layer0_outputs(7078) <= a and not b;
    layer0_outputs(7079) <= a and not b;
    layer0_outputs(7080) <= a xor b;
    layer0_outputs(7081) <= not (a xor b);
    layer0_outputs(7082) <= not a;
    layer0_outputs(7083) <= a or b;
    layer0_outputs(7084) <= not (a and b);
    layer0_outputs(7085) <= not (a or b);
    layer0_outputs(7086) <= not b;
    layer0_outputs(7087) <= b and not a;
    layer0_outputs(7088) <= 1'b0;
    layer0_outputs(7089) <= not b;
    layer0_outputs(7090) <= not (a or b);
    layer0_outputs(7091) <= a xor b;
    layer0_outputs(7092) <= not b or a;
    layer0_outputs(7093) <= not b or a;
    layer0_outputs(7094) <= a or b;
    layer0_outputs(7095) <= not (a xor b);
    layer0_outputs(7096) <= not a or b;
    layer0_outputs(7097) <= a xor b;
    layer0_outputs(7098) <= b;
    layer0_outputs(7099) <= not b or a;
    layer0_outputs(7100) <= a or b;
    layer0_outputs(7101) <= not (a or b);
    layer0_outputs(7102) <= 1'b1;
    layer0_outputs(7103) <= not a;
    layer0_outputs(7104) <= not b;
    layer0_outputs(7105) <= not a;
    layer0_outputs(7106) <= a and not b;
    layer0_outputs(7107) <= a;
    layer0_outputs(7108) <= not (a or b);
    layer0_outputs(7109) <= not a;
    layer0_outputs(7110) <= not (a xor b);
    layer0_outputs(7111) <= b and not a;
    layer0_outputs(7112) <= a or b;
    layer0_outputs(7113) <= b;
    layer0_outputs(7114) <= a and b;
    layer0_outputs(7115) <= not (a or b);
    layer0_outputs(7116) <= a;
    layer0_outputs(7117) <= b;
    layer0_outputs(7118) <= a;
    layer0_outputs(7119) <= a and not b;
    layer0_outputs(7120) <= not b;
    layer0_outputs(7121) <= b and not a;
    layer0_outputs(7122) <= not (a xor b);
    layer0_outputs(7123) <= a and not b;
    layer0_outputs(7124) <= not (a xor b);
    layer0_outputs(7125) <= b and not a;
    layer0_outputs(7126) <= a or b;
    layer0_outputs(7127) <= not b;
    layer0_outputs(7128) <= not (a xor b);
    layer0_outputs(7129) <= not b or a;
    layer0_outputs(7130) <= 1'b1;
    layer0_outputs(7131) <= not (a xor b);
    layer0_outputs(7132) <= 1'b1;
    layer0_outputs(7133) <= a or b;
    layer0_outputs(7134) <= a;
    layer0_outputs(7135) <= not a;
    layer0_outputs(7136) <= not b;
    layer0_outputs(7137) <= a and not b;
    layer0_outputs(7138) <= a and not b;
    layer0_outputs(7139) <= a or b;
    layer0_outputs(7140) <= 1'b1;
    layer0_outputs(7141) <= not b;
    layer0_outputs(7142) <= a or b;
    layer0_outputs(7143) <= a and not b;
    layer0_outputs(7144) <= a or b;
    layer0_outputs(7145) <= a and b;
    layer0_outputs(7146) <= not a;
    layer0_outputs(7147) <= a and not b;
    layer0_outputs(7148) <= 1'b1;
    layer0_outputs(7149) <= not b;
    layer0_outputs(7150) <= b;
    layer0_outputs(7151) <= not a or b;
    layer0_outputs(7152) <= a;
    layer0_outputs(7153) <= not (a xor b);
    layer0_outputs(7154) <= not b;
    layer0_outputs(7155) <= a and not b;
    layer0_outputs(7156) <= not b or a;
    layer0_outputs(7157) <= not (a and b);
    layer0_outputs(7158) <= a or b;
    layer0_outputs(7159) <= a xor b;
    layer0_outputs(7160) <= not (a xor b);
    layer0_outputs(7161) <= not b;
    layer0_outputs(7162) <= not a or b;
    layer0_outputs(7163) <= 1'b1;
    layer0_outputs(7164) <= a or b;
    layer0_outputs(7165) <= a or b;
    layer0_outputs(7166) <= not (a and b);
    layer0_outputs(7167) <= not a or b;
    layer0_outputs(7168) <= not (a or b);
    layer0_outputs(7169) <= a xor b;
    layer0_outputs(7170) <= not (a or b);
    layer0_outputs(7171) <= a;
    layer0_outputs(7172) <= not b or a;
    layer0_outputs(7173) <= a;
    layer0_outputs(7174) <= not a or b;
    layer0_outputs(7175) <= 1'b1;
    layer0_outputs(7176) <= not a;
    layer0_outputs(7177) <= a;
    layer0_outputs(7178) <= b;
    layer0_outputs(7179) <= 1'b0;
    layer0_outputs(7180) <= not b;
    layer0_outputs(7181) <= 1'b0;
    layer0_outputs(7182) <= b;
    layer0_outputs(7183) <= not (a or b);
    layer0_outputs(7184) <= a;
    layer0_outputs(7185) <= not (a or b);
    layer0_outputs(7186) <= a xor b;
    layer0_outputs(7187) <= not a;
    layer0_outputs(7188) <= not b;
    layer0_outputs(7189) <= 1'b1;
    layer0_outputs(7190) <= not (a or b);
    layer0_outputs(7191) <= not b or a;
    layer0_outputs(7192) <= a;
    layer0_outputs(7193) <= not (a or b);
    layer0_outputs(7194) <= a;
    layer0_outputs(7195) <= a xor b;
    layer0_outputs(7196) <= not a;
    layer0_outputs(7197) <= 1'b1;
    layer0_outputs(7198) <= not b or a;
    layer0_outputs(7199) <= not a;
    layer0_outputs(7200) <= a or b;
    layer0_outputs(7201) <= b and not a;
    layer0_outputs(7202) <= not b;
    layer0_outputs(7203) <= not (a xor b);
    layer0_outputs(7204) <= a or b;
    layer0_outputs(7205) <= a;
    layer0_outputs(7206) <= not b;
    layer0_outputs(7207) <= a or b;
    layer0_outputs(7208) <= 1'b0;
    layer0_outputs(7209) <= a and not b;
    layer0_outputs(7210) <= not (a or b);
    layer0_outputs(7211) <= not b;
    layer0_outputs(7212) <= a or b;
    layer0_outputs(7213) <= a xor b;
    layer0_outputs(7214) <= not a;
    layer0_outputs(7215) <= b and not a;
    layer0_outputs(7216) <= not a;
    layer0_outputs(7217) <= not (a and b);
    layer0_outputs(7218) <= not (a or b);
    layer0_outputs(7219) <= a xor b;
    layer0_outputs(7220) <= not (a or b);
    layer0_outputs(7221) <= 1'b0;
    layer0_outputs(7222) <= 1'b0;
    layer0_outputs(7223) <= a xor b;
    layer0_outputs(7224) <= a;
    layer0_outputs(7225) <= a;
    layer0_outputs(7226) <= a or b;
    layer0_outputs(7227) <= not b;
    layer0_outputs(7228) <= not (a or b);
    layer0_outputs(7229) <= a or b;
    layer0_outputs(7230) <= not (a or b);
    layer0_outputs(7231) <= not a or b;
    layer0_outputs(7232) <= b;
    layer0_outputs(7233) <= not a or b;
    layer0_outputs(7234) <= not (a or b);
    layer0_outputs(7235) <= not b;
    layer0_outputs(7236) <= a and not b;
    layer0_outputs(7237) <= b;
    layer0_outputs(7238) <= a and b;
    layer0_outputs(7239) <= not a;
    layer0_outputs(7240) <= a and b;
    layer0_outputs(7241) <= a and not b;
    layer0_outputs(7242) <= a or b;
    layer0_outputs(7243) <= not a;
    layer0_outputs(7244) <= not a or b;
    layer0_outputs(7245) <= 1'b1;
    layer0_outputs(7246) <= a or b;
    layer0_outputs(7247) <= not (a xor b);
    layer0_outputs(7248) <= not a;
    layer0_outputs(7249) <= not b;
    layer0_outputs(7250) <= not b or a;
    layer0_outputs(7251) <= not (a xor b);
    layer0_outputs(7252) <= a;
    layer0_outputs(7253) <= a;
    layer0_outputs(7254) <= a or b;
    layer0_outputs(7255) <= not (a xor b);
    layer0_outputs(7256) <= not (a and b);
    layer0_outputs(7257) <= b and not a;
    layer0_outputs(7258) <= not (a or b);
    layer0_outputs(7259) <= 1'b1;
    layer0_outputs(7260) <= a;
    layer0_outputs(7261) <= a or b;
    layer0_outputs(7262) <= b and not a;
    layer0_outputs(7263) <= not (a xor b);
    layer0_outputs(7264) <= 1'b0;
    layer0_outputs(7265) <= 1'b1;
    layer0_outputs(7266) <= not (a or b);
    layer0_outputs(7267) <= not (a xor b);
    layer0_outputs(7268) <= b;
    layer0_outputs(7269) <= 1'b0;
    layer0_outputs(7270) <= not b;
    layer0_outputs(7271) <= not (a xor b);
    layer0_outputs(7272) <= a and not b;
    layer0_outputs(7273) <= not a or b;
    layer0_outputs(7274) <= not (a and b);
    layer0_outputs(7275) <= b and not a;
    layer0_outputs(7276) <= not b;
    layer0_outputs(7277) <= a;
    layer0_outputs(7278) <= not (a or b);
    layer0_outputs(7279) <= not (a xor b);
    layer0_outputs(7280) <= not (a or b);
    layer0_outputs(7281) <= a and b;
    layer0_outputs(7282) <= not (a and b);
    layer0_outputs(7283) <= a xor b;
    layer0_outputs(7284) <= not (a or b);
    layer0_outputs(7285) <= not a;
    layer0_outputs(7286) <= not (a or b);
    layer0_outputs(7287) <= not (a and b);
    layer0_outputs(7288) <= not a or b;
    layer0_outputs(7289) <= not b;
    layer0_outputs(7290) <= a and b;
    layer0_outputs(7291) <= 1'b1;
    layer0_outputs(7292) <= not b or a;
    layer0_outputs(7293) <= a and b;
    layer0_outputs(7294) <= not a or b;
    layer0_outputs(7295) <= not (a or b);
    layer0_outputs(7296) <= not a or b;
    layer0_outputs(7297) <= a or b;
    layer0_outputs(7298) <= a;
    layer0_outputs(7299) <= not (a or b);
    layer0_outputs(7300) <= a and not b;
    layer0_outputs(7301) <= not (a xor b);
    layer0_outputs(7302) <= not (a and b);
    layer0_outputs(7303) <= not (a xor b);
    layer0_outputs(7304) <= 1'b1;
    layer0_outputs(7305) <= not a;
    layer0_outputs(7306) <= a;
    layer0_outputs(7307) <= a and b;
    layer0_outputs(7308) <= not (a and b);
    layer0_outputs(7309) <= a or b;
    layer0_outputs(7310) <= not a or b;
    layer0_outputs(7311) <= not b;
    layer0_outputs(7312) <= a;
    layer0_outputs(7313) <= not a or b;
    layer0_outputs(7314) <= a xor b;
    layer0_outputs(7315) <= not a;
    layer0_outputs(7316) <= a or b;
    layer0_outputs(7317) <= b;
    layer0_outputs(7318) <= a;
    layer0_outputs(7319) <= not (a xor b);
    layer0_outputs(7320) <= b;
    layer0_outputs(7321) <= not (a or b);
    layer0_outputs(7322) <= not b;
    layer0_outputs(7323) <= not b or a;
    layer0_outputs(7324) <= b;
    layer0_outputs(7325) <= not (a xor b);
    layer0_outputs(7326) <= a and not b;
    layer0_outputs(7327) <= b;
    layer0_outputs(7328) <= not (a or b);
    layer0_outputs(7329) <= a;
    layer0_outputs(7330) <= a;
    layer0_outputs(7331) <= a and b;
    layer0_outputs(7332) <= not (a or b);
    layer0_outputs(7333) <= b and not a;
    layer0_outputs(7334) <= a and not b;
    layer0_outputs(7335) <= a and not b;
    layer0_outputs(7336) <= not b;
    layer0_outputs(7337) <= b;
    layer0_outputs(7338) <= a and not b;
    layer0_outputs(7339) <= not (a or b);
    layer0_outputs(7340) <= a or b;
    layer0_outputs(7341) <= not b;
    layer0_outputs(7342) <= a;
    layer0_outputs(7343) <= a and not b;
    layer0_outputs(7344) <= a xor b;
    layer0_outputs(7345) <= b and not a;
    layer0_outputs(7346) <= 1'b0;
    layer0_outputs(7347) <= a or b;
    layer0_outputs(7348) <= 1'b0;
    layer0_outputs(7349) <= 1'b0;
    layer0_outputs(7350) <= not (a or b);
    layer0_outputs(7351) <= not a;
    layer0_outputs(7352) <= b and not a;
    layer0_outputs(7353) <= not b;
    layer0_outputs(7354) <= b;
    layer0_outputs(7355) <= a xor b;
    layer0_outputs(7356) <= b and not a;
    layer0_outputs(7357) <= a;
    layer0_outputs(7358) <= not b;
    layer0_outputs(7359) <= not (a and b);
    layer0_outputs(7360) <= a xor b;
    layer0_outputs(7361) <= a or b;
    layer0_outputs(7362) <= not b;
    layer0_outputs(7363) <= not b;
    layer0_outputs(7364) <= not b;
    layer0_outputs(7365) <= not b;
    layer0_outputs(7366) <= a xor b;
    layer0_outputs(7367) <= a or b;
    layer0_outputs(7368) <= not a or b;
    layer0_outputs(7369) <= a;
    layer0_outputs(7370) <= b;
    layer0_outputs(7371) <= not b;
    layer0_outputs(7372) <= not (a or b);
    layer0_outputs(7373) <= not (a xor b);
    layer0_outputs(7374) <= a or b;
    layer0_outputs(7375) <= a or b;
    layer0_outputs(7376) <= not a;
    layer0_outputs(7377) <= not a;
    layer0_outputs(7378) <= not b;
    layer0_outputs(7379) <= a or b;
    layer0_outputs(7380) <= not a;
    layer0_outputs(7381) <= a and b;
    layer0_outputs(7382) <= a and not b;
    layer0_outputs(7383) <= a xor b;
    layer0_outputs(7384) <= not a or b;
    layer0_outputs(7385) <= a or b;
    layer0_outputs(7386) <= b and not a;
    layer0_outputs(7387) <= a xor b;
    layer0_outputs(7388) <= not (a xor b);
    layer0_outputs(7389) <= not (a or b);
    layer0_outputs(7390) <= not b or a;
    layer0_outputs(7391) <= not (a or b);
    layer0_outputs(7392) <= a or b;
    layer0_outputs(7393) <= b;
    layer0_outputs(7394) <= not b;
    layer0_outputs(7395) <= not b;
    layer0_outputs(7396) <= a xor b;
    layer0_outputs(7397) <= not (a or b);
    layer0_outputs(7398) <= not b;
    layer0_outputs(7399) <= not (a or b);
    layer0_outputs(7400) <= not (a and b);
    layer0_outputs(7401) <= not b;
    layer0_outputs(7402) <= b and not a;
    layer0_outputs(7403) <= a and not b;
    layer0_outputs(7404) <= not (a or b);
    layer0_outputs(7405) <= not b;
    layer0_outputs(7406) <= not (a xor b);
    layer0_outputs(7407) <= b;
    layer0_outputs(7408) <= a;
    layer0_outputs(7409) <= not a or b;
    layer0_outputs(7410) <= not a or b;
    layer0_outputs(7411) <= b and not a;
    layer0_outputs(7412) <= not (a or b);
    layer0_outputs(7413) <= not a;
    layer0_outputs(7414) <= a and not b;
    layer0_outputs(7415) <= not (a or b);
    layer0_outputs(7416) <= not (a and b);
    layer0_outputs(7417) <= a and not b;
    layer0_outputs(7418) <= a and b;
    layer0_outputs(7419) <= not b or a;
    layer0_outputs(7420) <= a xor b;
    layer0_outputs(7421) <= not (a and b);
    layer0_outputs(7422) <= not a;
    layer0_outputs(7423) <= a and b;
    layer0_outputs(7424) <= 1'b0;
    layer0_outputs(7425) <= a and b;
    layer0_outputs(7426) <= not a;
    layer0_outputs(7427) <= b and not a;
    layer0_outputs(7428) <= not (a or b);
    layer0_outputs(7429) <= a and not b;
    layer0_outputs(7430) <= not (a xor b);
    layer0_outputs(7431) <= b;
    layer0_outputs(7432) <= not a or b;
    layer0_outputs(7433) <= not (a and b);
    layer0_outputs(7434) <= not (a or b);
    layer0_outputs(7435) <= a and not b;
    layer0_outputs(7436) <= a and not b;
    layer0_outputs(7437) <= b;
    layer0_outputs(7438) <= not a or b;
    layer0_outputs(7439) <= not (a or b);
    layer0_outputs(7440) <= a;
    layer0_outputs(7441) <= 1'b0;
    layer0_outputs(7442) <= not (a xor b);
    layer0_outputs(7443) <= not b;
    layer0_outputs(7444) <= a and not b;
    layer0_outputs(7445) <= not (a xor b);
    layer0_outputs(7446) <= b and not a;
    layer0_outputs(7447) <= not (a xor b);
    layer0_outputs(7448) <= not a or b;
    layer0_outputs(7449) <= not a or b;
    layer0_outputs(7450) <= not b;
    layer0_outputs(7451) <= not a;
    layer0_outputs(7452) <= a and not b;
    layer0_outputs(7453) <= not (a or b);
    layer0_outputs(7454) <= a;
    layer0_outputs(7455) <= b and not a;
    layer0_outputs(7456) <= not (a or b);
    layer0_outputs(7457) <= not (a xor b);
    layer0_outputs(7458) <= not a;
    layer0_outputs(7459) <= not (a and b);
    layer0_outputs(7460) <= a and b;
    layer0_outputs(7461) <= not a;
    layer0_outputs(7462) <= not (a and b);
    layer0_outputs(7463) <= not (a xor b);
    layer0_outputs(7464) <= not b or a;
    layer0_outputs(7465) <= a and not b;
    layer0_outputs(7466) <= not (a and b);
    layer0_outputs(7467) <= not b;
    layer0_outputs(7468) <= b and not a;
    layer0_outputs(7469) <= not b;
    layer0_outputs(7470) <= b;
    layer0_outputs(7471) <= not b;
    layer0_outputs(7472) <= not (a and b);
    layer0_outputs(7473) <= a;
    layer0_outputs(7474) <= 1'b0;
    layer0_outputs(7475) <= not (a and b);
    layer0_outputs(7476) <= a xor b;
    layer0_outputs(7477) <= b and not a;
    layer0_outputs(7478) <= not (a xor b);
    layer0_outputs(7479) <= a or b;
    layer0_outputs(7480) <= not b or a;
    layer0_outputs(7481) <= not a;
    layer0_outputs(7482) <= not (a or b);
    layer0_outputs(7483) <= a and not b;
    layer0_outputs(7484) <= b and not a;
    layer0_outputs(7485) <= b and not a;
    layer0_outputs(7486) <= b and not a;
    layer0_outputs(7487) <= not (a and b);
    layer0_outputs(7488) <= not (a xor b);
    layer0_outputs(7489) <= b;
    layer0_outputs(7490) <= a;
    layer0_outputs(7491) <= not b or a;
    layer0_outputs(7492) <= not a;
    layer0_outputs(7493) <= not b or a;
    layer0_outputs(7494) <= not (a xor b);
    layer0_outputs(7495) <= not a;
    layer0_outputs(7496) <= a and b;
    layer0_outputs(7497) <= a xor b;
    layer0_outputs(7498) <= a and not b;
    layer0_outputs(7499) <= a;
    layer0_outputs(7500) <= a;
    layer0_outputs(7501) <= b and not a;
    layer0_outputs(7502) <= not (a xor b);
    layer0_outputs(7503) <= not (a xor b);
    layer0_outputs(7504) <= a;
    layer0_outputs(7505) <= a xor b;
    layer0_outputs(7506) <= not b;
    layer0_outputs(7507) <= not (a or b);
    layer0_outputs(7508) <= a and not b;
    layer0_outputs(7509) <= a xor b;
    layer0_outputs(7510) <= not a;
    layer0_outputs(7511) <= b;
    layer0_outputs(7512) <= b and not a;
    layer0_outputs(7513) <= a and not b;
    layer0_outputs(7514) <= not (a xor b);
    layer0_outputs(7515) <= a and not b;
    layer0_outputs(7516) <= not (a or b);
    layer0_outputs(7517) <= not (a or b);
    layer0_outputs(7518) <= not (a and b);
    layer0_outputs(7519) <= not a or b;
    layer0_outputs(7520) <= a;
    layer0_outputs(7521) <= b and not a;
    layer0_outputs(7522) <= a and b;
    layer0_outputs(7523) <= not a;
    layer0_outputs(7524) <= a;
    layer0_outputs(7525) <= not a;
    layer0_outputs(7526) <= a or b;
    layer0_outputs(7527) <= a and not b;
    layer0_outputs(7528) <= not b or a;
    layer0_outputs(7529) <= a;
    layer0_outputs(7530) <= 1'b0;
    layer0_outputs(7531) <= b;
    layer0_outputs(7532) <= b and not a;
    layer0_outputs(7533) <= not b or a;
    layer0_outputs(7534) <= a xor b;
    layer0_outputs(7535) <= a and b;
    layer0_outputs(7536) <= a or b;
    layer0_outputs(7537) <= not (a and b);
    layer0_outputs(7538) <= a and not b;
    layer0_outputs(7539) <= not (a or b);
    layer0_outputs(7540) <= not a;
    layer0_outputs(7541) <= not a;
    layer0_outputs(7542) <= a or b;
    layer0_outputs(7543) <= not a or b;
    layer0_outputs(7544) <= b;
    layer0_outputs(7545) <= a xor b;
    layer0_outputs(7546) <= not (a or b);
    layer0_outputs(7547) <= not b or a;
    layer0_outputs(7548) <= not a or b;
    layer0_outputs(7549) <= a and not b;
    layer0_outputs(7550) <= not (a or b);
    layer0_outputs(7551) <= a;
    layer0_outputs(7552) <= b;
    layer0_outputs(7553) <= a and not b;
    layer0_outputs(7554) <= b and not a;
    layer0_outputs(7555) <= a or b;
    layer0_outputs(7556) <= not (a or b);
    layer0_outputs(7557) <= a and not b;
    layer0_outputs(7558) <= a or b;
    layer0_outputs(7559) <= b and not a;
    layer0_outputs(7560) <= not (a xor b);
    layer0_outputs(7561) <= a;
    layer0_outputs(7562) <= not (a xor b);
    layer0_outputs(7563) <= 1'b1;
    layer0_outputs(7564) <= not (a or b);
    layer0_outputs(7565) <= not a or b;
    layer0_outputs(7566) <= a and b;
    layer0_outputs(7567) <= a and b;
    layer0_outputs(7568) <= b and not a;
    layer0_outputs(7569) <= not (a or b);
    layer0_outputs(7570) <= not b or a;
    layer0_outputs(7571) <= not (a xor b);
    layer0_outputs(7572) <= a and b;
    layer0_outputs(7573) <= 1'b1;
    layer0_outputs(7574) <= a;
    layer0_outputs(7575) <= not (a and b);
    layer0_outputs(7576) <= b;
    layer0_outputs(7577) <= a xor b;
    layer0_outputs(7578) <= a xor b;
    layer0_outputs(7579) <= not a or b;
    layer0_outputs(7580) <= b and not a;
    layer0_outputs(7581) <= not a;
    layer0_outputs(7582) <= b;
    layer0_outputs(7583) <= not a;
    layer0_outputs(7584) <= not b;
    layer0_outputs(7585) <= not (a or b);
    layer0_outputs(7586) <= a and not b;
    layer0_outputs(7587) <= not a or b;
    layer0_outputs(7588) <= not a or b;
    layer0_outputs(7589) <= not a;
    layer0_outputs(7590) <= not b or a;
    layer0_outputs(7591) <= not (a or b);
    layer0_outputs(7592) <= a;
    layer0_outputs(7593) <= 1'b1;
    layer0_outputs(7594) <= a xor b;
    layer0_outputs(7595) <= not (a or b);
    layer0_outputs(7596) <= 1'b1;
    layer0_outputs(7597) <= 1'b1;
    layer0_outputs(7598) <= a and b;
    layer0_outputs(7599) <= 1'b1;
    layer0_outputs(7600) <= not a or b;
    layer0_outputs(7601) <= not a or b;
    layer0_outputs(7602) <= not a;
    layer0_outputs(7603) <= a or b;
    layer0_outputs(7604) <= not b;
    layer0_outputs(7605) <= a or b;
    layer0_outputs(7606) <= not (a or b);
    layer0_outputs(7607) <= not b or a;
    layer0_outputs(7608) <= not b;
    layer0_outputs(7609) <= not b;
    layer0_outputs(7610) <= a or b;
    layer0_outputs(7611) <= a and not b;
    layer0_outputs(7612) <= not b;
    layer0_outputs(7613) <= b;
    layer0_outputs(7614) <= not (a or b);
    layer0_outputs(7615) <= not (a xor b);
    layer0_outputs(7616) <= a;
    layer0_outputs(7617) <= not (a or b);
    layer0_outputs(7618) <= a;
    layer0_outputs(7619) <= a and b;
    layer0_outputs(7620) <= not a;
    layer0_outputs(7621) <= not a or b;
    layer0_outputs(7622) <= not (a xor b);
    layer0_outputs(7623) <= b and not a;
    layer0_outputs(7624) <= not (a xor b);
    layer0_outputs(7625) <= 1'b1;
    layer0_outputs(7626) <= not a or b;
    layer0_outputs(7627) <= not (a or b);
    layer0_outputs(7628) <= a;
    layer0_outputs(7629) <= not (a xor b);
    layer0_outputs(7630) <= a xor b;
    layer0_outputs(7631) <= not a or b;
    layer0_outputs(7632) <= not (a and b);
    layer0_outputs(7633) <= not a or b;
    layer0_outputs(7634) <= a and b;
    layer0_outputs(7635) <= a;
    layer0_outputs(7636) <= not (a or b);
    layer0_outputs(7637) <= not a;
    layer0_outputs(7638) <= not a;
    layer0_outputs(7639) <= not a;
    layer0_outputs(7640) <= b and not a;
    layer0_outputs(7641) <= a xor b;
    layer0_outputs(7642) <= 1'b1;
    layer0_outputs(7643) <= a and not b;
    layer0_outputs(7644) <= a and b;
    layer0_outputs(7645) <= a;
    layer0_outputs(7646) <= b;
    layer0_outputs(7647) <= not b;
    layer0_outputs(7648) <= b;
    layer0_outputs(7649) <= 1'b0;
    layer0_outputs(7650) <= a or b;
    layer0_outputs(7651) <= not a;
    layer0_outputs(7652) <= b and not a;
    layer0_outputs(7653) <= b and not a;
    layer0_outputs(7654) <= not b or a;
    layer0_outputs(7655) <= not b or a;
    layer0_outputs(7656) <= 1'b0;
    layer0_outputs(7657) <= b;
    layer0_outputs(7658) <= not a or b;
    layer0_outputs(7659) <= a and not b;
    layer0_outputs(7660) <= not (a or b);
    layer0_outputs(7661) <= not (a xor b);
    layer0_outputs(7662) <= not b;
    layer0_outputs(7663) <= a or b;
    layer0_outputs(7664) <= not a;
    layer0_outputs(7665) <= not b;
    layer0_outputs(7666) <= a and not b;
    layer0_outputs(7667) <= not (a and b);
    layer0_outputs(7668) <= a and not b;
    layer0_outputs(7669) <= b and not a;
    layer0_outputs(7670) <= 1'b0;
    layer0_outputs(7671) <= a or b;
    layer0_outputs(7672) <= a or b;
    layer0_outputs(7673) <= not b or a;
    layer0_outputs(7674) <= not a or b;
    layer0_outputs(7675) <= not a or b;
    layer0_outputs(7676) <= a and not b;
    layer0_outputs(7677) <= b;
    layer0_outputs(7678) <= b and not a;
    layer0_outputs(7679) <= a or b;
    layer0_outputs(7680) <= b and not a;
    layer0_outputs(7681) <= not b or a;
    layer0_outputs(7682) <= not b;
    layer0_outputs(7683) <= 1'b0;
    layer0_outputs(7684) <= not b or a;
    layer0_outputs(7685) <= not a or b;
    layer0_outputs(7686) <= not (a or b);
    layer0_outputs(7687) <= b and not a;
    layer0_outputs(7688) <= not b or a;
    layer0_outputs(7689) <= b and not a;
    layer0_outputs(7690) <= 1'b0;
    layer0_outputs(7691) <= a and not b;
    layer0_outputs(7692) <= b;
    layer0_outputs(7693) <= not (a xor b);
    layer0_outputs(7694) <= not a or b;
    layer0_outputs(7695) <= not a;
    layer0_outputs(7696) <= not (a xor b);
    layer0_outputs(7697) <= a or b;
    layer0_outputs(7698) <= not (a xor b);
    layer0_outputs(7699) <= not (a xor b);
    layer0_outputs(7700) <= b and not a;
    layer0_outputs(7701) <= a and not b;
    layer0_outputs(7702) <= a and b;
    layer0_outputs(7703) <= 1'b0;
    layer0_outputs(7704) <= not a;
    layer0_outputs(7705) <= not a;
    layer0_outputs(7706) <= b and not a;
    layer0_outputs(7707) <= a xor b;
    layer0_outputs(7708) <= b;
    layer0_outputs(7709) <= a;
    layer0_outputs(7710) <= a;
    layer0_outputs(7711) <= not a or b;
    layer0_outputs(7712) <= b;
    layer0_outputs(7713) <= a or b;
    layer0_outputs(7714) <= a;
    layer0_outputs(7715) <= b;
    layer0_outputs(7716) <= a;
    layer0_outputs(7717) <= 1'b0;
    layer0_outputs(7718) <= b and not a;
    layer0_outputs(7719) <= a;
    layer0_outputs(7720) <= a xor b;
    layer0_outputs(7721) <= not b;
    layer0_outputs(7722) <= not (a or b);
    layer0_outputs(7723) <= not (a or b);
    layer0_outputs(7724) <= not a or b;
    layer0_outputs(7725) <= 1'b1;
    layer0_outputs(7726) <= 1'b0;
    layer0_outputs(7727) <= not (a or b);
    layer0_outputs(7728) <= a or b;
    layer0_outputs(7729) <= a or b;
    layer0_outputs(7730) <= 1'b1;
    layer0_outputs(7731) <= a or b;
    layer0_outputs(7732) <= not b or a;
    layer0_outputs(7733) <= not (a xor b);
    layer0_outputs(7734) <= b and not a;
    layer0_outputs(7735) <= a;
    layer0_outputs(7736) <= a or b;
    layer0_outputs(7737) <= not (a and b);
    layer0_outputs(7738) <= not (a xor b);
    layer0_outputs(7739) <= a and b;
    layer0_outputs(7740) <= b and not a;
    layer0_outputs(7741) <= a and b;
    layer0_outputs(7742) <= not a or b;
    layer0_outputs(7743) <= not (a or b);
    layer0_outputs(7744) <= b;
    layer0_outputs(7745) <= a;
    layer0_outputs(7746) <= not (a and b);
    layer0_outputs(7747) <= not b or a;
    layer0_outputs(7748) <= a or b;
    layer0_outputs(7749) <= not (a xor b);
    layer0_outputs(7750) <= a xor b;
    layer0_outputs(7751) <= not b;
    layer0_outputs(7752) <= a xor b;
    layer0_outputs(7753) <= not b;
    layer0_outputs(7754) <= b and not a;
    layer0_outputs(7755) <= not b or a;
    layer0_outputs(7756) <= not a or b;
    layer0_outputs(7757) <= not a or b;
    layer0_outputs(7758) <= a and b;
    layer0_outputs(7759) <= a xor b;
    layer0_outputs(7760) <= not b or a;
    layer0_outputs(7761) <= 1'b1;
    layer0_outputs(7762) <= a and b;
    layer0_outputs(7763) <= 1'b1;
    layer0_outputs(7764) <= 1'b1;
    layer0_outputs(7765) <= a;
    layer0_outputs(7766) <= b;
    layer0_outputs(7767) <= a or b;
    layer0_outputs(7768) <= 1'b1;
    layer0_outputs(7769) <= not (a xor b);
    layer0_outputs(7770) <= not a;
    layer0_outputs(7771) <= not a or b;
    layer0_outputs(7772) <= not b or a;
    layer0_outputs(7773) <= a or b;
    layer0_outputs(7774) <= b;
    layer0_outputs(7775) <= 1'b0;
    layer0_outputs(7776) <= not a;
    layer0_outputs(7777) <= a and not b;
    layer0_outputs(7778) <= a or b;
    layer0_outputs(7779) <= a and b;
    layer0_outputs(7780) <= not a;
    layer0_outputs(7781) <= a;
    layer0_outputs(7782) <= not (a or b);
    layer0_outputs(7783) <= not (a or b);
    layer0_outputs(7784) <= not b;
    layer0_outputs(7785) <= not (a and b);
    layer0_outputs(7786) <= b and not a;
    layer0_outputs(7787) <= not a;
    layer0_outputs(7788) <= not b or a;
    layer0_outputs(7789) <= a or b;
    layer0_outputs(7790) <= not a or b;
    layer0_outputs(7791) <= b;
    layer0_outputs(7792) <= a;
    layer0_outputs(7793) <= a;
    layer0_outputs(7794) <= b;
    layer0_outputs(7795) <= a and not b;
    layer0_outputs(7796) <= not a or b;
    layer0_outputs(7797) <= b and not a;
    layer0_outputs(7798) <= not b or a;
    layer0_outputs(7799) <= b and not a;
    layer0_outputs(7800) <= a or b;
    layer0_outputs(7801) <= a or b;
    layer0_outputs(7802) <= not b;
    layer0_outputs(7803) <= b and not a;
    layer0_outputs(7804) <= 1'b1;
    layer0_outputs(7805) <= a and not b;
    layer0_outputs(7806) <= a xor b;
    layer0_outputs(7807) <= b;
    layer0_outputs(7808) <= b;
    layer0_outputs(7809) <= 1'b1;
    layer0_outputs(7810) <= not b or a;
    layer0_outputs(7811) <= a and not b;
    layer0_outputs(7812) <= 1'b0;
    layer0_outputs(7813) <= a;
    layer0_outputs(7814) <= not (a or b);
    layer0_outputs(7815) <= b and not a;
    layer0_outputs(7816) <= not a or b;
    layer0_outputs(7817) <= a;
    layer0_outputs(7818) <= not (a and b);
    layer0_outputs(7819) <= not b or a;
    layer0_outputs(7820) <= not a or b;
    layer0_outputs(7821) <= a xor b;
    layer0_outputs(7822) <= b and not a;
    layer0_outputs(7823) <= a;
    layer0_outputs(7824) <= a;
    layer0_outputs(7825) <= not b;
    layer0_outputs(7826) <= not b or a;
    layer0_outputs(7827) <= a and not b;
    layer0_outputs(7828) <= a or b;
    layer0_outputs(7829) <= b and not a;
    layer0_outputs(7830) <= a;
    layer0_outputs(7831) <= not (a or b);
    layer0_outputs(7832) <= not (a xor b);
    layer0_outputs(7833) <= not (a xor b);
    layer0_outputs(7834) <= not (a and b);
    layer0_outputs(7835) <= a and b;
    layer0_outputs(7836) <= a or b;
    layer0_outputs(7837) <= a and b;
    layer0_outputs(7838) <= not a or b;
    layer0_outputs(7839) <= a and not b;
    layer0_outputs(7840) <= not a;
    layer0_outputs(7841) <= b and not a;
    layer0_outputs(7842) <= a or b;
    layer0_outputs(7843) <= not b or a;
    layer0_outputs(7844) <= b and not a;
    layer0_outputs(7845) <= a;
    layer0_outputs(7846) <= not (a or b);
    layer0_outputs(7847) <= not a or b;
    layer0_outputs(7848) <= not b;
    layer0_outputs(7849) <= not a or b;
    layer0_outputs(7850) <= not (a or b);
    layer0_outputs(7851) <= not a or b;
    layer0_outputs(7852) <= not b;
    layer0_outputs(7853) <= 1'b1;
    layer0_outputs(7854) <= not (a and b);
    layer0_outputs(7855) <= not b;
    layer0_outputs(7856) <= not b;
    layer0_outputs(7857) <= b;
    layer0_outputs(7858) <= a and not b;
    layer0_outputs(7859) <= not b;
    layer0_outputs(7860) <= not b;
    layer0_outputs(7861) <= not (a or b);
    layer0_outputs(7862) <= b and not a;
    layer0_outputs(7863) <= not b or a;
    layer0_outputs(7864) <= a;
    layer0_outputs(7865) <= not a;
    layer0_outputs(7866) <= not (a and b);
    layer0_outputs(7867) <= a and not b;
    layer0_outputs(7868) <= b and not a;
    layer0_outputs(7869) <= not b;
    layer0_outputs(7870) <= not b or a;
    layer0_outputs(7871) <= not b or a;
    layer0_outputs(7872) <= a and b;
    layer0_outputs(7873) <= not b or a;
    layer0_outputs(7874) <= not (a and b);
    layer0_outputs(7875) <= a and not b;
    layer0_outputs(7876) <= not b or a;
    layer0_outputs(7877) <= a or b;
    layer0_outputs(7878) <= not (a or b);
    layer0_outputs(7879) <= a or b;
    layer0_outputs(7880) <= a and not b;
    layer0_outputs(7881) <= a and b;
    layer0_outputs(7882) <= a and not b;
    layer0_outputs(7883) <= not a;
    layer0_outputs(7884) <= a or b;
    layer0_outputs(7885) <= b and not a;
    layer0_outputs(7886) <= not (a xor b);
    layer0_outputs(7887) <= not a;
    layer0_outputs(7888) <= b;
    layer0_outputs(7889) <= not b;
    layer0_outputs(7890) <= not (a or b);
    layer0_outputs(7891) <= a or b;
    layer0_outputs(7892) <= a or b;
    layer0_outputs(7893) <= not (a and b);
    layer0_outputs(7894) <= a and b;
    layer0_outputs(7895) <= not (a or b);
    layer0_outputs(7896) <= not a;
    layer0_outputs(7897) <= not (a and b);
    layer0_outputs(7898) <= not a;
    layer0_outputs(7899) <= b;
    layer0_outputs(7900) <= not b or a;
    layer0_outputs(7901) <= a or b;
    layer0_outputs(7902) <= not a;
    layer0_outputs(7903) <= a;
    layer0_outputs(7904) <= a xor b;
    layer0_outputs(7905) <= a;
    layer0_outputs(7906) <= b and not a;
    layer0_outputs(7907) <= 1'b1;
    layer0_outputs(7908) <= not (a or b);
    layer0_outputs(7909) <= not a;
    layer0_outputs(7910) <= b;
    layer0_outputs(7911) <= not b;
    layer0_outputs(7912) <= a xor b;
    layer0_outputs(7913) <= a and b;
    layer0_outputs(7914) <= b;
    layer0_outputs(7915) <= not b or a;
    layer0_outputs(7916) <= 1'b0;
    layer0_outputs(7917) <= not a or b;
    layer0_outputs(7918) <= not (a or b);
    layer0_outputs(7919) <= not (a xor b);
    layer0_outputs(7920) <= not b or a;
    layer0_outputs(7921) <= not (a or b);
    layer0_outputs(7922) <= b;
    layer0_outputs(7923) <= not (a or b);
    layer0_outputs(7924) <= a and b;
    layer0_outputs(7925) <= a and b;
    layer0_outputs(7926) <= a and not b;
    layer0_outputs(7927) <= not (a or b);
    layer0_outputs(7928) <= not a or b;
    layer0_outputs(7929) <= a xor b;
    layer0_outputs(7930) <= b and not a;
    layer0_outputs(7931) <= not (a or b);
    layer0_outputs(7932) <= a;
    layer0_outputs(7933) <= a xor b;
    layer0_outputs(7934) <= not (a or b);
    layer0_outputs(7935) <= not b or a;
    layer0_outputs(7936) <= not b or a;
    layer0_outputs(7937) <= a or b;
    layer0_outputs(7938) <= a;
    layer0_outputs(7939) <= b;
    layer0_outputs(7940) <= not (a and b);
    layer0_outputs(7941) <= not (a or b);
    layer0_outputs(7942) <= not b;
    layer0_outputs(7943) <= not a or b;
    layer0_outputs(7944) <= a or b;
    layer0_outputs(7945) <= b and not a;
    layer0_outputs(7946) <= not a or b;
    layer0_outputs(7947) <= a;
    layer0_outputs(7948) <= b;
    layer0_outputs(7949) <= not a or b;
    layer0_outputs(7950) <= not (a or b);
    layer0_outputs(7951) <= not b;
    layer0_outputs(7952) <= not (a xor b);
    layer0_outputs(7953) <= a;
    layer0_outputs(7954) <= a or b;
    layer0_outputs(7955) <= b;
    layer0_outputs(7956) <= not b or a;
    layer0_outputs(7957) <= a or b;
    layer0_outputs(7958) <= b;
    layer0_outputs(7959) <= b and not a;
    layer0_outputs(7960) <= not b or a;
    layer0_outputs(7961) <= not b or a;
    layer0_outputs(7962) <= a xor b;
    layer0_outputs(7963) <= not b;
    layer0_outputs(7964) <= a and b;
    layer0_outputs(7965) <= b;
    layer0_outputs(7966) <= b;
    layer0_outputs(7967) <= 1'b1;
    layer0_outputs(7968) <= not b or a;
    layer0_outputs(7969) <= 1'b1;
    layer0_outputs(7970) <= a xor b;
    layer0_outputs(7971) <= not (a xor b);
    layer0_outputs(7972) <= 1'b1;
    layer0_outputs(7973) <= not a;
    layer0_outputs(7974) <= b and not a;
    layer0_outputs(7975) <= a;
    layer0_outputs(7976) <= not (a or b);
    layer0_outputs(7977) <= a and not b;
    layer0_outputs(7978) <= a;
    layer0_outputs(7979) <= not (a or b);
    layer0_outputs(7980) <= a;
    layer0_outputs(7981) <= b;
    layer0_outputs(7982) <= 1'b0;
    layer0_outputs(7983) <= not a;
    layer0_outputs(7984) <= b;
    layer0_outputs(7985) <= not (a or b);
    layer0_outputs(7986) <= 1'b1;
    layer0_outputs(7987) <= not b;
    layer0_outputs(7988) <= not (a or b);
    layer0_outputs(7989) <= not a;
    layer0_outputs(7990) <= not a or b;
    layer0_outputs(7991) <= not (a xor b);
    layer0_outputs(7992) <= not (a or b);
    layer0_outputs(7993) <= b;
    layer0_outputs(7994) <= not (a xor b);
    layer0_outputs(7995) <= not (a xor b);
    layer0_outputs(7996) <= a;
    layer0_outputs(7997) <= a and not b;
    layer0_outputs(7998) <= not (a xor b);
    layer0_outputs(7999) <= a or b;
    layer0_outputs(8000) <= a or b;
    layer0_outputs(8001) <= 1'b0;
    layer0_outputs(8002) <= not (a xor b);
    layer0_outputs(8003) <= not (a or b);
    layer0_outputs(8004) <= not b or a;
    layer0_outputs(8005) <= a or b;
    layer0_outputs(8006) <= a and not b;
    layer0_outputs(8007) <= a and b;
    layer0_outputs(8008) <= not b or a;
    layer0_outputs(8009) <= not (a xor b);
    layer0_outputs(8010) <= a and b;
    layer0_outputs(8011) <= not (a xor b);
    layer0_outputs(8012) <= a or b;
    layer0_outputs(8013) <= not a;
    layer0_outputs(8014) <= a xor b;
    layer0_outputs(8015) <= a and not b;
    layer0_outputs(8016) <= a or b;
    layer0_outputs(8017) <= 1'b1;
    layer0_outputs(8018) <= not a or b;
    layer0_outputs(8019) <= 1'b1;
    layer0_outputs(8020) <= 1'b1;
    layer0_outputs(8021) <= not (a xor b);
    layer0_outputs(8022) <= not b or a;
    layer0_outputs(8023) <= not a or b;
    layer0_outputs(8024) <= not a;
    layer0_outputs(8025) <= 1'b0;
    layer0_outputs(8026) <= not a or b;
    layer0_outputs(8027) <= a or b;
    layer0_outputs(8028) <= 1'b1;
    layer0_outputs(8029) <= a;
    layer0_outputs(8030) <= b and not a;
    layer0_outputs(8031) <= not b or a;
    layer0_outputs(8032) <= a;
    layer0_outputs(8033) <= b;
    layer0_outputs(8034) <= not b;
    layer0_outputs(8035) <= a;
    layer0_outputs(8036) <= not (a and b);
    layer0_outputs(8037) <= not (a or b);
    layer0_outputs(8038) <= a xor b;
    layer0_outputs(8039) <= a and b;
    layer0_outputs(8040) <= a xor b;
    layer0_outputs(8041) <= a or b;
    layer0_outputs(8042) <= not b or a;
    layer0_outputs(8043) <= not (a and b);
    layer0_outputs(8044) <= a;
    layer0_outputs(8045) <= b;
    layer0_outputs(8046) <= 1'b0;
    layer0_outputs(8047) <= a and not b;
    layer0_outputs(8048) <= b;
    layer0_outputs(8049) <= not a or b;
    layer0_outputs(8050) <= a;
    layer0_outputs(8051) <= not b or a;
    layer0_outputs(8052) <= not a;
    layer0_outputs(8053) <= not (a or b);
    layer0_outputs(8054) <= not a;
    layer0_outputs(8055) <= 1'b0;
    layer0_outputs(8056) <= b and not a;
    layer0_outputs(8057) <= a and b;
    layer0_outputs(8058) <= a or b;
    layer0_outputs(8059) <= not b;
    layer0_outputs(8060) <= a;
    layer0_outputs(8061) <= not b;
    layer0_outputs(8062) <= 1'b0;
    layer0_outputs(8063) <= a and not b;
    layer0_outputs(8064) <= a;
    layer0_outputs(8065) <= not a;
    layer0_outputs(8066) <= a and not b;
    layer0_outputs(8067) <= b and not a;
    layer0_outputs(8068) <= not a;
    layer0_outputs(8069) <= not a;
    layer0_outputs(8070) <= not b or a;
    layer0_outputs(8071) <= 1'b1;
    layer0_outputs(8072) <= b and not a;
    layer0_outputs(8073) <= b;
    layer0_outputs(8074) <= b and not a;
    layer0_outputs(8075) <= not b or a;
    layer0_outputs(8076) <= not b;
    layer0_outputs(8077) <= a xor b;
    layer0_outputs(8078) <= a xor b;
    layer0_outputs(8079) <= 1'b0;
    layer0_outputs(8080) <= a and not b;
    layer0_outputs(8081) <= a and b;
    layer0_outputs(8082) <= a or b;
    layer0_outputs(8083) <= not b or a;
    layer0_outputs(8084) <= b;
    layer0_outputs(8085) <= a and b;
    layer0_outputs(8086) <= not a;
    layer0_outputs(8087) <= a;
    layer0_outputs(8088) <= a or b;
    layer0_outputs(8089) <= not b;
    layer0_outputs(8090) <= a or b;
    layer0_outputs(8091) <= not (a xor b);
    layer0_outputs(8092) <= b;
    layer0_outputs(8093) <= not b;
    layer0_outputs(8094) <= a xor b;
    layer0_outputs(8095) <= not (a and b);
    layer0_outputs(8096) <= not (a and b);
    layer0_outputs(8097) <= a or b;
    layer0_outputs(8098) <= a;
    layer0_outputs(8099) <= not (a or b);
    layer0_outputs(8100) <= not (a xor b);
    layer0_outputs(8101) <= not a or b;
    layer0_outputs(8102) <= not b;
    layer0_outputs(8103) <= not (a xor b);
    layer0_outputs(8104) <= not b;
    layer0_outputs(8105) <= 1'b0;
    layer0_outputs(8106) <= b;
    layer0_outputs(8107) <= not b or a;
    layer0_outputs(8108) <= not a;
    layer0_outputs(8109) <= a xor b;
    layer0_outputs(8110) <= not (a or b);
    layer0_outputs(8111) <= 1'b1;
    layer0_outputs(8112) <= b;
    layer0_outputs(8113) <= not (a and b);
    layer0_outputs(8114) <= not a;
    layer0_outputs(8115) <= not b;
    layer0_outputs(8116) <= a;
    layer0_outputs(8117) <= 1'b0;
    layer0_outputs(8118) <= 1'b0;
    layer0_outputs(8119) <= a or b;
    layer0_outputs(8120) <= not a;
    layer0_outputs(8121) <= not (a or b);
    layer0_outputs(8122) <= not (a and b);
    layer0_outputs(8123) <= a and not b;
    layer0_outputs(8124) <= not a;
    layer0_outputs(8125) <= not a;
    layer0_outputs(8126) <= not (a and b);
    layer0_outputs(8127) <= a or b;
    layer0_outputs(8128) <= a and not b;
    layer0_outputs(8129) <= a or b;
    layer0_outputs(8130) <= not b;
    layer0_outputs(8131) <= a and b;
    layer0_outputs(8132) <= b and not a;
    layer0_outputs(8133) <= a;
    layer0_outputs(8134) <= not (a and b);
    layer0_outputs(8135) <= b;
    layer0_outputs(8136) <= not (a or b);
    layer0_outputs(8137) <= not b;
    layer0_outputs(8138) <= not (a xor b);
    layer0_outputs(8139) <= a xor b;
    layer0_outputs(8140) <= not a;
    layer0_outputs(8141) <= not a or b;
    layer0_outputs(8142) <= not (a xor b);
    layer0_outputs(8143) <= a xor b;
    layer0_outputs(8144) <= b and not a;
    layer0_outputs(8145) <= a or b;
    layer0_outputs(8146) <= not (a and b);
    layer0_outputs(8147) <= b and not a;
    layer0_outputs(8148) <= not a;
    layer0_outputs(8149) <= not (a xor b);
    layer0_outputs(8150) <= b and not a;
    layer0_outputs(8151) <= a;
    layer0_outputs(8152) <= a xor b;
    layer0_outputs(8153) <= a xor b;
    layer0_outputs(8154) <= 1'b0;
    layer0_outputs(8155) <= not (a and b);
    layer0_outputs(8156) <= 1'b0;
    layer0_outputs(8157) <= a xor b;
    layer0_outputs(8158) <= b and not a;
    layer0_outputs(8159) <= a xor b;
    layer0_outputs(8160) <= not (a or b);
    layer0_outputs(8161) <= b;
    layer0_outputs(8162) <= not (a or b);
    layer0_outputs(8163) <= not a;
    layer0_outputs(8164) <= not (a xor b);
    layer0_outputs(8165) <= a xor b;
    layer0_outputs(8166) <= not (a or b);
    layer0_outputs(8167) <= 1'b0;
    layer0_outputs(8168) <= not a or b;
    layer0_outputs(8169) <= b;
    layer0_outputs(8170) <= not (a or b);
    layer0_outputs(8171) <= not a or b;
    layer0_outputs(8172) <= not (a and b);
    layer0_outputs(8173) <= not b or a;
    layer0_outputs(8174) <= not a;
    layer0_outputs(8175) <= not b or a;
    layer0_outputs(8176) <= a xor b;
    layer0_outputs(8177) <= not (a xor b);
    layer0_outputs(8178) <= not (a or b);
    layer0_outputs(8179) <= a xor b;
    layer0_outputs(8180) <= a or b;
    layer0_outputs(8181) <= not b;
    layer0_outputs(8182) <= not a or b;
    layer0_outputs(8183) <= not (a or b);
    layer0_outputs(8184) <= not a or b;
    layer0_outputs(8185) <= a or b;
    layer0_outputs(8186) <= not (a xor b);
    layer0_outputs(8187) <= a or b;
    layer0_outputs(8188) <= not b;
    layer0_outputs(8189) <= 1'b0;
    layer0_outputs(8190) <= not (a or b);
    layer0_outputs(8191) <= not a;
    layer0_outputs(8192) <= not a;
    layer0_outputs(8193) <= not b or a;
    layer0_outputs(8194) <= a or b;
    layer0_outputs(8195) <= b and not a;
    layer0_outputs(8196) <= a;
    layer0_outputs(8197) <= not (a and b);
    layer0_outputs(8198) <= a and not b;
    layer0_outputs(8199) <= not a or b;
    layer0_outputs(8200) <= a and b;
    layer0_outputs(8201) <= a or b;
    layer0_outputs(8202) <= not a;
    layer0_outputs(8203) <= a;
    layer0_outputs(8204) <= not a or b;
    layer0_outputs(8205) <= not b or a;
    layer0_outputs(8206) <= a;
    layer0_outputs(8207) <= not a;
    layer0_outputs(8208) <= b and not a;
    layer0_outputs(8209) <= not (a xor b);
    layer0_outputs(8210) <= not (a or b);
    layer0_outputs(8211) <= not (a or b);
    layer0_outputs(8212) <= a or b;
    layer0_outputs(8213) <= a or b;
    layer0_outputs(8214) <= not b or a;
    layer0_outputs(8215) <= 1'b0;
    layer0_outputs(8216) <= a xor b;
    layer0_outputs(8217) <= not b or a;
    layer0_outputs(8218) <= not a;
    layer0_outputs(8219) <= not (a xor b);
    layer0_outputs(8220) <= not (a xor b);
    layer0_outputs(8221) <= not (a or b);
    layer0_outputs(8222) <= not b or a;
    layer0_outputs(8223) <= not (a or b);
    layer0_outputs(8224) <= not b or a;
    layer0_outputs(8225) <= b and not a;
    layer0_outputs(8226) <= b;
    layer0_outputs(8227) <= a xor b;
    layer0_outputs(8228) <= not (a and b);
    layer0_outputs(8229) <= not b or a;
    layer0_outputs(8230) <= not (a or b);
    layer0_outputs(8231) <= not (a and b);
    layer0_outputs(8232) <= b and not a;
    layer0_outputs(8233) <= not b or a;
    layer0_outputs(8234) <= b;
    layer0_outputs(8235) <= a;
    layer0_outputs(8236) <= not a;
    layer0_outputs(8237) <= a;
    layer0_outputs(8238) <= a and b;
    layer0_outputs(8239) <= a and not b;
    layer0_outputs(8240) <= a;
    layer0_outputs(8241) <= 1'b0;
    layer0_outputs(8242) <= not (a or b);
    layer0_outputs(8243) <= not a or b;
    layer0_outputs(8244) <= a and not b;
    layer0_outputs(8245) <= a and b;
    layer0_outputs(8246) <= a;
    layer0_outputs(8247) <= not b;
    layer0_outputs(8248) <= not a;
    layer0_outputs(8249) <= a or b;
    layer0_outputs(8250) <= a or b;
    layer0_outputs(8251) <= not (a and b);
    layer0_outputs(8252) <= 1'b0;
    layer0_outputs(8253) <= a and b;
    layer0_outputs(8254) <= a;
    layer0_outputs(8255) <= not (a and b);
    layer0_outputs(8256) <= 1'b1;
    layer0_outputs(8257) <= not b or a;
    layer0_outputs(8258) <= a;
    layer0_outputs(8259) <= a;
    layer0_outputs(8260) <= not a;
    layer0_outputs(8261) <= a or b;
    layer0_outputs(8262) <= not a or b;
    layer0_outputs(8263) <= not a or b;
    layer0_outputs(8264) <= a xor b;
    layer0_outputs(8265) <= not a;
    layer0_outputs(8266) <= a and b;
    layer0_outputs(8267) <= not a or b;
    layer0_outputs(8268) <= a or b;
    layer0_outputs(8269) <= not a;
    layer0_outputs(8270) <= not a or b;
    layer0_outputs(8271) <= not a;
    layer0_outputs(8272) <= a or b;
    layer0_outputs(8273) <= not b or a;
    layer0_outputs(8274) <= a;
    layer0_outputs(8275) <= not (a and b);
    layer0_outputs(8276) <= not a;
    layer0_outputs(8277) <= not (a xor b);
    layer0_outputs(8278) <= not (a or b);
    layer0_outputs(8279) <= 1'b1;
    layer0_outputs(8280) <= not (a or b);
    layer0_outputs(8281) <= not b;
    layer0_outputs(8282) <= not b;
    layer0_outputs(8283) <= not a or b;
    layer0_outputs(8284) <= not a;
    layer0_outputs(8285) <= not b;
    layer0_outputs(8286) <= a or b;
    layer0_outputs(8287) <= not a;
    layer0_outputs(8288) <= a;
    layer0_outputs(8289) <= not b;
    layer0_outputs(8290) <= a or b;
    layer0_outputs(8291) <= a xor b;
    layer0_outputs(8292) <= a;
    layer0_outputs(8293) <= a;
    layer0_outputs(8294) <= not (a xor b);
    layer0_outputs(8295) <= not a or b;
    layer0_outputs(8296) <= not a;
    layer0_outputs(8297) <= a and not b;
    layer0_outputs(8298) <= b;
    layer0_outputs(8299) <= a and not b;
    layer0_outputs(8300) <= not (a or b);
    layer0_outputs(8301) <= a or b;
    layer0_outputs(8302) <= not (a or b);
    layer0_outputs(8303) <= b;
    layer0_outputs(8304) <= a;
    layer0_outputs(8305) <= b;
    layer0_outputs(8306) <= a or b;
    layer0_outputs(8307) <= not a;
    layer0_outputs(8308) <= a xor b;
    layer0_outputs(8309) <= a and b;
    layer0_outputs(8310) <= not b;
    layer0_outputs(8311) <= not a or b;
    layer0_outputs(8312) <= a or b;
    layer0_outputs(8313) <= a xor b;
    layer0_outputs(8314) <= not (a and b);
    layer0_outputs(8315) <= not b or a;
    layer0_outputs(8316) <= a;
    layer0_outputs(8317) <= a or b;
    layer0_outputs(8318) <= a xor b;
    layer0_outputs(8319) <= b;
    layer0_outputs(8320) <= not a;
    layer0_outputs(8321) <= not b or a;
    layer0_outputs(8322) <= a or b;
    layer0_outputs(8323) <= a and b;
    layer0_outputs(8324) <= a or b;
    layer0_outputs(8325) <= not a or b;
    layer0_outputs(8326) <= not (a or b);
    layer0_outputs(8327) <= a xor b;
    layer0_outputs(8328) <= a and b;
    layer0_outputs(8329) <= 1'b0;
    layer0_outputs(8330) <= a xor b;
    layer0_outputs(8331) <= not (a xor b);
    layer0_outputs(8332) <= not b or a;
    layer0_outputs(8333) <= b and not a;
    layer0_outputs(8334) <= b;
    layer0_outputs(8335) <= a and b;
    layer0_outputs(8336) <= not a or b;
    layer0_outputs(8337) <= not a or b;
    layer0_outputs(8338) <= a and not b;
    layer0_outputs(8339) <= not b or a;
    layer0_outputs(8340) <= b;
    layer0_outputs(8341) <= b;
    layer0_outputs(8342) <= not b or a;
    layer0_outputs(8343) <= a xor b;
    layer0_outputs(8344) <= b and not a;
    layer0_outputs(8345) <= not b or a;
    layer0_outputs(8346) <= a or b;
    layer0_outputs(8347) <= a and b;
    layer0_outputs(8348) <= a and b;
    layer0_outputs(8349) <= not b;
    layer0_outputs(8350) <= not a;
    layer0_outputs(8351) <= a or b;
    layer0_outputs(8352) <= a and b;
    layer0_outputs(8353) <= not a;
    layer0_outputs(8354) <= not (a xor b);
    layer0_outputs(8355) <= a xor b;
    layer0_outputs(8356) <= b;
    layer0_outputs(8357) <= a xor b;
    layer0_outputs(8358) <= not (a or b);
    layer0_outputs(8359) <= b;
    layer0_outputs(8360) <= not a;
    layer0_outputs(8361) <= b and not a;
    layer0_outputs(8362) <= not (a or b);
    layer0_outputs(8363) <= not (a xor b);
    layer0_outputs(8364) <= not a;
    layer0_outputs(8365) <= a or b;
    layer0_outputs(8366) <= a xor b;
    layer0_outputs(8367) <= a xor b;
    layer0_outputs(8368) <= 1'b0;
    layer0_outputs(8369) <= a or b;
    layer0_outputs(8370) <= a and not b;
    layer0_outputs(8371) <= not (a or b);
    layer0_outputs(8372) <= not b;
    layer0_outputs(8373) <= not (a or b);
    layer0_outputs(8374) <= b;
    layer0_outputs(8375) <= b and not a;
    layer0_outputs(8376) <= a xor b;
    layer0_outputs(8377) <= a xor b;
    layer0_outputs(8378) <= not (a xor b);
    layer0_outputs(8379) <= not (a xor b);
    layer0_outputs(8380) <= a;
    layer0_outputs(8381) <= 1'b1;
    layer0_outputs(8382) <= not b or a;
    layer0_outputs(8383) <= b;
    layer0_outputs(8384) <= not a;
    layer0_outputs(8385) <= not (a xor b);
    layer0_outputs(8386) <= not a or b;
    layer0_outputs(8387) <= not b;
    layer0_outputs(8388) <= not (a or b);
    layer0_outputs(8389) <= not (a and b);
    layer0_outputs(8390) <= a or b;
    layer0_outputs(8391) <= not b or a;
    layer0_outputs(8392) <= not a or b;
    layer0_outputs(8393) <= not a or b;
    layer0_outputs(8394) <= a and not b;
    layer0_outputs(8395) <= 1'b1;
    layer0_outputs(8396) <= not (a or b);
    layer0_outputs(8397) <= not a;
    layer0_outputs(8398) <= a xor b;
    layer0_outputs(8399) <= a xor b;
    layer0_outputs(8400) <= a xor b;
    layer0_outputs(8401) <= not (a xor b);
    layer0_outputs(8402) <= not b or a;
    layer0_outputs(8403) <= not a or b;
    layer0_outputs(8404) <= not a or b;
    layer0_outputs(8405) <= a;
    layer0_outputs(8406) <= 1'b0;
    layer0_outputs(8407) <= not a;
    layer0_outputs(8408) <= not (a and b);
    layer0_outputs(8409) <= b;
    layer0_outputs(8410) <= a or b;
    layer0_outputs(8411) <= a or b;
    layer0_outputs(8412) <= a;
    layer0_outputs(8413) <= a;
    layer0_outputs(8414) <= not b;
    layer0_outputs(8415) <= not a;
    layer0_outputs(8416) <= 1'b1;
    layer0_outputs(8417) <= not a or b;
    layer0_outputs(8418) <= b and not a;
    layer0_outputs(8419) <= a or b;
    layer0_outputs(8420) <= a or b;
    layer0_outputs(8421) <= not (a xor b);
    layer0_outputs(8422) <= not a;
    layer0_outputs(8423) <= not (a xor b);
    layer0_outputs(8424) <= not a;
    layer0_outputs(8425) <= a or b;
    layer0_outputs(8426) <= a;
    layer0_outputs(8427) <= a or b;
    layer0_outputs(8428) <= not (a xor b);
    layer0_outputs(8429) <= not a or b;
    layer0_outputs(8430) <= a and not b;
    layer0_outputs(8431) <= not a;
    layer0_outputs(8432) <= b;
    layer0_outputs(8433) <= b and not a;
    layer0_outputs(8434) <= b and not a;
    layer0_outputs(8435) <= not a;
    layer0_outputs(8436) <= not (a or b);
    layer0_outputs(8437) <= b;
    layer0_outputs(8438) <= a;
    layer0_outputs(8439) <= not b or a;
    layer0_outputs(8440) <= not a;
    layer0_outputs(8441) <= not (a xor b);
    layer0_outputs(8442) <= not b or a;
    layer0_outputs(8443) <= not a;
    layer0_outputs(8444) <= b;
    layer0_outputs(8445) <= b and not a;
    layer0_outputs(8446) <= a;
    layer0_outputs(8447) <= a and not b;
    layer0_outputs(8448) <= not b;
    layer0_outputs(8449) <= a and not b;
    layer0_outputs(8450) <= a and b;
    layer0_outputs(8451) <= not a;
    layer0_outputs(8452) <= not a;
    layer0_outputs(8453) <= not b or a;
    layer0_outputs(8454) <= not a;
    layer0_outputs(8455) <= not b;
    layer0_outputs(8456) <= not a;
    layer0_outputs(8457) <= a xor b;
    layer0_outputs(8458) <= not b;
    layer0_outputs(8459) <= 1'b0;
    layer0_outputs(8460) <= a or b;
    layer0_outputs(8461) <= a or b;
    layer0_outputs(8462) <= not (a or b);
    layer0_outputs(8463) <= a xor b;
    layer0_outputs(8464) <= not b;
    layer0_outputs(8465) <= a and b;
    layer0_outputs(8466) <= not (a or b);
    layer0_outputs(8467) <= not b or a;
    layer0_outputs(8468) <= not (a xor b);
    layer0_outputs(8469) <= not (a xor b);
    layer0_outputs(8470) <= not a;
    layer0_outputs(8471) <= not (a or b);
    layer0_outputs(8472) <= 1'b0;
    layer0_outputs(8473) <= a and b;
    layer0_outputs(8474) <= not (a xor b);
    layer0_outputs(8475) <= a;
    layer0_outputs(8476) <= a xor b;
    layer0_outputs(8477) <= not a;
    layer0_outputs(8478) <= not b;
    layer0_outputs(8479) <= b and not a;
    layer0_outputs(8480) <= a and b;
    layer0_outputs(8481) <= a or b;
    layer0_outputs(8482) <= a or b;
    layer0_outputs(8483) <= not b or a;
    layer0_outputs(8484) <= not (a or b);
    layer0_outputs(8485) <= b and not a;
    layer0_outputs(8486) <= not (a or b);
    layer0_outputs(8487) <= not b or a;
    layer0_outputs(8488) <= b and not a;
    layer0_outputs(8489) <= not a or b;
    layer0_outputs(8490) <= not b;
    layer0_outputs(8491) <= b and not a;
    layer0_outputs(8492) <= a and not b;
    layer0_outputs(8493) <= a and b;
    layer0_outputs(8494) <= not (a or b);
    layer0_outputs(8495) <= b and not a;
    layer0_outputs(8496) <= a and not b;
    layer0_outputs(8497) <= a or b;
    layer0_outputs(8498) <= not a or b;
    layer0_outputs(8499) <= 1'b0;
    layer0_outputs(8500) <= not (a or b);
    layer0_outputs(8501) <= not a or b;
    layer0_outputs(8502) <= a;
    layer0_outputs(8503) <= not b or a;
    layer0_outputs(8504) <= b and not a;
    layer0_outputs(8505) <= not (a xor b);
    layer0_outputs(8506) <= b and not a;
    layer0_outputs(8507) <= a;
    layer0_outputs(8508) <= not a or b;
    layer0_outputs(8509) <= a and not b;
    layer0_outputs(8510) <= not b or a;
    layer0_outputs(8511) <= a or b;
    layer0_outputs(8512) <= not a or b;
    layer0_outputs(8513) <= not b or a;
    layer0_outputs(8514) <= not b;
    layer0_outputs(8515) <= a and not b;
    layer0_outputs(8516) <= 1'b1;
    layer0_outputs(8517) <= not (a and b);
    layer0_outputs(8518) <= not (a or b);
    layer0_outputs(8519) <= not b;
    layer0_outputs(8520) <= not (a or b);
    layer0_outputs(8521) <= a;
    layer0_outputs(8522) <= a xor b;
    layer0_outputs(8523) <= a and b;
    layer0_outputs(8524) <= a and not b;
    layer0_outputs(8525) <= a and not b;
    layer0_outputs(8526) <= b;
    layer0_outputs(8527) <= not (a or b);
    layer0_outputs(8528) <= not (a and b);
    layer0_outputs(8529) <= not a;
    layer0_outputs(8530) <= a or b;
    layer0_outputs(8531) <= 1'b0;
    layer0_outputs(8532) <= not a;
    layer0_outputs(8533) <= not b or a;
    layer0_outputs(8534) <= b;
    layer0_outputs(8535) <= not b;
    layer0_outputs(8536) <= a;
    layer0_outputs(8537) <= a;
    layer0_outputs(8538) <= not (a xor b);
    layer0_outputs(8539) <= b and not a;
    layer0_outputs(8540) <= 1'b1;
    layer0_outputs(8541) <= b and not a;
    layer0_outputs(8542) <= a and b;
    layer0_outputs(8543) <= a and not b;
    layer0_outputs(8544) <= not a or b;
    layer0_outputs(8545) <= a and b;
    layer0_outputs(8546) <= a or b;
    layer0_outputs(8547) <= not a or b;
    layer0_outputs(8548) <= not (a or b);
    layer0_outputs(8549) <= not a;
    layer0_outputs(8550) <= 1'b1;
    layer0_outputs(8551) <= not a or b;
    layer0_outputs(8552) <= not b;
    layer0_outputs(8553) <= not (a xor b);
    layer0_outputs(8554) <= a and not b;
    layer0_outputs(8555) <= not (a xor b);
    layer0_outputs(8556) <= not (a or b);
    layer0_outputs(8557) <= not a;
    layer0_outputs(8558) <= not (a and b);
    layer0_outputs(8559) <= 1'b0;
    layer0_outputs(8560) <= b;
    layer0_outputs(8561) <= 1'b1;
    layer0_outputs(8562) <= not (a xor b);
    layer0_outputs(8563) <= not b or a;
    layer0_outputs(8564) <= a xor b;
    layer0_outputs(8565) <= not (a or b);
    layer0_outputs(8566) <= b and not a;
    layer0_outputs(8567) <= a and not b;
    layer0_outputs(8568) <= a xor b;
    layer0_outputs(8569) <= b;
    layer0_outputs(8570) <= 1'b1;
    layer0_outputs(8571) <= a or b;
    layer0_outputs(8572) <= not b;
    layer0_outputs(8573) <= a xor b;
    layer0_outputs(8574) <= not b;
    layer0_outputs(8575) <= not (a or b);
    layer0_outputs(8576) <= not (a and b);
    layer0_outputs(8577) <= not a;
    layer0_outputs(8578) <= a and not b;
    layer0_outputs(8579) <= not b;
    layer0_outputs(8580) <= not (a or b);
    layer0_outputs(8581) <= not (a or b);
    layer0_outputs(8582) <= not a;
    layer0_outputs(8583) <= not a;
    layer0_outputs(8584) <= b and not a;
    layer0_outputs(8585) <= not a or b;
    layer0_outputs(8586) <= b;
    layer0_outputs(8587) <= b;
    layer0_outputs(8588) <= a xor b;
    layer0_outputs(8589) <= not a or b;
    layer0_outputs(8590) <= b;
    layer0_outputs(8591) <= not (a or b);
    layer0_outputs(8592) <= not (a or b);
    layer0_outputs(8593) <= not a;
    layer0_outputs(8594) <= not (a or b);
    layer0_outputs(8595) <= b and not a;
    layer0_outputs(8596) <= not a;
    layer0_outputs(8597) <= 1'b1;
    layer0_outputs(8598) <= not (a and b);
    layer0_outputs(8599) <= a and b;
    layer0_outputs(8600) <= not (a and b);
    layer0_outputs(8601) <= not b or a;
    layer0_outputs(8602) <= not a or b;
    layer0_outputs(8603) <= 1'b0;
    layer0_outputs(8604) <= b and not a;
    layer0_outputs(8605) <= a xor b;
    layer0_outputs(8606) <= not a;
    layer0_outputs(8607) <= a xor b;
    layer0_outputs(8608) <= not a;
    layer0_outputs(8609) <= b and not a;
    layer0_outputs(8610) <= a and not b;
    layer0_outputs(8611) <= not (a and b);
    layer0_outputs(8612) <= a xor b;
    layer0_outputs(8613) <= b;
    layer0_outputs(8614) <= a or b;
    layer0_outputs(8615) <= b;
    layer0_outputs(8616) <= a or b;
    layer0_outputs(8617) <= a xor b;
    layer0_outputs(8618) <= a xor b;
    layer0_outputs(8619) <= a or b;
    layer0_outputs(8620) <= a and not b;
    layer0_outputs(8621) <= a or b;
    layer0_outputs(8622) <= 1'b0;
    layer0_outputs(8623) <= not b;
    layer0_outputs(8624) <= not b;
    layer0_outputs(8625) <= not (a xor b);
    layer0_outputs(8626) <= not (a xor b);
    layer0_outputs(8627) <= not (a and b);
    layer0_outputs(8628) <= a and not b;
    layer0_outputs(8629) <= b and not a;
    layer0_outputs(8630) <= not (a xor b);
    layer0_outputs(8631) <= not b or a;
    layer0_outputs(8632) <= a and not b;
    layer0_outputs(8633) <= a or b;
    layer0_outputs(8634) <= a;
    layer0_outputs(8635) <= not (a xor b);
    layer0_outputs(8636) <= b and not a;
    layer0_outputs(8637) <= not (a xor b);
    layer0_outputs(8638) <= not b;
    layer0_outputs(8639) <= not a;
    layer0_outputs(8640) <= a;
    layer0_outputs(8641) <= a xor b;
    layer0_outputs(8642) <= b;
    layer0_outputs(8643) <= not (a and b);
    layer0_outputs(8644) <= b;
    layer0_outputs(8645) <= not b or a;
    layer0_outputs(8646) <= not a;
    layer0_outputs(8647) <= b and not a;
    layer0_outputs(8648) <= a;
    layer0_outputs(8649) <= a and b;
    layer0_outputs(8650) <= b;
    layer0_outputs(8651) <= a xor b;
    layer0_outputs(8652) <= b;
    layer0_outputs(8653) <= a or b;
    layer0_outputs(8654) <= not b;
    layer0_outputs(8655) <= a;
    layer0_outputs(8656) <= a or b;
    layer0_outputs(8657) <= 1'b1;
    layer0_outputs(8658) <= b and not a;
    layer0_outputs(8659) <= not a or b;
    layer0_outputs(8660) <= not a;
    layer0_outputs(8661) <= not a;
    layer0_outputs(8662) <= not (a or b);
    layer0_outputs(8663) <= not (a or b);
    layer0_outputs(8664) <= a and not b;
    layer0_outputs(8665) <= b and not a;
    layer0_outputs(8666) <= a;
    layer0_outputs(8667) <= a xor b;
    layer0_outputs(8668) <= not (a and b);
    layer0_outputs(8669) <= not (a or b);
    layer0_outputs(8670) <= a or b;
    layer0_outputs(8671) <= not (a or b);
    layer0_outputs(8672) <= not a;
    layer0_outputs(8673) <= not a;
    layer0_outputs(8674) <= a or b;
    layer0_outputs(8675) <= not (a or b);
    layer0_outputs(8676) <= b;
    layer0_outputs(8677) <= a or b;
    layer0_outputs(8678) <= 1'b1;
    layer0_outputs(8679) <= b and not a;
    layer0_outputs(8680) <= 1'b0;
    layer0_outputs(8681) <= not b;
    layer0_outputs(8682) <= not a;
    layer0_outputs(8683) <= 1'b1;
    layer0_outputs(8684) <= not (a xor b);
    layer0_outputs(8685) <= a;
    layer0_outputs(8686) <= a or b;
    layer0_outputs(8687) <= not (a xor b);
    layer0_outputs(8688) <= a xor b;
    layer0_outputs(8689) <= not (a or b);
    layer0_outputs(8690) <= 1'b1;
    layer0_outputs(8691) <= not (a or b);
    layer0_outputs(8692) <= b and not a;
    layer0_outputs(8693) <= 1'b0;
    layer0_outputs(8694) <= not (a or b);
    layer0_outputs(8695) <= a and b;
    layer0_outputs(8696) <= a or b;
    layer0_outputs(8697) <= a xor b;
    layer0_outputs(8698) <= b and not a;
    layer0_outputs(8699) <= not (a and b);
    layer0_outputs(8700) <= not a;
    layer0_outputs(8701) <= a or b;
    layer0_outputs(8702) <= not b or a;
    layer0_outputs(8703) <= not a;
    layer0_outputs(8704) <= not b or a;
    layer0_outputs(8705) <= a xor b;
    layer0_outputs(8706) <= b;
    layer0_outputs(8707) <= not b;
    layer0_outputs(8708) <= not a or b;
    layer0_outputs(8709) <= not b;
    layer0_outputs(8710) <= a and not b;
    layer0_outputs(8711) <= not (a or b);
    layer0_outputs(8712) <= not (a or b);
    layer0_outputs(8713) <= a or b;
    layer0_outputs(8714) <= not (a xor b);
    layer0_outputs(8715) <= not (a or b);
    layer0_outputs(8716) <= not a;
    layer0_outputs(8717) <= a;
    layer0_outputs(8718) <= a xor b;
    layer0_outputs(8719) <= not a or b;
    layer0_outputs(8720) <= a or b;
    layer0_outputs(8721) <= a;
    layer0_outputs(8722) <= b;
    layer0_outputs(8723) <= not b;
    layer0_outputs(8724) <= 1'b1;
    layer0_outputs(8725) <= a;
    layer0_outputs(8726) <= not (a or b);
    layer0_outputs(8727) <= a xor b;
    layer0_outputs(8728) <= a xor b;
    layer0_outputs(8729) <= not (a xor b);
    layer0_outputs(8730) <= a and not b;
    layer0_outputs(8731) <= a or b;
    layer0_outputs(8732) <= not a or b;
    layer0_outputs(8733) <= not b or a;
    layer0_outputs(8734) <= a and not b;
    layer0_outputs(8735) <= b;
    layer0_outputs(8736) <= not a or b;
    layer0_outputs(8737) <= not b or a;
    layer0_outputs(8738) <= not a;
    layer0_outputs(8739) <= not (a xor b);
    layer0_outputs(8740) <= not a;
    layer0_outputs(8741) <= a xor b;
    layer0_outputs(8742) <= b and not a;
    layer0_outputs(8743) <= not a;
    layer0_outputs(8744) <= 1'b1;
    layer0_outputs(8745) <= b and not a;
    layer0_outputs(8746) <= a and not b;
    layer0_outputs(8747) <= a and not b;
    layer0_outputs(8748) <= not a;
    layer0_outputs(8749) <= b;
    layer0_outputs(8750) <= 1'b0;
    layer0_outputs(8751) <= not a or b;
    layer0_outputs(8752) <= a or b;
    layer0_outputs(8753) <= a;
    layer0_outputs(8754) <= a or b;
    layer0_outputs(8755) <= not (a xor b);
    layer0_outputs(8756) <= not (a xor b);
    layer0_outputs(8757) <= not a or b;
    layer0_outputs(8758) <= a or b;
    layer0_outputs(8759) <= not (a xor b);
    layer0_outputs(8760) <= 1'b1;
    layer0_outputs(8761) <= a xor b;
    layer0_outputs(8762) <= b and not a;
    layer0_outputs(8763) <= b and not a;
    layer0_outputs(8764) <= a or b;
    layer0_outputs(8765) <= not (a or b);
    layer0_outputs(8766) <= b and not a;
    layer0_outputs(8767) <= 1'b0;
    layer0_outputs(8768) <= not b;
    layer0_outputs(8769) <= not a or b;
    layer0_outputs(8770) <= not a;
    layer0_outputs(8771) <= not a or b;
    layer0_outputs(8772) <= not (a or b);
    layer0_outputs(8773) <= 1'b1;
    layer0_outputs(8774) <= a and b;
    layer0_outputs(8775) <= a and b;
    layer0_outputs(8776) <= not a;
    layer0_outputs(8777) <= not b or a;
    layer0_outputs(8778) <= not b;
    layer0_outputs(8779) <= a and b;
    layer0_outputs(8780) <= 1'b1;
    layer0_outputs(8781) <= a;
    layer0_outputs(8782) <= 1'b1;
    layer0_outputs(8783) <= b and not a;
    layer0_outputs(8784) <= not a;
    layer0_outputs(8785) <= 1'b0;
    layer0_outputs(8786) <= a;
    layer0_outputs(8787) <= a xor b;
    layer0_outputs(8788) <= a or b;
    layer0_outputs(8789) <= 1'b0;
    layer0_outputs(8790) <= not a or b;
    layer0_outputs(8791) <= b;
    layer0_outputs(8792) <= not a;
    layer0_outputs(8793) <= not a or b;
    layer0_outputs(8794) <= a and not b;
    layer0_outputs(8795) <= 1'b0;
    layer0_outputs(8796) <= b;
    layer0_outputs(8797) <= not b or a;
    layer0_outputs(8798) <= a and b;
    layer0_outputs(8799) <= 1'b1;
    layer0_outputs(8800) <= 1'b1;
    layer0_outputs(8801) <= not (a xor b);
    layer0_outputs(8802) <= a and not b;
    layer0_outputs(8803) <= a xor b;
    layer0_outputs(8804) <= a;
    layer0_outputs(8805) <= a or b;
    layer0_outputs(8806) <= a xor b;
    layer0_outputs(8807) <= a;
    layer0_outputs(8808) <= not (a xor b);
    layer0_outputs(8809) <= not a or b;
    layer0_outputs(8810) <= not (a or b);
    layer0_outputs(8811) <= a and b;
    layer0_outputs(8812) <= b and not a;
    layer0_outputs(8813) <= a xor b;
    layer0_outputs(8814) <= not a or b;
    layer0_outputs(8815) <= not (a and b);
    layer0_outputs(8816) <= 1'b1;
    layer0_outputs(8817) <= not a;
    layer0_outputs(8818) <= b and not a;
    layer0_outputs(8819) <= not (a and b);
    layer0_outputs(8820) <= not (a and b);
    layer0_outputs(8821) <= not b or a;
    layer0_outputs(8822) <= 1'b1;
    layer0_outputs(8823) <= not (a or b);
    layer0_outputs(8824) <= a and not b;
    layer0_outputs(8825) <= not (a xor b);
    layer0_outputs(8826) <= b;
    layer0_outputs(8827) <= a and not b;
    layer0_outputs(8828) <= a or b;
    layer0_outputs(8829) <= b and not a;
    layer0_outputs(8830) <= not a;
    layer0_outputs(8831) <= not b or a;
    layer0_outputs(8832) <= not (a xor b);
    layer0_outputs(8833) <= b and not a;
    layer0_outputs(8834) <= b and not a;
    layer0_outputs(8835) <= a or b;
    layer0_outputs(8836) <= not a or b;
    layer0_outputs(8837) <= not (a or b);
    layer0_outputs(8838) <= not (a and b);
    layer0_outputs(8839) <= a or b;
    layer0_outputs(8840) <= a;
    layer0_outputs(8841) <= 1'b0;
    layer0_outputs(8842) <= b;
    layer0_outputs(8843) <= a or b;
    layer0_outputs(8844) <= b and not a;
    layer0_outputs(8845) <= b and not a;
    layer0_outputs(8846) <= a;
    layer0_outputs(8847) <= not b;
    layer0_outputs(8848) <= b and not a;
    layer0_outputs(8849) <= a or b;
    layer0_outputs(8850) <= not a or b;
    layer0_outputs(8851) <= 1'b1;
    layer0_outputs(8852) <= a and not b;
    layer0_outputs(8853) <= b;
    layer0_outputs(8854) <= not (a and b);
    layer0_outputs(8855) <= not a;
    layer0_outputs(8856) <= not b or a;
    layer0_outputs(8857) <= a and not b;
    layer0_outputs(8858) <= not (a or b);
    layer0_outputs(8859) <= not (a or b);
    layer0_outputs(8860) <= a and not b;
    layer0_outputs(8861) <= not b or a;
    layer0_outputs(8862) <= a and not b;
    layer0_outputs(8863) <= a;
    layer0_outputs(8864) <= not (a or b);
    layer0_outputs(8865) <= not a or b;
    layer0_outputs(8866) <= a;
    layer0_outputs(8867) <= b and not a;
    layer0_outputs(8868) <= a;
    layer0_outputs(8869) <= 1'b1;
    layer0_outputs(8870) <= not b or a;
    layer0_outputs(8871) <= not a;
    layer0_outputs(8872) <= not a;
    layer0_outputs(8873) <= not (a or b);
    layer0_outputs(8874) <= 1'b1;
    layer0_outputs(8875) <= b;
    layer0_outputs(8876) <= not b or a;
    layer0_outputs(8877) <= not (a or b);
    layer0_outputs(8878) <= not (a and b);
    layer0_outputs(8879) <= not (a xor b);
    layer0_outputs(8880) <= not a;
    layer0_outputs(8881) <= not b;
    layer0_outputs(8882) <= not a;
    layer0_outputs(8883) <= a or b;
    layer0_outputs(8884) <= a or b;
    layer0_outputs(8885) <= not a or b;
    layer0_outputs(8886) <= not a or b;
    layer0_outputs(8887) <= a and not b;
    layer0_outputs(8888) <= a xor b;
    layer0_outputs(8889) <= not a or b;
    layer0_outputs(8890) <= a or b;
    layer0_outputs(8891) <= 1'b1;
    layer0_outputs(8892) <= not b;
    layer0_outputs(8893) <= a;
    layer0_outputs(8894) <= 1'b0;
    layer0_outputs(8895) <= a or b;
    layer0_outputs(8896) <= not (a or b);
    layer0_outputs(8897) <= not b;
    layer0_outputs(8898) <= a;
    layer0_outputs(8899) <= not (a or b);
    layer0_outputs(8900) <= b and not a;
    layer0_outputs(8901) <= a;
    layer0_outputs(8902) <= not a or b;
    layer0_outputs(8903) <= not (a and b);
    layer0_outputs(8904) <= a or b;
    layer0_outputs(8905) <= a and not b;
    layer0_outputs(8906) <= not b;
    layer0_outputs(8907) <= 1'b0;
    layer0_outputs(8908) <= not (a or b);
    layer0_outputs(8909) <= b and not a;
    layer0_outputs(8910) <= a or b;
    layer0_outputs(8911) <= not b;
    layer0_outputs(8912) <= not a;
    layer0_outputs(8913) <= 1'b0;
    layer0_outputs(8914) <= 1'b0;
    layer0_outputs(8915) <= not (a or b);
    layer0_outputs(8916) <= b and not a;
    layer0_outputs(8917) <= not b;
    layer0_outputs(8918) <= a xor b;
    layer0_outputs(8919) <= a xor b;
    layer0_outputs(8920) <= not b or a;
    layer0_outputs(8921) <= a or b;
    layer0_outputs(8922) <= b and not a;
    layer0_outputs(8923) <= a;
    layer0_outputs(8924) <= not b or a;
    layer0_outputs(8925) <= b;
    layer0_outputs(8926) <= b;
    layer0_outputs(8927) <= not (a or b);
    layer0_outputs(8928) <= 1'b0;
    layer0_outputs(8929) <= b and not a;
    layer0_outputs(8930) <= a;
    layer0_outputs(8931) <= not b;
    layer0_outputs(8932) <= not (a or b);
    layer0_outputs(8933) <= not (a or b);
    layer0_outputs(8934) <= not a or b;
    layer0_outputs(8935) <= 1'b0;
    layer0_outputs(8936) <= not b;
    layer0_outputs(8937) <= a or b;
    layer0_outputs(8938) <= not a;
    layer0_outputs(8939) <= a;
    layer0_outputs(8940) <= b;
    layer0_outputs(8941) <= 1'b0;
    layer0_outputs(8942) <= not (a or b);
    layer0_outputs(8943) <= 1'b1;
    layer0_outputs(8944) <= a or b;
    layer0_outputs(8945) <= not b or a;
    layer0_outputs(8946) <= not a or b;
    layer0_outputs(8947) <= not a;
    layer0_outputs(8948) <= not a or b;
    layer0_outputs(8949) <= 1'b1;
    layer0_outputs(8950) <= a xor b;
    layer0_outputs(8951) <= 1'b0;
    layer0_outputs(8952) <= a xor b;
    layer0_outputs(8953) <= not (a and b);
    layer0_outputs(8954) <= not (a or b);
    layer0_outputs(8955) <= a or b;
    layer0_outputs(8956) <= not a or b;
    layer0_outputs(8957) <= not b or a;
    layer0_outputs(8958) <= not a;
    layer0_outputs(8959) <= not a;
    layer0_outputs(8960) <= b;
    layer0_outputs(8961) <= b and not a;
    layer0_outputs(8962) <= not (a or b);
    layer0_outputs(8963) <= not b or a;
    layer0_outputs(8964) <= a or b;
    layer0_outputs(8965) <= a;
    layer0_outputs(8966) <= 1'b0;
    layer0_outputs(8967) <= a or b;
    layer0_outputs(8968) <= not (a xor b);
    layer0_outputs(8969) <= a and not b;
    layer0_outputs(8970) <= a xor b;
    layer0_outputs(8971) <= a or b;
    layer0_outputs(8972) <= a xor b;
    layer0_outputs(8973) <= 1'b1;
    layer0_outputs(8974) <= not a;
    layer0_outputs(8975) <= a xor b;
    layer0_outputs(8976) <= a or b;
    layer0_outputs(8977) <= a or b;
    layer0_outputs(8978) <= not (a or b);
    layer0_outputs(8979) <= not b or a;
    layer0_outputs(8980) <= a and not b;
    layer0_outputs(8981) <= not b;
    layer0_outputs(8982) <= not a or b;
    layer0_outputs(8983) <= 1'b0;
    layer0_outputs(8984) <= b and not a;
    layer0_outputs(8985) <= not (a xor b);
    layer0_outputs(8986) <= b;
    layer0_outputs(8987) <= not (a or b);
    layer0_outputs(8988) <= not (a or b);
    layer0_outputs(8989) <= not (a xor b);
    layer0_outputs(8990) <= a and not b;
    layer0_outputs(8991) <= not (a and b);
    layer0_outputs(8992) <= not a;
    layer0_outputs(8993) <= not b or a;
    layer0_outputs(8994) <= a and not b;
    layer0_outputs(8995) <= not a;
    layer0_outputs(8996) <= not (a xor b);
    layer0_outputs(8997) <= 1'b0;
    layer0_outputs(8998) <= a xor b;
    layer0_outputs(8999) <= not b;
    layer0_outputs(9000) <= b;
    layer0_outputs(9001) <= not b;
    layer0_outputs(9002) <= not a;
    layer0_outputs(9003) <= a or b;
    layer0_outputs(9004) <= not (a or b);
    layer0_outputs(9005) <= b;
    layer0_outputs(9006) <= not b;
    layer0_outputs(9007) <= b;
    layer0_outputs(9008) <= not (a or b);
    layer0_outputs(9009) <= not a;
    layer0_outputs(9010) <= b and not a;
    layer0_outputs(9011) <= not (a xor b);
    layer0_outputs(9012) <= not b or a;
    layer0_outputs(9013) <= not a or b;
    layer0_outputs(9014) <= a and b;
    layer0_outputs(9015) <= not (a or b);
    layer0_outputs(9016) <= a and not b;
    layer0_outputs(9017) <= a and b;
    layer0_outputs(9018) <= not (a or b);
    layer0_outputs(9019) <= not b or a;
    layer0_outputs(9020) <= a and not b;
    layer0_outputs(9021) <= b;
    layer0_outputs(9022) <= b and not a;
    layer0_outputs(9023) <= 1'b0;
    layer0_outputs(9024) <= not (a xor b);
    layer0_outputs(9025) <= a;
    layer0_outputs(9026) <= b and not a;
    layer0_outputs(9027) <= a and not b;
    layer0_outputs(9028) <= not b;
    layer0_outputs(9029) <= b and not a;
    layer0_outputs(9030) <= not b or a;
    layer0_outputs(9031) <= b;
    layer0_outputs(9032) <= a;
    layer0_outputs(9033) <= a and b;
    layer0_outputs(9034) <= a or b;
    layer0_outputs(9035) <= a;
    layer0_outputs(9036) <= not b;
    layer0_outputs(9037) <= not a or b;
    layer0_outputs(9038) <= a xor b;
    layer0_outputs(9039) <= not (a or b);
    layer0_outputs(9040) <= not b;
    layer0_outputs(9041) <= not a;
    layer0_outputs(9042) <= a and not b;
    layer0_outputs(9043) <= a xor b;
    layer0_outputs(9044) <= not (a xor b);
    layer0_outputs(9045) <= b;
    layer0_outputs(9046) <= not (a or b);
    layer0_outputs(9047) <= a and not b;
    layer0_outputs(9048) <= a xor b;
    layer0_outputs(9049) <= a and not b;
    layer0_outputs(9050) <= 1'b0;
    layer0_outputs(9051) <= a xor b;
    layer0_outputs(9052) <= not (a or b);
    layer0_outputs(9053) <= not b;
    layer0_outputs(9054) <= a;
    layer0_outputs(9055) <= not (a or b);
    layer0_outputs(9056) <= a or b;
    layer0_outputs(9057) <= a;
    layer0_outputs(9058) <= not (a xor b);
    layer0_outputs(9059) <= a and not b;
    layer0_outputs(9060) <= 1'b1;
    layer0_outputs(9061) <= not (a and b);
    layer0_outputs(9062) <= not (a or b);
    layer0_outputs(9063) <= not (a or b);
    layer0_outputs(9064) <= b;
    layer0_outputs(9065) <= a;
    layer0_outputs(9066) <= 1'b1;
    layer0_outputs(9067) <= a xor b;
    layer0_outputs(9068) <= not b or a;
    layer0_outputs(9069) <= a;
    layer0_outputs(9070) <= a;
    layer0_outputs(9071) <= a or b;
    layer0_outputs(9072) <= 1'b1;
    layer0_outputs(9073) <= b and not a;
    layer0_outputs(9074) <= not (a or b);
    layer0_outputs(9075) <= not (a or b);
    layer0_outputs(9076) <= not (a or b);
    layer0_outputs(9077) <= a or b;
    layer0_outputs(9078) <= a and not b;
    layer0_outputs(9079) <= a and b;
    layer0_outputs(9080) <= 1'b1;
    layer0_outputs(9081) <= not a;
    layer0_outputs(9082) <= not b;
    layer0_outputs(9083) <= a;
    layer0_outputs(9084) <= 1'b0;
    layer0_outputs(9085) <= not a or b;
    layer0_outputs(9086) <= not b or a;
    layer0_outputs(9087) <= not (a and b);
    layer0_outputs(9088) <= not b;
    layer0_outputs(9089) <= not b or a;
    layer0_outputs(9090) <= not a;
    layer0_outputs(9091) <= b;
    layer0_outputs(9092) <= b;
    layer0_outputs(9093) <= not a;
    layer0_outputs(9094) <= a;
    layer0_outputs(9095) <= a;
    layer0_outputs(9096) <= b and not a;
    layer0_outputs(9097) <= not (a and b);
    layer0_outputs(9098) <= a and not b;
    layer0_outputs(9099) <= not (a or b);
    layer0_outputs(9100) <= b and not a;
    layer0_outputs(9101) <= not b;
    layer0_outputs(9102) <= a or b;
    layer0_outputs(9103) <= not a;
    layer0_outputs(9104) <= a or b;
    layer0_outputs(9105) <= not (a or b);
    layer0_outputs(9106) <= not (a or b);
    layer0_outputs(9107) <= b;
    layer0_outputs(9108) <= b and not a;
    layer0_outputs(9109) <= not b or a;
    layer0_outputs(9110) <= b;
    layer0_outputs(9111) <= b and not a;
    layer0_outputs(9112) <= a or b;
    layer0_outputs(9113) <= not (a and b);
    layer0_outputs(9114) <= not (a and b);
    layer0_outputs(9115) <= a xor b;
    layer0_outputs(9116) <= b;
    layer0_outputs(9117) <= a and not b;
    layer0_outputs(9118) <= a xor b;
    layer0_outputs(9119) <= a xor b;
    layer0_outputs(9120) <= not b or a;
    layer0_outputs(9121) <= a or b;
    layer0_outputs(9122) <= not b or a;
    layer0_outputs(9123) <= not (a xor b);
    layer0_outputs(9124) <= not (a or b);
    layer0_outputs(9125) <= a or b;
    layer0_outputs(9126) <= not b or a;
    layer0_outputs(9127) <= not a;
    layer0_outputs(9128) <= b and not a;
    layer0_outputs(9129) <= not a;
    layer0_outputs(9130) <= not (a xor b);
    layer0_outputs(9131) <= not (a or b);
    layer0_outputs(9132) <= not a;
    layer0_outputs(9133) <= a or b;
    layer0_outputs(9134) <= a;
    layer0_outputs(9135) <= a and b;
    layer0_outputs(9136) <= not (a or b);
    layer0_outputs(9137) <= a or b;
    layer0_outputs(9138) <= b;
    layer0_outputs(9139) <= not a;
    layer0_outputs(9140) <= not (a xor b);
    layer0_outputs(9141) <= b;
    layer0_outputs(9142) <= a or b;
    layer0_outputs(9143) <= a xor b;
    layer0_outputs(9144) <= b;
    layer0_outputs(9145) <= a and b;
    layer0_outputs(9146) <= not (a xor b);
    layer0_outputs(9147) <= not (a or b);
    layer0_outputs(9148) <= not a;
    layer0_outputs(9149) <= 1'b1;
    layer0_outputs(9150) <= not b;
    layer0_outputs(9151) <= not a;
    layer0_outputs(9152) <= b;
    layer0_outputs(9153) <= b and not a;
    layer0_outputs(9154) <= a xor b;
    layer0_outputs(9155) <= a xor b;
    layer0_outputs(9156) <= a and b;
    layer0_outputs(9157) <= not (a xor b);
    layer0_outputs(9158) <= a and b;
    layer0_outputs(9159) <= b and not a;
    layer0_outputs(9160) <= a xor b;
    layer0_outputs(9161) <= not (a or b);
    layer0_outputs(9162) <= not a;
    layer0_outputs(9163) <= a and b;
    layer0_outputs(9164) <= a;
    layer0_outputs(9165) <= a and b;
    layer0_outputs(9166) <= not b;
    layer0_outputs(9167) <= not b;
    layer0_outputs(9168) <= a and not b;
    layer0_outputs(9169) <= b and not a;
    layer0_outputs(9170) <= not a;
    layer0_outputs(9171) <= not (a or b);
    layer0_outputs(9172) <= a xor b;
    layer0_outputs(9173) <= b and not a;
    layer0_outputs(9174) <= a or b;
    layer0_outputs(9175) <= not (a xor b);
    layer0_outputs(9176) <= 1'b1;
    layer0_outputs(9177) <= a or b;
    layer0_outputs(9178) <= 1'b0;
    layer0_outputs(9179) <= a or b;
    layer0_outputs(9180) <= a or b;
    layer0_outputs(9181) <= 1'b1;
    layer0_outputs(9182) <= not b or a;
    layer0_outputs(9183) <= not (a or b);
    layer0_outputs(9184) <= a or b;
    layer0_outputs(9185) <= 1'b0;
    layer0_outputs(9186) <= b and not a;
    layer0_outputs(9187) <= a or b;
    layer0_outputs(9188) <= not (a or b);
    layer0_outputs(9189) <= not (a and b);
    layer0_outputs(9190) <= a;
    layer0_outputs(9191) <= not a or b;
    layer0_outputs(9192) <= a and not b;
    layer0_outputs(9193) <= not b or a;
    layer0_outputs(9194) <= not b;
    layer0_outputs(9195) <= not (a or b);
    layer0_outputs(9196) <= 1'b1;
    layer0_outputs(9197) <= a;
    layer0_outputs(9198) <= not a or b;
    layer0_outputs(9199) <= not (a xor b);
    layer0_outputs(9200) <= a and b;
    layer0_outputs(9201) <= b and not a;
    layer0_outputs(9202) <= not (a or b);
    layer0_outputs(9203) <= b and not a;
    layer0_outputs(9204) <= b;
    layer0_outputs(9205) <= a or b;
    layer0_outputs(9206) <= b and not a;
    layer0_outputs(9207) <= a or b;
    layer0_outputs(9208) <= not (a or b);
    layer0_outputs(9209) <= b;
    layer0_outputs(9210) <= not b;
    layer0_outputs(9211) <= not a;
    layer0_outputs(9212) <= not a or b;
    layer0_outputs(9213) <= not a;
    layer0_outputs(9214) <= not (a or b);
    layer0_outputs(9215) <= not a;
    layer0_outputs(9216) <= not (a xor b);
    layer0_outputs(9217) <= a;
    layer0_outputs(9218) <= not a or b;
    layer0_outputs(9219) <= b;
    layer0_outputs(9220) <= a or b;
    layer0_outputs(9221) <= 1'b0;
    layer0_outputs(9222) <= a;
    layer0_outputs(9223) <= not b;
    layer0_outputs(9224) <= b;
    layer0_outputs(9225) <= 1'b0;
    layer0_outputs(9226) <= not b;
    layer0_outputs(9227) <= not (a and b);
    layer0_outputs(9228) <= a and not b;
    layer0_outputs(9229) <= not (a or b);
    layer0_outputs(9230) <= not a;
    layer0_outputs(9231) <= b;
    layer0_outputs(9232) <= b;
    layer0_outputs(9233) <= b;
    layer0_outputs(9234) <= not a;
    layer0_outputs(9235) <= not a or b;
    layer0_outputs(9236) <= b and not a;
    layer0_outputs(9237) <= not (a xor b);
    layer0_outputs(9238) <= a;
    layer0_outputs(9239) <= a;
    layer0_outputs(9240) <= not a;
    layer0_outputs(9241) <= a xor b;
    layer0_outputs(9242) <= 1'b1;
    layer0_outputs(9243) <= not (a or b);
    layer0_outputs(9244) <= not a;
    layer0_outputs(9245) <= not a or b;
    layer0_outputs(9246) <= not (a or b);
    layer0_outputs(9247) <= not a or b;
    layer0_outputs(9248) <= not b or a;
    layer0_outputs(9249) <= not (a or b);
    layer0_outputs(9250) <= not (a xor b);
    layer0_outputs(9251) <= a and not b;
    layer0_outputs(9252) <= a and b;
    layer0_outputs(9253) <= not (a or b);
    layer0_outputs(9254) <= a xor b;
    layer0_outputs(9255) <= not a;
    layer0_outputs(9256) <= not b or a;
    layer0_outputs(9257) <= b;
    layer0_outputs(9258) <= not a or b;
    layer0_outputs(9259) <= not a;
    layer0_outputs(9260) <= not (a xor b);
    layer0_outputs(9261) <= a and not b;
    layer0_outputs(9262) <= not (a or b);
    layer0_outputs(9263) <= not b;
    layer0_outputs(9264) <= 1'b0;
    layer0_outputs(9265) <= b;
    layer0_outputs(9266) <= not (a xor b);
    layer0_outputs(9267) <= not b;
    layer0_outputs(9268) <= not (a or b);
    layer0_outputs(9269) <= a;
    layer0_outputs(9270) <= a xor b;
    layer0_outputs(9271) <= b and not a;
    layer0_outputs(9272) <= 1'b1;
    layer0_outputs(9273) <= not (a and b);
    layer0_outputs(9274) <= a xor b;
    layer0_outputs(9275) <= 1'b0;
    layer0_outputs(9276) <= not b or a;
    layer0_outputs(9277) <= a and b;
    layer0_outputs(9278) <= a or b;
    layer0_outputs(9279) <= not (a and b);
    layer0_outputs(9280) <= not (a and b);
    layer0_outputs(9281) <= not (a or b);
    layer0_outputs(9282) <= not a;
    layer0_outputs(9283) <= a xor b;
    layer0_outputs(9284) <= not a;
    layer0_outputs(9285) <= not a or b;
    layer0_outputs(9286) <= b and not a;
    layer0_outputs(9287) <= 1'b1;
    layer0_outputs(9288) <= a xor b;
    layer0_outputs(9289) <= a;
    layer0_outputs(9290) <= a or b;
    layer0_outputs(9291) <= 1'b1;
    layer0_outputs(9292) <= not (a or b);
    layer0_outputs(9293) <= a and not b;
    layer0_outputs(9294) <= not (a or b);
    layer0_outputs(9295) <= not b or a;
    layer0_outputs(9296) <= not a or b;
    layer0_outputs(9297) <= not b or a;
    layer0_outputs(9298) <= not a or b;
    layer0_outputs(9299) <= a;
    layer0_outputs(9300) <= not a;
    layer0_outputs(9301) <= a or b;
    layer0_outputs(9302) <= not (a or b);
    layer0_outputs(9303) <= not a or b;
    layer0_outputs(9304) <= not (a or b);
    layer0_outputs(9305) <= not b or a;
    layer0_outputs(9306) <= a xor b;
    layer0_outputs(9307) <= not a;
    layer0_outputs(9308) <= not (a or b);
    layer0_outputs(9309) <= not b;
    layer0_outputs(9310) <= a or b;
    layer0_outputs(9311) <= a or b;
    layer0_outputs(9312) <= a xor b;
    layer0_outputs(9313) <= not (a xor b);
    layer0_outputs(9314) <= not b or a;
    layer0_outputs(9315) <= not b or a;
    layer0_outputs(9316) <= b;
    layer0_outputs(9317) <= a or b;
    layer0_outputs(9318) <= a xor b;
    layer0_outputs(9319) <= not a or b;
    layer0_outputs(9320) <= b;
    layer0_outputs(9321) <= a and b;
    layer0_outputs(9322) <= a;
    layer0_outputs(9323) <= not a;
    layer0_outputs(9324) <= not (a xor b);
    layer0_outputs(9325) <= 1'b1;
    layer0_outputs(9326) <= not (a or b);
    layer0_outputs(9327) <= not b or a;
    layer0_outputs(9328) <= b;
    layer0_outputs(9329) <= b and not a;
    layer0_outputs(9330) <= not a;
    layer0_outputs(9331) <= b;
    layer0_outputs(9332) <= not a;
    layer0_outputs(9333) <= b and not a;
    layer0_outputs(9334) <= b and not a;
    layer0_outputs(9335) <= a or b;
    layer0_outputs(9336) <= b;
    layer0_outputs(9337) <= not b or a;
    layer0_outputs(9338) <= not (a or b);
    layer0_outputs(9339) <= not a;
    layer0_outputs(9340) <= a;
    layer0_outputs(9341) <= not a or b;
    layer0_outputs(9342) <= not a;
    layer0_outputs(9343) <= a or b;
    layer0_outputs(9344) <= b;
    layer0_outputs(9345) <= not a or b;
    layer0_outputs(9346) <= a or b;
    layer0_outputs(9347) <= not (a and b);
    layer0_outputs(9348) <= a and not b;
    layer0_outputs(9349) <= not (a and b);
    layer0_outputs(9350) <= a;
    layer0_outputs(9351) <= not (a xor b);
    layer0_outputs(9352) <= not b;
    layer0_outputs(9353) <= not a or b;
    layer0_outputs(9354) <= not (a or b);
    layer0_outputs(9355) <= b and not a;
    layer0_outputs(9356) <= a xor b;
    layer0_outputs(9357) <= b;
    layer0_outputs(9358) <= 1'b0;
    layer0_outputs(9359) <= not a or b;
    layer0_outputs(9360) <= a xor b;
    layer0_outputs(9361) <= not a or b;
    layer0_outputs(9362) <= not a or b;
    layer0_outputs(9363) <= not b;
    layer0_outputs(9364) <= not (a xor b);
    layer0_outputs(9365) <= not (a xor b);
    layer0_outputs(9366) <= a or b;
    layer0_outputs(9367) <= not a;
    layer0_outputs(9368) <= not a;
    layer0_outputs(9369) <= a or b;
    layer0_outputs(9370) <= 1'b1;
    layer0_outputs(9371) <= a;
    layer0_outputs(9372) <= 1'b0;
    layer0_outputs(9373) <= b;
    layer0_outputs(9374) <= a or b;
    layer0_outputs(9375) <= not a;
    layer0_outputs(9376) <= not (a or b);
    layer0_outputs(9377) <= not a or b;
    layer0_outputs(9378) <= not b or a;
    layer0_outputs(9379) <= a and not b;
    layer0_outputs(9380) <= b;
    layer0_outputs(9381) <= not (a and b);
    layer0_outputs(9382) <= not (a and b);
    layer0_outputs(9383) <= 1'b1;
    layer0_outputs(9384) <= not b or a;
    layer0_outputs(9385) <= not (a and b);
    layer0_outputs(9386) <= not (a xor b);
    layer0_outputs(9387) <= a or b;
    layer0_outputs(9388) <= a and not b;
    layer0_outputs(9389) <= not (a xor b);
    layer0_outputs(9390) <= a and not b;
    layer0_outputs(9391) <= 1'b1;
    layer0_outputs(9392) <= a or b;
    layer0_outputs(9393) <= 1'b0;
    layer0_outputs(9394) <= a or b;
    layer0_outputs(9395) <= not b;
    layer0_outputs(9396) <= b;
    layer0_outputs(9397) <= a xor b;
    layer0_outputs(9398) <= not (a or b);
    layer0_outputs(9399) <= a and b;
    layer0_outputs(9400) <= a xor b;
    layer0_outputs(9401) <= not (a or b);
    layer0_outputs(9402) <= not b;
    layer0_outputs(9403) <= a and not b;
    layer0_outputs(9404) <= not b or a;
    layer0_outputs(9405) <= a and not b;
    layer0_outputs(9406) <= a;
    layer0_outputs(9407) <= b and not a;
    layer0_outputs(9408) <= a and not b;
    layer0_outputs(9409) <= 1'b0;
    layer0_outputs(9410) <= not (a and b);
    layer0_outputs(9411) <= not b;
    layer0_outputs(9412) <= a or b;
    layer0_outputs(9413) <= a or b;
    layer0_outputs(9414) <= not (a xor b);
    layer0_outputs(9415) <= a;
    layer0_outputs(9416) <= a and not b;
    layer0_outputs(9417) <= not (a or b);
    layer0_outputs(9418) <= not (a or b);
    layer0_outputs(9419) <= a or b;
    layer0_outputs(9420) <= 1'b1;
    layer0_outputs(9421) <= not (a or b);
    layer0_outputs(9422) <= a xor b;
    layer0_outputs(9423) <= not a;
    layer0_outputs(9424) <= not a or b;
    layer0_outputs(9425) <= a and b;
    layer0_outputs(9426) <= b;
    layer0_outputs(9427) <= b and not a;
    layer0_outputs(9428) <= a and not b;
    layer0_outputs(9429) <= not (a xor b);
    layer0_outputs(9430) <= b;
    layer0_outputs(9431) <= 1'b1;
    layer0_outputs(9432) <= b;
    layer0_outputs(9433) <= not a or b;
    layer0_outputs(9434) <= b and not a;
    layer0_outputs(9435) <= 1'b0;
    layer0_outputs(9436) <= not a;
    layer0_outputs(9437) <= not (a or b);
    layer0_outputs(9438) <= a;
    layer0_outputs(9439) <= a or b;
    layer0_outputs(9440) <= b and not a;
    layer0_outputs(9441) <= a or b;
    layer0_outputs(9442) <= not (a xor b);
    layer0_outputs(9443) <= not b or a;
    layer0_outputs(9444) <= not a or b;
    layer0_outputs(9445) <= a or b;
    layer0_outputs(9446) <= not (a xor b);
    layer0_outputs(9447) <= a or b;
    layer0_outputs(9448) <= not (a or b);
    layer0_outputs(9449) <= not a or b;
    layer0_outputs(9450) <= a;
    layer0_outputs(9451) <= not (a and b);
    layer0_outputs(9452) <= not (a or b);
    layer0_outputs(9453) <= 1'b1;
    layer0_outputs(9454) <= a xor b;
    layer0_outputs(9455) <= b and not a;
    layer0_outputs(9456) <= not (a xor b);
    layer0_outputs(9457) <= b and not a;
    layer0_outputs(9458) <= a;
    layer0_outputs(9459) <= a or b;
    layer0_outputs(9460) <= not (a or b);
    layer0_outputs(9461) <= not a or b;
    layer0_outputs(9462) <= 1'b0;
    layer0_outputs(9463) <= not a or b;
    layer0_outputs(9464) <= a xor b;
    layer0_outputs(9465) <= b;
    layer0_outputs(9466) <= not (a or b);
    layer0_outputs(9467) <= a or b;
    layer0_outputs(9468) <= a and b;
    layer0_outputs(9469) <= a and b;
    layer0_outputs(9470) <= a or b;
    layer0_outputs(9471) <= 1'b1;
    layer0_outputs(9472) <= a or b;
    layer0_outputs(9473) <= 1'b1;
    layer0_outputs(9474) <= not (a or b);
    layer0_outputs(9475) <= not (a or b);
    layer0_outputs(9476) <= not (a or b);
    layer0_outputs(9477) <= not (a or b);
    layer0_outputs(9478) <= a or b;
    layer0_outputs(9479) <= a or b;
    layer0_outputs(9480) <= not (a or b);
    layer0_outputs(9481) <= not b;
    layer0_outputs(9482) <= not (a or b);
    layer0_outputs(9483) <= not (a or b);
    layer0_outputs(9484) <= a or b;
    layer0_outputs(9485) <= a and not b;
    layer0_outputs(9486) <= a xor b;
    layer0_outputs(9487) <= a;
    layer0_outputs(9488) <= not a or b;
    layer0_outputs(9489) <= a xor b;
    layer0_outputs(9490) <= not (a and b);
    layer0_outputs(9491) <= a and not b;
    layer0_outputs(9492) <= a and b;
    layer0_outputs(9493) <= not (a xor b);
    layer0_outputs(9494) <= not a;
    layer0_outputs(9495) <= a xor b;
    layer0_outputs(9496) <= not a;
    layer0_outputs(9497) <= a and not b;
    layer0_outputs(9498) <= not b or a;
    layer0_outputs(9499) <= a and not b;
    layer0_outputs(9500) <= a;
    layer0_outputs(9501) <= b;
    layer0_outputs(9502) <= not b;
    layer0_outputs(9503) <= not (a or b);
    layer0_outputs(9504) <= a and not b;
    layer0_outputs(9505) <= b and not a;
    layer0_outputs(9506) <= not (a or b);
    layer0_outputs(9507) <= not b;
    layer0_outputs(9508) <= not b or a;
    layer0_outputs(9509) <= not a or b;
    layer0_outputs(9510) <= a xor b;
    layer0_outputs(9511) <= not b or a;
    layer0_outputs(9512) <= not (a xor b);
    layer0_outputs(9513) <= not a or b;
    layer0_outputs(9514) <= not a;
    layer0_outputs(9515) <= a xor b;
    layer0_outputs(9516) <= a xor b;
    layer0_outputs(9517) <= a xor b;
    layer0_outputs(9518) <= not (a xor b);
    layer0_outputs(9519) <= not (a or b);
    layer0_outputs(9520) <= a xor b;
    layer0_outputs(9521) <= not (a xor b);
    layer0_outputs(9522) <= not (a and b);
    layer0_outputs(9523) <= a;
    layer0_outputs(9524) <= not (a xor b);
    layer0_outputs(9525) <= b;
    layer0_outputs(9526) <= b;
    layer0_outputs(9527) <= a and not b;
    layer0_outputs(9528) <= b;
    layer0_outputs(9529) <= not b;
    layer0_outputs(9530) <= a and b;
    layer0_outputs(9531) <= not b;
    layer0_outputs(9532) <= not b;
    layer0_outputs(9533) <= b;
    layer0_outputs(9534) <= not (a or b);
    layer0_outputs(9535) <= a or b;
    layer0_outputs(9536) <= a or b;
    layer0_outputs(9537) <= b;
    layer0_outputs(9538) <= 1'b1;
    layer0_outputs(9539) <= not b;
    layer0_outputs(9540) <= not a;
    layer0_outputs(9541) <= 1'b0;
    layer0_outputs(9542) <= not (a xor b);
    layer0_outputs(9543) <= not (a or b);
    layer0_outputs(9544) <= not a;
    layer0_outputs(9545) <= a and b;
    layer0_outputs(9546) <= b and not a;
    layer0_outputs(9547) <= b and not a;
    layer0_outputs(9548) <= not b or a;
    layer0_outputs(9549) <= not a or b;
    layer0_outputs(9550) <= a or b;
    layer0_outputs(9551) <= b;
    layer0_outputs(9552) <= not b or a;
    layer0_outputs(9553) <= not (a xor b);
    layer0_outputs(9554) <= a xor b;
    layer0_outputs(9555) <= 1'b1;
    layer0_outputs(9556) <= a and not b;
    layer0_outputs(9557) <= a xor b;
    layer0_outputs(9558) <= not a;
    layer0_outputs(9559) <= b and not a;
    layer0_outputs(9560) <= a xor b;
    layer0_outputs(9561) <= not b;
    layer0_outputs(9562) <= not b or a;
    layer0_outputs(9563) <= not a;
    layer0_outputs(9564) <= a and not b;
    layer0_outputs(9565) <= not a;
    layer0_outputs(9566) <= a or b;
    layer0_outputs(9567) <= not b;
    layer0_outputs(9568) <= b and not a;
    layer0_outputs(9569) <= not a;
    layer0_outputs(9570) <= not a or b;
    layer0_outputs(9571) <= not a;
    layer0_outputs(9572) <= a or b;
    layer0_outputs(9573) <= not (a or b);
    layer0_outputs(9574) <= b;
    layer0_outputs(9575) <= not (a or b);
    layer0_outputs(9576) <= not (a or b);
    layer0_outputs(9577) <= b and not a;
    layer0_outputs(9578) <= not (a or b);
    layer0_outputs(9579) <= not a;
    layer0_outputs(9580) <= not (a or b);
    layer0_outputs(9581) <= b and not a;
    layer0_outputs(9582) <= not (a or b);
    layer0_outputs(9583) <= a and not b;
    layer0_outputs(9584) <= not b;
    layer0_outputs(9585) <= not (a or b);
    layer0_outputs(9586) <= not a or b;
    layer0_outputs(9587) <= not (a or b);
    layer0_outputs(9588) <= not (a xor b);
    layer0_outputs(9589) <= not a or b;
    layer0_outputs(9590) <= not (a and b);
    layer0_outputs(9591) <= not a or b;
    layer0_outputs(9592) <= a or b;
    layer0_outputs(9593) <= not (a and b);
    layer0_outputs(9594) <= 1'b0;
    layer0_outputs(9595) <= not b;
    layer0_outputs(9596) <= b;
    layer0_outputs(9597) <= a or b;
    layer0_outputs(9598) <= b;
    layer0_outputs(9599) <= a xor b;
    layer0_outputs(9600) <= not b or a;
    layer0_outputs(9601) <= b and not a;
    layer0_outputs(9602) <= 1'b1;
    layer0_outputs(9603) <= not (a or b);
    layer0_outputs(9604) <= not (a xor b);
    layer0_outputs(9605) <= not (a xor b);
    layer0_outputs(9606) <= b;
    layer0_outputs(9607) <= a xor b;
    layer0_outputs(9608) <= b;
    layer0_outputs(9609) <= not (a or b);
    layer0_outputs(9610) <= not (a or b);
    layer0_outputs(9611) <= not b or a;
    layer0_outputs(9612) <= a and not b;
    layer0_outputs(9613) <= not (a or b);
    layer0_outputs(9614) <= b;
    layer0_outputs(9615) <= 1'b1;
    layer0_outputs(9616) <= b;
    layer0_outputs(9617) <= not (a xor b);
    layer0_outputs(9618) <= 1'b0;
    layer0_outputs(9619) <= a and b;
    layer0_outputs(9620) <= not (a xor b);
    layer0_outputs(9621) <= b;
    layer0_outputs(9622) <= a;
    layer0_outputs(9623) <= a or b;
    layer0_outputs(9624) <= not (a or b);
    layer0_outputs(9625) <= a and b;
    layer0_outputs(9626) <= 1'b1;
    layer0_outputs(9627) <= a xor b;
    layer0_outputs(9628) <= b and not a;
    layer0_outputs(9629) <= not (a or b);
    layer0_outputs(9630) <= not (a xor b);
    layer0_outputs(9631) <= not (a xor b);
    layer0_outputs(9632) <= not b or a;
    layer0_outputs(9633) <= b and not a;
    layer0_outputs(9634) <= a or b;
    layer0_outputs(9635) <= not b;
    layer0_outputs(9636) <= not (a or b);
    layer0_outputs(9637) <= not (a or b);
    layer0_outputs(9638) <= b;
    layer0_outputs(9639) <= not b;
    layer0_outputs(9640) <= not (a xor b);
    layer0_outputs(9641) <= not a or b;
    layer0_outputs(9642) <= not (a or b);
    layer0_outputs(9643) <= not (a and b);
    layer0_outputs(9644) <= not (a and b);
    layer0_outputs(9645) <= not (a and b);
    layer0_outputs(9646) <= b;
    layer0_outputs(9647) <= a xor b;
    layer0_outputs(9648) <= not a or b;
    layer0_outputs(9649) <= b and not a;
    layer0_outputs(9650) <= b;
    layer0_outputs(9651) <= not b;
    layer0_outputs(9652) <= not (a or b);
    layer0_outputs(9653) <= b and not a;
    layer0_outputs(9654) <= a or b;
    layer0_outputs(9655) <= b;
    layer0_outputs(9656) <= not b or a;
    layer0_outputs(9657) <= not (a or b);
    layer0_outputs(9658) <= a xor b;
    layer0_outputs(9659) <= not b;
    layer0_outputs(9660) <= b and not a;
    layer0_outputs(9661) <= not a or b;
    layer0_outputs(9662) <= not b or a;
    layer0_outputs(9663) <= b;
    layer0_outputs(9664) <= a and not b;
    layer0_outputs(9665) <= not (a xor b);
    layer0_outputs(9666) <= not b or a;
    layer0_outputs(9667) <= not (a and b);
    layer0_outputs(9668) <= a xor b;
    layer0_outputs(9669) <= not (a xor b);
    layer0_outputs(9670) <= 1'b0;
    layer0_outputs(9671) <= not a;
    layer0_outputs(9672) <= not a;
    layer0_outputs(9673) <= not a;
    layer0_outputs(9674) <= b;
    layer0_outputs(9675) <= not a;
    layer0_outputs(9676) <= not (a or b);
    layer0_outputs(9677) <= not (a xor b);
    layer0_outputs(9678) <= not a;
    layer0_outputs(9679) <= not a or b;
    layer0_outputs(9680) <= not (a or b);
    layer0_outputs(9681) <= b;
    layer0_outputs(9682) <= not (a and b);
    layer0_outputs(9683) <= not b or a;
    layer0_outputs(9684) <= not (a xor b);
    layer0_outputs(9685) <= a;
    layer0_outputs(9686) <= 1'b1;
    layer0_outputs(9687) <= not (a xor b);
    layer0_outputs(9688) <= b and not a;
    layer0_outputs(9689) <= not a or b;
    layer0_outputs(9690) <= not b or a;
    layer0_outputs(9691) <= not (a or b);
    layer0_outputs(9692) <= a or b;
    layer0_outputs(9693) <= a or b;
    layer0_outputs(9694) <= b;
    layer0_outputs(9695) <= not a;
    layer0_outputs(9696) <= not b or a;
    layer0_outputs(9697) <= not (a xor b);
    layer0_outputs(9698) <= a and not b;
    layer0_outputs(9699) <= not a;
    layer0_outputs(9700) <= not b or a;
    layer0_outputs(9701) <= a xor b;
    layer0_outputs(9702) <= not (a xor b);
    layer0_outputs(9703) <= a xor b;
    layer0_outputs(9704) <= not (a xor b);
    layer0_outputs(9705) <= 1'b0;
    layer0_outputs(9706) <= a and b;
    layer0_outputs(9707) <= not (a or b);
    layer0_outputs(9708) <= a and b;
    layer0_outputs(9709) <= a and not b;
    layer0_outputs(9710) <= b;
    layer0_outputs(9711) <= not b;
    layer0_outputs(9712) <= a xor b;
    layer0_outputs(9713) <= not b or a;
    layer0_outputs(9714) <= not a;
    layer0_outputs(9715) <= a;
    layer0_outputs(9716) <= not b or a;
    layer0_outputs(9717) <= not b;
    layer0_outputs(9718) <= not b or a;
    layer0_outputs(9719) <= not (a or b);
    layer0_outputs(9720) <= a;
    layer0_outputs(9721) <= not (a xor b);
    layer0_outputs(9722) <= a xor b;
    layer0_outputs(9723) <= not (a or b);
    layer0_outputs(9724) <= a xor b;
    layer0_outputs(9725) <= a and not b;
    layer0_outputs(9726) <= a or b;
    layer0_outputs(9727) <= a or b;
    layer0_outputs(9728) <= not a or b;
    layer0_outputs(9729) <= not a;
    layer0_outputs(9730) <= b and not a;
    layer0_outputs(9731) <= not a;
    layer0_outputs(9732) <= not (a or b);
    layer0_outputs(9733) <= a;
    layer0_outputs(9734) <= a xor b;
    layer0_outputs(9735) <= a and not b;
    layer0_outputs(9736) <= a xor b;
    layer0_outputs(9737) <= not a;
    layer0_outputs(9738) <= not b or a;
    layer0_outputs(9739) <= not (a or b);
    layer0_outputs(9740) <= a xor b;
    layer0_outputs(9741) <= not (a and b);
    layer0_outputs(9742) <= a xor b;
    layer0_outputs(9743) <= a xor b;
    layer0_outputs(9744) <= not b or a;
    layer0_outputs(9745) <= not b or a;
    layer0_outputs(9746) <= not a;
    layer0_outputs(9747) <= b;
    layer0_outputs(9748) <= a or b;
    layer0_outputs(9749) <= not a;
    layer0_outputs(9750) <= not b or a;
    layer0_outputs(9751) <= not (a xor b);
    layer0_outputs(9752) <= 1'b1;
    layer0_outputs(9753) <= not a;
    layer0_outputs(9754) <= not a or b;
    layer0_outputs(9755) <= not a or b;
    layer0_outputs(9756) <= not b or a;
    layer0_outputs(9757) <= a and not b;
    layer0_outputs(9758) <= 1'b0;
    layer0_outputs(9759) <= not (a or b);
    layer0_outputs(9760) <= not a;
    layer0_outputs(9761) <= not b or a;
    layer0_outputs(9762) <= not b;
    layer0_outputs(9763) <= not b;
    layer0_outputs(9764) <= not (a xor b);
    layer0_outputs(9765) <= a;
    layer0_outputs(9766) <= not b or a;
    layer0_outputs(9767) <= b and not a;
    layer0_outputs(9768) <= 1'b0;
    layer0_outputs(9769) <= a or b;
    layer0_outputs(9770) <= a or b;
    layer0_outputs(9771) <= not (a xor b);
    layer0_outputs(9772) <= a or b;
    layer0_outputs(9773) <= not a;
    layer0_outputs(9774) <= a or b;
    layer0_outputs(9775) <= a and b;
    layer0_outputs(9776) <= b;
    layer0_outputs(9777) <= b and not a;
    layer0_outputs(9778) <= not b;
    layer0_outputs(9779) <= b;
    layer0_outputs(9780) <= not b;
    layer0_outputs(9781) <= a or b;
    layer0_outputs(9782) <= 1'b0;
    layer0_outputs(9783) <= not (a xor b);
    layer0_outputs(9784) <= 1'b1;
    layer0_outputs(9785) <= a xor b;
    layer0_outputs(9786) <= not b;
    layer0_outputs(9787) <= b;
    layer0_outputs(9788) <= not b;
    layer0_outputs(9789) <= a and b;
    layer0_outputs(9790) <= a xor b;
    layer0_outputs(9791) <= not (a xor b);
    layer0_outputs(9792) <= a;
    layer0_outputs(9793) <= not (a or b);
    layer0_outputs(9794) <= a and b;
    layer0_outputs(9795) <= 1'b0;
    layer0_outputs(9796) <= a and not b;
    layer0_outputs(9797) <= b and not a;
    layer0_outputs(9798) <= not a;
    layer0_outputs(9799) <= 1'b1;
    layer0_outputs(9800) <= not b or a;
    layer0_outputs(9801) <= a;
    layer0_outputs(9802) <= b;
    layer0_outputs(9803) <= b and not a;
    layer0_outputs(9804) <= 1'b0;
    layer0_outputs(9805) <= not a;
    layer0_outputs(9806) <= a;
    layer0_outputs(9807) <= a or b;
    layer0_outputs(9808) <= not (a and b);
    layer0_outputs(9809) <= b;
    layer0_outputs(9810) <= not b or a;
    layer0_outputs(9811) <= a and not b;
    layer0_outputs(9812) <= a or b;
    layer0_outputs(9813) <= not b;
    layer0_outputs(9814) <= a or b;
    layer0_outputs(9815) <= a and b;
    layer0_outputs(9816) <= not b;
    layer0_outputs(9817) <= not b;
    layer0_outputs(9818) <= b;
    layer0_outputs(9819) <= not (a or b);
    layer0_outputs(9820) <= not a;
    layer0_outputs(9821) <= not b or a;
    layer0_outputs(9822) <= not a or b;
    layer0_outputs(9823) <= 1'b1;
    layer0_outputs(9824) <= not (a and b);
    layer0_outputs(9825) <= not a;
    layer0_outputs(9826) <= a or b;
    layer0_outputs(9827) <= not (a or b);
    layer0_outputs(9828) <= not (a xor b);
    layer0_outputs(9829) <= a and not b;
    layer0_outputs(9830) <= a or b;
    layer0_outputs(9831) <= 1'b1;
    layer0_outputs(9832) <= not b or a;
    layer0_outputs(9833) <= 1'b1;
    layer0_outputs(9834) <= 1'b1;
    layer0_outputs(9835) <= not (a xor b);
    layer0_outputs(9836) <= not (a or b);
    layer0_outputs(9837) <= not a or b;
    layer0_outputs(9838) <= not b;
    layer0_outputs(9839) <= b and not a;
    layer0_outputs(9840) <= a and not b;
    layer0_outputs(9841) <= not a or b;
    layer0_outputs(9842) <= not (a xor b);
    layer0_outputs(9843) <= not (a and b);
    layer0_outputs(9844) <= not b or a;
    layer0_outputs(9845) <= not b or a;
    layer0_outputs(9846) <= b;
    layer0_outputs(9847) <= b;
    layer0_outputs(9848) <= not b;
    layer0_outputs(9849) <= 1'b1;
    layer0_outputs(9850) <= not b or a;
    layer0_outputs(9851) <= not (a xor b);
    layer0_outputs(9852) <= b and not a;
    layer0_outputs(9853) <= a;
    layer0_outputs(9854) <= a and not b;
    layer0_outputs(9855) <= not b or a;
    layer0_outputs(9856) <= a xor b;
    layer0_outputs(9857) <= a or b;
    layer0_outputs(9858) <= not a;
    layer0_outputs(9859) <= not a or b;
    layer0_outputs(9860) <= not (a or b);
    layer0_outputs(9861) <= not (a xor b);
    layer0_outputs(9862) <= b and not a;
    layer0_outputs(9863) <= a xor b;
    layer0_outputs(9864) <= not (a or b);
    layer0_outputs(9865) <= not b;
    layer0_outputs(9866) <= a xor b;
    layer0_outputs(9867) <= not b or a;
    layer0_outputs(9868) <= not (a xor b);
    layer0_outputs(9869) <= a or b;
    layer0_outputs(9870) <= a or b;
    layer0_outputs(9871) <= a xor b;
    layer0_outputs(9872) <= not b;
    layer0_outputs(9873) <= b;
    layer0_outputs(9874) <= a and b;
    layer0_outputs(9875) <= not a;
    layer0_outputs(9876) <= not a or b;
    layer0_outputs(9877) <= not b;
    layer0_outputs(9878) <= a or b;
    layer0_outputs(9879) <= not (a or b);
    layer0_outputs(9880) <= not (a xor b);
    layer0_outputs(9881) <= not (a or b);
    layer0_outputs(9882) <= a or b;
    layer0_outputs(9883) <= not (a or b);
    layer0_outputs(9884) <= not a;
    layer0_outputs(9885) <= a and not b;
    layer0_outputs(9886) <= not b or a;
    layer0_outputs(9887) <= a or b;
    layer0_outputs(9888) <= 1'b1;
    layer0_outputs(9889) <= a and b;
    layer0_outputs(9890) <= a;
    layer0_outputs(9891) <= a or b;
    layer0_outputs(9892) <= not (a or b);
    layer0_outputs(9893) <= not a;
    layer0_outputs(9894) <= a and b;
    layer0_outputs(9895) <= a or b;
    layer0_outputs(9896) <= not (a or b);
    layer0_outputs(9897) <= b;
    layer0_outputs(9898) <= not (a and b);
    layer0_outputs(9899) <= b;
    layer0_outputs(9900) <= not (a and b);
    layer0_outputs(9901) <= not (a or b);
    layer0_outputs(9902) <= not (a or b);
    layer0_outputs(9903) <= not (a or b);
    layer0_outputs(9904) <= a or b;
    layer0_outputs(9905) <= 1'b0;
    layer0_outputs(9906) <= not (a or b);
    layer0_outputs(9907) <= not (a or b);
    layer0_outputs(9908) <= b and not a;
    layer0_outputs(9909) <= not (a or b);
    layer0_outputs(9910) <= 1'b1;
    layer0_outputs(9911) <= not b;
    layer0_outputs(9912) <= not b or a;
    layer0_outputs(9913) <= not b or a;
    layer0_outputs(9914) <= b and not a;
    layer0_outputs(9915) <= b and not a;
    layer0_outputs(9916) <= a or b;
    layer0_outputs(9917) <= not b;
    layer0_outputs(9918) <= not (a and b);
    layer0_outputs(9919) <= a and not b;
    layer0_outputs(9920) <= b and not a;
    layer0_outputs(9921) <= a and not b;
    layer0_outputs(9922) <= 1'b1;
    layer0_outputs(9923) <= a and not b;
    layer0_outputs(9924) <= a and not b;
    layer0_outputs(9925) <= not (a and b);
    layer0_outputs(9926) <= a and not b;
    layer0_outputs(9927) <= not (a and b);
    layer0_outputs(9928) <= not (a or b);
    layer0_outputs(9929) <= a or b;
    layer0_outputs(9930) <= not (a and b);
    layer0_outputs(9931) <= not (a xor b);
    layer0_outputs(9932) <= b;
    layer0_outputs(9933) <= not b;
    layer0_outputs(9934) <= a and not b;
    layer0_outputs(9935) <= not (a xor b);
    layer0_outputs(9936) <= a xor b;
    layer0_outputs(9937) <= a or b;
    layer0_outputs(9938) <= a or b;
    layer0_outputs(9939) <= a or b;
    layer0_outputs(9940) <= a and not b;
    layer0_outputs(9941) <= not (a or b);
    layer0_outputs(9942) <= not b or a;
    layer0_outputs(9943) <= a xor b;
    layer0_outputs(9944) <= a xor b;
    layer0_outputs(9945) <= not (a and b);
    layer0_outputs(9946) <= a or b;
    layer0_outputs(9947) <= not (a or b);
    layer0_outputs(9948) <= not a;
    layer0_outputs(9949) <= 1'b1;
    layer0_outputs(9950) <= b;
    layer0_outputs(9951) <= not (a xor b);
    layer0_outputs(9952) <= not (a or b);
    layer0_outputs(9953) <= 1'b1;
    layer0_outputs(9954) <= a;
    layer0_outputs(9955) <= a;
    layer0_outputs(9956) <= a xor b;
    layer0_outputs(9957) <= 1'b1;
    layer0_outputs(9958) <= not (a or b);
    layer0_outputs(9959) <= not (a xor b);
    layer0_outputs(9960) <= a xor b;
    layer0_outputs(9961) <= a;
    layer0_outputs(9962) <= a and not b;
    layer0_outputs(9963) <= a xor b;
    layer0_outputs(9964) <= b and not a;
    layer0_outputs(9965) <= not b;
    layer0_outputs(9966) <= b;
    layer0_outputs(9967) <= not (a or b);
    layer0_outputs(9968) <= not (a or b);
    layer0_outputs(9969) <= not a;
    layer0_outputs(9970) <= a or b;
    layer0_outputs(9971) <= a;
    layer0_outputs(9972) <= not a or b;
    layer0_outputs(9973) <= a and b;
    layer0_outputs(9974) <= not a or b;
    layer0_outputs(9975) <= not b or a;
    layer0_outputs(9976) <= not b;
    layer0_outputs(9977) <= not (a or b);
    layer0_outputs(9978) <= 1'b1;
    layer0_outputs(9979) <= a xor b;
    layer0_outputs(9980) <= not b;
    layer0_outputs(9981) <= b;
    layer0_outputs(9982) <= a or b;
    layer0_outputs(9983) <= not a;
    layer0_outputs(9984) <= b;
    layer0_outputs(9985) <= a;
    layer0_outputs(9986) <= a;
    layer0_outputs(9987) <= not a or b;
    layer0_outputs(9988) <= not a;
    layer0_outputs(9989) <= b and not a;
    layer0_outputs(9990) <= 1'b0;
    layer0_outputs(9991) <= a xor b;
    layer0_outputs(9992) <= a xor b;
    layer0_outputs(9993) <= not b or a;
    layer0_outputs(9994) <= not b or a;
    layer0_outputs(9995) <= not a or b;
    layer0_outputs(9996) <= b;
    layer0_outputs(9997) <= not (a xor b);
    layer0_outputs(9998) <= a xor b;
    layer0_outputs(9999) <= not a;
    layer0_outputs(10000) <= not (a xor b);
    layer0_outputs(10001) <= not (a xor b);
    layer0_outputs(10002) <= a or b;
    layer0_outputs(10003) <= b;
    layer0_outputs(10004) <= b;
    layer0_outputs(10005) <= not (a or b);
    layer0_outputs(10006) <= not a;
    layer0_outputs(10007) <= not a or b;
    layer0_outputs(10008) <= not (a xor b);
    layer0_outputs(10009) <= a or b;
    layer0_outputs(10010) <= not b or a;
    layer0_outputs(10011) <= 1'b1;
    layer0_outputs(10012) <= not b;
    layer0_outputs(10013) <= not (a or b);
    layer0_outputs(10014) <= not b or a;
    layer0_outputs(10015) <= 1'b1;
    layer0_outputs(10016) <= not a or b;
    layer0_outputs(10017) <= a or b;
    layer0_outputs(10018) <= 1'b1;
    layer0_outputs(10019) <= not (a or b);
    layer0_outputs(10020) <= a or b;
    layer0_outputs(10021) <= a and not b;
    layer0_outputs(10022) <= not a;
    layer0_outputs(10023) <= a and not b;
    layer0_outputs(10024) <= b;
    layer0_outputs(10025) <= not b;
    layer0_outputs(10026) <= b;
    layer0_outputs(10027) <= not (a and b);
    layer0_outputs(10028) <= a xor b;
    layer0_outputs(10029) <= a xor b;
    layer0_outputs(10030) <= not a;
    layer0_outputs(10031) <= not (a and b);
    layer0_outputs(10032) <= b;
    layer0_outputs(10033) <= not b or a;
    layer0_outputs(10034) <= a xor b;
    layer0_outputs(10035) <= not (a or b);
    layer0_outputs(10036) <= b;
    layer0_outputs(10037) <= b and not a;
    layer0_outputs(10038) <= a or b;
    layer0_outputs(10039) <= not b;
    layer0_outputs(10040) <= a and not b;
    layer0_outputs(10041) <= b and not a;
    layer0_outputs(10042) <= not a;
    layer0_outputs(10043) <= b and not a;
    layer0_outputs(10044) <= a;
    layer0_outputs(10045) <= b;
    layer0_outputs(10046) <= b and not a;
    layer0_outputs(10047) <= not (a or b);
    layer0_outputs(10048) <= not a or b;
    layer0_outputs(10049) <= a xor b;
    layer0_outputs(10050) <= b;
    layer0_outputs(10051) <= not (a xor b);
    layer0_outputs(10052) <= 1'b0;
    layer0_outputs(10053) <= a and not b;
    layer0_outputs(10054) <= 1'b0;
    layer0_outputs(10055) <= a xor b;
    layer0_outputs(10056) <= not a or b;
    layer0_outputs(10057) <= not a;
    layer0_outputs(10058) <= 1'b1;
    layer0_outputs(10059) <= a xor b;
    layer0_outputs(10060) <= a and b;
    layer0_outputs(10061) <= a and not b;
    layer0_outputs(10062) <= not b;
    layer0_outputs(10063) <= b;
    layer0_outputs(10064) <= a or b;
    layer0_outputs(10065) <= b and not a;
    layer0_outputs(10066) <= not (a or b);
    layer0_outputs(10067) <= not (a or b);
    layer0_outputs(10068) <= a;
    layer0_outputs(10069) <= 1'b1;
    layer0_outputs(10070) <= not b;
    layer0_outputs(10071) <= not (a or b);
    layer0_outputs(10072) <= 1'b0;
    layer0_outputs(10073) <= not a or b;
    layer0_outputs(10074) <= a xor b;
    layer0_outputs(10075) <= not (a or b);
    layer0_outputs(10076) <= 1'b0;
    layer0_outputs(10077) <= b and not a;
    layer0_outputs(10078) <= not b;
    layer0_outputs(10079) <= not (a and b);
    layer0_outputs(10080) <= not b or a;
    layer0_outputs(10081) <= b and not a;
    layer0_outputs(10082) <= not a;
    layer0_outputs(10083) <= b;
    layer0_outputs(10084) <= a xor b;
    layer0_outputs(10085) <= not (a or b);
    layer0_outputs(10086) <= a and b;
    layer0_outputs(10087) <= a xor b;
    layer0_outputs(10088) <= b and not a;
    layer0_outputs(10089) <= not b;
    layer0_outputs(10090) <= a and not b;
    layer0_outputs(10091) <= 1'b1;
    layer0_outputs(10092) <= b;
    layer0_outputs(10093) <= 1'b0;
    layer0_outputs(10094) <= not a;
    layer0_outputs(10095) <= a;
    layer0_outputs(10096) <= not (a xor b);
    layer0_outputs(10097) <= not a;
    layer0_outputs(10098) <= b;
    layer0_outputs(10099) <= not b;
    layer0_outputs(10100) <= not (a or b);
    layer0_outputs(10101) <= b and not a;
    layer0_outputs(10102) <= not (a or b);
    layer0_outputs(10103) <= a;
    layer0_outputs(10104) <= a xor b;
    layer0_outputs(10105) <= not (a or b);
    layer0_outputs(10106) <= a or b;
    layer0_outputs(10107) <= a or b;
    layer0_outputs(10108) <= 1'b1;
    layer0_outputs(10109) <= not a;
    layer0_outputs(10110) <= not b;
    layer0_outputs(10111) <= a and b;
    layer0_outputs(10112) <= a and not b;
    layer0_outputs(10113) <= b;
    layer0_outputs(10114) <= not b or a;
    layer0_outputs(10115) <= not b;
    layer0_outputs(10116) <= b and not a;
    layer0_outputs(10117) <= a;
    layer0_outputs(10118) <= a and b;
    layer0_outputs(10119) <= not a or b;
    layer0_outputs(10120) <= not (a or b);
    layer0_outputs(10121) <= not b;
    layer0_outputs(10122) <= not a;
    layer0_outputs(10123) <= not (a or b);
    layer0_outputs(10124) <= a or b;
    layer0_outputs(10125) <= a;
    layer0_outputs(10126) <= a or b;
    layer0_outputs(10127) <= a or b;
    layer0_outputs(10128) <= a and b;
    layer0_outputs(10129) <= b;
    layer0_outputs(10130) <= not (a xor b);
    layer0_outputs(10131) <= not (a or b);
    layer0_outputs(10132) <= a and b;
    layer0_outputs(10133) <= not a or b;
    layer0_outputs(10134) <= not (a and b);
    layer0_outputs(10135) <= 1'b1;
    layer0_outputs(10136) <= a xor b;
    layer0_outputs(10137) <= not b or a;
    layer0_outputs(10138) <= b;
    layer0_outputs(10139) <= not a;
    layer0_outputs(10140) <= not b or a;
    layer0_outputs(10141) <= not (a xor b);
    layer0_outputs(10142) <= not (a xor b);
    layer0_outputs(10143) <= a and b;
    layer0_outputs(10144) <= b and not a;
    layer0_outputs(10145) <= a;
    layer0_outputs(10146) <= not (a or b);
    layer0_outputs(10147) <= not b;
    layer0_outputs(10148) <= not a or b;
    layer0_outputs(10149) <= a;
    layer0_outputs(10150) <= b and not a;
    layer0_outputs(10151) <= not a or b;
    layer0_outputs(10152) <= not (a or b);
    layer0_outputs(10153) <= a;
    layer0_outputs(10154) <= a;
    layer0_outputs(10155) <= not a;
    layer0_outputs(10156) <= a or b;
    layer0_outputs(10157) <= not a;
    layer0_outputs(10158) <= not (a or b);
    layer0_outputs(10159) <= not b;
    layer0_outputs(10160) <= b and not a;
    layer0_outputs(10161) <= b and not a;
    layer0_outputs(10162) <= a or b;
    layer0_outputs(10163) <= a;
    layer0_outputs(10164) <= a and not b;
    layer0_outputs(10165) <= a and not b;
    layer0_outputs(10166) <= not (a xor b);
    layer0_outputs(10167) <= a and not b;
    layer0_outputs(10168) <= not (a or b);
    layer0_outputs(10169) <= not (a or b);
    layer0_outputs(10170) <= b and not a;
    layer0_outputs(10171) <= b;
    layer0_outputs(10172) <= not (a or b);
    layer0_outputs(10173) <= not a or b;
    layer0_outputs(10174) <= b;
    layer0_outputs(10175) <= b;
    layer0_outputs(10176) <= b and not a;
    layer0_outputs(10177) <= a or b;
    layer0_outputs(10178) <= a xor b;
    layer0_outputs(10179) <= a;
    layer0_outputs(10180) <= b and not a;
    layer0_outputs(10181) <= not (a xor b);
    layer0_outputs(10182) <= a or b;
    layer0_outputs(10183) <= 1'b0;
    layer0_outputs(10184) <= not b;
    layer0_outputs(10185) <= not (a and b);
    layer0_outputs(10186) <= a and not b;
    layer0_outputs(10187) <= a and not b;
    layer0_outputs(10188) <= not b or a;
    layer0_outputs(10189) <= a or b;
    layer0_outputs(10190) <= b;
    layer0_outputs(10191) <= not b;
    layer0_outputs(10192) <= not (a or b);
    layer0_outputs(10193) <= a;
    layer0_outputs(10194) <= a xor b;
    layer0_outputs(10195) <= a and not b;
    layer0_outputs(10196) <= not b or a;
    layer0_outputs(10197) <= not (a or b);
    layer0_outputs(10198) <= not a or b;
    layer0_outputs(10199) <= a and not b;
    layer0_outputs(10200) <= not a;
    layer0_outputs(10201) <= a or b;
    layer0_outputs(10202) <= not b;
    layer0_outputs(10203) <= not b or a;
    layer0_outputs(10204) <= a or b;
    layer0_outputs(10205) <= a or b;
    layer0_outputs(10206) <= not b or a;
    layer0_outputs(10207) <= a;
    layer0_outputs(10208) <= not (a xor b);
    layer0_outputs(10209) <= a xor b;
    layer0_outputs(10210) <= not a or b;
    layer0_outputs(10211) <= not (a or b);
    layer0_outputs(10212) <= b;
    layer0_outputs(10213) <= not a;
    layer0_outputs(10214) <= b;
    layer0_outputs(10215) <= not a;
    layer0_outputs(10216) <= a or b;
    layer0_outputs(10217) <= a;
    layer0_outputs(10218) <= not (a xor b);
    layer0_outputs(10219) <= not b or a;
    layer0_outputs(10220) <= a and not b;
    layer0_outputs(10221) <= not (a or b);
    layer0_outputs(10222) <= 1'b0;
    layer0_outputs(10223) <= not a;
    layer0_outputs(10224) <= not (a xor b);
    layer0_outputs(10225) <= not b or a;
    layer0_outputs(10226) <= not a;
    layer0_outputs(10227) <= b and not a;
    layer0_outputs(10228) <= a;
    layer0_outputs(10229) <= b and not a;
    layer0_outputs(10230) <= 1'b0;
    layer0_outputs(10231) <= a;
    layer0_outputs(10232) <= a and not b;
    layer0_outputs(10233) <= a and not b;
    layer0_outputs(10234) <= not (a or b);
    layer0_outputs(10235) <= 1'b0;
    layer0_outputs(10236) <= a xor b;
    layer0_outputs(10237) <= a and not b;
    layer0_outputs(10238) <= 1'b1;
    layer0_outputs(10239) <= 1'b0;
    layer1_outputs(0) <= a;
    layer1_outputs(1) <= a xor b;
    layer1_outputs(2) <= a;
    layer1_outputs(3) <= b and not a;
    layer1_outputs(4) <= not (a and b);
    layer1_outputs(5) <= not a or b;
    layer1_outputs(6) <= not (a xor b);
    layer1_outputs(7) <= not (a and b);
    layer1_outputs(8) <= a;
    layer1_outputs(9) <= not (a and b);
    layer1_outputs(10) <= b and not a;
    layer1_outputs(11) <= not b;
    layer1_outputs(12) <= not (a and b);
    layer1_outputs(13) <= not b;
    layer1_outputs(14) <= not (a xor b);
    layer1_outputs(15) <= not b;
    layer1_outputs(16) <= a;
    layer1_outputs(17) <= a;
    layer1_outputs(18) <= not a;
    layer1_outputs(19) <= not (a xor b);
    layer1_outputs(20) <= not a;
    layer1_outputs(21) <= not a;
    layer1_outputs(22) <= a and b;
    layer1_outputs(23) <= a;
    layer1_outputs(24) <= not (a and b);
    layer1_outputs(25) <= not a;
    layer1_outputs(26) <= b;
    layer1_outputs(27) <= not (a and b);
    layer1_outputs(28) <= not (a or b);
    layer1_outputs(29) <= a and b;
    layer1_outputs(30) <= a;
    layer1_outputs(31) <= 1'b1;
    layer1_outputs(32) <= a and b;
    layer1_outputs(33) <= 1'b1;
    layer1_outputs(34) <= not (a xor b);
    layer1_outputs(35) <= a and b;
    layer1_outputs(36) <= 1'b0;
    layer1_outputs(37) <= not a or b;
    layer1_outputs(38) <= not a or b;
    layer1_outputs(39) <= a and b;
    layer1_outputs(40) <= not b;
    layer1_outputs(41) <= 1'b1;
    layer1_outputs(42) <= 1'b0;
    layer1_outputs(43) <= not a;
    layer1_outputs(44) <= not a;
    layer1_outputs(45) <= b and not a;
    layer1_outputs(46) <= not a or b;
    layer1_outputs(47) <= b;
    layer1_outputs(48) <= a;
    layer1_outputs(49) <= b and not a;
    layer1_outputs(50) <= a and b;
    layer1_outputs(51) <= not b or a;
    layer1_outputs(52) <= not b;
    layer1_outputs(53) <= not b or a;
    layer1_outputs(54) <= not (a or b);
    layer1_outputs(55) <= not a;
    layer1_outputs(56) <= 1'b1;
    layer1_outputs(57) <= 1'b0;
    layer1_outputs(58) <= a or b;
    layer1_outputs(59) <= not a or b;
    layer1_outputs(60) <= 1'b0;
    layer1_outputs(61) <= a;
    layer1_outputs(62) <= not b;
    layer1_outputs(63) <= a xor b;
    layer1_outputs(64) <= a;
    layer1_outputs(65) <= a xor b;
    layer1_outputs(66) <= 1'b1;
    layer1_outputs(67) <= a xor b;
    layer1_outputs(68) <= not b;
    layer1_outputs(69) <= not b or a;
    layer1_outputs(70) <= not (a or b);
    layer1_outputs(71) <= b and not a;
    layer1_outputs(72) <= 1'b0;
    layer1_outputs(73) <= 1'b0;
    layer1_outputs(74) <= not a;
    layer1_outputs(75) <= 1'b1;
    layer1_outputs(76) <= a and b;
    layer1_outputs(77) <= a;
    layer1_outputs(78) <= a and b;
    layer1_outputs(79) <= not a;
    layer1_outputs(80) <= not b;
    layer1_outputs(81) <= a;
    layer1_outputs(82) <= not b or a;
    layer1_outputs(83) <= a;
    layer1_outputs(84) <= a;
    layer1_outputs(85) <= a and not b;
    layer1_outputs(86) <= a or b;
    layer1_outputs(87) <= a and not b;
    layer1_outputs(88) <= not (a and b);
    layer1_outputs(89) <= b and not a;
    layer1_outputs(90) <= not b;
    layer1_outputs(91) <= not a;
    layer1_outputs(92) <= not (a xor b);
    layer1_outputs(93) <= not b;
    layer1_outputs(94) <= b and not a;
    layer1_outputs(95) <= not b;
    layer1_outputs(96) <= not b;
    layer1_outputs(97) <= not b or a;
    layer1_outputs(98) <= not (a and b);
    layer1_outputs(99) <= a and not b;
    layer1_outputs(100) <= a;
    layer1_outputs(101) <= 1'b1;
    layer1_outputs(102) <= not a or b;
    layer1_outputs(103) <= not a;
    layer1_outputs(104) <= 1'b1;
    layer1_outputs(105) <= a xor b;
    layer1_outputs(106) <= b;
    layer1_outputs(107) <= not (a xor b);
    layer1_outputs(108) <= a or b;
    layer1_outputs(109) <= b;
    layer1_outputs(110) <= not b or a;
    layer1_outputs(111) <= a and not b;
    layer1_outputs(112) <= not (a or b);
    layer1_outputs(113) <= not a or b;
    layer1_outputs(114) <= not a or b;
    layer1_outputs(115) <= b and not a;
    layer1_outputs(116) <= 1'b0;
    layer1_outputs(117) <= not b;
    layer1_outputs(118) <= b and not a;
    layer1_outputs(119) <= not a or b;
    layer1_outputs(120) <= 1'b0;
    layer1_outputs(121) <= not a;
    layer1_outputs(122) <= b and not a;
    layer1_outputs(123) <= a and not b;
    layer1_outputs(124) <= not (a xor b);
    layer1_outputs(125) <= not a or b;
    layer1_outputs(126) <= not (a xor b);
    layer1_outputs(127) <= not (a xor b);
    layer1_outputs(128) <= a or b;
    layer1_outputs(129) <= not a or b;
    layer1_outputs(130) <= not b;
    layer1_outputs(131) <= a or b;
    layer1_outputs(132) <= a and b;
    layer1_outputs(133) <= a or b;
    layer1_outputs(134) <= a and b;
    layer1_outputs(135) <= b and not a;
    layer1_outputs(136) <= not b;
    layer1_outputs(137) <= not a;
    layer1_outputs(138) <= not a or b;
    layer1_outputs(139) <= a or b;
    layer1_outputs(140) <= not (a and b);
    layer1_outputs(141) <= not b;
    layer1_outputs(142) <= not (a xor b);
    layer1_outputs(143) <= a and b;
    layer1_outputs(144) <= a xor b;
    layer1_outputs(145) <= not a;
    layer1_outputs(146) <= b and not a;
    layer1_outputs(147) <= b and not a;
    layer1_outputs(148) <= a and b;
    layer1_outputs(149) <= a or b;
    layer1_outputs(150) <= not a;
    layer1_outputs(151) <= not (a or b);
    layer1_outputs(152) <= not (a xor b);
    layer1_outputs(153) <= a and b;
    layer1_outputs(154) <= not a;
    layer1_outputs(155) <= not b;
    layer1_outputs(156) <= not a;
    layer1_outputs(157) <= not a or b;
    layer1_outputs(158) <= b and not a;
    layer1_outputs(159) <= not (a or b);
    layer1_outputs(160) <= not (a or b);
    layer1_outputs(161) <= a or b;
    layer1_outputs(162) <= not a;
    layer1_outputs(163) <= not b or a;
    layer1_outputs(164) <= not (a or b);
    layer1_outputs(165) <= a or b;
    layer1_outputs(166) <= a or b;
    layer1_outputs(167) <= a xor b;
    layer1_outputs(168) <= not b or a;
    layer1_outputs(169) <= a and b;
    layer1_outputs(170) <= b;
    layer1_outputs(171) <= not (a or b);
    layer1_outputs(172) <= 1'b0;
    layer1_outputs(173) <= not b;
    layer1_outputs(174) <= a or b;
    layer1_outputs(175) <= a xor b;
    layer1_outputs(176) <= not b;
    layer1_outputs(177) <= not a;
    layer1_outputs(178) <= a and not b;
    layer1_outputs(179) <= b and not a;
    layer1_outputs(180) <= not b or a;
    layer1_outputs(181) <= not b;
    layer1_outputs(182) <= not a;
    layer1_outputs(183) <= a;
    layer1_outputs(184) <= b and not a;
    layer1_outputs(185) <= a and b;
    layer1_outputs(186) <= 1'b0;
    layer1_outputs(187) <= not a or b;
    layer1_outputs(188) <= b and not a;
    layer1_outputs(189) <= a or b;
    layer1_outputs(190) <= a;
    layer1_outputs(191) <= not (a or b);
    layer1_outputs(192) <= not a or b;
    layer1_outputs(193) <= not (a xor b);
    layer1_outputs(194) <= b;
    layer1_outputs(195) <= not (a and b);
    layer1_outputs(196) <= a and b;
    layer1_outputs(197) <= not a;
    layer1_outputs(198) <= not (a and b);
    layer1_outputs(199) <= a and b;
    layer1_outputs(200) <= b;
    layer1_outputs(201) <= not b;
    layer1_outputs(202) <= not b;
    layer1_outputs(203) <= not (a or b);
    layer1_outputs(204) <= b and not a;
    layer1_outputs(205) <= not a;
    layer1_outputs(206) <= a and not b;
    layer1_outputs(207) <= b and not a;
    layer1_outputs(208) <= b;
    layer1_outputs(209) <= not a;
    layer1_outputs(210) <= a xor b;
    layer1_outputs(211) <= not a;
    layer1_outputs(212) <= not b or a;
    layer1_outputs(213) <= not (a xor b);
    layer1_outputs(214) <= 1'b1;
    layer1_outputs(215) <= b;
    layer1_outputs(216) <= not a or b;
    layer1_outputs(217) <= a;
    layer1_outputs(218) <= 1'b1;
    layer1_outputs(219) <= not (a and b);
    layer1_outputs(220) <= a;
    layer1_outputs(221) <= b;
    layer1_outputs(222) <= a;
    layer1_outputs(223) <= a xor b;
    layer1_outputs(224) <= a and not b;
    layer1_outputs(225) <= a or b;
    layer1_outputs(226) <= a and not b;
    layer1_outputs(227) <= not b;
    layer1_outputs(228) <= not (a or b);
    layer1_outputs(229) <= not a or b;
    layer1_outputs(230) <= not b;
    layer1_outputs(231) <= not (a or b);
    layer1_outputs(232) <= a and not b;
    layer1_outputs(233) <= not (a or b);
    layer1_outputs(234) <= a and b;
    layer1_outputs(235) <= a and b;
    layer1_outputs(236) <= not (a xor b);
    layer1_outputs(237) <= a and not b;
    layer1_outputs(238) <= not a or b;
    layer1_outputs(239) <= 1'b1;
    layer1_outputs(240) <= a or b;
    layer1_outputs(241) <= b and not a;
    layer1_outputs(242) <= a;
    layer1_outputs(243) <= a or b;
    layer1_outputs(244) <= not a or b;
    layer1_outputs(245) <= not (a xor b);
    layer1_outputs(246) <= a;
    layer1_outputs(247) <= b and not a;
    layer1_outputs(248) <= 1'b1;
    layer1_outputs(249) <= not (a or b);
    layer1_outputs(250) <= b and not a;
    layer1_outputs(251) <= not (a xor b);
    layer1_outputs(252) <= not b or a;
    layer1_outputs(253) <= not (a or b);
    layer1_outputs(254) <= not (a and b);
    layer1_outputs(255) <= a or b;
    layer1_outputs(256) <= not a or b;
    layer1_outputs(257) <= b and not a;
    layer1_outputs(258) <= a and not b;
    layer1_outputs(259) <= a xor b;
    layer1_outputs(260) <= not a;
    layer1_outputs(261) <= not (a and b);
    layer1_outputs(262) <= not (a xor b);
    layer1_outputs(263) <= 1'b0;
    layer1_outputs(264) <= 1'b1;
    layer1_outputs(265) <= a and not b;
    layer1_outputs(266) <= a xor b;
    layer1_outputs(267) <= not (a and b);
    layer1_outputs(268) <= a and not b;
    layer1_outputs(269) <= not a;
    layer1_outputs(270) <= 1'b1;
    layer1_outputs(271) <= not b or a;
    layer1_outputs(272) <= not b;
    layer1_outputs(273) <= a and b;
    layer1_outputs(274) <= not a or b;
    layer1_outputs(275) <= not a;
    layer1_outputs(276) <= b;
    layer1_outputs(277) <= not b;
    layer1_outputs(278) <= not (a and b);
    layer1_outputs(279) <= not a;
    layer1_outputs(280) <= not (a and b);
    layer1_outputs(281) <= not (a and b);
    layer1_outputs(282) <= not (a and b);
    layer1_outputs(283) <= 1'b1;
    layer1_outputs(284) <= b and not a;
    layer1_outputs(285) <= a;
    layer1_outputs(286) <= not a;
    layer1_outputs(287) <= a and b;
    layer1_outputs(288) <= not a;
    layer1_outputs(289) <= 1'b0;
    layer1_outputs(290) <= 1'b1;
    layer1_outputs(291) <= not a or b;
    layer1_outputs(292) <= not b;
    layer1_outputs(293) <= not a;
    layer1_outputs(294) <= not b or a;
    layer1_outputs(295) <= a;
    layer1_outputs(296) <= a;
    layer1_outputs(297) <= not (a or b);
    layer1_outputs(298) <= not (a and b);
    layer1_outputs(299) <= not (a and b);
    layer1_outputs(300) <= a and not b;
    layer1_outputs(301) <= not b or a;
    layer1_outputs(302) <= a and not b;
    layer1_outputs(303) <= 1'b0;
    layer1_outputs(304) <= a and b;
    layer1_outputs(305) <= a;
    layer1_outputs(306) <= b;
    layer1_outputs(307) <= a xor b;
    layer1_outputs(308) <= a or b;
    layer1_outputs(309) <= not (a xor b);
    layer1_outputs(310) <= a and not b;
    layer1_outputs(311) <= b;
    layer1_outputs(312) <= a or b;
    layer1_outputs(313) <= a;
    layer1_outputs(314) <= b;
    layer1_outputs(315) <= not (a or b);
    layer1_outputs(316) <= not (a or b);
    layer1_outputs(317) <= not b;
    layer1_outputs(318) <= b and not a;
    layer1_outputs(319) <= not (a and b);
    layer1_outputs(320) <= a or b;
    layer1_outputs(321) <= a and b;
    layer1_outputs(322) <= b and not a;
    layer1_outputs(323) <= not b;
    layer1_outputs(324) <= a;
    layer1_outputs(325) <= not a;
    layer1_outputs(326) <= not (a and b);
    layer1_outputs(327) <= not a;
    layer1_outputs(328) <= not a;
    layer1_outputs(329) <= not a or b;
    layer1_outputs(330) <= 1'b0;
    layer1_outputs(331) <= a and b;
    layer1_outputs(332) <= not b;
    layer1_outputs(333) <= a;
    layer1_outputs(334) <= a or b;
    layer1_outputs(335) <= a and not b;
    layer1_outputs(336) <= a;
    layer1_outputs(337) <= not b;
    layer1_outputs(338) <= not b or a;
    layer1_outputs(339) <= not b or a;
    layer1_outputs(340) <= not (a xor b);
    layer1_outputs(341) <= not a;
    layer1_outputs(342) <= not (a and b);
    layer1_outputs(343) <= b and not a;
    layer1_outputs(344) <= a or b;
    layer1_outputs(345) <= not a or b;
    layer1_outputs(346) <= not b;
    layer1_outputs(347) <= not (a or b);
    layer1_outputs(348) <= a and b;
    layer1_outputs(349) <= not b or a;
    layer1_outputs(350) <= b and not a;
    layer1_outputs(351) <= not b;
    layer1_outputs(352) <= 1'b1;
    layer1_outputs(353) <= a and not b;
    layer1_outputs(354) <= not (a xor b);
    layer1_outputs(355) <= b;
    layer1_outputs(356) <= not b or a;
    layer1_outputs(357) <= a;
    layer1_outputs(358) <= not (a xor b);
    layer1_outputs(359) <= a and b;
    layer1_outputs(360) <= not (a and b);
    layer1_outputs(361) <= a;
    layer1_outputs(362) <= not a or b;
    layer1_outputs(363) <= b;
    layer1_outputs(364) <= a and not b;
    layer1_outputs(365) <= not b or a;
    layer1_outputs(366) <= a and b;
    layer1_outputs(367) <= not (a or b);
    layer1_outputs(368) <= not (a or b);
    layer1_outputs(369) <= a and b;
    layer1_outputs(370) <= b;
    layer1_outputs(371) <= a;
    layer1_outputs(372) <= not b;
    layer1_outputs(373) <= not a or b;
    layer1_outputs(374) <= not b;
    layer1_outputs(375) <= b;
    layer1_outputs(376) <= not b;
    layer1_outputs(377) <= not (a xor b);
    layer1_outputs(378) <= not b;
    layer1_outputs(379) <= a or b;
    layer1_outputs(380) <= a;
    layer1_outputs(381) <= not (a xor b);
    layer1_outputs(382) <= b;
    layer1_outputs(383) <= not (a or b);
    layer1_outputs(384) <= not (a or b);
    layer1_outputs(385) <= not a;
    layer1_outputs(386) <= a and b;
    layer1_outputs(387) <= a and not b;
    layer1_outputs(388) <= a;
    layer1_outputs(389) <= b;
    layer1_outputs(390) <= b and not a;
    layer1_outputs(391) <= a;
    layer1_outputs(392) <= not (a and b);
    layer1_outputs(393) <= b and not a;
    layer1_outputs(394) <= not (a and b);
    layer1_outputs(395) <= a and not b;
    layer1_outputs(396) <= a and b;
    layer1_outputs(397) <= not (a and b);
    layer1_outputs(398) <= not (a or b);
    layer1_outputs(399) <= not a or b;
    layer1_outputs(400) <= not (a or b);
    layer1_outputs(401) <= 1'b0;
    layer1_outputs(402) <= a xor b;
    layer1_outputs(403) <= a or b;
    layer1_outputs(404) <= not a;
    layer1_outputs(405) <= a;
    layer1_outputs(406) <= not a;
    layer1_outputs(407) <= b;
    layer1_outputs(408) <= a;
    layer1_outputs(409) <= not (a or b);
    layer1_outputs(410) <= not a;
    layer1_outputs(411) <= b;
    layer1_outputs(412) <= not a;
    layer1_outputs(413) <= not (a xor b);
    layer1_outputs(414) <= b and not a;
    layer1_outputs(415) <= not b;
    layer1_outputs(416) <= not (a or b);
    layer1_outputs(417) <= not (a and b);
    layer1_outputs(418) <= 1'b0;
    layer1_outputs(419) <= not (a or b);
    layer1_outputs(420) <= b;
    layer1_outputs(421) <= a xor b;
    layer1_outputs(422) <= not (a xor b);
    layer1_outputs(423) <= b and not a;
    layer1_outputs(424) <= not b;
    layer1_outputs(425) <= a;
    layer1_outputs(426) <= not (a or b);
    layer1_outputs(427) <= not (a or b);
    layer1_outputs(428) <= 1'b0;
    layer1_outputs(429) <= not (a xor b);
    layer1_outputs(430) <= b;
    layer1_outputs(431) <= not b;
    layer1_outputs(432) <= not a or b;
    layer1_outputs(433) <= not b;
    layer1_outputs(434) <= a and not b;
    layer1_outputs(435) <= a;
    layer1_outputs(436) <= a and not b;
    layer1_outputs(437) <= not (a or b);
    layer1_outputs(438) <= a and not b;
    layer1_outputs(439) <= not b;
    layer1_outputs(440) <= a and b;
    layer1_outputs(441) <= a or b;
    layer1_outputs(442) <= not b;
    layer1_outputs(443) <= b and not a;
    layer1_outputs(444) <= not a or b;
    layer1_outputs(445) <= not a or b;
    layer1_outputs(446) <= a;
    layer1_outputs(447) <= not a or b;
    layer1_outputs(448) <= not (a and b);
    layer1_outputs(449) <= a;
    layer1_outputs(450) <= a or b;
    layer1_outputs(451) <= not (a and b);
    layer1_outputs(452) <= not a or b;
    layer1_outputs(453) <= 1'b0;
    layer1_outputs(454) <= not a or b;
    layer1_outputs(455) <= not a;
    layer1_outputs(456) <= not (a or b);
    layer1_outputs(457) <= a;
    layer1_outputs(458) <= not (a or b);
    layer1_outputs(459) <= not (a or b);
    layer1_outputs(460) <= not a;
    layer1_outputs(461) <= 1'b0;
    layer1_outputs(462) <= not (a and b);
    layer1_outputs(463) <= b;
    layer1_outputs(464) <= a;
    layer1_outputs(465) <= not (a or b);
    layer1_outputs(466) <= not a or b;
    layer1_outputs(467) <= a or b;
    layer1_outputs(468) <= not a or b;
    layer1_outputs(469) <= not a;
    layer1_outputs(470) <= not (a and b);
    layer1_outputs(471) <= not a or b;
    layer1_outputs(472) <= a;
    layer1_outputs(473) <= not b or a;
    layer1_outputs(474) <= a and b;
    layer1_outputs(475) <= a and b;
    layer1_outputs(476) <= b and not a;
    layer1_outputs(477) <= not (a xor b);
    layer1_outputs(478) <= not b;
    layer1_outputs(479) <= not b;
    layer1_outputs(480) <= 1'b0;
    layer1_outputs(481) <= not (a and b);
    layer1_outputs(482) <= not (a xor b);
    layer1_outputs(483) <= not a;
    layer1_outputs(484) <= not a;
    layer1_outputs(485) <= not b;
    layer1_outputs(486) <= not (a or b);
    layer1_outputs(487) <= b;
    layer1_outputs(488) <= a;
    layer1_outputs(489) <= not b;
    layer1_outputs(490) <= a xor b;
    layer1_outputs(491) <= not (a or b);
    layer1_outputs(492) <= not b or a;
    layer1_outputs(493) <= a and b;
    layer1_outputs(494) <= a;
    layer1_outputs(495) <= a and b;
    layer1_outputs(496) <= not (a or b);
    layer1_outputs(497) <= not (a or b);
    layer1_outputs(498) <= not a;
    layer1_outputs(499) <= 1'b1;
    layer1_outputs(500) <= not (a or b);
    layer1_outputs(501) <= not a or b;
    layer1_outputs(502) <= a and not b;
    layer1_outputs(503) <= not a;
    layer1_outputs(504) <= a;
    layer1_outputs(505) <= b;
    layer1_outputs(506) <= not b;
    layer1_outputs(507) <= a;
    layer1_outputs(508) <= b and not a;
    layer1_outputs(509) <= a;
    layer1_outputs(510) <= not a;
    layer1_outputs(511) <= a or b;
    layer1_outputs(512) <= b;
    layer1_outputs(513) <= a xor b;
    layer1_outputs(514) <= not b;
    layer1_outputs(515) <= b;
    layer1_outputs(516) <= not (a and b);
    layer1_outputs(517) <= a and not b;
    layer1_outputs(518) <= a xor b;
    layer1_outputs(519) <= not a;
    layer1_outputs(520) <= a;
    layer1_outputs(521) <= b and not a;
    layer1_outputs(522) <= a or b;
    layer1_outputs(523) <= not a;
    layer1_outputs(524) <= a xor b;
    layer1_outputs(525) <= not b or a;
    layer1_outputs(526) <= not (a and b);
    layer1_outputs(527) <= not (a or b);
    layer1_outputs(528) <= not (a and b);
    layer1_outputs(529) <= b and not a;
    layer1_outputs(530) <= not b or a;
    layer1_outputs(531) <= not b;
    layer1_outputs(532) <= a and not b;
    layer1_outputs(533) <= not (a and b);
    layer1_outputs(534) <= not b;
    layer1_outputs(535) <= a or b;
    layer1_outputs(536) <= not a;
    layer1_outputs(537) <= a and b;
    layer1_outputs(538) <= a and not b;
    layer1_outputs(539) <= not (a and b);
    layer1_outputs(540) <= not b;
    layer1_outputs(541) <= b;
    layer1_outputs(542) <= a or b;
    layer1_outputs(543) <= not (a and b);
    layer1_outputs(544) <= not (a or b);
    layer1_outputs(545) <= 1'b1;
    layer1_outputs(546) <= b;
    layer1_outputs(547) <= not b;
    layer1_outputs(548) <= not a;
    layer1_outputs(549) <= not (a or b);
    layer1_outputs(550) <= not b or a;
    layer1_outputs(551) <= not (a or b);
    layer1_outputs(552) <= b and not a;
    layer1_outputs(553) <= not a;
    layer1_outputs(554) <= b;
    layer1_outputs(555) <= a or b;
    layer1_outputs(556) <= b;
    layer1_outputs(557) <= b and not a;
    layer1_outputs(558) <= not (a and b);
    layer1_outputs(559) <= not a or b;
    layer1_outputs(560) <= not a;
    layer1_outputs(561) <= 1'b1;
    layer1_outputs(562) <= 1'b1;
    layer1_outputs(563) <= not a;
    layer1_outputs(564) <= a and b;
    layer1_outputs(565) <= not b or a;
    layer1_outputs(566) <= 1'b0;
    layer1_outputs(567) <= a or b;
    layer1_outputs(568) <= a and not b;
    layer1_outputs(569) <= a and not b;
    layer1_outputs(570) <= b and not a;
    layer1_outputs(571) <= not a or b;
    layer1_outputs(572) <= b;
    layer1_outputs(573) <= a or b;
    layer1_outputs(574) <= not (a xor b);
    layer1_outputs(575) <= 1'b1;
    layer1_outputs(576) <= not b or a;
    layer1_outputs(577) <= not (a or b);
    layer1_outputs(578) <= not a or b;
    layer1_outputs(579) <= b and not a;
    layer1_outputs(580) <= not a or b;
    layer1_outputs(581) <= a and b;
    layer1_outputs(582) <= a and b;
    layer1_outputs(583) <= b;
    layer1_outputs(584) <= b;
    layer1_outputs(585) <= b;
    layer1_outputs(586) <= b;
    layer1_outputs(587) <= not (a and b);
    layer1_outputs(588) <= not a or b;
    layer1_outputs(589) <= a or b;
    layer1_outputs(590) <= not (a xor b);
    layer1_outputs(591) <= not b;
    layer1_outputs(592) <= b;
    layer1_outputs(593) <= b and not a;
    layer1_outputs(594) <= not a;
    layer1_outputs(595) <= a and b;
    layer1_outputs(596) <= a;
    layer1_outputs(597) <= a;
    layer1_outputs(598) <= not b;
    layer1_outputs(599) <= b;
    layer1_outputs(600) <= not a or b;
    layer1_outputs(601) <= a and b;
    layer1_outputs(602) <= a and not b;
    layer1_outputs(603) <= not b or a;
    layer1_outputs(604) <= not b;
    layer1_outputs(605) <= not (a and b);
    layer1_outputs(606) <= a or b;
    layer1_outputs(607) <= not (a or b);
    layer1_outputs(608) <= a and not b;
    layer1_outputs(609) <= b and not a;
    layer1_outputs(610) <= not a;
    layer1_outputs(611) <= not b;
    layer1_outputs(612) <= not a;
    layer1_outputs(613) <= b and not a;
    layer1_outputs(614) <= not b;
    layer1_outputs(615) <= a xor b;
    layer1_outputs(616) <= a xor b;
    layer1_outputs(617) <= 1'b1;
    layer1_outputs(618) <= not (a or b);
    layer1_outputs(619) <= 1'b1;
    layer1_outputs(620) <= b and not a;
    layer1_outputs(621) <= not b or a;
    layer1_outputs(622) <= 1'b1;
    layer1_outputs(623) <= not (a or b);
    layer1_outputs(624) <= not (a and b);
    layer1_outputs(625) <= not a;
    layer1_outputs(626) <= b;
    layer1_outputs(627) <= not b;
    layer1_outputs(628) <= a and not b;
    layer1_outputs(629) <= not a;
    layer1_outputs(630) <= not a or b;
    layer1_outputs(631) <= a or b;
    layer1_outputs(632) <= not b;
    layer1_outputs(633) <= not b;
    layer1_outputs(634) <= a;
    layer1_outputs(635) <= not (a or b);
    layer1_outputs(636) <= b;
    layer1_outputs(637) <= b;
    layer1_outputs(638) <= not (a or b);
    layer1_outputs(639) <= b;
    layer1_outputs(640) <= not b or a;
    layer1_outputs(641) <= a;
    layer1_outputs(642) <= not a;
    layer1_outputs(643) <= not (a or b);
    layer1_outputs(644) <= a;
    layer1_outputs(645) <= a and b;
    layer1_outputs(646) <= a;
    layer1_outputs(647) <= not (a or b);
    layer1_outputs(648) <= not b;
    layer1_outputs(649) <= a or b;
    layer1_outputs(650) <= b and not a;
    layer1_outputs(651) <= not (a and b);
    layer1_outputs(652) <= not a or b;
    layer1_outputs(653) <= a;
    layer1_outputs(654) <= not (a xor b);
    layer1_outputs(655) <= not a;
    layer1_outputs(656) <= a and b;
    layer1_outputs(657) <= 1'b0;
    layer1_outputs(658) <= not a or b;
    layer1_outputs(659) <= not b or a;
    layer1_outputs(660) <= a and b;
    layer1_outputs(661) <= not a;
    layer1_outputs(662) <= a;
    layer1_outputs(663) <= not a;
    layer1_outputs(664) <= a;
    layer1_outputs(665) <= a and not b;
    layer1_outputs(666) <= a xor b;
    layer1_outputs(667) <= not (a xor b);
    layer1_outputs(668) <= b and not a;
    layer1_outputs(669) <= a;
    layer1_outputs(670) <= not (a and b);
    layer1_outputs(671) <= not a;
    layer1_outputs(672) <= a and not b;
    layer1_outputs(673) <= a;
    layer1_outputs(674) <= b and not a;
    layer1_outputs(675) <= b;
    layer1_outputs(676) <= not (a xor b);
    layer1_outputs(677) <= not a or b;
    layer1_outputs(678) <= not (a or b);
    layer1_outputs(679) <= not (a and b);
    layer1_outputs(680) <= a and not b;
    layer1_outputs(681) <= not a or b;
    layer1_outputs(682) <= not a or b;
    layer1_outputs(683) <= not a;
    layer1_outputs(684) <= a and not b;
    layer1_outputs(685) <= 1'b1;
    layer1_outputs(686) <= 1'b0;
    layer1_outputs(687) <= a or b;
    layer1_outputs(688) <= b;
    layer1_outputs(689) <= b and not a;
    layer1_outputs(690) <= not b;
    layer1_outputs(691) <= a and b;
    layer1_outputs(692) <= not b;
    layer1_outputs(693) <= b and not a;
    layer1_outputs(694) <= a;
    layer1_outputs(695) <= not a;
    layer1_outputs(696) <= 1'b0;
    layer1_outputs(697) <= a or b;
    layer1_outputs(698) <= not (a and b);
    layer1_outputs(699) <= a or b;
    layer1_outputs(700) <= not b or a;
    layer1_outputs(701) <= a;
    layer1_outputs(702) <= 1'b1;
    layer1_outputs(703) <= not a or b;
    layer1_outputs(704) <= a or b;
    layer1_outputs(705) <= a and not b;
    layer1_outputs(706) <= b;
    layer1_outputs(707) <= not (a and b);
    layer1_outputs(708) <= 1'b0;
    layer1_outputs(709) <= 1'b0;
    layer1_outputs(710) <= not b or a;
    layer1_outputs(711) <= a and b;
    layer1_outputs(712) <= not (a and b);
    layer1_outputs(713) <= a xor b;
    layer1_outputs(714) <= not (a and b);
    layer1_outputs(715) <= a xor b;
    layer1_outputs(716) <= not b;
    layer1_outputs(717) <= not (a or b);
    layer1_outputs(718) <= not b or a;
    layer1_outputs(719) <= a or b;
    layer1_outputs(720) <= not a or b;
    layer1_outputs(721) <= not a or b;
    layer1_outputs(722) <= not a;
    layer1_outputs(723) <= not b;
    layer1_outputs(724) <= not a;
    layer1_outputs(725) <= not a;
    layer1_outputs(726) <= b and not a;
    layer1_outputs(727) <= b;
    layer1_outputs(728) <= not a or b;
    layer1_outputs(729) <= a xor b;
    layer1_outputs(730) <= a and not b;
    layer1_outputs(731) <= not b;
    layer1_outputs(732) <= a;
    layer1_outputs(733) <= a xor b;
    layer1_outputs(734) <= b and not a;
    layer1_outputs(735) <= not a or b;
    layer1_outputs(736) <= not b or a;
    layer1_outputs(737) <= not a;
    layer1_outputs(738) <= a;
    layer1_outputs(739) <= not b;
    layer1_outputs(740) <= not b;
    layer1_outputs(741) <= not b or a;
    layer1_outputs(742) <= a and not b;
    layer1_outputs(743) <= not b;
    layer1_outputs(744) <= not a;
    layer1_outputs(745) <= 1'b0;
    layer1_outputs(746) <= not b;
    layer1_outputs(747) <= not a;
    layer1_outputs(748) <= a and not b;
    layer1_outputs(749) <= b;
    layer1_outputs(750) <= a and not b;
    layer1_outputs(751) <= a xor b;
    layer1_outputs(752) <= not a or b;
    layer1_outputs(753) <= a and b;
    layer1_outputs(754) <= b and not a;
    layer1_outputs(755) <= a;
    layer1_outputs(756) <= not (a or b);
    layer1_outputs(757) <= b;
    layer1_outputs(758) <= not (a and b);
    layer1_outputs(759) <= not b;
    layer1_outputs(760) <= not (a or b);
    layer1_outputs(761) <= a and not b;
    layer1_outputs(762) <= a or b;
    layer1_outputs(763) <= not a or b;
    layer1_outputs(764) <= not a;
    layer1_outputs(765) <= not (a and b);
    layer1_outputs(766) <= b;
    layer1_outputs(767) <= 1'b0;
    layer1_outputs(768) <= not a;
    layer1_outputs(769) <= a and b;
    layer1_outputs(770) <= b;
    layer1_outputs(771) <= a and b;
    layer1_outputs(772) <= a and not b;
    layer1_outputs(773) <= b;
    layer1_outputs(774) <= a and not b;
    layer1_outputs(775) <= not b or a;
    layer1_outputs(776) <= 1'b0;
    layer1_outputs(777) <= not (a and b);
    layer1_outputs(778) <= not b;
    layer1_outputs(779) <= not (a or b);
    layer1_outputs(780) <= a;
    layer1_outputs(781) <= a and not b;
    layer1_outputs(782) <= a xor b;
    layer1_outputs(783) <= not (a or b);
    layer1_outputs(784) <= not (a and b);
    layer1_outputs(785) <= b;
    layer1_outputs(786) <= not (a or b);
    layer1_outputs(787) <= not b;
    layer1_outputs(788) <= b and not a;
    layer1_outputs(789) <= b and not a;
    layer1_outputs(790) <= a and not b;
    layer1_outputs(791) <= not b or a;
    layer1_outputs(792) <= not b or a;
    layer1_outputs(793) <= not (a and b);
    layer1_outputs(794) <= not (a xor b);
    layer1_outputs(795) <= a xor b;
    layer1_outputs(796) <= not a;
    layer1_outputs(797) <= a xor b;
    layer1_outputs(798) <= not a;
    layer1_outputs(799) <= b and not a;
    layer1_outputs(800) <= not b;
    layer1_outputs(801) <= not a or b;
    layer1_outputs(802) <= b and not a;
    layer1_outputs(803) <= a and not b;
    layer1_outputs(804) <= 1'b1;
    layer1_outputs(805) <= a or b;
    layer1_outputs(806) <= b and not a;
    layer1_outputs(807) <= not b;
    layer1_outputs(808) <= a and b;
    layer1_outputs(809) <= 1'b1;
    layer1_outputs(810) <= not a;
    layer1_outputs(811) <= a;
    layer1_outputs(812) <= a and not b;
    layer1_outputs(813) <= a or b;
    layer1_outputs(814) <= a and not b;
    layer1_outputs(815) <= not a or b;
    layer1_outputs(816) <= not a or b;
    layer1_outputs(817) <= not (a xor b);
    layer1_outputs(818) <= a and b;
    layer1_outputs(819) <= not b or a;
    layer1_outputs(820) <= not a;
    layer1_outputs(821) <= not (a or b);
    layer1_outputs(822) <= a;
    layer1_outputs(823) <= a or b;
    layer1_outputs(824) <= not a;
    layer1_outputs(825) <= a or b;
    layer1_outputs(826) <= not b or a;
    layer1_outputs(827) <= b;
    layer1_outputs(828) <= not b;
    layer1_outputs(829) <= not b;
    layer1_outputs(830) <= a or b;
    layer1_outputs(831) <= not b;
    layer1_outputs(832) <= a and not b;
    layer1_outputs(833) <= a and not b;
    layer1_outputs(834) <= not a;
    layer1_outputs(835) <= a and not b;
    layer1_outputs(836) <= not b or a;
    layer1_outputs(837) <= b and not a;
    layer1_outputs(838) <= not b;
    layer1_outputs(839) <= not a;
    layer1_outputs(840) <= not (a xor b);
    layer1_outputs(841) <= b and not a;
    layer1_outputs(842) <= a;
    layer1_outputs(843) <= not (a and b);
    layer1_outputs(844) <= not (a and b);
    layer1_outputs(845) <= 1'b0;
    layer1_outputs(846) <= a;
    layer1_outputs(847) <= b;
    layer1_outputs(848) <= a and not b;
    layer1_outputs(849) <= not a or b;
    layer1_outputs(850) <= not (a or b);
    layer1_outputs(851) <= not (a or b);
    layer1_outputs(852) <= a and b;
    layer1_outputs(853) <= not a or b;
    layer1_outputs(854) <= not a;
    layer1_outputs(855) <= a;
    layer1_outputs(856) <= b and not a;
    layer1_outputs(857) <= not b;
    layer1_outputs(858) <= not a or b;
    layer1_outputs(859) <= b and not a;
    layer1_outputs(860) <= b and not a;
    layer1_outputs(861) <= not (a or b);
    layer1_outputs(862) <= a;
    layer1_outputs(863) <= not a;
    layer1_outputs(864) <= not b;
    layer1_outputs(865) <= not (a or b);
    layer1_outputs(866) <= not b or a;
    layer1_outputs(867) <= a and b;
    layer1_outputs(868) <= a and not b;
    layer1_outputs(869) <= not a or b;
    layer1_outputs(870) <= b and not a;
    layer1_outputs(871) <= not (a and b);
    layer1_outputs(872) <= not b;
    layer1_outputs(873) <= not (a and b);
    layer1_outputs(874) <= a and not b;
    layer1_outputs(875) <= not a;
    layer1_outputs(876) <= a;
    layer1_outputs(877) <= not b or a;
    layer1_outputs(878) <= not a or b;
    layer1_outputs(879) <= b and not a;
    layer1_outputs(880) <= not (a and b);
    layer1_outputs(881) <= not (a and b);
    layer1_outputs(882) <= not a or b;
    layer1_outputs(883) <= a and b;
    layer1_outputs(884) <= b;
    layer1_outputs(885) <= not b;
    layer1_outputs(886) <= a;
    layer1_outputs(887) <= not (a and b);
    layer1_outputs(888) <= a or b;
    layer1_outputs(889) <= not a;
    layer1_outputs(890) <= not (a and b);
    layer1_outputs(891) <= not a;
    layer1_outputs(892) <= 1'b1;
    layer1_outputs(893) <= a;
    layer1_outputs(894) <= a xor b;
    layer1_outputs(895) <= not b;
    layer1_outputs(896) <= not (a and b);
    layer1_outputs(897) <= not (a xor b);
    layer1_outputs(898) <= not b or a;
    layer1_outputs(899) <= a or b;
    layer1_outputs(900) <= a;
    layer1_outputs(901) <= 1'b0;
    layer1_outputs(902) <= a;
    layer1_outputs(903) <= not a;
    layer1_outputs(904) <= not (a or b);
    layer1_outputs(905) <= a xor b;
    layer1_outputs(906) <= not (a and b);
    layer1_outputs(907) <= a or b;
    layer1_outputs(908) <= not (a or b);
    layer1_outputs(909) <= not (a xor b);
    layer1_outputs(910) <= not b;
    layer1_outputs(911) <= not b or a;
    layer1_outputs(912) <= not a or b;
    layer1_outputs(913) <= b and not a;
    layer1_outputs(914) <= a or b;
    layer1_outputs(915) <= not (a and b);
    layer1_outputs(916) <= a or b;
    layer1_outputs(917) <= not (a xor b);
    layer1_outputs(918) <= b;
    layer1_outputs(919) <= not b or a;
    layer1_outputs(920) <= not b or a;
    layer1_outputs(921) <= 1'b1;
    layer1_outputs(922) <= a;
    layer1_outputs(923) <= 1'b1;
    layer1_outputs(924) <= 1'b1;
    layer1_outputs(925) <= not a;
    layer1_outputs(926) <= b;
    layer1_outputs(927) <= not (a and b);
    layer1_outputs(928) <= not a or b;
    layer1_outputs(929) <= b;
    layer1_outputs(930) <= not b;
    layer1_outputs(931) <= a and not b;
    layer1_outputs(932) <= a and b;
    layer1_outputs(933) <= not b;
    layer1_outputs(934) <= a;
    layer1_outputs(935) <= a;
    layer1_outputs(936) <= not b;
    layer1_outputs(937) <= b;
    layer1_outputs(938) <= not b;
    layer1_outputs(939) <= not b;
    layer1_outputs(940) <= 1'b1;
    layer1_outputs(941) <= a;
    layer1_outputs(942) <= a or b;
    layer1_outputs(943) <= a;
    layer1_outputs(944) <= not (a and b);
    layer1_outputs(945) <= not (a or b);
    layer1_outputs(946) <= a;
    layer1_outputs(947) <= 1'b1;
    layer1_outputs(948) <= a;
    layer1_outputs(949) <= a;
    layer1_outputs(950) <= b and not a;
    layer1_outputs(951) <= 1'b1;
    layer1_outputs(952) <= 1'b0;
    layer1_outputs(953) <= a and b;
    layer1_outputs(954) <= b and not a;
    layer1_outputs(955) <= b and not a;
    layer1_outputs(956) <= 1'b0;
    layer1_outputs(957) <= not (a and b);
    layer1_outputs(958) <= not a;
    layer1_outputs(959) <= not (a xor b);
    layer1_outputs(960) <= a and b;
    layer1_outputs(961) <= b;
    layer1_outputs(962) <= not (a and b);
    layer1_outputs(963) <= a and b;
    layer1_outputs(964) <= not a or b;
    layer1_outputs(965) <= not (a xor b);
    layer1_outputs(966) <= 1'b0;
    layer1_outputs(967) <= a and b;
    layer1_outputs(968) <= b;
    layer1_outputs(969) <= a and not b;
    layer1_outputs(970) <= not (a and b);
    layer1_outputs(971) <= not b or a;
    layer1_outputs(972) <= a xor b;
    layer1_outputs(973) <= not b or a;
    layer1_outputs(974) <= a and b;
    layer1_outputs(975) <= not a;
    layer1_outputs(976) <= not (a xor b);
    layer1_outputs(977) <= not b or a;
    layer1_outputs(978) <= a xor b;
    layer1_outputs(979) <= a xor b;
    layer1_outputs(980) <= not a;
    layer1_outputs(981) <= a xor b;
    layer1_outputs(982) <= not a;
    layer1_outputs(983) <= not a;
    layer1_outputs(984) <= not a;
    layer1_outputs(985) <= 1'b0;
    layer1_outputs(986) <= a or b;
    layer1_outputs(987) <= a and b;
    layer1_outputs(988) <= not b;
    layer1_outputs(989) <= a and not b;
    layer1_outputs(990) <= not b;
    layer1_outputs(991) <= not (a or b);
    layer1_outputs(992) <= b;
    layer1_outputs(993) <= 1'b0;
    layer1_outputs(994) <= not a;
    layer1_outputs(995) <= b;
    layer1_outputs(996) <= not (a or b);
    layer1_outputs(997) <= not (a and b);
    layer1_outputs(998) <= a;
    layer1_outputs(999) <= b and not a;
    layer1_outputs(1000) <= a;
    layer1_outputs(1001) <= not (a and b);
    layer1_outputs(1002) <= a and not b;
    layer1_outputs(1003) <= not (a or b);
    layer1_outputs(1004) <= not b or a;
    layer1_outputs(1005) <= not b;
    layer1_outputs(1006) <= not a;
    layer1_outputs(1007) <= 1'b1;
    layer1_outputs(1008) <= a and not b;
    layer1_outputs(1009) <= not b;
    layer1_outputs(1010) <= not a or b;
    layer1_outputs(1011) <= not (a and b);
    layer1_outputs(1012) <= b;
    layer1_outputs(1013) <= a;
    layer1_outputs(1014) <= not a;
    layer1_outputs(1015) <= a xor b;
    layer1_outputs(1016) <= not a;
    layer1_outputs(1017) <= 1'b1;
    layer1_outputs(1018) <= 1'b0;
    layer1_outputs(1019) <= not a;
    layer1_outputs(1020) <= not a or b;
    layer1_outputs(1021) <= a xor b;
    layer1_outputs(1022) <= not (a or b);
    layer1_outputs(1023) <= not b or a;
    layer1_outputs(1024) <= a and not b;
    layer1_outputs(1025) <= a;
    layer1_outputs(1026) <= b and not a;
    layer1_outputs(1027) <= not b or a;
    layer1_outputs(1028) <= not a or b;
    layer1_outputs(1029) <= not (a and b);
    layer1_outputs(1030) <= a and b;
    layer1_outputs(1031) <= a or b;
    layer1_outputs(1032) <= a;
    layer1_outputs(1033) <= 1'b1;
    layer1_outputs(1034) <= b;
    layer1_outputs(1035) <= 1'b1;
    layer1_outputs(1036) <= b;
    layer1_outputs(1037) <= not a;
    layer1_outputs(1038) <= a;
    layer1_outputs(1039) <= a;
    layer1_outputs(1040) <= b;
    layer1_outputs(1041) <= a and not b;
    layer1_outputs(1042) <= a and not b;
    layer1_outputs(1043) <= not a;
    layer1_outputs(1044) <= b and not a;
    layer1_outputs(1045) <= a or b;
    layer1_outputs(1046) <= a;
    layer1_outputs(1047) <= not b or a;
    layer1_outputs(1048) <= not b or a;
    layer1_outputs(1049) <= a;
    layer1_outputs(1050) <= b;
    layer1_outputs(1051) <= not (a xor b);
    layer1_outputs(1052) <= a and b;
    layer1_outputs(1053) <= 1'b0;
    layer1_outputs(1054) <= not b;
    layer1_outputs(1055) <= not a;
    layer1_outputs(1056) <= not b or a;
    layer1_outputs(1057) <= b and not a;
    layer1_outputs(1058) <= not (a or b);
    layer1_outputs(1059) <= a and not b;
    layer1_outputs(1060) <= a;
    layer1_outputs(1061) <= b;
    layer1_outputs(1062) <= b;
    layer1_outputs(1063) <= not (a and b);
    layer1_outputs(1064) <= not (a and b);
    layer1_outputs(1065) <= 1'b0;
    layer1_outputs(1066) <= not a or b;
    layer1_outputs(1067) <= not b;
    layer1_outputs(1068) <= a;
    layer1_outputs(1069) <= not a or b;
    layer1_outputs(1070) <= not a;
    layer1_outputs(1071) <= not a or b;
    layer1_outputs(1072) <= not a or b;
    layer1_outputs(1073) <= a and b;
    layer1_outputs(1074) <= b;
    layer1_outputs(1075) <= a and not b;
    layer1_outputs(1076) <= a or b;
    layer1_outputs(1077) <= b and not a;
    layer1_outputs(1078) <= a and b;
    layer1_outputs(1079) <= not a or b;
    layer1_outputs(1080) <= not b;
    layer1_outputs(1081) <= b and not a;
    layer1_outputs(1082) <= a and b;
    layer1_outputs(1083) <= a or b;
    layer1_outputs(1084) <= a and b;
    layer1_outputs(1085) <= a;
    layer1_outputs(1086) <= a and b;
    layer1_outputs(1087) <= a;
    layer1_outputs(1088) <= a or b;
    layer1_outputs(1089) <= b and not a;
    layer1_outputs(1090) <= 1'b0;
    layer1_outputs(1091) <= not (a and b);
    layer1_outputs(1092) <= 1'b1;
    layer1_outputs(1093) <= not (a and b);
    layer1_outputs(1094) <= a or b;
    layer1_outputs(1095) <= a and not b;
    layer1_outputs(1096) <= 1'b1;
    layer1_outputs(1097) <= b and not a;
    layer1_outputs(1098) <= not b or a;
    layer1_outputs(1099) <= not (a and b);
    layer1_outputs(1100) <= not (a or b);
    layer1_outputs(1101) <= not (a or b);
    layer1_outputs(1102) <= a xor b;
    layer1_outputs(1103) <= not (a and b);
    layer1_outputs(1104) <= not b or a;
    layer1_outputs(1105) <= not a or b;
    layer1_outputs(1106) <= b and not a;
    layer1_outputs(1107) <= a xor b;
    layer1_outputs(1108) <= not b;
    layer1_outputs(1109) <= not b;
    layer1_outputs(1110) <= 1'b1;
    layer1_outputs(1111) <= not (a or b);
    layer1_outputs(1112) <= not (a and b);
    layer1_outputs(1113) <= not (a and b);
    layer1_outputs(1114) <= not b;
    layer1_outputs(1115) <= a and b;
    layer1_outputs(1116) <= not a;
    layer1_outputs(1117) <= a;
    layer1_outputs(1118) <= a or b;
    layer1_outputs(1119) <= not (a xor b);
    layer1_outputs(1120) <= not a;
    layer1_outputs(1121) <= 1'b0;
    layer1_outputs(1122) <= not a;
    layer1_outputs(1123) <= a xor b;
    layer1_outputs(1124) <= not (a xor b);
    layer1_outputs(1125) <= b and not a;
    layer1_outputs(1126) <= not a or b;
    layer1_outputs(1127) <= a and not b;
    layer1_outputs(1128) <= 1'b1;
    layer1_outputs(1129) <= not a;
    layer1_outputs(1130) <= a and b;
    layer1_outputs(1131) <= not (a or b);
    layer1_outputs(1132) <= not b;
    layer1_outputs(1133) <= b;
    layer1_outputs(1134) <= a;
    layer1_outputs(1135) <= not b;
    layer1_outputs(1136) <= not a;
    layer1_outputs(1137) <= a and b;
    layer1_outputs(1138) <= a or b;
    layer1_outputs(1139) <= a or b;
    layer1_outputs(1140) <= not b;
    layer1_outputs(1141) <= a xor b;
    layer1_outputs(1142) <= not b;
    layer1_outputs(1143) <= not a;
    layer1_outputs(1144) <= not b or a;
    layer1_outputs(1145) <= a and not b;
    layer1_outputs(1146) <= not (a and b);
    layer1_outputs(1147) <= not b;
    layer1_outputs(1148) <= b and not a;
    layer1_outputs(1149) <= not a or b;
    layer1_outputs(1150) <= a or b;
    layer1_outputs(1151) <= 1'b1;
    layer1_outputs(1152) <= not (a and b);
    layer1_outputs(1153) <= not b;
    layer1_outputs(1154) <= 1'b1;
    layer1_outputs(1155) <= not a or b;
    layer1_outputs(1156) <= 1'b1;
    layer1_outputs(1157) <= a;
    layer1_outputs(1158) <= not a or b;
    layer1_outputs(1159) <= not (a or b);
    layer1_outputs(1160) <= a xor b;
    layer1_outputs(1161) <= not (a and b);
    layer1_outputs(1162) <= not (a xor b);
    layer1_outputs(1163) <= not a;
    layer1_outputs(1164) <= not b or a;
    layer1_outputs(1165) <= not a or b;
    layer1_outputs(1166) <= not b;
    layer1_outputs(1167) <= not a;
    layer1_outputs(1168) <= a and not b;
    layer1_outputs(1169) <= 1'b1;
    layer1_outputs(1170) <= b and not a;
    layer1_outputs(1171) <= a or b;
    layer1_outputs(1172) <= a and b;
    layer1_outputs(1173) <= a;
    layer1_outputs(1174) <= 1'b1;
    layer1_outputs(1175) <= not b;
    layer1_outputs(1176) <= a and b;
    layer1_outputs(1177) <= a xor b;
    layer1_outputs(1178) <= not a or b;
    layer1_outputs(1179) <= not b;
    layer1_outputs(1180) <= 1'b1;
    layer1_outputs(1181) <= a;
    layer1_outputs(1182) <= not a;
    layer1_outputs(1183) <= not (a and b);
    layer1_outputs(1184) <= not (a xor b);
    layer1_outputs(1185) <= not (a or b);
    layer1_outputs(1186) <= a and b;
    layer1_outputs(1187) <= not a;
    layer1_outputs(1188) <= a xor b;
    layer1_outputs(1189) <= b and not a;
    layer1_outputs(1190) <= a xor b;
    layer1_outputs(1191) <= a and not b;
    layer1_outputs(1192) <= not (a or b);
    layer1_outputs(1193) <= not b;
    layer1_outputs(1194) <= not a;
    layer1_outputs(1195) <= 1'b0;
    layer1_outputs(1196) <= not b;
    layer1_outputs(1197) <= not (a or b);
    layer1_outputs(1198) <= a;
    layer1_outputs(1199) <= a;
    layer1_outputs(1200) <= not (a xor b);
    layer1_outputs(1201) <= b and not a;
    layer1_outputs(1202) <= not (a xor b);
    layer1_outputs(1203) <= a;
    layer1_outputs(1204) <= not a or b;
    layer1_outputs(1205) <= a xor b;
    layer1_outputs(1206) <= not (a or b);
    layer1_outputs(1207) <= b;
    layer1_outputs(1208) <= 1'b0;
    layer1_outputs(1209) <= not (a or b);
    layer1_outputs(1210) <= not a;
    layer1_outputs(1211) <= not a;
    layer1_outputs(1212) <= b;
    layer1_outputs(1213) <= not a;
    layer1_outputs(1214) <= b and not a;
    layer1_outputs(1215) <= b;
    layer1_outputs(1216) <= not b;
    layer1_outputs(1217) <= a or b;
    layer1_outputs(1218) <= not (a or b);
    layer1_outputs(1219) <= a;
    layer1_outputs(1220) <= b;
    layer1_outputs(1221) <= a xor b;
    layer1_outputs(1222) <= 1'b0;
    layer1_outputs(1223) <= b;
    layer1_outputs(1224) <= a and not b;
    layer1_outputs(1225) <= not b;
    layer1_outputs(1226) <= a;
    layer1_outputs(1227) <= b and not a;
    layer1_outputs(1228) <= a and b;
    layer1_outputs(1229) <= not (a and b);
    layer1_outputs(1230) <= a or b;
    layer1_outputs(1231) <= a and not b;
    layer1_outputs(1232) <= not b or a;
    layer1_outputs(1233) <= not b;
    layer1_outputs(1234) <= a;
    layer1_outputs(1235) <= a or b;
    layer1_outputs(1236) <= 1'b0;
    layer1_outputs(1237) <= not a or b;
    layer1_outputs(1238) <= b;
    layer1_outputs(1239) <= a or b;
    layer1_outputs(1240) <= a and b;
    layer1_outputs(1241) <= a;
    layer1_outputs(1242) <= a;
    layer1_outputs(1243) <= a and b;
    layer1_outputs(1244) <= a;
    layer1_outputs(1245) <= not (a and b);
    layer1_outputs(1246) <= a or b;
    layer1_outputs(1247) <= b;
    layer1_outputs(1248) <= b;
    layer1_outputs(1249) <= 1'b1;
    layer1_outputs(1250) <= b and not a;
    layer1_outputs(1251) <= b and not a;
    layer1_outputs(1252) <= 1'b1;
    layer1_outputs(1253) <= not a or b;
    layer1_outputs(1254) <= not a or b;
    layer1_outputs(1255) <= not a;
    layer1_outputs(1256) <= not (a xor b);
    layer1_outputs(1257) <= not (a xor b);
    layer1_outputs(1258) <= b;
    layer1_outputs(1259) <= b;
    layer1_outputs(1260) <= b and not a;
    layer1_outputs(1261) <= 1'b1;
    layer1_outputs(1262) <= b;
    layer1_outputs(1263) <= not (a and b);
    layer1_outputs(1264) <= a;
    layer1_outputs(1265) <= a and b;
    layer1_outputs(1266) <= a;
    layer1_outputs(1267) <= not (a xor b);
    layer1_outputs(1268) <= not (a and b);
    layer1_outputs(1269) <= a and b;
    layer1_outputs(1270) <= not a;
    layer1_outputs(1271) <= not b or a;
    layer1_outputs(1272) <= a or b;
    layer1_outputs(1273) <= not (a and b);
    layer1_outputs(1274) <= not a or b;
    layer1_outputs(1275) <= a;
    layer1_outputs(1276) <= not a;
    layer1_outputs(1277) <= a or b;
    layer1_outputs(1278) <= a;
    layer1_outputs(1279) <= not (a xor b);
    layer1_outputs(1280) <= not (a and b);
    layer1_outputs(1281) <= a xor b;
    layer1_outputs(1282) <= a and not b;
    layer1_outputs(1283) <= a and b;
    layer1_outputs(1284) <= b;
    layer1_outputs(1285) <= b and not a;
    layer1_outputs(1286) <= not (a xor b);
    layer1_outputs(1287) <= not a;
    layer1_outputs(1288) <= a or b;
    layer1_outputs(1289) <= a and not b;
    layer1_outputs(1290) <= a;
    layer1_outputs(1291) <= a and not b;
    layer1_outputs(1292) <= not (a or b);
    layer1_outputs(1293) <= a;
    layer1_outputs(1294) <= 1'b0;
    layer1_outputs(1295) <= a;
    layer1_outputs(1296) <= not b;
    layer1_outputs(1297) <= not a or b;
    layer1_outputs(1298) <= not b;
    layer1_outputs(1299) <= not b;
    layer1_outputs(1300) <= a xor b;
    layer1_outputs(1301) <= b and not a;
    layer1_outputs(1302) <= a xor b;
    layer1_outputs(1303) <= a or b;
    layer1_outputs(1304) <= not (a and b);
    layer1_outputs(1305) <= not a or b;
    layer1_outputs(1306) <= not (a xor b);
    layer1_outputs(1307) <= not b or a;
    layer1_outputs(1308) <= b;
    layer1_outputs(1309) <= not (a or b);
    layer1_outputs(1310) <= not (a xor b);
    layer1_outputs(1311) <= not b;
    layer1_outputs(1312) <= not b or a;
    layer1_outputs(1313) <= a and b;
    layer1_outputs(1314) <= not a;
    layer1_outputs(1315) <= b;
    layer1_outputs(1316) <= not a;
    layer1_outputs(1317) <= not a;
    layer1_outputs(1318) <= not (a xor b);
    layer1_outputs(1319) <= not b;
    layer1_outputs(1320) <= a and not b;
    layer1_outputs(1321) <= not a or b;
    layer1_outputs(1322) <= b;
    layer1_outputs(1323) <= not (a xor b);
    layer1_outputs(1324) <= not a;
    layer1_outputs(1325) <= b and not a;
    layer1_outputs(1326) <= not (a or b);
    layer1_outputs(1327) <= a;
    layer1_outputs(1328) <= not b;
    layer1_outputs(1329) <= not b or a;
    layer1_outputs(1330) <= a xor b;
    layer1_outputs(1331) <= a or b;
    layer1_outputs(1332) <= b;
    layer1_outputs(1333) <= not (a or b);
    layer1_outputs(1334) <= a;
    layer1_outputs(1335) <= not a;
    layer1_outputs(1336) <= not b;
    layer1_outputs(1337) <= a and b;
    layer1_outputs(1338) <= not b;
    layer1_outputs(1339) <= not (a or b);
    layer1_outputs(1340) <= not a;
    layer1_outputs(1341) <= a and not b;
    layer1_outputs(1342) <= a xor b;
    layer1_outputs(1343) <= a or b;
    layer1_outputs(1344) <= not a or b;
    layer1_outputs(1345) <= b;
    layer1_outputs(1346) <= a and not b;
    layer1_outputs(1347) <= a or b;
    layer1_outputs(1348) <= b and not a;
    layer1_outputs(1349) <= b;
    layer1_outputs(1350) <= a;
    layer1_outputs(1351) <= not (a or b);
    layer1_outputs(1352) <= not a or b;
    layer1_outputs(1353) <= a;
    layer1_outputs(1354) <= a and b;
    layer1_outputs(1355) <= not (a and b);
    layer1_outputs(1356) <= b;
    layer1_outputs(1357) <= not a or b;
    layer1_outputs(1358) <= a and b;
    layer1_outputs(1359) <= b and not a;
    layer1_outputs(1360) <= a;
    layer1_outputs(1361) <= b;
    layer1_outputs(1362) <= b;
    layer1_outputs(1363) <= b;
    layer1_outputs(1364) <= b and not a;
    layer1_outputs(1365) <= a and not b;
    layer1_outputs(1366) <= not a or b;
    layer1_outputs(1367) <= not a;
    layer1_outputs(1368) <= a or b;
    layer1_outputs(1369) <= not b;
    layer1_outputs(1370) <= not a;
    layer1_outputs(1371) <= b and not a;
    layer1_outputs(1372) <= a and b;
    layer1_outputs(1373) <= a;
    layer1_outputs(1374) <= b and not a;
    layer1_outputs(1375) <= 1'b0;
    layer1_outputs(1376) <= not (a and b);
    layer1_outputs(1377) <= a and b;
    layer1_outputs(1378) <= not (a and b);
    layer1_outputs(1379) <= a xor b;
    layer1_outputs(1380) <= 1'b1;
    layer1_outputs(1381) <= a or b;
    layer1_outputs(1382) <= not b;
    layer1_outputs(1383) <= not b or a;
    layer1_outputs(1384) <= a and b;
    layer1_outputs(1385) <= b;
    layer1_outputs(1386) <= b and not a;
    layer1_outputs(1387) <= not (a and b);
    layer1_outputs(1388) <= not a or b;
    layer1_outputs(1389) <= 1'b0;
    layer1_outputs(1390) <= a and b;
    layer1_outputs(1391) <= b;
    layer1_outputs(1392) <= not b or a;
    layer1_outputs(1393) <= not (a xor b);
    layer1_outputs(1394) <= a or b;
    layer1_outputs(1395) <= b;
    layer1_outputs(1396) <= b;
    layer1_outputs(1397) <= a;
    layer1_outputs(1398) <= a;
    layer1_outputs(1399) <= not (a and b);
    layer1_outputs(1400) <= not (a and b);
    layer1_outputs(1401) <= a and not b;
    layer1_outputs(1402) <= not (a xor b);
    layer1_outputs(1403) <= a;
    layer1_outputs(1404) <= b;
    layer1_outputs(1405) <= not b;
    layer1_outputs(1406) <= 1'b1;
    layer1_outputs(1407) <= not b;
    layer1_outputs(1408) <= not a or b;
    layer1_outputs(1409) <= a;
    layer1_outputs(1410) <= 1'b0;
    layer1_outputs(1411) <= a xor b;
    layer1_outputs(1412) <= b and not a;
    layer1_outputs(1413) <= b and not a;
    layer1_outputs(1414) <= a or b;
    layer1_outputs(1415) <= a or b;
    layer1_outputs(1416) <= not (a or b);
    layer1_outputs(1417) <= b;
    layer1_outputs(1418) <= a and not b;
    layer1_outputs(1419) <= b and not a;
    layer1_outputs(1420) <= a;
    layer1_outputs(1421) <= not a;
    layer1_outputs(1422) <= 1'b0;
    layer1_outputs(1423) <= not a or b;
    layer1_outputs(1424) <= a and b;
    layer1_outputs(1425) <= 1'b0;
    layer1_outputs(1426) <= not a or b;
    layer1_outputs(1427) <= a and b;
    layer1_outputs(1428) <= not a or b;
    layer1_outputs(1429) <= b;
    layer1_outputs(1430) <= b and not a;
    layer1_outputs(1431) <= not (a and b);
    layer1_outputs(1432) <= b;
    layer1_outputs(1433) <= b;
    layer1_outputs(1434) <= 1'b1;
    layer1_outputs(1435) <= not (a or b);
    layer1_outputs(1436) <= not (a or b);
    layer1_outputs(1437) <= a or b;
    layer1_outputs(1438) <= 1'b0;
    layer1_outputs(1439) <= not b or a;
    layer1_outputs(1440) <= not (a or b);
    layer1_outputs(1441) <= 1'b1;
    layer1_outputs(1442) <= not (a and b);
    layer1_outputs(1443) <= not (a xor b);
    layer1_outputs(1444) <= b and not a;
    layer1_outputs(1445) <= a or b;
    layer1_outputs(1446) <= b;
    layer1_outputs(1447) <= not (a or b);
    layer1_outputs(1448) <= b and not a;
    layer1_outputs(1449) <= a and b;
    layer1_outputs(1450) <= a or b;
    layer1_outputs(1451) <= not a;
    layer1_outputs(1452) <= not b;
    layer1_outputs(1453) <= b;
    layer1_outputs(1454) <= a and b;
    layer1_outputs(1455) <= not (a xor b);
    layer1_outputs(1456) <= 1'b0;
    layer1_outputs(1457) <= not a or b;
    layer1_outputs(1458) <= a and b;
    layer1_outputs(1459) <= a;
    layer1_outputs(1460) <= not (a and b);
    layer1_outputs(1461) <= not a;
    layer1_outputs(1462) <= not a;
    layer1_outputs(1463) <= not (a or b);
    layer1_outputs(1464) <= b;
    layer1_outputs(1465) <= not a;
    layer1_outputs(1466) <= not (a or b);
    layer1_outputs(1467) <= not (a and b);
    layer1_outputs(1468) <= a;
    layer1_outputs(1469) <= not (a or b);
    layer1_outputs(1470) <= not a or b;
    layer1_outputs(1471) <= 1'b1;
    layer1_outputs(1472) <= 1'b1;
    layer1_outputs(1473) <= not b or a;
    layer1_outputs(1474) <= not a or b;
    layer1_outputs(1475) <= 1'b0;
    layer1_outputs(1476) <= a;
    layer1_outputs(1477) <= b;
    layer1_outputs(1478) <= a and not b;
    layer1_outputs(1479) <= b and not a;
    layer1_outputs(1480) <= not b or a;
    layer1_outputs(1481) <= 1'b0;
    layer1_outputs(1482) <= not a or b;
    layer1_outputs(1483) <= not b;
    layer1_outputs(1484) <= b;
    layer1_outputs(1485) <= not b;
    layer1_outputs(1486) <= b;
    layer1_outputs(1487) <= not b;
    layer1_outputs(1488) <= not (a or b);
    layer1_outputs(1489) <= not (a xor b);
    layer1_outputs(1490) <= 1'b1;
    layer1_outputs(1491) <= 1'b0;
    layer1_outputs(1492) <= b;
    layer1_outputs(1493) <= b;
    layer1_outputs(1494) <= not (a or b);
    layer1_outputs(1495) <= a and b;
    layer1_outputs(1496) <= a or b;
    layer1_outputs(1497) <= not a or b;
    layer1_outputs(1498) <= not (a and b);
    layer1_outputs(1499) <= not (a and b);
    layer1_outputs(1500) <= not b or a;
    layer1_outputs(1501) <= a and b;
    layer1_outputs(1502) <= not (a and b);
    layer1_outputs(1503) <= not b;
    layer1_outputs(1504) <= not a;
    layer1_outputs(1505) <= a;
    layer1_outputs(1506) <= not (a or b);
    layer1_outputs(1507) <= not (a or b);
    layer1_outputs(1508) <= not (a and b);
    layer1_outputs(1509) <= a and b;
    layer1_outputs(1510) <= b and not a;
    layer1_outputs(1511) <= not b;
    layer1_outputs(1512) <= not a;
    layer1_outputs(1513) <= not (a or b);
    layer1_outputs(1514) <= not (a or b);
    layer1_outputs(1515) <= not b;
    layer1_outputs(1516) <= b;
    layer1_outputs(1517) <= not b or a;
    layer1_outputs(1518) <= a;
    layer1_outputs(1519) <= not a;
    layer1_outputs(1520) <= a xor b;
    layer1_outputs(1521) <= not b;
    layer1_outputs(1522) <= not (a and b);
    layer1_outputs(1523) <= a;
    layer1_outputs(1524) <= 1'b1;
    layer1_outputs(1525) <= not (a and b);
    layer1_outputs(1526) <= not (a or b);
    layer1_outputs(1527) <= not (a or b);
    layer1_outputs(1528) <= a and b;
    layer1_outputs(1529) <= a and b;
    layer1_outputs(1530) <= not a;
    layer1_outputs(1531) <= a and b;
    layer1_outputs(1532) <= a xor b;
    layer1_outputs(1533) <= a;
    layer1_outputs(1534) <= a and not b;
    layer1_outputs(1535) <= a or b;
    layer1_outputs(1536) <= not b;
    layer1_outputs(1537) <= a or b;
    layer1_outputs(1538) <= not (a and b);
    layer1_outputs(1539) <= a;
    layer1_outputs(1540) <= b;
    layer1_outputs(1541) <= not (a and b);
    layer1_outputs(1542) <= not (a or b);
    layer1_outputs(1543) <= b and not a;
    layer1_outputs(1544) <= a;
    layer1_outputs(1545) <= not (a xor b);
    layer1_outputs(1546) <= a;
    layer1_outputs(1547) <= not (a or b);
    layer1_outputs(1548) <= b;
    layer1_outputs(1549) <= not (a or b);
    layer1_outputs(1550) <= not (a and b);
    layer1_outputs(1551) <= not b or a;
    layer1_outputs(1552) <= not b or a;
    layer1_outputs(1553) <= not a;
    layer1_outputs(1554) <= not a;
    layer1_outputs(1555) <= 1'b0;
    layer1_outputs(1556) <= a;
    layer1_outputs(1557) <= not (a and b);
    layer1_outputs(1558) <= not (a xor b);
    layer1_outputs(1559) <= 1'b0;
    layer1_outputs(1560) <= a or b;
    layer1_outputs(1561) <= not a;
    layer1_outputs(1562) <= b and not a;
    layer1_outputs(1563) <= not (a and b);
    layer1_outputs(1564) <= a;
    layer1_outputs(1565) <= b;
    layer1_outputs(1566) <= b;
    layer1_outputs(1567) <= a and b;
    layer1_outputs(1568) <= a xor b;
    layer1_outputs(1569) <= not (a or b);
    layer1_outputs(1570) <= a or b;
    layer1_outputs(1571) <= not (a xor b);
    layer1_outputs(1572) <= b and not a;
    layer1_outputs(1573) <= a and not b;
    layer1_outputs(1574) <= not b or a;
    layer1_outputs(1575) <= b;
    layer1_outputs(1576) <= a and b;
    layer1_outputs(1577) <= a and not b;
    layer1_outputs(1578) <= a;
    layer1_outputs(1579) <= a;
    layer1_outputs(1580) <= b and not a;
    layer1_outputs(1581) <= b and not a;
    layer1_outputs(1582) <= not (a xor b);
    layer1_outputs(1583) <= not a;
    layer1_outputs(1584) <= not (a xor b);
    layer1_outputs(1585) <= a and not b;
    layer1_outputs(1586) <= not a;
    layer1_outputs(1587) <= not b or a;
    layer1_outputs(1588) <= not a;
    layer1_outputs(1589) <= not b;
    layer1_outputs(1590) <= b and not a;
    layer1_outputs(1591) <= not (a and b);
    layer1_outputs(1592) <= not b or a;
    layer1_outputs(1593) <= not (a xor b);
    layer1_outputs(1594) <= b and not a;
    layer1_outputs(1595) <= a and b;
    layer1_outputs(1596) <= not (a and b);
    layer1_outputs(1597) <= not (a xor b);
    layer1_outputs(1598) <= not a or b;
    layer1_outputs(1599) <= b;
    layer1_outputs(1600) <= 1'b0;
    layer1_outputs(1601) <= not (a or b);
    layer1_outputs(1602) <= b;
    layer1_outputs(1603) <= a and not b;
    layer1_outputs(1604) <= not (a and b);
    layer1_outputs(1605) <= 1'b0;
    layer1_outputs(1606) <= 1'b0;
    layer1_outputs(1607) <= not (a or b);
    layer1_outputs(1608) <= b;
    layer1_outputs(1609) <= a xor b;
    layer1_outputs(1610) <= a or b;
    layer1_outputs(1611) <= a xor b;
    layer1_outputs(1612) <= not a;
    layer1_outputs(1613) <= a or b;
    layer1_outputs(1614) <= not a or b;
    layer1_outputs(1615) <= a;
    layer1_outputs(1616) <= not b;
    layer1_outputs(1617) <= not b or a;
    layer1_outputs(1618) <= not b or a;
    layer1_outputs(1619) <= not (a and b);
    layer1_outputs(1620) <= 1'b1;
    layer1_outputs(1621) <= a;
    layer1_outputs(1622) <= a and b;
    layer1_outputs(1623) <= a;
    layer1_outputs(1624) <= b and not a;
    layer1_outputs(1625) <= not a or b;
    layer1_outputs(1626) <= not a or b;
    layer1_outputs(1627) <= not a or b;
    layer1_outputs(1628) <= a and b;
    layer1_outputs(1629) <= a and not b;
    layer1_outputs(1630) <= b and not a;
    layer1_outputs(1631) <= not b;
    layer1_outputs(1632) <= a or b;
    layer1_outputs(1633) <= a and b;
    layer1_outputs(1634) <= b;
    layer1_outputs(1635) <= not (a xor b);
    layer1_outputs(1636) <= not b or a;
    layer1_outputs(1637) <= not b or a;
    layer1_outputs(1638) <= a xor b;
    layer1_outputs(1639) <= a;
    layer1_outputs(1640) <= not a or b;
    layer1_outputs(1641) <= not a;
    layer1_outputs(1642) <= b and not a;
    layer1_outputs(1643) <= not a;
    layer1_outputs(1644) <= not b;
    layer1_outputs(1645) <= not a or b;
    layer1_outputs(1646) <= a or b;
    layer1_outputs(1647) <= a and not b;
    layer1_outputs(1648) <= not (a or b);
    layer1_outputs(1649) <= 1'b1;
    layer1_outputs(1650) <= a and not b;
    layer1_outputs(1651) <= a;
    layer1_outputs(1652) <= not b;
    layer1_outputs(1653) <= a or b;
    layer1_outputs(1654) <= b and not a;
    layer1_outputs(1655) <= not (a and b);
    layer1_outputs(1656) <= not (a or b);
    layer1_outputs(1657) <= 1'b0;
    layer1_outputs(1658) <= a and not b;
    layer1_outputs(1659) <= not b or a;
    layer1_outputs(1660) <= not a;
    layer1_outputs(1661) <= a;
    layer1_outputs(1662) <= not (a and b);
    layer1_outputs(1663) <= a and b;
    layer1_outputs(1664) <= a;
    layer1_outputs(1665) <= not a or b;
    layer1_outputs(1666) <= b;
    layer1_outputs(1667) <= 1'b1;
    layer1_outputs(1668) <= not (a or b);
    layer1_outputs(1669) <= a xor b;
    layer1_outputs(1670) <= a and not b;
    layer1_outputs(1671) <= b and not a;
    layer1_outputs(1672) <= b and not a;
    layer1_outputs(1673) <= b and not a;
    layer1_outputs(1674) <= not (a and b);
    layer1_outputs(1675) <= not (a and b);
    layer1_outputs(1676) <= not b;
    layer1_outputs(1677) <= not a or b;
    layer1_outputs(1678) <= b and not a;
    layer1_outputs(1679) <= a;
    layer1_outputs(1680) <= not b;
    layer1_outputs(1681) <= not b;
    layer1_outputs(1682) <= not (a or b);
    layer1_outputs(1683) <= not b;
    layer1_outputs(1684) <= not a or b;
    layer1_outputs(1685) <= not (a or b);
    layer1_outputs(1686) <= not (a or b);
    layer1_outputs(1687) <= a xor b;
    layer1_outputs(1688) <= not (a xor b);
    layer1_outputs(1689) <= a and b;
    layer1_outputs(1690) <= b;
    layer1_outputs(1691) <= b and not a;
    layer1_outputs(1692) <= a;
    layer1_outputs(1693) <= a xor b;
    layer1_outputs(1694) <= 1'b0;
    layer1_outputs(1695) <= not (a xor b);
    layer1_outputs(1696) <= not (a or b);
    layer1_outputs(1697) <= a and not b;
    layer1_outputs(1698) <= a;
    layer1_outputs(1699) <= a xor b;
    layer1_outputs(1700) <= a or b;
    layer1_outputs(1701) <= b and not a;
    layer1_outputs(1702) <= not a or b;
    layer1_outputs(1703) <= b;
    layer1_outputs(1704) <= not a or b;
    layer1_outputs(1705) <= not (a and b);
    layer1_outputs(1706) <= b;
    layer1_outputs(1707) <= b and not a;
    layer1_outputs(1708) <= 1'b1;
    layer1_outputs(1709) <= not (a xor b);
    layer1_outputs(1710) <= b;
    layer1_outputs(1711) <= not a;
    layer1_outputs(1712) <= not (a or b);
    layer1_outputs(1713) <= a and b;
    layer1_outputs(1714) <= 1'b0;
    layer1_outputs(1715) <= a xor b;
    layer1_outputs(1716) <= b and not a;
    layer1_outputs(1717) <= a;
    layer1_outputs(1718) <= 1'b0;
    layer1_outputs(1719) <= not (a or b);
    layer1_outputs(1720) <= a xor b;
    layer1_outputs(1721) <= 1'b1;
    layer1_outputs(1722) <= a and b;
    layer1_outputs(1723) <= not a or b;
    layer1_outputs(1724) <= 1'b1;
    layer1_outputs(1725) <= not a;
    layer1_outputs(1726) <= 1'b1;
    layer1_outputs(1727) <= b;
    layer1_outputs(1728) <= b;
    layer1_outputs(1729) <= a or b;
    layer1_outputs(1730) <= 1'b0;
    layer1_outputs(1731) <= not (a or b);
    layer1_outputs(1732) <= b;
    layer1_outputs(1733) <= b and not a;
    layer1_outputs(1734) <= a and not b;
    layer1_outputs(1735) <= not (a or b);
    layer1_outputs(1736) <= 1'b0;
    layer1_outputs(1737) <= not a;
    layer1_outputs(1738) <= a;
    layer1_outputs(1739) <= b and not a;
    layer1_outputs(1740) <= b and not a;
    layer1_outputs(1741) <= not (a xor b);
    layer1_outputs(1742) <= a and b;
    layer1_outputs(1743) <= a;
    layer1_outputs(1744) <= not a;
    layer1_outputs(1745) <= a or b;
    layer1_outputs(1746) <= a and b;
    layer1_outputs(1747) <= not (a or b);
    layer1_outputs(1748) <= b;
    layer1_outputs(1749) <= b;
    layer1_outputs(1750) <= b and not a;
    layer1_outputs(1751) <= not b or a;
    layer1_outputs(1752) <= a and b;
    layer1_outputs(1753) <= not a or b;
    layer1_outputs(1754) <= not a;
    layer1_outputs(1755) <= b and not a;
    layer1_outputs(1756) <= a;
    layer1_outputs(1757) <= a xor b;
    layer1_outputs(1758) <= not (a or b);
    layer1_outputs(1759) <= b;
    layer1_outputs(1760) <= b and not a;
    layer1_outputs(1761) <= not (a and b);
    layer1_outputs(1762) <= not b or a;
    layer1_outputs(1763) <= b;
    layer1_outputs(1764) <= not b or a;
    layer1_outputs(1765) <= not (a and b);
    layer1_outputs(1766) <= not a;
    layer1_outputs(1767) <= not b;
    layer1_outputs(1768) <= b and not a;
    layer1_outputs(1769) <= a and not b;
    layer1_outputs(1770) <= not b;
    layer1_outputs(1771) <= a or b;
    layer1_outputs(1772) <= a and b;
    layer1_outputs(1773) <= b and not a;
    layer1_outputs(1774) <= 1'b1;
    layer1_outputs(1775) <= b;
    layer1_outputs(1776) <= not b or a;
    layer1_outputs(1777) <= a or b;
    layer1_outputs(1778) <= 1'b0;
    layer1_outputs(1779) <= 1'b0;
    layer1_outputs(1780) <= b;
    layer1_outputs(1781) <= a and b;
    layer1_outputs(1782) <= not b or a;
    layer1_outputs(1783) <= a or b;
    layer1_outputs(1784) <= a or b;
    layer1_outputs(1785) <= a and b;
    layer1_outputs(1786) <= a;
    layer1_outputs(1787) <= not a;
    layer1_outputs(1788) <= 1'b0;
    layer1_outputs(1789) <= a;
    layer1_outputs(1790) <= a or b;
    layer1_outputs(1791) <= b and not a;
    layer1_outputs(1792) <= a;
    layer1_outputs(1793) <= not a or b;
    layer1_outputs(1794) <= not a;
    layer1_outputs(1795) <= b and not a;
    layer1_outputs(1796) <= b and not a;
    layer1_outputs(1797) <= not b;
    layer1_outputs(1798) <= not (a xor b);
    layer1_outputs(1799) <= a and not b;
    layer1_outputs(1800) <= not b;
    layer1_outputs(1801) <= a;
    layer1_outputs(1802) <= a;
    layer1_outputs(1803) <= a;
    layer1_outputs(1804) <= a;
    layer1_outputs(1805) <= not b or a;
    layer1_outputs(1806) <= not b;
    layer1_outputs(1807) <= not a or b;
    layer1_outputs(1808) <= not b;
    layer1_outputs(1809) <= a and not b;
    layer1_outputs(1810) <= b;
    layer1_outputs(1811) <= not (a and b);
    layer1_outputs(1812) <= a and not b;
    layer1_outputs(1813) <= not b or a;
    layer1_outputs(1814) <= not (a or b);
    layer1_outputs(1815) <= b;
    layer1_outputs(1816) <= a;
    layer1_outputs(1817) <= a;
    layer1_outputs(1818) <= not b or a;
    layer1_outputs(1819) <= not a or b;
    layer1_outputs(1820) <= not (a or b);
    layer1_outputs(1821) <= 1'b0;
    layer1_outputs(1822) <= not (a and b);
    layer1_outputs(1823) <= b;
    layer1_outputs(1824) <= not (a and b);
    layer1_outputs(1825) <= a and b;
    layer1_outputs(1826) <= not a or b;
    layer1_outputs(1827) <= not b or a;
    layer1_outputs(1828) <= b and not a;
    layer1_outputs(1829) <= 1'b1;
    layer1_outputs(1830) <= not (a xor b);
    layer1_outputs(1831) <= not (a and b);
    layer1_outputs(1832) <= a xor b;
    layer1_outputs(1833) <= not b;
    layer1_outputs(1834) <= a and b;
    layer1_outputs(1835) <= a xor b;
    layer1_outputs(1836) <= not (a xor b);
    layer1_outputs(1837) <= not b;
    layer1_outputs(1838) <= not a;
    layer1_outputs(1839) <= a xor b;
    layer1_outputs(1840) <= not a;
    layer1_outputs(1841) <= b;
    layer1_outputs(1842) <= not b;
    layer1_outputs(1843) <= a or b;
    layer1_outputs(1844) <= a or b;
    layer1_outputs(1845) <= not (a and b);
    layer1_outputs(1846) <= a;
    layer1_outputs(1847) <= b;
    layer1_outputs(1848) <= a or b;
    layer1_outputs(1849) <= 1'b0;
    layer1_outputs(1850) <= not a or b;
    layer1_outputs(1851) <= not b;
    layer1_outputs(1852) <= 1'b0;
    layer1_outputs(1853) <= b;
    layer1_outputs(1854) <= a;
    layer1_outputs(1855) <= b and not a;
    layer1_outputs(1856) <= not b or a;
    layer1_outputs(1857) <= not a;
    layer1_outputs(1858) <= not (a and b);
    layer1_outputs(1859) <= not (a and b);
    layer1_outputs(1860) <= not (a xor b);
    layer1_outputs(1861) <= a and b;
    layer1_outputs(1862) <= 1'b1;
    layer1_outputs(1863) <= 1'b1;
    layer1_outputs(1864) <= a and b;
    layer1_outputs(1865) <= 1'b0;
    layer1_outputs(1866) <= a or b;
    layer1_outputs(1867) <= not b or a;
    layer1_outputs(1868) <= 1'b1;
    layer1_outputs(1869) <= a;
    layer1_outputs(1870) <= not b or a;
    layer1_outputs(1871) <= not (a or b);
    layer1_outputs(1872) <= not (a xor b);
    layer1_outputs(1873) <= not b or a;
    layer1_outputs(1874) <= 1'b0;
    layer1_outputs(1875) <= b;
    layer1_outputs(1876) <= a and not b;
    layer1_outputs(1877) <= not b or a;
    layer1_outputs(1878) <= not (a and b);
    layer1_outputs(1879) <= a or b;
    layer1_outputs(1880) <= not b;
    layer1_outputs(1881) <= 1'b1;
    layer1_outputs(1882) <= a;
    layer1_outputs(1883) <= a and b;
    layer1_outputs(1884) <= not b or a;
    layer1_outputs(1885) <= not a;
    layer1_outputs(1886) <= not a or b;
    layer1_outputs(1887) <= a and b;
    layer1_outputs(1888) <= not b;
    layer1_outputs(1889) <= not (a and b);
    layer1_outputs(1890) <= not (a or b);
    layer1_outputs(1891) <= not (a xor b);
    layer1_outputs(1892) <= a and not b;
    layer1_outputs(1893) <= 1'b1;
    layer1_outputs(1894) <= not b;
    layer1_outputs(1895) <= not b;
    layer1_outputs(1896) <= a and not b;
    layer1_outputs(1897) <= not b or a;
    layer1_outputs(1898) <= not a;
    layer1_outputs(1899) <= not a;
    layer1_outputs(1900) <= not b;
    layer1_outputs(1901) <= not a;
    layer1_outputs(1902) <= not b;
    layer1_outputs(1903) <= not a or b;
    layer1_outputs(1904) <= 1'b1;
    layer1_outputs(1905) <= not b;
    layer1_outputs(1906) <= a xor b;
    layer1_outputs(1907) <= 1'b1;
    layer1_outputs(1908) <= b and not a;
    layer1_outputs(1909) <= not (a and b);
    layer1_outputs(1910) <= not (a or b);
    layer1_outputs(1911) <= a;
    layer1_outputs(1912) <= 1'b1;
    layer1_outputs(1913) <= not a;
    layer1_outputs(1914) <= b and not a;
    layer1_outputs(1915) <= 1'b1;
    layer1_outputs(1916) <= a and not b;
    layer1_outputs(1917) <= b and not a;
    layer1_outputs(1918) <= a and b;
    layer1_outputs(1919) <= not (a or b);
    layer1_outputs(1920) <= a or b;
    layer1_outputs(1921) <= not b;
    layer1_outputs(1922) <= b and not a;
    layer1_outputs(1923) <= not b or a;
    layer1_outputs(1924) <= 1'b0;
    layer1_outputs(1925) <= not (a or b);
    layer1_outputs(1926) <= b and not a;
    layer1_outputs(1927) <= not b or a;
    layer1_outputs(1928) <= b and not a;
    layer1_outputs(1929) <= b;
    layer1_outputs(1930) <= not (a or b);
    layer1_outputs(1931) <= 1'b1;
    layer1_outputs(1932) <= not (a and b);
    layer1_outputs(1933) <= a and not b;
    layer1_outputs(1934) <= b;
    layer1_outputs(1935) <= a;
    layer1_outputs(1936) <= a and b;
    layer1_outputs(1937) <= not a;
    layer1_outputs(1938) <= not b;
    layer1_outputs(1939) <= a xor b;
    layer1_outputs(1940) <= b and not a;
    layer1_outputs(1941) <= 1'b1;
    layer1_outputs(1942) <= b;
    layer1_outputs(1943) <= not (a and b);
    layer1_outputs(1944) <= a xor b;
    layer1_outputs(1945) <= a and not b;
    layer1_outputs(1946) <= b and not a;
    layer1_outputs(1947) <= not (a xor b);
    layer1_outputs(1948) <= not (a and b);
    layer1_outputs(1949) <= a and b;
    layer1_outputs(1950) <= a;
    layer1_outputs(1951) <= not (a or b);
    layer1_outputs(1952) <= a;
    layer1_outputs(1953) <= a;
    layer1_outputs(1954) <= a;
    layer1_outputs(1955) <= a and not b;
    layer1_outputs(1956) <= not (a and b);
    layer1_outputs(1957) <= not a or b;
    layer1_outputs(1958) <= not (a or b);
    layer1_outputs(1959) <= not b or a;
    layer1_outputs(1960) <= not (a or b);
    layer1_outputs(1961) <= b and not a;
    layer1_outputs(1962) <= not b;
    layer1_outputs(1963) <= not (a or b);
    layer1_outputs(1964) <= 1'b0;
    layer1_outputs(1965) <= not (a xor b);
    layer1_outputs(1966) <= a and b;
    layer1_outputs(1967) <= b and not a;
    layer1_outputs(1968) <= not b or a;
    layer1_outputs(1969) <= not (a or b);
    layer1_outputs(1970) <= b;
    layer1_outputs(1971) <= 1'b1;
    layer1_outputs(1972) <= not a or b;
    layer1_outputs(1973) <= a and not b;
    layer1_outputs(1974) <= not a;
    layer1_outputs(1975) <= a;
    layer1_outputs(1976) <= b and not a;
    layer1_outputs(1977) <= not (a and b);
    layer1_outputs(1978) <= a and not b;
    layer1_outputs(1979) <= a and not b;
    layer1_outputs(1980) <= a or b;
    layer1_outputs(1981) <= not a;
    layer1_outputs(1982) <= 1'b0;
    layer1_outputs(1983) <= not b or a;
    layer1_outputs(1984) <= 1'b1;
    layer1_outputs(1985) <= not b or a;
    layer1_outputs(1986) <= not (a and b);
    layer1_outputs(1987) <= a and b;
    layer1_outputs(1988) <= not b;
    layer1_outputs(1989) <= not a;
    layer1_outputs(1990) <= not a or b;
    layer1_outputs(1991) <= b and not a;
    layer1_outputs(1992) <= a and b;
    layer1_outputs(1993) <= a xor b;
    layer1_outputs(1994) <= a and b;
    layer1_outputs(1995) <= not b or a;
    layer1_outputs(1996) <= not a;
    layer1_outputs(1997) <= a xor b;
    layer1_outputs(1998) <= a xor b;
    layer1_outputs(1999) <= not a or b;
    layer1_outputs(2000) <= not b or a;
    layer1_outputs(2001) <= not a or b;
    layer1_outputs(2002) <= not b or a;
    layer1_outputs(2003) <= not (a and b);
    layer1_outputs(2004) <= 1'b0;
    layer1_outputs(2005) <= a and not b;
    layer1_outputs(2006) <= a xor b;
    layer1_outputs(2007) <= 1'b0;
    layer1_outputs(2008) <= a or b;
    layer1_outputs(2009) <= a and not b;
    layer1_outputs(2010) <= b and not a;
    layer1_outputs(2011) <= not a;
    layer1_outputs(2012) <= b;
    layer1_outputs(2013) <= a and b;
    layer1_outputs(2014) <= a;
    layer1_outputs(2015) <= a;
    layer1_outputs(2016) <= 1'b1;
    layer1_outputs(2017) <= a;
    layer1_outputs(2018) <= not b or a;
    layer1_outputs(2019) <= not (a and b);
    layer1_outputs(2020) <= 1'b1;
    layer1_outputs(2021) <= not (a or b);
    layer1_outputs(2022) <= b;
    layer1_outputs(2023) <= a or b;
    layer1_outputs(2024) <= not (a and b);
    layer1_outputs(2025) <= not (a and b);
    layer1_outputs(2026) <= not (a and b);
    layer1_outputs(2027) <= a and not b;
    layer1_outputs(2028) <= a or b;
    layer1_outputs(2029) <= b;
    layer1_outputs(2030) <= not (a and b);
    layer1_outputs(2031) <= a xor b;
    layer1_outputs(2032) <= b;
    layer1_outputs(2033) <= a and not b;
    layer1_outputs(2034) <= b and not a;
    layer1_outputs(2035) <= a xor b;
    layer1_outputs(2036) <= b;
    layer1_outputs(2037) <= a xor b;
    layer1_outputs(2038) <= a and b;
    layer1_outputs(2039) <= b;
    layer1_outputs(2040) <= not b;
    layer1_outputs(2041) <= not (a or b);
    layer1_outputs(2042) <= a and b;
    layer1_outputs(2043) <= not a;
    layer1_outputs(2044) <= not (a and b);
    layer1_outputs(2045) <= not b;
    layer1_outputs(2046) <= not b or a;
    layer1_outputs(2047) <= a or b;
    layer1_outputs(2048) <= a and not b;
    layer1_outputs(2049) <= not (a and b);
    layer1_outputs(2050) <= not (a or b);
    layer1_outputs(2051) <= not (a xor b);
    layer1_outputs(2052) <= a or b;
    layer1_outputs(2053) <= b;
    layer1_outputs(2054) <= b and not a;
    layer1_outputs(2055) <= b;
    layer1_outputs(2056) <= b and not a;
    layer1_outputs(2057) <= a and not b;
    layer1_outputs(2058) <= a xor b;
    layer1_outputs(2059) <= not (a and b);
    layer1_outputs(2060) <= not (a or b);
    layer1_outputs(2061) <= 1'b1;
    layer1_outputs(2062) <= not (a or b);
    layer1_outputs(2063) <= not b;
    layer1_outputs(2064) <= not (a and b);
    layer1_outputs(2065) <= a xor b;
    layer1_outputs(2066) <= not (a or b);
    layer1_outputs(2067) <= not a or b;
    layer1_outputs(2068) <= a xor b;
    layer1_outputs(2069) <= not (a xor b);
    layer1_outputs(2070) <= not a or b;
    layer1_outputs(2071) <= not b;
    layer1_outputs(2072) <= a;
    layer1_outputs(2073) <= a;
    layer1_outputs(2074) <= a and not b;
    layer1_outputs(2075) <= not b;
    layer1_outputs(2076) <= a xor b;
    layer1_outputs(2077) <= not a or b;
    layer1_outputs(2078) <= not (a and b);
    layer1_outputs(2079) <= not b or a;
    layer1_outputs(2080) <= a and not b;
    layer1_outputs(2081) <= not (a or b);
    layer1_outputs(2082) <= not b or a;
    layer1_outputs(2083) <= 1'b0;
    layer1_outputs(2084) <= a xor b;
    layer1_outputs(2085) <= b;
    layer1_outputs(2086) <= a;
    layer1_outputs(2087) <= not a;
    layer1_outputs(2088) <= not b;
    layer1_outputs(2089) <= a and b;
    layer1_outputs(2090) <= not a or b;
    layer1_outputs(2091) <= not (a xor b);
    layer1_outputs(2092) <= a xor b;
    layer1_outputs(2093) <= a and b;
    layer1_outputs(2094) <= not a or b;
    layer1_outputs(2095) <= 1'b0;
    layer1_outputs(2096) <= a xor b;
    layer1_outputs(2097) <= not (a or b);
    layer1_outputs(2098) <= not b;
    layer1_outputs(2099) <= not a or b;
    layer1_outputs(2100) <= not b or a;
    layer1_outputs(2101) <= a and b;
    layer1_outputs(2102) <= b;
    layer1_outputs(2103) <= not a or b;
    layer1_outputs(2104) <= a xor b;
    layer1_outputs(2105) <= a;
    layer1_outputs(2106) <= a or b;
    layer1_outputs(2107) <= a and not b;
    layer1_outputs(2108) <= not (a xor b);
    layer1_outputs(2109) <= 1'b1;
    layer1_outputs(2110) <= a;
    layer1_outputs(2111) <= not (a and b);
    layer1_outputs(2112) <= not a;
    layer1_outputs(2113) <= not (a xor b);
    layer1_outputs(2114) <= not b;
    layer1_outputs(2115) <= not b;
    layer1_outputs(2116) <= b;
    layer1_outputs(2117) <= not a;
    layer1_outputs(2118) <= 1'b0;
    layer1_outputs(2119) <= b;
    layer1_outputs(2120) <= not b or a;
    layer1_outputs(2121) <= not b or a;
    layer1_outputs(2122) <= a and b;
    layer1_outputs(2123) <= b;
    layer1_outputs(2124) <= not (a or b);
    layer1_outputs(2125) <= not (a xor b);
    layer1_outputs(2126) <= a;
    layer1_outputs(2127) <= a and not b;
    layer1_outputs(2128) <= not a;
    layer1_outputs(2129) <= a;
    layer1_outputs(2130) <= a and not b;
    layer1_outputs(2131) <= a or b;
    layer1_outputs(2132) <= a and b;
    layer1_outputs(2133) <= a;
    layer1_outputs(2134) <= not (a xor b);
    layer1_outputs(2135) <= not a or b;
    layer1_outputs(2136) <= a;
    layer1_outputs(2137) <= a;
    layer1_outputs(2138) <= 1'b1;
    layer1_outputs(2139) <= a xor b;
    layer1_outputs(2140) <= not b;
    layer1_outputs(2141) <= a;
    layer1_outputs(2142) <= not b;
    layer1_outputs(2143) <= a and not b;
    layer1_outputs(2144) <= a or b;
    layer1_outputs(2145) <= b and not a;
    layer1_outputs(2146) <= a xor b;
    layer1_outputs(2147) <= not a or b;
    layer1_outputs(2148) <= not (a and b);
    layer1_outputs(2149) <= 1'b0;
    layer1_outputs(2150) <= 1'b1;
    layer1_outputs(2151) <= not b;
    layer1_outputs(2152) <= b;
    layer1_outputs(2153) <= a or b;
    layer1_outputs(2154) <= b;
    layer1_outputs(2155) <= a;
    layer1_outputs(2156) <= not b;
    layer1_outputs(2157) <= a;
    layer1_outputs(2158) <= 1'b1;
    layer1_outputs(2159) <= not b;
    layer1_outputs(2160) <= a or b;
    layer1_outputs(2161) <= a and not b;
    layer1_outputs(2162) <= not a;
    layer1_outputs(2163) <= a and not b;
    layer1_outputs(2164) <= not a or b;
    layer1_outputs(2165) <= not a;
    layer1_outputs(2166) <= a and not b;
    layer1_outputs(2167) <= not (a and b);
    layer1_outputs(2168) <= a and b;
    layer1_outputs(2169) <= a xor b;
    layer1_outputs(2170) <= a xor b;
    layer1_outputs(2171) <= not (a xor b);
    layer1_outputs(2172) <= a;
    layer1_outputs(2173) <= 1'b1;
    layer1_outputs(2174) <= a and b;
    layer1_outputs(2175) <= a xor b;
    layer1_outputs(2176) <= b;
    layer1_outputs(2177) <= not (a xor b);
    layer1_outputs(2178) <= a and not b;
    layer1_outputs(2179) <= a;
    layer1_outputs(2180) <= not a;
    layer1_outputs(2181) <= a and not b;
    layer1_outputs(2182) <= b;
    layer1_outputs(2183) <= not b or a;
    layer1_outputs(2184) <= not a;
    layer1_outputs(2185) <= not (a or b);
    layer1_outputs(2186) <= not (a xor b);
    layer1_outputs(2187) <= not (a or b);
    layer1_outputs(2188) <= not b or a;
    layer1_outputs(2189) <= b;
    layer1_outputs(2190) <= a and not b;
    layer1_outputs(2191) <= a or b;
    layer1_outputs(2192) <= a;
    layer1_outputs(2193) <= a and not b;
    layer1_outputs(2194) <= not (a and b);
    layer1_outputs(2195) <= not b;
    layer1_outputs(2196) <= b;
    layer1_outputs(2197) <= a xor b;
    layer1_outputs(2198) <= not b or a;
    layer1_outputs(2199) <= 1'b1;
    layer1_outputs(2200) <= a;
    layer1_outputs(2201) <= a and not b;
    layer1_outputs(2202) <= not (a and b);
    layer1_outputs(2203) <= b and not a;
    layer1_outputs(2204) <= not a;
    layer1_outputs(2205) <= not b;
    layer1_outputs(2206) <= not b;
    layer1_outputs(2207) <= b;
    layer1_outputs(2208) <= not a;
    layer1_outputs(2209) <= a and not b;
    layer1_outputs(2210) <= not (a xor b);
    layer1_outputs(2211) <= not a;
    layer1_outputs(2212) <= a;
    layer1_outputs(2213) <= a and b;
    layer1_outputs(2214) <= a and not b;
    layer1_outputs(2215) <= not b or a;
    layer1_outputs(2216) <= b and not a;
    layer1_outputs(2217) <= not a;
    layer1_outputs(2218) <= not b;
    layer1_outputs(2219) <= b and not a;
    layer1_outputs(2220) <= a and not b;
    layer1_outputs(2221) <= a xor b;
    layer1_outputs(2222) <= a;
    layer1_outputs(2223) <= 1'b1;
    layer1_outputs(2224) <= b;
    layer1_outputs(2225) <= a or b;
    layer1_outputs(2226) <= a and not b;
    layer1_outputs(2227) <= b and not a;
    layer1_outputs(2228) <= not b or a;
    layer1_outputs(2229) <= not b;
    layer1_outputs(2230) <= a and not b;
    layer1_outputs(2231) <= a;
    layer1_outputs(2232) <= a;
    layer1_outputs(2233) <= a and b;
    layer1_outputs(2234) <= a and b;
    layer1_outputs(2235) <= b;
    layer1_outputs(2236) <= a and not b;
    layer1_outputs(2237) <= b;
    layer1_outputs(2238) <= a and not b;
    layer1_outputs(2239) <= not b or a;
    layer1_outputs(2240) <= a;
    layer1_outputs(2241) <= a xor b;
    layer1_outputs(2242) <= b;
    layer1_outputs(2243) <= not (a and b);
    layer1_outputs(2244) <= b;
    layer1_outputs(2245) <= a or b;
    layer1_outputs(2246) <= b and not a;
    layer1_outputs(2247) <= not a;
    layer1_outputs(2248) <= a;
    layer1_outputs(2249) <= a and b;
    layer1_outputs(2250) <= not b;
    layer1_outputs(2251) <= not (a or b);
    layer1_outputs(2252) <= not b or a;
    layer1_outputs(2253) <= a and not b;
    layer1_outputs(2254) <= not (a and b);
    layer1_outputs(2255) <= not a or b;
    layer1_outputs(2256) <= a and b;
    layer1_outputs(2257) <= b;
    layer1_outputs(2258) <= a and not b;
    layer1_outputs(2259) <= not (a or b);
    layer1_outputs(2260) <= not (a and b);
    layer1_outputs(2261) <= b;
    layer1_outputs(2262) <= not (a xor b);
    layer1_outputs(2263) <= not b;
    layer1_outputs(2264) <= a xor b;
    layer1_outputs(2265) <= not b;
    layer1_outputs(2266) <= 1'b0;
    layer1_outputs(2267) <= a xor b;
    layer1_outputs(2268) <= not b or a;
    layer1_outputs(2269) <= a and b;
    layer1_outputs(2270) <= b and not a;
    layer1_outputs(2271) <= not (a and b);
    layer1_outputs(2272) <= 1'b1;
    layer1_outputs(2273) <= b and not a;
    layer1_outputs(2274) <= a and not b;
    layer1_outputs(2275) <= not (a xor b);
    layer1_outputs(2276) <= not b;
    layer1_outputs(2277) <= not (a and b);
    layer1_outputs(2278) <= not b;
    layer1_outputs(2279) <= not (a xor b);
    layer1_outputs(2280) <= not (a xor b);
    layer1_outputs(2281) <= not (a and b);
    layer1_outputs(2282) <= not b or a;
    layer1_outputs(2283) <= not b;
    layer1_outputs(2284) <= a;
    layer1_outputs(2285) <= a xor b;
    layer1_outputs(2286) <= b;
    layer1_outputs(2287) <= not b;
    layer1_outputs(2288) <= not a or b;
    layer1_outputs(2289) <= not b;
    layer1_outputs(2290) <= a;
    layer1_outputs(2291) <= not b;
    layer1_outputs(2292) <= a and b;
    layer1_outputs(2293) <= not a or b;
    layer1_outputs(2294) <= b;
    layer1_outputs(2295) <= not (a and b);
    layer1_outputs(2296) <= not (a or b);
    layer1_outputs(2297) <= a and b;
    layer1_outputs(2298) <= not a or b;
    layer1_outputs(2299) <= not a;
    layer1_outputs(2300) <= b;
    layer1_outputs(2301) <= 1'b0;
    layer1_outputs(2302) <= a;
    layer1_outputs(2303) <= b;
    layer1_outputs(2304) <= not b or a;
    layer1_outputs(2305) <= not a or b;
    layer1_outputs(2306) <= b and not a;
    layer1_outputs(2307) <= 1'b1;
    layer1_outputs(2308) <= not a or b;
    layer1_outputs(2309) <= b;
    layer1_outputs(2310) <= a or b;
    layer1_outputs(2311) <= a and not b;
    layer1_outputs(2312) <= not a or b;
    layer1_outputs(2313) <= not a or b;
    layer1_outputs(2314) <= a and not b;
    layer1_outputs(2315) <= not a;
    layer1_outputs(2316) <= a and b;
    layer1_outputs(2317) <= a or b;
    layer1_outputs(2318) <= a or b;
    layer1_outputs(2319) <= 1'b0;
    layer1_outputs(2320) <= a and not b;
    layer1_outputs(2321) <= b and not a;
    layer1_outputs(2322) <= not (a or b);
    layer1_outputs(2323) <= not b;
    layer1_outputs(2324) <= a;
    layer1_outputs(2325) <= b;
    layer1_outputs(2326) <= a or b;
    layer1_outputs(2327) <= not b;
    layer1_outputs(2328) <= 1'b1;
    layer1_outputs(2329) <= b;
    layer1_outputs(2330) <= a;
    layer1_outputs(2331) <= a;
    layer1_outputs(2332) <= not (a xor b);
    layer1_outputs(2333) <= not (a or b);
    layer1_outputs(2334) <= not a or b;
    layer1_outputs(2335) <= not (a and b);
    layer1_outputs(2336) <= not (a xor b);
    layer1_outputs(2337) <= a;
    layer1_outputs(2338) <= not b or a;
    layer1_outputs(2339) <= not b;
    layer1_outputs(2340) <= not a;
    layer1_outputs(2341) <= a or b;
    layer1_outputs(2342) <= a xor b;
    layer1_outputs(2343) <= a and b;
    layer1_outputs(2344) <= not a or b;
    layer1_outputs(2345) <= a or b;
    layer1_outputs(2346) <= b;
    layer1_outputs(2347) <= not b;
    layer1_outputs(2348) <= a;
    layer1_outputs(2349) <= b and not a;
    layer1_outputs(2350) <= 1'b0;
    layer1_outputs(2351) <= 1'b1;
    layer1_outputs(2352) <= a;
    layer1_outputs(2353) <= not b;
    layer1_outputs(2354) <= a or b;
    layer1_outputs(2355) <= not b or a;
    layer1_outputs(2356) <= not (a or b);
    layer1_outputs(2357) <= not a or b;
    layer1_outputs(2358) <= b and not a;
    layer1_outputs(2359) <= not b or a;
    layer1_outputs(2360) <= a and not b;
    layer1_outputs(2361) <= a and not b;
    layer1_outputs(2362) <= a and b;
    layer1_outputs(2363) <= a and not b;
    layer1_outputs(2364) <= a and not b;
    layer1_outputs(2365) <= a and not b;
    layer1_outputs(2366) <= b;
    layer1_outputs(2367) <= a;
    layer1_outputs(2368) <= a and not b;
    layer1_outputs(2369) <= 1'b0;
    layer1_outputs(2370) <= 1'b1;
    layer1_outputs(2371) <= a;
    layer1_outputs(2372) <= not b or a;
    layer1_outputs(2373) <= not a;
    layer1_outputs(2374) <= a xor b;
    layer1_outputs(2375) <= b and not a;
    layer1_outputs(2376) <= not (a and b);
    layer1_outputs(2377) <= not (a and b);
    layer1_outputs(2378) <= not a;
    layer1_outputs(2379) <= not b;
    layer1_outputs(2380) <= a and not b;
    layer1_outputs(2381) <= a;
    layer1_outputs(2382) <= 1'b0;
    layer1_outputs(2383) <= not a;
    layer1_outputs(2384) <= not a or b;
    layer1_outputs(2385) <= a;
    layer1_outputs(2386) <= not b or a;
    layer1_outputs(2387) <= not b or a;
    layer1_outputs(2388) <= not a or b;
    layer1_outputs(2389) <= not (a or b);
    layer1_outputs(2390) <= not b;
    layer1_outputs(2391) <= b and not a;
    layer1_outputs(2392) <= a;
    layer1_outputs(2393) <= not (a xor b);
    layer1_outputs(2394) <= a and b;
    layer1_outputs(2395) <= not (a or b);
    layer1_outputs(2396) <= a xor b;
    layer1_outputs(2397) <= 1'b1;
    layer1_outputs(2398) <= not (a or b);
    layer1_outputs(2399) <= not (a or b);
    layer1_outputs(2400) <= not (a xor b);
    layer1_outputs(2401) <= not (a and b);
    layer1_outputs(2402) <= a xor b;
    layer1_outputs(2403) <= not a;
    layer1_outputs(2404) <= not b;
    layer1_outputs(2405) <= a and b;
    layer1_outputs(2406) <= b and not a;
    layer1_outputs(2407) <= 1'b1;
    layer1_outputs(2408) <= not b or a;
    layer1_outputs(2409) <= a;
    layer1_outputs(2410) <= 1'b1;
    layer1_outputs(2411) <= b and not a;
    layer1_outputs(2412) <= not a or b;
    layer1_outputs(2413) <= a;
    layer1_outputs(2414) <= a or b;
    layer1_outputs(2415) <= not (a xor b);
    layer1_outputs(2416) <= not b;
    layer1_outputs(2417) <= not (a or b);
    layer1_outputs(2418) <= a and b;
    layer1_outputs(2419) <= a and not b;
    layer1_outputs(2420) <= 1'b0;
    layer1_outputs(2421) <= a or b;
    layer1_outputs(2422) <= a or b;
    layer1_outputs(2423) <= a and not b;
    layer1_outputs(2424) <= a;
    layer1_outputs(2425) <= not (a and b);
    layer1_outputs(2426) <= not (a and b);
    layer1_outputs(2427) <= a;
    layer1_outputs(2428) <= not a or b;
    layer1_outputs(2429) <= a and not b;
    layer1_outputs(2430) <= not b;
    layer1_outputs(2431) <= a xor b;
    layer1_outputs(2432) <= a xor b;
    layer1_outputs(2433) <= not b or a;
    layer1_outputs(2434) <= b;
    layer1_outputs(2435) <= 1'b1;
    layer1_outputs(2436) <= 1'b0;
    layer1_outputs(2437) <= a and b;
    layer1_outputs(2438) <= not b;
    layer1_outputs(2439) <= not (a and b);
    layer1_outputs(2440) <= not a or b;
    layer1_outputs(2441) <= not (a xor b);
    layer1_outputs(2442) <= not a or b;
    layer1_outputs(2443) <= b and not a;
    layer1_outputs(2444) <= not b;
    layer1_outputs(2445) <= not b;
    layer1_outputs(2446) <= a and b;
    layer1_outputs(2447) <= not b;
    layer1_outputs(2448) <= b;
    layer1_outputs(2449) <= b;
    layer1_outputs(2450) <= not b or a;
    layer1_outputs(2451) <= not b or a;
    layer1_outputs(2452) <= a and not b;
    layer1_outputs(2453) <= not (a or b);
    layer1_outputs(2454) <= not (a xor b);
    layer1_outputs(2455) <= not (a or b);
    layer1_outputs(2456) <= a;
    layer1_outputs(2457) <= a and b;
    layer1_outputs(2458) <= 1'b0;
    layer1_outputs(2459) <= not b;
    layer1_outputs(2460) <= not b;
    layer1_outputs(2461) <= b;
    layer1_outputs(2462) <= a or b;
    layer1_outputs(2463) <= not b;
    layer1_outputs(2464) <= a and not b;
    layer1_outputs(2465) <= a;
    layer1_outputs(2466) <= a;
    layer1_outputs(2467) <= a;
    layer1_outputs(2468) <= a xor b;
    layer1_outputs(2469) <= a and not b;
    layer1_outputs(2470) <= 1'b1;
    layer1_outputs(2471) <= not b;
    layer1_outputs(2472) <= not b or a;
    layer1_outputs(2473) <= not b or a;
    layer1_outputs(2474) <= not a;
    layer1_outputs(2475) <= not b or a;
    layer1_outputs(2476) <= b;
    layer1_outputs(2477) <= not a;
    layer1_outputs(2478) <= not (a and b);
    layer1_outputs(2479) <= not b;
    layer1_outputs(2480) <= a;
    layer1_outputs(2481) <= b and not a;
    layer1_outputs(2482) <= b and not a;
    layer1_outputs(2483) <= b and not a;
    layer1_outputs(2484) <= a;
    layer1_outputs(2485) <= not b;
    layer1_outputs(2486) <= not a;
    layer1_outputs(2487) <= b;
    layer1_outputs(2488) <= a and not b;
    layer1_outputs(2489) <= a xor b;
    layer1_outputs(2490) <= a and b;
    layer1_outputs(2491) <= not b;
    layer1_outputs(2492) <= not b;
    layer1_outputs(2493) <= not a or b;
    layer1_outputs(2494) <= 1'b1;
    layer1_outputs(2495) <= b and not a;
    layer1_outputs(2496) <= not b;
    layer1_outputs(2497) <= a;
    layer1_outputs(2498) <= a;
    layer1_outputs(2499) <= b and not a;
    layer1_outputs(2500) <= a and not b;
    layer1_outputs(2501) <= a and b;
    layer1_outputs(2502) <= 1'b1;
    layer1_outputs(2503) <= a and not b;
    layer1_outputs(2504) <= a;
    layer1_outputs(2505) <= a xor b;
    layer1_outputs(2506) <= a and b;
    layer1_outputs(2507) <= not a or b;
    layer1_outputs(2508) <= not (a xor b);
    layer1_outputs(2509) <= b and not a;
    layer1_outputs(2510) <= not a or b;
    layer1_outputs(2511) <= not a or b;
    layer1_outputs(2512) <= not b or a;
    layer1_outputs(2513) <= a and not b;
    layer1_outputs(2514) <= not b;
    layer1_outputs(2515) <= not (a or b);
    layer1_outputs(2516) <= a or b;
    layer1_outputs(2517) <= b;
    layer1_outputs(2518) <= b and not a;
    layer1_outputs(2519) <= a and not b;
    layer1_outputs(2520) <= b and not a;
    layer1_outputs(2521) <= a xor b;
    layer1_outputs(2522) <= a and b;
    layer1_outputs(2523) <= not a;
    layer1_outputs(2524) <= 1'b1;
    layer1_outputs(2525) <= b and not a;
    layer1_outputs(2526) <= a or b;
    layer1_outputs(2527) <= 1'b1;
    layer1_outputs(2528) <= not a or b;
    layer1_outputs(2529) <= b;
    layer1_outputs(2530) <= b;
    layer1_outputs(2531) <= a xor b;
    layer1_outputs(2532) <= a and b;
    layer1_outputs(2533) <= not (a or b);
    layer1_outputs(2534) <= not b or a;
    layer1_outputs(2535) <= not a;
    layer1_outputs(2536) <= not a;
    layer1_outputs(2537) <= a;
    layer1_outputs(2538) <= a and not b;
    layer1_outputs(2539) <= not (a and b);
    layer1_outputs(2540) <= not (a and b);
    layer1_outputs(2541) <= a and b;
    layer1_outputs(2542) <= not (a or b);
    layer1_outputs(2543) <= a and b;
    layer1_outputs(2544) <= a or b;
    layer1_outputs(2545) <= not (a or b);
    layer1_outputs(2546) <= a;
    layer1_outputs(2547) <= b and not a;
    layer1_outputs(2548) <= not a;
    layer1_outputs(2549) <= a or b;
    layer1_outputs(2550) <= a;
    layer1_outputs(2551) <= a;
    layer1_outputs(2552) <= a and b;
    layer1_outputs(2553) <= a and b;
    layer1_outputs(2554) <= not (a and b);
    layer1_outputs(2555) <= b;
    layer1_outputs(2556) <= a or b;
    layer1_outputs(2557) <= not b or a;
    layer1_outputs(2558) <= a and not b;
    layer1_outputs(2559) <= 1'b1;
    layer1_outputs(2560) <= a and b;
    layer1_outputs(2561) <= not (a and b);
    layer1_outputs(2562) <= a or b;
    layer1_outputs(2563) <= a;
    layer1_outputs(2564) <= not b;
    layer1_outputs(2565) <= a;
    layer1_outputs(2566) <= not (a and b);
    layer1_outputs(2567) <= b;
    layer1_outputs(2568) <= a or b;
    layer1_outputs(2569) <= not (a xor b);
    layer1_outputs(2570) <= b;
    layer1_outputs(2571) <= b;
    layer1_outputs(2572) <= a xor b;
    layer1_outputs(2573) <= not (a xor b);
    layer1_outputs(2574) <= a xor b;
    layer1_outputs(2575) <= not (a xor b);
    layer1_outputs(2576) <= not b;
    layer1_outputs(2577) <= b;
    layer1_outputs(2578) <= not b;
    layer1_outputs(2579) <= a or b;
    layer1_outputs(2580) <= a and b;
    layer1_outputs(2581) <= a and b;
    layer1_outputs(2582) <= not b;
    layer1_outputs(2583) <= not (a or b);
    layer1_outputs(2584) <= 1'b0;
    layer1_outputs(2585) <= 1'b1;
    layer1_outputs(2586) <= b and not a;
    layer1_outputs(2587) <= 1'b0;
    layer1_outputs(2588) <= not (a and b);
    layer1_outputs(2589) <= not a;
    layer1_outputs(2590) <= a;
    layer1_outputs(2591) <= a and b;
    layer1_outputs(2592) <= not a or b;
    layer1_outputs(2593) <= b;
    layer1_outputs(2594) <= a xor b;
    layer1_outputs(2595) <= a or b;
    layer1_outputs(2596) <= a;
    layer1_outputs(2597) <= not a;
    layer1_outputs(2598) <= a;
    layer1_outputs(2599) <= not (a or b);
    layer1_outputs(2600) <= a or b;
    layer1_outputs(2601) <= a;
    layer1_outputs(2602) <= a or b;
    layer1_outputs(2603) <= a;
    layer1_outputs(2604) <= not b;
    layer1_outputs(2605) <= b;
    layer1_outputs(2606) <= not (a xor b);
    layer1_outputs(2607) <= a or b;
    layer1_outputs(2608) <= b;
    layer1_outputs(2609) <= b;
    layer1_outputs(2610) <= not (a or b);
    layer1_outputs(2611) <= a and b;
    layer1_outputs(2612) <= not (a or b);
    layer1_outputs(2613) <= not b;
    layer1_outputs(2614) <= b;
    layer1_outputs(2615) <= a or b;
    layer1_outputs(2616) <= not a;
    layer1_outputs(2617) <= not b or a;
    layer1_outputs(2618) <= a xor b;
    layer1_outputs(2619) <= not b;
    layer1_outputs(2620) <= not (a and b);
    layer1_outputs(2621) <= a and b;
    layer1_outputs(2622) <= not a;
    layer1_outputs(2623) <= 1'b0;
    layer1_outputs(2624) <= not b or a;
    layer1_outputs(2625) <= not b;
    layer1_outputs(2626) <= not b or a;
    layer1_outputs(2627) <= a;
    layer1_outputs(2628) <= a and not b;
    layer1_outputs(2629) <= b and not a;
    layer1_outputs(2630) <= not b;
    layer1_outputs(2631) <= 1'b0;
    layer1_outputs(2632) <= b;
    layer1_outputs(2633) <= not (a or b);
    layer1_outputs(2634) <= a;
    layer1_outputs(2635) <= 1'b0;
    layer1_outputs(2636) <= not (a xor b);
    layer1_outputs(2637) <= 1'b1;
    layer1_outputs(2638) <= not b or a;
    layer1_outputs(2639) <= not a or b;
    layer1_outputs(2640) <= not (a xor b);
    layer1_outputs(2641) <= not (a xor b);
    layer1_outputs(2642) <= a and b;
    layer1_outputs(2643) <= b and not a;
    layer1_outputs(2644) <= 1'b1;
    layer1_outputs(2645) <= b and not a;
    layer1_outputs(2646) <= not a;
    layer1_outputs(2647) <= a or b;
    layer1_outputs(2648) <= a;
    layer1_outputs(2649) <= 1'b1;
    layer1_outputs(2650) <= not a;
    layer1_outputs(2651) <= not (a and b);
    layer1_outputs(2652) <= b;
    layer1_outputs(2653) <= a and b;
    layer1_outputs(2654) <= not b or a;
    layer1_outputs(2655) <= a and not b;
    layer1_outputs(2656) <= not a;
    layer1_outputs(2657) <= a or b;
    layer1_outputs(2658) <= a and not b;
    layer1_outputs(2659) <= a and b;
    layer1_outputs(2660) <= not b or a;
    layer1_outputs(2661) <= b and not a;
    layer1_outputs(2662) <= a or b;
    layer1_outputs(2663) <= not (a and b);
    layer1_outputs(2664) <= a or b;
    layer1_outputs(2665) <= not a or b;
    layer1_outputs(2666) <= not a or b;
    layer1_outputs(2667) <= b and not a;
    layer1_outputs(2668) <= not b;
    layer1_outputs(2669) <= not (a or b);
    layer1_outputs(2670) <= b and not a;
    layer1_outputs(2671) <= a xor b;
    layer1_outputs(2672) <= a;
    layer1_outputs(2673) <= a and b;
    layer1_outputs(2674) <= 1'b0;
    layer1_outputs(2675) <= b and not a;
    layer1_outputs(2676) <= b;
    layer1_outputs(2677) <= not b;
    layer1_outputs(2678) <= b and not a;
    layer1_outputs(2679) <= not a;
    layer1_outputs(2680) <= not b;
    layer1_outputs(2681) <= b;
    layer1_outputs(2682) <= not (a xor b);
    layer1_outputs(2683) <= not (a or b);
    layer1_outputs(2684) <= b;
    layer1_outputs(2685) <= not a;
    layer1_outputs(2686) <= a;
    layer1_outputs(2687) <= not b;
    layer1_outputs(2688) <= a;
    layer1_outputs(2689) <= not (a xor b);
    layer1_outputs(2690) <= not a;
    layer1_outputs(2691) <= a;
    layer1_outputs(2692) <= 1'b0;
    layer1_outputs(2693) <= not (a and b);
    layer1_outputs(2694) <= b;
    layer1_outputs(2695) <= not (a and b);
    layer1_outputs(2696) <= not b;
    layer1_outputs(2697) <= a and b;
    layer1_outputs(2698) <= not a or b;
    layer1_outputs(2699) <= a and b;
    layer1_outputs(2700) <= a;
    layer1_outputs(2701) <= 1'b1;
    layer1_outputs(2702) <= not b;
    layer1_outputs(2703) <= a xor b;
    layer1_outputs(2704) <= a;
    layer1_outputs(2705) <= 1'b0;
    layer1_outputs(2706) <= a xor b;
    layer1_outputs(2707) <= not b or a;
    layer1_outputs(2708) <= a or b;
    layer1_outputs(2709) <= a and b;
    layer1_outputs(2710) <= 1'b0;
    layer1_outputs(2711) <= a or b;
    layer1_outputs(2712) <= not a or b;
    layer1_outputs(2713) <= a;
    layer1_outputs(2714) <= a or b;
    layer1_outputs(2715) <= not a;
    layer1_outputs(2716) <= not a;
    layer1_outputs(2717) <= not b or a;
    layer1_outputs(2718) <= not a;
    layer1_outputs(2719) <= not a or b;
    layer1_outputs(2720) <= not b;
    layer1_outputs(2721) <= 1'b0;
    layer1_outputs(2722) <= not (a or b);
    layer1_outputs(2723) <= 1'b1;
    layer1_outputs(2724) <= b;
    layer1_outputs(2725) <= not (a or b);
    layer1_outputs(2726) <= b and not a;
    layer1_outputs(2727) <= a;
    layer1_outputs(2728) <= not a;
    layer1_outputs(2729) <= a or b;
    layer1_outputs(2730) <= 1'b0;
    layer1_outputs(2731) <= 1'b1;
    layer1_outputs(2732) <= a xor b;
    layer1_outputs(2733) <= a;
    layer1_outputs(2734) <= not a;
    layer1_outputs(2735) <= not (a or b);
    layer1_outputs(2736) <= 1'b1;
    layer1_outputs(2737) <= a;
    layer1_outputs(2738) <= 1'b1;
    layer1_outputs(2739) <= not (a xor b);
    layer1_outputs(2740) <= b and not a;
    layer1_outputs(2741) <= not a or b;
    layer1_outputs(2742) <= b and not a;
    layer1_outputs(2743) <= not a or b;
    layer1_outputs(2744) <= not b;
    layer1_outputs(2745) <= a;
    layer1_outputs(2746) <= not (a and b);
    layer1_outputs(2747) <= 1'b1;
    layer1_outputs(2748) <= a or b;
    layer1_outputs(2749) <= not (a or b);
    layer1_outputs(2750) <= not b;
    layer1_outputs(2751) <= not (a xor b);
    layer1_outputs(2752) <= not b or a;
    layer1_outputs(2753) <= a and not b;
    layer1_outputs(2754) <= 1'b0;
    layer1_outputs(2755) <= not a;
    layer1_outputs(2756) <= not (a or b);
    layer1_outputs(2757) <= 1'b1;
    layer1_outputs(2758) <= a xor b;
    layer1_outputs(2759) <= b;
    layer1_outputs(2760) <= not (a or b);
    layer1_outputs(2761) <= a and not b;
    layer1_outputs(2762) <= not a;
    layer1_outputs(2763) <= a and not b;
    layer1_outputs(2764) <= not a or b;
    layer1_outputs(2765) <= not (a and b);
    layer1_outputs(2766) <= not (a and b);
    layer1_outputs(2767) <= b and not a;
    layer1_outputs(2768) <= a and not b;
    layer1_outputs(2769) <= a and not b;
    layer1_outputs(2770) <= not b;
    layer1_outputs(2771) <= not (a and b);
    layer1_outputs(2772) <= not a or b;
    layer1_outputs(2773) <= a and not b;
    layer1_outputs(2774) <= not b or a;
    layer1_outputs(2775) <= a;
    layer1_outputs(2776) <= not b or a;
    layer1_outputs(2777) <= a and not b;
    layer1_outputs(2778) <= b;
    layer1_outputs(2779) <= a and b;
    layer1_outputs(2780) <= not b or a;
    layer1_outputs(2781) <= not b or a;
    layer1_outputs(2782) <= a;
    layer1_outputs(2783) <= not b or a;
    layer1_outputs(2784) <= a and b;
    layer1_outputs(2785) <= a or b;
    layer1_outputs(2786) <= b;
    layer1_outputs(2787) <= not a;
    layer1_outputs(2788) <= a;
    layer1_outputs(2789) <= not a or b;
    layer1_outputs(2790) <= not (a xor b);
    layer1_outputs(2791) <= b;
    layer1_outputs(2792) <= not b;
    layer1_outputs(2793) <= not a or b;
    layer1_outputs(2794) <= not b;
    layer1_outputs(2795) <= not (a or b);
    layer1_outputs(2796) <= not a;
    layer1_outputs(2797) <= not (a and b);
    layer1_outputs(2798) <= b and not a;
    layer1_outputs(2799) <= not b or a;
    layer1_outputs(2800) <= not (a or b);
    layer1_outputs(2801) <= not b;
    layer1_outputs(2802) <= not (a and b);
    layer1_outputs(2803) <= 1'b1;
    layer1_outputs(2804) <= b and not a;
    layer1_outputs(2805) <= not (a or b);
    layer1_outputs(2806) <= a and not b;
    layer1_outputs(2807) <= not a;
    layer1_outputs(2808) <= a xor b;
    layer1_outputs(2809) <= not b or a;
    layer1_outputs(2810) <= not (a and b);
    layer1_outputs(2811) <= not (a or b);
    layer1_outputs(2812) <= a or b;
    layer1_outputs(2813) <= b and not a;
    layer1_outputs(2814) <= a and b;
    layer1_outputs(2815) <= not (a or b);
    layer1_outputs(2816) <= not b;
    layer1_outputs(2817) <= 1'b1;
    layer1_outputs(2818) <= not b;
    layer1_outputs(2819) <= not a;
    layer1_outputs(2820) <= a or b;
    layer1_outputs(2821) <= b and not a;
    layer1_outputs(2822) <= not b;
    layer1_outputs(2823) <= not a or b;
    layer1_outputs(2824) <= a;
    layer1_outputs(2825) <= 1'b0;
    layer1_outputs(2826) <= b;
    layer1_outputs(2827) <= a;
    layer1_outputs(2828) <= not (a xor b);
    layer1_outputs(2829) <= not a;
    layer1_outputs(2830) <= a and b;
    layer1_outputs(2831) <= not b;
    layer1_outputs(2832) <= a;
    layer1_outputs(2833) <= not a or b;
    layer1_outputs(2834) <= 1'b0;
    layer1_outputs(2835) <= not (a or b);
    layer1_outputs(2836) <= 1'b1;
    layer1_outputs(2837) <= b and not a;
    layer1_outputs(2838) <= not b or a;
    layer1_outputs(2839) <= not (a or b);
    layer1_outputs(2840) <= a and not b;
    layer1_outputs(2841) <= 1'b0;
    layer1_outputs(2842) <= a;
    layer1_outputs(2843) <= not b;
    layer1_outputs(2844) <= 1'b1;
    layer1_outputs(2845) <= not b or a;
    layer1_outputs(2846) <= a or b;
    layer1_outputs(2847) <= not (a or b);
    layer1_outputs(2848) <= not a;
    layer1_outputs(2849) <= not b;
    layer1_outputs(2850) <= not b or a;
    layer1_outputs(2851) <= not (a or b);
    layer1_outputs(2852) <= a and b;
    layer1_outputs(2853) <= not (a or b);
    layer1_outputs(2854) <= a;
    layer1_outputs(2855) <= not (a and b);
    layer1_outputs(2856) <= a xor b;
    layer1_outputs(2857) <= a and not b;
    layer1_outputs(2858) <= not (a and b);
    layer1_outputs(2859) <= a;
    layer1_outputs(2860) <= b and not a;
    layer1_outputs(2861) <= b;
    layer1_outputs(2862) <= not b or a;
    layer1_outputs(2863) <= not (a xor b);
    layer1_outputs(2864) <= not (a xor b);
    layer1_outputs(2865) <= not (a and b);
    layer1_outputs(2866) <= not a;
    layer1_outputs(2867) <= a and not b;
    layer1_outputs(2868) <= a xor b;
    layer1_outputs(2869) <= a xor b;
    layer1_outputs(2870) <= b;
    layer1_outputs(2871) <= not (a and b);
    layer1_outputs(2872) <= not (a or b);
    layer1_outputs(2873) <= not a or b;
    layer1_outputs(2874) <= a xor b;
    layer1_outputs(2875) <= not a;
    layer1_outputs(2876) <= not (a and b);
    layer1_outputs(2877) <= a xor b;
    layer1_outputs(2878) <= a;
    layer1_outputs(2879) <= a and not b;
    layer1_outputs(2880) <= b;
    layer1_outputs(2881) <= a;
    layer1_outputs(2882) <= not a;
    layer1_outputs(2883) <= b;
    layer1_outputs(2884) <= not (a or b);
    layer1_outputs(2885) <= a;
    layer1_outputs(2886) <= a or b;
    layer1_outputs(2887) <= not (a or b);
    layer1_outputs(2888) <= not (a or b);
    layer1_outputs(2889) <= not a;
    layer1_outputs(2890) <= b;
    layer1_outputs(2891) <= not (a and b);
    layer1_outputs(2892) <= not b or a;
    layer1_outputs(2893) <= b;
    layer1_outputs(2894) <= not (a and b);
    layer1_outputs(2895) <= not b;
    layer1_outputs(2896) <= a;
    layer1_outputs(2897) <= a xor b;
    layer1_outputs(2898) <= not (a or b);
    layer1_outputs(2899) <= a xor b;
    layer1_outputs(2900) <= not a or b;
    layer1_outputs(2901) <= a or b;
    layer1_outputs(2902) <= a;
    layer1_outputs(2903) <= not b or a;
    layer1_outputs(2904) <= b and not a;
    layer1_outputs(2905) <= not (a or b);
    layer1_outputs(2906) <= not b;
    layer1_outputs(2907) <= not (a xor b);
    layer1_outputs(2908) <= not b or a;
    layer1_outputs(2909) <= a xor b;
    layer1_outputs(2910) <= not b;
    layer1_outputs(2911) <= not (a xor b);
    layer1_outputs(2912) <= not a;
    layer1_outputs(2913) <= not b or a;
    layer1_outputs(2914) <= a or b;
    layer1_outputs(2915) <= a and b;
    layer1_outputs(2916) <= a xor b;
    layer1_outputs(2917) <= a;
    layer1_outputs(2918) <= not b;
    layer1_outputs(2919) <= not a;
    layer1_outputs(2920) <= a;
    layer1_outputs(2921) <= a or b;
    layer1_outputs(2922) <= a and not b;
    layer1_outputs(2923) <= not b or a;
    layer1_outputs(2924) <= 1'b1;
    layer1_outputs(2925) <= 1'b0;
    layer1_outputs(2926) <= a and not b;
    layer1_outputs(2927) <= b and not a;
    layer1_outputs(2928) <= not (a and b);
    layer1_outputs(2929) <= a xor b;
    layer1_outputs(2930) <= not b or a;
    layer1_outputs(2931) <= not b;
    layer1_outputs(2932) <= not a;
    layer1_outputs(2933) <= not (a xor b);
    layer1_outputs(2934) <= b and not a;
    layer1_outputs(2935) <= not a;
    layer1_outputs(2936) <= not a or b;
    layer1_outputs(2937) <= 1'b1;
    layer1_outputs(2938) <= a or b;
    layer1_outputs(2939) <= not (a and b);
    layer1_outputs(2940) <= not b or a;
    layer1_outputs(2941) <= not (a or b);
    layer1_outputs(2942) <= b and not a;
    layer1_outputs(2943) <= a;
    layer1_outputs(2944) <= not (a xor b);
    layer1_outputs(2945) <= not a;
    layer1_outputs(2946) <= not a or b;
    layer1_outputs(2947) <= not a;
    layer1_outputs(2948) <= not (a or b);
    layer1_outputs(2949) <= not a or b;
    layer1_outputs(2950) <= not a;
    layer1_outputs(2951) <= a and not b;
    layer1_outputs(2952) <= 1'b1;
    layer1_outputs(2953) <= a or b;
    layer1_outputs(2954) <= not a or b;
    layer1_outputs(2955) <= b;
    layer1_outputs(2956) <= not (a xor b);
    layer1_outputs(2957) <= not (a or b);
    layer1_outputs(2958) <= not (a xor b);
    layer1_outputs(2959) <= a;
    layer1_outputs(2960) <= a and not b;
    layer1_outputs(2961) <= a;
    layer1_outputs(2962) <= not a or b;
    layer1_outputs(2963) <= not a;
    layer1_outputs(2964) <= b;
    layer1_outputs(2965) <= a and b;
    layer1_outputs(2966) <= 1'b1;
    layer1_outputs(2967) <= b;
    layer1_outputs(2968) <= not a;
    layer1_outputs(2969) <= not a or b;
    layer1_outputs(2970) <= a;
    layer1_outputs(2971) <= a xor b;
    layer1_outputs(2972) <= a;
    layer1_outputs(2973) <= not (a xor b);
    layer1_outputs(2974) <= not b or a;
    layer1_outputs(2975) <= not (a and b);
    layer1_outputs(2976) <= not a or b;
    layer1_outputs(2977) <= not a or b;
    layer1_outputs(2978) <= not b;
    layer1_outputs(2979) <= a xor b;
    layer1_outputs(2980) <= b;
    layer1_outputs(2981) <= 1'b0;
    layer1_outputs(2982) <= b;
    layer1_outputs(2983) <= not (a or b);
    layer1_outputs(2984) <= a and not b;
    layer1_outputs(2985) <= not (a and b);
    layer1_outputs(2986) <= not a;
    layer1_outputs(2987) <= not a;
    layer1_outputs(2988) <= b;
    layer1_outputs(2989) <= not (a xor b);
    layer1_outputs(2990) <= a and not b;
    layer1_outputs(2991) <= a and b;
    layer1_outputs(2992) <= not a;
    layer1_outputs(2993) <= not (a and b);
    layer1_outputs(2994) <= a or b;
    layer1_outputs(2995) <= not a or b;
    layer1_outputs(2996) <= not (a and b);
    layer1_outputs(2997) <= b and not a;
    layer1_outputs(2998) <= a xor b;
    layer1_outputs(2999) <= a or b;
    layer1_outputs(3000) <= a;
    layer1_outputs(3001) <= 1'b1;
    layer1_outputs(3002) <= a and not b;
    layer1_outputs(3003) <= a or b;
    layer1_outputs(3004) <= a and not b;
    layer1_outputs(3005) <= a and not b;
    layer1_outputs(3006) <= b;
    layer1_outputs(3007) <= b;
    layer1_outputs(3008) <= b;
    layer1_outputs(3009) <= not (a or b);
    layer1_outputs(3010) <= not a;
    layer1_outputs(3011) <= not (a and b);
    layer1_outputs(3012) <= a and b;
    layer1_outputs(3013) <= b and not a;
    layer1_outputs(3014) <= a and not b;
    layer1_outputs(3015) <= not (a xor b);
    layer1_outputs(3016) <= b;
    layer1_outputs(3017) <= b;
    layer1_outputs(3018) <= not a;
    layer1_outputs(3019) <= a and not b;
    layer1_outputs(3020) <= a and not b;
    layer1_outputs(3021) <= 1'b0;
    layer1_outputs(3022) <= a and b;
    layer1_outputs(3023) <= b;
    layer1_outputs(3024) <= b;
    layer1_outputs(3025) <= not a;
    layer1_outputs(3026) <= not (a or b);
    layer1_outputs(3027) <= not a;
    layer1_outputs(3028) <= not b or a;
    layer1_outputs(3029) <= a or b;
    layer1_outputs(3030) <= a xor b;
    layer1_outputs(3031) <= not (a xor b);
    layer1_outputs(3032) <= b and not a;
    layer1_outputs(3033) <= a and not b;
    layer1_outputs(3034) <= not a;
    layer1_outputs(3035) <= a and not b;
    layer1_outputs(3036) <= a and not b;
    layer1_outputs(3037) <= not b or a;
    layer1_outputs(3038) <= a and b;
    layer1_outputs(3039) <= not (a and b);
    layer1_outputs(3040) <= not a or b;
    layer1_outputs(3041) <= not (a xor b);
    layer1_outputs(3042) <= not (a xor b);
    layer1_outputs(3043) <= b;
    layer1_outputs(3044) <= a and b;
    layer1_outputs(3045) <= b;
    layer1_outputs(3046) <= not a;
    layer1_outputs(3047) <= not (a or b);
    layer1_outputs(3048) <= not b;
    layer1_outputs(3049) <= b;
    layer1_outputs(3050) <= not a or b;
    layer1_outputs(3051) <= 1'b0;
    layer1_outputs(3052) <= b and not a;
    layer1_outputs(3053) <= not b or a;
    layer1_outputs(3054) <= not (a or b);
    layer1_outputs(3055) <= not (a xor b);
    layer1_outputs(3056) <= not b;
    layer1_outputs(3057) <= a and not b;
    layer1_outputs(3058) <= b and not a;
    layer1_outputs(3059) <= 1'b1;
    layer1_outputs(3060) <= not a or b;
    layer1_outputs(3061) <= not (a or b);
    layer1_outputs(3062) <= not b or a;
    layer1_outputs(3063) <= a or b;
    layer1_outputs(3064) <= a and b;
    layer1_outputs(3065) <= 1'b0;
    layer1_outputs(3066) <= not a or b;
    layer1_outputs(3067) <= a;
    layer1_outputs(3068) <= not a or b;
    layer1_outputs(3069) <= not b;
    layer1_outputs(3070) <= not (a and b);
    layer1_outputs(3071) <= a and b;
    layer1_outputs(3072) <= not a;
    layer1_outputs(3073) <= not a;
    layer1_outputs(3074) <= a and not b;
    layer1_outputs(3075) <= not (a and b);
    layer1_outputs(3076) <= not a or b;
    layer1_outputs(3077) <= not (a or b);
    layer1_outputs(3078) <= not (a and b);
    layer1_outputs(3079) <= b;
    layer1_outputs(3080) <= not a;
    layer1_outputs(3081) <= b and not a;
    layer1_outputs(3082) <= a and b;
    layer1_outputs(3083) <= 1'b1;
    layer1_outputs(3084) <= not a;
    layer1_outputs(3085) <= not a or b;
    layer1_outputs(3086) <= a and not b;
    layer1_outputs(3087) <= b and not a;
    layer1_outputs(3088) <= a;
    layer1_outputs(3089) <= a and not b;
    layer1_outputs(3090) <= a or b;
    layer1_outputs(3091) <= not a or b;
    layer1_outputs(3092) <= not b or a;
    layer1_outputs(3093) <= b;
    layer1_outputs(3094) <= b;
    layer1_outputs(3095) <= not b or a;
    layer1_outputs(3096) <= not a;
    layer1_outputs(3097) <= not (a and b);
    layer1_outputs(3098) <= a xor b;
    layer1_outputs(3099) <= not a;
    layer1_outputs(3100) <= a and not b;
    layer1_outputs(3101) <= not (a and b);
    layer1_outputs(3102) <= b and not a;
    layer1_outputs(3103) <= a and not b;
    layer1_outputs(3104) <= a or b;
    layer1_outputs(3105) <= not b or a;
    layer1_outputs(3106) <= not (a xor b);
    layer1_outputs(3107) <= not (a xor b);
    layer1_outputs(3108) <= a and b;
    layer1_outputs(3109) <= not (a and b);
    layer1_outputs(3110) <= b;
    layer1_outputs(3111) <= not a;
    layer1_outputs(3112) <= b and not a;
    layer1_outputs(3113) <= b and not a;
    layer1_outputs(3114) <= not (a and b);
    layer1_outputs(3115) <= b;
    layer1_outputs(3116) <= not b;
    layer1_outputs(3117) <= a xor b;
    layer1_outputs(3118) <= not (a and b);
    layer1_outputs(3119) <= not b or a;
    layer1_outputs(3120) <= b and not a;
    layer1_outputs(3121) <= a and b;
    layer1_outputs(3122) <= not a;
    layer1_outputs(3123) <= not (a or b);
    layer1_outputs(3124) <= not (a or b);
    layer1_outputs(3125) <= b;
    layer1_outputs(3126) <= a or b;
    layer1_outputs(3127) <= not (a or b);
    layer1_outputs(3128) <= b;
    layer1_outputs(3129) <= 1'b1;
    layer1_outputs(3130) <= not (a or b);
    layer1_outputs(3131) <= a and b;
    layer1_outputs(3132) <= not (a or b);
    layer1_outputs(3133) <= a or b;
    layer1_outputs(3134) <= not (a or b);
    layer1_outputs(3135) <= a;
    layer1_outputs(3136) <= not a;
    layer1_outputs(3137) <= a or b;
    layer1_outputs(3138) <= not a or b;
    layer1_outputs(3139) <= b and not a;
    layer1_outputs(3140) <= b;
    layer1_outputs(3141) <= not a or b;
    layer1_outputs(3142) <= not b;
    layer1_outputs(3143) <= not a or b;
    layer1_outputs(3144) <= not b;
    layer1_outputs(3145) <= not a or b;
    layer1_outputs(3146) <= not b;
    layer1_outputs(3147) <= not b or a;
    layer1_outputs(3148) <= not (a and b);
    layer1_outputs(3149) <= not a or b;
    layer1_outputs(3150) <= not b or a;
    layer1_outputs(3151) <= 1'b0;
    layer1_outputs(3152) <= not a;
    layer1_outputs(3153) <= a;
    layer1_outputs(3154) <= 1'b0;
    layer1_outputs(3155) <= not a or b;
    layer1_outputs(3156) <= a or b;
    layer1_outputs(3157) <= not b or a;
    layer1_outputs(3158) <= a xor b;
    layer1_outputs(3159) <= 1'b0;
    layer1_outputs(3160) <= not (a or b);
    layer1_outputs(3161) <= a or b;
    layer1_outputs(3162) <= 1'b0;
    layer1_outputs(3163) <= not b or a;
    layer1_outputs(3164) <= not (a and b);
    layer1_outputs(3165) <= not a;
    layer1_outputs(3166) <= a;
    layer1_outputs(3167) <= a and b;
    layer1_outputs(3168) <= not (a or b);
    layer1_outputs(3169) <= a and not b;
    layer1_outputs(3170) <= b and not a;
    layer1_outputs(3171) <= not (a and b);
    layer1_outputs(3172) <= not a;
    layer1_outputs(3173) <= a and not b;
    layer1_outputs(3174) <= b;
    layer1_outputs(3175) <= a;
    layer1_outputs(3176) <= a and not b;
    layer1_outputs(3177) <= not (a or b);
    layer1_outputs(3178) <= b and not a;
    layer1_outputs(3179) <= a;
    layer1_outputs(3180) <= not b;
    layer1_outputs(3181) <= not b;
    layer1_outputs(3182) <= b;
    layer1_outputs(3183) <= a or b;
    layer1_outputs(3184) <= a;
    layer1_outputs(3185) <= a and b;
    layer1_outputs(3186) <= b;
    layer1_outputs(3187) <= not b;
    layer1_outputs(3188) <= b and not a;
    layer1_outputs(3189) <= a and not b;
    layer1_outputs(3190) <= not a;
    layer1_outputs(3191) <= not a or b;
    layer1_outputs(3192) <= a or b;
    layer1_outputs(3193) <= a and b;
    layer1_outputs(3194) <= a;
    layer1_outputs(3195) <= not b;
    layer1_outputs(3196) <= a and b;
    layer1_outputs(3197) <= not b;
    layer1_outputs(3198) <= not a;
    layer1_outputs(3199) <= not b;
    layer1_outputs(3200) <= not a;
    layer1_outputs(3201) <= a;
    layer1_outputs(3202) <= not a;
    layer1_outputs(3203) <= not a or b;
    layer1_outputs(3204) <= b;
    layer1_outputs(3205) <= not a or b;
    layer1_outputs(3206) <= not a;
    layer1_outputs(3207) <= a;
    layer1_outputs(3208) <= not b or a;
    layer1_outputs(3209) <= 1'b1;
    layer1_outputs(3210) <= a and b;
    layer1_outputs(3211) <= b;
    layer1_outputs(3212) <= not b or a;
    layer1_outputs(3213) <= b;
    layer1_outputs(3214) <= not b;
    layer1_outputs(3215) <= not a or b;
    layer1_outputs(3216) <= not (a or b);
    layer1_outputs(3217) <= a and not b;
    layer1_outputs(3218) <= b and not a;
    layer1_outputs(3219) <= not (a or b);
    layer1_outputs(3220) <= a and b;
    layer1_outputs(3221) <= not a or b;
    layer1_outputs(3222) <= a xor b;
    layer1_outputs(3223) <= not b;
    layer1_outputs(3224) <= not (a xor b);
    layer1_outputs(3225) <= a;
    layer1_outputs(3226) <= not a or b;
    layer1_outputs(3227) <= not (a and b);
    layer1_outputs(3228) <= not a;
    layer1_outputs(3229) <= a;
    layer1_outputs(3230) <= a;
    layer1_outputs(3231) <= 1'b0;
    layer1_outputs(3232) <= a and not b;
    layer1_outputs(3233) <= b;
    layer1_outputs(3234) <= a;
    layer1_outputs(3235) <= not a or b;
    layer1_outputs(3236) <= not (a or b);
    layer1_outputs(3237) <= a and not b;
    layer1_outputs(3238) <= a;
    layer1_outputs(3239) <= not b;
    layer1_outputs(3240) <= a xor b;
    layer1_outputs(3241) <= not (a xor b);
    layer1_outputs(3242) <= not (a and b);
    layer1_outputs(3243) <= a and not b;
    layer1_outputs(3244) <= not (a or b);
    layer1_outputs(3245) <= a and not b;
    layer1_outputs(3246) <= a and b;
    layer1_outputs(3247) <= a or b;
    layer1_outputs(3248) <= not b;
    layer1_outputs(3249) <= 1'b1;
    layer1_outputs(3250) <= 1'b0;
    layer1_outputs(3251) <= a or b;
    layer1_outputs(3252) <= not b;
    layer1_outputs(3253) <= a and b;
    layer1_outputs(3254) <= not a or b;
    layer1_outputs(3255) <= not b;
    layer1_outputs(3256) <= a and b;
    layer1_outputs(3257) <= not a;
    layer1_outputs(3258) <= not a or b;
    layer1_outputs(3259) <= 1'b0;
    layer1_outputs(3260) <= b and not a;
    layer1_outputs(3261) <= not b or a;
    layer1_outputs(3262) <= a xor b;
    layer1_outputs(3263) <= not (a and b);
    layer1_outputs(3264) <= a;
    layer1_outputs(3265) <= a;
    layer1_outputs(3266) <= not (a and b);
    layer1_outputs(3267) <= b and not a;
    layer1_outputs(3268) <= not (a or b);
    layer1_outputs(3269) <= not a;
    layer1_outputs(3270) <= b and not a;
    layer1_outputs(3271) <= b and not a;
    layer1_outputs(3272) <= a and b;
    layer1_outputs(3273) <= a;
    layer1_outputs(3274) <= not a;
    layer1_outputs(3275) <= a;
    layer1_outputs(3276) <= not b or a;
    layer1_outputs(3277) <= b and not a;
    layer1_outputs(3278) <= not a;
    layer1_outputs(3279) <= a xor b;
    layer1_outputs(3280) <= not a;
    layer1_outputs(3281) <= a;
    layer1_outputs(3282) <= not (a xor b);
    layer1_outputs(3283) <= b and not a;
    layer1_outputs(3284) <= not b;
    layer1_outputs(3285) <= b;
    layer1_outputs(3286) <= not a or b;
    layer1_outputs(3287) <= a;
    layer1_outputs(3288) <= not b;
    layer1_outputs(3289) <= not (a and b);
    layer1_outputs(3290) <= b and not a;
    layer1_outputs(3291) <= a xor b;
    layer1_outputs(3292) <= not (a and b);
    layer1_outputs(3293) <= not a or b;
    layer1_outputs(3294) <= b and not a;
    layer1_outputs(3295) <= 1'b0;
    layer1_outputs(3296) <= b and not a;
    layer1_outputs(3297) <= a and not b;
    layer1_outputs(3298) <= not (a or b);
    layer1_outputs(3299) <= b and not a;
    layer1_outputs(3300) <= not b;
    layer1_outputs(3301) <= not a or b;
    layer1_outputs(3302) <= not (a and b);
    layer1_outputs(3303) <= a;
    layer1_outputs(3304) <= b and not a;
    layer1_outputs(3305) <= a xor b;
    layer1_outputs(3306) <= a and b;
    layer1_outputs(3307) <= not (a or b);
    layer1_outputs(3308) <= not (a xor b);
    layer1_outputs(3309) <= b and not a;
    layer1_outputs(3310) <= b;
    layer1_outputs(3311) <= not b or a;
    layer1_outputs(3312) <= a and not b;
    layer1_outputs(3313) <= a or b;
    layer1_outputs(3314) <= not a;
    layer1_outputs(3315) <= a and b;
    layer1_outputs(3316) <= not a;
    layer1_outputs(3317) <= 1'b0;
    layer1_outputs(3318) <= 1'b0;
    layer1_outputs(3319) <= not a or b;
    layer1_outputs(3320) <= not a;
    layer1_outputs(3321) <= not (a and b);
    layer1_outputs(3322) <= a;
    layer1_outputs(3323) <= 1'b1;
    layer1_outputs(3324) <= not b;
    layer1_outputs(3325) <= not (a xor b);
    layer1_outputs(3326) <= not (a or b);
    layer1_outputs(3327) <= not a or b;
    layer1_outputs(3328) <= a and not b;
    layer1_outputs(3329) <= not b or a;
    layer1_outputs(3330) <= not b or a;
    layer1_outputs(3331) <= a;
    layer1_outputs(3332) <= not b;
    layer1_outputs(3333) <= a or b;
    layer1_outputs(3334) <= a and b;
    layer1_outputs(3335) <= 1'b0;
    layer1_outputs(3336) <= b and not a;
    layer1_outputs(3337) <= a and b;
    layer1_outputs(3338) <= a;
    layer1_outputs(3339) <= not b or a;
    layer1_outputs(3340) <= not a or b;
    layer1_outputs(3341) <= not a;
    layer1_outputs(3342) <= a and b;
    layer1_outputs(3343) <= not b;
    layer1_outputs(3344) <= a or b;
    layer1_outputs(3345) <= not (a xor b);
    layer1_outputs(3346) <= a or b;
    layer1_outputs(3347) <= not b or a;
    layer1_outputs(3348) <= not (a xor b);
    layer1_outputs(3349) <= 1'b0;
    layer1_outputs(3350) <= b;
    layer1_outputs(3351) <= a;
    layer1_outputs(3352) <= not b or a;
    layer1_outputs(3353) <= b and not a;
    layer1_outputs(3354) <= a and b;
    layer1_outputs(3355) <= not b or a;
    layer1_outputs(3356) <= a;
    layer1_outputs(3357) <= 1'b0;
    layer1_outputs(3358) <= not a;
    layer1_outputs(3359) <= b;
    layer1_outputs(3360) <= a;
    layer1_outputs(3361) <= not a;
    layer1_outputs(3362) <= b;
    layer1_outputs(3363) <= 1'b0;
    layer1_outputs(3364) <= b;
    layer1_outputs(3365) <= a or b;
    layer1_outputs(3366) <= not (a and b);
    layer1_outputs(3367) <= not (a xor b);
    layer1_outputs(3368) <= b;
    layer1_outputs(3369) <= a and b;
    layer1_outputs(3370) <= not (a xor b);
    layer1_outputs(3371) <= not b;
    layer1_outputs(3372) <= a or b;
    layer1_outputs(3373) <= not b;
    layer1_outputs(3374) <= a and b;
    layer1_outputs(3375) <= b;
    layer1_outputs(3376) <= b;
    layer1_outputs(3377) <= not b or a;
    layer1_outputs(3378) <= not b or a;
    layer1_outputs(3379) <= not b;
    layer1_outputs(3380) <= not b;
    layer1_outputs(3381) <= not (a or b);
    layer1_outputs(3382) <= 1'b1;
    layer1_outputs(3383) <= not (a and b);
    layer1_outputs(3384) <= not a or b;
    layer1_outputs(3385) <= not b or a;
    layer1_outputs(3386) <= a and b;
    layer1_outputs(3387) <= not a;
    layer1_outputs(3388) <= not a or b;
    layer1_outputs(3389) <= not (a and b);
    layer1_outputs(3390) <= b;
    layer1_outputs(3391) <= not (a xor b);
    layer1_outputs(3392) <= not a;
    layer1_outputs(3393) <= a;
    layer1_outputs(3394) <= not (a or b);
    layer1_outputs(3395) <= a;
    layer1_outputs(3396) <= 1'b0;
    layer1_outputs(3397) <= a;
    layer1_outputs(3398) <= not (a and b);
    layer1_outputs(3399) <= a and not b;
    layer1_outputs(3400) <= not b or a;
    layer1_outputs(3401) <= a and not b;
    layer1_outputs(3402) <= not a;
    layer1_outputs(3403) <= not (a and b);
    layer1_outputs(3404) <= not a or b;
    layer1_outputs(3405) <= not b;
    layer1_outputs(3406) <= not a;
    layer1_outputs(3407) <= b and not a;
    layer1_outputs(3408) <= not (a or b);
    layer1_outputs(3409) <= not b;
    layer1_outputs(3410) <= not (a or b);
    layer1_outputs(3411) <= not a or b;
    layer1_outputs(3412) <= a xor b;
    layer1_outputs(3413) <= b;
    layer1_outputs(3414) <= b;
    layer1_outputs(3415) <= not a;
    layer1_outputs(3416) <= a and b;
    layer1_outputs(3417) <= 1'b0;
    layer1_outputs(3418) <= not a or b;
    layer1_outputs(3419) <= not (a or b);
    layer1_outputs(3420) <= b;
    layer1_outputs(3421) <= b;
    layer1_outputs(3422) <= not b;
    layer1_outputs(3423) <= b;
    layer1_outputs(3424) <= a and b;
    layer1_outputs(3425) <= 1'b0;
    layer1_outputs(3426) <= a and b;
    layer1_outputs(3427) <= a;
    layer1_outputs(3428) <= 1'b0;
    layer1_outputs(3429) <= not a;
    layer1_outputs(3430) <= a xor b;
    layer1_outputs(3431) <= not (a and b);
    layer1_outputs(3432) <= not a;
    layer1_outputs(3433) <= 1'b1;
    layer1_outputs(3434) <= a or b;
    layer1_outputs(3435) <= a;
    layer1_outputs(3436) <= a and b;
    layer1_outputs(3437) <= not b;
    layer1_outputs(3438) <= not (a or b);
    layer1_outputs(3439) <= 1'b0;
    layer1_outputs(3440) <= not b or a;
    layer1_outputs(3441) <= not b;
    layer1_outputs(3442) <= b and not a;
    layer1_outputs(3443) <= not b;
    layer1_outputs(3444) <= a and b;
    layer1_outputs(3445) <= not a;
    layer1_outputs(3446) <= 1'b1;
    layer1_outputs(3447) <= a xor b;
    layer1_outputs(3448) <= b;
    layer1_outputs(3449) <= a;
    layer1_outputs(3450) <= a or b;
    layer1_outputs(3451) <= not a or b;
    layer1_outputs(3452) <= a and not b;
    layer1_outputs(3453) <= not (a xor b);
    layer1_outputs(3454) <= not a;
    layer1_outputs(3455) <= a or b;
    layer1_outputs(3456) <= not (a xor b);
    layer1_outputs(3457) <= 1'b1;
    layer1_outputs(3458) <= not (a xor b);
    layer1_outputs(3459) <= b;
    layer1_outputs(3460) <= a or b;
    layer1_outputs(3461) <= not b;
    layer1_outputs(3462) <= a and b;
    layer1_outputs(3463) <= not a;
    layer1_outputs(3464) <= not a;
    layer1_outputs(3465) <= b;
    layer1_outputs(3466) <= not b;
    layer1_outputs(3467) <= b;
    layer1_outputs(3468) <= b;
    layer1_outputs(3469) <= a;
    layer1_outputs(3470) <= 1'b0;
    layer1_outputs(3471) <= not a;
    layer1_outputs(3472) <= not (a and b);
    layer1_outputs(3473) <= not b;
    layer1_outputs(3474) <= not a;
    layer1_outputs(3475) <= b;
    layer1_outputs(3476) <= a or b;
    layer1_outputs(3477) <= not a;
    layer1_outputs(3478) <= b;
    layer1_outputs(3479) <= not a;
    layer1_outputs(3480) <= 1'b1;
    layer1_outputs(3481) <= not (a xor b);
    layer1_outputs(3482) <= not b or a;
    layer1_outputs(3483) <= a and b;
    layer1_outputs(3484) <= not b;
    layer1_outputs(3485) <= not (a or b);
    layer1_outputs(3486) <= not (a and b);
    layer1_outputs(3487) <= 1'b0;
    layer1_outputs(3488) <= not b;
    layer1_outputs(3489) <= not (a or b);
    layer1_outputs(3490) <= not (a xor b);
    layer1_outputs(3491) <= b;
    layer1_outputs(3492) <= not b or a;
    layer1_outputs(3493) <= a;
    layer1_outputs(3494) <= not a;
    layer1_outputs(3495) <= a or b;
    layer1_outputs(3496) <= b and not a;
    layer1_outputs(3497) <= not b;
    layer1_outputs(3498) <= a and b;
    layer1_outputs(3499) <= a and b;
    layer1_outputs(3500) <= not a;
    layer1_outputs(3501) <= not b or a;
    layer1_outputs(3502) <= not b;
    layer1_outputs(3503) <= a xor b;
    layer1_outputs(3504) <= a and not b;
    layer1_outputs(3505) <= a xor b;
    layer1_outputs(3506) <= not (a or b);
    layer1_outputs(3507) <= not a;
    layer1_outputs(3508) <= a and not b;
    layer1_outputs(3509) <= not a or b;
    layer1_outputs(3510) <= not a or b;
    layer1_outputs(3511) <= not b or a;
    layer1_outputs(3512) <= not b or a;
    layer1_outputs(3513) <= b;
    layer1_outputs(3514) <= b;
    layer1_outputs(3515) <= b;
    layer1_outputs(3516) <= 1'b0;
    layer1_outputs(3517) <= a and b;
    layer1_outputs(3518) <= not a or b;
    layer1_outputs(3519) <= not a or b;
    layer1_outputs(3520) <= not b or a;
    layer1_outputs(3521) <= 1'b0;
    layer1_outputs(3522) <= 1'b0;
    layer1_outputs(3523) <= a and b;
    layer1_outputs(3524) <= not a;
    layer1_outputs(3525) <= b;
    layer1_outputs(3526) <= b;
    layer1_outputs(3527) <= b and not a;
    layer1_outputs(3528) <= not b;
    layer1_outputs(3529) <= b;
    layer1_outputs(3530) <= 1'b0;
    layer1_outputs(3531) <= 1'b1;
    layer1_outputs(3532) <= 1'b1;
    layer1_outputs(3533) <= b;
    layer1_outputs(3534) <= b;
    layer1_outputs(3535) <= a and not b;
    layer1_outputs(3536) <= b;
    layer1_outputs(3537) <= not b or a;
    layer1_outputs(3538) <= not (a or b);
    layer1_outputs(3539) <= not a or b;
    layer1_outputs(3540) <= b;
    layer1_outputs(3541) <= b;
    layer1_outputs(3542) <= not b;
    layer1_outputs(3543) <= not a or b;
    layer1_outputs(3544) <= not b;
    layer1_outputs(3545) <= a;
    layer1_outputs(3546) <= not (a or b);
    layer1_outputs(3547) <= not a;
    layer1_outputs(3548) <= not (a or b);
    layer1_outputs(3549) <= 1'b1;
    layer1_outputs(3550) <= not a;
    layer1_outputs(3551) <= a;
    layer1_outputs(3552) <= not b or a;
    layer1_outputs(3553) <= not b or a;
    layer1_outputs(3554) <= not a or b;
    layer1_outputs(3555) <= a xor b;
    layer1_outputs(3556) <= a and b;
    layer1_outputs(3557) <= a xor b;
    layer1_outputs(3558) <= a or b;
    layer1_outputs(3559) <= a or b;
    layer1_outputs(3560) <= not b or a;
    layer1_outputs(3561) <= b;
    layer1_outputs(3562) <= 1'b0;
    layer1_outputs(3563) <= not b or a;
    layer1_outputs(3564) <= not (a or b);
    layer1_outputs(3565) <= a and not b;
    layer1_outputs(3566) <= a;
    layer1_outputs(3567) <= not b;
    layer1_outputs(3568) <= not (a or b);
    layer1_outputs(3569) <= b and not a;
    layer1_outputs(3570) <= a;
    layer1_outputs(3571) <= not (a xor b);
    layer1_outputs(3572) <= a or b;
    layer1_outputs(3573) <= not (a or b);
    layer1_outputs(3574) <= not a;
    layer1_outputs(3575) <= not b;
    layer1_outputs(3576) <= not b;
    layer1_outputs(3577) <= a or b;
    layer1_outputs(3578) <= not (a xor b);
    layer1_outputs(3579) <= not a;
    layer1_outputs(3580) <= a and b;
    layer1_outputs(3581) <= a and b;
    layer1_outputs(3582) <= a or b;
    layer1_outputs(3583) <= not (a xor b);
    layer1_outputs(3584) <= not a;
    layer1_outputs(3585) <= b;
    layer1_outputs(3586) <= not b or a;
    layer1_outputs(3587) <= not (a xor b);
    layer1_outputs(3588) <= a xor b;
    layer1_outputs(3589) <= b and not a;
    layer1_outputs(3590) <= b and not a;
    layer1_outputs(3591) <= not (a and b);
    layer1_outputs(3592) <= a xor b;
    layer1_outputs(3593) <= not a;
    layer1_outputs(3594) <= a and not b;
    layer1_outputs(3595) <= not (a xor b);
    layer1_outputs(3596) <= not a;
    layer1_outputs(3597) <= not a;
    layer1_outputs(3598) <= not a;
    layer1_outputs(3599) <= not (a xor b);
    layer1_outputs(3600) <= not a or b;
    layer1_outputs(3601) <= a and b;
    layer1_outputs(3602) <= not a or b;
    layer1_outputs(3603) <= a and not b;
    layer1_outputs(3604) <= not (a or b);
    layer1_outputs(3605) <= b;
    layer1_outputs(3606) <= not b;
    layer1_outputs(3607) <= a xor b;
    layer1_outputs(3608) <= a and not b;
    layer1_outputs(3609) <= not (a and b);
    layer1_outputs(3610) <= a and b;
    layer1_outputs(3611) <= a and b;
    layer1_outputs(3612) <= a or b;
    layer1_outputs(3613) <= a;
    layer1_outputs(3614) <= a and b;
    layer1_outputs(3615) <= b;
    layer1_outputs(3616) <= not b or a;
    layer1_outputs(3617) <= a and not b;
    layer1_outputs(3618) <= a or b;
    layer1_outputs(3619) <= not (a or b);
    layer1_outputs(3620) <= 1'b1;
    layer1_outputs(3621) <= b;
    layer1_outputs(3622) <= not b;
    layer1_outputs(3623) <= not b or a;
    layer1_outputs(3624) <= b;
    layer1_outputs(3625) <= 1'b0;
    layer1_outputs(3626) <= a and not b;
    layer1_outputs(3627) <= not a or b;
    layer1_outputs(3628) <= a and b;
    layer1_outputs(3629) <= 1'b1;
    layer1_outputs(3630) <= a;
    layer1_outputs(3631) <= 1'b1;
    layer1_outputs(3632) <= not b or a;
    layer1_outputs(3633) <= not b or a;
    layer1_outputs(3634) <= not b;
    layer1_outputs(3635) <= a xor b;
    layer1_outputs(3636) <= not (a xor b);
    layer1_outputs(3637) <= not b or a;
    layer1_outputs(3638) <= not (a and b);
    layer1_outputs(3639) <= a and not b;
    layer1_outputs(3640) <= not b;
    layer1_outputs(3641) <= not b;
    layer1_outputs(3642) <= not a;
    layer1_outputs(3643) <= not (a or b);
    layer1_outputs(3644) <= not a;
    layer1_outputs(3645) <= a and not b;
    layer1_outputs(3646) <= 1'b1;
    layer1_outputs(3647) <= not a;
    layer1_outputs(3648) <= b and not a;
    layer1_outputs(3649) <= not a;
    layer1_outputs(3650) <= not b or a;
    layer1_outputs(3651) <= not (a or b);
    layer1_outputs(3652) <= 1'b0;
    layer1_outputs(3653) <= a;
    layer1_outputs(3654) <= b;
    layer1_outputs(3655) <= not b or a;
    layer1_outputs(3656) <= b;
    layer1_outputs(3657) <= a and b;
    layer1_outputs(3658) <= not b;
    layer1_outputs(3659) <= 1'b0;
    layer1_outputs(3660) <= not a or b;
    layer1_outputs(3661) <= a or b;
    layer1_outputs(3662) <= not b;
    layer1_outputs(3663) <= a xor b;
    layer1_outputs(3664) <= not a;
    layer1_outputs(3665) <= not (a or b);
    layer1_outputs(3666) <= not (a xor b);
    layer1_outputs(3667) <= not b or a;
    layer1_outputs(3668) <= not b;
    layer1_outputs(3669) <= a xor b;
    layer1_outputs(3670) <= not b or a;
    layer1_outputs(3671) <= b and not a;
    layer1_outputs(3672) <= a or b;
    layer1_outputs(3673) <= b and not a;
    layer1_outputs(3674) <= a and not b;
    layer1_outputs(3675) <= b and not a;
    layer1_outputs(3676) <= b;
    layer1_outputs(3677) <= not a;
    layer1_outputs(3678) <= not b or a;
    layer1_outputs(3679) <= not a;
    layer1_outputs(3680) <= 1'b1;
    layer1_outputs(3681) <= b and not a;
    layer1_outputs(3682) <= a;
    layer1_outputs(3683) <= a and not b;
    layer1_outputs(3684) <= not b;
    layer1_outputs(3685) <= not (a or b);
    layer1_outputs(3686) <= not a;
    layer1_outputs(3687) <= b;
    layer1_outputs(3688) <= not (a or b);
    layer1_outputs(3689) <= not b or a;
    layer1_outputs(3690) <= not b or a;
    layer1_outputs(3691) <= not a;
    layer1_outputs(3692) <= a and not b;
    layer1_outputs(3693) <= not (a or b);
    layer1_outputs(3694) <= a;
    layer1_outputs(3695) <= b;
    layer1_outputs(3696) <= b;
    layer1_outputs(3697) <= a and b;
    layer1_outputs(3698) <= not b;
    layer1_outputs(3699) <= 1'b0;
    layer1_outputs(3700) <= not (a xor b);
    layer1_outputs(3701) <= b and not a;
    layer1_outputs(3702) <= not b;
    layer1_outputs(3703) <= a xor b;
    layer1_outputs(3704) <= not b;
    layer1_outputs(3705) <= b and not a;
    layer1_outputs(3706) <= not b or a;
    layer1_outputs(3707) <= a xor b;
    layer1_outputs(3708) <= not (a xor b);
    layer1_outputs(3709) <= b;
    layer1_outputs(3710) <= 1'b1;
    layer1_outputs(3711) <= a and b;
    layer1_outputs(3712) <= b;
    layer1_outputs(3713) <= a or b;
    layer1_outputs(3714) <= a and not b;
    layer1_outputs(3715) <= a;
    layer1_outputs(3716) <= not b;
    layer1_outputs(3717) <= not (a or b);
    layer1_outputs(3718) <= not a or b;
    layer1_outputs(3719) <= 1'b1;
    layer1_outputs(3720) <= not a or b;
    layer1_outputs(3721) <= not b;
    layer1_outputs(3722) <= a and b;
    layer1_outputs(3723) <= b and not a;
    layer1_outputs(3724) <= b and not a;
    layer1_outputs(3725) <= a;
    layer1_outputs(3726) <= not (a xor b);
    layer1_outputs(3727) <= not b;
    layer1_outputs(3728) <= b;
    layer1_outputs(3729) <= b;
    layer1_outputs(3730) <= b;
    layer1_outputs(3731) <= a or b;
    layer1_outputs(3732) <= not (a or b);
    layer1_outputs(3733) <= not (a xor b);
    layer1_outputs(3734) <= not a;
    layer1_outputs(3735) <= not (a or b);
    layer1_outputs(3736) <= a or b;
    layer1_outputs(3737) <= not b or a;
    layer1_outputs(3738) <= not b;
    layer1_outputs(3739) <= not (a xor b);
    layer1_outputs(3740) <= b;
    layer1_outputs(3741) <= a and not b;
    layer1_outputs(3742) <= a xor b;
    layer1_outputs(3743) <= b;
    layer1_outputs(3744) <= not b or a;
    layer1_outputs(3745) <= not b;
    layer1_outputs(3746) <= a and b;
    layer1_outputs(3747) <= not (a and b);
    layer1_outputs(3748) <= a and not b;
    layer1_outputs(3749) <= a or b;
    layer1_outputs(3750) <= a or b;
    layer1_outputs(3751) <= not b;
    layer1_outputs(3752) <= 1'b1;
    layer1_outputs(3753) <= 1'b1;
    layer1_outputs(3754) <= a and b;
    layer1_outputs(3755) <= not (a xor b);
    layer1_outputs(3756) <= not a or b;
    layer1_outputs(3757) <= 1'b1;
    layer1_outputs(3758) <= b;
    layer1_outputs(3759) <= b;
    layer1_outputs(3760) <= a and b;
    layer1_outputs(3761) <= not b or a;
    layer1_outputs(3762) <= 1'b0;
    layer1_outputs(3763) <= a and not b;
    layer1_outputs(3764) <= not a or b;
    layer1_outputs(3765) <= not b;
    layer1_outputs(3766) <= b;
    layer1_outputs(3767) <= not b;
    layer1_outputs(3768) <= b;
    layer1_outputs(3769) <= not (a and b);
    layer1_outputs(3770) <= not b or a;
    layer1_outputs(3771) <= a and not b;
    layer1_outputs(3772) <= a;
    layer1_outputs(3773) <= a and not b;
    layer1_outputs(3774) <= not (a and b);
    layer1_outputs(3775) <= not b;
    layer1_outputs(3776) <= not (a or b);
    layer1_outputs(3777) <= not a or b;
    layer1_outputs(3778) <= a and not b;
    layer1_outputs(3779) <= b;
    layer1_outputs(3780) <= not (a or b);
    layer1_outputs(3781) <= 1'b0;
    layer1_outputs(3782) <= not b;
    layer1_outputs(3783) <= a or b;
    layer1_outputs(3784) <= b;
    layer1_outputs(3785) <= 1'b0;
    layer1_outputs(3786) <= b and not a;
    layer1_outputs(3787) <= 1'b1;
    layer1_outputs(3788) <= not (a xor b);
    layer1_outputs(3789) <= b;
    layer1_outputs(3790) <= b;
    layer1_outputs(3791) <= a or b;
    layer1_outputs(3792) <= b;
    layer1_outputs(3793) <= a xor b;
    layer1_outputs(3794) <= a and b;
    layer1_outputs(3795) <= a and b;
    layer1_outputs(3796) <= not (a or b);
    layer1_outputs(3797) <= a or b;
    layer1_outputs(3798) <= not b;
    layer1_outputs(3799) <= not a or b;
    layer1_outputs(3800) <= a xor b;
    layer1_outputs(3801) <= a or b;
    layer1_outputs(3802) <= a and b;
    layer1_outputs(3803) <= not a or b;
    layer1_outputs(3804) <= a and not b;
    layer1_outputs(3805) <= not a or b;
    layer1_outputs(3806) <= b;
    layer1_outputs(3807) <= not a;
    layer1_outputs(3808) <= not (a and b);
    layer1_outputs(3809) <= a xor b;
    layer1_outputs(3810) <= not (a and b);
    layer1_outputs(3811) <= a and not b;
    layer1_outputs(3812) <= not b;
    layer1_outputs(3813) <= a xor b;
    layer1_outputs(3814) <= not (a and b);
    layer1_outputs(3815) <= a;
    layer1_outputs(3816) <= not b;
    layer1_outputs(3817) <= a and b;
    layer1_outputs(3818) <= not a;
    layer1_outputs(3819) <= not a;
    layer1_outputs(3820) <= not a;
    layer1_outputs(3821) <= a and b;
    layer1_outputs(3822) <= a and b;
    layer1_outputs(3823) <= 1'b0;
    layer1_outputs(3824) <= not (a and b);
    layer1_outputs(3825) <= a;
    layer1_outputs(3826) <= not (a xor b);
    layer1_outputs(3827) <= not (a and b);
    layer1_outputs(3828) <= b;
    layer1_outputs(3829) <= a or b;
    layer1_outputs(3830) <= not a;
    layer1_outputs(3831) <= not (a and b);
    layer1_outputs(3832) <= not a;
    layer1_outputs(3833) <= a and b;
    layer1_outputs(3834) <= not b;
    layer1_outputs(3835) <= a;
    layer1_outputs(3836) <= a;
    layer1_outputs(3837) <= not a;
    layer1_outputs(3838) <= b;
    layer1_outputs(3839) <= not a;
    layer1_outputs(3840) <= not b or a;
    layer1_outputs(3841) <= 1'b1;
    layer1_outputs(3842) <= a xor b;
    layer1_outputs(3843) <= a xor b;
    layer1_outputs(3844) <= b;
    layer1_outputs(3845) <= not b;
    layer1_outputs(3846) <= not a;
    layer1_outputs(3847) <= not a or b;
    layer1_outputs(3848) <= not a;
    layer1_outputs(3849) <= 1'b0;
    layer1_outputs(3850) <= b and not a;
    layer1_outputs(3851) <= a xor b;
    layer1_outputs(3852) <= not b;
    layer1_outputs(3853) <= a xor b;
    layer1_outputs(3854) <= not a;
    layer1_outputs(3855) <= b;
    layer1_outputs(3856) <= not a;
    layer1_outputs(3857) <= b;
    layer1_outputs(3858) <= not (a or b);
    layer1_outputs(3859) <= not a or b;
    layer1_outputs(3860) <= not (a or b);
    layer1_outputs(3861) <= a xor b;
    layer1_outputs(3862) <= not (a xor b);
    layer1_outputs(3863) <= a xor b;
    layer1_outputs(3864) <= a and not b;
    layer1_outputs(3865) <= b;
    layer1_outputs(3866) <= not b or a;
    layer1_outputs(3867) <= b;
    layer1_outputs(3868) <= a;
    layer1_outputs(3869) <= not (a and b);
    layer1_outputs(3870) <= not b;
    layer1_outputs(3871) <= not (a and b);
    layer1_outputs(3872) <= b and not a;
    layer1_outputs(3873) <= not b;
    layer1_outputs(3874) <= b and not a;
    layer1_outputs(3875) <= not a or b;
    layer1_outputs(3876) <= 1'b1;
    layer1_outputs(3877) <= a;
    layer1_outputs(3878) <= 1'b0;
    layer1_outputs(3879) <= a;
    layer1_outputs(3880) <= b;
    layer1_outputs(3881) <= a and b;
    layer1_outputs(3882) <= b and not a;
    layer1_outputs(3883) <= not b or a;
    layer1_outputs(3884) <= not b;
    layer1_outputs(3885) <= not a or b;
    layer1_outputs(3886) <= a and not b;
    layer1_outputs(3887) <= b;
    layer1_outputs(3888) <= not (a and b);
    layer1_outputs(3889) <= a or b;
    layer1_outputs(3890) <= a and not b;
    layer1_outputs(3891) <= not (a or b);
    layer1_outputs(3892) <= not b;
    layer1_outputs(3893) <= a and b;
    layer1_outputs(3894) <= a;
    layer1_outputs(3895) <= a or b;
    layer1_outputs(3896) <= a;
    layer1_outputs(3897) <= not (a and b);
    layer1_outputs(3898) <= a;
    layer1_outputs(3899) <= a xor b;
    layer1_outputs(3900) <= not (a xor b);
    layer1_outputs(3901) <= a and not b;
    layer1_outputs(3902) <= a or b;
    layer1_outputs(3903) <= b and not a;
    layer1_outputs(3904) <= not (a xor b);
    layer1_outputs(3905) <= not (a or b);
    layer1_outputs(3906) <= a or b;
    layer1_outputs(3907) <= 1'b1;
    layer1_outputs(3908) <= not b or a;
    layer1_outputs(3909) <= not b or a;
    layer1_outputs(3910) <= a xor b;
    layer1_outputs(3911) <= 1'b0;
    layer1_outputs(3912) <= a or b;
    layer1_outputs(3913) <= not a or b;
    layer1_outputs(3914) <= a xor b;
    layer1_outputs(3915) <= not (a and b);
    layer1_outputs(3916) <= not b;
    layer1_outputs(3917) <= a or b;
    layer1_outputs(3918) <= a xor b;
    layer1_outputs(3919) <= 1'b0;
    layer1_outputs(3920) <= a and b;
    layer1_outputs(3921) <= not b;
    layer1_outputs(3922) <= a;
    layer1_outputs(3923) <= 1'b0;
    layer1_outputs(3924) <= not b;
    layer1_outputs(3925) <= a or b;
    layer1_outputs(3926) <= not (a xor b);
    layer1_outputs(3927) <= b;
    layer1_outputs(3928) <= a and b;
    layer1_outputs(3929) <= 1'b0;
    layer1_outputs(3930) <= not a or b;
    layer1_outputs(3931) <= a xor b;
    layer1_outputs(3932) <= a and not b;
    layer1_outputs(3933) <= not (a or b);
    layer1_outputs(3934) <= not a or b;
    layer1_outputs(3935) <= b;
    layer1_outputs(3936) <= a and not b;
    layer1_outputs(3937) <= not a;
    layer1_outputs(3938) <= not b;
    layer1_outputs(3939) <= not a;
    layer1_outputs(3940) <= not b;
    layer1_outputs(3941) <= a and not b;
    layer1_outputs(3942) <= b and not a;
    layer1_outputs(3943) <= a;
    layer1_outputs(3944) <= not a;
    layer1_outputs(3945) <= a;
    layer1_outputs(3946) <= a xor b;
    layer1_outputs(3947) <= not (a or b);
    layer1_outputs(3948) <= a and b;
    layer1_outputs(3949) <= 1'b1;
    layer1_outputs(3950) <= not (a xor b);
    layer1_outputs(3951) <= not (a and b);
    layer1_outputs(3952) <= b;
    layer1_outputs(3953) <= 1'b0;
    layer1_outputs(3954) <= not b;
    layer1_outputs(3955) <= not a or b;
    layer1_outputs(3956) <= not (a or b);
    layer1_outputs(3957) <= a xor b;
    layer1_outputs(3958) <= not a or b;
    layer1_outputs(3959) <= not b or a;
    layer1_outputs(3960) <= b;
    layer1_outputs(3961) <= not b;
    layer1_outputs(3962) <= a;
    layer1_outputs(3963) <= not a;
    layer1_outputs(3964) <= a and not b;
    layer1_outputs(3965) <= not a;
    layer1_outputs(3966) <= a and b;
    layer1_outputs(3967) <= not a or b;
    layer1_outputs(3968) <= not b;
    layer1_outputs(3969) <= not a;
    layer1_outputs(3970) <= not (a and b);
    layer1_outputs(3971) <= not a;
    layer1_outputs(3972) <= a;
    layer1_outputs(3973) <= not (a xor b);
    layer1_outputs(3974) <= a and not b;
    layer1_outputs(3975) <= not a or b;
    layer1_outputs(3976) <= a xor b;
    layer1_outputs(3977) <= a xor b;
    layer1_outputs(3978) <= not b;
    layer1_outputs(3979) <= a or b;
    layer1_outputs(3980) <= not (a or b);
    layer1_outputs(3981) <= a;
    layer1_outputs(3982) <= not a or b;
    layer1_outputs(3983) <= not (a and b);
    layer1_outputs(3984) <= 1'b1;
    layer1_outputs(3985) <= a and not b;
    layer1_outputs(3986) <= not b or a;
    layer1_outputs(3987) <= a;
    layer1_outputs(3988) <= not b or a;
    layer1_outputs(3989) <= not (a and b);
    layer1_outputs(3990) <= not b or a;
    layer1_outputs(3991) <= not (a or b);
    layer1_outputs(3992) <= not (a and b);
    layer1_outputs(3993) <= 1'b0;
    layer1_outputs(3994) <= not a;
    layer1_outputs(3995) <= not b;
    layer1_outputs(3996) <= not a or b;
    layer1_outputs(3997) <= a and b;
    layer1_outputs(3998) <= not a or b;
    layer1_outputs(3999) <= a and not b;
    layer1_outputs(4000) <= 1'b0;
    layer1_outputs(4001) <= a xor b;
    layer1_outputs(4002) <= not (a or b);
    layer1_outputs(4003) <= b and not a;
    layer1_outputs(4004) <= not (a and b);
    layer1_outputs(4005) <= b;
    layer1_outputs(4006) <= a and not b;
    layer1_outputs(4007) <= not b;
    layer1_outputs(4008) <= 1'b1;
    layer1_outputs(4009) <= b;
    layer1_outputs(4010) <= not (a xor b);
    layer1_outputs(4011) <= not (a and b);
    layer1_outputs(4012) <= a or b;
    layer1_outputs(4013) <= a and b;
    layer1_outputs(4014) <= a or b;
    layer1_outputs(4015) <= 1'b1;
    layer1_outputs(4016) <= b and not a;
    layer1_outputs(4017) <= not b;
    layer1_outputs(4018) <= not a or b;
    layer1_outputs(4019) <= b;
    layer1_outputs(4020) <= a or b;
    layer1_outputs(4021) <= 1'b0;
    layer1_outputs(4022) <= not (a and b);
    layer1_outputs(4023) <= not a or b;
    layer1_outputs(4024) <= a;
    layer1_outputs(4025) <= 1'b1;
    layer1_outputs(4026) <= a and b;
    layer1_outputs(4027) <= not (a xor b);
    layer1_outputs(4028) <= not a or b;
    layer1_outputs(4029) <= not (a and b);
    layer1_outputs(4030) <= b;
    layer1_outputs(4031) <= a or b;
    layer1_outputs(4032) <= a xor b;
    layer1_outputs(4033) <= b and not a;
    layer1_outputs(4034) <= not b;
    layer1_outputs(4035) <= 1'b0;
    layer1_outputs(4036) <= 1'b0;
    layer1_outputs(4037) <= b;
    layer1_outputs(4038) <= a and not b;
    layer1_outputs(4039) <= not b;
    layer1_outputs(4040) <= b and not a;
    layer1_outputs(4041) <= not a or b;
    layer1_outputs(4042) <= b;
    layer1_outputs(4043) <= b;
    layer1_outputs(4044) <= not b or a;
    layer1_outputs(4045) <= a and not b;
    layer1_outputs(4046) <= a xor b;
    layer1_outputs(4047) <= b and not a;
    layer1_outputs(4048) <= a and not b;
    layer1_outputs(4049) <= 1'b0;
    layer1_outputs(4050) <= a xor b;
    layer1_outputs(4051) <= a or b;
    layer1_outputs(4052) <= not b;
    layer1_outputs(4053) <= b and not a;
    layer1_outputs(4054) <= a;
    layer1_outputs(4055) <= a or b;
    layer1_outputs(4056) <= not b;
    layer1_outputs(4057) <= 1'b0;
    layer1_outputs(4058) <= not a or b;
    layer1_outputs(4059) <= a and not b;
    layer1_outputs(4060) <= 1'b0;
    layer1_outputs(4061) <= not a;
    layer1_outputs(4062) <= a and b;
    layer1_outputs(4063) <= b;
    layer1_outputs(4064) <= a xor b;
    layer1_outputs(4065) <= b;
    layer1_outputs(4066) <= a and not b;
    layer1_outputs(4067) <= b;
    layer1_outputs(4068) <= a and not b;
    layer1_outputs(4069) <= b and not a;
    layer1_outputs(4070) <= a and b;
    layer1_outputs(4071) <= not (a or b);
    layer1_outputs(4072) <= not a;
    layer1_outputs(4073) <= 1'b1;
    layer1_outputs(4074) <= 1'b1;
    layer1_outputs(4075) <= b;
    layer1_outputs(4076) <= not (a or b);
    layer1_outputs(4077) <= 1'b1;
    layer1_outputs(4078) <= not b;
    layer1_outputs(4079) <= 1'b0;
    layer1_outputs(4080) <= a;
    layer1_outputs(4081) <= a and b;
    layer1_outputs(4082) <= a;
    layer1_outputs(4083) <= not (a or b);
    layer1_outputs(4084) <= a and not b;
    layer1_outputs(4085) <= a;
    layer1_outputs(4086) <= 1'b1;
    layer1_outputs(4087) <= a and b;
    layer1_outputs(4088) <= b and not a;
    layer1_outputs(4089) <= b and not a;
    layer1_outputs(4090) <= a and b;
    layer1_outputs(4091) <= a and b;
    layer1_outputs(4092) <= not a;
    layer1_outputs(4093) <= a and not b;
    layer1_outputs(4094) <= a or b;
    layer1_outputs(4095) <= b;
    layer1_outputs(4096) <= 1'b0;
    layer1_outputs(4097) <= b and not a;
    layer1_outputs(4098) <= not (a and b);
    layer1_outputs(4099) <= not a;
    layer1_outputs(4100) <= not b;
    layer1_outputs(4101) <= b;
    layer1_outputs(4102) <= b;
    layer1_outputs(4103) <= not (a and b);
    layer1_outputs(4104) <= a;
    layer1_outputs(4105) <= not b or a;
    layer1_outputs(4106) <= a;
    layer1_outputs(4107) <= not a;
    layer1_outputs(4108) <= not b or a;
    layer1_outputs(4109) <= a and b;
    layer1_outputs(4110) <= not b or a;
    layer1_outputs(4111) <= not b;
    layer1_outputs(4112) <= b;
    layer1_outputs(4113) <= a and not b;
    layer1_outputs(4114) <= not a or b;
    layer1_outputs(4115) <= not b or a;
    layer1_outputs(4116) <= a and b;
    layer1_outputs(4117) <= a;
    layer1_outputs(4118) <= 1'b0;
    layer1_outputs(4119) <= b and not a;
    layer1_outputs(4120) <= not (a and b);
    layer1_outputs(4121) <= a xor b;
    layer1_outputs(4122) <= b and not a;
    layer1_outputs(4123) <= b;
    layer1_outputs(4124) <= 1'b1;
    layer1_outputs(4125) <= a or b;
    layer1_outputs(4126) <= b and not a;
    layer1_outputs(4127) <= a and b;
    layer1_outputs(4128) <= a and b;
    layer1_outputs(4129) <= not a;
    layer1_outputs(4130) <= 1'b1;
    layer1_outputs(4131) <= a;
    layer1_outputs(4132) <= not (a xor b);
    layer1_outputs(4133) <= not a or b;
    layer1_outputs(4134) <= a xor b;
    layer1_outputs(4135) <= not a or b;
    layer1_outputs(4136) <= b;
    layer1_outputs(4137) <= a and b;
    layer1_outputs(4138) <= a and b;
    layer1_outputs(4139) <= not b;
    layer1_outputs(4140) <= b and not a;
    layer1_outputs(4141) <= not b or a;
    layer1_outputs(4142) <= a or b;
    layer1_outputs(4143) <= 1'b1;
    layer1_outputs(4144) <= not b;
    layer1_outputs(4145) <= not a or b;
    layer1_outputs(4146) <= b;
    layer1_outputs(4147) <= not a or b;
    layer1_outputs(4148) <= b and not a;
    layer1_outputs(4149) <= a;
    layer1_outputs(4150) <= not a;
    layer1_outputs(4151) <= not a or b;
    layer1_outputs(4152) <= a or b;
    layer1_outputs(4153) <= a xor b;
    layer1_outputs(4154) <= not b or a;
    layer1_outputs(4155) <= not (a or b);
    layer1_outputs(4156) <= 1'b1;
    layer1_outputs(4157) <= not b or a;
    layer1_outputs(4158) <= 1'b1;
    layer1_outputs(4159) <= not (a or b);
    layer1_outputs(4160) <= 1'b1;
    layer1_outputs(4161) <= a and b;
    layer1_outputs(4162) <= a and not b;
    layer1_outputs(4163) <= 1'b1;
    layer1_outputs(4164) <= not a or b;
    layer1_outputs(4165) <= not (a and b);
    layer1_outputs(4166) <= a or b;
    layer1_outputs(4167) <= not b or a;
    layer1_outputs(4168) <= b;
    layer1_outputs(4169) <= b;
    layer1_outputs(4170) <= not b;
    layer1_outputs(4171) <= a;
    layer1_outputs(4172) <= not (a and b);
    layer1_outputs(4173) <= not b;
    layer1_outputs(4174) <= a and not b;
    layer1_outputs(4175) <= b;
    layer1_outputs(4176) <= a;
    layer1_outputs(4177) <= not a or b;
    layer1_outputs(4178) <= not (a and b);
    layer1_outputs(4179) <= b and not a;
    layer1_outputs(4180) <= not b;
    layer1_outputs(4181) <= not b or a;
    layer1_outputs(4182) <= not b or a;
    layer1_outputs(4183) <= not a;
    layer1_outputs(4184) <= not (a and b);
    layer1_outputs(4185) <= not b;
    layer1_outputs(4186) <= a;
    layer1_outputs(4187) <= 1'b0;
    layer1_outputs(4188) <= not a or b;
    layer1_outputs(4189) <= 1'b0;
    layer1_outputs(4190) <= not (a xor b);
    layer1_outputs(4191) <= not a;
    layer1_outputs(4192) <= a;
    layer1_outputs(4193) <= not a;
    layer1_outputs(4194) <= a or b;
    layer1_outputs(4195) <= a or b;
    layer1_outputs(4196) <= not b;
    layer1_outputs(4197) <= not b or a;
    layer1_outputs(4198) <= a or b;
    layer1_outputs(4199) <= not b or a;
    layer1_outputs(4200) <= not a;
    layer1_outputs(4201) <= not (a and b);
    layer1_outputs(4202) <= a and not b;
    layer1_outputs(4203) <= not a;
    layer1_outputs(4204) <= b and not a;
    layer1_outputs(4205) <= 1'b0;
    layer1_outputs(4206) <= a or b;
    layer1_outputs(4207) <= not a or b;
    layer1_outputs(4208) <= b and not a;
    layer1_outputs(4209) <= a and not b;
    layer1_outputs(4210) <= a and b;
    layer1_outputs(4211) <= a or b;
    layer1_outputs(4212) <= b;
    layer1_outputs(4213) <= not a or b;
    layer1_outputs(4214) <= b and not a;
    layer1_outputs(4215) <= not (a xor b);
    layer1_outputs(4216) <= a xor b;
    layer1_outputs(4217) <= not a or b;
    layer1_outputs(4218) <= not b;
    layer1_outputs(4219) <= not b;
    layer1_outputs(4220) <= a;
    layer1_outputs(4221) <= a and b;
    layer1_outputs(4222) <= a or b;
    layer1_outputs(4223) <= a;
    layer1_outputs(4224) <= a and not b;
    layer1_outputs(4225) <= not (a xor b);
    layer1_outputs(4226) <= not a;
    layer1_outputs(4227) <= a and b;
    layer1_outputs(4228) <= a and b;
    layer1_outputs(4229) <= a;
    layer1_outputs(4230) <= a and b;
    layer1_outputs(4231) <= not a;
    layer1_outputs(4232) <= b and not a;
    layer1_outputs(4233) <= a and not b;
    layer1_outputs(4234) <= b;
    layer1_outputs(4235) <= b;
    layer1_outputs(4236) <= b;
    layer1_outputs(4237) <= not b;
    layer1_outputs(4238) <= not a;
    layer1_outputs(4239) <= a or b;
    layer1_outputs(4240) <= b;
    layer1_outputs(4241) <= b and not a;
    layer1_outputs(4242) <= b;
    layer1_outputs(4243) <= not b or a;
    layer1_outputs(4244) <= a;
    layer1_outputs(4245) <= 1'b1;
    layer1_outputs(4246) <= not (a or b);
    layer1_outputs(4247) <= not a or b;
    layer1_outputs(4248) <= not a;
    layer1_outputs(4249) <= a xor b;
    layer1_outputs(4250) <= not (a xor b);
    layer1_outputs(4251) <= not (a xor b);
    layer1_outputs(4252) <= not a;
    layer1_outputs(4253) <= b;
    layer1_outputs(4254) <= a and b;
    layer1_outputs(4255) <= not (a xor b);
    layer1_outputs(4256) <= not (a and b);
    layer1_outputs(4257) <= not b;
    layer1_outputs(4258) <= not a or b;
    layer1_outputs(4259) <= b;
    layer1_outputs(4260) <= b and not a;
    layer1_outputs(4261) <= not (a xor b);
    layer1_outputs(4262) <= 1'b0;
    layer1_outputs(4263) <= not a;
    layer1_outputs(4264) <= a and b;
    layer1_outputs(4265) <= a and not b;
    layer1_outputs(4266) <= a xor b;
    layer1_outputs(4267) <= not a;
    layer1_outputs(4268) <= 1'b0;
    layer1_outputs(4269) <= a;
    layer1_outputs(4270) <= not (a and b);
    layer1_outputs(4271) <= not (a or b);
    layer1_outputs(4272) <= b and not a;
    layer1_outputs(4273) <= a and not b;
    layer1_outputs(4274) <= a;
    layer1_outputs(4275) <= b;
    layer1_outputs(4276) <= 1'b0;
    layer1_outputs(4277) <= not b;
    layer1_outputs(4278) <= a or b;
    layer1_outputs(4279) <= not a;
    layer1_outputs(4280) <= 1'b1;
    layer1_outputs(4281) <= b;
    layer1_outputs(4282) <= a or b;
    layer1_outputs(4283) <= 1'b1;
    layer1_outputs(4284) <= not a or b;
    layer1_outputs(4285) <= a;
    layer1_outputs(4286) <= a xor b;
    layer1_outputs(4287) <= b and not a;
    layer1_outputs(4288) <= b and not a;
    layer1_outputs(4289) <= 1'b1;
    layer1_outputs(4290) <= a and b;
    layer1_outputs(4291) <= 1'b0;
    layer1_outputs(4292) <= a;
    layer1_outputs(4293) <= not b;
    layer1_outputs(4294) <= not a;
    layer1_outputs(4295) <= not a;
    layer1_outputs(4296) <= a or b;
    layer1_outputs(4297) <= a;
    layer1_outputs(4298) <= b;
    layer1_outputs(4299) <= not (a or b);
    layer1_outputs(4300) <= not a;
    layer1_outputs(4301) <= not b;
    layer1_outputs(4302) <= not a or b;
    layer1_outputs(4303) <= not b or a;
    layer1_outputs(4304) <= not b or a;
    layer1_outputs(4305) <= not (a xor b);
    layer1_outputs(4306) <= b and not a;
    layer1_outputs(4307) <= 1'b0;
    layer1_outputs(4308) <= not a;
    layer1_outputs(4309) <= a xor b;
    layer1_outputs(4310) <= not a;
    layer1_outputs(4311) <= a xor b;
    layer1_outputs(4312) <= not b;
    layer1_outputs(4313) <= a or b;
    layer1_outputs(4314) <= a or b;
    layer1_outputs(4315) <= a;
    layer1_outputs(4316) <= a xor b;
    layer1_outputs(4317) <= a and not b;
    layer1_outputs(4318) <= a and not b;
    layer1_outputs(4319) <= not (a xor b);
    layer1_outputs(4320) <= 1'b1;
    layer1_outputs(4321) <= not b;
    layer1_outputs(4322) <= not b or a;
    layer1_outputs(4323) <= b and not a;
    layer1_outputs(4324) <= a and not b;
    layer1_outputs(4325) <= not (a or b);
    layer1_outputs(4326) <= 1'b0;
    layer1_outputs(4327) <= a and not b;
    layer1_outputs(4328) <= not (a xor b);
    layer1_outputs(4329) <= b and not a;
    layer1_outputs(4330) <= b and not a;
    layer1_outputs(4331) <= b and not a;
    layer1_outputs(4332) <= not (a and b);
    layer1_outputs(4333) <= not b;
    layer1_outputs(4334) <= not a;
    layer1_outputs(4335) <= b;
    layer1_outputs(4336) <= a xor b;
    layer1_outputs(4337) <= b;
    layer1_outputs(4338) <= not (a or b);
    layer1_outputs(4339) <= not b or a;
    layer1_outputs(4340) <= b and not a;
    layer1_outputs(4341) <= not (a or b);
    layer1_outputs(4342) <= a;
    layer1_outputs(4343) <= not (a or b);
    layer1_outputs(4344) <= not (a and b);
    layer1_outputs(4345) <= not b;
    layer1_outputs(4346) <= b;
    layer1_outputs(4347) <= a;
    layer1_outputs(4348) <= not a;
    layer1_outputs(4349) <= 1'b0;
    layer1_outputs(4350) <= b and not a;
    layer1_outputs(4351) <= b;
    layer1_outputs(4352) <= a;
    layer1_outputs(4353) <= not b;
    layer1_outputs(4354) <= a or b;
    layer1_outputs(4355) <= a;
    layer1_outputs(4356) <= a and not b;
    layer1_outputs(4357) <= a or b;
    layer1_outputs(4358) <= a and not b;
    layer1_outputs(4359) <= 1'b1;
    layer1_outputs(4360) <= b;
    layer1_outputs(4361) <= a and not b;
    layer1_outputs(4362) <= not a;
    layer1_outputs(4363) <= not b;
    layer1_outputs(4364) <= a or b;
    layer1_outputs(4365) <= a and b;
    layer1_outputs(4366) <= b;
    layer1_outputs(4367) <= b and not a;
    layer1_outputs(4368) <= a or b;
    layer1_outputs(4369) <= a or b;
    layer1_outputs(4370) <= a and b;
    layer1_outputs(4371) <= not b or a;
    layer1_outputs(4372) <= a or b;
    layer1_outputs(4373) <= not b;
    layer1_outputs(4374) <= not b;
    layer1_outputs(4375) <= not b or a;
    layer1_outputs(4376) <= a or b;
    layer1_outputs(4377) <= a and not b;
    layer1_outputs(4378) <= b;
    layer1_outputs(4379) <= a or b;
    layer1_outputs(4380) <= 1'b0;
    layer1_outputs(4381) <= not b;
    layer1_outputs(4382) <= not b or a;
    layer1_outputs(4383) <= a;
    layer1_outputs(4384) <= not a;
    layer1_outputs(4385) <= a or b;
    layer1_outputs(4386) <= b;
    layer1_outputs(4387) <= 1'b0;
    layer1_outputs(4388) <= 1'b1;
    layer1_outputs(4389) <= not a;
    layer1_outputs(4390) <= b;
    layer1_outputs(4391) <= 1'b0;
    layer1_outputs(4392) <= a or b;
    layer1_outputs(4393) <= 1'b1;
    layer1_outputs(4394) <= not b or a;
    layer1_outputs(4395) <= not b or a;
    layer1_outputs(4396) <= a or b;
    layer1_outputs(4397) <= a or b;
    layer1_outputs(4398) <= a;
    layer1_outputs(4399) <= not (a xor b);
    layer1_outputs(4400) <= not (a and b);
    layer1_outputs(4401) <= a and b;
    layer1_outputs(4402) <= not a or b;
    layer1_outputs(4403) <= a and b;
    layer1_outputs(4404) <= a or b;
    layer1_outputs(4405) <= not (a or b);
    layer1_outputs(4406) <= 1'b0;
    layer1_outputs(4407) <= 1'b0;
    layer1_outputs(4408) <= a;
    layer1_outputs(4409) <= a xor b;
    layer1_outputs(4410) <= 1'b1;
    layer1_outputs(4411) <= a xor b;
    layer1_outputs(4412) <= b and not a;
    layer1_outputs(4413) <= 1'b0;
    layer1_outputs(4414) <= a and b;
    layer1_outputs(4415) <= 1'b0;
    layer1_outputs(4416) <= not (a xor b);
    layer1_outputs(4417) <= 1'b0;
    layer1_outputs(4418) <= a;
    layer1_outputs(4419) <= 1'b0;
    layer1_outputs(4420) <= a;
    layer1_outputs(4421) <= b and not a;
    layer1_outputs(4422) <= 1'b1;
    layer1_outputs(4423) <= b and not a;
    layer1_outputs(4424) <= not b or a;
    layer1_outputs(4425) <= 1'b1;
    layer1_outputs(4426) <= not b or a;
    layer1_outputs(4427) <= not b;
    layer1_outputs(4428) <= not (a and b);
    layer1_outputs(4429) <= not b or a;
    layer1_outputs(4430) <= a or b;
    layer1_outputs(4431) <= 1'b1;
    layer1_outputs(4432) <= not (a and b);
    layer1_outputs(4433) <= not a or b;
    layer1_outputs(4434) <= b;
    layer1_outputs(4435) <= not (a and b);
    layer1_outputs(4436) <= not b or a;
    layer1_outputs(4437) <= b and not a;
    layer1_outputs(4438) <= not a;
    layer1_outputs(4439) <= b and not a;
    layer1_outputs(4440) <= not b or a;
    layer1_outputs(4441) <= a;
    layer1_outputs(4442) <= not (a or b);
    layer1_outputs(4443) <= not a or b;
    layer1_outputs(4444) <= not a or b;
    layer1_outputs(4445) <= not (a and b);
    layer1_outputs(4446) <= a;
    layer1_outputs(4447) <= not (a xor b);
    layer1_outputs(4448) <= not (a xor b);
    layer1_outputs(4449) <= not b;
    layer1_outputs(4450) <= b and not a;
    layer1_outputs(4451) <= a;
    layer1_outputs(4452) <= not b or a;
    layer1_outputs(4453) <= 1'b1;
    layer1_outputs(4454) <= a;
    layer1_outputs(4455) <= not b;
    layer1_outputs(4456) <= not a;
    layer1_outputs(4457) <= not b;
    layer1_outputs(4458) <= a and b;
    layer1_outputs(4459) <= a and not b;
    layer1_outputs(4460) <= a xor b;
    layer1_outputs(4461) <= not a;
    layer1_outputs(4462) <= a or b;
    layer1_outputs(4463) <= a and not b;
    layer1_outputs(4464) <= not (a and b);
    layer1_outputs(4465) <= not b;
    layer1_outputs(4466) <= a xor b;
    layer1_outputs(4467) <= not b;
    layer1_outputs(4468) <= not (a and b);
    layer1_outputs(4469) <= not a;
    layer1_outputs(4470) <= not b or a;
    layer1_outputs(4471) <= b;
    layer1_outputs(4472) <= not a or b;
    layer1_outputs(4473) <= a and b;
    layer1_outputs(4474) <= 1'b1;
    layer1_outputs(4475) <= not (a or b);
    layer1_outputs(4476) <= a and not b;
    layer1_outputs(4477) <= not a or b;
    layer1_outputs(4478) <= 1'b1;
    layer1_outputs(4479) <= a xor b;
    layer1_outputs(4480) <= not (a or b);
    layer1_outputs(4481) <= not b or a;
    layer1_outputs(4482) <= a;
    layer1_outputs(4483) <= a or b;
    layer1_outputs(4484) <= b;
    layer1_outputs(4485) <= a;
    layer1_outputs(4486) <= not (a and b);
    layer1_outputs(4487) <= a and not b;
    layer1_outputs(4488) <= not b or a;
    layer1_outputs(4489) <= b;
    layer1_outputs(4490) <= a xor b;
    layer1_outputs(4491) <= a and b;
    layer1_outputs(4492) <= a and b;
    layer1_outputs(4493) <= not b or a;
    layer1_outputs(4494) <= a;
    layer1_outputs(4495) <= a and not b;
    layer1_outputs(4496) <= a and not b;
    layer1_outputs(4497) <= not b or a;
    layer1_outputs(4498) <= not (a or b);
    layer1_outputs(4499) <= not b;
    layer1_outputs(4500) <= a or b;
    layer1_outputs(4501) <= not (a or b);
    layer1_outputs(4502) <= a;
    layer1_outputs(4503) <= not a;
    layer1_outputs(4504) <= not b;
    layer1_outputs(4505) <= a;
    layer1_outputs(4506) <= a or b;
    layer1_outputs(4507) <= not b or a;
    layer1_outputs(4508) <= not a;
    layer1_outputs(4509) <= not b or a;
    layer1_outputs(4510) <= a and b;
    layer1_outputs(4511) <= not a;
    layer1_outputs(4512) <= a or b;
    layer1_outputs(4513) <= a and not b;
    layer1_outputs(4514) <= not b;
    layer1_outputs(4515) <= not b;
    layer1_outputs(4516) <= a and b;
    layer1_outputs(4517) <= not b or a;
    layer1_outputs(4518) <= not (a xor b);
    layer1_outputs(4519) <= not b;
    layer1_outputs(4520) <= b;
    layer1_outputs(4521) <= b and not a;
    layer1_outputs(4522) <= a and not b;
    layer1_outputs(4523) <= b;
    layer1_outputs(4524) <= not a;
    layer1_outputs(4525) <= 1'b0;
    layer1_outputs(4526) <= b;
    layer1_outputs(4527) <= b and not a;
    layer1_outputs(4528) <= b;
    layer1_outputs(4529) <= not b;
    layer1_outputs(4530) <= not a;
    layer1_outputs(4531) <= not b;
    layer1_outputs(4532) <= a and not b;
    layer1_outputs(4533) <= b;
    layer1_outputs(4534) <= a or b;
    layer1_outputs(4535) <= not (a and b);
    layer1_outputs(4536) <= a;
    layer1_outputs(4537) <= not (a or b);
    layer1_outputs(4538) <= 1'b1;
    layer1_outputs(4539) <= not (a or b);
    layer1_outputs(4540) <= not a;
    layer1_outputs(4541) <= not b;
    layer1_outputs(4542) <= a and not b;
    layer1_outputs(4543) <= not b;
    layer1_outputs(4544) <= not (a and b);
    layer1_outputs(4545) <= b;
    layer1_outputs(4546) <= b;
    layer1_outputs(4547) <= not a;
    layer1_outputs(4548) <= a and b;
    layer1_outputs(4549) <= a and b;
    layer1_outputs(4550) <= not b;
    layer1_outputs(4551) <= 1'b0;
    layer1_outputs(4552) <= not (a xor b);
    layer1_outputs(4553) <= not (a and b);
    layer1_outputs(4554) <= not (a xor b);
    layer1_outputs(4555) <= a;
    layer1_outputs(4556) <= a and not b;
    layer1_outputs(4557) <= b;
    layer1_outputs(4558) <= 1'b0;
    layer1_outputs(4559) <= not a;
    layer1_outputs(4560) <= not a or b;
    layer1_outputs(4561) <= not a or b;
    layer1_outputs(4562) <= a and b;
    layer1_outputs(4563) <= not a;
    layer1_outputs(4564) <= b and not a;
    layer1_outputs(4565) <= b;
    layer1_outputs(4566) <= 1'b1;
    layer1_outputs(4567) <= a and b;
    layer1_outputs(4568) <= not (a or b);
    layer1_outputs(4569) <= not b;
    layer1_outputs(4570) <= a;
    layer1_outputs(4571) <= not (a and b);
    layer1_outputs(4572) <= not a;
    layer1_outputs(4573) <= 1'b0;
    layer1_outputs(4574) <= a and not b;
    layer1_outputs(4575) <= a xor b;
    layer1_outputs(4576) <= a;
    layer1_outputs(4577) <= not (a and b);
    layer1_outputs(4578) <= not b;
    layer1_outputs(4579) <= b;
    layer1_outputs(4580) <= not b;
    layer1_outputs(4581) <= 1'b1;
    layer1_outputs(4582) <= not b;
    layer1_outputs(4583) <= not a;
    layer1_outputs(4584) <= not b;
    layer1_outputs(4585) <= not a or b;
    layer1_outputs(4586) <= not a or b;
    layer1_outputs(4587) <= not a;
    layer1_outputs(4588) <= a and b;
    layer1_outputs(4589) <= 1'b0;
    layer1_outputs(4590) <= not a;
    layer1_outputs(4591) <= a;
    layer1_outputs(4592) <= not (a xor b);
    layer1_outputs(4593) <= not a;
    layer1_outputs(4594) <= a xor b;
    layer1_outputs(4595) <= b and not a;
    layer1_outputs(4596) <= not a or b;
    layer1_outputs(4597) <= b and not a;
    layer1_outputs(4598) <= not a or b;
    layer1_outputs(4599) <= a;
    layer1_outputs(4600) <= 1'b1;
    layer1_outputs(4601) <= b;
    layer1_outputs(4602) <= a xor b;
    layer1_outputs(4603) <= a and not b;
    layer1_outputs(4604) <= not a or b;
    layer1_outputs(4605) <= not b or a;
    layer1_outputs(4606) <= not a or b;
    layer1_outputs(4607) <= not (a and b);
    layer1_outputs(4608) <= a xor b;
    layer1_outputs(4609) <= not a or b;
    layer1_outputs(4610) <= a;
    layer1_outputs(4611) <= a;
    layer1_outputs(4612) <= not a or b;
    layer1_outputs(4613) <= a;
    layer1_outputs(4614) <= b;
    layer1_outputs(4615) <= 1'b1;
    layer1_outputs(4616) <= not (a or b);
    layer1_outputs(4617) <= a and b;
    layer1_outputs(4618) <= a;
    layer1_outputs(4619) <= not a;
    layer1_outputs(4620) <= b;
    layer1_outputs(4621) <= a;
    layer1_outputs(4622) <= not (a and b);
    layer1_outputs(4623) <= 1'b0;
    layer1_outputs(4624) <= b and not a;
    layer1_outputs(4625) <= a and b;
    layer1_outputs(4626) <= a;
    layer1_outputs(4627) <= a or b;
    layer1_outputs(4628) <= b;
    layer1_outputs(4629) <= 1'b1;
    layer1_outputs(4630) <= a or b;
    layer1_outputs(4631) <= not b or a;
    layer1_outputs(4632) <= not (a or b);
    layer1_outputs(4633) <= not a;
    layer1_outputs(4634) <= not a;
    layer1_outputs(4635) <= not b or a;
    layer1_outputs(4636) <= not b or a;
    layer1_outputs(4637) <= a;
    layer1_outputs(4638) <= b and not a;
    layer1_outputs(4639) <= not a or b;
    layer1_outputs(4640) <= not (a and b);
    layer1_outputs(4641) <= b;
    layer1_outputs(4642) <= not b;
    layer1_outputs(4643) <= a;
    layer1_outputs(4644) <= not b;
    layer1_outputs(4645) <= a and not b;
    layer1_outputs(4646) <= not b;
    layer1_outputs(4647) <= a;
    layer1_outputs(4648) <= a xor b;
    layer1_outputs(4649) <= a;
    layer1_outputs(4650) <= a;
    layer1_outputs(4651) <= a and not b;
    layer1_outputs(4652) <= not (a or b);
    layer1_outputs(4653) <= not (a or b);
    layer1_outputs(4654) <= b;
    layer1_outputs(4655) <= 1'b1;
    layer1_outputs(4656) <= not b or a;
    layer1_outputs(4657) <= not b;
    layer1_outputs(4658) <= a;
    layer1_outputs(4659) <= not a;
    layer1_outputs(4660) <= a and b;
    layer1_outputs(4661) <= a or b;
    layer1_outputs(4662) <= 1'b0;
    layer1_outputs(4663) <= not b;
    layer1_outputs(4664) <= not b;
    layer1_outputs(4665) <= a;
    layer1_outputs(4666) <= not a or b;
    layer1_outputs(4667) <= a and not b;
    layer1_outputs(4668) <= not b;
    layer1_outputs(4669) <= not b or a;
    layer1_outputs(4670) <= not a or b;
    layer1_outputs(4671) <= not a or b;
    layer1_outputs(4672) <= not b;
    layer1_outputs(4673) <= b;
    layer1_outputs(4674) <= a and b;
    layer1_outputs(4675) <= not b or a;
    layer1_outputs(4676) <= not (a xor b);
    layer1_outputs(4677) <= a and not b;
    layer1_outputs(4678) <= a;
    layer1_outputs(4679) <= not a;
    layer1_outputs(4680) <= a and not b;
    layer1_outputs(4681) <= b;
    layer1_outputs(4682) <= b;
    layer1_outputs(4683) <= a;
    layer1_outputs(4684) <= a;
    layer1_outputs(4685) <= not b or a;
    layer1_outputs(4686) <= 1'b1;
    layer1_outputs(4687) <= a or b;
    layer1_outputs(4688) <= not a or b;
    layer1_outputs(4689) <= a and b;
    layer1_outputs(4690) <= a and not b;
    layer1_outputs(4691) <= a and b;
    layer1_outputs(4692) <= b;
    layer1_outputs(4693) <= 1'b0;
    layer1_outputs(4694) <= not b;
    layer1_outputs(4695) <= not b;
    layer1_outputs(4696) <= b and not a;
    layer1_outputs(4697) <= not (a or b);
    layer1_outputs(4698) <= 1'b1;
    layer1_outputs(4699) <= not (a xor b);
    layer1_outputs(4700) <= a and not b;
    layer1_outputs(4701) <= not (a xor b);
    layer1_outputs(4702) <= not (a and b);
    layer1_outputs(4703) <= a and not b;
    layer1_outputs(4704) <= a;
    layer1_outputs(4705) <= not a or b;
    layer1_outputs(4706) <= a and not b;
    layer1_outputs(4707) <= 1'b0;
    layer1_outputs(4708) <= a or b;
    layer1_outputs(4709) <= b;
    layer1_outputs(4710) <= b and not a;
    layer1_outputs(4711) <= a xor b;
    layer1_outputs(4712) <= not b or a;
    layer1_outputs(4713) <= not b;
    layer1_outputs(4714) <= not b or a;
    layer1_outputs(4715) <= not (a xor b);
    layer1_outputs(4716) <= not a;
    layer1_outputs(4717) <= not b;
    layer1_outputs(4718) <= not (a or b);
    layer1_outputs(4719) <= a or b;
    layer1_outputs(4720) <= not a;
    layer1_outputs(4721) <= a and not b;
    layer1_outputs(4722) <= a and not b;
    layer1_outputs(4723) <= not (a xor b);
    layer1_outputs(4724) <= a xor b;
    layer1_outputs(4725) <= not (a and b);
    layer1_outputs(4726) <= b;
    layer1_outputs(4727) <= not a or b;
    layer1_outputs(4728) <= not b or a;
    layer1_outputs(4729) <= a and b;
    layer1_outputs(4730) <= b;
    layer1_outputs(4731) <= not (a xor b);
    layer1_outputs(4732) <= not a;
    layer1_outputs(4733) <= not (a or b);
    layer1_outputs(4734) <= a or b;
    layer1_outputs(4735) <= 1'b0;
    layer1_outputs(4736) <= a and not b;
    layer1_outputs(4737) <= a or b;
    layer1_outputs(4738) <= a and not b;
    layer1_outputs(4739) <= a xor b;
    layer1_outputs(4740) <= not (a or b);
    layer1_outputs(4741) <= b;
    layer1_outputs(4742) <= not (a or b);
    layer1_outputs(4743) <= 1'b0;
    layer1_outputs(4744) <= not b or a;
    layer1_outputs(4745) <= 1'b0;
    layer1_outputs(4746) <= not a or b;
    layer1_outputs(4747) <= not a;
    layer1_outputs(4748) <= a or b;
    layer1_outputs(4749) <= not b or a;
    layer1_outputs(4750) <= a;
    layer1_outputs(4751) <= 1'b1;
    layer1_outputs(4752) <= a or b;
    layer1_outputs(4753) <= a;
    layer1_outputs(4754) <= a and not b;
    layer1_outputs(4755) <= a and b;
    layer1_outputs(4756) <= a and not b;
    layer1_outputs(4757) <= not a;
    layer1_outputs(4758) <= not b;
    layer1_outputs(4759) <= a xor b;
    layer1_outputs(4760) <= a or b;
    layer1_outputs(4761) <= not b or a;
    layer1_outputs(4762) <= a or b;
    layer1_outputs(4763) <= not b or a;
    layer1_outputs(4764) <= not (a and b);
    layer1_outputs(4765) <= a and not b;
    layer1_outputs(4766) <= 1'b0;
    layer1_outputs(4767) <= not a or b;
    layer1_outputs(4768) <= b;
    layer1_outputs(4769) <= a and b;
    layer1_outputs(4770) <= a;
    layer1_outputs(4771) <= a and not b;
    layer1_outputs(4772) <= not b or a;
    layer1_outputs(4773) <= not a or b;
    layer1_outputs(4774) <= a and b;
    layer1_outputs(4775) <= b;
    layer1_outputs(4776) <= 1'b0;
    layer1_outputs(4777) <= a;
    layer1_outputs(4778) <= not a;
    layer1_outputs(4779) <= a;
    layer1_outputs(4780) <= not b;
    layer1_outputs(4781) <= not a;
    layer1_outputs(4782) <= a;
    layer1_outputs(4783) <= 1'b1;
    layer1_outputs(4784) <= a xor b;
    layer1_outputs(4785) <= not a;
    layer1_outputs(4786) <= a;
    layer1_outputs(4787) <= a and b;
    layer1_outputs(4788) <= a xor b;
    layer1_outputs(4789) <= not (a and b);
    layer1_outputs(4790) <= not (a and b);
    layer1_outputs(4791) <= 1'b0;
    layer1_outputs(4792) <= 1'b0;
    layer1_outputs(4793) <= not (a or b);
    layer1_outputs(4794) <= not (a xor b);
    layer1_outputs(4795) <= b;
    layer1_outputs(4796) <= not b;
    layer1_outputs(4797) <= not a or b;
    layer1_outputs(4798) <= not b or a;
    layer1_outputs(4799) <= a and not b;
    layer1_outputs(4800) <= not b;
    layer1_outputs(4801) <= a and b;
    layer1_outputs(4802) <= not a;
    layer1_outputs(4803) <= not b;
    layer1_outputs(4804) <= b;
    layer1_outputs(4805) <= not b;
    layer1_outputs(4806) <= not (a or b);
    layer1_outputs(4807) <= not a;
    layer1_outputs(4808) <= not a;
    layer1_outputs(4809) <= not a or b;
    layer1_outputs(4810) <= a and b;
    layer1_outputs(4811) <= not b or a;
    layer1_outputs(4812) <= not a or b;
    layer1_outputs(4813) <= b and not a;
    layer1_outputs(4814) <= b and not a;
    layer1_outputs(4815) <= not a;
    layer1_outputs(4816) <= not (a and b);
    layer1_outputs(4817) <= 1'b1;
    layer1_outputs(4818) <= a and not b;
    layer1_outputs(4819) <= not (a or b);
    layer1_outputs(4820) <= a or b;
    layer1_outputs(4821) <= a or b;
    layer1_outputs(4822) <= b;
    layer1_outputs(4823) <= b and not a;
    layer1_outputs(4824) <= a;
    layer1_outputs(4825) <= a;
    layer1_outputs(4826) <= b and not a;
    layer1_outputs(4827) <= b;
    layer1_outputs(4828) <= b and not a;
    layer1_outputs(4829) <= not a or b;
    layer1_outputs(4830) <= not b;
    layer1_outputs(4831) <= not (a or b);
    layer1_outputs(4832) <= b and not a;
    layer1_outputs(4833) <= a;
    layer1_outputs(4834) <= a xor b;
    layer1_outputs(4835) <= b;
    layer1_outputs(4836) <= not (a or b);
    layer1_outputs(4837) <= a;
    layer1_outputs(4838) <= not (a and b);
    layer1_outputs(4839) <= b;
    layer1_outputs(4840) <= a and b;
    layer1_outputs(4841) <= not (a and b);
    layer1_outputs(4842) <= b;
    layer1_outputs(4843) <= not b or a;
    layer1_outputs(4844) <= a xor b;
    layer1_outputs(4845) <= not b;
    layer1_outputs(4846) <= a and not b;
    layer1_outputs(4847) <= b;
    layer1_outputs(4848) <= 1'b1;
    layer1_outputs(4849) <= not a or b;
    layer1_outputs(4850) <= not (a xor b);
    layer1_outputs(4851) <= a or b;
    layer1_outputs(4852) <= not (a and b);
    layer1_outputs(4853) <= a;
    layer1_outputs(4854) <= not a or b;
    layer1_outputs(4855) <= a and b;
    layer1_outputs(4856) <= a;
    layer1_outputs(4857) <= not a or b;
    layer1_outputs(4858) <= not (a and b);
    layer1_outputs(4859) <= b;
    layer1_outputs(4860) <= b;
    layer1_outputs(4861) <= a or b;
    layer1_outputs(4862) <= b;
    layer1_outputs(4863) <= a;
    layer1_outputs(4864) <= b;
    layer1_outputs(4865) <= not a or b;
    layer1_outputs(4866) <= 1'b0;
    layer1_outputs(4867) <= not b or a;
    layer1_outputs(4868) <= not a;
    layer1_outputs(4869) <= not a;
    layer1_outputs(4870) <= a xor b;
    layer1_outputs(4871) <= a xor b;
    layer1_outputs(4872) <= a;
    layer1_outputs(4873) <= not a;
    layer1_outputs(4874) <= not (a and b);
    layer1_outputs(4875) <= not b;
    layer1_outputs(4876) <= not b;
    layer1_outputs(4877) <= not (a xor b);
    layer1_outputs(4878) <= not (a xor b);
    layer1_outputs(4879) <= a or b;
    layer1_outputs(4880) <= not b or a;
    layer1_outputs(4881) <= 1'b0;
    layer1_outputs(4882) <= not (a or b);
    layer1_outputs(4883) <= a;
    layer1_outputs(4884) <= not (a or b);
    layer1_outputs(4885) <= b and not a;
    layer1_outputs(4886) <= not a or b;
    layer1_outputs(4887) <= not (a or b);
    layer1_outputs(4888) <= a and b;
    layer1_outputs(4889) <= a and b;
    layer1_outputs(4890) <= a and b;
    layer1_outputs(4891) <= not (a xor b);
    layer1_outputs(4892) <= a and b;
    layer1_outputs(4893) <= a and not b;
    layer1_outputs(4894) <= not a or b;
    layer1_outputs(4895) <= a or b;
    layer1_outputs(4896) <= 1'b1;
    layer1_outputs(4897) <= b;
    layer1_outputs(4898) <= not (a and b);
    layer1_outputs(4899) <= a;
    layer1_outputs(4900) <= b and not a;
    layer1_outputs(4901) <= 1'b1;
    layer1_outputs(4902) <= not (a and b);
    layer1_outputs(4903) <= not (a xor b);
    layer1_outputs(4904) <= b;
    layer1_outputs(4905) <= a;
    layer1_outputs(4906) <= a or b;
    layer1_outputs(4907) <= b;
    layer1_outputs(4908) <= a;
    layer1_outputs(4909) <= a or b;
    layer1_outputs(4910) <= not b;
    layer1_outputs(4911) <= a and b;
    layer1_outputs(4912) <= b and not a;
    layer1_outputs(4913) <= a or b;
    layer1_outputs(4914) <= a and b;
    layer1_outputs(4915) <= a and b;
    layer1_outputs(4916) <= not a or b;
    layer1_outputs(4917) <= a and b;
    layer1_outputs(4918) <= a and b;
    layer1_outputs(4919) <= 1'b0;
    layer1_outputs(4920) <= a xor b;
    layer1_outputs(4921) <= a or b;
    layer1_outputs(4922) <= not (a or b);
    layer1_outputs(4923) <= a;
    layer1_outputs(4924) <= not b or a;
    layer1_outputs(4925) <= not b or a;
    layer1_outputs(4926) <= not a;
    layer1_outputs(4927) <= not b or a;
    layer1_outputs(4928) <= not a or b;
    layer1_outputs(4929) <= a;
    layer1_outputs(4930) <= not b;
    layer1_outputs(4931) <= a xor b;
    layer1_outputs(4932) <= not a or b;
    layer1_outputs(4933) <= b;
    layer1_outputs(4934) <= a;
    layer1_outputs(4935) <= b and not a;
    layer1_outputs(4936) <= a;
    layer1_outputs(4937) <= not (a or b);
    layer1_outputs(4938) <= b;
    layer1_outputs(4939) <= a xor b;
    layer1_outputs(4940) <= b;
    layer1_outputs(4941) <= not b;
    layer1_outputs(4942) <= a and not b;
    layer1_outputs(4943) <= a xor b;
    layer1_outputs(4944) <= not (a xor b);
    layer1_outputs(4945) <= not (a or b);
    layer1_outputs(4946) <= a xor b;
    layer1_outputs(4947) <= a xor b;
    layer1_outputs(4948) <= b;
    layer1_outputs(4949) <= not (a and b);
    layer1_outputs(4950) <= not a or b;
    layer1_outputs(4951) <= a;
    layer1_outputs(4952) <= b;
    layer1_outputs(4953) <= not b or a;
    layer1_outputs(4954) <= not b;
    layer1_outputs(4955) <= not a;
    layer1_outputs(4956) <= not a or b;
    layer1_outputs(4957) <= not (a and b);
    layer1_outputs(4958) <= 1'b0;
    layer1_outputs(4959) <= a;
    layer1_outputs(4960) <= not a;
    layer1_outputs(4961) <= not (a and b);
    layer1_outputs(4962) <= not (a or b);
    layer1_outputs(4963) <= b and not a;
    layer1_outputs(4964) <= a and not b;
    layer1_outputs(4965) <= a or b;
    layer1_outputs(4966) <= not (a or b);
    layer1_outputs(4967) <= a xor b;
    layer1_outputs(4968) <= not (a or b);
    layer1_outputs(4969) <= not b;
    layer1_outputs(4970) <= not b or a;
    layer1_outputs(4971) <= a;
    layer1_outputs(4972) <= a;
    layer1_outputs(4973) <= not b or a;
    layer1_outputs(4974) <= b and not a;
    layer1_outputs(4975) <= a;
    layer1_outputs(4976) <= not a or b;
    layer1_outputs(4977) <= a or b;
    layer1_outputs(4978) <= not a;
    layer1_outputs(4979) <= not (a and b);
    layer1_outputs(4980) <= not (a xor b);
    layer1_outputs(4981) <= a;
    layer1_outputs(4982) <= a and b;
    layer1_outputs(4983) <= not b or a;
    layer1_outputs(4984) <= a or b;
    layer1_outputs(4985) <= not a;
    layer1_outputs(4986) <= not (a and b);
    layer1_outputs(4987) <= a and not b;
    layer1_outputs(4988) <= a;
    layer1_outputs(4989) <= not b;
    layer1_outputs(4990) <= a and not b;
    layer1_outputs(4991) <= not a or b;
    layer1_outputs(4992) <= not b;
    layer1_outputs(4993) <= not a;
    layer1_outputs(4994) <= not b;
    layer1_outputs(4995) <= b and not a;
    layer1_outputs(4996) <= not b or a;
    layer1_outputs(4997) <= not (a or b);
    layer1_outputs(4998) <= not a;
    layer1_outputs(4999) <= b;
    layer1_outputs(5000) <= not (a or b);
    layer1_outputs(5001) <= a or b;
    layer1_outputs(5002) <= a;
    layer1_outputs(5003) <= not b or a;
    layer1_outputs(5004) <= not a or b;
    layer1_outputs(5005) <= 1'b1;
    layer1_outputs(5006) <= a;
    layer1_outputs(5007) <= b;
    layer1_outputs(5008) <= not b or a;
    layer1_outputs(5009) <= not b;
    layer1_outputs(5010) <= a;
    layer1_outputs(5011) <= a and b;
    layer1_outputs(5012) <= b;
    layer1_outputs(5013) <= not (a and b);
    layer1_outputs(5014) <= a xor b;
    layer1_outputs(5015) <= b and not a;
    layer1_outputs(5016) <= b and not a;
    layer1_outputs(5017) <= a;
    layer1_outputs(5018) <= 1'b0;
    layer1_outputs(5019) <= not a;
    layer1_outputs(5020) <= b and not a;
    layer1_outputs(5021) <= a or b;
    layer1_outputs(5022) <= a;
    layer1_outputs(5023) <= a and b;
    layer1_outputs(5024) <= not b or a;
    layer1_outputs(5025) <= a and not b;
    layer1_outputs(5026) <= a;
    layer1_outputs(5027) <= 1'b0;
    layer1_outputs(5028) <= b;
    layer1_outputs(5029) <= not a;
    layer1_outputs(5030) <= not b;
    layer1_outputs(5031) <= a and b;
    layer1_outputs(5032) <= not a;
    layer1_outputs(5033) <= not a;
    layer1_outputs(5034) <= not a;
    layer1_outputs(5035) <= not a or b;
    layer1_outputs(5036) <= b;
    layer1_outputs(5037) <= a and b;
    layer1_outputs(5038) <= a and not b;
    layer1_outputs(5039) <= not (a and b);
    layer1_outputs(5040) <= not a;
    layer1_outputs(5041) <= a and b;
    layer1_outputs(5042) <= 1'b1;
    layer1_outputs(5043) <= not a;
    layer1_outputs(5044) <= not (a or b);
    layer1_outputs(5045) <= not (a or b);
    layer1_outputs(5046) <= a;
    layer1_outputs(5047) <= a;
    layer1_outputs(5048) <= not (a xor b);
    layer1_outputs(5049) <= not b or a;
    layer1_outputs(5050) <= not b or a;
    layer1_outputs(5051) <= b;
    layer1_outputs(5052) <= b;
    layer1_outputs(5053) <= not (a or b);
    layer1_outputs(5054) <= not b;
    layer1_outputs(5055) <= 1'b0;
    layer1_outputs(5056) <= not a;
    layer1_outputs(5057) <= not a;
    layer1_outputs(5058) <= b;
    layer1_outputs(5059) <= not (a or b);
    layer1_outputs(5060) <= b;
    layer1_outputs(5061) <= not a;
    layer1_outputs(5062) <= not b;
    layer1_outputs(5063) <= a and b;
    layer1_outputs(5064) <= b;
    layer1_outputs(5065) <= not (a or b);
    layer1_outputs(5066) <= not (a and b);
    layer1_outputs(5067) <= not (a xor b);
    layer1_outputs(5068) <= a xor b;
    layer1_outputs(5069) <= a or b;
    layer1_outputs(5070) <= not (a and b);
    layer1_outputs(5071) <= not a;
    layer1_outputs(5072) <= not a;
    layer1_outputs(5073) <= a or b;
    layer1_outputs(5074) <= a xor b;
    layer1_outputs(5075) <= not (a xor b);
    layer1_outputs(5076) <= not a;
    layer1_outputs(5077) <= not a or b;
    layer1_outputs(5078) <= not a;
    layer1_outputs(5079) <= a xor b;
    layer1_outputs(5080) <= not a or b;
    layer1_outputs(5081) <= b;
    layer1_outputs(5082) <= a and b;
    layer1_outputs(5083) <= b;
    layer1_outputs(5084) <= not b;
    layer1_outputs(5085) <= not (a or b);
    layer1_outputs(5086) <= a and b;
    layer1_outputs(5087) <= a;
    layer1_outputs(5088) <= not b;
    layer1_outputs(5089) <= not a or b;
    layer1_outputs(5090) <= not (a and b);
    layer1_outputs(5091) <= not a or b;
    layer1_outputs(5092) <= b;
    layer1_outputs(5093) <= not a or b;
    layer1_outputs(5094) <= a or b;
    layer1_outputs(5095) <= not a or b;
    layer1_outputs(5096) <= a;
    layer1_outputs(5097) <= a or b;
    layer1_outputs(5098) <= not b;
    layer1_outputs(5099) <= not a or b;
    layer1_outputs(5100) <= not (a or b);
    layer1_outputs(5101) <= a or b;
    layer1_outputs(5102) <= not (a or b);
    layer1_outputs(5103) <= not (a and b);
    layer1_outputs(5104) <= not b or a;
    layer1_outputs(5105) <= not (a and b);
    layer1_outputs(5106) <= 1'b1;
    layer1_outputs(5107) <= a xor b;
    layer1_outputs(5108) <= not b;
    layer1_outputs(5109) <= not b or a;
    layer1_outputs(5110) <= b and not a;
    layer1_outputs(5111) <= a;
    layer1_outputs(5112) <= not a or b;
    layer1_outputs(5113) <= a and b;
    layer1_outputs(5114) <= not (a and b);
    layer1_outputs(5115) <= not (a and b);
    layer1_outputs(5116) <= not b or a;
    layer1_outputs(5117) <= not (a and b);
    layer1_outputs(5118) <= a and b;
    layer1_outputs(5119) <= b and not a;
    layer1_outputs(5120) <= not a or b;
    layer1_outputs(5121) <= not a or b;
    layer1_outputs(5122) <= not a;
    layer1_outputs(5123) <= not a;
    layer1_outputs(5124) <= 1'b0;
    layer1_outputs(5125) <= not a;
    layer1_outputs(5126) <= not b or a;
    layer1_outputs(5127) <= b and not a;
    layer1_outputs(5128) <= b and not a;
    layer1_outputs(5129) <= not b;
    layer1_outputs(5130) <= a;
    layer1_outputs(5131) <= not a or b;
    layer1_outputs(5132) <= b;
    layer1_outputs(5133) <= a and b;
    layer1_outputs(5134) <= not (a and b);
    layer1_outputs(5135) <= a;
    layer1_outputs(5136) <= not (a xor b);
    layer1_outputs(5137) <= a and b;
    layer1_outputs(5138) <= not b;
    layer1_outputs(5139) <= a and not b;
    layer1_outputs(5140) <= not a;
    layer1_outputs(5141) <= not a or b;
    layer1_outputs(5142) <= not b or a;
    layer1_outputs(5143) <= a xor b;
    layer1_outputs(5144) <= not b;
    layer1_outputs(5145) <= not (a xor b);
    layer1_outputs(5146) <= b;
    layer1_outputs(5147) <= a;
    layer1_outputs(5148) <= not a;
    layer1_outputs(5149) <= not (a xor b);
    layer1_outputs(5150) <= a or b;
    layer1_outputs(5151) <= not b;
    layer1_outputs(5152) <= not a or b;
    layer1_outputs(5153) <= not a or b;
    layer1_outputs(5154) <= a xor b;
    layer1_outputs(5155) <= not (a and b);
    layer1_outputs(5156) <= b;
    layer1_outputs(5157) <= not b;
    layer1_outputs(5158) <= not b;
    layer1_outputs(5159) <= a xor b;
    layer1_outputs(5160) <= a and b;
    layer1_outputs(5161) <= a or b;
    layer1_outputs(5162) <= a;
    layer1_outputs(5163) <= not (a or b);
    layer1_outputs(5164) <= not (a xor b);
    layer1_outputs(5165) <= not b;
    layer1_outputs(5166) <= not (a or b);
    layer1_outputs(5167) <= a or b;
    layer1_outputs(5168) <= a;
    layer1_outputs(5169) <= a and b;
    layer1_outputs(5170) <= a or b;
    layer1_outputs(5171) <= not (a and b);
    layer1_outputs(5172) <= a and not b;
    layer1_outputs(5173) <= not b or a;
    layer1_outputs(5174) <= b and not a;
    layer1_outputs(5175) <= b and not a;
    layer1_outputs(5176) <= 1'b1;
    layer1_outputs(5177) <= a;
    layer1_outputs(5178) <= not b or a;
    layer1_outputs(5179) <= not (a or b);
    layer1_outputs(5180) <= a and b;
    layer1_outputs(5181) <= not (a or b);
    layer1_outputs(5182) <= b and not a;
    layer1_outputs(5183) <= a or b;
    layer1_outputs(5184) <= not a or b;
    layer1_outputs(5185) <= 1'b0;
    layer1_outputs(5186) <= not (a or b);
    layer1_outputs(5187) <= b;
    layer1_outputs(5188) <= not a or b;
    layer1_outputs(5189) <= a;
    layer1_outputs(5190) <= not a or b;
    layer1_outputs(5191) <= not (a and b);
    layer1_outputs(5192) <= a or b;
    layer1_outputs(5193) <= not a;
    layer1_outputs(5194) <= not b;
    layer1_outputs(5195) <= 1'b1;
    layer1_outputs(5196) <= 1'b0;
    layer1_outputs(5197) <= a;
    layer1_outputs(5198) <= b;
    layer1_outputs(5199) <= not (a or b);
    layer1_outputs(5200) <= a;
    layer1_outputs(5201) <= a xor b;
    layer1_outputs(5202) <= not a;
    layer1_outputs(5203) <= not a or b;
    layer1_outputs(5204) <= not (a and b);
    layer1_outputs(5205) <= not a;
    layer1_outputs(5206) <= not (a or b);
    layer1_outputs(5207) <= not b;
    layer1_outputs(5208) <= not (a xor b);
    layer1_outputs(5209) <= not (a and b);
    layer1_outputs(5210) <= a xor b;
    layer1_outputs(5211) <= not a or b;
    layer1_outputs(5212) <= a and b;
    layer1_outputs(5213) <= a;
    layer1_outputs(5214) <= not b;
    layer1_outputs(5215) <= not (a and b);
    layer1_outputs(5216) <= not (a and b);
    layer1_outputs(5217) <= not a or b;
    layer1_outputs(5218) <= not a or b;
    layer1_outputs(5219) <= a and not b;
    layer1_outputs(5220) <= a and b;
    layer1_outputs(5221) <= 1'b0;
    layer1_outputs(5222) <= not a or b;
    layer1_outputs(5223) <= not a;
    layer1_outputs(5224) <= not b;
    layer1_outputs(5225) <= b;
    layer1_outputs(5226) <= b;
    layer1_outputs(5227) <= not a;
    layer1_outputs(5228) <= not b;
    layer1_outputs(5229) <= not b;
    layer1_outputs(5230) <= a and b;
    layer1_outputs(5231) <= a xor b;
    layer1_outputs(5232) <= 1'b0;
    layer1_outputs(5233) <= not (a and b);
    layer1_outputs(5234) <= a;
    layer1_outputs(5235) <= not a or b;
    layer1_outputs(5236) <= a xor b;
    layer1_outputs(5237) <= a;
    layer1_outputs(5238) <= b;
    layer1_outputs(5239) <= not (a and b);
    layer1_outputs(5240) <= b;
    layer1_outputs(5241) <= a or b;
    layer1_outputs(5242) <= 1'b0;
    layer1_outputs(5243) <= not b;
    layer1_outputs(5244) <= a and b;
    layer1_outputs(5245) <= a or b;
    layer1_outputs(5246) <= a or b;
    layer1_outputs(5247) <= a or b;
    layer1_outputs(5248) <= a;
    layer1_outputs(5249) <= a and b;
    layer1_outputs(5250) <= not a;
    layer1_outputs(5251) <= a and not b;
    layer1_outputs(5252) <= not b;
    layer1_outputs(5253) <= not b;
    layer1_outputs(5254) <= b and not a;
    layer1_outputs(5255) <= not b or a;
    layer1_outputs(5256) <= a and not b;
    layer1_outputs(5257) <= a or b;
    layer1_outputs(5258) <= a;
    layer1_outputs(5259) <= b;
    layer1_outputs(5260) <= 1'b0;
    layer1_outputs(5261) <= 1'b0;
    layer1_outputs(5262) <= not (a and b);
    layer1_outputs(5263) <= a and not b;
    layer1_outputs(5264) <= not a or b;
    layer1_outputs(5265) <= not a or b;
    layer1_outputs(5266) <= a or b;
    layer1_outputs(5267) <= a;
    layer1_outputs(5268) <= not a or b;
    layer1_outputs(5269) <= 1'b1;
    layer1_outputs(5270) <= not a or b;
    layer1_outputs(5271) <= a;
    layer1_outputs(5272) <= not (a xor b);
    layer1_outputs(5273) <= not a;
    layer1_outputs(5274) <= b;
    layer1_outputs(5275) <= a;
    layer1_outputs(5276) <= not a;
    layer1_outputs(5277) <= a xor b;
    layer1_outputs(5278) <= not a;
    layer1_outputs(5279) <= not b;
    layer1_outputs(5280) <= a;
    layer1_outputs(5281) <= not (a or b);
    layer1_outputs(5282) <= a or b;
    layer1_outputs(5283) <= not b or a;
    layer1_outputs(5284) <= not a;
    layer1_outputs(5285) <= b;
    layer1_outputs(5286) <= a and b;
    layer1_outputs(5287) <= b;
    layer1_outputs(5288) <= a;
    layer1_outputs(5289) <= a and b;
    layer1_outputs(5290) <= a and not b;
    layer1_outputs(5291) <= a or b;
    layer1_outputs(5292) <= not a;
    layer1_outputs(5293) <= not a or b;
    layer1_outputs(5294) <= not a;
    layer1_outputs(5295) <= not (a xor b);
    layer1_outputs(5296) <= 1'b0;
    layer1_outputs(5297) <= not b;
    layer1_outputs(5298) <= a;
    layer1_outputs(5299) <= not (a or b);
    layer1_outputs(5300) <= not (a or b);
    layer1_outputs(5301) <= not (a or b);
    layer1_outputs(5302) <= b and not a;
    layer1_outputs(5303) <= b and not a;
    layer1_outputs(5304) <= not a or b;
    layer1_outputs(5305) <= a;
    layer1_outputs(5306) <= a;
    layer1_outputs(5307) <= b;
    layer1_outputs(5308) <= a;
    layer1_outputs(5309) <= a and b;
    layer1_outputs(5310) <= not b;
    layer1_outputs(5311) <= not a or b;
    layer1_outputs(5312) <= not a;
    layer1_outputs(5313) <= b;
    layer1_outputs(5314) <= not a or b;
    layer1_outputs(5315) <= a;
    layer1_outputs(5316) <= b and not a;
    layer1_outputs(5317) <= b and not a;
    layer1_outputs(5318) <= b and not a;
    layer1_outputs(5319) <= not b;
    layer1_outputs(5320) <= 1'b1;
    layer1_outputs(5321) <= not a or b;
    layer1_outputs(5322) <= not b;
    layer1_outputs(5323) <= not (a and b);
    layer1_outputs(5324) <= a xor b;
    layer1_outputs(5325) <= not (a or b);
    layer1_outputs(5326) <= b;
    layer1_outputs(5327) <= not b or a;
    layer1_outputs(5328) <= not a;
    layer1_outputs(5329) <= not b;
    layer1_outputs(5330) <= a and b;
    layer1_outputs(5331) <= a or b;
    layer1_outputs(5332) <= a or b;
    layer1_outputs(5333) <= a and b;
    layer1_outputs(5334) <= b;
    layer1_outputs(5335) <= not a;
    layer1_outputs(5336) <= not (a and b);
    layer1_outputs(5337) <= a xor b;
    layer1_outputs(5338) <= a and b;
    layer1_outputs(5339) <= a and b;
    layer1_outputs(5340) <= not b or a;
    layer1_outputs(5341) <= a and b;
    layer1_outputs(5342) <= not a;
    layer1_outputs(5343) <= not a;
    layer1_outputs(5344) <= a and b;
    layer1_outputs(5345) <= 1'b0;
    layer1_outputs(5346) <= 1'b0;
    layer1_outputs(5347) <= not b;
    layer1_outputs(5348) <= a xor b;
    layer1_outputs(5349) <= a and not b;
    layer1_outputs(5350) <= not a;
    layer1_outputs(5351) <= not (a xor b);
    layer1_outputs(5352) <= a;
    layer1_outputs(5353) <= not (a or b);
    layer1_outputs(5354) <= not b;
    layer1_outputs(5355) <= a and not b;
    layer1_outputs(5356) <= not b;
    layer1_outputs(5357) <= not (a or b);
    layer1_outputs(5358) <= b;
    layer1_outputs(5359) <= not b;
    layer1_outputs(5360) <= b and not a;
    layer1_outputs(5361) <= a and not b;
    layer1_outputs(5362) <= b;
    layer1_outputs(5363) <= not (a or b);
    layer1_outputs(5364) <= not b;
    layer1_outputs(5365) <= 1'b1;
    layer1_outputs(5366) <= a;
    layer1_outputs(5367) <= a and not b;
    layer1_outputs(5368) <= 1'b1;
    layer1_outputs(5369) <= a and not b;
    layer1_outputs(5370) <= a and not b;
    layer1_outputs(5371) <= b and not a;
    layer1_outputs(5372) <= b and not a;
    layer1_outputs(5373) <= not (a and b);
    layer1_outputs(5374) <= not (a xor b);
    layer1_outputs(5375) <= not (a xor b);
    layer1_outputs(5376) <= a and b;
    layer1_outputs(5377) <= not a;
    layer1_outputs(5378) <= not a;
    layer1_outputs(5379) <= b;
    layer1_outputs(5380) <= not a or b;
    layer1_outputs(5381) <= not a or b;
    layer1_outputs(5382) <= not a or b;
    layer1_outputs(5383) <= not (a and b);
    layer1_outputs(5384) <= not b or a;
    layer1_outputs(5385) <= a or b;
    layer1_outputs(5386) <= a or b;
    layer1_outputs(5387) <= a xor b;
    layer1_outputs(5388) <= a and b;
    layer1_outputs(5389) <= not b or a;
    layer1_outputs(5390) <= not b or a;
    layer1_outputs(5391) <= not a or b;
    layer1_outputs(5392) <= b;
    layer1_outputs(5393) <= a;
    layer1_outputs(5394) <= a and not b;
    layer1_outputs(5395) <= not b;
    layer1_outputs(5396) <= a or b;
    layer1_outputs(5397) <= a and not b;
    layer1_outputs(5398) <= a xor b;
    layer1_outputs(5399) <= a;
    layer1_outputs(5400) <= b;
    layer1_outputs(5401) <= not (a xor b);
    layer1_outputs(5402) <= a or b;
    layer1_outputs(5403) <= not a;
    layer1_outputs(5404) <= a;
    layer1_outputs(5405) <= not b;
    layer1_outputs(5406) <= b;
    layer1_outputs(5407) <= not (a or b);
    layer1_outputs(5408) <= 1'b1;
    layer1_outputs(5409) <= not a or b;
    layer1_outputs(5410) <= a;
    layer1_outputs(5411) <= b;
    layer1_outputs(5412) <= 1'b1;
    layer1_outputs(5413) <= not b;
    layer1_outputs(5414) <= not a;
    layer1_outputs(5415) <= a or b;
    layer1_outputs(5416) <= a;
    layer1_outputs(5417) <= not (a and b);
    layer1_outputs(5418) <= 1'b0;
    layer1_outputs(5419) <= b;
    layer1_outputs(5420) <= a xor b;
    layer1_outputs(5421) <= a and not b;
    layer1_outputs(5422) <= not b;
    layer1_outputs(5423) <= not b or a;
    layer1_outputs(5424) <= not (a and b);
    layer1_outputs(5425) <= not (a xor b);
    layer1_outputs(5426) <= a;
    layer1_outputs(5427) <= 1'b1;
    layer1_outputs(5428) <= b;
    layer1_outputs(5429) <= not (a xor b);
    layer1_outputs(5430) <= 1'b0;
    layer1_outputs(5431) <= not (a and b);
    layer1_outputs(5432) <= not a;
    layer1_outputs(5433) <= a and not b;
    layer1_outputs(5434) <= a;
    layer1_outputs(5435) <= a and not b;
    layer1_outputs(5436) <= a xor b;
    layer1_outputs(5437) <= 1'b0;
    layer1_outputs(5438) <= b;
    layer1_outputs(5439) <= a and not b;
    layer1_outputs(5440) <= a and b;
    layer1_outputs(5441) <= b and not a;
    layer1_outputs(5442) <= 1'b0;
    layer1_outputs(5443) <= 1'b0;
    layer1_outputs(5444) <= b;
    layer1_outputs(5445) <= not b;
    layer1_outputs(5446) <= not b;
    layer1_outputs(5447) <= not (a and b);
    layer1_outputs(5448) <= b;
    layer1_outputs(5449) <= not (a or b);
    layer1_outputs(5450) <= a and not b;
    layer1_outputs(5451) <= not a or b;
    layer1_outputs(5452) <= b and not a;
    layer1_outputs(5453) <= a and not b;
    layer1_outputs(5454) <= not a;
    layer1_outputs(5455) <= b;
    layer1_outputs(5456) <= b;
    layer1_outputs(5457) <= not a or b;
    layer1_outputs(5458) <= not (a or b);
    layer1_outputs(5459) <= not (a and b);
    layer1_outputs(5460) <= not (a xor b);
    layer1_outputs(5461) <= a xor b;
    layer1_outputs(5462) <= not (a xor b);
    layer1_outputs(5463) <= b and not a;
    layer1_outputs(5464) <= a;
    layer1_outputs(5465) <= a xor b;
    layer1_outputs(5466) <= not a or b;
    layer1_outputs(5467) <= a xor b;
    layer1_outputs(5468) <= b and not a;
    layer1_outputs(5469) <= a or b;
    layer1_outputs(5470) <= not (a or b);
    layer1_outputs(5471) <= not a or b;
    layer1_outputs(5472) <= b;
    layer1_outputs(5473) <= not (a and b);
    layer1_outputs(5474) <= not a or b;
    layer1_outputs(5475) <= not b;
    layer1_outputs(5476) <= a or b;
    layer1_outputs(5477) <= not b or a;
    layer1_outputs(5478) <= not a or b;
    layer1_outputs(5479) <= a or b;
    layer1_outputs(5480) <= 1'b1;
    layer1_outputs(5481) <= a xor b;
    layer1_outputs(5482) <= 1'b0;
    layer1_outputs(5483) <= not (a and b);
    layer1_outputs(5484) <= a and not b;
    layer1_outputs(5485) <= not a;
    layer1_outputs(5486) <= not (a xor b);
    layer1_outputs(5487) <= b and not a;
    layer1_outputs(5488) <= not a or b;
    layer1_outputs(5489) <= not a;
    layer1_outputs(5490) <= 1'b1;
    layer1_outputs(5491) <= b;
    layer1_outputs(5492) <= b;
    layer1_outputs(5493) <= a xor b;
    layer1_outputs(5494) <= not a or b;
    layer1_outputs(5495) <= b and not a;
    layer1_outputs(5496) <= not a or b;
    layer1_outputs(5497) <= b and not a;
    layer1_outputs(5498) <= not (a or b);
    layer1_outputs(5499) <= b;
    layer1_outputs(5500) <= a or b;
    layer1_outputs(5501) <= not (a or b);
    layer1_outputs(5502) <= not a or b;
    layer1_outputs(5503) <= not a or b;
    layer1_outputs(5504) <= not (a or b);
    layer1_outputs(5505) <= not a;
    layer1_outputs(5506) <= not b;
    layer1_outputs(5507) <= a;
    layer1_outputs(5508) <= 1'b0;
    layer1_outputs(5509) <= not b or a;
    layer1_outputs(5510) <= b;
    layer1_outputs(5511) <= a;
    layer1_outputs(5512) <= not a or b;
    layer1_outputs(5513) <= b;
    layer1_outputs(5514) <= a;
    layer1_outputs(5515) <= b and not a;
    layer1_outputs(5516) <= b;
    layer1_outputs(5517) <= a and b;
    layer1_outputs(5518) <= a or b;
    layer1_outputs(5519) <= not b or a;
    layer1_outputs(5520) <= 1'b1;
    layer1_outputs(5521) <= a and not b;
    layer1_outputs(5522) <= 1'b0;
    layer1_outputs(5523) <= not b;
    layer1_outputs(5524) <= a or b;
    layer1_outputs(5525) <= not a;
    layer1_outputs(5526) <= not (a or b);
    layer1_outputs(5527) <= not a or b;
    layer1_outputs(5528) <= not a;
    layer1_outputs(5529) <= a xor b;
    layer1_outputs(5530) <= a;
    layer1_outputs(5531) <= b and not a;
    layer1_outputs(5532) <= not (a xor b);
    layer1_outputs(5533) <= not (a xor b);
    layer1_outputs(5534) <= not a;
    layer1_outputs(5535) <= not b or a;
    layer1_outputs(5536) <= b and not a;
    layer1_outputs(5537) <= b and not a;
    layer1_outputs(5538) <= not a or b;
    layer1_outputs(5539) <= not a;
    layer1_outputs(5540) <= not (a or b);
    layer1_outputs(5541) <= not (a and b);
    layer1_outputs(5542) <= a xor b;
    layer1_outputs(5543) <= a and b;
    layer1_outputs(5544) <= a;
    layer1_outputs(5545) <= not (a and b);
    layer1_outputs(5546) <= a and b;
    layer1_outputs(5547) <= b and not a;
    layer1_outputs(5548) <= not a or b;
    layer1_outputs(5549) <= a and not b;
    layer1_outputs(5550) <= not b or a;
    layer1_outputs(5551) <= not a;
    layer1_outputs(5552) <= not b or a;
    layer1_outputs(5553) <= a or b;
    layer1_outputs(5554) <= not (a and b);
    layer1_outputs(5555) <= b and not a;
    layer1_outputs(5556) <= not b;
    layer1_outputs(5557) <= a or b;
    layer1_outputs(5558) <= a and not b;
    layer1_outputs(5559) <= b;
    layer1_outputs(5560) <= a xor b;
    layer1_outputs(5561) <= a and not b;
    layer1_outputs(5562) <= not (a or b);
    layer1_outputs(5563) <= a or b;
    layer1_outputs(5564) <= a;
    layer1_outputs(5565) <= not b or a;
    layer1_outputs(5566) <= a or b;
    layer1_outputs(5567) <= a and b;
    layer1_outputs(5568) <= not a;
    layer1_outputs(5569) <= a or b;
    layer1_outputs(5570) <= not b;
    layer1_outputs(5571) <= a and b;
    layer1_outputs(5572) <= not a;
    layer1_outputs(5573) <= not (a and b);
    layer1_outputs(5574) <= not (a and b);
    layer1_outputs(5575) <= a and b;
    layer1_outputs(5576) <= a xor b;
    layer1_outputs(5577) <= a and b;
    layer1_outputs(5578) <= a xor b;
    layer1_outputs(5579) <= not b;
    layer1_outputs(5580) <= not b;
    layer1_outputs(5581) <= 1'b1;
    layer1_outputs(5582) <= b and not a;
    layer1_outputs(5583) <= a or b;
    layer1_outputs(5584) <= a and not b;
    layer1_outputs(5585) <= not a;
    layer1_outputs(5586) <= a;
    layer1_outputs(5587) <= a;
    layer1_outputs(5588) <= b;
    layer1_outputs(5589) <= not b;
    layer1_outputs(5590) <= b;
    layer1_outputs(5591) <= a and not b;
    layer1_outputs(5592) <= b and not a;
    layer1_outputs(5593) <= a and not b;
    layer1_outputs(5594) <= a and b;
    layer1_outputs(5595) <= a or b;
    layer1_outputs(5596) <= a and not b;
    layer1_outputs(5597) <= a and b;
    layer1_outputs(5598) <= b and not a;
    layer1_outputs(5599) <= not a;
    layer1_outputs(5600) <= not a;
    layer1_outputs(5601) <= a;
    layer1_outputs(5602) <= a or b;
    layer1_outputs(5603) <= not b;
    layer1_outputs(5604) <= not b;
    layer1_outputs(5605) <= b and not a;
    layer1_outputs(5606) <= 1'b1;
    layer1_outputs(5607) <= not b;
    layer1_outputs(5608) <= a or b;
    layer1_outputs(5609) <= a or b;
    layer1_outputs(5610) <= not (a xor b);
    layer1_outputs(5611) <= b;
    layer1_outputs(5612) <= not a;
    layer1_outputs(5613) <= 1'b0;
    layer1_outputs(5614) <= not a or b;
    layer1_outputs(5615) <= a;
    layer1_outputs(5616) <= not (a or b);
    layer1_outputs(5617) <= not (a and b);
    layer1_outputs(5618) <= a and b;
    layer1_outputs(5619) <= not (a xor b);
    layer1_outputs(5620) <= not a;
    layer1_outputs(5621) <= b;
    layer1_outputs(5622) <= a and not b;
    layer1_outputs(5623) <= a;
    layer1_outputs(5624) <= not b or a;
    layer1_outputs(5625) <= 1'b1;
    layer1_outputs(5626) <= not b or a;
    layer1_outputs(5627) <= a and not b;
    layer1_outputs(5628) <= a;
    layer1_outputs(5629) <= a xor b;
    layer1_outputs(5630) <= not b;
    layer1_outputs(5631) <= not b or a;
    layer1_outputs(5632) <= b and not a;
    layer1_outputs(5633) <= a xor b;
    layer1_outputs(5634) <= not a or b;
    layer1_outputs(5635) <= b;
    layer1_outputs(5636) <= a and b;
    layer1_outputs(5637) <= not (a or b);
    layer1_outputs(5638) <= a and b;
    layer1_outputs(5639) <= not b;
    layer1_outputs(5640) <= b and not a;
    layer1_outputs(5641) <= not (a or b);
    layer1_outputs(5642) <= not b or a;
    layer1_outputs(5643) <= not b;
    layer1_outputs(5644) <= a and b;
    layer1_outputs(5645) <= b;
    layer1_outputs(5646) <= a xor b;
    layer1_outputs(5647) <= not a;
    layer1_outputs(5648) <= 1'b0;
    layer1_outputs(5649) <= a xor b;
    layer1_outputs(5650) <= not (a and b);
    layer1_outputs(5651) <= not a or b;
    layer1_outputs(5652) <= not (a xor b);
    layer1_outputs(5653) <= a;
    layer1_outputs(5654) <= b;
    layer1_outputs(5655) <= a and b;
    layer1_outputs(5656) <= 1'b1;
    layer1_outputs(5657) <= a;
    layer1_outputs(5658) <= 1'b0;
    layer1_outputs(5659) <= 1'b1;
    layer1_outputs(5660) <= b;
    layer1_outputs(5661) <= a xor b;
    layer1_outputs(5662) <= not b or a;
    layer1_outputs(5663) <= b and not a;
    layer1_outputs(5664) <= not b or a;
    layer1_outputs(5665) <= not b or a;
    layer1_outputs(5666) <= a or b;
    layer1_outputs(5667) <= a;
    layer1_outputs(5668) <= not a;
    layer1_outputs(5669) <= not (a or b);
    layer1_outputs(5670) <= b;
    layer1_outputs(5671) <= 1'b0;
    layer1_outputs(5672) <= a and not b;
    layer1_outputs(5673) <= not b;
    layer1_outputs(5674) <= not a or b;
    layer1_outputs(5675) <= a and not b;
    layer1_outputs(5676) <= a and not b;
    layer1_outputs(5677) <= a or b;
    layer1_outputs(5678) <= not a;
    layer1_outputs(5679) <= not (a xor b);
    layer1_outputs(5680) <= a and b;
    layer1_outputs(5681) <= b;
    layer1_outputs(5682) <= not (a or b);
    layer1_outputs(5683) <= a or b;
    layer1_outputs(5684) <= a xor b;
    layer1_outputs(5685) <= a and b;
    layer1_outputs(5686) <= not b;
    layer1_outputs(5687) <= 1'b1;
    layer1_outputs(5688) <= not b;
    layer1_outputs(5689) <= not (a or b);
    layer1_outputs(5690) <= b;
    layer1_outputs(5691) <= not (a xor b);
    layer1_outputs(5692) <= not a;
    layer1_outputs(5693) <= not a or b;
    layer1_outputs(5694) <= not (a xor b);
    layer1_outputs(5695) <= not b;
    layer1_outputs(5696) <= a xor b;
    layer1_outputs(5697) <= b;
    layer1_outputs(5698) <= a and b;
    layer1_outputs(5699) <= 1'b1;
    layer1_outputs(5700) <= not a;
    layer1_outputs(5701) <= not a;
    layer1_outputs(5702) <= not b;
    layer1_outputs(5703) <= not a;
    layer1_outputs(5704) <= a;
    layer1_outputs(5705) <= a;
    layer1_outputs(5706) <= a and b;
    layer1_outputs(5707) <= not (a xor b);
    layer1_outputs(5708) <= a or b;
    layer1_outputs(5709) <= b;
    layer1_outputs(5710) <= a and b;
    layer1_outputs(5711) <= a and not b;
    layer1_outputs(5712) <= a xor b;
    layer1_outputs(5713) <= not (a and b);
    layer1_outputs(5714) <= b;
    layer1_outputs(5715) <= not b;
    layer1_outputs(5716) <= not b;
    layer1_outputs(5717) <= not (a and b);
    layer1_outputs(5718) <= not b or a;
    layer1_outputs(5719) <= a;
    layer1_outputs(5720) <= not b;
    layer1_outputs(5721) <= not b;
    layer1_outputs(5722) <= a and not b;
    layer1_outputs(5723) <= not b or a;
    layer1_outputs(5724) <= b;
    layer1_outputs(5725) <= not b;
    layer1_outputs(5726) <= not b or a;
    layer1_outputs(5727) <= not (a or b);
    layer1_outputs(5728) <= a and b;
    layer1_outputs(5729) <= b and not a;
    layer1_outputs(5730) <= a;
    layer1_outputs(5731) <= not b;
    layer1_outputs(5732) <= not a or b;
    layer1_outputs(5733) <= b;
    layer1_outputs(5734) <= b and not a;
    layer1_outputs(5735) <= b;
    layer1_outputs(5736) <= b;
    layer1_outputs(5737) <= not (a or b);
    layer1_outputs(5738) <= not (a xor b);
    layer1_outputs(5739) <= not (a and b);
    layer1_outputs(5740) <= not a;
    layer1_outputs(5741) <= not (a and b);
    layer1_outputs(5742) <= a and b;
    layer1_outputs(5743) <= b;
    layer1_outputs(5744) <= a xor b;
    layer1_outputs(5745) <= not (a or b);
    layer1_outputs(5746) <= b;
    layer1_outputs(5747) <= not (a or b);
    layer1_outputs(5748) <= b;
    layer1_outputs(5749) <= a;
    layer1_outputs(5750) <= a and b;
    layer1_outputs(5751) <= not (a and b);
    layer1_outputs(5752) <= not a;
    layer1_outputs(5753) <= a and not b;
    layer1_outputs(5754) <= a or b;
    layer1_outputs(5755) <= not b or a;
    layer1_outputs(5756) <= not (a and b);
    layer1_outputs(5757) <= a or b;
    layer1_outputs(5758) <= a xor b;
    layer1_outputs(5759) <= a and not b;
    layer1_outputs(5760) <= b and not a;
    layer1_outputs(5761) <= b and not a;
    layer1_outputs(5762) <= b and not a;
    layer1_outputs(5763) <= 1'b1;
    layer1_outputs(5764) <= b and not a;
    layer1_outputs(5765) <= not a or b;
    layer1_outputs(5766) <= a and b;
    layer1_outputs(5767) <= b and not a;
    layer1_outputs(5768) <= b;
    layer1_outputs(5769) <= 1'b0;
    layer1_outputs(5770) <= not b or a;
    layer1_outputs(5771) <= a;
    layer1_outputs(5772) <= a;
    layer1_outputs(5773) <= a xor b;
    layer1_outputs(5774) <= a and not b;
    layer1_outputs(5775) <= not b;
    layer1_outputs(5776) <= not b or a;
    layer1_outputs(5777) <= 1'b1;
    layer1_outputs(5778) <= not b;
    layer1_outputs(5779) <= not (a and b);
    layer1_outputs(5780) <= b;
    layer1_outputs(5781) <= 1'b1;
    layer1_outputs(5782) <= not a or b;
    layer1_outputs(5783) <= a;
    layer1_outputs(5784) <= not (a and b);
    layer1_outputs(5785) <= not (a and b);
    layer1_outputs(5786) <= not b or a;
    layer1_outputs(5787) <= a;
    layer1_outputs(5788) <= a and not b;
    layer1_outputs(5789) <= a xor b;
    layer1_outputs(5790) <= a xor b;
    layer1_outputs(5791) <= a;
    layer1_outputs(5792) <= not (a or b);
    layer1_outputs(5793) <= not b;
    layer1_outputs(5794) <= not b;
    layer1_outputs(5795) <= not b or a;
    layer1_outputs(5796) <= not a;
    layer1_outputs(5797) <= not (a and b);
    layer1_outputs(5798) <= a;
    layer1_outputs(5799) <= a;
    layer1_outputs(5800) <= a or b;
    layer1_outputs(5801) <= a xor b;
    layer1_outputs(5802) <= b and not a;
    layer1_outputs(5803) <= a;
    layer1_outputs(5804) <= b;
    layer1_outputs(5805) <= a and not b;
    layer1_outputs(5806) <= b;
    layer1_outputs(5807) <= not a or b;
    layer1_outputs(5808) <= not b;
    layer1_outputs(5809) <= not (a and b);
    layer1_outputs(5810) <= not b;
    layer1_outputs(5811) <= b and not a;
    layer1_outputs(5812) <= not b or a;
    layer1_outputs(5813) <= a or b;
    layer1_outputs(5814) <= b and not a;
    layer1_outputs(5815) <= not (a or b);
    layer1_outputs(5816) <= not a;
    layer1_outputs(5817) <= not (a xor b);
    layer1_outputs(5818) <= not (a or b);
    layer1_outputs(5819) <= not b or a;
    layer1_outputs(5820) <= b;
    layer1_outputs(5821) <= not (a xor b);
    layer1_outputs(5822) <= b;
    layer1_outputs(5823) <= a xor b;
    layer1_outputs(5824) <= a or b;
    layer1_outputs(5825) <= a and b;
    layer1_outputs(5826) <= not (a and b);
    layer1_outputs(5827) <= not (a and b);
    layer1_outputs(5828) <= b;
    layer1_outputs(5829) <= not b or a;
    layer1_outputs(5830) <= a or b;
    layer1_outputs(5831) <= not a or b;
    layer1_outputs(5832) <= not b or a;
    layer1_outputs(5833) <= b and not a;
    layer1_outputs(5834) <= a or b;
    layer1_outputs(5835) <= not (a and b);
    layer1_outputs(5836) <= not b or a;
    layer1_outputs(5837) <= 1'b1;
    layer1_outputs(5838) <= 1'b1;
    layer1_outputs(5839) <= b;
    layer1_outputs(5840) <= 1'b0;
    layer1_outputs(5841) <= a;
    layer1_outputs(5842) <= b and not a;
    layer1_outputs(5843) <= not b;
    layer1_outputs(5844) <= not b;
    layer1_outputs(5845) <= 1'b1;
    layer1_outputs(5846) <= not a;
    layer1_outputs(5847) <= not a;
    layer1_outputs(5848) <= not a;
    layer1_outputs(5849) <= not a;
    layer1_outputs(5850) <= a and b;
    layer1_outputs(5851) <= b;
    layer1_outputs(5852) <= a;
    layer1_outputs(5853) <= a and b;
    layer1_outputs(5854) <= not b;
    layer1_outputs(5855) <= a and not b;
    layer1_outputs(5856) <= a;
    layer1_outputs(5857) <= not b or a;
    layer1_outputs(5858) <= not b;
    layer1_outputs(5859) <= not (a or b);
    layer1_outputs(5860) <= b;
    layer1_outputs(5861) <= a xor b;
    layer1_outputs(5862) <= 1'b1;
    layer1_outputs(5863) <= b and not a;
    layer1_outputs(5864) <= b;
    layer1_outputs(5865) <= 1'b0;
    layer1_outputs(5866) <= not a;
    layer1_outputs(5867) <= b;
    layer1_outputs(5868) <= a xor b;
    layer1_outputs(5869) <= not b or a;
    layer1_outputs(5870) <= b;
    layer1_outputs(5871) <= b;
    layer1_outputs(5872) <= 1'b0;
    layer1_outputs(5873) <= b and not a;
    layer1_outputs(5874) <= b;
    layer1_outputs(5875) <= not b or a;
    layer1_outputs(5876) <= b and not a;
    layer1_outputs(5877) <= a or b;
    layer1_outputs(5878) <= not (a xor b);
    layer1_outputs(5879) <= a xor b;
    layer1_outputs(5880) <= b;
    layer1_outputs(5881) <= a and not b;
    layer1_outputs(5882) <= a and not b;
    layer1_outputs(5883) <= not (a or b);
    layer1_outputs(5884) <= b and not a;
    layer1_outputs(5885) <= not b or a;
    layer1_outputs(5886) <= b;
    layer1_outputs(5887) <= not (a xor b);
    layer1_outputs(5888) <= a and b;
    layer1_outputs(5889) <= a and not b;
    layer1_outputs(5890) <= b;
    layer1_outputs(5891) <= a;
    layer1_outputs(5892) <= b and not a;
    layer1_outputs(5893) <= not (a or b);
    layer1_outputs(5894) <= b and not a;
    layer1_outputs(5895) <= not (a or b);
    layer1_outputs(5896) <= not b or a;
    layer1_outputs(5897) <= a;
    layer1_outputs(5898) <= not b or a;
    layer1_outputs(5899) <= a and b;
    layer1_outputs(5900) <= not (a and b);
    layer1_outputs(5901) <= a and b;
    layer1_outputs(5902) <= not (a and b);
    layer1_outputs(5903) <= 1'b1;
    layer1_outputs(5904) <= a or b;
    layer1_outputs(5905) <= a;
    layer1_outputs(5906) <= a or b;
    layer1_outputs(5907) <= not (a and b);
    layer1_outputs(5908) <= not a or b;
    layer1_outputs(5909) <= b and not a;
    layer1_outputs(5910) <= not a or b;
    layer1_outputs(5911) <= not a;
    layer1_outputs(5912) <= not (a and b);
    layer1_outputs(5913) <= not b;
    layer1_outputs(5914) <= a or b;
    layer1_outputs(5915) <= 1'b1;
    layer1_outputs(5916) <= a;
    layer1_outputs(5917) <= not (a and b);
    layer1_outputs(5918) <= 1'b0;
    layer1_outputs(5919) <= not b;
    layer1_outputs(5920) <= a and not b;
    layer1_outputs(5921) <= a and not b;
    layer1_outputs(5922) <= not b;
    layer1_outputs(5923) <= not a or b;
    layer1_outputs(5924) <= not (a xor b);
    layer1_outputs(5925) <= not b;
    layer1_outputs(5926) <= a or b;
    layer1_outputs(5927) <= b and not a;
    layer1_outputs(5928) <= not b or a;
    layer1_outputs(5929) <= a or b;
    layer1_outputs(5930) <= a xor b;
    layer1_outputs(5931) <= not b;
    layer1_outputs(5932) <= not (a or b);
    layer1_outputs(5933) <= not a or b;
    layer1_outputs(5934) <= a and b;
    layer1_outputs(5935) <= not a;
    layer1_outputs(5936) <= a xor b;
    layer1_outputs(5937) <= not a or b;
    layer1_outputs(5938) <= not a;
    layer1_outputs(5939) <= a;
    layer1_outputs(5940) <= a;
    layer1_outputs(5941) <= not b;
    layer1_outputs(5942) <= a;
    layer1_outputs(5943) <= a or b;
    layer1_outputs(5944) <= a;
    layer1_outputs(5945) <= a and not b;
    layer1_outputs(5946) <= a and not b;
    layer1_outputs(5947) <= a and not b;
    layer1_outputs(5948) <= not b;
    layer1_outputs(5949) <= b and not a;
    layer1_outputs(5950) <= a xor b;
    layer1_outputs(5951) <= not a;
    layer1_outputs(5952) <= not (a or b);
    layer1_outputs(5953) <= not b or a;
    layer1_outputs(5954) <= 1'b0;
    layer1_outputs(5955) <= not b;
    layer1_outputs(5956) <= not a or b;
    layer1_outputs(5957) <= a and b;
    layer1_outputs(5958) <= a and b;
    layer1_outputs(5959) <= a xor b;
    layer1_outputs(5960) <= 1'b1;
    layer1_outputs(5961) <= b and not a;
    layer1_outputs(5962) <= a;
    layer1_outputs(5963) <= not b or a;
    layer1_outputs(5964) <= not (a or b);
    layer1_outputs(5965) <= not b or a;
    layer1_outputs(5966) <= not b or a;
    layer1_outputs(5967) <= a and not b;
    layer1_outputs(5968) <= not a;
    layer1_outputs(5969) <= not (a and b);
    layer1_outputs(5970) <= a;
    layer1_outputs(5971) <= a;
    layer1_outputs(5972) <= a;
    layer1_outputs(5973) <= a xor b;
    layer1_outputs(5974) <= not b or a;
    layer1_outputs(5975) <= not b or a;
    layer1_outputs(5976) <= a;
    layer1_outputs(5977) <= 1'b1;
    layer1_outputs(5978) <= not (a xor b);
    layer1_outputs(5979) <= not a;
    layer1_outputs(5980) <= b and not a;
    layer1_outputs(5981) <= not b;
    layer1_outputs(5982) <= a;
    layer1_outputs(5983) <= not b;
    layer1_outputs(5984) <= not (a xor b);
    layer1_outputs(5985) <= not a;
    layer1_outputs(5986) <= not b or a;
    layer1_outputs(5987) <= not (a and b);
    layer1_outputs(5988) <= not a or b;
    layer1_outputs(5989) <= not (a and b);
    layer1_outputs(5990) <= a or b;
    layer1_outputs(5991) <= a and b;
    layer1_outputs(5992) <= not a or b;
    layer1_outputs(5993) <= a and not b;
    layer1_outputs(5994) <= not a or b;
    layer1_outputs(5995) <= a;
    layer1_outputs(5996) <= a and b;
    layer1_outputs(5997) <= b;
    layer1_outputs(5998) <= b;
    layer1_outputs(5999) <= not a or b;
    layer1_outputs(6000) <= a and not b;
    layer1_outputs(6001) <= a and not b;
    layer1_outputs(6002) <= not a;
    layer1_outputs(6003) <= a and b;
    layer1_outputs(6004) <= not b;
    layer1_outputs(6005) <= not a;
    layer1_outputs(6006) <= not b;
    layer1_outputs(6007) <= a or b;
    layer1_outputs(6008) <= a xor b;
    layer1_outputs(6009) <= not a;
    layer1_outputs(6010) <= a and not b;
    layer1_outputs(6011) <= not b;
    layer1_outputs(6012) <= not b;
    layer1_outputs(6013) <= a;
    layer1_outputs(6014) <= 1'b1;
    layer1_outputs(6015) <= a or b;
    layer1_outputs(6016) <= not b;
    layer1_outputs(6017) <= not b;
    layer1_outputs(6018) <= a;
    layer1_outputs(6019) <= not a or b;
    layer1_outputs(6020) <= not a or b;
    layer1_outputs(6021) <= not b or a;
    layer1_outputs(6022) <= a and not b;
    layer1_outputs(6023) <= 1'b1;
    layer1_outputs(6024) <= not a or b;
    layer1_outputs(6025) <= a and b;
    layer1_outputs(6026) <= a and not b;
    layer1_outputs(6027) <= a and b;
    layer1_outputs(6028) <= a and b;
    layer1_outputs(6029) <= 1'b1;
    layer1_outputs(6030) <= a or b;
    layer1_outputs(6031) <= b;
    layer1_outputs(6032) <= not (a and b);
    layer1_outputs(6033) <= not (a or b);
    layer1_outputs(6034) <= a or b;
    layer1_outputs(6035) <= 1'b0;
    layer1_outputs(6036) <= a and b;
    layer1_outputs(6037) <= not b or a;
    layer1_outputs(6038) <= not b;
    layer1_outputs(6039) <= a;
    layer1_outputs(6040) <= not (a xor b);
    layer1_outputs(6041) <= b and not a;
    layer1_outputs(6042) <= not (a and b);
    layer1_outputs(6043) <= a xor b;
    layer1_outputs(6044) <= a and b;
    layer1_outputs(6045) <= a;
    layer1_outputs(6046) <= a and not b;
    layer1_outputs(6047) <= a and b;
    layer1_outputs(6048) <= b and not a;
    layer1_outputs(6049) <= a and b;
    layer1_outputs(6050) <= a and not b;
    layer1_outputs(6051) <= not b or a;
    layer1_outputs(6052) <= b and not a;
    layer1_outputs(6053) <= not b;
    layer1_outputs(6054) <= not b;
    layer1_outputs(6055) <= a and not b;
    layer1_outputs(6056) <= 1'b1;
    layer1_outputs(6057) <= a and not b;
    layer1_outputs(6058) <= a and b;
    layer1_outputs(6059) <= b and not a;
    layer1_outputs(6060) <= not b;
    layer1_outputs(6061) <= b;
    layer1_outputs(6062) <= not b;
    layer1_outputs(6063) <= not b;
    layer1_outputs(6064) <= b;
    layer1_outputs(6065) <= a and not b;
    layer1_outputs(6066) <= a and not b;
    layer1_outputs(6067) <= not (a xor b);
    layer1_outputs(6068) <= not b or a;
    layer1_outputs(6069) <= a and b;
    layer1_outputs(6070) <= b;
    layer1_outputs(6071) <= a and not b;
    layer1_outputs(6072) <= not a or b;
    layer1_outputs(6073) <= not b;
    layer1_outputs(6074) <= not b;
    layer1_outputs(6075) <= a;
    layer1_outputs(6076) <= a;
    layer1_outputs(6077) <= not a or b;
    layer1_outputs(6078) <= a;
    layer1_outputs(6079) <= a or b;
    layer1_outputs(6080) <= a xor b;
    layer1_outputs(6081) <= not (a and b);
    layer1_outputs(6082) <= b and not a;
    layer1_outputs(6083) <= not (a or b);
    layer1_outputs(6084) <= not (a xor b);
    layer1_outputs(6085) <= not a;
    layer1_outputs(6086) <= not a or b;
    layer1_outputs(6087) <= a xor b;
    layer1_outputs(6088) <= a and not b;
    layer1_outputs(6089) <= a;
    layer1_outputs(6090) <= 1'b1;
    layer1_outputs(6091) <= a xor b;
    layer1_outputs(6092) <= not a;
    layer1_outputs(6093) <= not b;
    layer1_outputs(6094) <= not a;
    layer1_outputs(6095) <= a and not b;
    layer1_outputs(6096) <= b;
    layer1_outputs(6097) <= a or b;
    layer1_outputs(6098) <= b and not a;
    layer1_outputs(6099) <= b and not a;
    layer1_outputs(6100) <= a and not b;
    layer1_outputs(6101) <= not a;
    layer1_outputs(6102) <= b;
    layer1_outputs(6103) <= b;
    layer1_outputs(6104) <= not b;
    layer1_outputs(6105) <= not (a and b);
    layer1_outputs(6106) <= not a or b;
    layer1_outputs(6107) <= b and not a;
    layer1_outputs(6108) <= a;
    layer1_outputs(6109) <= not (a and b);
    layer1_outputs(6110) <= 1'b0;
    layer1_outputs(6111) <= not b;
    layer1_outputs(6112) <= not a;
    layer1_outputs(6113) <= not a;
    layer1_outputs(6114) <= a;
    layer1_outputs(6115) <= not (a or b);
    layer1_outputs(6116) <= a xor b;
    layer1_outputs(6117) <= a or b;
    layer1_outputs(6118) <= a and b;
    layer1_outputs(6119) <= not (a xor b);
    layer1_outputs(6120) <= not a;
    layer1_outputs(6121) <= a;
    layer1_outputs(6122) <= not (a or b);
    layer1_outputs(6123) <= not a or b;
    layer1_outputs(6124) <= 1'b1;
    layer1_outputs(6125) <= not a or b;
    layer1_outputs(6126) <= not (a and b);
    layer1_outputs(6127) <= not a;
    layer1_outputs(6128) <= a;
    layer1_outputs(6129) <= a xor b;
    layer1_outputs(6130) <= a and b;
    layer1_outputs(6131) <= not (a xor b);
    layer1_outputs(6132) <= a;
    layer1_outputs(6133) <= a and b;
    layer1_outputs(6134) <= not (a and b);
    layer1_outputs(6135) <= not a;
    layer1_outputs(6136) <= not (a or b);
    layer1_outputs(6137) <= not b;
    layer1_outputs(6138) <= not (a and b);
    layer1_outputs(6139) <= not b or a;
    layer1_outputs(6140) <= not b;
    layer1_outputs(6141) <= b and not a;
    layer1_outputs(6142) <= not a;
    layer1_outputs(6143) <= not a;
    layer1_outputs(6144) <= not (a and b);
    layer1_outputs(6145) <= b;
    layer1_outputs(6146) <= b;
    layer1_outputs(6147) <= b and not a;
    layer1_outputs(6148) <= a xor b;
    layer1_outputs(6149) <= a and not b;
    layer1_outputs(6150) <= b;
    layer1_outputs(6151) <= not a;
    layer1_outputs(6152) <= 1'b1;
    layer1_outputs(6153) <= not (a or b);
    layer1_outputs(6154) <= not b or a;
    layer1_outputs(6155) <= a and b;
    layer1_outputs(6156) <= a and b;
    layer1_outputs(6157) <= a and not b;
    layer1_outputs(6158) <= b;
    layer1_outputs(6159) <= 1'b0;
    layer1_outputs(6160) <= 1'b1;
    layer1_outputs(6161) <= not (a xor b);
    layer1_outputs(6162) <= not (a and b);
    layer1_outputs(6163) <= not b;
    layer1_outputs(6164) <= not b;
    layer1_outputs(6165) <= not (a or b);
    layer1_outputs(6166) <= a and b;
    layer1_outputs(6167) <= a or b;
    layer1_outputs(6168) <= a xor b;
    layer1_outputs(6169) <= not (a or b);
    layer1_outputs(6170) <= not b;
    layer1_outputs(6171) <= a;
    layer1_outputs(6172) <= a xor b;
    layer1_outputs(6173) <= not (a and b);
    layer1_outputs(6174) <= a xor b;
    layer1_outputs(6175) <= not a;
    layer1_outputs(6176) <= not b;
    layer1_outputs(6177) <= b and not a;
    layer1_outputs(6178) <= b;
    layer1_outputs(6179) <= not a;
    layer1_outputs(6180) <= not (a or b);
    layer1_outputs(6181) <= a and b;
    layer1_outputs(6182) <= a or b;
    layer1_outputs(6183) <= b;
    layer1_outputs(6184) <= not (a or b);
    layer1_outputs(6185) <= not b;
    layer1_outputs(6186) <= not (a or b);
    layer1_outputs(6187) <= 1'b1;
    layer1_outputs(6188) <= a and b;
    layer1_outputs(6189) <= not (a or b);
    layer1_outputs(6190) <= 1'b1;
    layer1_outputs(6191) <= a;
    layer1_outputs(6192) <= not a or b;
    layer1_outputs(6193) <= not (a or b);
    layer1_outputs(6194) <= a;
    layer1_outputs(6195) <= not a;
    layer1_outputs(6196) <= b;
    layer1_outputs(6197) <= b and not a;
    layer1_outputs(6198) <= not (a and b);
    layer1_outputs(6199) <= 1'b0;
    layer1_outputs(6200) <= b;
    layer1_outputs(6201) <= a or b;
    layer1_outputs(6202) <= a xor b;
    layer1_outputs(6203) <= a and not b;
    layer1_outputs(6204) <= not b or a;
    layer1_outputs(6205) <= not a;
    layer1_outputs(6206) <= not (a or b);
    layer1_outputs(6207) <= a;
    layer1_outputs(6208) <= not (a or b);
    layer1_outputs(6209) <= not (a and b);
    layer1_outputs(6210) <= a xor b;
    layer1_outputs(6211) <= not a;
    layer1_outputs(6212) <= a;
    layer1_outputs(6213) <= a and b;
    layer1_outputs(6214) <= not a;
    layer1_outputs(6215) <= not a or b;
    layer1_outputs(6216) <= a or b;
    layer1_outputs(6217) <= not b;
    layer1_outputs(6218) <= not a;
    layer1_outputs(6219) <= a;
    layer1_outputs(6220) <= a or b;
    layer1_outputs(6221) <= b;
    layer1_outputs(6222) <= b and not a;
    layer1_outputs(6223) <= not b or a;
    layer1_outputs(6224) <= a and b;
    layer1_outputs(6225) <= not b;
    layer1_outputs(6226) <= a xor b;
    layer1_outputs(6227) <= not a or b;
    layer1_outputs(6228) <= a or b;
    layer1_outputs(6229) <= b;
    layer1_outputs(6230) <= not a or b;
    layer1_outputs(6231) <= not (a and b);
    layer1_outputs(6232) <= b and not a;
    layer1_outputs(6233) <= a xor b;
    layer1_outputs(6234) <= not b or a;
    layer1_outputs(6235) <= 1'b1;
    layer1_outputs(6236) <= not b;
    layer1_outputs(6237) <= a and not b;
    layer1_outputs(6238) <= not b;
    layer1_outputs(6239) <= not b;
    layer1_outputs(6240) <= not (a or b);
    layer1_outputs(6241) <= a;
    layer1_outputs(6242) <= b;
    layer1_outputs(6243) <= a and b;
    layer1_outputs(6244) <= a or b;
    layer1_outputs(6245) <= a xor b;
    layer1_outputs(6246) <= a and not b;
    layer1_outputs(6247) <= not a or b;
    layer1_outputs(6248) <= not b;
    layer1_outputs(6249) <= not b or a;
    layer1_outputs(6250) <= not (a or b);
    layer1_outputs(6251) <= not b;
    layer1_outputs(6252) <= not (a xor b);
    layer1_outputs(6253) <= 1'b0;
    layer1_outputs(6254) <= 1'b0;
    layer1_outputs(6255) <= a or b;
    layer1_outputs(6256) <= not (a or b);
    layer1_outputs(6257) <= a and not b;
    layer1_outputs(6258) <= a and not b;
    layer1_outputs(6259) <= not (a or b);
    layer1_outputs(6260) <= a or b;
    layer1_outputs(6261) <= not (a and b);
    layer1_outputs(6262) <= b;
    layer1_outputs(6263) <= b and not a;
    layer1_outputs(6264) <= not a;
    layer1_outputs(6265) <= a or b;
    layer1_outputs(6266) <= not (a and b);
    layer1_outputs(6267) <= not a;
    layer1_outputs(6268) <= b;
    layer1_outputs(6269) <= not a or b;
    layer1_outputs(6270) <= 1'b0;
    layer1_outputs(6271) <= not a;
    layer1_outputs(6272) <= a and not b;
    layer1_outputs(6273) <= not (a and b);
    layer1_outputs(6274) <= a;
    layer1_outputs(6275) <= a and not b;
    layer1_outputs(6276) <= a or b;
    layer1_outputs(6277) <= not (a xor b);
    layer1_outputs(6278) <= b;
    layer1_outputs(6279) <= not (a and b);
    layer1_outputs(6280) <= not (a xor b);
    layer1_outputs(6281) <= not a;
    layer1_outputs(6282) <= not (a or b);
    layer1_outputs(6283) <= not a;
    layer1_outputs(6284) <= not b;
    layer1_outputs(6285) <= a and b;
    layer1_outputs(6286) <= not b;
    layer1_outputs(6287) <= a or b;
    layer1_outputs(6288) <= not (a xor b);
    layer1_outputs(6289) <= 1'b0;
    layer1_outputs(6290) <= a and not b;
    layer1_outputs(6291) <= not a or b;
    layer1_outputs(6292) <= b;
    layer1_outputs(6293) <= not b;
    layer1_outputs(6294) <= a and not b;
    layer1_outputs(6295) <= a or b;
    layer1_outputs(6296) <= not (a and b);
    layer1_outputs(6297) <= a;
    layer1_outputs(6298) <= b and not a;
    layer1_outputs(6299) <= a;
    layer1_outputs(6300) <= a xor b;
    layer1_outputs(6301) <= a and not b;
    layer1_outputs(6302) <= 1'b1;
    layer1_outputs(6303) <= not a or b;
    layer1_outputs(6304) <= a;
    layer1_outputs(6305) <= a xor b;
    layer1_outputs(6306) <= not a or b;
    layer1_outputs(6307) <= a or b;
    layer1_outputs(6308) <= not b or a;
    layer1_outputs(6309) <= not b;
    layer1_outputs(6310) <= not (a and b);
    layer1_outputs(6311) <= b;
    layer1_outputs(6312) <= b;
    layer1_outputs(6313) <= a;
    layer1_outputs(6314) <= b and not a;
    layer1_outputs(6315) <= a;
    layer1_outputs(6316) <= not b;
    layer1_outputs(6317) <= not a or b;
    layer1_outputs(6318) <= a and b;
    layer1_outputs(6319) <= a or b;
    layer1_outputs(6320) <= not b or a;
    layer1_outputs(6321) <= not b;
    layer1_outputs(6322) <= not (a and b);
    layer1_outputs(6323) <= b;
    layer1_outputs(6324) <= not b;
    layer1_outputs(6325) <= not a;
    layer1_outputs(6326) <= a xor b;
    layer1_outputs(6327) <= a;
    layer1_outputs(6328) <= a or b;
    layer1_outputs(6329) <= 1'b1;
    layer1_outputs(6330) <= not b or a;
    layer1_outputs(6331) <= not a or b;
    layer1_outputs(6332) <= b;
    layer1_outputs(6333) <= a or b;
    layer1_outputs(6334) <= not (a xor b);
    layer1_outputs(6335) <= a;
    layer1_outputs(6336) <= 1'b0;
    layer1_outputs(6337) <= not (a xor b);
    layer1_outputs(6338) <= 1'b1;
    layer1_outputs(6339) <= a or b;
    layer1_outputs(6340) <= b;
    layer1_outputs(6341) <= a and b;
    layer1_outputs(6342) <= not (a or b);
    layer1_outputs(6343) <= not b;
    layer1_outputs(6344) <= not a;
    layer1_outputs(6345) <= a and not b;
    layer1_outputs(6346) <= not b;
    layer1_outputs(6347) <= not b;
    layer1_outputs(6348) <= not b or a;
    layer1_outputs(6349) <= a;
    layer1_outputs(6350) <= a and b;
    layer1_outputs(6351) <= not a;
    layer1_outputs(6352) <= not b;
    layer1_outputs(6353) <= not (a xor b);
    layer1_outputs(6354) <= a or b;
    layer1_outputs(6355) <= not (a or b);
    layer1_outputs(6356) <= not (a and b);
    layer1_outputs(6357) <= a;
    layer1_outputs(6358) <= 1'b0;
    layer1_outputs(6359) <= b;
    layer1_outputs(6360) <= a or b;
    layer1_outputs(6361) <= not b;
    layer1_outputs(6362) <= not b;
    layer1_outputs(6363) <= not a;
    layer1_outputs(6364) <= a;
    layer1_outputs(6365) <= not a;
    layer1_outputs(6366) <= not (a or b);
    layer1_outputs(6367) <= not (a or b);
    layer1_outputs(6368) <= 1'b0;
    layer1_outputs(6369) <= a and not b;
    layer1_outputs(6370) <= b;
    layer1_outputs(6371) <= a;
    layer1_outputs(6372) <= not a;
    layer1_outputs(6373) <= not a;
    layer1_outputs(6374) <= not b or a;
    layer1_outputs(6375) <= not a;
    layer1_outputs(6376) <= not (a xor b);
    layer1_outputs(6377) <= a or b;
    layer1_outputs(6378) <= b and not a;
    layer1_outputs(6379) <= not (a or b);
    layer1_outputs(6380) <= not (a or b);
    layer1_outputs(6381) <= b and not a;
    layer1_outputs(6382) <= not a;
    layer1_outputs(6383) <= not (a and b);
    layer1_outputs(6384) <= not a;
    layer1_outputs(6385) <= not (a and b);
    layer1_outputs(6386) <= a or b;
    layer1_outputs(6387) <= not (a and b);
    layer1_outputs(6388) <= a and b;
    layer1_outputs(6389) <= not a or b;
    layer1_outputs(6390) <= not a;
    layer1_outputs(6391) <= b;
    layer1_outputs(6392) <= not b or a;
    layer1_outputs(6393) <= a;
    layer1_outputs(6394) <= not b or a;
    layer1_outputs(6395) <= 1'b0;
    layer1_outputs(6396) <= not a;
    layer1_outputs(6397) <= b and not a;
    layer1_outputs(6398) <= b and not a;
    layer1_outputs(6399) <= not (a and b);
    layer1_outputs(6400) <= not b;
    layer1_outputs(6401) <= not a;
    layer1_outputs(6402) <= not (a xor b);
    layer1_outputs(6403) <= a and not b;
    layer1_outputs(6404) <= b and not a;
    layer1_outputs(6405) <= b;
    layer1_outputs(6406) <= a and b;
    layer1_outputs(6407) <= not a;
    layer1_outputs(6408) <= 1'b0;
    layer1_outputs(6409) <= not (a and b);
    layer1_outputs(6410) <= not b or a;
    layer1_outputs(6411) <= not b or a;
    layer1_outputs(6412) <= not a or b;
    layer1_outputs(6413) <= not a or b;
    layer1_outputs(6414) <= not (a or b);
    layer1_outputs(6415) <= a or b;
    layer1_outputs(6416) <= not (a and b);
    layer1_outputs(6417) <= not (a and b);
    layer1_outputs(6418) <= b;
    layer1_outputs(6419) <= not a;
    layer1_outputs(6420) <= 1'b1;
    layer1_outputs(6421) <= a xor b;
    layer1_outputs(6422) <= not b;
    layer1_outputs(6423) <= b;
    layer1_outputs(6424) <= a and b;
    layer1_outputs(6425) <= not (a and b);
    layer1_outputs(6426) <= a;
    layer1_outputs(6427) <= b;
    layer1_outputs(6428) <= a xor b;
    layer1_outputs(6429) <= not (a xor b);
    layer1_outputs(6430) <= not (a or b);
    layer1_outputs(6431) <= not b;
    layer1_outputs(6432) <= a or b;
    layer1_outputs(6433) <= b and not a;
    layer1_outputs(6434) <= not b;
    layer1_outputs(6435) <= not (a or b);
    layer1_outputs(6436) <= a;
    layer1_outputs(6437) <= a and b;
    layer1_outputs(6438) <= not b or a;
    layer1_outputs(6439) <= not a;
    layer1_outputs(6440) <= not (a or b);
    layer1_outputs(6441) <= 1'b0;
    layer1_outputs(6442) <= a and not b;
    layer1_outputs(6443) <= 1'b0;
    layer1_outputs(6444) <= a xor b;
    layer1_outputs(6445) <= 1'b1;
    layer1_outputs(6446) <= not a;
    layer1_outputs(6447) <= a;
    layer1_outputs(6448) <= b;
    layer1_outputs(6449) <= 1'b0;
    layer1_outputs(6450) <= b;
    layer1_outputs(6451) <= b and not a;
    layer1_outputs(6452) <= not b;
    layer1_outputs(6453) <= 1'b0;
    layer1_outputs(6454) <= not (a and b);
    layer1_outputs(6455) <= b;
    layer1_outputs(6456) <= not (a or b);
    layer1_outputs(6457) <= not (a xor b);
    layer1_outputs(6458) <= not (a and b);
    layer1_outputs(6459) <= b;
    layer1_outputs(6460) <= not a or b;
    layer1_outputs(6461) <= a and b;
    layer1_outputs(6462) <= a xor b;
    layer1_outputs(6463) <= not a;
    layer1_outputs(6464) <= a and not b;
    layer1_outputs(6465) <= a or b;
    layer1_outputs(6466) <= a;
    layer1_outputs(6467) <= a or b;
    layer1_outputs(6468) <= not a or b;
    layer1_outputs(6469) <= 1'b0;
    layer1_outputs(6470) <= not b;
    layer1_outputs(6471) <= not b;
    layer1_outputs(6472) <= 1'b0;
    layer1_outputs(6473) <= b and not a;
    layer1_outputs(6474) <= a;
    layer1_outputs(6475) <= not a;
    layer1_outputs(6476) <= 1'b0;
    layer1_outputs(6477) <= a and not b;
    layer1_outputs(6478) <= a;
    layer1_outputs(6479) <= 1'b0;
    layer1_outputs(6480) <= 1'b1;
    layer1_outputs(6481) <= b;
    layer1_outputs(6482) <= not b;
    layer1_outputs(6483) <= a;
    layer1_outputs(6484) <= not a;
    layer1_outputs(6485) <= not (a or b);
    layer1_outputs(6486) <= not a or b;
    layer1_outputs(6487) <= a or b;
    layer1_outputs(6488) <= not (a or b);
    layer1_outputs(6489) <= not a or b;
    layer1_outputs(6490) <= not a;
    layer1_outputs(6491) <= b and not a;
    layer1_outputs(6492) <= a or b;
    layer1_outputs(6493) <= not a or b;
    layer1_outputs(6494) <= a xor b;
    layer1_outputs(6495) <= not (a and b);
    layer1_outputs(6496) <= b;
    layer1_outputs(6497) <= a and not b;
    layer1_outputs(6498) <= a and not b;
    layer1_outputs(6499) <= b and not a;
    layer1_outputs(6500) <= not b;
    layer1_outputs(6501) <= b;
    layer1_outputs(6502) <= not (a and b);
    layer1_outputs(6503) <= not (a and b);
    layer1_outputs(6504) <= a xor b;
    layer1_outputs(6505) <= not (a and b);
    layer1_outputs(6506) <= not a;
    layer1_outputs(6507) <= not (a and b);
    layer1_outputs(6508) <= a;
    layer1_outputs(6509) <= not a;
    layer1_outputs(6510) <= not a;
    layer1_outputs(6511) <= a;
    layer1_outputs(6512) <= a and not b;
    layer1_outputs(6513) <= a and not b;
    layer1_outputs(6514) <= a xor b;
    layer1_outputs(6515) <= not (a xor b);
    layer1_outputs(6516) <= a xor b;
    layer1_outputs(6517) <= a or b;
    layer1_outputs(6518) <= not (a xor b);
    layer1_outputs(6519) <= b and not a;
    layer1_outputs(6520) <= not a or b;
    layer1_outputs(6521) <= not a;
    layer1_outputs(6522) <= b and not a;
    layer1_outputs(6523) <= a and not b;
    layer1_outputs(6524) <= not a or b;
    layer1_outputs(6525) <= a or b;
    layer1_outputs(6526) <= not (a and b);
    layer1_outputs(6527) <= b;
    layer1_outputs(6528) <= a and b;
    layer1_outputs(6529) <= a and not b;
    layer1_outputs(6530) <= b;
    layer1_outputs(6531) <= not (a or b);
    layer1_outputs(6532) <= not b or a;
    layer1_outputs(6533) <= not a or b;
    layer1_outputs(6534) <= not b or a;
    layer1_outputs(6535) <= not (a and b);
    layer1_outputs(6536) <= not a or b;
    layer1_outputs(6537) <= a and b;
    layer1_outputs(6538) <= 1'b1;
    layer1_outputs(6539) <= 1'b0;
    layer1_outputs(6540) <= a and not b;
    layer1_outputs(6541) <= not a;
    layer1_outputs(6542) <= not a or b;
    layer1_outputs(6543) <= a and not b;
    layer1_outputs(6544) <= 1'b1;
    layer1_outputs(6545) <= a or b;
    layer1_outputs(6546) <= 1'b1;
    layer1_outputs(6547) <= not b or a;
    layer1_outputs(6548) <= not (a xor b);
    layer1_outputs(6549) <= a or b;
    layer1_outputs(6550) <= not (a and b);
    layer1_outputs(6551) <= a and not b;
    layer1_outputs(6552) <= a xor b;
    layer1_outputs(6553) <= not b;
    layer1_outputs(6554) <= not (a or b);
    layer1_outputs(6555) <= not a;
    layer1_outputs(6556) <= not b;
    layer1_outputs(6557) <= a or b;
    layer1_outputs(6558) <= a and not b;
    layer1_outputs(6559) <= not (a or b);
    layer1_outputs(6560) <= not (a or b);
    layer1_outputs(6561) <= not (a or b);
    layer1_outputs(6562) <= a;
    layer1_outputs(6563) <= 1'b0;
    layer1_outputs(6564) <= not (a or b);
    layer1_outputs(6565) <= not (a or b);
    layer1_outputs(6566) <= not (a or b);
    layer1_outputs(6567) <= not a;
    layer1_outputs(6568) <= not a or b;
    layer1_outputs(6569) <= not (a xor b);
    layer1_outputs(6570) <= b;
    layer1_outputs(6571) <= b;
    layer1_outputs(6572) <= a;
    layer1_outputs(6573) <= not b;
    layer1_outputs(6574) <= not b;
    layer1_outputs(6575) <= not a or b;
    layer1_outputs(6576) <= a;
    layer1_outputs(6577) <= a xor b;
    layer1_outputs(6578) <= a and not b;
    layer1_outputs(6579) <= 1'b1;
    layer1_outputs(6580) <= 1'b1;
    layer1_outputs(6581) <= not (a and b);
    layer1_outputs(6582) <= b and not a;
    layer1_outputs(6583) <= not b;
    layer1_outputs(6584) <= a or b;
    layer1_outputs(6585) <= not (a and b);
    layer1_outputs(6586) <= not a or b;
    layer1_outputs(6587) <= a xor b;
    layer1_outputs(6588) <= not (a or b);
    layer1_outputs(6589) <= b and not a;
    layer1_outputs(6590) <= b;
    layer1_outputs(6591) <= b;
    layer1_outputs(6592) <= a and b;
    layer1_outputs(6593) <= a;
    layer1_outputs(6594) <= not (a xor b);
    layer1_outputs(6595) <= b;
    layer1_outputs(6596) <= a and b;
    layer1_outputs(6597) <= a xor b;
    layer1_outputs(6598) <= not (a or b);
    layer1_outputs(6599) <= not (a and b);
    layer1_outputs(6600) <= b and not a;
    layer1_outputs(6601) <= 1'b1;
    layer1_outputs(6602) <= b and not a;
    layer1_outputs(6603) <= a;
    layer1_outputs(6604) <= a xor b;
    layer1_outputs(6605) <= 1'b1;
    layer1_outputs(6606) <= 1'b0;
    layer1_outputs(6607) <= a;
    layer1_outputs(6608) <= not (a xor b);
    layer1_outputs(6609) <= a and not b;
    layer1_outputs(6610) <= b;
    layer1_outputs(6611) <= 1'b1;
    layer1_outputs(6612) <= not (a and b);
    layer1_outputs(6613) <= a;
    layer1_outputs(6614) <= a xor b;
    layer1_outputs(6615) <= a and b;
    layer1_outputs(6616) <= a and b;
    layer1_outputs(6617) <= a;
    layer1_outputs(6618) <= b and not a;
    layer1_outputs(6619) <= 1'b0;
    layer1_outputs(6620) <= not b or a;
    layer1_outputs(6621) <= a or b;
    layer1_outputs(6622) <= b and not a;
    layer1_outputs(6623) <= not b or a;
    layer1_outputs(6624) <= not b or a;
    layer1_outputs(6625) <= not a;
    layer1_outputs(6626) <= 1'b0;
    layer1_outputs(6627) <= not a;
    layer1_outputs(6628) <= not (a or b);
    layer1_outputs(6629) <= 1'b1;
    layer1_outputs(6630) <= a;
    layer1_outputs(6631) <= a and not b;
    layer1_outputs(6632) <= a and b;
    layer1_outputs(6633) <= not a;
    layer1_outputs(6634) <= not a;
    layer1_outputs(6635) <= not (a xor b);
    layer1_outputs(6636) <= a;
    layer1_outputs(6637) <= a and b;
    layer1_outputs(6638) <= a;
    layer1_outputs(6639) <= b;
    layer1_outputs(6640) <= not b or a;
    layer1_outputs(6641) <= not (a or b);
    layer1_outputs(6642) <= b and not a;
    layer1_outputs(6643) <= b;
    layer1_outputs(6644) <= not (a and b);
    layer1_outputs(6645) <= not (a and b);
    layer1_outputs(6646) <= not (a and b);
    layer1_outputs(6647) <= not a;
    layer1_outputs(6648) <= b;
    layer1_outputs(6649) <= b;
    layer1_outputs(6650) <= not (a xor b);
    layer1_outputs(6651) <= not (a or b);
    layer1_outputs(6652) <= not b;
    layer1_outputs(6653) <= not b or a;
    layer1_outputs(6654) <= a or b;
    layer1_outputs(6655) <= not (a or b);
    layer1_outputs(6656) <= a and b;
    layer1_outputs(6657) <= not a or b;
    layer1_outputs(6658) <= a;
    layer1_outputs(6659) <= not b or a;
    layer1_outputs(6660) <= not a;
    layer1_outputs(6661) <= not (a and b);
    layer1_outputs(6662) <= not (a xor b);
    layer1_outputs(6663) <= a or b;
    layer1_outputs(6664) <= a or b;
    layer1_outputs(6665) <= a and b;
    layer1_outputs(6666) <= not b;
    layer1_outputs(6667) <= not (a and b);
    layer1_outputs(6668) <= not a or b;
    layer1_outputs(6669) <= not b;
    layer1_outputs(6670) <= not (a or b);
    layer1_outputs(6671) <= not b or a;
    layer1_outputs(6672) <= not (a xor b);
    layer1_outputs(6673) <= not a;
    layer1_outputs(6674) <= b;
    layer1_outputs(6675) <= a;
    layer1_outputs(6676) <= not b or a;
    layer1_outputs(6677) <= not (a and b);
    layer1_outputs(6678) <= not (a and b);
    layer1_outputs(6679) <= b and not a;
    layer1_outputs(6680) <= not (a and b);
    layer1_outputs(6681) <= 1'b0;
    layer1_outputs(6682) <= a and b;
    layer1_outputs(6683) <= not a or b;
    layer1_outputs(6684) <= a;
    layer1_outputs(6685) <= not b or a;
    layer1_outputs(6686) <= b and not a;
    layer1_outputs(6687) <= not b or a;
    layer1_outputs(6688) <= a and b;
    layer1_outputs(6689) <= a or b;
    layer1_outputs(6690) <= 1'b1;
    layer1_outputs(6691) <= not (a xor b);
    layer1_outputs(6692) <= a;
    layer1_outputs(6693) <= not (a xor b);
    layer1_outputs(6694) <= not (a or b);
    layer1_outputs(6695) <= a xor b;
    layer1_outputs(6696) <= a and not b;
    layer1_outputs(6697) <= not (a and b);
    layer1_outputs(6698) <= not a or b;
    layer1_outputs(6699) <= a and not b;
    layer1_outputs(6700) <= not (a xor b);
    layer1_outputs(6701) <= a or b;
    layer1_outputs(6702) <= a and not b;
    layer1_outputs(6703) <= b;
    layer1_outputs(6704) <= not b;
    layer1_outputs(6705) <= not b;
    layer1_outputs(6706) <= not b;
    layer1_outputs(6707) <= b and not a;
    layer1_outputs(6708) <= not (a xor b);
    layer1_outputs(6709) <= not (a or b);
    layer1_outputs(6710) <= a;
    layer1_outputs(6711) <= a;
    layer1_outputs(6712) <= b and not a;
    layer1_outputs(6713) <= a and not b;
    layer1_outputs(6714) <= b and not a;
    layer1_outputs(6715) <= a or b;
    layer1_outputs(6716) <= 1'b0;
    layer1_outputs(6717) <= not b or a;
    layer1_outputs(6718) <= b and not a;
    layer1_outputs(6719) <= not (a and b);
    layer1_outputs(6720) <= not (a xor b);
    layer1_outputs(6721) <= not a or b;
    layer1_outputs(6722) <= not b;
    layer1_outputs(6723) <= a xor b;
    layer1_outputs(6724) <= not b or a;
    layer1_outputs(6725) <= not b;
    layer1_outputs(6726) <= b and not a;
    layer1_outputs(6727) <= not b or a;
    layer1_outputs(6728) <= not (a or b);
    layer1_outputs(6729) <= a xor b;
    layer1_outputs(6730) <= not a;
    layer1_outputs(6731) <= not b;
    layer1_outputs(6732) <= not (a and b);
    layer1_outputs(6733) <= not (a xor b);
    layer1_outputs(6734) <= not (a xor b);
    layer1_outputs(6735) <= b;
    layer1_outputs(6736) <= not a or b;
    layer1_outputs(6737) <= not (a xor b);
    layer1_outputs(6738) <= not (a xor b);
    layer1_outputs(6739) <= not b or a;
    layer1_outputs(6740) <= b and not a;
    layer1_outputs(6741) <= a or b;
    layer1_outputs(6742) <= b;
    layer1_outputs(6743) <= a;
    layer1_outputs(6744) <= not b;
    layer1_outputs(6745) <= not (a or b);
    layer1_outputs(6746) <= not (a and b);
    layer1_outputs(6747) <= not a;
    layer1_outputs(6748) <= 1'b1;
    layer1_outputs(6749) <= a and b;
    layer1_outputs(6750) <= a;
    layer1_outputs(6751) <= not (a and b);
    layer1_outputs(6752) <= not (a xor b);
    layer1_outputs(6753) <= not b or a;
    layer1_outputs(6754) <= not (a and b);
    layer1_outputs(6755) <= not a or b;
    layer1_outputs(6756) <= b;
    layer1_outputs(6757) <= a or b;
    layer1_outputs(6758) <= not (a and b);
    layer1_outputs(6759) <= not b or a;
    layer1_outputs(6760) <= not (a and b);
    layer1_outputs(6761) <= not b or a;
    layer1_outputs(6762) <= a;
    layer1_outputs(6763) <= a and not b;
    layer1_outputs(6764) <= not b;
    layer1_outputs(6765) <= not a;
    layer1_outputs(6766) <= a or b;
    layer1_outputs(6767) <= b and not a;
    layer1_outputs(6768) <= not (a xor b);
    layer1_outputs(6769) <= not (a xor b);
    layer1_outputs(6770) <= not b;
    layer1_outputs(6771) <= not a or b;
    layer1_outputs(6772) <= 1'b0;
    layer1_outputs(6773) <= a and b;
    layer1_outputs(6774) <= a and not b;
    layer1_outputs(6775) <= a and not b;
    layer1_outputs(6776) <= a;
    layer1_outputs(6777) <= a;
    layer1_outputs(6778) <= b;
    layer1_outputs(6779) <= not (a or b);
    layer1_outputs(6780) <= a xor b;
    layer1_outputs(6781) <= b;
    layer1_outputs(6782) <= not (a and b);
    layer1_outputs(6783) <= not b;
    layer1_outputs(6784) <= 1'b1;
    layer1_outputs(6785) <= 1'b1;
    layer1_outputs(6786) <= not b;
    layer1_outputs(6787) <= not (a xor b);
    layer1_outputs(6788) <= 1'b1;
    layer1_outputs(6789) <= b and not a;
    layer1_outputs(6790) <= b;
    layer1_outputs(6791) <= not b;
    layer1_outputs(6792) <= 1'b1;
    layer1_outputs(6793) <= not a or b;
    layer1_outputs(6794) <= not b;
    layer1_outputs(6795) <= not (a xor b);
    layer1_outputs(6796) <= a and not b;
    layer1_outputs(6797) <= not a;
    layer1_outputs(6798) <= b and not a;
    layer1_outputs(6799) <= a and not b;
    layer1_outputs(6800) <= not a;
    layer1_outputs(6801) <= a xor b;
    layer1_outputs(6802) <= not a;
    layer1_outputs(6803) <= a;
    layer1_outputs(6804) <= b;
    layer1_outputs(6805) <= a xor b;
    layer1_outputs(6806) <= a xor b;
    layer1_outputs(6807) <= not a;
    layer1_outputs(6808) <= not b or a;
    layer1_outputs(6809) <= not b;
    layer1_outputs(6810) <= a xor b;
    layer1_outputs(6811) <= not a;
    layer1_outputs(6812) <= a and b;
    layer1_outputs(6813) <= not b;
    layer1_outputs(6814) <= not a;
    layer1_outputs(6815) <= not b or a;
    layer1_outputs(6816) <= a xor b;
    layer1_outputs(6817) <= a and b;
    layer1_outputs(6818) <= not a;
    layer1_outputs(6819) <= b and not a;
    layer1_outputs(6820) <= a and b;
    layer1_outputs(6821) <= a xor b;
    layer1_outputs(6822) <= not a or b;
    layer1_outputs(6823) <= a;
    layer1_outputs(6824) <= not b;
    layer1_outputs(6825) <= a and b;
    layer1_outputs(6826) <= not b;
    layer1_outputs(6827) <= a xor b;
    layer1_outputs(6828) <= a and b;
    layer1_outputs(6829) <= not (a or b);
    layer1_outputs(6830) <= not b;
    layer1_outputs(6831) <= a or b;
    layer1_outputs(6832) <= a or b;
    layer1_outputs(6833) <= b and not a;
    layer1_outputs(6834) <= a;
    layer1_outputs(6835) <= a or b;
    layer1_outputs(6836) <= not a;
    layer1_outputs(6837) <= not b;
    layer1_outputs(6838) <= b;
    layer1_outputs(6839) <= not a;
    layer1_outputs(6840) <= b;
    layer1_outputs(6841) <= a and not b;
    layer1_outputs(6842) <= b and not a;
    layer1_outputs(6843) <= a xor b;
    layer1_outputs(6844) <= not a or b;
    layer1_outputs(6845) <= not a;
    layer1_outputs(6846) <= not (a or b);
    layer1_outputs(6847) <= a xor b;
    layer1_outputs(6848) <= not a;
    layer1_outputs(6849) <= a or b;
    layer1_outputs(6850) <= b and not a;
    layer1_outputs(6851) <= a and b;
    layer1_outputs(6852) <= a xor b;
    layer1_outputs(6853) <= a or b;
    layer1_outputs(6854) <= not b or a;
    layer1_outputs(6855) <= not (a xor b);
    layer1_outputs(6856) <= not b;
    layer1_outputs(6857) <= b and not a;
    layer1_outputs(6858) <= a and b;
    layer1_outputs(6859) <= a and b;
    layer1_outputs(6860) <= not a or b;
    layer1_outputs(6861) <= a or b;
    layer1_outputs(6862) <= a xor b;
    layer1_outputs(6863) <= not (a or b);
    layer1_outputs(6864) <= a and b;
    layer1_outputs(6865) <= a xor b;
    layer1_outputs(6866) <= not (a and b);
    layer1_outputs(6867) <= not a or b;
    layer1_outputs(6868) <= a and b;
    layer1_outputs(6869) <= b;
    layer1_outputs(6870) <= not a or b;
    layer1_outputs(6871) <= b;
    layer1_outputs(6872) <= not b;
    layer1_outputs(6873) <= b and not a;
    layer1_outputs(6874) <= a xor b;
    layer1_outputs(6875) <= a;
    layer1_outputs(6876) <= not (a xor b);
    layer1_outputs(6877) <= not a;
    layer1_outputs(6878) <= a;
    layer1_outputs(6879) <= not a or b;
    layer1_outputs(6880) <= not a or b;
    layer1_outputs(6881) <= 1'b1;
    layer1_outputs(6882) <= 1'b0;
    layer1_outputs(6883) <= not b;
    layer1_outputs(6884) <= a and b;
    layer1_outputs(6885) <= b and not a;
    layer1_outputs(6886) <= a and b;
    layer1_outputs(6887) <= a;
    layer1_outputs(6888) <= not a or b;
    layer1_outputs(6889) <= not b or a;
    layer1_outputs(6890) <= b;
    layer1_outputs(6891) <= not a or b;
    layer1_outputs(6892) <= not (a or b);
    layer1_outputs(6893) <= a or b;
    layer1_outputs(6894) <= not a;
    layer1_outputs(6895) <= not (a and b);
    layer1_outputs(6896) <= 1'b0;
    layer1_outputs(6897) <= not a;
    layer1_outputs(6898) <= a;
    layer1_outputs(6899) <= a or b;
    layer1_outputs(6900) <= a or b;
    layer1_outputs(6901) <= 1'b0;
    layer1_outputs(6902) <= a and not b;
    layer1_outputs(6903) <= not a;
    layer1_outputs(6904) <= a xor b;
    layer1_outputs(6905) <= not (a xor b);
    layer1_outputs(6906) <= not a;
    layer1_outputs(6907) <= not a;
    layer1_outputs(6908) <= not a;
    layer1_outputs(6909) <= not (a or b);
    layer1_outputs(6910) <= a and not b;
    layer1_outputs(6911) <= not (a or b);
    layer1_outputs(6912) <= 1'b0;
    layer1_outputs(6913) <= not (a and b);
    layer1_outputs(6914) <= b and not a;
    layer1_outputs(6915) <= not a;
    layer1_outputs(6916) <= not a;
    layer1_outputs(6917) <= not a or b;
    layer1_outputs(6918) <= a;
    layer1_outputs(6919) <= a and b;
    layer1_outputs(6920) <= not a;
    layer1_outputs(6921) <= not (a xor b);
    layer1_outputs(6922) <= b;
    layer1_outputs(6923) <= a and not b;
    layer1_outputs(6924) <= a or b;
    layer1_outputs(6925) <= not b;
    layer1_outputs(6926) <= a xor b;
    layer1_outputs(6927) <= a;
    layer1_outputs(6928) <= b and not a;
    layer1_outputs(6929) <= not (a and b);
    layer1_outputs(6930) <= not a or b;
    layer1_outputs(6931) <= a and not b;
    layer1_outputs(6932) <= a;
    layer1_outputs(6933) <= not (a or b);
    layer1_outputs(6934) <= a or b;
    layer1_outputs(6935) <= b;
    layer1_outputs(6936) <= a;
    layer1_outputs(6937) <= not (a xor b);
    layer1_outputs(6938) <= not a or b;
    layer1_outputs(6939) <= a and not b;
    layer1_outputs(6940) <= b;
    layer1_outputs(6941) <= b and not a;
    layer1_outputs(6942) <= b and not a;
    layer1_outputs(6943) <= b;
    layer1_outputs(6944) <= not b or a;
    layer1_outputs(6945) <= not (a or b);
    layer1_outputs(6946) <= a and b;
    layer1_outputs(6947) <= b;
    layer1_outputs(6948) <= not a;
    layer1_outputs(6949) <= not (a or b);
    layer1_outputs(6950) <= a;
    layer1_outputs(6951) <= b and not a;
    layer1_outputs(6952) <= not b;
    layer1_outputs(6953) <= not a;
    layer1_outputs(6954) <= a;
    layer1_outputs(6955) <= a and b;
    layer1_outputs(6956) <= b;
    layer1_outputs(6957) <= not (a xor b);
    layer1_outputs(6958) <= 1'b1;
    layer1_outputs(6959) <= not a;
    layer1_outputs(6960) <= not a;
    layer1_outputs(6961) <= not b;
    layer1_outputs(6962) <= a or b;
    layer1_outputs(6963) <= not b;
    layer1_outputs(6964) <= a or b;
    layer1_outputs(6965) <= a and b;
    layer1_outputs(6966) <= b;
    layer1_outputs(6967) <= not b;
    layer1_outputs(6968) <= not a or b;
    layer1_outputs(6969) <= a and b;
    layer1_outputs(6970) <= not b or a;
    layer1_outputs(6971) <= 1'b0;
    layer1_outputs(6972) <= a or b;
    layer1_outputs(6973) <= not (a xor b);
    layer1_outputs(6974) <= not (a or b);
    layer1_outputs(6975) <= not b;
    layer1_outputs(6976) <= b and not a;
    layer1_outputs(6977) <= 1'b1;
    layer1_outputs(6978) <= not b or a;
    layer1_outputs(6979) <= b and not a;
    layer1_outputs(6980) <= a and b;
    layer1_outputs(6981) <= b and not a;
    layer1_outputs(6982) <= not a;
    layer1_outputs(6983) <= not b or a;
    layer1_outputs(6984) <= a and b;
    layer1_outputs(6985) <= b and not a;
    layer1_outputs(6986) <= not a or b;
    layer1_outputs(6987) <= a xor b;
    layer1_outputs(6988) <= b;
    layer1_outputs(6989) <= b and not a;
    layer1_outputs(6990) <= not b;
    layer1_outputs(6991) <= not a;
    layer1_outputs(6992) <= not (a xor b);
    layer1_outputs(6993) <= a;
    layer1_outputs(6994) <= 1'b0;
    layer1_outputs(6995) <= not b;
    layer1_outputs(6996) <= not a;
    layer1_outputs(6997) <= a;
    layer1_outputs(6998) <= not b;
    layer1_outputs(6999) <= not (a and b);
    layer1_outputs(7000) <= a;
    layer1_outputs(7001) <= not a;
    layer1_outputs(7002) <= not b or a;
    layer1_outputs(7003) <= not (a xor b);
    layer1_outputs(7004) <= b;
    layer1_outputs(7005) <= b and not a;
    layer1_outputs(7006) <= not a or b;
    layer1_outputs(7007) <= b and not a;
    layer1_outputs(7008) <= 1'b0;
    layer1_outputs(7009) <= a or b;
    layer1_outputs(7010) <= not (a and b);
    layer1_outputs(7011) <= not b;
    layer1_outputs(7012) <= 1'b0;
    layer1_outputs(7013) <= not (a or b);
    layer1_outputs(7014) <= a and b;
    layer1_outputs(7015) <= a;
    layer1_outputs(7016) <= a;
    layer1_outputs(7017) <= a and b;
    layer1_outputs(7018) <= a and b;
    layer1_outputs(7019) <= 1'b1;
    layer1_outputs(7020) <= a xor b;
    layer1_outputs(7021) <= a and b;
    layer1_outputs(7022) <= a and not b;
    layer1_outputs(7023) <= a xor b;
    layer1_outputs(7024) <= b and not a;
    layer1_outputs(7025) <= b and not a;
    layer1_outputs(7026) <= b;
    layer1_outputs(7027) <= not b;
    layer1_outputs(7028) <= not (a and b);
    layer1_outputs(7029) <= a and not b;
    layer1_outputs(7030) <= not (a or b);
    layer1_outputs(7031) <= not (a xor b);
    layer1_outputs(7032) <= b;
    layer1_outputs(7033) <= a;
    layer1_outputs(7034) <= not (a and b);
    layer1_outputs(7035) <= not a or b;
    layer1_outputs(7036) <= not b or a;
    layer1_outputs(7037) <= not a or b;
    layer1_outputs(7038) <= not b;
    layer1_outputs(7039) <= a and b;
    layer1_outputs(7040) <= b and not a;
    layer1_outputs(7041) <= b and not a;
    layer1_outputs(7042) <= not b;
    layer1_outputs(7043) <= not a;
    layer1_outputs(7044) <= a xor b;
    layer1_outputs(7045) <= not a;
    layer1_outputs(7046) <= not (a or b);
    layer1_outputs(7047) <= not (a xor b);
    layer1_outputs(7048) <= a xor b;
    layer1_outputs(7049) <= not (a or b);
    layer1_outputs(7050) <= not (a or b);
    layer1_outputs(7051) <= not b;
    layer1_outputs(7052) <= a and b;
    layer1_outputs(7053) <= not (a xor b);
    layer1_outputs(7054) <= 1'b0;
    layer1_outputs(7055) <= a or b;
    layer1_outputs(7056) <= a;
    layer1_outputs(7057) <= a and b;
    layer1_outputs(7058) <= a;
    layer1_outputs(7059) <= not (a and b);
    layer1_outputs(7060) <= b and not a;
    layer1_outputs(7061) <= a;
    layer1_outputs(7062) <= b and not a;
    layer1_outputs(7063) <= not b;
    layer1_outputs(7064) <= not (a or b);
    layer1_outputs(7065) <= not (a xor b);
    layer1_outputs(7066) <= b;
    layer1_outputs(7067) <= not b;
    layer1_outputs(7068) <= not a or b;
    layer1_outputs(7069) <= not (a or b);
    layer1_outputs(7070) <= b;
    layer1_outputs(7071) <= b;
    layer1_outputs(7072) <= not a or b;
    layer1_outputs(7073) <= a and b;
    layer1_outputs(7074) <= not b;
    layer1_outputs(7075) <= b;
    layer1_outputs(7076) <= not b;
    layer1_outputs(7077) <= not (a and b);
    layer1_outputs(7078) <= not (a xor b);
    layer1_outputs(7079) <= a and b;
    layer1_outputs(7080) <= b;
    layer1_outputs(7081) <= 1'b1;
    layer1_outputs(7082) <= b;
    layer1_outputs(7083) <= a and b;
    layer1_outputs(7084) <= b and not a;
    layer1_outputs(7085) <= not b or a;
    layer1_outputs(7086) <= not b or a;
    layer1_outputs(7087) <= a and not b;
    layer1_outputs(7088) <= not (a and b);
    layer1_outputs(7089) <= not b or a;
    layer1_outputs(7090) <= not a or b;
    layer1_outputs(7091) <= not b;
    layer1_outputs(7092) <= b and not a;
    layer1_outputs(7093) <= not a;
    layer1_outputs(7094) <= not b or a;
    layer1_outputs(7095) <= a or b;
    layer1_outputs(7096) <= a and b;
    layer1_outputs(7097) <= b;
    layer1_outputs(7098) <= not (a xor b);
    layer1_outputs(7099) <= not b or a;
    layer1_outputs(7100) <= a or b;
    layer1_outputs(7101) <= 1'b1;
    layer1_outputs(7102) <= a;
    layer1_outputs(7103) <= a and b;
    layer1_outputs(7104) <= not b;
    layer1_outputs(7105) <= a and not b;
    layer1_outputs(7106) <= a or b;
    layer1_outputs(7107) <= not a or b;
    layer1_outputs(7108) <= a;
    layer1_outputs(7109) <= 1'b0;
    layer1_outputs(7110) <= b;
    layer1_outputs(7111) <= b and not a;
    layer1_outputs(7112) <= not a;
    layer1_outputs(7113) <= a;
    layer1_outputs(7114) <= a;
    layer1_outputs(7115) <= a and not b;
    layer1_outputs(7116) <= not a;
    layer1_outputs(7117) <= not a or b;
    layer1_outputs(7118) <= not b;
    layer1_outputs(7119) <= b;
    layer1_outputs(7120) <= not b;
    layer1_outputs(7121) <= a or b;
    layer1_outputs(7122) <= a and not b;
    layer1_outputs(7123) <= a xor b;
    layer1_outputs(7124) <= not (a and b);
    layer1_outputs(7125) <= not a;
    layer1_outputs(7126) <= a and not b;
    layer1_outputs(7127) <= a and b;
    layer1_outputs(7128) <= a xor b;
    layer1_outputs(7129) <= a;
    layer1_outputs(7130) <= 1'b0;
    layer1_outputs(7131) <= not a or b;
    layer1_outputs(7132) <= a xor b;
    layer1_outputs(7133) <= a or b;
    layer1_outputs(7134) <= 1'b0;
    layer1_outputs(7135) <= b;
    layer1_outputs(7136) <= a and b;
    layer1_outputs(7137) <= 1'b0;
    layer1_outputs(7138) <= b;
    layer1_outputs(7139) <= a and not b;
    layer1_outputs(7140) <= a xor b;
    layer1_outputs(7141) <= a xor b;
    layer1_outputs(7142) <= a or b;
    layer1_outputs(7143) <= a and not b;
    layer1_outputs(7144) <= not a or b;
    layer1_outputs(7145) <= b;
    layer1_outputs(7146) <= b;
    layer1_outputs(7147) <= a and not b;
    layer1_outputs(7148) <= not (a or b);
    layer1_outputs(7149) <= 1'b0;
    layer1_outputs(7150) <= a or b;
    layer1_outputs(7151) <= not (a and b);
    layer1_outputs(7152) <= not b or a;
    layer1_outputs(7153) <= a;
    layer1_outputs(7154) <= b;
    layer1_outputs(7155) <= not (a and b);
    layer1_outputs(7156) <= not a or b;
    layer1_outputs(7157) <= a or b;
    layer1_outputs(7158) <= a xor b;
    layer1_outputs(7159) <= not (a or b);
    layer1_outputs(7160) <= a;
    layer1_outputs(7161) <= not (a xor b);
    layer1_outputs(7162) <= a xor b;
    layer1_outputs(7163) <= a and b;
    layer1_outputs(7164) <= not (a and b);
    layer1_outputs(7165) <= b;
    layer1_outputs(7166) <= not a or b;
    layer1_outputs(7167) <= not (a or b);
    layer1_outputs(7168) <= not (a xor b);
    layer1_outputs(7169) <= 1'b0;
    layer1_outputs(7170) <= b;
    layer1_outputs(7171) <= b and not a;
    layer1_outputs(7172) <= not (a and b);
    layer1_outputs(7173) <= b and not a;
    layer1_outputs(7174) <= not a;
    layer1_outputs(7175) <= not a or b;
    layer1_outputs(7176) <= not (a and b);
    layer1_outputs(7177) <= a or b;
    layer1_outputs(7178) <= b and not a;
    layer1_outputs(7179) <= not a;
    layer1_outputs(7180) <= 1'b1;
    layer1_outputs(7181) <= not b;
    layer1_outputs(7182) <= a or b;
    layer1_outputs(7183) <= not b;
    layer1_outputs(7184) <= not (a or b);
    layer1_outputs(7185) <= a xor b;
    layer1_outputs(7186) <= b;
    layer1_outputs(7187) <= a or b;
    layer1_outputs(7188) <= a or b;
    layer1_outputs(7189) <= not (a and b);
    layer1_outputs(7190) <= not b or a;
    layer1_outputs(7191) <= a and not b;
    layer1_outputs(7192) <= not (a or b);
    layer1_outputs(7193) <= not a;
    layer1_outputs(7194) <= a and not b;
    layer1_outputs(7195) <= a and not b;
    layer1_outputs(7196) <= not (a xor b);
    layer1_outputs(7197) <= a;
    layer1_outputs(7198) <= a;
    layer1_outputs(7199) <= not (a or b);
    layer1_outputs(7200) <= a;
    layer1_outputs(7201) <= not (a and b);
    layer1_outputs(7202) <= not b or a;
    layer1_outputs(7203) <= not b or a;
    layer1_outputs(7204) <= not b or a;
    layer1_outputs(7205) <= b and not a;
    layer1_outputs(7206) <= 1'b1;
    layer1_outputs(7207) <= not (a xor b);
    layer1_outputs(7208) <= 1'b0;
    layer1_outputs(7209) <= a and b;
    layer1_outputs(7210) <= a;
    layer1_outputs(7211) <= not (a xor b);
    layer1_outputs(7212) <= not (a and b);
    layer1_outputs(7213) <= 1'b1;
    layer1_outputs(7214) <= not (a or b);
    layer1_outputs(7215) <= a;
    layer1_outputs(7216) <= not a;
    layer1_outputs(7217) <= not a or b;
    layer1_outputs(7218) <= b and not a;
    layer1_outputs(7219) <= not a;
    layer1_outputs(7220) <= b and not a;
    layer1_outputs(7221) <= not (a xor b);
    layer1_outputs(7222) <= not (a or b);
    layer1_outputs(7223) <= a or b;
    layer1_outputs(7224) <= a and not b;
    layer1_outputs(7225) <= not a;
    layer1_outputs(7226) <= not a;
    layer1_outputs(7227) <= not b;
    layer1_outputs(7228) <= not a;
    layer1_outputs(7229) <= a;
    layer1_outputs(7230) <= not a;
    layer1_outputs(7231) <= b;
    layer1_outputs(7232) <= a or b;
    layer1_outputs(7233) <= 1'b0;
    layer1_outputs(7234) <= not (a and b);
    layer1_outputs(7235) <= a or b;
    layer1_outputs(7236) <= b;
    layer1_outputs(7237) <= 1'b1;
    layer1_outputs(7238) <= not (a and b);
    layer1_outputs(7239) <= a;
    layer1_outputs(7240) <= a;
    layer1_outputs(7241) <= not b;
    layer1_outputs(7242) <= a and not b;
    layer1_outputs(7243) <= not a;
    layer1_outputs(7244) <= a;
    layer1_outputs(7245) <= not b or a;
    layer1_outputs(7246) <= b and not a;
    layer1_outputs(7247) <= 1'b0;
    layer1_outputs(7248) <= not b or a;
    layer1_outputs(7249) <= b;
    layer1_outputs(7250) <= b;
    layer1_outputs(7251) <= not b or a;
    layer1_outputs(7252) <= b;
    layer1_outputs(7253) <= a;
    layer1_outputs(7254) <= a;
    layer1_outputs(7255) <= 1'b1;
    layer1_outputs(7256) <= 1'b0;
    layer1_outputs(7257) <= a or b;
    layer1_outputs(7258) <= 1'b1;
    layer1_outputs(7259) <= a or b;
    layer1_outputs(7260) <= not b;
    layer1_outputs(7261) <= not (a or b);
    layer1_outputs(7262) <= not a or b;
    layer1_outputs(7263) <= a and b;
    layer1_outputs(7264) <= a;
    layer1_outputs(7265) <= a or b;
    layer1_outputs(7266) <= b;
    layer1_outputs(7267) <= not (a and b);
    layer1_outputs(7268) <= not (a or b);
    layer1_outputs(7269) <= a or b;
    layer1_outputs(7270) <= 1'b0;
    layer1_outputs(7271) <= not (a and b);
    layer1_outputs(7272) <= a xor b;
    layer1_outputs(7273) <= not (a or b);
    layer1_outputs(7274) <= a xor b;
    layer1_outputs(7275) <= not b or a;
    layer1_outputs(7276) <= not a or b;
    layer1_outputs(7277) <= not (a or b);
    layer1_outputs(7278) <= b;
    layer1_outputs(7279) <= not b or a;
    layer1_outputs(7280) <= b;
    layer1_outputs(7281) <= not a or b;
    layer1_outputs(7282) <= b and not a;
    layer1_outputs(7283) <= a;
    layer1_outputs(7284) <= not b or a;
    layer1_outputs(7285) <= a or b;
    layer1_outputs(7286) <= b and not a;
    layer1_outputs(7287) <= not (a and b);
    layer1_outputs(7288) <= not (a xor b);
    layer1_outputs(7289) <= a or b;
    layer1_outputs(7290) <= a or b;
    layer1_outputs(7291) <= not (a xor b);
    layer1_outputs(7292) <= not (a and b);
    layer1_outputs(7293) <= b;
    layer1_outputs(7294) <= not b;
    layer1_outputs(7295) <= not b;
    layer1_outputs(7296) <= not (a or b);
    layer1_outputs(7297) <= not (a or b);
    layer1_outputs(7298) <= not a or b;
    layer1_outputs(7299) <= not (a and b);
    layer1_outputs(7300) <= not b or a;
    layer1_outputs(7301) <= not (a and b);
    layer1_outputs(7302) <= a xor b;
    layer1_outputs(7303) <= not b or a;
    layer1_outputs(7304) <= b and not a;
    layer1_outputs(7305) <= a and not b;
    layer1_outputs(7306) <= 1'b0;
    layer1_outputs(7307) <= b;
    layer1_outputs(7308) <= 1'b1;
    layer1_outputs(7309) <= a xor b;
    layer1_outputs(7310) <= b;
    layer1_outputs(7311) <= not a;
    layer1_outputs(7312) <= 1'b0;
    layer1_outputs(7313) <= b;
    layer1_outputs(7314) <= not a or b;
    layer1_outputs(7315) <= not (a xor b);
    layer1_outputs(7316) <= not b or a;
    layer1_outputs(7317) <= a and not b;
    layer1_outputs(7318) <= a;
    layer1_outputs(7319) <= a;
    layer1_outputs(7320) <= not a or b;
    layer1_outputs(7321) <= a;
    layer1_outputs(7322) <= a and not b;
    layer1_outputs(7323) <= a or b;
    layer1_outputs(7324) <= 1'b0;
    layer1_outputs(7325) <= not (a or b);
    layer1_outputs(7326) <= a or b;
    layer1_outputs(7327) <= not b or a;
    layer1_outputs(7328) <= b and not a;
    layer1_outputs(7329) <= not a;
    layer1_outputs(7330) <= b and not a;
    layer1_outputs(7331) <= not a or b;
    layer1_outputs(7332) <= a xor b;
    layer1_outputs(7333) <= not b;
    layer1_outputs(7334) <= not (a xor b);
    layer1_outputs(7335) <= b and not a;
    layer1_outputs(7336) <= a xor b;
    layer1_outputs(7337) <= b;
    layer1_outputs(7338) <= not a or b;
    layer1_outputs(7339) <= a;
    layer1_outputs(7340) <= a and b;
    layer1_outputs(7341) <= a;
    layer1_outputs(7342) <= not b or a;
    layer1_outputs(7343) <= not (a xor b);
    layer1_outputs(7344) <= not (a and b);
    layer1_outputs(7345) <= a or b;
    layer1_outputs(7346) <= not (a xor b);
    layer1_outputs(7347) <= not a or b;
    layer1_outputs(7348) <= not b or a;
    layer1_outputs(7349) <= a or b;
    layer1_outputs(7350) <= not b;
    layer1_outputs(7351) <= not b;
    layer1_outputs(7352) <= not (a and b);
    layer1_outputs(7353) <= b;
    layer1_outputs(7354) <= a and b;
    layer1_outputs(7355) <= 1'b0;
    layer1_outputs(7356) <= not (a and b);
    layer1_outputs(7357) <= b;
    layer1_outputs(7358) <= not (a or b);
    layer1_outputs(7359) <= not b or a;
    layer1_outputs(7360) <= b;
    layer1_outputs(7361) <= a or b;
    layer1_outputs(7362) <= 1'b0;
    layer1_outputs(7363) <= a;
    layer1_outputs(7364) <= not (a or b);
    layer1_outputs(7365) <= a xor b;
    layer1_outputs(7366) <= a;
    layer1_outputs(7367) <= not (a and b);
    layer1_outputs(7368) <= a and b;
    layer1_outputs(7369) <= b and not a;
    layer1_outputs(7370) <= not a;
    layer1_outputs(7371) <= a;
    layer1_outputs(7372) <= a xor b;
    layer1_outputs(7373) <= a or b;
    layer1_outputs(7374) <= a and not b;
    layer1_outputs(7375) <= b;
    layer1_outputs(7376) <= a;
    layer1_outputs(7377) <= b;
    layer1_outputs(7378) <= not b or a;
    layer1_outputs(7379) <= not a or b;
    layer1_outputs(7380) <= not (a xor b);
    layer1_outputs(7381) <= b;
    layer1_outputs(7382) <= not (a and b);
    layer1_outputs(7383) <= b;
    layer1_outputs(7384) <= not b;
    layer1_outputs(7385) <= a or b;
    layer1_outputs(7386) <= 1'b1;
    layer1_outputs(7387) <= a and not b;
    layer1_outputs(7388) <= not b;
    layer1_outputs(7389) <= a;
    layer1_outputs(7390) <= not (a xor b);
    layer1_outputs(7391) <= not b or a;
    layer1_outputs(7392) <= not (a xor b);
    layer1_outputs(7393) <= a or b;
    layer1_outputs(7394) <= a and b;
    layer1_outputs(7395) <= not b;
    layer1_outputs(7396) <= a;
    layer1_outputs(7397) <= b and not a;
    layer1_outputs(7398) <= a and not b;
    layer1_outputs(7399) <= a or b;
    layer1_outputs(7400) <= b;
    layer1_outputs(7401) <= not b or a;
    layer1_outputs(7402) <= not b;
    layer1_outputs(7403) <= not b;
    layer1_outputs(7404) <= b and not a;
    layer1_outputs(7405) <= not (a or b);
    layer1_outputs(7406) <= not (a and b);
    layer1_outputs(7407) <= a;
    layer1_outputs(7408) <= not a;
    layer1_outputs(7409) <= not a or b;
    layer1_outputs(7410) <= a;
    layer1_outputs(7411) <= not (a or b);
    layer1_outputs(7412) <= 1'b0;
    layer1_outputs(7413) <= a or b;
    layer1_outputs(7414) <= b;
    layer1_outputs(7415) <= 1'b1;
    layer1_outputs(7416) <= not (a xor b);
    layer1_outputs(7417) <= not (a and b);
    layer1_outputs(7418) <= a and not b;
    layer1_outputs(7419) <= b;
    layer1_outputs(7420) <= a or b;
    layer1_outputs(7421) <= a;
    layer1_outputs(7422) <= a;
    layer1_outputs(7423) <= a and not b;
    layer1_outputs(7424) <= not (a and b);
    layer1_outputs(7425) <= not b;
    layer1_outputs(7426) <= 1'b0;
    layer1_outputs(7427) <= a and not b;
    layer1_outputs(7428) <= not (a and b);
    layer1_outputs(7429) <= not b;
    layer1_outputs(7430) <= not b or a;
    layer1_outputs(7431) <= not b;
    layer1_outputs(7432) <= not b;
    layer1_outputs(7433) <= 1'b1;
    layer1_outputs(7434) <= not a;
    layer1_outputs(7435) <= not b or a;
    layer1_outputs(7436) <= a or b;
    layer1_outputs(7437) <= not a or b;
    layer1_outputs(7438) <= a or b;
    layer1_outputs(7439) <= not b or a;
    layer1_outputs(7440) <= b;
    layer1_outputs(7441) <= a and b;
    layer1_outputs(7442) <= not a;
    layer1_outputs(7443) <= not b;
    layer1_outputs(7444) <= a or b;
    layer1_outputs(7445) <= not b;
    layer1_outputs(7446) <= not a or b;
    layer1_outputs(7447) <= not (a or b);
    layer1_outputs(7448) <= a or b;
    layer1_outputs(7449) <= a or b;
    layer1_outputs(7450) <= not b;
    layer1_outputs(7451) <= not b or a;
    layer1_outputs(7452) <= not (a xor b);
    layer1_outputs(7453) <= not b or a;
    layer1_outputs(7454) <= a and b;
    layer1_outputs(7455) <= not (a and b);
    layer1_outputs(7456) <= not b or a;
    layer1_outputs(7457) <= not a;
    layer1_outputs(7458) <= not (a xor b);
    layer1_outputs(7459) <= a;
    layer1_outputs(7460) <= a xor b;
    layer1_outputs(7461) <= not b;
    layer1_outputs(7462) <= b and not a;
    layer1_outputs(7463) <= not a;
    layer1_outputs(7464) <= a and b;
    layer1_outputs(7465) <= not b;
    layer1_outputs(7466) <= not a or b;
    layer1_outputs(7467) <= not a;
    layer1_outputs(7468) <= a xor b;
    layer1_outputs(7469) <= not b;
    layer1_outputs(7470) <= 1'b0;
    layer1_outputs(7471) <= b;
    layer1_outputs(7472) <= a;
    layer1_outputs(7473) <= b;
    layer1_outputs(7474) <= not a;
    layer1_outputs(7475) <= b and not a;
    layer1_outputs(7476) <= not a;
    layer1_outputs(7477) <= not a;
    layer1_outputs(7478) <= not b;
    layer1_outputs(7479) <= a xor b;
    layer1_outputs(7480) <= not a;
    layer1_outputs(7481) <= not b;
    layer1_outputs(7482) <= 1'b1;
    layer1_outputs(7483) <= a and b;
    layer1_outputs(7484) <= a or b;
    layer1_outputs(7485) <= a and b;
    layer1_outputs(7486) <= b and not a;
    layer1_outputs(7487) <= a and b;
    layer1_outputs(7488) <= a or b;
    layer1_outputs(7489) <= not b;
    layer1_outputs(7490) <= not (a or b);
    layer1_outputs(7491) <= a and b;
    layer1_outputs(7492) <= not (a or b);
    layer1_outputs(7493) <= not (a xor b);
    layer1_outputs(7494) <= not b;
    layer1_outputs(7495) <= not (a xor b);
    layer1_outputs(7496) <= a or b;
    layer1_outputs(7497) <= not a;
    layer1_outputs(7498) <= a;
    layer1_outputs(7499) <= not a;
    layer1_outputs(7500) <= b and not a;
    layer1_outputs(7501) <= 1'b0;
    layer1_outputs(7502) <= not b or a;
    layer1_outputs(7503) <= not a;
    layer1_outputs(7504) <= not a;
    layer1_outputs(7505) <= not b;
    layer1_outputs(7506) <= not b;
    layer1_outputs(7507) <= not a;
    layer1_outputs(7508) <= b and not a;
    layer1_outputs(7509) <= a;
    layer1_outputs(7510) <= not a;
    layer1_outputs(7511) <= a and not b;
    layer1_outputs(7512) <= not (a and b);
    layer1_outputs(7513) <= a or b;
    layer1_outputs(7514) <= b;
    layer1_outputs(7515) <= not (a or b);
    layer1_outputs(7516) <= a and b;
    layer1_outputs(7517) <= b;
    layer1_outputs(7518) <= not b;
    layer1_outputs(7519) <= a and b;
    layer1_outputs(7520) <= a;
    layer1_outputs(7521) <= a;
    layer1_outputs(7522) <= a and b;
    layer1_outputs(7523) <= b;
    layer1_outputs(7524) <= 1'b1;
    layer1_outputs(7525) <= a;
    layer1_outputs(7526) <= not a;
    layer1_outputs(7527) <= a and not b;
    layer1_outputs(7528) <= b and not a;
    layer1_outputs(7529) <= not a or b;
    layer1_outputs(7530) <= b;
    layer1_outputs(7531) <= not a;
    layer1_outputs(7532) <= not a or b;
    layer1_outputs(7533) <= a xor b;
    layer1_outputs(7534) <= not a or b;
    layer1_outputs(7535) <= a or b;
    layer1_outputs(7536) <= a;
    layer1_outputs(7537) <= not (a and b);
    layer1_outputs(7538) <= not (a xor b);
    layer1_outputs(7539) <= a xor b;
    layer1_outputs(7540) <= a and b;
    layer1_outputs(7541) <= a or b;
    layer1_outputs(7542) <= not b;
    layer1_outputs(7543) <= not b;
    layer1_outputs(7544) <= not b or a;
    layer1_outputs(7545) <= not b or a;
    layer1_outputs(7546) <= not (a or b);
    layer1_outputs(7547) <= a or b;
    layer1_outputs(7548) <= a;
    layer1_outputs(7549) <= not (a xor b);
    layer1_outputs(7550) <= not a;
    layer1_outputs(7551) <= not (a or b);
    layer1_outputs(7552) <= not (a xor b);
    layer1_outputs(7553) <= not (a or b);
    layer1_outputs(7554) <= not (a and b);
    layer1_outputs(7555) <= not a;
    layer1_outputs(7556) <= a or b;
    layer1_outputs(7557) <= not a;
    layer1_outputs(7558) <= a and b;
    layer1_outputs(7559) <= not b;
    layer1_outputs(7560) <= a or b;
    layer1_outputs(7561) <= not b;
    layer1_outputs(7562) <= not (a and b);
    layer1_outputs(7563) <= b and not a;
    layer1_outputs(7564) <= not b;
    layer1_outputs(7565) <= b;
    layer1_outputs(7566) <= not (a xor b);
    layer1_outputs(7567) <= not (a or b);
    layer1_outputs(7568) <= a or b;
    layer1_outputs(7569) <= not a or b;
    layer1_outputs(7570) <= not a;
    layer1_outputs(7571) <= a and b;
    layer1_outputs(7572) <= not a;
    layer1_outputs(7573) <= a;
    layer1_outputs(7574) <= a or b;
    layer1_outputs(7575) <= not a;
    layer1_outputs(7576) <= not (a and b);
    layer1_outputs(7577) <= 1'b0;
    layer1_outputs(7578) <= not b;
    layer1_outputs(7579) <= not a or b;
    layer1_outputs(7580) <= a;
    layer1_outputs(7581) <= a;
    layer1_outputs(7582) <= b;
    layer1_outputs(7583) <= a or b;
    layer1_outputs(7584) <= a;
    layer1_outputs(7585) <= 1'b0;
    layer1_outputs(7586) <= not a or b;
    layer1_outputs(7587) <= b;
    layer1_outputs(7588) <= not b or a;
    layer1_outputs(7589) <= not b;
    layer1_outputs(7590) <= not a;
    layer1_outputs(7591) <= a;
    layer1_outputs(7592) <= b and not a;
    layer1_outputs(7593) <= a and b;
    layer1_outputs(7594) <= not b;
    layer1_outputs(7595) <= not (a or b);
    layer1_outputs(7596) <= not a;
    layer1_outputs(7597) <= not b;
    layer1_outputs(7598) <= not b;
    layer1_outputs(7599) <= b;
    layer1_outputs(7600) <= a;
    layer1_outputs(7601) <= 1'b0;
    layer1_outputs(7602) <= a;
    layer1_outputs(7603) <= not (a or b);
    layer1_outputs(7604) <= not b or a;
    layer1_outputs(7605) <= not b or a;
    layer1_outputs(7606) <= not a;
    layer1_outputs(7607) <= a;
    layer1_outputs(7608) <= not (a and b);
    layer1_outputs(7609) <= b;
    layer1_outputs(7610) <= not (a or b);
    layer1_outputs(7611) <= b and not a;
    layer1_outputs(7612) <= not (a and b);
    layer1_outputs(7613) <= 1'b1;
    layer1_outputs(7614) <= a;
    layer1_outputs(7615) <= a;
    layer1_outputs(7616) <= not b;
    layer1_outputs(7617) <= b and not a;
    layer1_outputs(7618) <= a and b;
    layer1_outputs(7619) <= a or b;
    layer1_outputs(7620) <= not a;
    layer1_outputs(7621) <= b;
    layer1_outputs(7622) <= a and b;
    layer1_outputs(7623) <= not a;
    layer1_outputs(7624) <= a xor b;
    layer1_outputs(7625) <= b and not a;
    layer1_outputs(7626) <= a and b;
    layer1_outputs(7627) <= a;
    layer1_outputs(7628) <= not (a or b);
    layer1_outputs(7629) <= a and b;
    layer1_outputs(7630) <= b and not a;
    layer1_outputs(7631) <= b;
    layer1_outputs(7632) <= 1'b1;
    layer1_outputs(7633) <= not b;
    layer1_outputs(7634) <= not b;
    layer1_outputs(7635) <= a xor b;
    layer1_outputs(7636) <= not a or b;
    layer1_outputs(7637) <= not (a and b);
    layer1_outputs(7638) <= a and b;
    layer1_outputs(7639) <= a or b;
    layer1_outputs(7640) <= not (a or b);
    layer1_outputs(7641) <= not (a and b);
    layer1_outputs(7642) <= not (a xor b);
    layer1_outputs(7643) <= not b;
    layer1_outputs(7644) <= b;
    layer1_outputs(7645) <= not b or a;
    layer1_outputs(7646) <= not b;
    layer1_outputs(7647) <= a or b;
    layer1_outputs(7648) <= 1'b0;
    layer1_outputs(7649) <= not (a xor b);
    layer1_outputs(7650) <= a and not b;
    layer1_outputs(7651) <= a or b;
    layer1_outputs(7652) <= 1'b0;
    layer1_outputs(7653) <= 1'b1;
    layer1_outputs(7654) <= a;
    layer1_outputs(7655) <= a;
    layer1_outputs(7656) <= a and not b;
    layer1_outputs(7657) <= b;
    layer1_outputs(7658) <= not b;
    layer1_outputs(7659) <= 1'b0;
    layer1_outputs(7660) <= not b or a;
    layer1_outputs(7661) <= a and not b;
    layer1_outputs(7662) <= not a or b;
    layer1_outputs(7663) <= not (a or b);
    layer1_outputs(7664) <= not b or a;
    layer1_outputs(7665) <= a or b;
    layer1_outputs(7666) <= not b;
    layer1_outputs(7667) <= a and not b;
    layer1_outputs(7668) <= b;
    layer1_outputs(7669) <= not b;
    layer1_outputs(7670) <= a and not b;
    layer1_outputs(7671) <= b;
    layer1_outputs(7672) <= 1'b1;
    layer1_outputs(7673) <= not a;
    layer1_outputs(7674) <= not b;
    layer1_outputs(7675) <= not (a or b);
    layer1_outputs(7676) <= not (a and b);
    layer1_outputs(7677) <= not a or b;
    layer1_outputs(7678) <= a or b;
    layer1_outputs(7679) <= a and b;
    layer1_outputs(7680) <= a and b;
    layer1_outputs(7681) <= b and not a;
    layer1_outputs(7682) <= a;
    layer1_outputs(7683) <= a and b;
    layer1_outputs(7684) <= not (a or b);
    layer1_outputs(7685) <= a;
    layer1_outputs(7686) <= not b;
    layer1_outputs(7687) <= b;
    layer1_outputs(7688) <= a xor b;
    layer1_outputs(7689) <= not (a or b);
    layer1_outputs(7690) <= not b or a;
    layer1_outputs(7691) <= not b or a;
    layer1_outputs(7692) <= not a or b;
    layer1_outputs(7693) <= not (a and b);
    layer1_outputs(7694) <= 1'b0;
    layer1_outputs(7695) <= 1'b1;
    layer1_outputs(7696) <= a or b;
    layer1_outputs(7697) <= not a;
    layer1_outputs(7698) <= a or b;
    layer1_outputs(7699) <= 1'b0;
    layer1_outputs(7700) <= not (a and b);
    layer1_outputs(7701) <= not (a and b);
    layer1_outputs(7702) <= a;
    layer1_outputs(7703) <= a and b;
    layer1_outputs(7704) <= a and not b;
    layer1_outputs(7705) <= a or b;
    layer1_outputs(7706) <= not (a xor b);
    layer1_outputs(7707) <= not (a and b);
    layer1_outputs(7708) <= not b;
    layer1_outputs(7709) <= not (a and b);
    layer1_outputs(7710) <= not a;
    layer1_outputs(7711) <= b;
    layer1_outputs(7712) <= not b or a;
    layer1_outputs(7713) <= a xor b;
    layer1_outputs(7714) <= not (a and b);
    layer1_outputs(7715) <= a or b;
    layer1_outputs(7716) <= not b;
    layer1_outputs(7717) <= not (a and b);
    layer1_outputs(7718) <= not a or b;
    layer1_outputs(7719) <= not a or b;
    layer1_outputs(7720) <= not (a xor b);
    layer1_outputs(7721) <= b;
    layer1_outputs(7722) <= not b or a;
    layer1_outputs(7723) <= not a or b;
    layer1_outputs(7724) <= not b;
    layer1_outputs(7725) <= b and not a;
    layer1_outputs(7726) <= not b;
    layer1_outputs(7727) <= a or b;
    layer1_outputs(7728) <= not a or b;
    layer1_outputs(7729) <= not a;
    layer1_outputs(7730) <= not b;
    layer1_outputs(7731) <= a and b;
    layer1_outputs(7732) <= b;
    layer1_outputs(7733) <= b and not a;
    layer1_outputs(7734) <= not a or b;
    layer1_outputs(7735) <= not b;
    layer1_outputs(7736) <= not b or a;
    layer1_outputs(7737) <= not b or a;
    layer1_outputs(7738) <= not b;
    layer1_outputs(7739) <= not b or a;
    layer1_outputs(7740) <= b and not a;
    layer1_outputs(7741) <= 1'b1;
    layer1_outputs(7742) <= not (a and b);
    layer1_outputs(7743) <= not (a xor b);
    layer1_outputs(7744) <= 1'b0;
    layer1_outputs(7745) <= 1'b0;
    layer1_outputs(7746) <= not b;
    layer1_outputs(7747) <= b and not a;
    layer1_outputs(7748) <= a and not b;
    layer1_outputs(7749) <= not (a and b);
    layer1_outputs(7750) <= 1'b0;
    layer1_outputs(7751) <= 1'b1;
    layer1_outputs(7752) <= not a;
    layer1_outputs(7753) <= 1'b1;
    layer1_outputs(7754) <= not (a xor b);
    layer1_outputs(7755) <= b and not a;
    layer1_outputs(7756) <= not (a and b);
    layer1_outputs(7757) <= a;
    layer1_outputs(7758) <= 1'b0;
    layer1_outputs(7759) <= not (a and b);
    layer1_outputs(7760) <= not (a and b);
    layer1_outputs(7761) <= not b;
    layer1_outputs(7762) <= 1'b0;
    layer1_outputs(7763) <= not a or b;
    layer1_outputs(7764) <= not (a or b);
    layer1_outputs(7765) <= not a or b;
    layer1_outputs(7766) <= a and b;
    layer1_outputs(7767) <= a and not b;
    layer1_outputs(7768) <= b and not a;
    layer1_outputs(7769) <= a xor b;
    layer1_outputs(7770) <= not a or b;
    layer1_outputs(7771) <= not b or a;
    layer1_outputs(7772) <= 1'b0;
    layer1_outputs(7773) <= a xor b;
    layer1_outputs(7774) <= not b;
    layer1_outputs(7775) <= not b;
    layer1_outputs(7776) <= a and not b;
    layer1_outputs(7777) <= a and b;
    layer1_outputs(7778) <= a or b;
    layer1_outputs(7779) <= not b;
    layer1_outputs(7780) <= not (a and b);
    layer1_outputs(7781) <= not a;
    layer1_outputs(7782) <= 1'b0;
    layer1_outputs(7783) <= not b;
    layer1_outputs(7784) <= a or b;
    layer1_outputs(7785) <= b and not a;
    layer1_outputs(7786) <= not (a and b);
    layer1_outputs(7787) <= not a or b;
    layer1_outputs(7788) <= not a or b;
    layer1_outputs(7789) <= not b;
    layer1_outputs(7790) <= a and b;
    layer1_outputs(7791) <= not a or b;
    layer1_outputs(7792) <= not (a xor b);
    layer1_outputs(7793) <= a;
    layer1_outputs(7794) <= a and b;
    layer1_outputs(7795) <= not b;
    layer1_outputs(7796) <= a and b;
    layer1_outputs(7797) <= not b;
    layer1_outputs(7798) <= not a or b;
    layer1_outputs(7799) <= not b;
    layer1_outputs(7800) <= a and not b;
    layer1_outputs(7801) <= b;
    layer1_outputs(7802) <= b;
    layer1_outputs(7803) <= not b or a;
    layer1_outputs(7804) <= not a or b;
    layer1_outputs(7805) <= not b;
    layer1_outputs(7806) <= b;
    layer1_outputs(7807) <= not (a or b);
    layer1_outputs(7808) <= not a or b;
    layer1_outputs(7809) <= a;
    layer1_outputs(7810) <= not (a or b);
    layer1_outputs(7811) <= a and not b;
    layer1_outputs(7812) <= a xor b;
    layer1_outputs(7813) <= not b or a;
    layer1_outputs(7814) <= b;
    layer1_outputs(7815) <= not b;
    layer1_outputs(7816) <= not b;
    layer1_outputs(7817) <= not (a and b);
    layer1_outputs(7818) <= a and not b;
    layer1_outputs(7819) <= a xor b;
    layer1_outputs(7820) <= a and b;
    layer1_outputs(7821) <= a xor b;
    layer1_outputs(7822) <= b;
    layer1_outputs(7823) <= b;
    layer1_outputs(7824) <= 1'b0;
    layer1_outputs(7825) <= not (a or b);
    layer1_outputs(7826) <= not (a or b);
    layer1_outputs(7827) <= b;
    layer1_outputs(7828) <= not a or b;
    layer1_outputs(7829) <= not a or b;
    layer1_outputs(7830) <= not a or b;
    layer1_outputs(7831) <= a and not b;
    layer1_outputs(7832) <= b and not a;
    layer1_outputs(7833) <= not (a and b);
    layer1_outputs(7834) <= not b or a;
    layer1_outputs(7835) <= not b or a;
    layer1_outputs(7836) <= a and b;
    layer1_outputs(7837) <= not b or a;
    layer1_outputs(7838) <= a xor b;
    layer1_outputs(7839) <= a;
    layer1_outputs(7840) <= not a;
    layer1_outputs(7841) <= a;
    layer1_outputs(7842) <= 1'b1;
    layer1_outputs(7843) <= not (a or b);
    layer1_outputs(7844) <= not (a or b);
    layer1_outputs(7845) <= a xor b;
    layer1_outputs(7846) <= not b;
    layer1_outputs(7847) <= a;
    layer1_outputs(7848) <= b and not a;
    layer1_outputs(7849) <= a;
    layer1_outputs(7850) <= not a;
    layer1_outputs(7851) <= a or b;
    layer1_outputs(7852) <= b and not a;
    layer1_outputs(7853) <= not a or b;
    layer1_outputs(7854) <= not a or b;
    layer1_outputs(7855) <= not a or b;
    layer1_outputs(7856) <= a or b;
    layer1_outputs(7857) <= a and b;
    layer1_outputs(7858) <= not b or a;
    layer1_outputs(7859) <= not (a or b);
    layer1_outputs(7860) <= a;
    layer1_outputs(7861) <= not (a and b);
    layer1_outputs(7862) <= not a or b;
    layer1_outputs(7863) <= not (a and b);
    layer1_outputs(7864) <= a and b;
    layer1_outputs(7865) <= not b or a;
    layer1_outputs(7866) <= not b;
    layer1_outputs(7867) <= b and not a;
    layer1_outputs(7868) <= a xor b;
    layer1_outputs(7869) <= 1'b1;
    layer1_outputs(7870) <= not a or b;
    layer1_outputs(7871) <= not b or a;
    layer1_outputs(7872) <= not (a xor b);
    layer1_outputs(7873) <= not b;
    layer1_outputs(7874) <= not b;
    layer1_outputs(7875) <= not (a or b);
    layer1_outputs(7876) <= b;
    layer1_outputs(7877) <= a or b;
    layer1_outputs(7878) <= b and not a;
    layer1_outputs(7879) <= a and not b;
    layer1_outputs(7880) <= not a or b;
    layer1_outputs(7881) <= a xor b;
    layer1_outputs(7882) <= not (a or b);
    layer1_outputs(7883) <= not a;
    layer1_outputs(7884) <= a and not b;
    layer1_outputs(7885) <= 1'b1;
    layer1_outputs(7886) <= not a or b;
    layer1_outputs(7887) <= a and not b;
    layer1_outputs(7888) <= not a or b;
    layer1_outputs(7889) <= a;
    layer1_outputs(7890) <= not b;
    layer1_outputs(7891) <= a;
    layer1_outputs(7892) <= a and b;
    layer1_outputs(7893) <= not (a and b);
    layer1_outputs(7894) <= not a;
    layer1_outputs(7895) <= not (a and b);
    layer1_outputs(7896) <= not a or b;
    layer1_outputs(7897) <= 1'b1;
    layer1_outputs(7898) <= not b;
    layer1_outputs(7899) <= not b or a;
    layer1_outputs(7900) <= not (a or b);
    layer1_outputs(7901) <= not (a or b);
    layer1_outputs(7902) <= not (a and b);
    layer1_outputs(7903) <= not b;
    layer1_outputs(7904) <= 1'b0;
    layer1_outputs(7905) <= a;
    layer1_outputs(7906) <= not b;
    layer1_outputs(7907) <= a;
    layer1_outputs(7908) <= not a;
    layer1_outputs(7909) <= not a or b;
    layer1_outputs(7910) <= not a;
    layer1_outputs(7911) <= not a;
    layer1_outputs(7912) <= not b or a;
    layer1_outputs(7913) <= not a;
    layer1_outputs(7914) <= not (a and b);
    layer1_outputs(7915) <= b;
    layer1_outputs(7916) <= not b or a;
    layer1_outputs(7917) <= not b or a;
    layer1_outputs(7918) <= b;
    layer1_outputs(7919) <= not (a and b);
    layer1_outputs(7920) <= b and not a;
    layer1_outputs(7921) <= a or b;
    layer1_outputs(7922) <= a xor b;
    layer1_outputs(7923) <= not (a or b);
    layer1_outputs(7924) <= b;
    layer1_outputs(7925) <= not b;
    layer1_outputs(7926) <= a or b;
    layer1_outputs(7927) <= a and b;
    layer1_outputs(7928) <= a and b;
    layer1_outputs(7929) <= a xor b;
    layer1_outputs(7930) <= 1'b0;
    layer1_outputs(7931) <= a;
    layer1_outputs(7932) <= not a or b;
    layer1_outputs(7933) <= a;
    layer1_outputs(7934) <= not (a or b);
    layer1_outputs(7935) <= a and b;
    layer1_outputs(7936) <= not a or b;
    layer1_outputs(7937) <= a and not b;
    layer1_outputs(7938) <= not (a or b);
    layer1_outputs(7939) <= b;
    layer1_outputs(7940) <= a xor b;
    layer1_outputs(7941) <= a xor b;
    layer1_outputs(7942) <= not (a and b);
    layer1_outputs(7943) <= b and not a;
    layer1_outputs(7944) <= not b;
    layer1_outputs(7945) <= not (a and b);
    layer1_outputs(7946) <= not a;
    layer1_outputs(7947) <= 1'b0;
    layer1_outputs(7948) <= not a or b;
    layer1_outputs(7949) <= a and b;
    layer1_outputs(7950) <= a xor b;
    layer1_outputs(7951) <= not b or a;
    layer1_outputs(7952) <= not b;
    layer1_outputs(7953) <= not b or a;
    layer1_outputs(7954) <= a and not b;
    layer1_outputs(7955) <= not a;
    layer1_outputs(7956) <= a or b;
    layer1_outputs(7957) <= not b;
    layer1_outputs(7958) <= not (a and b);
    layer1_outputs(7959) <= b;
    layer1_outputs(7960) <= a xor b;
    layer1_outputs(7961) <= not a or b;
    layer1_outputs(7962) <= a and b;
    layer1_outputs(7963) <= a xor b;
    layer1_outputs(7964) <= a or b;
    layer1_outputs(7965) <= 1'b1;
    layer1_outputs(7966) <= b;
    layer1_outputs(7967) <= not (a or b);
    layer1_outputs(7968) <= a;
    layer1_outputs(7969) <= a;
    layer1_outputs(7970) <= not a;
    layer1_outputs(7971) <= a and b;
    layer1_outputs(7972) <= b;
    layer1_outputs(7973) <= not a;
    layer1_outputs(7974) <= a or b;
    layer1_outputs(7975) <= b and not a;
    layer1_outputs(7976) <= a or b;
    layer1_outputs(7977) <= a and b;
    layer1_outputs(7978) <= a;
    layer1_outputs(7979) <= a or b;
    layer1_outputs(7980) <= not (a or b);
    layer1_outputs(7981) <= b;
    layer1_outputs(7982) <= not a;
    layer1_outputs(7983) <= b and not a;
    layer1_outputs(7984) <= not (a or b);
    layer1_outputs(7985) <= not (a and b);
    layer1_outputs(7986) <= a;
    layer1_outputs(7987) <= not (a xor b);
    layer1_outputs(7988) <= not a or b;
    layer1_outputs(7989) <= not a;
    layer1_outputs(7990) <= a and b;
    layer1_outputs(7991) <= not a or b;
    layer1_outputs(7992) <= not b;
    layer1_outputs(7993) <= not a;
    layer1_outputs(7994) <= a;
    layer1_outputs(7995) <= not b or a;
    layer1_outputs(7996) <= not b;
    layer1_outputs(7997) <= not (a xor b);
    layer1_outputs(7998) <= a;
    layer1_outputs(7999) <= not b or a;
    layer1_outputs(8000) <= not b;
    layer1_outputs(8001) <= not a;
    layer1_outputs(8002) <= not a or b;
    layer1_outputs(8003) <= not a or b;
    layer1_outputs(8004) <= b and not a;
    layer1_outputs(8005) <= a;
    layer1_outputs(8006) <= not a;
    layer1_outputs(8007) <= a or b;
    layer1_outputs(8008) <= not b or a;
    layer1_outputs(8009) <= not (a and b);
    layer1_outputs(8010) <= not (a and b);
    layer1_outputs(8011) <= a or b;
    layer1_outputs(8012) <= not a;
    layer1_outputs(8013) <= not (a xor b);
    layer1_outputs(8014) <= not (a or b);
    layer1_outputs(8015) <= not a or b;
    layer1_outputs(8016) <= not a;
    layer1_outputs(8017) <= not (a and b);
    layer1_outputs(8018) <= not b or a;
    layer1_outputs(8019) <= not (a xor b);
    layer1_outputs(8020) <= 1'b1;
    layer1_outputs(8021) <= a or b;
    layer1_outputs(8022) <= b and not a;
    layer1_outputs(8023) <= not (a xor b);
    layer1_outputs(8024) <= b and not a;
    layer1_outputs(8025) <= a xor b;
    layer1_outputs(8026) <= a xor b;
    layer1_outputs(8027) <= not b;
    layer1_outputs(8028) <= not a;
    layer1_outputs(8029) <= not b;
    layer1_outputs(8030) <= not b;
    layer1_outputs(8031) <= a and b;
    layer1_outputs(8032) <= not b or a;
    layer1_outputs(8033) <= a;
    layer1_outputs(8034) <= not a;
    layer1_outputs(8035) <= not (a or b);
    layer1_outputs(8036) <= not a or b;
    layer1_outputs(8037) <= not b or a;
    layer1_outputs(8038) <= b;
    layer1_outputs(8039) <= not (a and b);
    layer1_outputs(8040) <= not b;
    layer1_outputs(8041) <= not b;
    layer1_outputs(8042) <= a and not b;
    layer1_outputs(8043) <= not b;
    layer1_outputs(8044) <= a;
    layer1_outputs(8045) <= a or b;
    layer1_outputs(8046) <= a xor b;
    layer1_outputs(8047) <= not (a or b);
    layer1_outputs(8048) <= b;
    layer1_outputs(8049) <= a;
    layer1_outputs(8050) <= not (a xor b);
    layer1_outputs(8051) <= not a;
    layer1_outputs(8052) <= not a or b;
    layer1_outputs(8053) <= not (a and b);
    layer1_outputs(8054) <= not a or b;
    layer1_outputs(8055) <= not b or a;
    layer1_outputs(8056) <= not b;
    layer1_outputs(8057) <= b;
    layer1_outputs(8058) <= b;
    layer1_outputs(8059) <= not (a and b);
    layer1_outputs(8060) <= b and not a;
    layer1_outputs(8061) <= not b or a;
    layer1_outputs(8062) <= 1'b0;
    layer1_outputs(8063) <= a and not b;
    layer1_outputs(8064) <= a and b;
    layer1_outputs(8065) <= not a;
    layer1_outputs(8066) <= not b or a;
    layer1_outputs(8067) <= b and not a;
    layer1_outputs(8068) <= a;
    layer1_outputs(8069) <= a and b;
    layer1_outputs(8070) <= not a or b;
    layer1_outputs(8071) <= a;
    layer1_outputs(8072) <= a and b;
    layer1_outputs(8073) <= a or b;
    layer1_outputs(8074) <= not (a and b);
    layer1_outputs(8075) <= a;
    layer1_outputs(8076) <= not (a xor b);
    layer1_outputs(8077) <= b;
    layer1_outputs(8078) <= a and not b;
    layer1_outputs(8079) <= not b;
    layer1_outputs(8080) <= 1'b0;
    layer1_outputs(8081) <= not a or b;
    layer1_outputs(8082) <= 1'b1;
    layer1_outputs(8083) <= 1'b1;
    layer1_outputs(8084) <= a or b;
    layer1_outputs(8085) <= b;
    layer1_outputs(8086) <= a and b;
    layer1_outputs(8087) <= not a;
    layer1_outputs(8088) <= b and not a;
    layer1_outputs(8089) <= not a;
    layer1_outputs(8090) <= a or b;
    layer1_outputs(8091) <= not (a xor b);
    layer1_outputs(8092) <= b and not a;
    layer1_outputs(8093) <= not a or b;
    layer1_outputs(8094) <= b and not a;
    layer1_outputs(8095) <= a xor b;
    layer1_outputs(8096) <= not b;
    layer1_outputs(8097) <= not (a and b);
    layer1_outputs(8098) <= a or b;
    layer1_outputs(8099) <= not (a and b);
    layer1_outputs(8100) <= a and b;
    layer1_outputs(8101) <= a;
    layer1_outputs(8102) <= a and not b;
    layer1_outputs(8103) <= not a;
    layer1_outputs(8104) <= not a or b;
    layer1_outputs(8105) <= not a;
    layer1_outputs(8106) <= not a;
    layer1_outputs(8107) <= a;
    layer1_outputs(8108) <= not b or a;
    layer1_outputs(8109) <= 1'b1;
    layer1_outputs(8110) <= not b or a;
    layer1_outputs(8111) <= a and not b;
    layer1_outputs(8112) <= a and not b;
    layer1_outputs(8113) <= not b;
    layer1_outputs(8114) <= not a;
    layer1_outputs(8115) <= not (a or b);
    layer1_outputs(8116) <= not (a or b);
    layer1_outputs(8117) <= not b or a;
    layer1_outputs(8118) <= a and not b;
    layer1_outputs(8119) <= a;
    layer1_outputs(8120) <= a xor b;
    layer1_outputs(8121) <= a and b;
    layer1_outputs(8122) <= a or b;
    layer1_outputs(8123) <= not a;
    layer1_outputs(8124) <= a;
    layer1_outputs(8125) <= a and b;
    layer1_outputs(8126) <= a;
    layer1_outputs(8127) <= b;
    layer1_outputs(8128) <= not (a or b);
    layer1_outputs(8129) <= not (a and b);
    layer1_outputs(8130) <= 1'b1;
    layer1_outputs(8131) <= not b;
    layer1_outputs(8132) <= a xor b;
    layer1_outputs(8133) <= b;
    layer1_outputs(8134) <= a and b;
    layer1_outputs(8135) <= not (a xor b);
    layer1_outputs(8136) <= 1'b1;
    layer1_outputs(8137) <= not a or b;
    layer1_outputs(8138) <= not b or a;
    layer1_outputs(8139) <= not (a xor b);
    layer1_outputs(8140) <= a;
    layer1_outputs(8141) <= a xor b;
    layer1_outputs(8142) <= a;
    layer1_outputs(8143) <= not b or a;
    layer1_outputs(8144) <= not (a and b);
    layer1_outputs(8145) <= a and not b;
    layer1_outputs(8146) <= 1'b0;
    layer1_outputs(8147) <= not a;
    layer1_outputs(8148) <= not (a xor b);
    layer1_outputs(8149) <= b and not a;
    layer1_outputs(8150) <= a or b;
    layer1_outputs(8151) <= not (a or b);
    layer1_outputs(8152) <= a;
    layer1_outputs(8153) <= not a;
    layer1_outputs(8154) <= b;
    layer1_outputs(8155) <= not (a and b);
    layer1_outputs(8156) <= not (a or b);
    layer1_outputs(8157) <= not (a xor b);
    layer1_outputs(8158) <= not b;
    layer1_outputs(8159) <= 1'b0;
    layer1_outputs(8160) <= not b or a;
    layer1_outputs(8161) <= not (a and b);
    layer1_outputs(8162) <= not (a xor b);
    layer1_outputs(8163) <= not a or b;
    layer1_outputs(8164) <= a;
    layer1_outputs(8165) <= not (a or b);
    layer1_outputs(8166) <= not a;
    layer1_outputs(8167) <= not a;
    layer1_outputs(8168) <= a and b;
    layer1_outputs(8169) <= a and not b;
    layer1_outputs(8170) <= a xor b;
    layer1_outputs(8171) <= not (a or b);
    layer1_outputs(8172) <= not b;
    layer1_outputs(8173) <= a and b;
    layer1_outputs(8174) <= b and not a;
    layer1_outputs(8175) <= a and b;
    layer1_outputs(8176) <= not a or b;
    layer1_outputs(8177) <= not b;
    layer1_outputs(8178) <= not a;
    layer1_outputs(8179) <= b;
    layer1_outputs(8180) <= 1'b0;
    layer1_outputs(8181) <= not b;
    layer1_outputs(8182) <= 1'b1;
    layer1_outputs(8183) <= b;
    layer1_outputs(8184) <= not b or a;
    layer1_outputs(8185) <= a and b;
    layer1_outputs(8186) <= b and not a;
    layer1_outputs(8187) <= not (a or b);
    layer1_outputs(8188) <= not b;
    layer1_outputs(8189) <= not (a or b);
    layer1_outputs(8190) <= not a or b;
    layer1_outputs(8191) <= a;
    layer1_outputs(8192) <= b;
    layer1_outputs(8193) <= 1'b1;
    layer1_outputs(8194) <= a or b;
    layer1_outputs(8195) <= b;
    layer1_outputs(8196) <= not a;
    layer1_outputs(8197) <= a and not b;
    layer1_outputs(8198) <= a or b;
    layer1_outputs(8199) <= a;
    layer1_outputs(8200) <= not a;
    layer1_outputs(8201) <= b and not a;
    layer1_outputs(8202) <= b;
    layer1_outputs(8203) <= a and not b;
    layer1_outputs(8204) <= a and not b;
    layer1_outputs(8205) <= not (a xor b);
    layer1_outputs(8206) <= a and not b;
    layer1_outputs(8207) <= not a;
    layer1_outputs(8208) <= not (a or b);
    layer1_outputs(8209) <= not b;
    layer1_outputs(8210) <= a xor b;
    layer1_outputs(8211) <= not a or b;
    layer1_outputs(8212) <= not b;
    layer1_outputs(8213) <= a and not b;
    layer1_outputs(8214) <= not b;
    layer1_outputs(8215) <= 1'b1;
    layer1_outputs(8216) <= b and not a;
    layer1_outputs(8217) <= a or b;
    layer1_outputs(8218) <= not (a or b);
    layer1_outputs(8219) <= not a;
    layer1_outputs(8220) <= b and not a;
    layer1_outputs(8221) <= a and b;
    layer1_outputs(8222) <= a;
    layer1_outputs(8223) <= a;
    layer1_outputs(8224) <= b;
    layer1_outputs(8225) <= a and b;
    layer1_outputs(8226) <= a and not b;
    layer1_outputs(8227) <= a or b;
    layer1_outputs(8228) <= a and b;
    layer1_outputs(8229) <= not (a or b);
    layer1_outputs(8230) <= a and b;
    layer1_outputs(8231) <= not (a xor b);
    layer1_outputs(8232) <= not b;
    layer1_outputs(8233) <= not b;
    layer1_outputs(8234) <= b;
    layer1_outputs(8235) <= b and not a;
    layer1_outputs(8236) <= a;
    layer1_outputs(8237) <= b;
    layer1_outputs(8238) <= not a or b;
    layer1_outputs(8239) <= a or b;
    layer1_outputs(8240) <= a or b;
    layer1_outputs(8241) <= not b;
    layer1_outputs(8242) <= not b or a;
    layer1_outputs(8243) <= b;
    layer1_outputs(8244) <= b;
    layer1_outputs(8245) <= a and not b;
    layer1_outputs(8246) <= not (a xor b);
    layer1_outputs(8247) <= a and not b;
    layer1_outputs(8248) <= a and b;
    layer1_outputs(8249) <= 1'b0;
    layer1_outputs(8250) <= b;
    layer1_outputs(8251) <= 1'b0;
    layer1_outputs(8252) <= a xor b;
    layer1_outputs(8253) <= a and b;
    layer1_outputs(8254) <= not (a or b);
    layer1_outputs(8255) <= a and b;
    layer1_outputs(8256) <= not (a and b);
    layer1_outputs(8257) <= not b;
    layer1_outputs(8258) <= a and not b;
    layer1_outputs(8259) <= a;
    layer1_outputs(8260) <= b and not a;
    layer1_outputs(8261) <= b and not a;
    layer1_outputs(8262) <= a or b;
    layer1_outputs(8263) <= not a;
    layer1_outputs(8264) <= not b or a;
    layer1_outputs(8265) <= a;
    layer1_outputs(8266) <= a and b;
    layer1_outputs(8267) <= a;
    layer1_outputs(8268) <= not a;
    layer1_outputs(8269) <= 1'b0;
    layer1_outputs(8270) <= 1'b0;
    layer1_outputs(8271) <= a and not b;
    layer1_outputs(8272) <= not (a or b);
    layer1_outputs(8273) <= not a;
    layer1_outputs(8274) <= a;
    layer1_outputs(8275) <= a;
    layer1_outputs(8276) <= b;
    layer1_outputs(8277) <= not (a or b);
    layer1_outputs(8278) <= a;
    layer1_outputs(8279) <= a or b;
    layer1_outputs(8280) <= 1'b1;
    layer1_outputs(8281) <= a and b;
    layer1_outputs(8282) <= not (a or b);
    layer1_outputs(8283) <= not b or a;
    layer1_outputs(8284) <= not (a or b);
    layer1_outputs(8285) <= a;
    layer1_outputs(8286) <= not (a or b);
    layer1_outputs(8287) <= not a;
    layer1_outputs(8288) <= a and b;
    layer1_outputs(8289) <= not a or b;
    layer1_outputs(8290) <= not b;
    layer1_outputs(8291) <= b and not a;
    layer1_outputs(8292) <= not b or a;
    layer1_outputs(8293) <= 1'b1;
    layer1_outputs(8294) <= a xor b;
    layer1_outputs(8295) <= not a or b;
    layer1_outputs(8296) <= not (a or b);
    layer1_outputs(8297) <= a;
    layer1_outputs(8298) <= not b;
    layer1_outputs(8299) <= a and not b;
    layer1_outputs(8300) <= not (a xor b);
    layer1_outputs(8301) <= not a or b;
    layer1_outputs(8302) <= a;
    layer1_outputs(8303) <= not (a and b);
    layer1_outputs(8304) <= a;
    layer1_outputs(8305) <= b and not a;
    layer1_outputs(8306) <= a;
    layer1_outputs(8307) <= a and not b;
    layer1_outputs(8308) <= not a;
    layer1_outputs(8309) <= not a;
    layer1_outputs(8310) <= b and not a;
    layer1_outputs(8311) <= not b;
    layer1_outputs(8312) <= b and not a;
    layer1_outputs(8313) <= not b;
    layer1_outputs(8314) <= a and b;
    layer1_outputs(8315) <= a;
    layer1_outputs(8316) <= a or b;
    layer1_outputs(8317) <= not (a or b);
    layer1_outputs(8318) <= a and not b;
    layer1_outputs(8319) <= not a or b;
    layer1_outputs(8320) <= not (a and b);
    layer1_outputs(8321) <= not (a and b);
    layer1_outputs(8322) <= b;
    layer1_outputs(8323) <= b;
    layer1_outputs(8324) <= not a;
    layer1_outputs(8325) <= not a or b;
    layer1_outputs(8326) <= b;
    layer1_outputs(8327) <= not (a xor b);
    layer1_outputs(8328) <= not b or a;
    layer1_outputs(8329) <= not (a xor b);
    layer1_outputs(8330) <= b;
    layer1_outputs(8331) <= not a;
    layer1_outputs(8332) <= a;
    layer1_outputs(8333) <= not a;
    layer1_outputs(8334) <= not a or b;
    layer1_outputs(8335) <= 1'b0;
    layer1_outputs(8336) <= a;
    layer1_outputs(8337) <= b and not a;
    layer1_outputs(8338) <= a and b;
    layer1_outputs(8339) <= a and not b;
    layer1_outputs(8340) <= not b;
    layer1_outputs(8341) <= not (a or b);
    layer1_outputs(8342) <= a or b;
    layer1_outputs(8343) <= not a or b;
    layer1_outputs(8344) <= a xor b;
    layer1_outputs(8345) <= not a;
    layer1_outputs(8346) <= a or b;
    layer1_outputs(8347) <= a;
    layer1_outputs(8348) <= 1'b0;
    layer1_outputs(8349) <= not b or a;
    layer1_outputs(8350) <= b and not a;
    layer1_outputs(8351) <= a xor b;
    layer1_outputs(8352) <= a and b;
    layer1_outputs(8353) <= not (a xor b);
    layer1_outputs(8354) <= 1'b1;
    layer1_outputs(8355) <= a xor b;
    layer1_outputs(8356) <= a xor b;
    layer1_outputs(8357) <= not a or b;
    layer1_outputs(8358) <= b;
    layer1_outputs(8359) <= a;
    layer1_outputs(8360) <= not a or b;
    layer1_outputs(8361) <= not b or a;
    layer1_outputs(8362) <= 1'b1;
    layer1_outputs(8363) <= a xor b;
    layer1_outputs(8364) <= not b;
    layer1_outputs(8365) <= not a or b;
    layer1_outputs(8366) <= not a;
    layer1_outputs(8367) <= a;
    layer1_outputs(8368) <= a and not b;
    layer1_outputs(8369) <= a and not b;
    layer1_outputs(8370) <= 1'b1;
    layer1_outputs(8371) <= not (a xor b);
    layer1_outputs(8372) <= b and not a;
    layer1_outputs(8373) <= a xor b;
    layer1_outputs(8374) <= not b;
    layer1_outputs(8375) <= not b or a;
    layer1_outputs(8376) <= 1'b1;
    layer1_outputs(8377) <= not a;
    layer1_outputs(8378) <= not b;
    layer1_outputs(8379) <= not (a and b);
    layer1_outputs(8380) <= not a or b;
    layer1_outputs(8381) <= b and not a;
    layer1_outputs(8382) <= a xor b;
    layer1_outputs(8383) <= a and b;
    layer1_outputs(8384) <= b;
    layer1_outputs(8385) <= 1'b0;
    layer1_outputs(8386) <= not a or b;
    layer1_outputs(8387) <= 1'b1;
    layer1_outputs(8388) <= not (a xor b);
    layer1_outputs(8389) <= b and not a;
    layer1_outputs(8390) <= not b;
    layer1_outputs(8391) <= b and not a;
    layer1_outputs(8392) <= a or b;
    layer1_outputs(8393) <= not (a or b);
    layer1_outputs(8394) <= not (a and b);
    layer1_outputs(8395) <= not a or b;
    layer1_outputs(8396) <= 1'b1;
    layer1_outputs(8397) <= not (a and b);
    layer1_outputs(8398) <= a and not b;
    layer1_outputs(8399) <= not a;
    layer1_outputs(8400) <= a xor b;
    layer1_outputs(8401) <= a;
    layer1_outputs(8402) <= not b;
    layer1_outputs(8403) <= not a;
    layer1_outputs(8404) <= not (a and b);
    layer1_outputs(8405) <= not a;
    layer1_outputs(8406) <= not a;
    layer1_outputs(8407) <= a and not b;
    layer1_outputs(8408) <= not b or a;
    layer1_outputs(8409) <= b;
    layer1_outputs(8410) <= a;
    layer1_outputs(8411) <= 1'b0;
    layer1_outputs(8412) <= not b or a;
    layer1_outputs(8413) <= not b;
    layer1_outputs(8414) <= not (a or b);
    layer1_outputs(8415) <= a and b;
    layer1_outputs(8416) <= not (a xor b);
    layer1_outputs(8417) <= 1'b1;
    layer1_outputs(8418) <= not a or b;
    layer1_outputs(8419) <= a and b;
    layer1_outputs(8420) <= not b or a;
    layer1_outputs(8421) <= a xor b;
    layer1_outputs(8422) <= not a;
    layer1_outputs(8423) <= not a;
    layer1_outputs(8424) <= not (a and b);
    layer1_outputs(8425) <= not (a and b);
    layer1_outputs(8426) <= not b or a;
    layer1_outputs(8427) <= not (a and b);
    layer1_outputs(8428) <= not (a or b);
    layer1_outputs(8429) <= b and not a;
    layer1_outputs(8430) <= not (a or b);
    layer1_outputs(8431) <= not b;
    layer1_outputs(8432) <= not a;
    layer1_outputs(8433) <= not (a or b);
    layer1_outputs(8434) <= 1'b1;
    layer1_outputs(8435) <= a and b;
    layer1_outputs(8436) <= not b;
    layer1_outputs(8437) <= not (a and b);
    layer1_outputs(8438) <= not (a or b);
    layer1_outputs(8439) <= 1'b1;
    layer1_outputs(8440) <= not (a and b);
    layer1_outputs(8441) <= a and b;
    layer1_outputs(8442) <= a and not b;
    layer1_outputs(8443) <= not (a or b);
    layer1_outputs(8444) <= not (a and b);
    layer1_outputs(8445) <= not (a or b);
    layer1_outputs(8446) <= b;
    layer1_outputs(8447) <= not b or a;
    layer1_outputs(8448) <= not b;
    layer1_outputs(8449) <= a;
    layer1_outputs(8450) <= a;
    layer1_outputs(8451) <= not (a or b);
    layer1_outputs(8452) <= not a;
    layer1_outputs(8453) <= b and not a;
    layer1_outputs(8454) <= not (a and b);
    layer1_outputs(8455) <= 1'b1;
    layer1_outputs(8456) <= not a;
    layer1_outputs(8457) <= not a or b;
    layer1_outputs(8458) <= not (a and b);
    layer1_outputs(8459) <= a;
    layer1_outputs(8460) <= not (a and b);
    layer1_outputs(8461) <= not a;
    layer1_outputs(8462) <= not a;
    layer1_outputs(8463) <= a and b;
    layer1_outputs(8464) <= not b or a;
    layer1_outputs(8465) <= not (a xor b);
    layer1_outputs(8466) <= not a or b;
    layer1_outputs(8467) <= a;
    layer1_outputs(8468) <= b;
    layer1_outputs(8469) <= not b;
    layer1_outputs(8470) <= not b or a;
    layer1_outputs(8471) <= not b;
    layer1_outputs(8472) <= not (a xor b);
    layer1_outputs(8473) <= a and not b;
    layer1_outputs(8474) <= not b or a;
    layer1_outputs(8475) <= a or b;
    layer1_outputs(8476) <= not b;
    layer1_outputs(8477) <= not (a or b);
    layer1_outputs(8478) <= 1'b0;
    layer1_outputs(8479) <= not b;
    layer1_outputs(8480) <= not a or b;
    layer1_outputs(8481) <= a xor b;
    layer1_outputs(8482) <= a and b;
    layer1_outputs(8483) <= b;
    layer1_outputs(8484) <= not a;
    layer1_outputs(8485) <= a or b;
    layer1_outputs(8486) <= a;
    layer1_outputs(8487) <= not a or b;
    layer1_outputs(8488) <= not a or b;
    layer1_outputs(8489) <= b;
    layer1_outputs(8490) <= b and not a;
    layer1_outputs(8491) <= not (a and b);
    layer1_outputs(8492) <= a or b;
    layer1_outputs(8493) <= a and not b;
    layer1_outputs(8494) <= not b;
    layer1_outputs(8495) <= a or b;
    layer1_outputs(8496) <= not (a or b);
    layer1_outputs(8497) <= not a or b;
    layer1_outputs(8498) <= 1'b1;
    layer1_outputs(8499) <= not b;
    layer1_outputs(8500) <= a or b;
    layer1_outputs(8501) <= a and b;
    layer1_outputs(8502) <= not b;
    layer1_outputs(8503) <= a and b;
    layer1_outputs(8504) <= not (a xor b);
    layer1_outputs(8505) <= not (a or b);
    layer1_outputs(8506) <= not (a or b);
    layer1_outputs(8507) <= not (a xor b);
    layer1_outputs(8508) <= b;
    layer1_outputs(8509) <= not (a xor b);
    layer1_outputs(8510) <= b and not a;
    layer1_outputs(8511) <= a and not b;
    layer1_outputs(8512) <= not a or b;
    layer1_outputs(8513) <= not a or b;
    layer1_outputs(8514) <= not b;
    layer1_outputs(8515) <= not a;
    layer1_outputs(8516) <= a;
    layer1_outputs(8517) <= b and not a;
    layer1_outputs(8518) <= b and not a;
    layer1_outputs(8519) <= b;
    layer1_outputs(8520) <= not b or a;
    layer1_outputs(8521) <= a xor b;
    layer1_outputs(8522) <= not (a or b);
    layer1_outputs(8523) <= a and not b;
    layer1_outputs(8524) <= a xor b;
    layer1_outputs(8525) <= a xor b;
    layer1_outputs(8526) <= not a or b;
    layer1_outputs(8527) <= not a;
    layer1_outputs(8528) <= b;
    layer1_outputs(8529) <= not b;
    layer1_outputs(8530) <= not b or a;
    layer1_outputs(8531) <= a or b;
    layer1_outputs(8532) <= not b;
    layer1_outputs(8533) <= a and not b;
    layer1_outputs(8534) <= not (a or b);
    layer1_outputs(8535) <= 1'b1;
    layer1_outputs(8536) <= not a or b;
    layer1_outputs(8537) <= a;
    layer1_outputs(8538) <= not b;
    layer1_outputs(8539) <= not a or b;
    layer1_outputs(8540) <= not (a and b);
    layer1_outputs(8541) <= not (a and b);
    layer1_outputs(8542) <= b;
    layer1_outputs(8543) <= not b;
    layer1_outputs(8544) <= not b or a;
    layer1_outputs(8545) <= not (a or b);
    layer1_outputs(8546) <= a or b;
    layer1_outputs(8547) <= a or b;
    layer1_outputs(8548) <= not b or a;
    layer1_outputs(8549) <= 1'b1;
    layer1_outputs(8550) <= not (a xor b);
    layer1_outputs(8551) <= not b;
    layer1_outputs(8552) <= a and not b;
    layer1_outputs(8553) <= b;
    layer1_outputs(8554) <= a;
    layer1_outputs(8555) <= a and b;
    layer1_outputs(8556) <= not (a or b);
    layer1_outputs(8557) <= not b or a;
    layer1_outputs(8558) <= not (a xor b);
    layer1_outputs(8559) <= b;
    layer1_outputs(8560) <= a and not b;
    layer1_outputs(8561) <= not a;
    layer1_outputs(8562) <= b and not a;
    layer1_outputs(8563) <= not b;
    layer1_outputs(8564) <= not b;
    layer1_outputs(8565) <= 1'b0;
    layer1_outputs(8566) <= not (a or b);
    layer1_outputs(8567) <= not b or a;
    layer1_outputs(8568) <= b and not a;
    layer1_outputs(8569) <= not a;
    layer1_outputs(8570) <= not a or b;
    layer1_outputs(8571) <= not (a xor b);
    layer1_outputs(8572) <= not a or b;
    layer1_outputs(8573) <= b and not a;
    layer1_outputs(8574) <= a;
    layer1_outputs(8575) <= a and b;
    layer1_outputs(8576) <= not a;
    layer1_outputs(8577) <= b;
    layer1_outputs(8578) <= not b;
    layer1_outputs(8579) <= a or b;
    layer1_outputs(8580) <= a;
    layer1_outputs(8581) <= not (a and b);
    layer1_outputs(8582) <= a;
    layer1_outputs(8583) <= a or b;
    layer1_outputs(8584) <= a and not b;
    layer1_outputs(8585) <= b and not a;
    layer1_outputs(8586) <= a;
    layer1_outputs(8587) <= not b;
    layer1_outputs(8588) <= a or b;
    layer1_outputs(8589) <= a;
    layer1_outputs(8590) <= not b or a;
    layer1_outputs(8591) <= not a or b;
    layer1_outputs(8592) <= not a or b;
    layer1_outputs(8593) <= a and not b;
    layer1_outputs(8594) <= a and b;
    layer1_outputs(8595) <= a;
    layer1_outputs(8596) <= not b or a;
    layer1_outputs(8597) <= b;
    layer1_outputs(8598) <= not b;
    layer1_outputs(8599) <= not a;
    layer1_outputs(8600) <= a and not b;
    layer1_outputs(8601) <= a and not b;
    layer1_outputs(8602) <= a xor b;
    layer1_outputs(8603) <= b;
    layer1_outputs(8604) <= a xor b;
    layer1_outputs(8605) <= not b or a;
    layer1_outputs(8606) <= not (a and b);
    layer1_outputs(8607) <= not a or b;
    layer1_outputs(8608) <= not (a or b);
    layer1_outputs(8609) <= b;
    layer1_outputs(8610) <= not (a or b);
    layer1_outputs(8611) <= not (a and b);
    layer1_outputs(8612) <= not b;
    layer1_outputs(8613) <= not b;
    layer1_outputs(8614) <= b and not a;
    layer1_outputs(8615) <= a xor b;
    layer1_outputs(8616) <= not (a xor b);
    layer1_outputs(8617) <= not a;
    layer1_outputs(8618) <= 1'b1;
    layer1_outputs(8619) <= not a;
    layer1_outputs(8620) <= a and not b;
    layer1_outputs(8621) <= not a;
    layer1_outputs(8622) <= not b or a;
    layer1_outputs(8623) <= not (a or b);
    layer1_outputs(8624) <= not (a or b);
    layer1_outputs(8625) <= not (a xor b);
    layer1_outputs(8626) <= not (a or b);
    layer1_outputs(8627) <= a and b;
    layer1_outputs(8628) <= a or b;
    layer1_outputs(8629) <= a or b;
    layer1_outputs(8630) <= a;
    layer1_outputs(8631) <= not a;
    layer1_outputs(8632) <= not (a and b);
    layer1_outputs(8633) <= not b;
    layer1_outputs(8634) <= a xor b;
    layer1_outputs(8635) <= a and b;
    layer1_outputs(8636) <= a and b;
    layer1_outputs(8637) <= not (a or b);
    layer1_outputs(8638) <= b and not a;
    layer1_outputs(8639) <= 1'b1;
    layer1_outputs(8640) <= not b;
    layer1_outputs(8641) <= not b;
    layer1_outputs(8642) <= a xor b;
    layer1_outputs(8643) <= not (a and b);
    layer1_outputs(8644) <= 1'b0;
    layer1_outputs(8645) <= a and b;
    layer1_outputs(8646) <= not a or b;
    layer1_outputs(8647) <= a and not b;
    layer1_outputs(8648) <= b and not a;
    layer1_outputs(8649) <= b and not a;
    layer1_outputs(8650) <= a or b;
    layer1_outputs(8651) <= not b;
    layer1_outputs(8652) <= not a;
    layer1_outputs(8653) <= not a or b;
    layer1_outputs(8654) <= not b or a;
    layer1_outputs(8655) <= a;
    layer1_outputs(8656) <= b and not a;
    layer1_outputs(8657) <= not b;
    layer1_outputs(8658) <= a and not b;
    layer1_outputs(8659) <= a and not b;
    layer1_outputs(8660) <= b;
    layer1_outputs(8661) <= 1'b1;
    layer1_outputs(8662) <= not a or b;
    layer1_outputs(8663) <= a and not b;
    layer1_outputs(8664) <= a or b;
    layer1_outputs(8665) <= not a;
    layer1_outputs(8666) <= b;
    layer1_outputs(8667) <= not b or a;
    layer1_outputs(8668) <= b;
    layer1_outputs(8669) <= not a;
    layer1_outputs(8670) <= a and b;
    layer1_outputs(8671) <= a or b;
    layer1_outputs(8672) <= not a or b;
    layer1_outputs(8673) <= not (a or b);
    layer1_outputs(8674) <= not (a or b);
    layer1_outputs(8675) <= a and not b;
    layer1_outputs(8676) <= not b;
    layer1_outputs(8677) <= not b;
    layer1_outputs(8678) <= not a;
    layer1_outputs(8679) <= a and b;
    layer1_outputs(8680) <= a and not b;
    layer1_outputs(8681) <= a xor b;
    layer1_outputs(8682) <= b;
    layer1_outputs(8683) <= a and b;
    layer1_outputs(8684) <= a and not b;
    layer1_outputs(8685) <= not a;
    layer1_outputs(8686) <= not (a or b);
    layer1_outputs(8687) <= not (a or b);
    layer1_outputs(8688) <= a xor b;
    layer1_outputs(8689) <= not a;
    layer1_outputs(8690) <= a or b;
    layer1_outputs(8691) <= a;
    layer1_outputs(8692) <= b;
    layer1_outputs(8693) <= not b or a;
    layer1_outputs(8694) <= not (a and b);
    layer1_outputs(8695) <= not b or a;
    layer1_outputs(8696) <= not a or b;
    layer1_outputs(8697) <= not (a or b);
    layer1_outputs(8698) <= 1'b1;
    layer1_outputs(8699) <= a or b;
    layer1_outputs(8700) <= not (a or b);
    layer1_outputs(8701) <= not (a and b);
    layer1_outputs(8702) <= 1'b1;
    layer1_outputs(8703) <= a xor b;
    layer1_outputs(8704) <= a or b;
    layer1_outputs(8705) <= b;
    layer1_outputs(8706) <= not a or b;
    layer1_outputs(8707) <= b;
    layer1_outputs(8708) <= not b or a;
    layer1_outputs(8709) <= 1'b1;
    layer1_outputs(8710) <= b;
    layer1_outputs(8711) <= a and not b;
    layer1_outputs(8712) <= not (a and b);
    layer1_outputs(8713) <= not a;
    layer1_outputs(8714) <= not b;
    layer1_outputs(8715) <= b;
    layer1_outputs(8716) <= a and not b;
    layer1_outputs(8717) <= not b or a;
    layer1_outputs(8718) <= 1'b0;
    layer1_outputs(8719) <= a xor b;
    layer1_outputs(8720) <= 1'b1;
    layer1_outputs(8721) <= not a;
    layer1_outputs(8722) <= not a;
    layer1_outputs(8723) <= not (a xor b);
    layer1_outputs(8724) <= a or b;
    layer1_outputs(8725) <= not b;
    layer1_outputs(8726) <= a xor b;
    layer1_outputs(8727) <= a;
    layer1_outputs(8728) <= a;
    layer1_outputs(8729) <= not (a or b);
    layer1_outputs(8730) <= b;
    layer1_outputs(8731) <= a xor b;
    layer1_outputs(8732) <= a and not b;
    layer1_outputs(8733) <= not (a and b);
    layer1_outputs(8734) <= not a;
    layer1_outputs(8735) <= not a;
    layer1_outputs(8736) <= a or b;
    layer1_outputs(8737) <= b;
    layer1_outputs(8738) <= b;
    layer1_outputs(8739) <= not a or b;
    layer1_outputs(8740) <= b and not a;
    layer1_outputs(8741) <= not a or b;
    layer1_outputs(8742) <= a;
    layer1_outputs(8743) <= not a or b;
    layer1_outputs(8744) <= not (a and b);
    layer1_outputs(8745) <= a and not b;
    layer1_outputs(8746) <= not (a or b);
    layer1_outputs(8747) <= not (a xor b);
    layer1_outputs(8748) <= a and not b;
    layer1_outputs(8749) <= not b or a;
    layer1_outputs(8750) <= a or b;
    layer1_outputs(8751) <= a and b;
    layer1_outputs(8752) <= a and b;
    layer1_outputs(8753) <= not (a or b);
    layer1_outputs(8754) <= not b;
    layer1_outputs(8755) <= not (a or b);
    layer1_outputs(8756) <= 1'b1;
    layer1_outputs(8757) <= a and b;
    layer1_outputs(8758) <= a and not b;
    layer1_outputs(8759) <= not b or a;
    layer1_outputs(8760) <= not a or b;
    layer1_outputs(8761) <= b;
    layer1_outputs(8762) <= a or b;
    layer1_outputs(8763) <= not (a and b);
    layer1_outputs(8764) <= not a;
    layer1_outputs(8765) <= 1'b1;
    layer1_outputs(8766) <= not b;
    layer1_outputs(8767) <= 1'b1;
    layer1_outputs(8768) <= not a or b;
    layer1_outputs(8769) <= a and not b;
    layer1_outputs(8770) <= not b or a;
    layer1_outputs(8771) <= a or b;
    layer1_outputs(8772) <= a xor b;
    layer1_outputs(8773) <= b;
    layer1_outputs(8774) <= not b;
    layer1_outputs(8775) <= not a;
    layer1_outputs(8776) <= not (a or b);
    layer1_outputs(8777) <= not b;
    layer1_outputs(8778) <= not a;
    layer1_outputs(8779) <= not (a xor b);
    layer1_outputs(8780) <= a and b;
    layer1_outputs(8781) <= 1'b0;
    layer1_outputs(8782) <= not b or a;
    layer1_outputs(8783) <= not (a and b);
    layer1_outputs(8784) <= not a;
    layer1_outputs(8785) <= not (a or b);
    layer1_outputs(8786) <= not a or b;
    layer1_outputs(8787) <= 1'b1;
    layer1_outputs(8788) <= a and b;
    layer1_outputs(8789) <= a and not b;
    layer1_outputs(8790) <= not b;
    layer1_outputs(8791) <= not (a and b);
    layer1_outputs(8792) <= not (a and b);
    layer1_outputs(8793) <= 1'b0;
    layer1_outputs(8794) <= b;
    layer1_outputs(8795) <= not (a or b);
    layer1_outputs(8796) <= not (a xor b);
    layer1_outputs(8797) <= a and b;
    layer1_outputs(8798) <= not a;
    layer1_outputs(8799) <= not a or b;
    layer1_outputs(8800) <= 1'b0;
    layer1_outputs(8801) <= not a;
    layer1_outputs(8802) <= b;
    layer1_outputs(8803) <= b;
    layer1_outputs(8804) <= b and not a;
    layer1_outputs(8805) <= not (a or b);
    layer1_outputs(8806) <= not a or b;
    layer1_outputs(8807) <= b and not a;
    layer1_outputs(8808) <= not a;
    layer1_outputs(8809) <= not a;
    layer1_outputs(8810) <= a and not b;
    layer1_outputs(8811) <= not a;
    layer1_outputs(8812) <= a and b;
    layer1_outputs(8813) <= not b;
    layer1_outputs(8814) <= b;
    layer1_outputs(8815) <= not (a or b);
    layer1_outputs(8816) <= 1'b0;
    layer1_outputs(8817) <= a and not b;
    layer1_outputs(8818) <= a;
    layer1_outputs(8819) <= b;
    layer1_outputs(8820) <= not a or b;
    layer1_outputs(8821) <= not a or b;
    layer1_outputs(8822) <= a or b;
    layer1_outputs(8823) <= a and b;
    layer1_outputs(8824) <= a and b;
    layer1_outputs(8825) <= not a;
    layer1_outputs(8826) <= not (a or b);
    layer1_outputs(8827) <= not (a xor b);
    layer1_outputs(8828) <= b;
    layer1_outputs(8829) <= not (a and b);
    layer1_outputs(8830) <= not b or a;
    layer1_outputs(8831) <= b and not a;
    layer1_outputs(8832) <= not (a and b);
    layer1_outputs(8833) <= not b;
    layer1_outputs(8834) <= not (a and b);
    layer1_outputs(8835) <= a xor b;
    layer1_outputs(8836) <= not b;
    layer1_outputs(8837) <= b;
    layer1_outputs(8838) <= not (a and b);
    layer1_outputs(8839) <= a or b;
    layer1_outputs(8840) <= a xor b;
    layer1_outputs(8841) <= not b;
    layer1_outputs(8842) <= b and not a;
    layer1_outputs(8843) <= a xor b;
    layer1_outputs(8844) <= not (a xor b);
    layer1_outputs(8845) <= a;
    layer1_outputs(8846) <= not (a xor b);
    layer1_outputs(8847) <= b and not a;
    layer1_outputs(8848) <= not a;
    layer1_outputs(8849) <= not b or a;
    layer1_outputs(8850) <= not b or a;
    layer1_outputs(8851) <= b and not a;
    layer1_outputs(8852) <= 1'b0;
    layer1_outputs(8853) <= a;
    layer1_outputs(8854) <= b;
    layer1_outputs(8855) <= not b;
    layer1_outputs(8856) <= not b;
    layer1_outputs(8857) <= not (a or b);
    layer1_outputs(8858) <= a;
    layer1_outputs(8859) <= a and not b;
    layer1_outputs(8860) <= 1'b0;
    layer1_outputs(8861) <= a and b;
    layer1_outputs(8862) <= 1'b1;
    layer1_outputs(8863) <= a or b;
    layer1_outputs(8864) <= not (a xor b);
    layer1_outputs(8865) <= not a;
    layer1_outputs(8866) <= a or b;
    layer1_outputs(8867) <= not (a or b);
    layer1_outputs(8868) <= not b or a;
    layer1_outputs(8869) <= a or b;
    layer1_outputs(8870) <= not (a xor b);
    layer1_outputs(8871) <= a or b;
    layer1_outputs(8872) <= a;
    layer1_outputs(8873) <= b;
    layer1_outputs(8874) <= not b or a;
    layer1_outputs(8875) <= a;
    layer1_outputs(8876) <= not a;
    layer1_outputs(8877) <= a xor b;
    layer1_outputs(8878) <= b;
    layer1_outputs(8879) <= a;
    layer1_outputs(8880) <= not b;
    layer1_outputs(8881) <= not (a or b);
    layer1_outputs(8882) <= a;
    layer1_outputs(8883) <= not (a xor b);
    layer1_outputs(8884) <= not b;
    layer1_outputs(8885) <= not a;
    layer1_outputs(8886) <= not (a and b);
    layer1_outputs(8887) <= not b;
    layer1_outputs(8888) <= b;
    layer1_outputs(8889) <= b;
    layer1_outputs(8890) <= a or b;
    layer1_outputs(8891) <= not b or a;
    layer1_outputs(8892) <= 1'b1;
    layer1_outputs(8893) <= not (a or b);
    layer1_outputs(8894) <= 1'b1;
    layer1_outputs(8895) <= not a;
    layer1_outputs(8896) <= not b or a;
    layer1_outputs(8897) <= a;
    layer1_outputs(8898) <= a or b;
    layer1_outputs(8899) <= a;
    layer1_outputs(8900) <= not b;
    layer1_outputs(8901) <= not b;
    layer1_outputs(8902) <= a and b;
    layer1_outputs(8903) <= a;
    layer1_outputs(8904) <= not a;
    layer1_outputs(8905) <= not (a xor b);
    layer1_outputs(8906) <= not b;
    layer1_outputs(8907) <= not b or a;
    layer1_outputs(8908) <= not a;
    layer1_outputs(8909) <= a xor b;
    layer1_outputs(8910) <= a and not b;
    layer1_outputs(8911) <= a or b;
    layer1_outputs(8912) <= a xor b;
    layer1_outputs(8913) <= not (a or b);
    layer1_outputs(8914) <= b and not a;
    layer1_outputs(8915) <= not a;
    layer1_outputs(8916) <= a xor b;
    layer1_outputs(8917) <= not b or a;
    layer1_outputs(8918) <= b;
    layer1_outputs(8919) <= b;
    layer1_outputs(8920) <= not (a xor b);
    layer1_outputs(8921) <= not b or a;
    layer1_outputs(8922) <= not a;
    layer1_outputs(8923) <= a or b;
    layer1_outputs(8924) <= a;
    layer1_outputs(8925) <= b;
    layer1_outputs(8926) <= not b;
    layer1_outputs(8927) <= a and b;
    layer1_outputs(8928) <= not (a or b);
    layer1_outputs(8929) <= 1'b1;
    layer1_outputs(8930) <= not a or b;
    layer1_outputs(8931) <= a and not b;
    layer1_outputs(8932) <= a and not b;
    layer1_outputs(8933) <= b;
    layer1_outputs(8934) <= not a;
    layer1_outputs(8935) <= not b;
    layer1_outputs(8936) <= not (a xor b);
    layer1_outputs(8937) <= a;
    layer1_outputs(8938) <= not b or a;
    layer1_outputs(8939) <= 1'b1;
    layer1_outputs(8940) <= b and not a;
    layer1_outputs(8941) <= 1'b0;
    layer1_outputs(8942) <= not b;
    layer1_outputs(8943) <= a;
    layer1_outputs(8944) <= b;
    layer1_outputs(8945) <= not (a or b);
    layer1_outputs(8946) <= a and not b;
    layer1_outputs(8947) <= not a;
    layer1_outputs(8948) <= 1'b1;
    layer1_outputs(8949) <= not a;
    layer1_outputs(8950) <= b and not a;
    layer1_outputs(8951) <= a or b;
    layer1_outputs(8952) <= b;
    layer1_outputs(8953) <= b;
    layer1_outputs(8954) <= not a;
    layer1_outputs(8955) <= not a;
    layer1_outputs(8956) <= a xor b;
    layer1_outputs(8957) <= a or b;
    layer1_outputs(8958) <= not a or b;
    layer1_outputs(8959) <= not (a and b);
    layer1_outputs(8960) <= b;
    layer1_outputs(8961) <= not (a or b);
    layer1_outputs(8962) <= a;
    layer1_outputs(8963) <= not b or a;
    layer1_outputs(8964) <= 1'b0;
    layer1_outputs(8965) <= a or b;
    layer1_outputs(8966) <= b and not a;
    layer1_outputs(8967) <= a and b;
    layer1_outputs(8968) <= 1'b1;
    layer1_outputs(8969) <= not (a xor b);
    layer1_outputs(8970) <= a xor b;
    layer1_outputs(8971) <= a and b;
    layer1_outputs(8972) <= a;
    layer1_outputs(8973) <= b;
    layer1_outputs(8974) <= b;
    layer1_outputs(8975) <= 1'b1;
    layer1_outputs(8976) <= b and not a;
    layer1_outputs(8977) <= not b or a;
    layer1_outputs(8978) <= a xor b;
    layer1_outputs(8979) <= a xor b;
    layer1_outputs(8980) <= a xor b;
    layer1_outputs(8981) <= a or b;
    layer1_outputs(8982) <= not (a xor b);
    layer1_outputs(8983) <= b;
    layer1_outputs(8984) <= a xor b;
    layer1_outputs(8985) <= 1'b1;
    layer1_outputs(8986) <= a;
    layer1_outputs(8987) <= b and not a;
    layer1_outputs(8988) <= a xor b;
    layer1_outputs(8989) <= not a;
    layer1_outputs(8990) <= b;
    layer1_outputs(8991) <= b;
    layer1_outputs(8992) <= a and b;
    layer1_outputs(8993) <= a and b;
    layer1_outputs(8994) <= a or b;
    layer1_outputs(8995) <= a or b;
    layer1_outputs(8996) <= a xor b;
    layer1_outputs(8997) <= not a or b;
    layer1_outputs(8998) <= not (a xor b);
    layer1_outputs(8999) <= not a;
    layer1_outputs(9000) <= a and not b;
    layer1_outputs(9001) <= b and not a;
    layer1_outputs(9002) <= 1'b0;
    layer1_outputs(9003) <= a;
    layer1_outputs(9004) <= b and not a;
    layer1_outputs(9005) <= a or b;
    layer1_outputs(9006) <= not (a xor b);
    layer1_outputs(9007) <= not (a xor b);
    layer1_outputs(9008) <= not b or a;
    layer1_outputs(9009) <= b;
    layer1_outputs(9010) <= b;
    layer1_outputs(9011) <= a or b;
    layer1_outputs(9012) <= not (a and b);
    layer1_outputs(9013) <= a or b;
    layer1_outputs(9014) <= a xor b;
    layer1_outputs(9015) <= a and b;
    layer1_outputs(9016) <= not b;
    layer1_outputs(9017) <= not b;
    layer1_outputs(9018) <= not a;
    layer1_outputs(9019) <= b and not a;
    layer1_outputs(9020) <= not a or b;
    layer1_outputs(9021) <= not a;
    layer1_outputs(9022) <= not a;
    layer1_outputs(9023) <= not a;
    layer1_outputs(9024) <= not b;
    layer1_outputs(9025) <= b;
    layer1_outputs(9026) <= not a or b;
    layer1_outputs(9027) <= a and b;
    layer1_outputs(9028) <= not (a xor b);
    layer1_outputs(9029) <= a;
    layer1_outputs(9030) <= a or b;
    layer1_outputs(9031) <= a;
    layer1_outputs(9032) <= not b;
    layer1_outputs(9033) <= not (a and b);
    layer1_outputs(9034) <= not b;
    layer1_outputs(9035) <= a or b;
    layer1_outputs(9036) <= not b;
    layer1_outputs(9037) <= not b or a;
    layer1_outputs(9038) <= not a;
    layer1_outputs(9039) <= not a;
    layer1_outputs(9040) <= not b;
    layer1_outputs(9041) <= not a or b;
    layer1_outputs(9042) <= a;
    layer1_outputs(9043) <= a or b;
    layer1_outputs(9044) <= a and b;
    layer1_outputs(9045) <= not b or a;
    layer1_outputs(9046) <= not (a or b);
    layer1_outputs(9047) <= not a;
    layer1_outputs(9048) <= a and not b;
    layer1_outputs(9049) <= 1'b0;
    layer1_outputs(9050) <= a or b;
    layer1_outputs(9051) <= not a;
    layer1_outputs(9052) <= b;
    layer1_outputs(9053) <= not b or a;
    layer1_outputs(9054) <= a xor b;
    layer1_outputs(9055) <= b;
    layer1_outputs(9056) <= a and b;
    layer1_outputs(9057) <= not b;
    layer1_outputs(9058) <= not a;
    layer1_outputs(9059) <= 1'b0;
    layer1_outputs(9060) <= not (a xor b);
    layer1_outputs(9061) <= b and not a;
    layer1_outputs(9062) <= b and not a;
    layer1_outputs(9063) <= not (a or b);
    layer1_outputs(9064) <= not b;
    layer1_outputs(9065) <= not (a and b);
    layer1_outputs(9066) <= b and not a;
    layer1_outputs(9067) <= a and b;
    layer1_outputs(9068) <= a or b;
    layer1_outputs(9069) <= a and not b;
    layer1_outputs(9070) <= not (a or b);
    layer1_outputs(9071) <= not a;
    layer1_outputs(9072) <= not b or a;
    layer1_outputs(9073) <= 1'b1;
    layer1_outputs(9074) <= b;
    layer1_outputs(9075) <= not (a or b);
    layer1_outputs(9076) <= a and not b;
    layer1_outputs(9077) <= not b;
    layer1_outputs(9078) <= not b or a;
    layer1_outputs(9079) <= not b;
    layer1_outputs(9080) <= not (a and b);
    layer1_outputs(9081) <= a or b;
    layer1_outputs(9082) <= a;
    layer1_outputs(9083) <= a and b;
    layer1_outputs(9084) <= not (a and b);
    layer1_outputs(9085) <= a and not b;
    layer1_outputs(9086) <= not (a or b);
    layer1_outputs(9087) <= not b;
    layer1_outputs(9088) <= a or b;
    layer1_outputs(9089) <= not a;
    layer1_outputs(9090) <= a xor b;
    layer1_outputs(9091) <= 1'b0;
    layer1_outputs(9092) <= a or b;
    layer1_outputs(9093) <= not (a and b);
    layer1_outputs(9094) <= a and b;
    layer1_outputs(9095) <= a;
    layer1_outputs(9096) <= b;
    layer1_outputs(9097) <= not (a or b);
    layer1_outputs(9098) <= b and not a;
    layer1_outputs(9099) <= a xor b;
    layer1_outputs(9100) <= b and not a;
    layer1_outputs(9101) <= 1'b1;
    layer1_outputs(9102) <= not b;
    layer1_outputs(9103) <= a;
    layer1_outputs(9104) <= a xor b;
    layer1_outputs(9105) <= not a or b;
    layer1_outputs(9106) <= not b or a;
    layer1_outputs(9107) <= not (a xor b);
    layer1_outputs(9108) <= not (a or b);
    layer1_outputs(9109) <= a;
    layer1_outputs(9110) <= not a;
    layer1_outputs(9111) <= a;
    layer1_outputs(9112) <= a and not b;
    layer1_outputs(9113) <= not a;
    layer1_outputs(9114) <= a and b;
    layer1_outputs(9115) <= not a or b;
    layer1_outputs(9116) <= a;
    layer1_outputs(9117) <= b and not a;
    layer1_outputs(9118) <= a or b;
    layer1_outputs(9119) <= b and not a;
    layer1_outputs(9120) <= a and b;
    layer1_outputs(9121) <= not a;
    layer1_outputs(9122) <= not a or b;
    layer1_outputs(9123) <= a or b;
    layer1_outputs(9124) <= a xor b;
    layer1_outputs(9125) <= not a;
    layer1_outputs(9126) <= not (a xor b);
    layer1_outputs(9127) <= not b or a;
    layer1_outputs(9128) <= not a;
    layer1_outputs(9129) <= not b;
    layer1_outputs(9130) <= not (a xor b);
    layer1_outputs(9131) <= b;
    layer1_outputs(9132) <= not b or a;
    layer1_outputs(9133) <= a xor b;
    layer1_outputs(9134) <= b;
    layer1_outputs(9135) <= not a or b;
    layer1_outputs(9136) <= a and b;
    layer1_outputs(9137) <= a xor b;
    layer1_outputs(9138) <= not (a and b);
    layer1_outputs(9139) <= not (a and b);
    layer1_outputs(9140) <= a and b;
    layer1_outputs(9141) <= not a;
    layer1_outputs(9142) <= a and b;
    layer1_outputs(9143) <= not a;
    layer1_outputs(9144) <= not a or b;
    layer1_outputs(9145) <= b;
    layer1_outputs(9146) <= 1'b0;
    layer1_outputs(9147) <= a and b;
    layer1_outputs(9148) <= a;
    layer1_outputs(9149) <= 1'b1;
    layer1_outputs(9150) <= b;
    layer1_outputs(9151) <= a or b;
    layer1_outputs(9152) <= b;
    layer1_outputs(9153) <= 1'b0;
    layer1_outputs(9154) <= a and b;
    layer1_outputs(9155) <= b;
    layer1_outputs(9156) <= a and not b;
    layer1_outputs(9157) <= 1'b1;
    layer1_outputs(9158) <= not (a or b);
    layer1_outputs(9159) <= a and not b;
    layer1_outputs(9160) <= not b;
    layer1_outputs(9161) <= not b;
    layer1_outputs(9162) <= not (a or b);
    layer1_outputs(9163) <= a and b;
    layer1_outputs(9164) <= not a;
    layer1_outputs(9165) <= not a or b;
    layer1_outputs(9166) <= b;
    layer1_outputs(9167) <= a and b;
    layer1_outputs(9168) <= not (a and b);
    layer1_outputs(9169) <= not a;
    layer1_outputs(9170) <= a xor b;
    layer1_outputs(9171) <= not b;
    layer1_outputs(9172) <= not (a or b);
    layer1_outputs(9173) <= 1'b1;
    layer1_outputs(9174) <= a xor b;
    layer1_outputs(9175) <= 1'b1;
    layer1_outputs(9176) <= a;
    layer1_outputs(9177) <= b;
    layer1_outputs(9178) <= not b;
    layer1_outputs(9179) <= not b;
    layer1_outputs(9180) <= not (a and b);
    layer1_outputs(9181) <= a xor b;
    layer1_outputs(9182) <= 1'b1;
    layer1_outputs(9183) <= not b or a;
    layer1_outputs(9184) <= b;
    layer1_outputs(9185) <= a and b;
    layer1_outputs(9186) <= not a or b;
    layer1_outputs(9187) <= a and not b;
    layer1_outputs(9188) <= not (a xor b);
    layer1_outputs(9189) <= not a;
    layer1_outputs(9190) <= not (a and b);
    layer1_outputs(9191) <= a or b;
    layer1_outputs(9192) <= a and b;
    layer1_outputs(9193) <= 1'b1;
    layer1_outputs(9194) <= a or b;
    layer1_outputs(9195) <= b;
    layer1_outputs(9196) <= a and not b;
    layer1_outputs(9197) <= a and b;
    layer1_outputs(9198) <= not a;
    layer1_outputs(9199) <= not b or a;
    layer1_outputs(9200) <= b;
    layer1_outputs(9201) <= a or b;
    layer1_outputs(9202) <= not (a xor b);
    layer1_outputs(9203) <= not a;
    layer1_outputs(9204) <= not a or b;
    layer1_outputs(9205) <= b;
    layer1_outputs(9206) <= not a;
    layer1_outputs(9207) <= a and not b;
    layer1_outputs(9208) <= a;
    layer1_outputs(9209) <= a xor b;
    layer1_outputs(9210) <= not b;
    layer1_outputs(9211) <= b and not a;
    layer1_outputs(9212) <= not b;
    layer1_outputs(9213) <= not a;
    layer1_outputs(9214) <= not b;
    layer1_outputs(9215) <= not b;
    layer1_outputs(9216) <= b and not a;
    layer1_outputs(9217) <= not a;
    layer1_outputs(9218) <= not b or a;
    layer1_outputs(9219) <= a xor b;
    layer1_outputs(9220) <= not b or a;
    layer1_outputs(9221) <= not (a and b);
    layer1_outputs(9222) <= b;
    layer1_outputs(9223) <= not b;
    layer1_outputs(9224) <= not (a or b);
    layer1_outputs(9225) <= a and not b;
    layer1_outputs(9226) <= not (a and b);
    layer1_outputs(9227) <= not b;
    layer1_outputs(9228) <= b;
    layer1_outputs(9229) <= a and not b;
    layer1_outputs(9230) <= a;
    layer1_outputs(9231) <= b;
    layer1_outputs(9232) <= a and not b;
    layer1_outputs(9233) <= not (a or b);
    layer1_outputs(9234) <= a;
    layer1_outputs(9235) <= not a or b;
    layer1_outputs(9236) <= b and not a;
    layer1_outputs(9237) <= a xor b;
    layer1_outputs(9238) <= not b or a;
    layer1_outputs(9239) <= a and not b;
    layer1_outputs(9240) <= b and not a;
    layer1_outputs(9241) <= not a or b;
    layer1_outputs(9242) <= a xor b;
    layer1_outputs(9243) <= a;
    layer1_outputs(9244) <= not (a or b);
    layer1_outputs(9245) <= not a;
    layer1_outputs(9246) <= not a or b;
    layer1_outputs(9247) <= not a or b;
    layer1_outputs(9248) <= 1'b1;
    layer1_outputs(9249) <= a and b;
    layer1_outputs(9250) <= a and not b;
    layer1_outputs(9251) <= not b;
    layer1_outputs(9252) <= a and b;
    layer1_outputs(9253) <= not (a or b);
    layer1_outputs(9254) <= not b or a;
    layer1_outputs(9255) <= b;
    layer1_outputs(9256) <= a and b;
    layer1_outputs(9257) <= not (a and b);
    layer1_outputs(9258) <= not a;
    layer1_outputs(9259) <= a;
    layer1_outputs(9260) <= not a or b;
    layer1_outputs(9261) <= not a;
    layer1_outputs(9262) <= not b;
    layer1_outputs(9263) <= a;
    layer1_outputs(9264) <= a or b;
    layer1_outputs(9265) <= not a or b;
    layer1_outputs(9266) <= not a;
    layer1_outputs(9267) <= not (a xor b);
    layer1_outputs(9268) <= not (a xor b);
    layer1_outputs(9269) <= not a;
    layer1_outputs(9270) <= a or b;
    layer1_outputs(9271) <= not (a or b);
    layer1_outputs(9272) <= a xor b;
    layer1_outputs(9273) <= 1'b1;
    layer1_outputs(9274) <= not b;
    layer1_outputs(9275) <= b and not a;
    layer1_outputs(9276) <= not (a xor b);
    layer1_outputs(9277) <= not a or b;
    layer1_outputs(9278) <= a;
    layer1_outputs(9279) <= a and b;
    layer1_outputs(9280) <= not a or b;
    layer1_outputs(9281) <= not (a or b);
    layer1_outputs(9282) <= not (a and b);
    layer1_outputs(9283) <= a or b;
    layer1_outputs(9284) <= not (a xor b);
    layer1_outputs(9285) <= not (a or b);
    layer1_outputs(9286) <= not (a or b);
    layer1_outputs(9287) <= a and not b;
    layer1_outputs(9288) <= b;
    layer1_outputs(9289) <= b and not a;
    layer1_outputs(9290) <= a;
    layer1_outputs(9291) <= a and not b;
    layer1_outputs(9292) <= a;
    layer1_outputs(9293) <= a or b;
    layer1_outputs(9294) <= not (a or b);
    layer1_outputs(9295) <= not b;
    layer1_outputs(9296) <= a or b;
    layer1_outputs(9297) <= 1'b0;
    layer1_outputs(9298) <= a and not b;
    layer1_outputs(9299) <= not b;
    layer1_outputs(9300) <= a or b;
    layer1_outputs(9301) <= a or b;
    layer1_outputs(9302) <= a and not b;
    layer1_outputs(9303) <= not a or b;
    layer1_outputs(9304) <= a or b;
    layer1_outputs(9305) <= not b;
    layer1_outputs(9306) <= a and b;
    layer1_outputs(9307) <= a and b;
    layer1_outputs(9308) <= 1'b1;
    layer1_outputs(9309) <= not (a or b);
    layer1_outputs(9310) <= a and b;
    layer1_outputs(9311) <= not a;
    layer1_outputs(9312) <= a;
    layer1_outputs(9313) <= 1'b1;
    layer1_outputs(9314) <= a;
    layer1_outputs(9315) <= not (a or b);
    layer1_outputs(9316) <= b;
    layer1_outputs(9317) <= not (a and b);
    layer1_outputs(9318) <= a;
    layer1_outputs(9319) <= 1'b1;
    layer1_outputs(9320) <= a;
    layer1_outputs(9321) <= 1'b0;
    layer1_outputs(9322) <= a;
    layer1_outputs(9323) <= a and b;
    layer1_outputs(9324) <= b and not a;
    layer1_outputs(9325) <= a and b;
    layer1_outputs(9326) <= not (a xor b);
    layer1_outputs(9327) <= not (a or b);
    layer1_outputs(9328) <= b;
    layer1_outputs(9329) <= a and not b;
    layer1_outputs(9330) <= a and b;
    layer1_outputs(9331) <= not b or a;
    layer1_outputs(9332) <= not (a xor b);
    layer1_outputs(9333) <= not (a or b);
    layer1_outputs(9334) <= not (a and b);
    layer1_outputs(9335) <= b and not a;
    layer1_outputs(9336) <= not a;
    layer1_outputs(9337) <= not b;
    layer1_outputs(9338) <= a or b;
    layer1_outputs(9339) <= 1'b1;
    layer1_outputs(9340) <= a;
    layer1_outputs(9341) <= a xor b;
    layer1_outputs(9342) <= a and not b;
    layer1_outputs(9343) <= a;
    layer1_outputs(9344) <= not a;
    layer1_outputs(9345) <= a or b;
    layer1_outputs(9346) <= a or b;
    layer1_outputs(9347) <= a xor b;
    layer1_outputs(9348) <= b;
    layer1_outputs(9349) <= b;
    layer1_outputs(9350) <= not (a and b);
    layer1_outputs(9351) <= not (a or b);
    layer1_outputs(9352) <= not b or a;
    layer1_outputs(9353) <= 1'b1;
    layer1_outputs(9354) <= not (a and b);
    layer1_outputs(9355) <= not (a and b);
    layer1_outputs(9356) <= a and not b;
    layer1_outputs(9357) <= a;
    layer1_outputs(9358) <= a and b;
    layer1_outputs(9359) <= not a;
    layer1_outputs(9360) <= b and not a;
    layer1_outputs(9361) <= a;
    layer1_outputs(9362) <= a and not b;
    layer1_outputs(9363) <= not (a xor b);
    layer1_outputs(9364) <= a or b;
    layer1_outputs(9365) <= a or b;
    layer1_outputs(9366) <= not b or a;
    layer1_outputs(9367) <= a;
    layer1_outputs(9368) <= not (a and b);
    layer1_outputs(9369) <= a or b;
    layer1_outputs(9370) <= not (a and b);
    layer1_outputs(9371) <= not b or a;
    layer1_outputs(9372) <= b;
    layer1_outputs(9373) <= b and not a;
    layer1_outputs(9374) <= not a or b;
    layer1_outputs(9375) <= a xor b;
    layer1_outputs(9376) <= 1'b0;
    layer1_outputs(9377) <= a;
    layer1_outputs(9378) <= not b or a;
    layer1_outputs(9379) <= not b;
    layer1_outputs(9380) <= not b or a;
    layer1_outputs(9381) <= a and b;
    layer1_outputs(9382) <= 1'b1;
    layer1_outputs(9383) <= not a;
    layer1_outputs(9384) <= not b or a;
    layer1_outputs(9385) <= a and b;
    layer1_outputs(9386) <= a;
    layer1_outputs(9387) <= a and not b;
    layer1_outputs(9388) <= not b;
    layer1_outputs(9389) <= 1'b0;
    layer1_outputs(9390) <= not b;
    layer1_outputs(9391) <= not a;
    layer1_outputs(9392) <= a;
    layer1_outputs(9393) <= not (a and b);
    layer1_outputs(9394) <= b and not a;
    layer1_outputs(9395) <= not b;
    layer1_outputs(9396) <= not a;
    layer1_outputs(9397) <= not a or b;
    layer1_outputs(9398) <= a or b;
    layer1_outputs(9399) <= not a or b;
    layer1_outputs(9400) <= 1'b0;
    layer1_outputs(9401) <= not (a xor b);
    layer1_outputs(9402) <= not b or a;
    layer1_outputs(9403) <= a;
    layer1_outputs(9404) <= a and not b;
    layer1_outputs(9405) <= b;
    layer1_outputs(9406) <= not (a and b);
    layer1_outputs(9407) <= not b;
    layer1_outputs(9408) <= b;
    layer1_outputs(9409) <= not (a or b);
    layer1_outputs(9410) <= not a or b;
    layer1_outputs(9411) <= not b or a;
    layer1_outputs(9412) <= not (a or b);
    layer1_outputs(9413) <= not b or a;
    layer1_outputs(9414) <= not (a xor b);
    layer1_outputs(9415) <= not b;
    layer1_outputs(9416) <= not (a or b);
    layer1_outputs(9417) <= a and not b;
    layer1_outputs(9418) <= not (a and b);
    layer1_outputs(9419) <= a;
    layer1_outputs(9420) <= a and b;
    layer1_outputs(9421) <= not a or b;
    layer1_outputs(9422) <= not a;
    layer1_outputs(9423) <= not b or a;
    layer1_outputs(9424) <= a xor b;
    layer1_outputs(9425) <= a and b;
    layer1_outputs(9426) <= a;
    layer1_outputs(9427) <= a and not b;
    layer1_outputs(9428) <= 1'b0;
    layer1_outputs(9429) <= not (a and b);
    layer1_outputs(9430) <= not (a or b);
    layer1_outputs(9431) <= b;
    layer1_outputs(9432) <= not b;
    layer1_outputs(9433) <= 1'b0;
    layer1_outputs(9434) <= b;
    layer1_outputs(9435) <= a;
    layer1_outputs(9436) <= a;
    layer1_outputs(9437) <= b;
    layer1_outputs(9438) <= a and b;
    layer1_outputs(9439) <= not (a xor b);
    layer1_outputs(9440) <= not (a and b);
    layer1_outputs(9441) <= not a;
    layer1_outputs(9442) <= not (a and b);
    layer1_outputs(9443) <= not b;
    layer1_outputs(9444) <= not (a or b);
    layer1_outputs(9445) <= not (a xor b);
    layer1_outputs(9446) <= not (a and b);
    layer1_outputs(9447) <= not a;
    layer1_outputs(9448) <= 1'b1;
    layer1_outputs(9449) <= b and not a;
    layer1_outputs(9450) <= not (a xor b);
    layer1_outputs(9451) <= not (a or b);
    layer1_outputs(9452) <= not a or b;
    layer1_outputs(9453) <= not b or a;
    layer1_outputs(9454) <= a and b;
    layer1_outputs(9455) <= not (a or b);
    layer1_outputs(9456) <= not b;
    layer1_outputs(9457) <= a xor b;
    layer1_outputs(9458) <= not (a or b);
    layer1_outputs(9459) <= not b;
    layer1_outputs(9460) <= 1'b1;
    layer1_outputs(9461) <= not b or a;
    layer1_outputs(9462) <= a and b;
    layer1_outputs(9463) <= not a;
    layer1_outputs(9464) <= a and b;
    layer1_outputs(9465) <= a or b;
    layer1_outputs(9466) <= not a;
    layer1_outputs(9467) <= a and not b;
    layer1_outputs(9468) <= not a;
    layer1_outputs(9469) <= a and not b;
    layer1_outputs(9470) <= not b or a;
    layer1_outputs(9471) <= a and b;
    layer1_outputs(9472) <= not (a or b);
    layer1_outputs(9473) <= a and b;
    layer1_outputs(9474) <= b;
    layer1_outputs(9475) <= not (a xor b);
    layer1_outputs(9476) <= a;
    layer1_outputs(9477) <= b;
    layer1_outputs(9478) <= not (a and b);
    layer1_outputs(9479) <= a and not b;
    layer1_outputs(9480) <= b;
    layer1_outputs(9481) <= not a or b;
    layer1_outputs(9482) <= a;
    layer1_outputs(9483) <= 1'b1;
    layer1_outputs(9484) <= not (a or b);
    layer1_outputs(9485) <= not (a and b);
    layer1_outputs(9486) <= not b;
    layer1_outputs(9487) <= not (a and b);
    layer1_outputs(9488) <= not a;
    layer1_outputs(9489) <= b;
    layer1_outputs(9490) <= not b;
    layer1_outputs(9491) <= a;
    layer1_outputs(9492) <= a and not b;
    layer1_outputs(9493) <= not (a and b);
    layer1_outputs(9494) <= not a or b;
    layer1_outputs(9495) <= a and not b;
    layer1_outputs(9496) <= not (a or b);
    layer1_outputs(9497) <= not (a or b);
    layer1_outputs(9498) <= a and b;
    layer1_outputs(9499) <= not b or a;
    layer1_outputs(9500) <= not a or b;
    layer1_outputs(9501) <= not (a or b);
    layer1_outputs(9502) <= not (a and b);
    layer1_outputs(9503) <= a or b;
    layer1_outputs(9504) <= a and not b;
    layer1_outputs(9505) <= not (a and b);
    layer1_outputs(9506) <= not b;
    layer1_outputs(9507) <= a;
    layer1_outputs(9508) <= not a;
    layer1_outputs(9509) <= not (a or b);
    layer1_outputs(9510) <= b;
    layer1_outputs(9511) <= a or b;
    layer1_outputs(9512) <= not (a or b);
    layer1_outputs(9513) <= not (a or b);
    layer1_outputs(9514) <= a xor b;
    layer1_outputs(9515) <= a;
    layer1_outputs(9516) <= 1'b1;
    layer1_outputs(9517) <= a and not b;
    layer1_outputs(9518) <= not (a and b);
    layer1_outputs(9519) <= a and b;
    layer1_outputs(9520) <= not (a or b);
    layer1_outputs(9521) <= 1'b1;
    layer1_outputs(9522) <= not a;
    layer1_outputs(9523) <= a xor b;
    layer1_outputs(9524) <= a and not b;
    layer1_outputs(9525) <= a and b;
    layer1_outputs(9526) <= not b or a;
    layer1_outputs(9527) <= not b or a;
    layer1_outputs(9528) <= not a;
    layer1_outputs(9529) <= b;
    layer1_outputs(9530) <= not (a xor b);
    layer1_outputs(9531) <= a and not b;
    layer1_outputs(9532) <= a xor b;
    layer1_outputs(9533) <= not (a xor b);
    layer1_outputs(9534) <= b and not a;
    layer1_outputs(9535) <= b;
    layer1_outputs(9536) <= not a or b;
    layer1_outputs(9537) <= a;
    layer1_outputs(9538) <= a and not b;
    layer1_outputs(9539) <= a and not b;
    layer1_outputs(9540) <= not (a xor b);
    layer1_outputs(9541) <= a;
    layer1_outputs(9542) <= a;
    layer1_outputs(9543) <= b;
    layer1_outputs(9544) <= not a or b;
    layer1_outputs(9545) <= b;
    layer1_outputs(9546) <= b and not a;
    layer1_outputs(9547) <= 1'b0;
    layer1_outputs(9548) <= b and not a;
    layer1_outputs(9549) <= not a;
    layer1_outputs(9550) <= a xor b;
    layer1_outputs(9551) <= a;
    layer1_outputs(9552) <= a or b;
    layer1_outputs(9553) <= a or b;
    layer1_outputs(9554) <= b;
    layer1_outputs(9555) <= a;
    layer1_outputs(9556) <= not a;
    layer1_outputs(9557) <= a;
    layer1_outputs(9558) <= not b;
    layer1_outputs(9559) <= a and not b;
    layer1_outputs(9560) <= not a;
    layer1_outputs(9561) <= not (a xor b);
    layer1_outputs(9562) <= b;
    layer1_outputs(9563) <= not (a xor b);
    layer1_outputs(9564) <= b and not a;
    layer1_outputs(9565) <= not b;
    layer1_outputs(9566) <= not a;
    layer1_outputs(9567) <= a or b;
    layer1_outputs(9568) <= b and not a;
    layer1_outputs(9569) <= a;
    layer1_outputs(9570) <= a;
    layer1_outputs(9571) <= a and b;
    layer1_outputs(9572) <= a xor b;
    layer1_outputs(9573) <= not a;
    layer1_outputs(9574) <= a;
    layer1_outputs(9575) <= a and b;
    layer1_outputs(9576) <= not (a xor b);
    layer1_outputs(9577) <= b and not a;
    layer1_outputs(9578) <= not a or b;
    layer1_outputs(9579) <= a and b;
    layer1_outputs(9580) <= 1'b0;
    layer1_outputs(9581) <= not (a and b);
    layer1_outputs(9582) <= not b;
    layer1_outputs(9583) <= not a;
    layer1_outputs(9584) <= not b;
    layer1_outputs(9585) <= b and not a;
    layer1_outputs(9586) <= not b;
    layer1_outputs(9587) <= 1'b0;
    layer1_outputs(9588) <= a;
    layer1_outputs(9589) <= not (a or b);
    layer1_outputs(9590) <= b;
    layer1_outputs(9591) <= b and not a;
    layer1_outputs(9592) <= not (a xor b);
    layer1_outputs(9593) <= b and not a;
    layer1_outputs(9594) <= not b;
    layer1_outputs(9595) <= not (a or b);
    layer1_outputs(9596) <= not a;
    layer1_outputs(9597) <= not b;
    layer1_outputs(9598) <= not (a and b);
    layer1_outputs(9599) <= not (a and b);
    layer1_outputs(9600) <= not a or b;
    layer1_outputs(9601) <= b and not a;
    layer1_outputs(9602) <= b;
    layer1_outputs(9603) <= not a;
    layer1_outputs(9604) <= a xor b;
    layer1_outputs(9605) <= b;
    layer1_outputs(9606) <= not b;
    layer1_outputs(9607) <= 1'b0;
    layer1_outputs(9608) <= a or b;
    layer1_outputs(9609) <= not a or b;
    layer1_outputs(9610) <= not a or b;
    layer1_outputs(9611) <= b and not a;
    layer1_outputs(9612) <= not b;
    layer1_outputs(9613) <= b;
    layer1_outputs(9614) <= not (a or b);
    layer1_outputs(9615) <= a and not b;
    layer1_outputs(9616) <= a;
    layer1_outputs(9617) <= not b;
    layer1_outputs(9618) <= a and not b;
    layer1_outputs(9619) <= not a or b;
    layer1_outputs(9620) <= a and not b;
    layer1_outputs(9621) <= not a;
    layer1_outputs(9622) <= not (a xor b);
    layer1_outputs(9623) <= b;
    layer1_outputs(9624) <= not b;
    layer1_outputs(9625) <= not b;
    layer1_outputs(9626) <= b;
    layer1_outputs(9627) <= not (a or b);
    layer1_outputs(9628) <= a xor b;
    layer1_outputs(9629) <= 1'b0;
    layer1_outputs(9630) <= not b;
    layer1_outputs(9631) <= not a or b;
    layer1_outputs(9632) <= not b;
    layer1_outputs(9633) <= a or b;
    layer1_outputs(9634) <= a;
    layer1_outputs(9635) <= not a or b;
    layer1_outputs(9636) <= b;
    layer1_outputs(9637) <= not a;
    layer1_outputs(9638) <= a and not b;
    layer1_outputs(9639) <= a or b;
    layer1_outputs(9640) <= not b or a;
    layer1_outputs(9641) <= not (a and b);
    layer1_outputs(9642) <= not (a or b);
    layer1_outputs(9643) <= b and not a;
    layer1_outputs(9644) <= a;
    layer1_outputs(9645) <= b;
    layer1_outputs(9646) <= not a;
    layer1_outputs(9647) <= a;
    layer1_outputs(9648) <= not b or a;
    layer1_outputs(9649) <= not (a or b);
    layer1_outputs(9650) <= b;
    layer1_outputs(9651) <= not a or b;
    layer1_outputs(9652) <= not b or a;
    layer1_outputs(9653) <= a;
    layer1_outputs(9654) <= a and b;
    layer1_outputs(9655) <= not (a or b);
    layer1_outputs(9656) <= a and not b;
    layer1_outputs(9657) <= a;
    layer1_outputs(9658) <= not b;
    layer1_outputs(9659) <= a xor b;
    layer1_outputs(9660) <= 1'b0;
    layer1_outputs(9661) <= not b or a;
    layer1_outputs(9662) <= b and not a;
    layer1_outputs(9663) <= a and b;
    layer1_outputs(9664) <= a and not b;
    layer1_outputs(9665) <= a;
    layer1_outputs(9666) <= a and not b;
    layer1_outputs(9667) <= a xor b;
    layer1_outputs(9668) <= a or b;
    layer1_outputs(9669) <= not b;
    layer1_outputs(9670) <= not (a and b);
    layer1_outputs(9671) <= a xor b;
    layer1_outputs(9672) <= not a;
    layer1_outputs(9673) <= b;
    layer1_outputs(9674) <= not a;
    layer1_outputs(9675) <= a;
    layer1_outputs(9676) <= 1'b0;
    layer1_outputs(9677) <= a and not b;
    layer1_outputs(9678) <= not a or b;
    layer1_outputs(9679) <= 1'b1;
    layer1_outputs(9680) <= not (a or b);
    layer1_outputs(9681) <= 1'b1;
    layer1_outputs(9682) <= b;
    layer1_outputs(9683) <= not b or a;
    layer1_outputs(9684) <= not (a or b);
    layer1_outputs(9685) <= a and b;
    layer1_outputs(9686) <= a;
    layer1_outputs(9687) <= not b;
    layer1_outputs(9688) <= b;
    layer1_outputs(9689) <= b;
    layer1_outputs(9690) <= not (a and b);
    layer1_outputs(9691) <= b;
    layer1_outputs(9692) <= not (a or b);
    layer1_outputs(9693) <= b and not a;
    layer1_outputs(9694) <= not a or b;
    layer1_outputs(9695) <= b and not a;
    layer1_outputs(9696) <= b;
    layer1_outputs(9697) <= not a or b;
    layer1_outputs(9698) <= not b;
    layer1_outputs(9699) <= not b;
    layer1_outputs(9700) <= 1'b0;
    layer1_outputs(9701) <= not b;
    layer1_outputs(9702) <= not b or a;
    layer1_outputs(9703) <= 1'b0;
    layer1_outputs(9704) <= a and not b;
    layer1_outputs(9705) <= a;
    layer1_outputs(9706) <= a and not b;
    layer1_outputs(9707) <= b;
    layer1_outputs(9708) <= b and not a;
    layer1_outputs(9709) <= a or b;
    layer1_outputs(9710) <= a;
    layer1_outputs(9711) <= not b;
    layer1_outputs(9712) <= not b or a;
    layer1_outputs(9713) <= not b or a;
    layer1_outputs(9714) <= not a;
    layer1_outputs(9715) <= a;
    layer1_outputs(9716) <= not (a xor b);
    layer1_outputs(9717) <= a;
    layer1_outputs(9718) <= b;
    layer1_outputs(9719) <= not (a and b);
    layer1_outputs(9720) <= not b or a;
    layer1_outputs(9721) <= not a;
    layer1_outputs(9722) <= not (a xor b);
    layer1_outputs(9723) <= not (a xor b);
    layer1_outputs(9724) <= not (a xor b);
    layer1_outputs(9725) <= a or b;
    layer1_outputs(9726) <= not b or a;
    layer1_outputs(9727) <= not b;
    layer1_outputs(9728) <= a;
    layer1_outputs(9729) <= b;
    layer1_outputs(9730) <= a and not b;
    layer1_outputs(9731) <= a or b;
    layer1_outputs(9732) <= b;
    layer1_outputs(9733) <= not (a xor b);
    layer1_outputs(9734) <= 1'b0;
    layer1_outputs(9735) <= b;
    layer1_outputs(9736) <= b;
    layer1_outputs(9737) <= b;
    layer1_outputs(9738) <= not (a and b);
    layer1_outputs(9739) <= not (a or b);
    layer1_outputs(9740) <= not (a or b);
    layer1_outputs(9741) <= a xor b;
    layer1_outputs(9742) <= not b;
    layer1_outputs(9743) <= a and not b;
    layer1_outputs(9744) <= not (a and b);
    layer1_outputs(9745) <= b and not a;
    layer1_outputs(9746) <= a;
    layer1_outputs(9747) <= not (a or b);
    layer1_outputs(9748) <= not (a xor b);
    layer1_outputs(9749) <= not a or b;
    layer1_outputs(9750) <= b;
    layer1_outputs(9751) <= a and not b;
    layer1_outputs(9752) <= not a;
    layer1_outputs(9753) <= not a or b;
    layer1_outputs(9754) <= not (a or b);
    layer1_outputs(9755) <= not b;
    layer1_outputs(9756) <= a and b;
    layer1_outputs(9757) <= not (a and b);
    layer1_outputs(9758) <= a;
    layer1_outputs(9759) <= a;
    layer1_outputs(9760) <= not a;
    layer1_outputs(9761) <= a and b;
    layer1_outputs(9762) <= a or b;
    layer1_outputs(9763) <= b;
    layer1_outputs(9764) <= 1'b1;
    layer1_outputs(9765) <= not a or b;
    layer1_outputs(9766) <= 1'b1;
    layer1_outputs(9767) <= not (a or b);
    layer1_outputs(9768) <= not a;
    layer1_outputs(9769) <= a and b;
    layer1_outputs(9770) <= b and not a;
    layer1_outputs(9771) <= not a or b;
    layer1_outputs(9772) <= b and not a;
    layer1_outputs(9773) <= a;
    layer1_outputs(9774) <= b;
    layer1_outputs(9775) <= a;
    layer1_outputs(9776) <= not a or b;
    layer1_outputs(9777) <= not b;
    layer1_outputs(9778) <= not b;
    layer1_outputs(9779) <= not b;
    layer1_outputs(9780) <= a and b;
    layer1_outputs(9781) <= not (a and b);
    layer1_outputs(9782) <= not b;
    layer1_outputs(9783) <= a;
    layer1_outputs(9784) <= a or b;
    layer1_outputs(9785) <= not (a or b);
    layer1_outputs(9786) <= b;
    layer1_outputs(9787) <= a and b;
    layer1_outputs(9788) <= not a or b;
    layer1_outputs(9789) <= not (a and b);
    layer1_outputs(9790) <= a;
    layer1_outputs(9791) <= a;
    layer1_outputs(9792) <= not a or b;
    layer1_outputs(9793) <= a;
    layer1_outputs(9794) <= not a;
    layer1_outputs(9795) <= a and b;
    layer1_outputs(9796) <= a xor b;
    layer1_outputs(9797) <= not b;
    layer1_outputs(9798) <= not b;
    layer1_outputs(9799) <= a;
    layer1_outputs(9800) <= not (a and b);
    layer1_outputs(9801) <= a;
    layer1_outputs(9802) <= not b or a;
    layer1_outputs(9803) <= a and b;
    layer1_outputs(9804) <= b;
    layer1_outputs(9805) <= b and not a;
    layer1_outputs(9806) <= not a;
    layer1_outputs(9807) <= not (a and b);
    layer1_outputs(9808) <= not a or b;
    layer1_outputs(9809) <= a and not b;
    layer1_outputs(9810) <= a or b;
    layer1_outputs(9811) <= not a or b;
    layer1_outputs(9812) <= a and b;
    layer1_outputs(9813) <= not b;
    layer1_outputs(9814) <= a and b;
    layer1_outputs(9815) <= b and not a;
    layer1_outputs(9816) <= b and not a;
    layer1_outputs(9817) <= a and not b;
    layer1_outputs(9818) <= b;
    layer1_outputs(9819) <= b;
    layer1_outputs(9820) <= a;
    layer1_outputs(9821) <= not (a xor b);
    layer1_outputs(9822) <= not (a or b);
    layer1_outputs(9823) <= not (a and b);
    layer1_outputs(9824) <= a;
    layer1_outputs(9825) <= b;
    layer1_outputs(9826) <= not (a and b);
    layer1_outputs(9827) <= a;
    layer1_outputs(9828) <= a and b;
    layer1_outputs(9829) <= a xor b;
    layer1_outputs(9830) <= a;
    layer1_outputs(9831) <= not a;
    layer1_outputs(9832) <= a;
    layer1_outputs(9833) <= b and not a;
    layer1_outputs(9834) <= not b;
    layer1_outputs(9835) <= not (a or b);
    layer1_outputs(9836) <= 1'b1;
    layer1_outputs(9837) <= a and not b;
    layer1_outputs(9838) <= not b or a;
    layer1_outputs(9839) <= b;
    layer1_outputs(9840) <= not b or a;
    layer1_outputs(9841) <= not b or a;
    layer1_outputs(9842) <= a or b;
    layer1_outputs(9843) <= not (a and b);
    layer1_outputs(9844) <= not b;
    layer1_outputs(9845) <= a and not b;
    layer1_outputs(9846) <= a or b;
    layer1_outputs(9847) <= not a;
    layer1_outputs(9848) <= not (a or b);
    layer1_outputs(9849) <= 1'b1;
    layer1_outputs(9850) <= b;
    layer1_outputs(9851) <= not b;
    layer1_outputs(9852) <= a and not b;
    layer1_outputs(9853) <= not (a and b);
    layer1_outputs(9854) <= a xor b;
    layer1_outputs(9855) <= not b or a;
    layer1_outputs(9856) <= not (a and b);
    layer1_outputs(9857) <= not (a or b);
    layer1_outputs(9858) <= not (a or b);
    layer1_outputs(9859) <= not b or a;
    layer1_outputs(9860) <= not a or b;
    layer1_outputs(9861) <= a;
    layer1_outputs(9862) <= a and b;
    layer1_outputs(9863) <= not b or a;
    layer1_outputs(9864) <= not (a xor b);
    layer1_outputs(9865) <= not a;
    layer1_outputs(9866) <= not a;
    layer1_outputs(9867) <= not (a or b);
    layer1_outputs(9868) <= not a;
    layer1_outputs(9869) <= b and not a;
    layer1_outputs(9870) <= not a or b;
    layer1_outputs(9871) <= a and not b;
    layer1_outputs(9872) <= a;
    layer1_outputs(9873) <= not a;
    layer1_outputs(9874) <= not a or b;
    layer1_outputs(9875) <= not (a or b);
    layer1_outputs(9876) <= b;
    layer1_outputs(9877) <= not (a or b);
    layer1_outputs(9878) <= a;
    layer1_outputs(9879) <= not a or b;
    layer1_outputs(9880) <= a;
    layer1_outputs(9881) <= b and not a;
    layer1_outputs(9882) <= not (a or b);
    layer1_outputs(9883) <= b and not a;
    layer1_outputs(9884) <= not a;
    layer1_outputs(9885) <= not (a and b);
    layer1_outputs(9886) <= not b;
    layer1_outputs(9887) <= 1'b0;
    layer1_outputs(9888) <= b and not a;
    layer1_outputs(9889) <= 1'b0;
    layer1_outputs(9890) <= a xor b;
    layer1_outputs(9891) <= not (a xor b);
    layer1_outputs(9892) <= b and not a;
    layer1_outputs(9893) <= not b or a;
    layer1_outputs(9894) <= a and b;
    layer1_outputs(9895) <= b and not a;
    layer1_outputs(9896) <= not (a or b);
    layer1_outputs(9897) <= not (a and b);
    layer1_outputs(9898) <= a;
    layer1_outputs(9899) <= not a or b;
    layer1_outputs(9900) <= a or b;
    layer1_outputs(9901) <= 1'b1;
    layer1_outputs(9902) <= a or b;
    layer1_outputs(9903) <= a and b;
    layer1_outputs(9904) <= b and not a;
    layer1_outputs(9905) <= not b or a;
    layer1_outputs(9906) <= not b or a;
    layer1_outputs(9907) <= not a;
    layer1_outputs(9908) <= a;
    layer1_outputs(9909) <= not b;
    layer1_outputs(9910) <= a or b;
    layer1_outputs(9911) <= not b or a;
    layer1_outputs(9912) <= not b or a;
    layer1_outputs(9913) <= not b or a;
    layer1_outputs(9914) <= a and not b;
    layer1_outputs(9915) <= not a;
    layer1_outputs(9916) <= not b;
    layer1_outputs(9917) <= not a;
    layer1_outputs(9918) <= 1'b1;
    layer1_outputs(9919) <= not (a xor b);
    layer1_outputs(9920) <= not b;
    layer1_outputs(9921) <= a and not b;
    layer1_outputs(9922) <= not (a and b);
    layer1_outputs(9923) <= not b or a;
    layer1_outputs(9924) <= not b or a;
    layer1_outputs(9925) <= a;
    layer1_outputs(9926) <= a and not b;
    layer1_outputs(9927) <= not b;
    layer1_outputs(9928) <= b and not a;
    layer1_outputs(9929) <= not (a xor b);
    layer1_outputs(9930) <= not (a and b);
    layer1_outputs(9931) <= a xor b;
    layer1_outputs(9932) <= not a;
    layer1_outputs(9933) <= not b;
    layer1_outputs(9934) <= a and not b;
    layer1_outputs(9935) <= not b or a;
    layer1_outputs(9936) <= a and not b;
    layer1_outputs(9937) <= not b;
    layer1_outputs(9938) <= a;
    layer1_outputs(9939) <= b and not a;
    layer1_outputs(9940) <= a;
    layer1_outputs(9941) <= not (a or b);
    layer1_outputs(9942) <= not a or b;
    layer1_outputs(9943) <= b;
    layer1_outputs(9944) <= 1'b0;
    layer1_outputs(9945) <= a and b;
    layer1_outputs(9946) <= not b;
    layer1_outputs(9947) <= 1'b1;
    layer1_outputs(9948) <= a;
    layer1_outputs(9949) <= not a or b;
    layer1_outputs(9950) <= not a or b;
    layer1_outputs(9951) <= not (a and b);
    layer1_outputs(9952) <= not (a or b);
    layer1_outputs(9953) <= a and not b;
    layer1_outputs(9954) <= not (a and b);
    layer1_outputs(9955) <= not b;
    layer1_outputs(9956) <= not (a xor b);
    layer1_outputs(9957) <= a xor b;
    layer1_outputs(9958) <= b;
    layer1_outputs(9959) <= 1'b0;
    layer1_outputs(9960) <= not a or b;
    layer1_outputs(9961) <= a xor b;
    layer1_outputs(9962) <= not (a or b);
    layer1_outputs(9963) <= a;
    layer1_outputs(9964) <= a or b;
    layer1_outputs(9965) <= b and not a;
    layer1_outputs(9966) <= a and b;
    layer1_outputs(9967) <= b;
    layer1_outputs(9968) <= a;
    layer1_outputs(9969) <= not b or a;
    layer1_outputs(9970) <= a or b;
    layer1_outputs(9971) <= b and not a;
    layer1_outputs(9972) <= 1'b0;
    layer1_outputs(9973) <= b;
    layer1_outputs(9974) <= a xor b;
    layer1_outputs(9975) <= a and b;
    layer1_outputs(9976) <= 1'b0;
    layer1_outputs(9977) <= a and not b;
    layer1_outputs(9978) <= 1'b1;
    layer1_outputs(9979) <= a xor b;
    layer1_outputs(9980) <= a;
    layer1_outputs(9981) <= a;
    layer1_outputs(9982) <= not b;
    layer1_outputs(9983) <= a or b;
    layer1_outputs(9984) <= not a;
    layer1_outputs(9985) <= not b or a;
    layer1_outputs(9986) <= not a;
    layer1_outputs(9987) <= not b;
    layer1_outputs(9988) <= not (a or b);
    layer1_outputs(9989) <= not a or b;
    layer1_outputs(9990) <= not (a or b);
    layer1_outputs(9991) <= 1'b0;
    layer1_outputs(9992) <= a or b;
    layer1_outputs(9993) <= not a;
    layer1_outputs(9994) <= a xor b;
    layer1_outputs(9995) <= a or b;
    layer1_outputs(9996) <= b and not a;
    layer1_outputs(9997) <= a or b;
    layer1_outputs(9998) <= not b or a;
    layer1_outputs(9999) <= not b or a;
    layer1_outputs(10000) <= a;
    layer1_outputs(10001) <= a;
    layer1_outputs(10002) <= not a or b;
    layer1_outputs(10003) <= a and b;
    layer1_outputs(10004) <= not a;
    layer1_outputs(10005) <= not b or a;
    layer1_outputs(10006) <= not b or a;
    layer1_outputs(10007) <= not (a xor b);
    layer1_outputs(10008) <= b;
    layer1_outputs(10009) <= a and not b;
    layer1_outputs(10010) <= not (a xor b);
    layer1_outputs(10011) <= not (a and b);
    layer1_outputs(10012) <= a or b;
    layer1_outputs(10013) <= not a;
    layer1_outputs(10014) <= a xor b;
    layer1_outputs(10015) <= a or b;
    layer1_outputs(10016) <= b and not a;
    layer1_outputs(10017) <= not (a and b);
    layer1_outputs(10018) <= not b or a;
    layer1_outputs(10019) <= not b or a;
    layer1_outputs(10020) <= a;
    layer1_outputs(10021) <= a;
    layer1_outputs(10022) <= a;
    layer1_outputs(10023) <= not b;
    layer1_outputs(10024) <= 1'b1;
    layer1_outputs(10025) <= b;
    layer1_outputs(10026) <= a xor b;
    layer1_outputs(10027) <= not a or b;
    layer1_outputs(10028) <= not (a or b);
    layer1_outputs(10029) <= a;
    layer1_outputs(10030) <= not (a or b);
    layer1_outputs(10031) <= a and b;
    layer1_outputs(10032) <= a and b;
    layer1_outputs(10033) <= not b or a;
    layer1_outputs(10034) <= a and b;
    layer1_outputs(10035) <= not a or b;
    layer1_outputs(10036) <= not (a and b);
    layer1_outputs(10037) <= 1'b0;
    layer1_outputs(10038) <= a;
    layer1_outputs(10039) <= a xor b;
    layer1_outputs(10040) <= not b or a;
    layer1_outputs(10041) <= not (a and b);
    layer1_outputs(10042) <= a xor b;
    layer1_outputs(10043) <= not b;
    layer1_outputs(10044) <= b;
    layer1_outputs(10045) <= not (a xor b);
    layer1_outputs(10046) <= a and not b;
    layer1_outputs(10047) <= not b;
    layer1_outputs(10048) <= b;
    layer1_outputs(10049) <= not a;
    layer1_outputs(10050) <= b;
    layer1_outputs(10051) <= b and not a;
    layer1_outputs(10052) <= b and not a;
    layer1_outputs(10053) <= not a;
    layer1_outputs(10054) <= b and not a;
    layer1_outputs(10055) <= not (a xor b);
    layer1_outputs(10056) <= not (a and b);
    layer1_outputs(10057) <= b and not a;
    layer1_outputs(10058) <= not (a xor b);
    layer1_outputs(10059) <= 1'b0;
    layer1_outputs(10060) <= not b;
    layer1_outputs(10061) <= a and not b;
    layer1_outputs(10062) <= not a;
    layer1_outputs(10063) <= a;
    layer1_outputs(10064) <= b and not a;
    layer1_outputs(10065) <= a;
    layer1_outputs(10066) <= a or b;
    layer1_outputs(10067) <= a and not b;
    layer1_outputs(10068) <= not b;
    layer1_outputs(10069) <= not b;
    layer1_outputs(10070) <= not (a and b);
    layer1_outputs(10071) <= not a;
    layer1_outputs(10072) <= a and not b;
    layer1_outputs(10073) <= not a or b;
    layer1_outputs(10074) <= a and b;
    layer1_outputs(10075) <= a;
    layer1_outputs(10076) <= not b;
    layer1_outputs(10077) <= not a or b;
    layer1_outputs(10078) <= not (a xor b);
    layer1_outputs(10079) <= not a or b;
    layer1_outputs(10080) <= a and b;
    layer1_outputs(10081) <= 1'b1;
    layer1_outputs(10082) <= a;
    layer1_outputs(10083) <= b;
    layer1_outputs(10084) <= not b or a;
    layer1_outputs(10085) <= a or b;
    layer1_outputs(10086) <= b and not a;
    layer1_outputs(10087) <= not (a or b);
    layer1_outputs(10088) <= a;
    layer1_outputs(10089) <= a;
    layer1_outputs(10090) <= a xor b;
    layer1_outputs(10091) <= not a or b;
    layer1_outputs(10092) <= b;
    layer1_outputs(10093) <= not b;
    layer1_outputs(10094) <= a and b;
    layer1_outputs(10095) <= not (a xor b);
    layer1_outputs(10096) <= 1'b1;
    layer1_outputs(10097) <= a and b;
    layer1_outputs(10098) <= not a;
    layer1_outputs(10099) <= a and not b;
    layer1_outputs(10100) <= a and not b;
    layer1_outputs(10101) <= not a;
    layer1_outputs(10102) <= b;
    layer1_outputs(10103) <= a xor b;
    layer1_outputs(10104) <= not (a xor b);
    layer1_outputs(10105) <= a or b;
    layer1_outputs(10106) <= a;
    layer1_outputs(10107) <= a and b;
    layer1_outputs(10108) <= b and not a;
    layer1_outputs(10109) <= not (a or b);
    layer1_outputs(10110) <= b;
    layer1_outputs(10111) <= b and not a;
    layer1_outputs(10112) <= not (a xor b);
    layer1_outputs(10113) <= 1'b1;
    layer1_outputs(10114) <= not a;
    layer1_outputs(10115) <= not a or b;
    layer1_outputs(10116) <= b;
    layer1_outputs(10117) <= a and not b;
    layer1_outputs(10118) <= a and not b;
    layer1_outputs(10119) <= a and not b;
    layer1_outputs(10120) <= b and not a;
    layer1_outputs(10121) <= not b or a;
    layer1_outputs(10122) <= 1'b0;
    layer1_outputs(10123) <= not (a or b);
    layer1_outputs(10124) <= not (a or b);
    layer1_outputs(10125) <= 1'b0;
    layer1_outputs(10126) <= not (a xor b);
    layer1_outputs(10127) <= not a or b;
    layer1_outputs(10128) <= a and b;
    layer1_outputs(10129) <= not a;
    layer1_outputs(10130) <= 1'b1;
    layer1_outputs(10131) <= not (a xor b);
    layer1_outputs(10132) <= a xor b;
    layer1_outputs(10133) <= not a;
    layer1_outputs(10134) <= not (a and b);
    layer1_outputs(10135) <= not (a or b);
    layer1_outputs(10136) <= b and not a;
    layer1_outputs(10137) <= 1'b0;
    layer1_outputs(10138) <= not a or b;
    layer1_outputs(10139) <= not b;
    layer1_outputs(10140) <= not (a or b);
    layer1_outputs(10141) <= not (a or b);
    layer1_outputs(10142) <= b;
    layer1_outputs(10143) <= b;
    layer1_outputs(10144) <= a and not b;
    layer1_outputs(10145) <= b and not a;
    layer1_outputs(10146) <= a or b;
    layer1_outputs(10147) <= b and not a;
    layer1_outputs(10148) <= not a or b;
    layer1_outputs(10149) <= a or b;
    layer1_outputs(10150) <= not b;
    layer1_outputs(10151) <= a;
    layer1_outputs(10152) <= not b;
    layer1_outputs(10153) <= not b;
    layer1_outputs(10154) <= not a or b;
    layer1_outputs(10155) <= 1'b0;
    layer1_outputs(10156) <= not (a xor b);
    layer1_outputs(10157) <= a xor b;
    layer1_outputs(10158) <= not (a or b);
    layer1_outputs(10159) <= a or b;
    layer1_outputs(10160) <= not a;
    layer1_outputs(10161) <= not b or a;
    layer1_outputs(10162) <= b;
    layer1_outputs(10163) <= not a;
    layer1_outputs(10164) <= a and b;
    layer1_outputs(10165) <= a and not b;
    layer1_outputs(10166) <= not a;
    layer1_outputs(10167) <= not b;
    layer1_outputs(10168) <= not b;
    layer1_outputs(10169) <= not (a or b);
    layer1_outputs(10170) <= a;
    layer1_outputs(10171) <= not a or b;
    layer1_outputs(10172) <= a and b;
    layer1_outputs(10173) <= a;
    layer1_outputs(10174) <= not a or b;
    layer1_outputs(10175) <= not (a or b);
    layer1_outputs(10176) <= not a or b;
    layer1_outputs(10177) <= not a or b;
    layer1_outputs(10178) <= a and b;
    layer1_outputs(10179) <= b;
    layer1_outputs(10180) <= not (a and b);
    layer1_outputs(10181) <= a or b;
    layer1_outputs(10182) <= not b or a;
    layer1_outputs(10183) <= a and not b;
    layer1_outputs(10184) <= not a;
    layer1_outputs(10185) <= b and not a;
    layer1_outputs(10186) <= a or b;
    layer1_outputs(10187) <= not (a or b);
    layer1_outputs(10188) <= b;
    layer1_outputs(10189) <= not (a and b);
    layer1_outputs(10190) <= b and not a;
    layer1_outputs(10191) <= a or b;
    layer1_outputs(10192) <= not (a and b);
    layer1_outputs(10193) <= not b or a;
    layer1_outputs(10194) <= not (a or b);
    layer1_outputs(10195) <= not (a or b);
    layer1_outputs(10196) <= not b or a;
    layer1_outputs(10197) <= not a or b;
    layer1_outputs(10198) <= not b or a;
    layer1_outputs(10199) <= not b or a;
    layer1_outputs(10200) <= not b;
    layer1_outputs(10201) <= a and not b;
    layer1_outputs(10202) <= not b;
    layer1_outputs(10203) <= a and not b;
    layer1_outputs(10204) <= a;
    layer1_outputs(10205) <= not a or b;
    layer1_outputs(10206) <= not b;
    layer1_outputs(10207) <= 1'b1;
    layer1_outputs(10208) <= a and not b;
    layer1_outputs(10209) <= not b or a;
    layer1_outputs(10210) <= not (a xor b);
    layer1_outputs(10211) <= a and b;
    layer1_outputs(10212) <= 1'b0;
    layer1_outputs(10213) <= not (a or b);
    layer1_outputs(10214) <= a and b;
    layer1_outputs(10215) <= not b or a;
    layer1_outputs(10216) <= a;
    layer1_outputs(10217) <= a and b;
    layer1_outputs(10218) <= not b or a;
    layer1_outputs(10219) <= not b or a;
    layer1_outputs(10220) <= a;
    layer1_outputs(10221) <= b;
    layer1_outputs(10222) <= 1'b1;
    layer1_outputs(10223) <= a or b;
    layer1_outputs(10224) <= a and b;
    layer1_outputs(10225) <= a and b;
    layer1_outputs(10226) <= b;
    layer1_outputs(10227) <= not (a xor b);
    layer1_outputs(10228) <= not (a and b);
    layer1_outputs(10229) <= b;
    layer1_outputs(10230) <= not b;
    layer1_outputs(10231) <= not (a or b);
    layer1_outputs(10232) <= not a;
    layer1_outputs(10233) <= a and not b;
    layer1_outputs(10234) <= a and b;
    layer1_outputs(10235) <= not (a or b);
    layer1_outputs(10236) <= not (a or b);
    layer1_outputs(10237) <= not (a and b);
    layer1_outputs(10238) <= not (a or b);
    layer1_outputs(10239) <= not b or a;
    layer2_outputs(0) <= not (a or b);
    layer2_outputs(1) <= not a;
    layer2_outputs(2) <= b;
    layer2_outputs(3) <= 1'b1;
    layer2_outputs(4) <= a and b;
    layer2_outputs(5) <= a and not b;
    layer2_outputs(6) <= not (a and b);
    layer2_outputs(7) <= a xor b;
    layer2_outputs(8) <= not a or b;
    layer2_outputs(9) <= a;
    layer2_outputs(10) <= b and not a;
    layer2_outputs(11) <= not a or b;
    layer2_outputs(12) <= not b or a;
    layer2_outputs(13) <= not (a and b);
    layer2_outputs(14) <= not (a xor b);
    layer2_outputs(15) <= a and not b;
    layer2_outputs(16) <= not (a or b);
    layer2_outputs(17) <= not (a and b);
    layer2_outputs(18) <= b and not a;
    layer2_outputs(19) <= not (a or b);
    layer2_outputs(20) <= not (a xor b);
    layer2_outputs(21) <= a xor b;
    layer2_outputs(22) <= not b;
    layer2_outputs(23) <= not a;
    layer2_outputs(24) <= not b;
    layer2_outputs(25) <= not (a and b);
    layer2_outputs(26) <= not b;
    layer2_outputs(27) <= not (a and b);
    layer2_outputs(28) <= b and not a;
    layer2_outputs(29) <= b and not a;
    layer2_outputs(30) <= not a;
    layer2_outputs(31) <= b;
    layer2_outputs(32) <= not a or b;
    layer2_outputs(33) <= a xor b;
    layer2_outputs(34) <= not (a or b);
    layer2_outputs(35) <= not b;
    layer2_outputs(36) <= a or b;
    layer2_outputs(37) <= b;
    layer2_outputs(38) <= 1'b0;
    layer2_outputs(39) <= b;
    layer2_outputs(40) <= a or b;
    layer2_outputs(41) <= a xor b;
    layer2_outputs(42) <= b;
    layer2_outputs(43) <= not (a or b);
    layer2_outputs(44) <= not (a xor b);
    layer2_outputs(45) <= b;
    layer2_outputs(46) <= a;
    layer2_outputs(47) <= a or b;
    layer2_outputs(48) <= a;
    layer2_outputs(49) <= a and b;
    layer2_outputs(50) <= a and b;
    layer2_outputs(51) <= not b or a;
    layer2_outputs(52) <= a and b;
    layer2_outputs(53) <= not a;
    layer2_outputs(54) <= not (a or b);
    layer2_outputs(55) <= a and not b;
    layer2_outputs(56) <= not (a and b);
    layer2_outputs(57) <= not (a and b);
    layer2_outputs(58) <= b;
    layer2_outputs(59) <= a;
    layer2_outputs(60) <= a and b;
    layer2_outputs(61) <= not (a and b);
    layer2_outputs(62) <= not b or a;
    layer2_outputs(63) <= not b or a;
    layer2_outputs(64) <= a xor b;
    layer2_outputs(65) <= not (a and b);
    layer2_outputs(66) <= b and not a;
    layer2_outputs(67) <= not b or a;
    layer2_outputs(68) <= not b;
    layer2_outputs(69) <= not (a xor b);
    layer2_outputs(70) <= not b;
    layer2_outputs(71) <= not (a xor b);
    layer2_outputs(72) <= a xor b;
    layer2_outputs(73) <= b;
    layer2_outputs(74) <= not (a or b);
    layer2_outputs(75) <= not (a or b);
    layer2_outputs(76) <= b;
    layer2_outputs(77) <= not a;
    layer2_outputs(78) <= not b;
    layer2_outputs(79) <= b;
    layer2_outputs(80) <= not b;
    layer2_outputs(81) <= b;
    layer2_outputs(82) <= b;
    layer2_outputs(83) <= b;
    layer2_outputs(84) <= not (a and b);
    layer2_outputs(85) <= a xor b;
    layer2_outputs(86) <= not (a and b);
    layer2_outputs(87) <= not a;
    layer2_outputs(88) <= not (a or b);
    layer2_outputs(89) <= a;
    layer2_outputs(90) <= not (a xor b);
    layer2_outputs(91) <= 1'b0;
    layer2_outputs(92) <= not (a xor b);
    layer2_outputs(93) <= not b;
    layer2_outputs(94) <= a and b;
    layer2_outputs(95) <= not b or a;
    layer2_outputs(96) <= a and b;
    layer2_outputs(97) <= not b;
    layer2_outputs(98) <= not a;
    layer2_outputs(99) <= not b;
    layer2_outputs(100) <= a;
    layer2_outputs(101) <= a or b;
    layer2_outputs(102) <= not a or b;
    layer2_outputs(103) <= not b;
    layer2_outputs(104) <= a xor b;
    layer2_outputs(105) <= not (a xor b);
    layer2_outputs(106) <= not a;
    layer2_outputs(107) <= not (a xor b);
    layer2_outputs(108) <= a or b;
    layer2_outputs(109) <= a and not b;
    layer2_outputs(110) <= a or b;
    layer2_outputs(111) <= not b;
    layer2_outputs(112) <= b and not a;
    layer2_outputs(113) <= b and not a;
    layer2_outputs(114) <= not (a or b);
    layer2_outputs(115) <= a or b;
    layer2_outputs(116) <= a;
    layer2_outputs(117) <= a and not b;
    layer2_outputs(118) <= 1'b1;
    layer2_outputs(119) <= a;
    layer2_outputs(120) <= a xor b;
    layer2_outputs(121) <= a;
    layer2_outputs(122) <= a;
    layer2_outputs(123) <= b and not a;
    layer2_outputs(124) <= a and b;
    layer2_outputs(125) <= b;
    layer2_outputs(126) <= not b;
    layer2_outputs(127) <= not a or b;
    layer2_outputs(128) <= b and not a;
    layer2_outputs(129) <= not b or a;
    layer2_outputs(130) <= not b;
    layer2_outputs(131) <= not a;
    layer2_outputs(132) <= 1'b1;
    layer2_outputs(133) <= 1'b1;
    layer2_outputs(134) <= not b;
    layer2_outputs(135) <= a;
    layer2_outputs(136) <= not (a and b);
    layer2_outputs(137) <= a xor b;
    layer2_outputs(138) <= not (a and b);
    layer2_outputs(139) <= b;
    layer2_outputs(140) <= not (a or b);
    layer2_outputs(141) <= a;
    layer2_outputs(142) <= a xor b;
    layer2_outputs(143) <= a;
    layer2_outputs(144) <= not a;
    layer2_outputs(145) <= not (a or b);
    layer2_outputs(146) <= not a or b;
    layer2_outputs(147) <= not (a xor b);
    layer2_outputs(148) <= not b or a;
    layer2_outputs(149) <= not a;
    layer2_outputs(150) <= not (a or b);
    layer2_outputs(151) <= not b;
    layer2_outputs(152) <= a or b;
    layer2_outputs(153) <= not a;
    layer2_outputs(154) <= not a or b;
    layer2_outputs(155) <= 1'b0;
    layer2_outputs(156) <= a and b;
    layer2_outputs(157) <= not b or a;
    layer2_outputs(158) <= b;
    layer2_outputs(159) <= not (a or b);
    layer2_outputs(160) <= a and b;
    layer2_outputs(161) <= a and b;
    layer2_outputs(162) <= not a;
    layer2_outputs(163) <= not (a xor b);
    layer2_outputs(164) <= b;
    layer2_outputs(165) <= a;
    layer2_outputs(166) <= a or b;
    layer2_outputs(167) <= a;
    layer2_outputs(168) <= a and b;
    layer2_outputs(169) <= b and not a;
    layer2_outputs(170) <= a;
    layer2_outputs(171) <= a;
    layer2_outputs(172) <= 1'b1;
    layer2_outputs(173) <= not b;
    layer2_outputs(174) <= not b;
    layer2_outputs(175) <= b;
    layer2_outputs(176) <= a xor b;
    layer2_outputs(177) <= a and b;
    layer2_outputs(178) <= a;
    layer2_outputs(179) <= a and b;
    layer2_outputs(180) <= a;
    layer2_outputs(181) <= b and not a;
    layer2_outputs(182) <= not (a or b);
    layer2_outputs(183) <= not b;
    layer2_outputs(184) <= a and b;
    layer2_outputs(185) <= not b;
    layer2_outputs(186) <= a and not b;
    layer2_outputs(187) <= not b;
    layer2_outputs(188) <= b and not a;
    layer2_outputs(189) <= a and b;
    layer2_outputs(190) <= a;
    layer2_outputs(191) <= 1'b0;
    layer2_outputs(192) <= a;
    layer2_outputs(193) <= b;
    layer2_outputs(194) <= a;
    layer2_outputs(195) <= not b or a;
    layer2_outputs(196) <= not a or b;
    layer2_outputs(197) <= not b;
    layer2_outputs(198) <= not b;
    layer2_outputs(199) <= b;
    layer2_outputs(200) <= not a or b;
    layer2_outputs(201) <= not a;
    layer2_outputs(202) <= not a;
    layer2_outputs(203) <= not b;
    layer2_outputs(204) <= not (a and b);
    layer2_outputs(205) <= b;
    layer2_outputs(206) <= not a;
    layer2_outputs(207) <= not b or a;
    layer2_outputs(208) <= a;
    layer2_outputs(209) <= not a;
    layer2_outputs(210) <= not (a or b);
    layer2_outputs(211) <= b;
    layer2_outputs(212) <= a;
    layer2_outputs(213) <= a or b;
    layer2_outputs(214) <= a and b;
    layer2_outputs(215) <= b and not a;
    layer2_outputs(216) <= a;
    layer2_outputs(217) <= a and not b;
    layer2_outputs(218) <= a xor b;
    layer2_outputs(219) <= b and not a;
    layer2_outputs(220) <= not (a and b);
    layer2_outputs(221) <= a or b;
    layer2_outputs(222) <= not a;
    layer2_outputs(223) <= not b or a;
    layer2_outputs(224) <= not (a and b);
    layer2_outputs(225) <= 1'b1;
    layer2_outputs(226) <= a xor b;
    layer2_outputs(227) <= not a or b;
    layer2_outputs(228) <= not (a xor b);
    layer2_outputs(229) <= not (a and b);
    layer2_outputs(230) <= a or b;
    layer2_outputs(231) <= 1'b0;
    layer2_outputs(232) <= a and not b;
    layer2_outputs(233) <= a or b;
    layer2_outputs(234) <= b and not a;
    layer2_outputs(235) <= not (a xor b);
    layer2_outputs(236) <= not b or a;
    layer2_outputs(237) <= not a or b;
    layer2_outputs(238) <= a or b;
    layer2_outputs(239) <= b;
    layer2_outputs(240) <= not b;
    layer2_outputs(241) <= b and not a;
    layer2_outputs(242) <= not a;
    layer2_outputs(243) <= not b or a;
    layer2_outputs(244) <= a and b;
    layer2_outputs(245) <= not b or a;
    layer2_outputs(246) <= a or b;
    layer2_outputs(247) <= 1'b1;
    layer2_outputs(248) <= b;
    layer2_outputs(249) <= not (a xor b);
    layer2_outputs(250) <= b;
    layer2_outputs(251) <= a and b;
    layer2_outputs(252) <= a and not b;
    layer2_outputs(253) <= not a;
    layer2_outputs(254) <= 1'b1;
    layer2_outputs(255) <= a and b;
    layer2_outputs(256) <= 1'b0;
    layer2_outputs(257) <= not b;
    layer2_outputs(258) <= not b;
    layer2_outputs(259) <= not a;
    layer2_outputs(260) <= b;
    layer2_outputs(261) <= b;
    layer2_outputs(262) <= 1'b1;
    layer2_outputs(263) <= 1'b0;
    layer2_outputs(264) <= a or b;
    layer2_outputs(265) <= a;
    layer2_outputs(266) <= a and not b;
    layer2_outputs(267) <= not (a xor b);
    layer2_outputs(268) <= not (a and b);
    layer2_outputs(269) <= a;
    layer2_outputs(270) <= 1'b0;
    layer2_outputs(271) <= b;
    layer2_outputs(272) <= b and not a;
    layer2_outputs(273) <= a and not b;
    layer2_outputs(274) <= b;
    layer2_outputs(275) <= not a;
    layer2_outputs(276) <= a or b;
    layer2_outputs(277) <= b;
    layer2_outputs(278) <= b;
    layer2_outputs(279) <= not a;
    layer2_outputs(280) <= not a or b;
    layer2_outputs(281) <= not a or b;
    layer2_outputs(282) <= a and not b;
    layer2_outputs(283) <= not a;
    layer2_outputs(284) <= not b or a;
    layer2_outputs(285) <= not (a or b);
    layer2_outputs(286) <= not a;
    layer2_outputs(287) <= not b or a;
    layer2_outputs(288) <= not a;
    layer2_outputs(289) <= not (a and b);
    layer2_outputs(290) <= b;
    layer2_outputs(291) <= not b or a;
    layer2_outputs(292) <= not b;
    layer2_outputs(293) <= not b or a;
    layer2_outputs(294) <= b and not a;
    layer2_outputs(295) <= not (a xor b);
    layer2_outputs(296) <= a and b;
    layer2_outputs(297) <= not a;
    layer2_outputs(298) <= b;
    layer2_outputs(299) <= a;
    layer2_outputs(300) <= a xor b;
    layer2_outputs(301) <= not a;
    layer2_outputs(302) <= a;
    layer2_outputs(303) <= not (a and b);
    layer2_outputs(304) <= not a;
    layer2_outputs(305) <= a;
    layer2_outputs(306) <= b and not a;
    layer2_outputs(307) <= a or b;
    layer2_outputs(308) <= 1'b1;
    layer2_outputs(309) <= not (a or b);
    layer2_outputs(310) <= not a;
    layer2_outputs(311) <= 1'b0;
    layer2_outputs(312) <= not b or a;
    layer2_outputs(313) <= b and not a;
    layer2_outputs(314) <= not (a or b);
    layer2_outputs(315) <= a or b;
    layer2_outputs(316) <= a;
    layer2_outputs(317) <= a;
    layer2_outputs(318) <= b;
    layer2_outputs(319) <= b and not a;
    layer2_outputs(320) <= not a or b;
    layer2_outputs(321) <= b and not a;
    layer2_outputs(322) <= a and b;
    layer2_outputs(323) <= b;
    layer2_outputs(324) <= not b or a;
    layer2_outputs(325) <= 1'b1;
    layer2_outputs(326) <= a;
    layer2_outputs(327) <= not (a xor b);
    layer2_outputs(328) <= b and not a;
    layer2_outputs(329) <= not a;
    layer2_outputs(330) <= not (a or b);
    layer2_outputs(331) <= a;
    layer2_outputs(332) <= not a;
    layer2_outputs(333) <= b and not a;
    layer2_outputs(334) <= not b;
    layer2_outputs(335) <= a or b;
    layer2_outputs(336) <= not b or a;
    layer2_outputs(337) <= 1'b1;
    layer2_outputs(338) <= a;
    layer2_outputs(339) <= b;
    layer2_outputs(340) <= b and not a;
    layer2_outputs(341) <= b and not a;
    layer2_outputs(342) <= a and b;
    layer2_outputs(343) <= b;
    layer2_outputs(344) <= not a;
    layer2_outputs(345) <= not b;
    layer2_outputs(346) <= a and b;
    layer2_outputs(347) <= not a or b;
    layer2_outputs(348) <= not a;
    layer2_outputs(349) <= b and not a;
    layer2_outputs(350) <= a;
    layer2_outputs(351) <= not b or a;
    layer2_outputs(352) <= b;
    layer2_outputs(353) <= a;
    layer2_outputs(354) <= not b or a;
    layer2_outputs(355) <= a;
    layer2_outputs(356) <= not b or a;
    layer2_outputs(357) <= not (a or b);
    layer2_outputs(358) <= not a or b;
    layer2_outputs(359) <= b and not a;
    layer2_outputs(360) <= a;
    layer2_outputs(361) <= b and not a;
    layer2_outputs(362) <= not (a and b);
    layer2_outputs(363) <= a;
    layer2_outputs(364) <= b;
    layer2_outputs(365) <= not a;
    layer2_outputs(366) <= a and not b;
    layer2_outputs(367) <= not b;
    layer2_outputs(368) <= not b or a;
    layer2_outputs(369) <= not a or b;
    layer2_outputs(370) <= not a;
    layer2_outputs(371) <= not (a xor b);
    layer2_outputs(372) <= a;
    layer2_outputs(373) <= not a;
    layer2_outputs(374) <= a xor b;
    layer2_outputs(375) <= a and not b;
    layer2_outputs(376) <= a and b;
    layer2_outputs(377) <= not b or a;
    layer2_outputs(378) <= b;
    layer2_outputs(379) <= not a;
    layer2_outputs(380) <= a xor b;
    layer2_outputs(381) <= not b or a;
    layer2_outputs(382) <= b;
    layer2_outputs(383) <= not b;
    layer2_outputs(384) <= a or b;
    layer2_outputs(385) <= not (a and b);
    layer2_outputs(386) <= not b;
    layer2_outputs(387) <= a;
    layer2_outputs(388) <= not (a and b);
    layer2_outputs(389) <= a;
    layer2_outputs(390) <= not a;
    layer2_outputs(391) <= not (a xor b);
    layer2_outputs(392) <= not b or a;
    layer2_outputs(393) <= a and b;
    layer2_outputs(394) <= not (a or b);
    layer2_outputs(395) <= a;
    layer2_outputs(396) <= a xor b;
    layer2_outputs(397) <= 1'b0;
    layer2_outputs(398) <= b;
    layer2_outputs(399) <= not a;
    layer2_outputs(400) <= not a;
    layer2_outputs(401) <= not (a and b);
    layer2_outputs(402) <= a and not b;
    layer2_outputs(403) <= not a;
    layer2_outputs(404) <= not b;
    layer2_outputs(405) <= not a or b;
    layer2_outputs(406) <= not (a and b);
    layer2_outputs(407) <= a or b;
    layer2_outputs(408) <= not (a or b);
    layer2_outputs(409) <= 1'b0;
    layer2_outputs(410) <= not (a or b);
    layer2_outputs(411) <= 1'b0;
    layer2_outputs(412) <= b;
    layer2_outputs(413) <= not a or b;
    layer2_outputs(414) <= not b;
    layer2_outputs(415) <= b and not a;
    layer2_outputs(416) <= a and b;
    layer2_outputs(417) <= not b or a;
    layer2_outputs(418) <= a and not b;
    layer2_outputs(419) <= not (a or b);
    layer2_outputs(420) <= a and b;
    layer2_outputs(421) <= b and not a;
    layer2_outputs(422) <= not a or b;
    layer2_outputs(423) <= 1'b0;
    layer2_outputs(424) <= a xor b;
    layer2_outputs(425) <= a xor b;
    layer2_outputs(426) <= not a;
    layer2_outputs(427) <= not a or b;
    layer2_outputs(428) <= not (a and b);
    layer2_outputs(429) <= not (a xor b);
    layer2_outputs(430) <= b;
    layer2_outputs(431) <= b;
    layer2_outputs(432) <= a;
    layer2_outputs(433) <= a xor b;
    layer2_outputs(434) <= a;
    layer2_outputs(435) <= a;
    layer2_outputs(436) <= a and not b;
    layer2_outputs(437) <= b and not a;
    layer2_outputs(438) <= not a;
    layer2_outputs(439) <= a and b;
    layer2_outputs(440) <= not a or b;
    layer2_outputs(441) <= not b;
    layer2_outputs(442) <= a and b;
    layer2_outputs(443) <= a and not b;
    layer2_outputs(444) <= 1'b0;
    layer2_outputs(445) <= a or b;
    layer2_outputs(446) <= b;
    layer2_outputs(447) <= b and not a;
    layer2_outputs(448) <= 1'b0;
    layer2_outputs(449) <= not a;
    layer2_outputs(450) <= not b;
    layer2_outputs(451) <= b and not a;
    layer2_outputs(452) <= a;
    layer2_outputs(453) <= not b;
    layer2_outputs(454) <= not a;
    layer2_outputs(455) <= 1'b0;
    layer2_outputs(456) <= b and not a;
    layer2_outputs(457) <= not b;
    layer2_outputs(458) <= a;
    layer2_outputs(459) <= a and not b;
    layer2_outputs(460) <= b;
    layer2_outputs(461) <= a or b;
    layer2_outputs(462) <= b and not a;
    layer2_outputs(463) <= 1'b0;
    layer2_outputs(464) <= not b or a;
    layer2_outputs(465) <= b;
    layer2_outputs(466) <= not a;
    layer2_outputs(467) <= not b;
    layer2_outputs(468) <= a or b;
    layer2_outputs(469) <= 1'b0;
    layer2_outputs(470) <= not a;
    layer2_outputs(471) <= a and b;
    layer2_outputs(472) <= a;
    layer2_outputs(473) <= a and not b;
    layer2_outputs(474) <= 1'b1;
    layer2_outputs(475) <= b;
    layer2_outputs(476) <= b and not a;
    layer2_outputs(477) <= not b;
    layer2_outputs(478) <= not (a xor b);
    layer2_outputs(479) <= a;
    layer2_outputs(480) <= a xor b;
    layer2_outputs(481) <= b;
    layer2_outputs(482) <= not a;
    layer2_outputs(483) <= a and not b;
    layer2_outputs(484) <= a xor b;
    layer2_outputs(485) <= b;
    layer2_outputs(486) <= not (a xor b);
    layer2_outputs(487) <= not b or a;
    layer2_outputs(488) <= not b;
    layer2_outputs(489) <= a and b;
    layer2_outputs(490) <= a;
    layer2_outputs(491) <= b and not a;
    layer2_outputs(492) <= a;
    layer2_outputs(493) <= not a;
    layer2_outputs(494) <= a and b;
    layer2_outputs(495) <= a or b;
    layer2_outputs(496) <= not b or a;
    layer2_outputs(497) <= not (a xor b);
    layer2_outputs(498) <= not a;
    layer2_outputs(499) <= not a;
    layer2_outputs(500) <= not (a and b);
    layer2_outputs(501) <= a and not b;
    layer2_outputs(502) <= b;
    layer2_outputs(503) <= not b;
    layer2_outputs(504) <= a;
    layer2_outputs(505) <= not (a and b);
    layer2_outputs(506) <= not a;
    layer2_outputs(507) <= not (a xor b);
    layer2_outputs(508) <= not (a or b);
    layer2_outputs(509) <= not a;
    layer2_outputs(510) <= not b or a;
    layer2_outputs(511) <= a;
    layer2_outputs(512) <= not a or b;
    layer2_outputs(513) <= a and b;
    layer2_outputs(514) <= a;
    layer2_outputs(515) <= not a;
    layer2_outputs(516) <= b and not a;
    layer2_outputs(517) <= b and not a;
    layer2_outputs(518) <= not a;
    layer2_outputs(519) <= not a;
    layer2_outputs(520) <= a xor b;
    layer2_outputs(521) <= a;
    layer2_outputs(522) <= a;
    layer2_outputs(523) <= not b;
    layer2_outputs(524) <= not a or b;
    layer2_outputs(525) <= a and not b;
    layer2_outputs(526) <= not a or b;
    layer2_outputs(527) <= b;
    layer2_outputs(528) <= not a or b;
    layer2_outputs(529) <= not (a and b);
    layer2_outputs(530) <= not (a and b);
    layer2_outputs(531) <= a xor b;
    layer2_outputs(532) <= a;
    layer2_outputs(533) <= a and not b;
    layer2_outputs(534) <= not a;
    layer2_outputs(535) <= not b;
    layer2_outputs(536) <= not (a xor b);
    layer2_outputs(537) <= not a or b;
    layer2_outputs(538) <= not (a and b);
    layer2_outputs(539) <= b and not a;
    layer2_outputs(540) <= b;
    layer2_outputs(541) <= not a;
    layer2_outputs(542) <= a;
    layer2_outputs(543) <= not b;
    layer2_outputs(544) <= a;
    layer2_outputs(545) <= a and b;
    layer2_outputs(546) <= b and not a;
    layer2_outputs(547) <= a xor b;
    layer2_outputs(548) <= b;
    layer2_outputs(549) <= b;
    layer2_outputs(550) <= not (a or b);
    layer2_outputs(551) <= a and not b;
    layer2_outputs(552) <= a and b;
    layer2_outputs(553) <= a;
    layer2_outputs(554) <= b and not a;
    layer2_outputs(555) <= not b;
    layer2_outputs(556) <= a xor b;
    layer2_outputs(557) <= a and b;
    layer2_outputs(558) <= 1'b0;
    layer2_outputs(559) <= not (a xor b);
    layer2_outputs(560) <= b;
    layer2_outputs(561) <= not b or a;
    layer2_outputs(562) <= a;
    layer2_outputs(563) <= a xor b;
    layer2_outputs(564) <= b and not a;
    layer2_outputs(565) <= b;
    layer2_outputs(566) <= not (a and b);
    layer2_outputs(567) <= not (a or b);
    layer2_outputs(568) <= b;
    layer2_outputs(569) <= b;
    layer2_outputs(570) <= a xor b;
    layer2_outputs(571) <= a;
    layer2_outputs(572) <= b;
    layer2_outputs(573) <= not (a or b);
    layer2_outputs(574) <= not a;
    layer2_outputs(575) <= a;
    layer2_outputs(576) <= a;
    layer2_outputs(577) <= a;
    layer2_outputs(578) <= not a or b;
    layer2_outputs(579) <= not b or a;
    layer2_outputs(580) <= not (a xor b);
    layer2_outputs(581) <= a;
    layer2_outputs(582) <= b;
    layer2_outputs(583) <= not a;
    layer2_outputs(584) <= not a or b;
    layer2_outputs(585) <= not b or a;
    layer2_outputs(586) <= b and not a;
    layer2_outputs(587) <= b;
    layer2_outputs(588) <= not a;
    layer2_outputs(589) <= a;
    layer2_outputs(590) <= not b or a;
    layer2_outputs(591) <= a and b;
    layer2_outputs(592) <= 1'b0;
    layer2_outputs(593) <= a or b;
    layer2_outputs(594) <= a and not b;
    layer2_outputs(595) <= not b;
    layer2_outputs(596) <= a;
    layer2_outputs(597) <= not a or b;
    layer2_outputs(598) <= not a or b;
    layer2_outputs(599) <= not (a xor b);
    layer2_outputs(600) <= not (a or b);
    layer2_outputs(601) <= a and b;
    layer2_outputs(602) <= a;
    layer2_outputs(603) <= a xor b;
    layer2_outputs(604) <= not (a and b);
    layer2_outputs(605) <= not b;
    layer2_outputs(606) <= a and not b;
    layer2_outputs(607) <= not b;
    layer2_outputs(608) <= b;
    layer2_outputs(609) <= not (a and b);
    layer2_outputs(610) <= b;
    layer2_outputs(611) <= not b;
    layer2_outputs(612) <= not (a xor b);
    layer2_outputs(613) <= not a;
    layer2_outputs(614) <= not (a or b);
    layer2_outputs(615) <= b and not a;
    layer2_outputs(616) <= not b;
    layer2_outputs(617) <= not a;
    layer2_outputs(618) <= not (a or b);
    layer2_outputs(619) <= a;
    layer2_outputs(620) <= a or b;
    layer2_outputs(621) <= b;
    layer2_outputs(622) <= a;
    layer2_outputs(623) <= not b;
    layer2_outputs(624) <= not b or a;
    layer2_outputs(625) <= not (a or b);
    layer2_outputs(626) <= a and b;
    layer2_outputs(627) <= a and b;
    layer2_outputs(628) <= b;
    layer2_outputs(629) <= a and b;
    layer2_outputs(630) <= not b;
    layer2_outputs(631) <= not a;
    layer2_outputs(632) <= b;
    layer2_outputs(633) <= b and not a;
    layer2_outputs(634) <= not a;
    layer2_outputs(635) <= not a;
    layer2_outputs(636) <= b and not a;
    layer2_outputs(637) <= not b or a;
    layer2_outputs(638) <= a and b;
    layer2_outputs(639) <= not b;
    layer2_outputs(640) <= not b;
    layer2_outputs(641) <= not a;
    layer2_outputs(642) <= not (a and b);
    layer2_outputs(643) <= not b;
    layer2_outputs(644) <= not (a and b);
    layer2_outputs(645) <= not b;
    layer2_outputs(646) <= not (a and b);
    layer2_outputs(647) <= not (a xor b);
    layer2_outputs(648) <= not b or a;
    layer2_outputs(649) <= a;
    layer2_outputs(650) <= not a or b;
    layer2_outputs(651) <= not (a xor b);
    layer2_outputs(652) <= 1'b0;
    layer2_outputs(653) <= not b;
    layer2_outputs(654) <= not b;
    layer2_outputs(655) <= a xor b;
    layer2_outputs(656) <= not (a and b);
    layer2_outputs(657) <= not (a or b);
    layer2_outputs(658) <= a;
    layer2_outputs(659) <= a;
    layer2_outputs(660) <= not (a and b);
    layer2_outputs(661) <= b and not a;
    layer2_outputs(662) <= not (a or b);
    layer2_outputs(663) <= a;
    layer2_outputs(664) <= b;
    layer2_outputs(665) <= a xor b;
    layer2_outputs(666) <= b;
    layer2_outputs(667) <= a;
    layer2_outputs(668) <= b;
    layer2_outputs(669) <= 1'b1;
    layer2_outputs(670) <= 1'b0;
    layer2_outputs(671) <= not (a and b);
    layer2_outputs(672) <= not (a and b);
    layer2_outputs(673) <= a;
    layer2_outputs(674) <= not b or a;
    layer2_outputs(675) <= not (a and b);
    layer2_outputs(676) <= not (a or b);
    layer2_outputs(677) <= not a;
    layer2_outputs(678) <= not a;
    layer2_outputs(679) <= not a;
    layer2_outputs(680) <= b;
    layer2_outputs(681) <= not b or a;
    layer2_outputs(682) <= a;
    layer2_outputs(683) <= not a;
    layer2_outputs(684) <= a and not b;
    layer2_outputs(685) <= a and b;
    layer2_outputs(686) <= not a or b;
    layer2_outputs(687) <= a xor b;
    layer2_outputs(688) <= not (a or b);
    layer2_outputs(689) <= a;
    layer2_outputs(690) <= a and b;
    layer2_outputs(691) <= not b;
    layer2_outputs(692) <= not b;
    layer2_outputs(693) <= a or b;
    layer2_outputs(694) <= 1'b1;
    layer2_outputs(695) <= a or b;
    layer2_outputs(696) <= a or b;
    layer2_outputs(697) <= b;
    layer2_outputs(698) <= a;
    layer2_outputs(699) <= not (a or b);
    layer2_outputs(700) <= a or b;
    layer2_outputs(701) <= not a;
    layer2_outputs(702) <= a or b;
    layer2_outputs(703) <= not b;
    layer2_outputs(704) <= not (a and b);
    layer2_outputs(705) <= a and b;
    layer2_outputs(706) <= 1'b0;
    layer2_outputs(707) <= b and not a;
    layer2_outputs(708) <= not a or b;
    layer2_outputs(709) <= not a or b;
    layer2_outputs(710) <= not (a xor b);
    layer2_outputs(711) <= not (a or b);
    layer2_outputs(712) <= a or b;
    layer2_outputs(713) <= b;
    layer2_outputs(714) <= a;
    layer2_outputs(715) <= not a or b;
    layer2_outputs(716) <= not b;
    layer2_outputs(717) <= not a or b;
    layer2_outputs(718) <= not (a xor b);
    layer2_outputs(719) <= a;
    layer2_outputs(720) <= b and not a;
    layer2_outputs(721) <= a and b;
    layer2_outputs(722) <= a;
    layer2_outputs(723) <= not (a or b);
    layer2_outputs(724) <= a;
    layer2_outputs(725) <= not a or b;
    layer2_outputs(726) <= not (a or b);
    layer2_outputs(727) <= not a;
    layer2_outputs(728) <= b;
    layer2_outputs(729) <= a;
    layer2_outputs(730) <= not b;
    layer2_outputs(731) <= a or b;
    layer2_outputs(732) <= not b;
    layer2_outputs(733) <= not b;
    layer2_outputs(734) <= not a or b;
    layer2_outputs(735) <= a xor b;
    layer2_outputs(736) <= a and not b;
    layer2_outputs(737) <= b;
    layer2_outputs(738) <= not b;
    layer2_outputs(739) <= a;
    layer2_outputs(740) <= a xor b;
    layer2_outputs(741) <= a xor b;
    layer2_outputs(742) <= a and not b;
    layer2_outputs(743) <= not a or b;
    layer2_outputs(744) <= not b;
    layer2_outputs(745) <= not b;
    layer2_outputs(746) <= a;
    layer2_outputs(747) <= a and b;
    layer2_outputs(748) <= a xor b;
    layer2_outputs(749) <= a;
    layer2_outputs(750) <= not (a xor b);
    layer2_outputs(751) <= not a or b;
    layer2_outputs(752) <= not (a and b);
    layer2_outputs(753) <= not b;
    layer2_outputs(754) <= a or b;
    layer2_outputs(755) <= a and not b;
    layer2_outputs(756) <= not a;
    layer2_outputs(757) <= b;
    layer2_outputs(758) <= a and not b;
    layer2_outputs(759) <= b;
    layer2_outputs(760) <= not b or a;
    layer2_outputs(761) <= not (a or b);
    layer2_outputs(762) <= a;
    layer2_outputs(763) <= not a;
    layer2_outputs(764) <= b;
    layer2_outputs(765) <= 1'b0;
    layer2_outputs(766) <= not (a or b);
    layer2_outputs(767) <= a;
    layer2_outputs(768) <= a xor b;
    layer2_outputs(769) <= a and b;
    layer2_outputs(770) <= a;
    layer2_outputs(771) <= not a;
    layer2_outputs(772) <= a or b;
    layer2_outputs(773) <= not (a or b);
    layer2_outputs(774) <= b;
    layer2_outputs(775) <= not (a or b);
    layer2_outputs(776) <= b and not a;
    layer2_outputs(777) <= not b or a;
    layer2_outputs(778) <= a and b;
    layer2_outputs(779) <= not a;
    layer2_outputs(780) <= b;
    layer2_outputs(781) <= not b or a;
    layer2_outputs(782) <= not a;
    layer2_outputs(783) <= not a;
    layer2_outputs(784) <= not b;
    layer2_outputs(785) <= not b or a;
    layer2_outputs(786) <= not (a and b);
    layer2_outputs(787) <= a;
    layer2_outputs(788) <= a and b;
    layer2_outputs(789) <= not a;
    layer2_outputs(790) <= not b;
    layer2_outputs(791) <= not a or b;
    layer2_outputs(792) <= b;
    layer2_outputs(793) <= not b;
    layer2_outputs(794) <= not b or a;
    layer2_outputs(795) <= not (a or b);
    layer2_outputs(796) <= not b;
    layer2_outputs(797) <= not b or a;
    layer2_outputs(798) <= a and not b;
    layer2_outputs(799) <= b;
    layer2_outputs(800) <= a xor b;
    layer2_outputs(801) <= a xor b;
    layer2_outputs(802) <= a or b;
    layer2_outputs(803) <= a and not b;
    layer2_outputs(804) <= not a;
    layer2_outputs(805) <= not b or a;
    layer2_outputs(806) <= not (a xor b);
    layer2_outputs(807) <= 1'b1;
    layer2_outputs(808) <= not (a or b);
    layer2_outputs(809) <= not a or b;
    layer2_outputs(810) <= a or b;
    layer2_outputs(811) <= not b;
    layer2_outputs(812) <= b;
    layer2_outputs(813) <= not b;
    layer2_outputs(814) <= not a or b;
    layer2_outputs(815) <= not (a and b);
    layer2_outputs(816) <= not a or b;
    layer2_outputs(817) <= not (a and b);
    layer2_outputs(818) <= a;
    layer2_outputs(819) <= not a or b;
    layer2_outputs(820) <= a;
    layer2_outputs(821) <= not a;
    layer2_outputs(822) <= a;
    layer2_outputs(823) <= a or b;
    layer2_outputs(824) <= a and b;
    layer2_outputs(825) <= not (a and b);
    layer2_outputs(826) <= not b;
    layer2_outputs(827) <= not (a and b);
    layer2_outputs(828) <= b;
    layer2_outputs(829) <= a;
    layer2_outputs(830) <= not b;
    layer2_outputs(831) <= not b;
    layer2_outputs(832) <= a and b;
    layer2_outputs(833) <= a;
    layer2_outputs(834) <= not a or b;
    layer2_outputs(835) <= not b;
    layer2_outputs(836) <= not a;
    layer2_outputs(837) <= a and b;
    layer2_outputs(838) <= a;
    layer2_outputs(839) <= 1'b0;
    layer2_outputs(840) <= not a;
    layer2_outputs(841) <= not b;
    layer2_outputs(842) <= not a;
    layer2_outputs(843) <= not a or b;
    layer2_outputs(844) <= not (a or b);
    layer2_outputs(845) <= not b;
    layer2_outputs(846) <= not a or b;
    layer2_outputs(847) <= a xor b;
    layer2_outputs(848) <= b;
    layer2_outputs(849) <= a;
    layer2_outputs(850) <= not a;
    layer2_outputs(851) <= a and b;
    layer2_outputs(852) <= not a;
    layer2_outputs(853) <= a xor b;
    layer2_outputs(854) <= b;
    layer2_outputs(855) <= a;
    layer2_outputs(856) <= b;
    layer2_outputs(857) <= not a;
    layer2_outputs(858) <= not a or b;
    layer2_outputs(859) <= not a;
    layer2_outputs(860) <= a xor b;
    layer2_outputs(861) <= not b;
    layer2_outputs(862) <= b and not a;
    layer2_outputs(863) <= b and not a;
    layer2_outputs(864) <= a;
    layer2_outputs(865) <= a xor b;
    layer2_outputs(866) <= a xor b;
    layer2_outputs(867) <= not a;
    layer2_outputs(868) <= a and b;
    layer2_outputs(869) <= a or b;
    layer2_outputs(870) <= not b or a;
    layer2_outputs(871) <= a and b;
    layer2_outputs(872) <= not a;
    layer2_outputs(873) <= not b or a;
    layer2_outputs(874) <= not a or b;
    layer2_outputs(875) <= a or b;
    layer2_outputs(876) <= not a;
    layer2_outputs(877) <= b;
    layer2_outputs(878) <= a xor b;
    layer2_outputs(879) <= a;
    layer2_outputs(880) <= not b;
    layer2_outputs(881) <= a and b;
    layer2_outputs(882) <= not (a xor b);
    layer2_outputs(883) <= a or b;
    layer2_outputs(884) <= not (a xor b);
    layer2_outputs(885) <= b;
    layer2_outputs(886) <= b;
    layer2_outputs(887) <= a;
    layer2_outputs(888) <= not (a xor b);
    layer2_outputs(889) <= a xor b;
    layer2_outputs(890) <= a;
    layer2_outputs(891) <= not a or b;
    layer2_outputs(892) <= a and not b;
    layer2_outputs(893) <= not (a xor b);
    layer2_outputs(894) <= not b;
    layer2_outputs(895) <= not b;
    layer2_outputs(896) <= b;
    layer2_outputs(897) <= not a or b;
    layer2_outputs(898) <= not (a or b);
    layer2_outputs(899) <= not (a xor b);
    layer2_outputs(900) <= not a or b;
    layer2_outputs(901) <= a and not b;
    layer2_outputs(902) <= a and b;
    layer2_outputs(903) <= 1'b1;
    layer2_outputs(904) <= a;
    layer2_outputs(905) <= a xor b;
    layer2_outputs(906) <= not (a or b);
    layer2_outputs(907) <= not a or b;
    layer2_outputs(908) <= b and not a;
    layer2_outputs(909) <= not a or b;
    layer2_outputs(910) <= a and b;
    layer2_outputs(911) <= a;
    layer2_outputs(912) <= not a;
    layer2_outputs(913) <= not a or b;
    layer2_outputs(914) <= a and b;
    layer2_outputs(915) <= a;
    layer2_outputs(916) <= a xor b;
    layer2_outputs(917) <= b;
    layer2_outputs(918) <= a and b;
    layer2_outputs(919) <= a xor b;
    layer2_outputs(920) <= a and not b;
    layer2_outputs(921) <= not b or a;
    layer2_outputs(922) <= not b or a;
    layer2_outputs(923) <= not b or a;
    layer2_outputs(924) <= a or b;
    layer2_outputs(925) <= b;
    layer2_outputs(926) <= a;
    layer2_outputs(927) <= not (a or b);
    layer2_outputs(928) <= a or b;
    layer2_outputs(929) <= b;
    layer2_outputs(930) <= a;
    layer2_outputs(931) <= a or b;
    layer2_outputs(932) <= a xor b;
    layer2_outputs(933) <= not (a and b);
    layer2_outputs(934) <= 1'b0;
    layer2_outputs(935) <= not (a or b);
    layer2_outputs(936) <= not a;
    layer2_outputs(937) <= a;
    layer2_outputs(938) <= a;
    layer2_outputs(939) <= not b;
    layer2_outputs(940) <= not (a and b);
    layer2_outputs(941) <= not b or a;
    layer2_outputs(942) <= a;
    layer2_outputs(943) <= not a;
    layer2_outputs(944) <= a and b;
    layer2_outputs(945) <= b;
    layer2_outputs(946) <= a and not b;
    layer2_outputs(947) <= b;
    layer2_outputs(948) <= not (a or b);
    layer2_outputs(949) <= not (a and b);
    layer2_outputs(950) <= not a;
    layer2_outputs(951) <= not b or a;
    layer2_outputs(952) <= a and b;
    layer2_outputs(953) <= a;
    layer2_outputs(954) <= a and b;
    layer2_outputs(955) <= a;
    layer2_outputs(956) <= not a;
    layer2_outputs(957) <= not b;
    layer2_outputs(958) <= not (a or b);
    layer2_outputs(959) <= b and not a;
    layer2_outputs(960) <= not (a and b);
    layer2_outputs(961) <= not a or b;
    layer2_outputs(962) <= a and b;
    layer2_outputs(963) <= not b or a;
    layer2_outputs(964) <= a;
    layer2_outputs(965) <= not a;
    layer2_outputs(966) <= not (a and b);
    layer2_outputs(967) <= not (a and b);
    layer2_outputs(968) <= not b or a;
    layer2_outputs(969) <= 1'b0;
    layer2_outputs(970) <= a and not b;
    layer2_outputs(971) <= not b;
    layer2_outputs(972) <= not b;
    layer2_outputs(973) <= a and not b;
    layer2_outputs(974) <= not a;
    layer2_outputs(975) <= a or b;
    layer2_outputs(976) <= a;
    layer2_outputs(977) <= a or b;
    layer2_outputs(978) <= b;
    layer2_outputs(979) <= not (a or b);
    layer2_outputs(980) <= a;
    layer2_outputs(981) <= a;
    layer2_outputs(982) <= a;
    layer2_outputs(983) <= a or b;
    layer2_outputs(984) <= a and not b;
    layer2_outputs(985) <= a or b;
    layer2_outputs(986) <= b;
    layer2_outputs(987) <= not a;
    layer2_outputs(988) <= not a;
    layer2_outputs(989) <= not (a or b);
    layer2_outputs(990) <= a and b;
    layer2_outputs(991) <= not b or a;
    layer2_outputs(992) <= a or b;
    layer2_outputs(993) <= a and not b;
    layer2_outputs(994) <= a or b;
    layer2_outputs(995) <= a;
    layer2_outputs(996) <= a xor b;
    layer2_outputs(997) <= not a or b;
    layer2_outputs(998) <= not (a xor b);
    layer2_outputs(999) <= a or b;
    layer2_outputs(1000) <= not b;
    layer2_outputs(1001) <= not a;
    layer2_outputs(1002) <= not a;
    layer2_outputs(1003) <= a;
    layer2_outputs(1004) <= not (a and b);
    layer2_outputs(1005) <= not a;
    layer2_outputs(1006) <= a or b;
    layer2_outputs(1007) <= a and b;
    layer2_outputs(1008) <= not b;
    layer2_outputs(1009) <= a;
    layer2_outputs(1010) <= not a or b;
    layer2_outputs(1011) <= not (a xor b);
    layer2_outputs(1012) <= a;
    layer2_outputs(1013) <= a;
    layer2_outputs(1014) <= not b;
    layer2_outputs(1015) <= not b;
    layer2_outputs(1016) <= b;
    layer2_outputs(1017) <= not b;
    layer2_outputs(1018) <= b;
    layer2_outputs(1019) <= a;
    layer2_outputs(1020) <= b;
    layer2_outputs(1021) <= a and b;
    layer2_outputs(1022) <= not b;
    layer2_outputs(1023) <= not a or b;
    layer2_outputs(1024) <= a and b;
    layer2_outputs(1025) <= a or b;
    layer2_outputs(1026) <= 1'b0;
    layer2_outputs(1027) <= b;
    layer2_outputs(1028) <= not (a and b);
    layer2_outputs(1029) <= a and not b;
    layer2_outputs(1030) <= b and not a;
    layer2_outputs(1031) <= not a;
    layer2_outputs(1032) <= not a or b;
    layer2_outputs(1033) <= not (a xor b);
    layer2_outputs(1034) <= a;
    layer2_outputs(1035) <= not b;
    layer2_outputs(1036) <= not a;
    layer2_outputs(1037) <= b;
    layer2_outputs(1038) <= not a;
    layer2_outputs(1039) <= a;
    layer2_outputs(1040) <= not b or a;
    layer2_outputs(1041) <= b and not a;
    layer2_outputs(1042) <= not b;
    layer2_outputs(1043) <= not b;
    layer2_outputs(1044) <= not b or a;
    layer2_outputs(1045) <= not b;
    layer2_outputs(1046) <= b;
    layer2_outputs(1047) <= not (a or b);
    layer2_outputs(1048) <= a;
    layer2_outputs(1049) <= a;
    layer2_outputs(1050) <= a xor b;
    layer2_outputs(1051) <= 1'b1;
    layer2_outputs(1052) <= a;
    layer2_outputs(1053) <= not (a and b);
    layer2_outputs(1054) <= a or b;
    layer2_outputs(1055) <= a or b;
    layer2_outputs(1056) <= not a;
    layer2_outputs(1057) <= b;
    layer2_outputs(1058) <= a and b;
    layer2_outputs(1059) <= not b or a;
    layer2_outputs(1060) <= a or b;
    layer2_outputs(1061) <= 1'b0;
    layer2_outputs(1062) <= a xor b;
    layer2_outputs(1063) <= not b;
    layer2_outputs(1064) <= a or b;
    layer2_outputs(1065) <= not b or a;
    layer2_outputs(1066) <= a or b;
    layer2_outputs(1067) <= not a;
    layer2_outputs(1068) <= b;
    layer2_outputs(1069) <= b and not a;
    layer2_outputs(1070) <= 1'b1;
    layer2_outputs(1071) <= b;
    layer2_outputs(1072) <= a and not b;
    layer2_outputs(1073) <= 1'b0;
    layer2_outputs(1074) <= not b or a;
    layer2_outputs(1075) <= not a or b;
    layer2_outputs(1076) <= not a;
    layer2_outputs(1077) <= not a;
    layer2_outputs(1078) <= b and not a;
    layer2_outputs(1079) <= a;
    layer2_outputs(1080) <= b and not a;
    layer2_outputs(1081) <= not b;
    layer2_outputs(1082) <= b;
    layer2_outputs(1083) <= b;
    layer2_outputs(1084) <= b;
    layer2_outputs(1085) <= not a;
    layer2_outputs(1086) <= 1'b0;
    layer2_outputs(1087) <= not b or a;
    layer2_outputs(1088) <= not a or b;
    layer2_outputs(1089) <= not a or b;
    layer2_outputs(1090) <= not b;
    layer2_outputs(1091) <= a or b;
    layer2_outputs(1092) <= not (a and b);
    layer2_outputs(1093) <= not a;
    layer2_outputs(1094) <= not b or a;
    layer2_outputs(1095) <= a;
    layer2_outputs(1096) <= a and not b;
    layer2_outputs(1097) <= 1'b1;
    layer2_outputs(1098) <= a and b;
    layer2_outputs(1099) <= b;
    layer2_outputs(1100) <= not a;
    layer2_outputs(1101) <= a and not b;
    layer2_outputs(1102) <= not a or b;
    layer2_outputs(1103) <= a;
    layer2_outputs(1104) <= b and not a;
    layer2_outputs(1105) <= not a;
    layer2_outputs(1106) <= not b or a;
    layer2_outputs(1107) <= not (a xor b);
    layer2_outputs(1108) <= b and not a;
    layer2_outputs(1109) <= not b;
    layer2_outputs(1110) <= a;
    layer2_outputs(1111) <= not a or b;
    layer2_outputs(1112) <= not (a and b);
    layer2_outputs(1113) <= not a;
    layer2_outputs(1114) <= a xor b;
    layer2_outputs(1115) <= not b or a;
    layer2_outputs(1116) <= b and not a;
    layer2_outputs(1117) <= a;
    layer2_outputs(1118) <= not b;
    layer2_outputs(1119) <= a;
    layer2_outputs(1120) <= not (a and b);
    layer2_outputs(1121) <= b and not a;
    layer2_outputs(1122) <= a;
    layer2_outputs(1123) <= not b;
    layer2_outputs(1124) <= a and b;
    layer2_outputs(1125) <= a or b;
    layer2_outputs(1126) <= a or b;
    layer2_outputs(1127) <= not b;
    layer2_outputs(1128) <= not b or a;
    layer2_outputs(1129) <= not b;
    layer2_outputs(1130) <= not a;
    layer2_outputs(1131) <= not a or b;
    layer2_outputs(1132) <= 1'b1;
    layer2_outputs(1133) <= not b or a;
    layer2_outputs(1134) <= not a or b;
    layer2_outputs(1135) <= a or b;
    layer2_outputs(1136) <= not a;
    layer2_outputs(1137) <= a;
    layer2_outputs(1138) <= b;
    layer2_outputs(1139) <= a or b;
    layer2_outputs(1140) <= b and not a;
    layer2_outputs(1141) <= 1'b0;
    layer2_outputs(1142) <= a xor b;
    layer2_outputs(1143) <= b;
    layer2_outputs(1144) <= not (a and b);
    layer2_outputs(1145) <= not a or b;
    layer2_outputs(1146) <= not (a or b);
    layer2_outputs(1147) <= not (a and b);
    layer2_outputs(1148) <= a and not b;
    layer2_outputs(1149) <= not b;
    layer2_outputs(1150) <= not b;
    layer2_outputs(1151) <= a and not b;
    layer2_outputs(1152) <= b;
    layer2_outputs(1153) <= b and not a;
    layer2_outputs(1154) <= not (a xor b);
    layer2_outputs(1155) <= not a;
    layer2_outputs(1156) <= not a or b;
    layer2_outputs(1157) <= not b or a;
    layer2_outputs(1158) <= b and not a;
    layer2_outputs(1159) <= a and not b;
    layer2_outputs(1160) <= b;
    layer2_outputs(1161) <= 1'b0;
    layer2_outputs(1162) <= not a or b;
    layer2_outputs(1163) <= a xor b;
    layer2_outputs(1164) <= not (a xor b);
    layer2_outputs(1165) <= a and not b;
    layer2_outputs(1166) <= not a;
    layer2_outputs(1167) <= a;
    layer2_outputs(1168) <= a;
    layer2_outputs(1169) <= not b;
    layer2_outputs(1170) <= a;
    layer2_outputs(1171) <= a and not b;
    layer2_outputs(1172) <= b;
    layer2_outputs(1173) <= a and not b;
    layer2_outputs(1174) <= not b;
    layer2_outputs(1175) <= b;
    layer2_outputs(1176) <= not a;
    layer2_outputs(1177) <= not (a and b);
    layer2_outputs(1178) <= b and not a;
    layer2_outputs(1179) <= a xor b;
    layer2_outputs(1180) <= b and not a;
    layer2_outputs(1181) <= b;
    layer2_outputs(1182) <= b and not a;
    layer2_outputs(1183) <= b;
    layer2_outputs(1184) <= not (a or b);
    layer2_outputs(1185) <= a and b;
    layer2_outputs(1186) <= a;
    layer2_outputs(1187) <= not b;
    layer2_outputs(1188) <= not a or b;
    layer2_outputs(1189) <= not b;
    layer2_outputs(1190) <= 1'b0;
    layer2_outputs(1191) <= 1'b1;
    layer2_outputs(1192) <= not a;
    layer2_outputs(1193) <= not (a or b);
    layer2_outputs(1194) <= a;
    layer2_outputs(1195) <= not (a xor b);
    layer2_outputs(1196) <= not a;
    layer2_outputs(1197) <= not b or a;
    layer2_outputs(1198) <= not a;
    layer2_outputs(1199) <= a or b;
    layer2_outputs(1200) <= not (a or b);
    layer2_outputs(1201) <= a or b;
    layer2_outputs(1202) <= not a;
    layer2_outputs(1203) <= a;
    layer2_outputs(1204) <= not (a or b);
    layer2_outputs(1205) <= a and b;
    layer2_outputs(1206) <= not a or b;
    layer2_outputs(1207) <= a;
    layer2_outputs(1208) <= a or b;
    layer2_outputs(1209) <= a or b;
    layer2_outputs(1210) <= b;
    layer2_outputs(1211) <= a;
    layer2_outputs(1212) <= not (a and b);
    layer2_outputs(1213) <= not (a or b);
    layer2_outputs(1214) <= a and b;
    layer2_outputs(1215) <= b;
    layer2_outputs(1216) <= a xor b;
    layer2_outputs(1217) <= b;
    layer2_outputs(1218) <= not b;
    layer2_outputs(1219) <= a xor b;
    layer2_outputs(1220) <= a;
    layer2_outputs(1221) <= not (a xor b);
    layer2_outputs(1222) <= not a;
    layer2_outputs(1223) <= not b or a;
    layer2_outputs(1224) <= a and b;
    layer2_outputs(1225) <= not a;
    layer2_outputs(1226) <= not a;
    layer2_outputs(1227) <= a;
    layer2_outputs(1228) <= a;
    layer2_outputs(1229) <= 1'b0;
    layer2_outputs(1230) <= not (a and b);
    layer2_outputs(1231) <= 1'b0;
    layer2_outputs(1232) <= b and not a;
    layer2_outputs(1233) <= a and not b;
    layer2_outputs(1234) <= not a;
    layer2_outputs(1235) <= a and not b;
    layer2_outputs(1236) <= a and not b;
    layer2_outputs(1237) <= not b or a;
    layer2_outputs(1238) <= b and not a;
    layer2_outputs(1239) <= a and not b;
    layer2_outputs(1240) <= a;
    layer2_outputs(1241) <= not b or a;
    layer2_outputs(1242) <= b;
    layer2_outputs(1243) <= b and not a;
    layer2_outputs(1244) <= not b;
    layer2_outputs(1245) <= not a;
    layer2_outputs(1246) <= not b;
    layer2_outputs(1247) <= b and not a;
    layer2_outputs(1248) <= a and b;
    layer2_outputs(1249) <= not a;
    layer2_outputs(1250) <= a and not b;
    layer2_outputs(1251) <= not b or a;
    layer2_outputs(1252) <= not (a and b);
    layer2_outputs(1253) <= not a or b;
    layer2_outputs(1254) <= a;
    layer2_outputs(1255) <= not b or a;
    layer2_outputs(1256) <= b and not a;
    layer2_outputs(1257) <= b and not a;
    layer2_outputs(1258) <= not a;
    layer2_outputs(1259) <= not b or a;
    layer2_outputs(1260) <= not (a and b);
    layer2_outputs(1261) <= not (a and b);
    layer2_outputs(1262) <= not b;
    layer2_outputs(1263) <= not (a or b);
    layer2_outputs(1264) <= b;
    layer2_outputs(1265) <= a and not b;
    layer2_outputs(1266) <= not b;
    layer2_outputs(1267) <= not b or a;
    layer2_outputs(1268) <= not (a xor b);
    layer2_outputs(1269) <= 1'b0;
    layer2_outputs(1270) <= a;
    layer2_outputs(1271) <= not b or a;
    layer2_outputs(1272) <= a xor b;
    layer2_outputs(1273) <= not a;
    layer2_outputs(1274) <= a and b;
    layer2_outputs(1275) <= not (a or b);
    layer2_outputs(1276) <= a;
    layer2_outputs(1277) <= not b;
    layer2_outputs(1278) <= not a;
    layer2_outputs(1279) <= not (a xor b);
    layer2_outputs(1280) <= 1'b1;
    layer2_outputs(1281) <= not b;
    layer2_outputs(1282) <= not (a or b);
    layer2_outputs(1283) <= not b;
    layer2_outputs(1284) <= a and b;
    layer2_outputs(1285) <= not b;
    layer2_outputs(1286) <= a xor b;
    layer2_outputs(1287) <= not a;
    layer2_outputs(1288) <= b and not a;
    layer2_outputs(1289) <= a;
    layer2_outputs(1290) <= not a or b;
    layer2_outputs(1291) <= not (a and b);
    layer2_outputs(1292) <= not a;
    layer2_outputs(1293) <= not b or a;
    layer2_outputs(1294) <= b and not a;
    layer2_outputs(1295) <= a;
    layer2_outputs(1296) <= a or b;
    layer2_outputs(1297) <= a and b;
    layer2_outputs(1298) <= not (a xor b);
    layer2_outputs(1299) <= a xor b;
    layer2_outputs(1300) <= not (a and b);
    layer2_outputs(1301) <= not (a or b);
    layer2_outputs(1302) <= not b or a;
    layer2_outputs(1303) <= a and not b;
    layer2_outputs(1304) <= a xor b;
    layer2_outputs(1305) <= a or b;
    layer2_outputs(1306) <= a;
    layer2_outputs(1307) <= 1'b0;
    layer2_outputs(1308) <= not a;
    layer2_outputs(1309) <= not a;
    layer2_outputs(1310) <= not (a or b);
    layer2_outputs(1311) <= not a;
    layer2_outputs(1312) <= not a;
    layer2_outputs(1313) <= a and b;
    layer2_outputs(1314) <= not a;
    layer2_outputs(1315) <= a xor b;
    layer2_outputs(1316) <= not a;
    layer2_outputs(1317) <= 1'b0;
    layer2_outputs(1318) <= a;
    layer2_outputs(1319) <= not a or b;
    layer2_outputs(1320) <= a xor b;
    layer2_outputs(1321) <= a and not b;
    layer2_outputs(1322) <= not (a xor b);
    layer2_outputs(1323) <= not a or b;
    layer2_outputs(1324) <= not (a and b);
    layer2_outputs(1325) <= not (a or b);
    layer2_outputs(1326) <= a or b;
    layer2_outputs(1327) <= a and b;
    layer2_outputs(1328) <= not b;
    layer2_outputs(1329) <= a xor b;
    layer2_outputs(1330) <= 1'b0;
    layer2_outputs(1331) <= a;
    layer2_outputs(1332) <= a;
    layer2_outputs(1333) <= b and not a;
    layer2_outputs(1334) <= 1'b0;
    layer2_outputs(1335) <= not a;
    layer2_outputs(1336) <= b;
    layer2_outputs(1337) <= a;
    layer2_outputs(1338) <= b and not a;
    layer2_outputs(1339) <= 1'b1;
    layer2_outputs(1340) <= b and not a;
    layer2_outputs(1341) <= not b;
    layer2_outputs(1342) <= a xor b;
    layer2_outputs(1343) <= a and b;
    layer2_outputs(1344) <= b and not a;
    layer2_outputs(1345) <= a;
    layer2_outputs(1346) <= b and not a;
    layer2_outputs(1347) <= b;
    layer2_outputs(1348) <= not b;
    layer2_outputs(1349) <= a and b;
    layer2_outputs(1350) <= not a or b;
    layer2_outputs(1351) <= a and b;
    layer2_outputs(1352) <= a;
    layer2_outputs(1353) <= a and not b;
    layer2_outputs(1354) <= not b or a;
    layer2_outputs(1355) <= not a;
    layer2_outputs(1356) <= not (a and b);
    layer2_outputs(1357) <= a or b;
    layer2_outputs(1358) <= a;
    layer2_outputs(1359) <= 1'b0;
    layer2_outputs(1360) <= not b or a;
    layer2_outputs(1361) <= a and b;
    layer2_outputs(1362) <= b;
    layer2_outputs(1363) <= a;
    layer2_outputs(1364) <= not (a or b);
    layer2_outputs(1365) <= not (a or b);
    layer2_outputs(1366) <= not a;
    layer2_outputs(1367) <= a;
    layer2_outputs(1368) <= b;
    layer2_outputs(1369) <= not a or b;
    layer2_outputs(1370) <= not (a and b);
    layer2_outputs(1371) <= not a;
    layer2_outputs(1372) <= not b or a;
    layer2_outputs(1373) <= not a or b;
    layer2_outputs(1374) <= 1'b0;
    layer2_outputs(1375) <= a;
    layer2_outputs(1376) <= b;
    layer2_outputs(1377) <= not b;
    layer2_outputs(1378) <= not b or a;
    layer2_outputs(1379) <= 1'b0;
    layer2_outputs(1380) <= a or b;
    layer2_outputs(1381) <= a or b;
    layer2_outputs(1382) <= b;
    layer2_outputs(1383) <= a or b;
    layer2_outputs(1384) <= a and not b;
    layer2_outputs(1385) <= a or b;
    layer2_outputs(1386) <= a and not b;
    layer2_outputs(1387) <= not (a or b);
    layer2_outputs(1388) <= b and not a;
    layer2_outputs(1389) <= not a;
    layer2_outputs(1390) <= a;
    layer2_outputs(1391) <= not a or b;
    layer2_outputs(1392) <= b;
    layer2_outputs(1393) <= a and not b;
    layer2_outputs(1394) <= not b;
    layer2_outputs(1395) <= a and b;
    layer2_outputs(1396) <= b and not a;
    layer2_outputs(1397) <= not b or a;
    layer2_outputs(1398) <= not (a or b);
    layer2_outputs(1399) <= not a;
    layer2_outputs(1400) <= not a;
    layer2_outputs(1401) <= 1'b0;
    layer2_outputs(1402) <= a and b;
    layer2_outputs(1403) <= a xor b;
    layer2_outputs(1404) <= not a or b;
    layer2_outputs(1405) <= not b;
    layer2_outputs(1406) <= not b;
    layer2_outputs(1407) <= 1'b0;
    layer2_outputs(1408) <= not (a or b);
    layer2_outputs(1409) <= not b;
    layer2_outputs(1410) <= not a;
    layer2_outputs(1411) <= b;
    layer2_outputs(1412) <= not a;
    layer2_outputs(1413) <= b;
    layer2_outputs(1414) <= a;
    layer2_outputs(1415) <= 1'b0;
    layer2_outputs(1416) <= a;
    layer2_outputs(1417) <= not (a and b);
    layer2_outputs(1418) <= not b or a;
    layer2_outputs(1419) <= a and b;
    layer2_outputs(1420) <= not b;
    layer2_outputs(1421) <= b and not a;
    layer2_outputs(1422) <= b;
    layer2_outputs(1423) <= not b or a;
    layer2_outputs(1424) <= not b;
    layer2_outputs(1425) <= a;
    layer2_outputs(1426) <= not b or a;
    layer2_outputs(1427) <= not a;
    layer2_outputs(1428) <= not b or a;
    layer2_outputs(1429) <= not b;
    layer2_outputs(1430) <= a and not b;
    layer2_outputs(1431) <= a and not b;
    layer2_outputs(1432) <= not b;
    layer2_outputs(1433) <= b;
    layer2_outputs(1434) <= not (a xor b);
    layer2_outputs(1435) <= not (a or b);
    layer2_outputs(1436) <= not b;
    layer2_outputs(1437) <= b;
    layer2_outputs(1438) <= a or b;
    layer2_outputs(1439) <= a and not b;
    layer2_outputs(1440) <= not (a or b);
    layer2_outputs(1441) <= not (a xor b);
    layer2_outputs(1442) <= 1'b1;
    layer2_outputs(1443) <= not a or b;
    layer2_outputs(1444) <= not b or a;
    layer2_outputs(1445) <= not b;
    layer2_outputs(1446) <= a or b;
    layer2_outputs(1447) <= a and b;
    layer2_outputs(1448) <= a;
    layer2_outputs(1449) <= 1'b1;
    layer2_outputs(1450) <= b;
    layer2_outputs(1451) <= b;
    layer2_outputs(1452) <= not (a or b);
    layer2_outputs(1453) <= a and b;
    layer2_outputs(1454) <= b and not a;
    layer2_outputs(1455) <= b;
    layer2_outputs(1456) <= b and not a;
    layer2_outputs(1457) <= a;
    layer2_outputs(1458) <= not b or a;
    layer2_outputs(1459) <= b and not a;
    layer2_outputs(1460) <= a and b;
    layer2_outputs(1461) <= not a;
    layer2_outputs(1462) <= not (a and b);
    layer2_outputs(1463) <= a;
    layer2_outputs(1464) <= not b or a;
    layer2_outputs(1465) <= a and b;
    layer2_outputs(1466) <= not a;
    layer2_outputs(1467) <= a and b;
    layer2_outputs(1468) <= a xor b;
    layer2_outputs(1469) <= not (a or b);
    layer2_outputs(1470) <= a and not b;
    layer2_outputs(1471) <= b;
    layer2_outputs(1472) <= 1'b0;
    layer2_outputs(1473) <= not b or a;
    layer2_outputs(1474) <= b;
    layer2_outputs(1475) <= a and b;
    layer2_outputs(1476) <= a;
    layer2_outputs(1477) <= not a;
    layer2_outputs(1478) <= not b or a;
    layer2_outputs(1479) <= not a or b;
    layer2_outputs(1480) <= a and not b;
    layer2_outputs(1481) <= not a;
    layer2_outputs(1482) <= a and b;
    layer2_outputs(1483) <= b and not a;
    layer2_outputs(1484) <= not b or a;
    layer2_outputs(1485) <= a;
    layer2_outputs(1486) <= b;
    layer2_outputs(1487) <= not b;
    layer2_outputs(1488) <= a or b;
    layer2_outputs(1489) <= 1'b1;
    layer2_outputs(1490) <= a;
    layer2_outputs(1491) <= not a;
    layer2_outputs(1492) <= not a or b;
    layer2_outputs(1493) <= a;
    layer2_outputs(1494) <= not a or b;
    layer2_outputs(1495) <= not a or b;
    layer2_outputs(1496) <= not (a and b);
    layer2_outputs(1497) <= b and not a;
    layer2_outputs(1498) <= not a;
    layer2_outputs(1499) <= a and b;
    layer2_outputs(1500) <= not b or a;
    layer2_outputs(1501) <= not (a xor b);
    layer2_outputs(1502) <= not (a or b);
    layer2_outputs(1503) <= not (a and b);
    layer2_outputs(1504) <= not a;
    layer2_outputs(1505) <= b;
    layer2_outputs(1506) <= b;
    layer2_outputs(1507) <= not b or a;
    layer2_outputs(1508) <= not b;
    layer2_outputs(1509) <= not a;
    layer2_outputs(1510) <= b;
    layer2_outputs(1511) <= a and b;
    layer2_outputs(1512) <= not b or a;
    layer2_outputs(1513) <= not (a or b);
    layer2_outputs(1514) <= a and not b;
    layer2_outputs(1515) <= b and not a;
    layer2_outputs(1516) <= a and b;
    layer2_outputs(1517) <= not a;
    layer2_outputs(1518) <= not (a xor b);
    layer2_outputs(1519) <= not (a or b);
    layer2_outputs(1520) <= not b;
    layer2_outputs(1521) <= a and b;
    layer2_outputs(1522) <= a and b;
    layer2_outputs(1523) <= not b;
    layer2_outputs(1524) <= not a;
    layer2_outputs(1525) <= not b;
    layer2_outputs(1526) <= b and not a;
    layer2_outputs(1527) <= a;
    layer2_outputs(1528) <= not a;
    layer2_outputs(1529) <= not (a xor b);
    layer2_outputs(1530) <= a or b;
    layer2_outputs(1531) <= not b;
    layer2_outputs(1532) <= not (a and b);
    layer2_outputs(1533) <= a or b;
    layer2_outputs(1534) <= a and not b;
    layer2_outputs(1535) <= a xor b;
    layer2_outputs(1536) <= not a;
    layer2_outputs(1537) <= not (a or b);
    layer2_outputs(1538) <= b and not a;
    layer2_outputs(1539) <= not a or b;
    layer2_outputs(1540) <= a and b;
    layer2_outputs(1541) <= not b or a;
    layer2_outputs(1542) <= a and b;
    layer2_outputs(1543) <= b;
    layer2_outputs(1544) <= b and not a;
    layer2_outputs(1545) <= b and not a;
    layer2_outputs(1546) <= not b;
    layer2_outputs(1547) <= b and not a;
    layer2_outputs(1548) <= not a or b;
    layer2_outputs(1549) <= not a or b;
    layer2_outputs(1550) <= a xor b;
    layer2_outputs(1551) <= not b or a;
    layer2_outputs(1552) <= a or b;
    layer2_outputs(1553) <= not a or b;
    layer2_outputs(1554) <= not (a or b);
    layer2_outputs(1555) <= a or b;
    layer2_outputs(1556) <= not (a xor b);
    layer2_outputs(1557) <= a;
    layer2_outputs(1558) <= a and not b;
    layer2_outputs(1559) <= a and not b;
    layer2_outputs(1560) <= not b or a;
    layer2_outputs(1561) <= b and not a;
    layer2_outputs(1562) <= a and not b;
    layer2_outputs(1563) <= a;
    layer2_outputs(1564) <= b and not a;
    layer2_outputs(1565) <= not a;
    layer2_outputs(1566) <= not (a xor b);
    layer2_outputs(1567) <= b;
    layer2_outputs(1568) <= b;
    layer2_outputs(1569) <= b and not a;
    layer2_outputs(1570) <= a and not b;
    layer2_outputs(1571) <= b;
    layer2_outputs(1572) <= not (a xor b);
    layer2_outputs(1573) <= not b;
    layer2_outputs(1574) <= not b or a;
    layer2_outputs(1575) <= a or b;
    layer2_outputs(1576) <= not a;
    layer2_outputs(1577) <= not b or a;
    layer2_outputs(1578) <= a;
    layer2_outputs(1579) <= not a;
    layer2_outputs(1580) <= not b or a;
    layer2_outputs(1581) <= b and not a;
    layer2_outputs(1582) <= a;
    layer2_outputs(1583) <= not (a or b);
    layer2_outputs(1584) <= a;
    layer2_outputs(1585) <= a and b;
    layer2_outputs(1586) <= 1'b1;
    layer2_outputs(1587) <= b and not a;
    layer2_outputs(1588) <= not a;
    layer2_outputs(1589) <= not a;
    layer2_outputs(1590) <= a;
    layer2_outputs(1591) <= a and b;
    layer2_outputs(1592) <= not a or b;
    layer2_outputs(1593) <= a xor b;
    layer2_outputs(1594) <= not a;
    layer2_outputs(1595) <= a and b;
    layer2_outputs(1596) <= not b;
    layer2_outputs(1597) <= not b or a;
    layer2_outputs(1598) <= a xor b;
    layer2_outputs(1599) <= not a;
    layer2_outputs(1600) <= not (a and b);
    layer2_outputs(1601) <= not a or b;
    layer2_outputs(1602) <= b and not a;
    layer2_outputs(1603) <= a and b;
    layer2_outputs(1604) <= a or b;
    layer2_outputs(1605) <= a xor b;
    layer2_outputs(1606) <= a or b;
    layer2_outputs(1607) <= 1'b0;
    layer2_outputs(1608) <= b and not a;
    layer2_outputs(1609) <= b and not a;
    layer2_outputs(1610) <= not a or b;
    layer2_outputs(1611) <= a;
    layer2_outputs(1612) <= not b;
    layer2_outputs(1613) <= 1'b0;
    layer2_outputs(1614) <= b and not a;
    layer2_outputs(1615) <= a;
    layer2_outputs(1616) <= a or b;
    layer2_outputs(1617) <= a and not b;
    layer2_outputs(1618) <= a;
    layer2_outputs(1619) <= a and b;
    layer2_outputs(1620) <= a and not b;
    layer2_outputs(1621) <= not (a and b);
    layer2_outputs(1622) <= b and not a;
    layer2_outputs(1623) <= not (a xor b);
    layer2_outputs(1624) <= not a;
    layer2_outputs(1625) <= not a;
    layer2_outputs(1626) <= a;
    layer2_outputs(1627) <= not b or a;
    layer2_outputs(1628) <= a or b;
    layer2_outputs(1629) <= not b or a;
    layer2_outputs(1630) <= not a or b;
    layer2_outputs(1631) <= not b or a;
    layer2_outputs(1632) <= a and b;
    layer2_outputs(1633) <= not a;
    layer2_outputs(1634) <= not (a xor b);
    layer2_outputs(1635) <= not (a or b);
    layer2_outputs(1636) <= not b;
    layer2_outputs(1637) <= not b or a;
    layer2_outputs(1638) <= not b;
    layer2_outputs(1639) <= 1'b0;
    layer2_outputs(1640) <= a and b;
    layer2_outputs(1641) <= not b;
    layer2_outputs(1642) <= a;
    layer2_outputs(1643) <= a and not b;
    layer2_outputs(1644) <= b;
    layer2_outputs(1645) <= not b or a;
    layer2_outputs(1646) <= a;
    layer2_outputs(1647) <= not b;
    layer2_outputs(1648) <= not (a or b);
    layer2_outputs(1649) <= not (a or b);
    layer2_outputs(1650) <= not a or b;
    layer2_outputs(1651) <= not a or b;
    layer2_outputs(1652) <= not a;
    layer2_outputs(1653) <= b;
    layer2_outputs(1654) <= not a;
    layer2_outputs(1655) <= not b;
    layer2_outputs(1656) <= not a;
    layer2_outputs(1657) <= a and b;
    layer2_outputs(1658) <= a;
    layer2_outputs(1659) <= not (a and b);
    layer2_outputs(1660) <= not (a xor b);
    layer2_outputs(1661) <= a;
    layer2_outputs(1662) <= not (a or b);
    layer2_outputs(1663) <= b;
    layer2_outputs(1664) <= a;
    layer2_outputs(1665) <= b;
    layer2_outputs(1666) <= not (a or b);
    layer2_outputs(1667) <= a;
    layer2_outputs(1668) <= not (a and b);
    layer2_outputs(1669) <= not (a or b);
    layer2_outputs(1670) <= not (a or b);
    layer2_outputs(1671) <= a xor b;
    layer2_outputs(1672) <= not b or a;
    layer2_outputs(1673) <= not (a or b);
    layer2_outputs(1674) <= not b or a;
    layer2_outputs(1675) <= not a;
    layer2_outputs(1676) <= not (a xor b);
    layer2_outputs(1677) <= not a;
    layer2_outputs(1678) <= b;
    layer2_outputs(1679) <= a xor b;
    layer2_outputs(1680) <= a;
    layer2_outputs(1681) <= not (a and b);
    layer2_outputs(1682) <= b;
    layer2_outputs(1683) <= not (a or b);
    layer2_outputs(1684) <= a;
    layer2_outputs(1685) <= a;
    layer2_outputs(1686) <= 1'b0;
    layer2_outputs(1687) <= not a;
    layer2_outputs(1688) <= a and not b;
    layer2_outputs(1689) <= a;
    layer2_outputs(1690) <= a;
    layer2_outputs(1691) <= not a;
    layer2_outputs(1692) <= not b or a;
    layer2_outputs(1693) <= not a;
    layer2_outputs(1694) <= a;
    layer2_outputs(1695) <= b;
    layer2_outputs(1696) <= not b;
    layer2_outputs(1697) <= not a;
    layer2_outputs(1698) <= 1'b0;
    layer2_outputs(1699) <= not (a xor b);
    layer2_outputs(1700) <= not a;
    layer2_outputs(1701) <= b;
    layer2_outputs(1702) <= not (a and b);
    layer2_outputs(1703) <= a and b;
    layer2_outputs(1704) <= a and not b;
    layer2_outputs(1705) <= b;
    layer2_outputs(1706) <= not (a xor b);
    layer2_outputs(1707) <= not (a xor b);
    layer2_outputs(1708) <= not a;
    layer2_outputs(1709) <= a xor b;
    layer2_outputs(1710) <= a or b;
    layer2_outputs(1711) <= a and not b;
    layer2_outputs(1712) <= not b;
    layer2_outputs(1713) <= a xor b;
    layer2_outputs(1714) <= a;
    layer2_outputs(1715) <= a and b;
    layer2_outputs(1716) <= a and not b;
    layer2_outputs(1717) <= not a;
    layer2_outputs(1718) <= a and not b;
    layer2_outputs(1719) <= not a;
    layer2_outputs(1720) <= b;
    layer2_outputs(1721) <= a and not b;
    layer2_outputs(1722) <= not b;
    layer2_outputs(1723) <= 1'b1;
    layer2_outputs(1724) <= b and not a;
    layer2_outputs(1725) <= b and not a;
    layer2_outputs(1726) <= not a;
    layer2_outputs(1727) <= a or b;
    layer2_outputs(1728) <= a;
    layer2_outputs(1729) <= a and b;
    layer2_outputs(1730) <= not a;
    layer2_outputs(1731) <= a and not b;
    layer2_outputs(1732) <= a and not b;
    layer2_outputs(1733) <= b and not a;
    layer2_outputs(1734) <= a and b;
    layer2_outputs(1735) <= b and not a;
    layer2_outputs(1736) <= not a or b;
    layer2_outputs(1737) <= b and not a;
    layer2_outputs(1738) <= not a;
    layer2_outputs(1739) <= a or b;
    layer2_outputs(1740) <= not a;
    layer2_outputs(1741) <= a and not b;
    layer2_outputs(1742) <= not b or a;
    layer2_outputs(1743) <= not a;
    layer2_outputs(1744) <= not b;
    layer2_outputs(1745) <= not (a xor b);
    layer2_outputs(1746) <= a;
    layer2_outputs(1747) <= a;
    layer2_outputs(1748) <= not b or a;
    layer2_outputs(1749) <= not (a or b);
    layer2_outputs(1750) <= not a;
    layer2_outputs(1751) <= not a or b;
    layer2_outputs(1752) <= not b;
    layer2_outputs(1753) <= b;
    layer2_outputs(1754) <= a;
    layer2_outputs(1755) <= a xor b;
    layer2_outputs(1756) <= b;
    layer2_outputs(1757) <= not a or b;
    layer2_outputs(1758) <= not b;
    layer2_outputs(1759) <= not a or b;
    layer2_outputs(1760) <= not (a and b);
    layer2_outputs(1761) <= b;
    layer2_outputs(1762) <= not b;
    layer2_outputs(1763) <= not (a xor b);
    layer2_outputs(1764) <= not b or a;
    layer2_outputs(1765) <= not b;
    layer2_outputs(1766) <= not a;
    layer2_outputs(1767) <= a and b;
    layer2_outputs(1768) <= not a or b;
    layer2_outputs(1769) <= not a;
    layer2_outputs(1770) <= 1'b1;
    layer2_outputs(1771) <= not (a or b);
    layer2_outputs(1772) <= a xor b;
    layer2_outputs(1773) <= 1'b1;
    layer2_outputs(1774) <= not (a or b);
    layer2_outputs(1775) <= not b;
    layer2_outputs(1776) <= not a;
    layer2_outputs(1777) <= b;
    layer2_outputs(1778) <= a and not b;
    layer2_outputs(1779) <= a or b;
    layer2_outputs(1780) <= b;
    layer2_outputs(1781) <= not a or b;
    layer2_outputs(1782) <= not b or a;
    layer2_outputs(1783) <= not (a or b);
    layer2_outputs(1784) <= a;
    layer2_outputs(1785) <= b and not a;
    layer2_outputs(1786) <= a and b;
    layer2_outputs(1787) <= not a or b;
    layer2_outputs(1788) <= not b or a;
    layer2_outputs(1789) <= not (a xor b);
    layer2_outputs(1790) <= not b;
    layer2_outputs(1791) <= not (a and b);
    layer2_outputs(1792) <= a;
    layer2_outputs(1793) <= b;
    layer2_outputs(1794) <= a;
    layer2_outputs(1795) <= not b;
    layer2_outputs(1796) <= not (a xor b);
    layer2_outputs(1797) <= not b;
    layer2_outputs(1798) <= a or b;
    layer2_outputs(1799) <= not a;
    layer2_outputs(1800) <= not (a and b);
    layer2_outputs(1801) <= a xor b;
    layer2_outputs(1802) <= not (a and b);
    layer2_outputs(1803) <= a xor b;
    layer2_outputs(1804) <= a;
    layer2_outputs(1805) <= not (a xor b);
    layer2_outputs(1806) <= not b;
    layer2_outputs(1807) <= not (a xor b);
    layer2_outputs(1808) <= a;
    layer2_outputs(1809) <= a or b;
    layer2_outputs(1810) <= not a or b;
    layer2_outputs(1811) <= not b;
    layer2_outputs(1812) <= a;
    layer2_outputs(1813) <= not b;
    layer2_outputs(1814) <= not a;
    layer2_outputs(1815) <= not (a xor b);
    layer2_outputs(1816) <= not a;
    layer2_outputs(1817) <= a and b;
    layer2_outputs(1818) <= b;
    layer2_outputs(1819) <= b;
    layer2_outputs(1820) <= not (a and b);
    layer2_outputs(1821) <= not a or b;
    layer2_outputs(1822) <= not (a and b);
    layer2_outputs(1823) <= a xor b;
    layer2_outputs(1824) <= b;
    layer2_outputs(1825) <= not a or b;
    layer2_outputs(1826) <= a and not b;
    layer2_outputs(1827) <= not (a or b);
    layer2_outputs(1828) <= b;
    layer2_outputs(1829) <= b and not a;
    layer2_outputs(1830) <= not (a and b);
    layer2_outputs(1831) <= not a;
    layer2_outputs(1832) <= not (a and b);
    layer2_outputs(1833) <= a and b;
    layer2_outputs(1834) <= not a;
    layer2_outputs(1835) <= not (a xor b);
    layer2_outputs(1836) <= not b or a;
    layer2_outputs(1837) <= a xor b;
    layer2_outputs(1838) <= not b or a;
    layer2_outputs(1839) <= a;
    layer2_outputs(1840) <= a and b;
    layer2_outputs(1841) <= a and not b;
    layer2_outputs(1842) <= 1'b1;
    layer2_outputs(1843) <= not (a and b);
    layer2_outputs(1844) <= not a;
    layer2_outputs(1845) <= 1'b1;
    layer2_outputs(1846) <= not b;
    layer2_outputs(1847) <= 1'b1;
    layer2_outputs(1848) <= not b;
    layer2_outputs(1849) <= not b;
    layer2_outputs(1850) <= a;
    layer2_outputs(1851) <= a and b;
    layer2_outputs(1852) <= not (a xor b);
    layer2_outputs(1853) <= not a;
    layer2_outputs(1854) <= not b;
    layer2_outputs(1855) <= a or b;
    layer2_outputs(1856) <= not a;
    layer2_outputs(1857) <= not (a and b);
    layer2_outputs(1858) <= not b or a;
    layer2_outputs(1859) <= b;
    layer2_outputs(1860) <= not (a and b);
    layer2_outputs(1861) <= a and not b;
    layer2_outputs(1862) <= b;
    layer2_outputs(1863) <= not a;
    layer2_outputs(1864) <= not a or b;
    layer2_outputs(1865) <= not b;
    layer2_outputs(1866) <= a and not b;
    layer2_outputs(1867) <= not a or b;
    layer2_outputs(1868) <= a and not b;
    layer2_outputs(1869) <= not (a or b);
    layer2_outputs(1870) <= not b;
    layer2_outputs(1871) <= 1'b0;
    layer2_outputs(1872) <= a or b;
    layer2_outputs(1873) <= not (a or b);
    layer2_outputs(1874) <= not b or a;
    layer2_outputs(1875) <= not b or a;
    layer2_outputs(1876) <= not b or a;
    layer2_outputs(1877) <= not a;
    layer2_outputs(1878) <= a or b;
    layer2_outputs(1879) <= b;
    layer2_outputs(1880) <= a;
    layer2_outputs(1881) <= b;
    layer2_outputs(1882) <= not b;
    layer2_outputs(1883) <= not b or a;
    layer2_outputs(1884) <= a and b;
    layer2_outputs(1885) <= not b;
    layer2_outputs(1886) <= not (a and b);
    layer2_outputs(1887) <= not b;
    layer2_outputs(1888) <= not a;
    layer2_outputs(1889) <= not (a xor b);
    layer2_outputs(1890) <= not a or b;
    layer2_outputs(1891) <= a and b;
    layer2_outputs(1892) <= not (a xor b);
    layer2_outputs(1893) <= not a;
    layer2_outputs(1894) <= a and not b;
    layer2_outputs(1895) <= a and not b;
    layer2_outputs(1896) <= not (a and b);
    layer2_outputs(1897) <= not (a xor b);
    layer2_outputs(1898) <= not b;
    layer2_outputs(1899) <= 1'b0;
    layer2_outputs(1900) <= not b;
    layer2_outputs(1901) <= not b or a;
    layer2_outputs(1902) <= not b or a;
    layer2_outputs(1903) <= a and not b;
    layer2_outputs(1904) <= a and not b;
    layer2_outputs(1905) <= a and b;
    layer2_outputs(1906) <= not a;
    layer2_outputs(1907) <= not (a or b);
    layer2_outputs(1908) <= not b or a;
    layer2_outputs(1909) <= not b;
    layer2_outputs(1910) <= a or b;
    layer2_outputs(1911) <= not b;
    layer2_outputs(1912) <= not a or b;
    layer2_outputs(1913) <= a and not b;
    layer2_outputs(1914) <= a and not b;
    layer2_outputs(1915) <= a;
    layer2_outputs(1916) <= not a;
    layer2_outputs(1917) <= a and not b;
    layer2_outputs(1918) <= not a;
    layer2_outputs(1919) <= not a or b;
    layer2_outputs(1920) <= b;
    layer2_outputs(1921) <= a;
    layer2_outputs(1922) <= not a;
    layer2_outputs(1923) <= a and b;
    layer2_outputs(1924) <= a;
    layer2_outputs(1925) <= b;
    layer2_outputs(1926) <= not (a and b);
    layer2_outputs(1927) <= not a;
    layer2_outputs(1928) <= not a or b;
    layer2_outputs(1929) <= not a;
    layer2_outputs(1930) <= a and not b;
    layer2_outputs(1931) <= not a;
    layer2_outputs(1932) <= not (a and b);
    layer2_outputs(1933) <= not a or b;
    layer2_outputs(1934) <= a;
    layer2_outputs(1935) <= a or b;
    layer2_outputs(1936) <= a or b;
    layer2_outputs(1937) <= not a or b;
    layer2_outputs(1938) <= not a;
    layer2_outputs(1939) <= a;
    layer2_outputs(1940) <= not b;
    layer2_outputs(1941) <= not a;
    layer2_outputs(1942) <= not b;
    layer2_outputs(1943) <= a and not b;
    layer2_outputs(1944) <= not (a or b);
    layer2_outputs(1945) <= b;
    layer2_outputs(1946) <= a or b;
    layer2_outputs(1947) <= a or b;
    layer2_outputs(1948) <= not b;
    layer2_outputs(1949) <= b and not a;
    layer2_outputs(1950) <= a xor b;
    layer2_outputs(1951) <= 1'b0;
    layer2_outputs(1952) <= not b;
    layer2_outputs(1953) <= not b or a;
    layer2_outputs(1954) <= not b;
    layer2_outputs(1955) <= a;
    layer2_outputs(1956) <= b;
    layer2_outputs(1957) <= not a or b;
    layer2_outputs(1958) <= not a;
    layer2_outputs(1959) <= a;
    layer2_outputs(1960) <= not b;
    layer2_outputs(1961) <= a and not b;
    layer2_outputs(1962) <= b and not a;
    layer2_outputs(1963) <= not b or a;
    layer2_outputs(1964) <= not a or b;
    layer2_outputs(1965) <= not (a or b);
    layer2_outputs(1966) <= not b or a;
    layer2_outputs(1967) <= a and b;
    layer2_outputs(1968) <= b and not a;
    layer2_outputs(1969) <= a xor b;
    layer2_outputs(1970) <= a or b;
    layer2_outputs(1971) <= 1'b0;
    layer2_outputs(1972) <= not b;
    layer2_outputs(1973) <= a and b;
    layer2_outputs(1974) <= not b or a;
    layer2_outputs(1975) <= not (a and b);
    layer2_outputs(1976) <= not a;
    layer2_outputs(1977) <= a or b;
    layer2_outputs(1978) <= a;
    layer2_outputs(1979) <= not (a xor b);
    layer2_outputs(1980) <= a;
    layer2_outputs(1981) <= b;
    layer2_outputs(1982) <= not b or a;
    layer2_outputs(1983) <= not (a or b);
    layer2_outputs(1984) <= b;
    layer2_outputs(1985) <= not b;
    layer2_outputs(1986) <= not b;
    layer2_outputs(1987) <= a xor b;
    layer2_outputs(1988) <= not b;
    layer2_outputs(1989) <= not a;
    layer2_outputs(1990) <= not (a xor b);
    layer2_outputs(1991) <= not (a xor b);
    layer2_outputs(1992) <= not (a or b);
    layer2_outputs(1993) <= a;
    layer2_outputs(1994) <= not (a or b);
    layer2_outputs(1995) <= not (a or b);
    layer2_outputs(1996) <= a and not b;
    layer2_outputs(1997) <= b;
    layer2_outputs(1998) <= not b;
    layer2_outputs(1999) <= b and not a;
    layer2_outputs(2000) <= not (a and b);
    layer2_outputs(2001) <= not a;
    layer2_outputs(2002) <= not (a and b);
    layer2_outputs(2003) <= b and not a;
    layer2_outputs(2004) <= not (a or b);
    layer2_outputs(2005) <= a or b;
    layer2_outputs(2006) <= not a or b;
    layer2_outputs(2007) <= not b;
    layer2_outputs(2008) <= not b;
    layer2_outputs(2009) <= b and not a;
    layer2_outputs(2010) <= a;
    layer2_outputs(2011) <= not b;
    layer2_outputs(2012) <= not b;
    layer2_outputs(2013) <= a;
    layer2_outputs(2014) <= not a;
    layer2_outputs(2015) <= a;
    layer2_outputs(2016) <= not a;
    layer2_outputs(2017) <= a and b;
    layer2_outputs(2018) <= a or b;
    layer2_outputs(2019) <= not (a and b);
    layer2_outputs(2020) <= a xor b;
    layer2_outputs(2021) <= a and b;
    layer2_outputs(2022) <= not (a xor b);
    layer2_outputs(2023) <= not b;
    layer2_outputs(2024) <= a or b;
    layer2_outputs(2025) <= not a;
    layer2_outputs(2026) <= b;
    layer2_outputs(2027) <= not (a or b);
    layer2_outputs(2028) <= a and not b;
    layer2_outputs(2029) <= not a;
    layer2_outputs(2030) <= not (a and b);
    layer2_outputs(2031) <= not (a or b);
    layer2_outputs(2032) <= not b or a;
    layer2_outputs(2033) <= 1'b1;
    layer2_outputs(2034) <= a;
    layer2_outputs(2035) <= a;
    layer2_outputs(2036) <= not (a and b);
    layer2_outputs(2037) <= a;
    layer2_outputs(2038) <= a;
    layer2_outputs(2039) <= b;
    layer2_outputs(2040) <= a or b;
    layer2_outputs(2041) <= not a or b;
    layer2_outputs(2042) <= not (a and b);
    layer2_outputs(2043) <= not a;
    layer2_outputs(2044) <= b;
    layer2_outputs(2045) <= b;
    layer2_outputs(2046) <= b;
    layer2_outputs(2047) <= b and not a;
    layer2_outputs(2048) <= not (a xor b);
    layer2_outputs(2049) <= not a;
    layer2_outputs(2050) <= a and not b;
    layer2_outputs(2051) <= a and not b;
    layer2_outputs(2052) <= not a;
    layer2_outputs(2053) <= b;
    layer2_outputs(2054) <= not (a or b);
    layer2_outputs(2055) <= a or b;
    layer2_outputs(2056) <= not a;
    layer2_outputs(2057) <= a and b;
    layer2_outputs(2058) <= not (a and b);
    layer2_outputs(2059) <= a or b;
    layer2_outputs(2060) <= a and b;
    layer2_outputs(2061) <= not a;
    layer2_outputs(2062) <= a;
    layer2_outputs(2063) <= b;
    layer2_outputs(2064) <= b;
    layer2_outputs(2065) <= not b or a;
    layer2_outputs(2066) <= 1'b0;
    layer2_outputs(2067) <= not b or a;
    layer2_outputs(2068) <= b;
    layer2_outputs(2069) <= a;
    layer2_outputs(2070) <= a xor b;
    layer2_outputs(2071) <= b;
    layer2_outputs(2072) <= not b or a;
    layer2_outputs(2073) <= not b or a;
    layer2_outputs(2074) <= not a or b;
    layer2_outputs(2075) <= not b;
    layer2_outputs(2076) <= not a;
    layer2_outputs(2077) <= not b or a;
    layer2_outputs(2078) <= a;
    layer2_outputs(2079) <= not b;
    layer2_outputs(2080) <= a or b;
    layer2_outputs(2081) <= not (a or b);
    layer2_outputs(2082) <= not a;
    layer2_outputs(2083) <= not a;
    layer2_outputs(2084) <= b;
    layer2_outputs(2085) <= a and not b;
    layer2_outputs(2086) <= not b or a;
    layer2_outputs(2087) <= not a or b;
    layer2_outputs(2088) <= not a;
    layer2_outputs(2089) <= not (a or b);
    layer2_outputs(2090) <= not a;
    layer2_outputs(2091) <= a;
    layer2_outputs(2092) <= not b;
    layer2_outputs(2093) <= not (a and b);
    layer2_outputs(2094) <= not a;
    layer2_outputs(2095) <= a;
    layer2_outputs(2096) <= not a or b;
    layer2_outputs(2097) <= a;
    layer2_outputs(2098) <= not (a and b);
    layer2_outputs(2099) <= a and b;
    layer2_outputs(2100) <= not (a xor b);
    layer2_outputs(2101) <= not a or b;
    layer2_outputs(2102) <= not a;
    layer2_outputs(2103) <= b;
    layer2_outputs(2104) <= a and not b;
    layer2_outputs(2105) <= a xor b;
    layer2_outputs(2106) <= b and not a;
    layer2_outputs(2107) <= not a;
    layer2_outputs(2108) <= not b or a;
    layer2_outputs(2109) <= not (a and b);
    layer2_outputs(2110) <= not a or b;
    layer2_outputs(2111) <= not a;
    layer2_outputs(2112) <= a and not b;
    layer2_outputs(2113) <= a xor b;
    layer2_outputs(2114) <= not b or a;
    layer2_outputs(2115) <= a;
    layer2_outputs(2116) <= a and not b;
    layer2_outputs(2117) <= not b or a;
    layer2_outputs(2118) <= a or b;
    layer2_outputs(2119) <= a and b;
    layer2_outputs(2120) <= not a or b;
    layer2_outputs(2121) <= not a or b;
    layer2_outputs(2122) <= not a;
    layer2_outputs(2123) <= b;
    layer2_outputs(2124) <= a and b;
    layer2_outputs(2125) <= a or b;
    layer2_outputs(2126) <= not b or a;
    layer2_outputs(2127) <= a;
    layer2_outputs(2128) <= a;
    layer2_outputs(2129) <= b and not a;
    layer2_outputs(2130) <= not (a xor b);
    layer2_outputs(2131) <= a and not b;
    layer2_outputs(2132) <= b and not a;
    layer2_outputs(2133) <= a or b;
    layer2_outputs(2134) <= a;
    layer2_outputs(2135) <= a or b;
    layer2_outputs(2136) <= b;
    layer2_outputs(2137) <= not (a xor b);
    layer2_outputs(2138) <= not b;
    layer2_outputs(2139) <= not b;
    layer2_outputs(2140) <= not (a and b);
    layer2_outputs(2141) <= not a or b;
    layer2_outputs(2142) <= a and not b;
    layer2_outputs(2143) <= 1'b1;
    layer2_outputs(2144) <= not b;
    layer2_outputs(2145) <= not a;
    layer2_outputs(2146) <= not (a or b);
    layer2_outputs(2147) <= not (a or b);
    layer2_outputs(2148) <= not (a and b);
    layer2_outputs(2149) <= not (a xor b);
    layer2_outputs(2150) <= not b or a;
    layer2_outputs(2151) <= not (a or b);
    layer2_outputs(2152) <= b;
    layer2_outputs(2153) <= a xor b;
    layer2_outputs(2154) <= a;
    layer2_outputs(2155) <= not (a xor b);
    layer2_outputs(2156) <= b;
    layer2_outputs(2157) <= a or b;
    layer2_outputs(2158) <= a or b;
    layer2_outputs(2159) <= a;
    layer2_outputs(2160) <= not b;
    layer2_outputs(2161) <= a and not b;
    layer2_outputs(2162) <= not a;
    layer2_outputs(2163) <= 1'b1;
    layer2_outputs(2164) <= a or b;
    layer2_outputs(2165) <= not b;
    layer2_outputs(2166) <= 1'b0;
    layer2_outputs(2167) <= b and not a;
    layer2_outputs(2168) <= b and not a;
    layer2_outputs(2169) <= a and not b;
    layer2_outputs(2170) <= not b;
    layer2_outputs(2171) <= not b;
    layer2_outputs(2172) <= a;
    layer2_outputs(2173) <= a;
    layer2_outputs(2174) <= b;
    layer2_outputs(2175) <= not b;
    layer2_outputs(2176) <= not (a or b);
    layer2_outputs(2177) <= not a;
    layer2_outputs(2178) <= a and b;
    layer2_outputs(2179) <= not b;
    layer2_outputs(2180) <= a or b;
    layer2_outputs(2181) <= a xor b;
    layer2_outputs(2182) <= a;
    layer2_outputs(2183) <= not b;
    layer2_outputs(2184) <= not b;
    layer2_outputs(2185) <= not a;
    layer2_outputs(2186) <= a and b;
    layer2_outputs(2187) <= not a;
    layer2_outputs(2188) <= not a;
    layer2_outputs(2189) <= a or b;
    layer2_outputs(2190) <= not b;
    layer2_outputs(2191) <= a;
    layer2_outputs(2192) <= not a or b;
    layer2_outputs(2193) <= a and not b;
    layer2_outputs(2194) <= b;
    layer2_outputs(2195) <= 1'b0;
    layer2_outputs(2196) <= b and not a;
    layer2_outputs(2197) <= not a or b;
    layer2_outputs(2198) <= not b;
    layer2_outputs(2199) <= not a or b;
    layer2_outputs(2200) <= a and b;
    layer2_outputs(2201) <= a or b;
    layer2_outputs(2202) <= not a or b;
    layer2_outputs(2203) <= b;
    layer2_outputs(2204) <= 1'b0;
    layer2_outputs(2205) <= a;
    layer2_outputs(2206) <= a xor b;
    layer2_outputs(2207) <= a and not b;
    layer2_outputs(2208) <= a xor b;
    layer2_outputs(2209) <= a and not b;
    layer2_outputs(2210) <= b and not a;
    layer2_outputs(2211) <= a;
    layer2_outputs(2212) <= not a;
    layer2_outputs(2213) <= not b;
    layer2_outputs(2214) <= b;
    layer2_outputs(2215) <= not b or a;
    layer2_outputs(2216) <= a or b;
    layer2_outputs(2217) <= a and not b;
    layer2_outputs(2218) <= 1'b1;
    layer2_outputs(2219) <= not b;
    layer2_outputs(2220) <= not b;
    layer2_outputs(2221) <= not (a and b);
    layer2_outputs(2222) <= a;
    layer2_outputs(2223) <= not (a xor b);
    layer2_outputs(2224) <= a or b;
    layer2_outputs(2225) <= b;
    layer2_outputs(2226) <= not (a or b);
    layer2_outputs(2227) <= b and not a;
    layer2_outputs(2228) <= not a;
    layer2_outputs(2229) <= not (a or b);
    layer2_outputs(2230) <= not a;
    layer2_outputs(2231) <= not (a or b);
    layer2_outputs(2232) <= b;
    layer2_outputs(2233) <= a;
    layer2_outputs(2234) <= not b;
    layer2_outputs(2235) <= a and b;
    layer2_outputs(2236) <= a;
    layer2_outputs(2237) <= not (a and b);
    layer2_outputs(2238) <= a and not b;
    layer2_outputs(2239) <= not b;
    layer2_outputs(2240) <= not a;
    layer2_outputs(2241) <= not a;
    layer2_outputs(2242) <= a xor b;
    layer2_outputs(2243) <= a;
    layer2_outputs(2244) <= not a;
    layer2_outputs(2245) <= not (a or b);
    layer2_outputs(2246) <= b and not a;
    layer2_outputs(2247) <= a or b;
    layer2_outputs(2248) <= not (a or b);
    layer2_outputs(2249) <= a and b;
    layer2_outputs(2250) <= a or b;
    layer2_outputs(2251) <= not a or b;
    layer2_outputs(2252) <= not (a or b);
    layer2_outputs(2253) <= a and b;
    layer2_outputs(2254) <= not a or b;
    layer2_outputs(2255) <= b;
    layer2_outputs(2256) <= not a or b;
    layer2_outputs(2257) <= not b;
    layer2_outputs(2258) <= not b or a;
    layer2_outputs(2259) <= a;
    layer2_outputs(2260) <= not b or a;
    layer2_outputs(2261) <= not b;
    layer2_outputs(2262) <= a;
    layer2_outputs(2263) <= not (a and b);
    layer2_outputs(2264) <= not a or b;
    layer2_outputs(2265) <= not (a or b);
    layer2_outputs(2266) <= not a or b;
    layer2_outputs(2267) <= not b or a;
    layer2_outputs(2268) <= b;
    layer2_outputs(2269) <= not b;
    layer2_outputs(2270) <= not (a or b);
    layer2_outputs(2271) <= 1'b0;
    layer2_outputs(2272) <= 1'b1;
    layer2_outputs(2273) <= a and b;
    layer2_outputs(2274) <= not (a or b);
    layer2_outputs(2275) <= not b;
    layer2_outputs(2276) <= not b;
    layer2_outputs(2277) <= not a or b;
    layer2_outputs(2278) <= a and b;
    layer2_outputs(2279) <= b and not a;
    layer2_outputs(2280) <= b;
    layer2_outputs(2281) <= a or b;
    layer2_outputs(2282) <= b and not a;
    layer2_outputs(2283) <= a and not b;
    layer2_outputs(2284) <= not b;
    layer2_outputs(2285) <= not (a or b);
    layer2_outputs(2286) <= a and b;
    layer2_outputs(2287) <= b and not a;
    layer2_outputs(2288) <= not (a and b);
    layer2_outputs(2289) <= a or b;
    layer2_outputs(2290) <= not b or a;
    layer2_outputs(2291) <= not (a and b);
    layer2_outputs(2292) <= not a;
    layer2_outputs(2293) <= not a;
    layer2_outputs(2294) <= not b or a;
    layer2_outputs(2295) <= not b or a;
    layer2_outputs(2296) <= not (a and b);
    layer2_outputs(2297) <= not b;
    layer2_outputs(2298) <= not (a and b);
    layer2_outputs(2299) <= not a;
    layer2_outputs(2300) <= a xor b;
    layer2_outputs(2301) <= a xor b;
    layer2_outputs(2302) <= b;
    layer2_outputs(2303) <= not a;
    layer2_outputs(2304) <= not a or b;
    layer2_outputs(2305) <= not a or b;
    layer2_outputs(2306) <= a and not b;
    layer2_outputs(2307) <= not b;
    layer2_outputs(2308) <= not a;
    layer2_outputs(2309) <= b;
    layer2_outputs(2310) <= not (a and b);
    layer2_outputs(2311) <= not b;
    layer2_outputs(2312) <= a;
    layer2_outputs(2313) <= a and not b;
    layer2_outputs(2314) <= not a or b;
    layer2_outputs(2315) <= a;
    layer2_outputs(2316) <= not b;
    layer2_outputs(2317) <= a;
    layer2_outputs(2318) <= not (a and b);
    layer2_outputs(2319) <= a;
    layer2_outputs(2320) <= not (a and b);
    layer2_outputs(2321) <= not (a xor b);
    layer2_outputs(2322) <= b and not a;
    layer2_outputs(2323) <= a or b;
    layer2_outputs(2324) <= not (a and b);
    layer2_outputs(2325) <= not (a and b);
    layer2_outputs(2326) <= a and not b;
    layer2_outputs(2327) <= not a;
    layer2_outputs(2328) <= 1'b1;
    layer2_outputs(2329) <= not a;
    layer2_outputs(2330) <= not b or a;
    layer2_outputs(2331) <= not b;
    layer2_outputs(2332) <= not b;
    layer2_outputs(2333) <= a and not b;
    layer2_outputs(2334) <= not (a xor b);
    layer2_outputs(2335) <= not (a or b);
    layer2_outputs(2336) <= not a;
    layer2_outputs(2337) <= not (a or b);
    layer2_outputs(2338) <= not a;
    layer2_outputs(2339) <= not (a or b);
    layer2_outputs(2340) <= b;
    layer2_outputs(2341) <= b and not a;
    layer2_outputs(2342) <= a and not b;
    layer2_outputs(2343) <= not b;
    layer2_outputs(2344) <= not (a or b);
    layer2_outputs(2345) <= not b;
    layer2_outputs(2346) <= not b;
    layer2_outputs(2347) <= a;
    layer2_outputs(2348) <= a;
    layer2_outputs(2349) <= not b or a;
    layer2_outputs(2350) <= not a;
    layer2_outputs(2351) <= not b;
    layer2_outputs(2352) <= b and not a;
    layer2_outputs(2353) <= not (a and b);
    layer2_outputs(2354) <= not a;
    layer2_outputs(2355) <= b;
    layer2_outputs(2356) <= not (a and b);
    layer2_outputs(2357) <= a and not b;
    layer2_outputs(2358) <= not (a xor b);
    layer2_outputs(2359) <= not a or b;
    layer2_outputs(2360) <= 1'b1;
    layer2_outputs(2361) <= not b;
    layer2_outputs(2362) <= not a;
    layer2_outputs(2363) <= a or b;
    layer2_outputs(2364) <= not (a or b);
    layer2_outputs(2365) <= b;
    layer2_outputs(2366) <= a xor b;
    layer2_outputs(2367) <= a;
    layer2_outputs(2368) <= not (a xor b);
    layer2_outputs(2369) <= a and b;
    layer2_outputs(2370) <= not a;
    layer2_outputs(2371) <= 1'b1;
    layer2_outputs(2372) <= a and not b;
    layer2_outputs(2373) <= a;
    layer2_outputs(2374) <= a;
    layer2_outputs(2375) <= a and b;
    layer2_outputs(2376) <= b;
    layer2_outputs(2377) <= a;
    layer2_outputs(2378) <= a and not b;
    layer2_outputs(2379) <= not (a and b);
    layer2_outputs(2380) <= b;
    layer2_outputs(2381) <= not a or b;
    layer2_outputs(2382) <= a or b;
    layer2_outputs(2383) <= not b or a;
    layer2_outputs(2384) <= a and not b;
    layer2_outputs(2385) <= not (a and b);
    layer2_outputs(2386) <= not b or a;
    layer2_outputs(2387) <= a and not b;
    layer2_outputs(2388) <= a or b;
    layer2_outputs(2389) <= 1'b1;
    layer2_outputs(2390) <= b;
    layer2_outputs(2391) <= 1'b0;
    layer2_outputs(2392) <= b;
    layer2_outputs(2393) <= a;
    layer2_outputs(2394) <= a xor b;
    layer2_outputs(2395) <= not b or a;
    layer2_outputs(2396) <= b;
    layer2_outputs(2397) <= a and b;
    layer2_outputs(2398) <= not (a or b);
    layer2_outputs(2399) <= not a;
    layer2_outputs(2400) <= not a;
    layer2_outputs(2401) <= a and b;
    layer2_outputs(2402) <= not a;
    layer2_outputs(2403) <= 1'b1;
    layer2_outputs(2404) <= not a;
    layer2_outputs(2405) <= b;
    layer2_outputs(2406) <= 1'b0;
    layer2_outputs(2407) <= a;
    layer2_outputs(2408) <= 1'b0;
    layer2_outputs(2409) <= b;
    layer2_outputs(2410) <= a xor b;
    layer2_outputs(2411) <= a xor b;
    layer2_outputs(2412) <= 1'b0;
    layer2_outputs(2413) <= not (a and b);
    layer2_outputs(2414) <= not a;
    layer2_outputs(2415) <= not b;
    layer2_outputs(2416) <= not (a or b);
    layer2_outputs(2417) <= a;
    layer2_outputs(2418) <= a;
    layer2_outputs(2419) <= not (a or b);
    layer2_outputs(2420) <= not (a or b);
    layer2_outputs(2421) <= a xor b;
    layer2_outputs(2422) <= not a or b;
    layer2_outputs(2423) <= not b or a;
    layer2_outputs(2424) <= not a;
    layer2_outputs(2425) <= b;
    layer2_outputs(2426) <= not a or b;
    layer2_outputs(2427) <= b;
    layer2_outputs(2428) <= not (a or b);
    layer2_outputs(2429) <= a xor b;
    layer2_outputs(2430) <= a;
    layer2_outputs(2431) <= not a;
    layer2_outputs(2432) <= 1'b1;
    layer2_outputs(2433) <= a;
    layer2_outputs(2434) <= a;
    layer2_outputs(2435) <= 1'b1;
    layer2_outputs(2436) <= not (a or b);
    layer2_outputs(2437) <= not (a or b);
    layer2_outputs(2438) <= not a;
    layer2_outputs(2439) <= b;
    layer2_outputs(2440) <= b and not a;
    layer2_outputs(2441) <= a;
    layer2_outputs(2442) <= b and not a;
    layer2_outputs(2443) <= not a;
    layer2_outputs(2444) <= b;
    layer2_outputs(2445) <= not a;
    layer2_outputs(2446) <= a and b;
    layer2_outputs(2447) <= a;
    layer2_outputs(2448) <= b and not a;
    layer2_outputs(2449) <= a xor b;
    layer2_outputs(2450) <= not a or b;
    layer2_outputs(2451) <= b;
    layer2_outputs(2452) <= a;
    layer2_outputs(2453) <= b;
    layer2_outputs(2454) <= a;
    layer2_outputs(2455) <= a and b;
    layer2_outputs(2456) <= not (a or b);
    layer2_outputs(2457) <= b and not a;
    layer2_outputs(2458) <= a;
    layer2_outputs(2459) <= not (a xor b);
    layer2_outputs(2460) <= not (a or b);
    layer2_outputs(2461) <= a and b;
    layer2_outputs(2462) <= a or b;
    layer2_outputs(2463) <= not a;
    layer2_outputs(2464) <= not (a and b);
    layer2_outputs(2465) <= not (a xor b);
    layer2_outputs(2466) <= not a or b;
    layer2_outputs(2467) <= not (a xor b);
    layer2_outputs(2468) <= a xor b;
    layer2_outputs(2469) <= a xor b;
    layer2_outputs(2470) <= not a;
    layer2_outputs(2471) <= a and not b;
    layer2_outputs(2472) <= a or b;
    layer2_outputs(2473) <= b;
    layer2_outputs(2474) <= a and b;
    layer2_outputs(2475) <= 1'b1;
    layer2_outputs(2476) <= 1'b0;
    layer2_outputs(2477) <= not a;
    layer2_outputs(2478) <= not a;
    layer2_outputs(2479) <= a and not b;
    layer2_outputs(2480) <= b and not a;
    layer2_outputs(2481) <= not a or b;
    layer2_outputs(2482) <= a xor b;
    layer2_outputs(2483) <= b;
    layer2_outputs(2484) <= b and not a;
    layer2_outputs(2485) <= b;
    layer2_outputs(2486) <= not (a xor b);
    layer2_outputs(2487) <= not a or b;
    layer2_outputs(2488) <= a xor b;
    layer2_outputs(2489) <= a xor b;
    layer2_outputs(2490) <= a and not b;
    layer2_outputs(2491) <= a xor b;
    layer2_outputs(2492) <= not b or a;
    layer2_outputs(2493) <= a and not b;
    layer2_outputs(2494) <= a and b;
    layer2_outputs(2495) <= not b or a;
    layer2_outputs(2496) <= not a;
    layer2_outputs(2497) <= not b or a;
    layer2_outputs(2498) <= a;
    layer2_outputs(2499) <= not b;
    layer2_outputs(2500) <= a xor b;
    layer2_outputs(2501) <= b and not a;
    layer2_outputs(2502) <= a;
    layer2_outputs(2503) <= a;
    layer2_outputs(2504) <= not a or b;
    layer2_outputs(2505) <= not a or b;
    layer2_outputs(2506) <= a and not b;
    layer2_outputs(2507) <= b and not a;
    layer2_outputs(2508) <= not a;
    layer2_outputs(2509) <= a and not b;
    layer2_outputs(2510) <= not (a or b);
    layer2_outputs(2511) <= not b;
    layer2_outputs(2512) <= not a;
    layer2_outputs(2513) <= b;
    layer2_outputs(2514) <= not b;
    layer2_outputs(2515) <= not a or b;
    layer2_outputs(2516) <= not (a or b);
    layer2_outputs(2517) <= not b or a;
    layer2_outputs(2518) <= 1'b0;
    layer2_outputs(2519) <= not a or b;
    layer2_outputs(2520) <= b and not a;
    layer2_outputs(2521) <= a and not b;
    layer2_outputs(2522) <= a;
    layer2_outputs(2523) <= a or b;
    layer2_outputs(2524) <= not (a and b);
    layer2_outputs(2525) <= not b;
    layer2_outputs(2526) <= not a;
    layer2_outputs(2527) <= not a or b;
    layer2_outputs(2528) <= not (a and b);
    layer2_outputs(2529) <= a and b;
    layer2_outputs(2530) <= a;
    layer2_outputs(2531) <= 1'b0;
    layer2_outputs(2532) <= a and b;
    layer2_outputs(2533) <= b;
    layer2_outputs(2534) <= a or b;
    layer2_outputs(2535) <= a;
    layer2_outputs(2536) <= not a;
    layer2_outputs(2537) <= a;
    layer2_outputs(2538) <= not (a and b);
    layer2_outputs(2539) <= not (a or b);
    layer2_outputs(2540) <= b and not a;
    layer2_outputs(2541) <= a or b;
    layer2_outputs(2542) <= a xor b;
    layer2_outputs(2543) <= b and not a;
    layer2_outputs(2544) <= not a or b;
    layer2_outputs(2545) <= not (a or b);
    layer2_outputs(2546) <= b;
    layer2_outputs(2547) <= b and not a;
    layer2_outputs(2548) <= a and b;
    layer2_outputs(2549) <= a and not b;
    layer2_outputs(2550) <= a and b;
    layer2_outputs(2551) <= a;
    layer2_outputs(2552) <= a;
    layer2_outputs(2553) <= not a or b;
    layer2_outputs(2554) <= a and b;
    layer2_outputs(2555) <= not b or a;
    layer2_outputs(2556) <= a xor b;
    layer2_outputs(2557) <= b;
    layer2_outputs(2558) <= not b;
    layer2_outputs(2559) <= not (a xor b);
    layer2_outputs(2560) <= not a;
    layer2_outputs(2561) <= a and not b;
    layer2_outputs(2562) <= 1'b1;
    layer2_outputs(2563) <= a;
    layer2_outputs(2564) <= a or b;
    layer2_outputs(2565) <= a xor b;
    layer2_outputs(2566) <= not b or a;
    layer2_outputs(2567) <= not (a or b);
    layer2_outputs(2568) <= not (a and b);
    layer2_outputs(2569) <= a and b;
    layer2_outputs(2570) <= not (a and b);
    layer2_outputs(2571) <= not (a and b);
    layer2_outputs(2572) <= a xor b;
    layer2_outputs(2573) <= not (a or b);
    layer2_outputs(2574) <= not (a or b);
    layer2_outputs(2575) <= not (a and b);
    layer2_outputs(2576) <= a and b;
    layer2_outputs(2577) <= not (a or b);
    layer2_outputs(2578) <= a and not b;
    layer2_outputs(2579) <= b and not a;
    layer2_outputs(2580) <= 1'b1;
    layer2_outputs(2581) <= not b;
    layer2_outputs(2582) <= not (a and b);
    layer2_outputs(2583) <= not b;
    layer2_outputs(2584) <= not (a and b);
    layer2_outputs(2585) <= a;
    layer2_outputs(2586) <= not a;
    layer2_outputs(2587) <= b;
    layer2_outputs(2588) <= a;
    layer2_outputs(2589) <= not b or a;
    layer2_outputs(2590) <= a or b;
    layer2_outputs(2591) <= not b;
    layer2_outputs(2592) <= b;
    layer2_outputs(2593) <= not (a or b);
    layer2_outputs(2594) <= b and not a;
    layer2_outputs(2595) <= a or b;
    layer2_outputs(2596) <= 1'b1;
    layer2_outputs(2597) <= b and not a;
    layer2_outputs(2598) <= a or b;
    layer2_outputs(2599) <= not b or a;
    layer2_outputs(2600) <= not (a or b);
    layer2_outputs(2601) <= not b;
    layer2_outputs(2602) <= a;
    layer2_outputs(2603) <= a and b;
    layer2_outputs(2604) <= not b;
    layer2_outputs(2605) <= a;
    layer2_outputs(2606) <= a and not b;
    layer2_outputs(2607) <= not a;
    layer2_outputs(2608) <= a;
    layer2_outputs(2609) <= a xor b;
    layer2_outputs(2610) <= b;
    layer2_outputs(2611) <= not (a xor b);
    layer2_outputs(2612) <= b;
    layer2_outputs(2613) <= a and b;
    layer2_outputs(2614) <= not (a xor b);
    layer2_outputs(2615) <= b and not a;
    layer2_outputs(2616) <= b;
    layer2_outputs(2617) <= not a or b;
    layer2_outputs(2618) <= b and not a;
    layer2_outputs(2619) <= a and not b;
    layer2_outputs(2620) <= not b or a;
    layer2_outputs(2621) <= b;
    layer2_outputs(2622) <= a xor b;
    layer2_outputs(2623) <= a;
    layer2_outputs(2624) <= not (a or b);
    layer2_outputs(2625) <= a;
    layer2_outputs(2626) <= not a or b;
    layer2_outputs(2627) <= b;
    layer2_outputs(2628) <= a and not b;
    layer2_outputs(2629) <= b;
    layer2_outputs(2630) <= b and not a;
    layer2_outputs(2631) <= not a;
    layer2_outputs(2632) <= a;
    layer2_outputs(2633) <= not a or b;
    layer2_outputs(2634) <= a and not b;
    layer2_outputs(2635) <= b and not a;
    layer2_outputs(2636) <= b;
    layer2_outputs(2637) <= not b;
    layer2_outputs(2638) <= a xor b;
    layer2_outputs(2639) <= b;
    layer2_outputs(2640) <= b;
    layer2_outputs(2641) <= not b;
    layer2_outputs(2642) <= b;
    layer2_outputs(2643) <= not (a and b);
    layer2_outputs(2644) <= a;
    layer2_outputs(2645) <= not (a or b);
    layer2_outputs(2646) <= not (a or b);
    layer2_outputs(2647) <= a and b;
    layer2_outputs(2648) <= a and b;
    layer2_outputs(2649) <= a and b;
    layer2_outputs(2650) <= 1'b0;
    layer2_outputs(2651) <= not a;
    layer2_outputs(2652) <= not a or b;
    layer2_outputs(2653) <= not (a xor b);
    layer2_outputs(2654) <= b;
    layer2_outputs(2655) <= a;
    layer2_outputs(2656) <= b;
    layer2_outputs(2657) <= a and not b;
    layer2_outputs(2658) <= not (a and b);
    layer2_outputs(2659) <= a xor b;
    layer2_outputs(2660) <= b;
    layer2_outputs(2661) <= not a;
    layer2_outputs(2662) <= not b;
    layer2_outputs(2663) <= not b or a;
    layer2_outputs(2664) <= a and b;
    layer2_outputs(2665) <= b;
    layer2_outputs(2666) <= not b;
    layer2_outputs(2667) <= not a or b;
    layer2_outputs(2668) <= b;
    layer2_outputs(2669) <= a or b;
    layer2_outputs(2670) <= b;
    layer2_outputs(2671) <= not (a and b);
    layer2_outputs(2672) <= not (a and b);
    layer2_outputs(2673) <= not b;
    layer2_outputs(2674) <= not (a and b);
    layer2_outputs(2675) <= not a;
    layer2_outputs(2676) <= a;
    layer2_outputs(2677) <= a;
    layer2_outputs(2678) <= b;
    layer2_outputs(2679) <= not a;
    layer2_outputs(2680) <= not (a and b);
    layer2_outputs(2681) <= a or b;
    layer2_outputs(2682) <= not b;
    layer2_outputs(2683) <= b;
    layer2_outputs(2684) <= not b or a;
    layer2_outputs(2685) <= b;
    layer2_outputs(2686) <= b;
    layer2_outputs(2687) <= a or b;
    layer2_outputs(2688) <= not (a or b);
    layer2_outputs(2689) <= a and b;
    layer2_outputs(2690) <= not (a and b);
    layer2_outputs(2691) <= not b;
    layer2_outputs(2692) <= a;
    layer2_outputs(2693) <= not b;
    layer2_outputs(2694) <= not b;
    layer2_outputs(2695) <= b and not a;
    layer2_outputs(2696) <= a;
    layer2_outputs(2697) <= not (a and b);
    layer2_outputs(2698) <= a;
    layer2_outputs(2699) <= 1'b1;
    layer2_outputs(2700) <= a;
    layer2_outputs(2701) <= a or b;
    layer2_outputs(2702) <= not b;
    layer2_outputs(2703) <= not (a xor b);
    layer2_outputs(2704) <= not a or b;
    layer2_outputs(2705) <= a or b;
    layer2_outputs(2706) <= not b;
    layer2_outputs(2707) <= 1'b0;
    layer2_outputs(2708) <= not (a xor b);
    layer2_outputs(2709) <= a and b;
    layer2_outputs(2710) <= a or b;
    layer2_outputs(2711) <= a and b;
    layer2_outputs(2712) <= not a;
    layer2_outputs(2713) <= not (a and b);
    layer2_outputs(2714) <= a and not b;
    layer2_outputs(2715) <= a and b;
    layer2_outputs(2716) <= a and b;
    layer2_outputs(2717) <= not b;
    layer2_outputs(2718) <= not (a xor b);
    layer2_outputs(2719) <= a;
    layer2_outputs(2720) <= not (a or b);
    layer2_outputs(2721) <= not b or a;
    layer2_outputs(2722) <= not a;
    layer2_outputs(2723) <= not (a and b);
    layer2_outputs(2724) <= not (a or b);
    layer2_outputs(2725) <= not (a xor b);
    layer2_outputs(2726) <= not b;
    layer2_outputs(2727) <= a xor b;
    layer2_outputs(2728) <= not (a xor b);
    layer2_outputs(2729) <= not (a or b);
    layer2_outputs(2730) <= not (a or b);
    layer2_outputs(2731) <= b;
    layer2_outputs(2732) <= not a or b;
    layer2_outputs(2733) <= not a;
    layer2_outputs(2734) <= 1'b0;
    layer2_outputs(2735) <= a or b;
    layer2_outputs(2736) <= not (a xor b);
    layer2_outputs(2737) <= not (a xor b);
    layer2_outputs(2738) <= not (a and b);
    layer2_outputs(2739) <= a;
    layer2_outputs(2740) <= not (a xor b);
    layer2_outputs(2741) <= a;
    layer2_outputs(2742) <= not b;
    layer2_outputs(2743) <= a;
    layer2_outputs(2744) <= a;
    layer2_outputs(2745) <= a and b;
    layer2_outputs(2746) <= not b;
    layer2_outputs(2747) <= a and b;
    layer2_outputs(2748) <= a and b;
    layer2_outputs(2749) <= a and b;
    layer2_outputs(2750) <= b;
    layer2_outputs(2751) <= a xor b;
    layer2_outputs(2752) <= a;
    layer2_outputs(2753) <= a and b;
    layer2_outputs(2754) <= b and not a;
    layer2_outputs(2755) <= a xor b;
    layer2_outputs(2756) <= not (a and b);
    layer2_outputs(2757) <= 1'b1;
    layer2_outputs(2758) <= a and b;
    layer2_outputs(2759) <= a and b;
    layer2_outputs(2760) <= not a or b;
    layer2_outputs(2761) <= not a or b;
    layer2_outputs(2762) <= a;
    layer2_outputs(2763) <= not (a xor b);
    layer2_outputs(2764) <= a and b;
    layer2_outputs(2765) <= b;
    layer2_outputs(2766) <= a and b;
    layer2_outputs(2767) <= not (a or b);
    layer2_outputs(2768) <= b;
    layer2_outputs(2769) <= not a;
    layer2_outputs(2770) <= not a;
    layer2_outputs(2771) <= b and not a;
    layer2_outputs(2772) <= not a;
    layer2_outputs(2773) <= b and not a;
    layer2_outputs(2774) <= b and not a;
    layer2_outputs(2775) <= not (a or b);
    layer2_outputs(2776) <= b and not a;
    layer2_outputs(2777) <= not a;
    layer2_outputs(2778) <= not (a and b);
    layer2_outputs(2779) <= a;
    layer2_outputs(2780) <= 1'b1;
    layer2_outputs(2781) <= b;
    layer2_outputs(2782) <= not a;
    layer2_outputs(2783) <= not b or a;
    layer2_outputs(2784) <= not b or a;
    layer2_outputs(2785) <= not (a xor b);
    layer2_outputs(2786) <= a and not b;
    layer2_outputs(2787) <= b;
    layer2_outputs(2788) <= not b or a;
    layer2_outputs(2789) <= not a;
    layer2_outputs(2790) <= not (a or b);
    layer2_outputs(2791) <= not (a or b);
    layer2_outputs(2792) <= not b;
    layer2_outputs(2793) <= a xor b;
    layer2_outputs(2794) <= a and not b;
    layer2_outputs(2795) <= 1'b0;
    layer2_outputs(2796) <= not (a xor b);
    layer2_outputs(2797) <= b;
    layer2_outputs(2798) <= not b or a;
    layer2_outputs(2799) <= b and not a;
    layer2_outputs(2800) <= not a;
    layer2_outputs(2801) <= 1'b0;
    layer2_outputs(2802) <= not (a xor b);
    layer2_outputs(2803) <= a and b;
    layer2_outputs(2804) <= a and b;
    layer2_outputs(2805) <= 1'b1;
    layer2_outputs(2806) <= a xor b;
    layer2_outputs(2807) <= a or b;
    layer2_outputs(2808) <= not b;
    layer2_outputs(2809) <= not a or b;
    layer2_outputs(2810) <= a;
    layer2_outputs(2811) <= b and not a;
    layer2_outputs(2812) <= a;
    layer2_outputs(2813) <= not (a xor b);
    layer2_outputs(2814) <= b;
    layer2_outputs(2815) <= not (a xor b);
    layer2_outputs(2816) <= not (a or b);
    layer2_outputs(2817) <= a xor b;
    layer2_outputs(2818) <= not b or a;
    layer2_outputs(2819) <= not b;
    layer2_outputs(2820) <= a and not b;
    layer2_outputs(2821) <= a;
    layer2_outputs(2822) <= 1'b1;
    layer2_outputs(2823) <= not b;
    layer2_outputs(2824) <= a;
    layer2_outputs(2825) <= b and not a;
    layer2_outputs(2826) <= a and not b;
    layer2_outputs(2827) <= not b or a;
    layer2_outputs(2828) <= not b or a;
    layer2_outputs(2829) <= not a;
    layer2_outputs(2830) <= b;
    layer2_outputs(2831) <= not (a and b);
    layer2_outputs(2832) <= a and not b;
    layer2_outputs(2833) <= not a or b;
    layer2_outputs(2834) <= not b;
    layer2_outputs(2835) <= not b;
    layer2_outputs(2836) <= a;
    layer2_outputs(2837) <= not a or b;
    layer2_outputs(2838) <= not (a xor b);
    layer2_outputs(2839) <= not (a xor b);
    layer2_outputs(2840) <= not b or a;
    layer2_outputs(2841) <= b;
    layer2_outputs(2842) <= not a;
    layer2_outputs(2843) <= not b or a;
    layer2_outputs(2844) <= not b;
    layer2_outputs(2845) <= not (a or b);
    layer2_outputs(2846) <= not a or b;
    layer2_outputs(2847) <= a and b;
    layer2_outputs(2848) <= b;
    layer2_outputs(2849) <= a;
    layer2_outputs(2850) <= a or b;
    layer2_outputs(2851) <= not b or a;
    layer2_outputs(2852) <= not a;
    layer2_outputs(2853) <= not b;
    layer2_outputs(2854) <= not a or b;
    layer2_outputs(2855) <= a;
    layer2_outputs(2856) <= not b or a;
    layer2_outputs(2857) <= a;
    layer2_outputs(2858) <= not b;
    layer2_outputs(2859) <= not b;
    layer2_outputs(2860) <= not (a or b);
    layer2_outputs(2861) <= a and not b;
    layer2_outputs(2862) <= a and b;
    layer2_outputs(2863) <= not (a and b);
    layer2_outputs(2864) <= not a or b;
    layer2_outputs(2865) <= not b;
    layer2_outputs(2866) <= not b;
    layer2_outputs(2867) <= not b;
    layer2_outputs(2868) <= not (a and b);
    layer2_outputs(2869) <= a or b;
    layer2_outputs(2870) <= a and not b;
    layer2_outputs(2871) <= b and not a;
    layer2_outputs(2872) <= not a or b;
    layer2_outputs(2873) <= b;
    layer2_outputs(2874) <= a and not b;
    layer2_outputs(2875) <= b and not a;
    layer2_outputs(2876) <= not a;
    layer2_outputs(2877) <= 1'b0;
    layer2_outputs(2878) <= a;
    layer2_outputs(2879) <= b and not a;
    layer2_outputs(2880) <= a and not b;
    layer2_outputs(2881) <= a xor b;
    layer2_outputs(2882) <= not a;
    layer2_outputs(2883) <= not (a or b);
    layer2_outputs(2884) <= a;
    layer2_outputs(2885) <= a and not b;
    layer2_outputs(2886) <= not a;
    layer2_outputs(2887) <= not a;
    layer2_outputs(2888) <= not (a and b);
    layer2_outputs(2889) <= not a;
    layer2_outputs(2890) <= not a or b;
    layer2_outputs(2891) <= b and not a;
    layer2_outputs(2892) <= a and b;
    layer2_outputs(2893) <= not (a and b);
    layer2_outputs(2894) <= 1'b1;
    layer2_outputs(2895) <= a and b;
    layer2_outputs(2896) <= not b;
    layer2_outputs(2897) <= a;
    layer2_outputs(2898) <= not (a and b);
    layer2_outputs(2899) <= not a or b;
    layer2_outputs(2900) <= a;
    layer2_outputs(2901) <= not b or a;
    layer2_outputs(2902) <= a or b;
    layer2_outputs(2903) <= not (a xor b);
    layer2_outputs(2904) <= not b;
    layer2_outputs(2905) <= a or b;
    layer2_outputs(2906) <= not b;
    layer2_outputs(2907) <= not (a or b);
    layer2_outputs(2908) <= a and not b;
    layer2_outputs(2909) <= not b;
    layer2_outputs(2910) <= 1'b0;
    layer2_outputs(2911) <= a or b;
    layer2_outputs(2912) <= a;
    layer2_outputs(2913) <= not b;
    layer2_outputs(2914) <= not (a or b);
    layer2_outputs(2915) <= not a;
    layer2_outputs(2916) <= not a;
    layer2_outputs(2917) <= not (a xor b);
    layer2_outputs(2918) <= not a;
    layer2_outputs(2919) <= not b;
    layer2_outputs(2920) <= not (a and b);
    layer2_outputs(2921) <= a;
    layer2_outputs(2922) <= a or b;
    layer2_outputs(2923) <= a and not b;
    layer2_outputs(2924) <= b and not a;
    layer2_outputs(2925) <= a and b;
    layer2_outputs(2926) <= not a;
    layer2_outputs(2927) <= b;
    layer2_outputs(2928) <= not (a xor b);
    layer2_outputs(2929) <= a;
    layer2_outputs(2930) <= not (a and b);
    layer2_outputs(2931) <= b and not a;
    layer2_outputs(2932) <= a and not b;
    layer2_outputs(2933) <= a;
    layer2_outputs(2934) <= b;
    layer2_outputs(2935) <= a and b;
    layer2_outputs(2936) <= a;
    layer2_outputs(2937) <= not a or b;
    layer2_outputs(2938) <= a xor b;
    layer2_outputs(2939) <= b;
    layer2_outputs(2940) <= a or b;
    layer2_outputs(2941) <= not b;
    layer2_outputs(2942) <= not a;
    layer2_outputs(2943) <= a xor b;
    layer2_outputs(2944) <= not (a and b);
    layer2_outputs(2945) <= b and not a;
    layer2_outputs(2946) <= not (a or b);
    layer2_outputs(2947) <= not b;
    layer2_outputs(2948) <= not (a xor b);
    layer2_outputs(2949) <= not b;
    layer2_outputs(2950) <= not (a or b);
    layer2_outputs(2951) <= a;
    layer2_outputs(2952) <= a and b;
    layer2_outputs(2953) <= b;
    layer2_outputs(2954) <= a or b;
    layer2_outputs(2955) <= b;
    layer2_outputs(2956) <= b;
    layer2_outputs(2957) <= not b;
    layer2_outputs(2958) <= not a or b;
    layer2_outputs(2959) <= not (a and b);
    layer2_outputs(2960) <= not (a xor b);
    layer2_outputs(2961) <= not (a or b);
    layer2_outputs(2962) <= not (a or b);
    layer2_outputs(2963) <= not b;
    layer2_outputs(2964) <= 1'b0;
    layer2_outputs(2965) <= a xor b;
    layer2_outputs(2966) <= a and b;
    layer2_outputs(2967) <= a and b;
    layer2_outputs(2968) <= 1'b0;
    layer2_outputs(2969) <= not a or b;
    layer2_outputs(2970) <= not a;
    layer2_outputs(2971) <= a or b;
    layer2_outputs(2972) <= a and not b;
    layer2_outputs(2973) <= not a;
    layer2_outputs(2974) <= a or b;
    layer2_outputs(2975) <= 1'b1;
    layer2_outputs(2976) <= not b;
    layer2_outputs(2977) <= b;
    layer2_outputs(2978) <= not (a xor b);
    layer2_outputs(2979) <= b;
    layer2_outputs(2980) <= not (a xor b);
    layer2_outputs(2981) <= not (a and b);
    layer2_outputs(2982) <= a;
    layer2_outputs(2983) <= 1'b0;
    layer2_outputs(2984) <= not b;
    layer2_outputs(2985) <= not a or b;
    layer2_outputs(2986) <= a and b;
    layer2_outputs(2987) <= a;
    layer2_outputs(2988) <= b;
    layer2_outputs(2989) <= a and b;
    layer2_outputs(2990) <= a and not b;
    layer2_outputs(2991) <= b;
    layer2_outputs(2992) <= not (a or b);
    layer2_outputs(2993) <= b;
    layer2_outputs(2994) <= b;
    layer2_outputs(2995) <= a xor b;
    layer2_outputs(2996) <= a or b;
    layer2_outputs(2997) <= not (a or b);
    layer2_outputs(2998) <= not b;
    layer2_outputs(2999) <= b;
    layer2_outputs(3000) <= not b;
    layer2_outputs(3001) <= a and not b;
    layer2_outputs(3002) <= a or b;
    layer2_outputs(3003) <= b and not a;
    layer2_outputs(3004) <= a;
    layer2_outputs(3005) <= a and b;
    layer2_outputs(3006) <= b and not a;
    layer2_outputs(3007) <= b;
    layer2_outputs(3008) <= a and not b;
    layer2_outputs(3009) <= not b;
    layer2_outputs(3010) <= not a or b;
    layer2_outputs(3011) <= 1'b1;
    layer2_outputs(3012) <= a or b;
    layer2_outputs(3013) <= a;
    layer2_outputs(3014) <= a or b;
    layer2_outputs(3015) <= a and not b;
    layer2_outputs(3016) <= not (a xor b);
    layer2_outputs(3017) <= not b;
    layer2_outputs(3018) <= not (a xor b);
    layer2_outputs(3019) <= not b;
    layer2_outputs(3020) <= b;
    layer2_outputs(3021) <= not b;
    layer2_outputs(3022) <= a and not b;
    layer2_outputs(3023) <= b and not a;
    layer2_outputs(3024) <= a and not b;
    layer2_outputs(3025) <= 1'b0;
    layer2_outputs(3026) <= 1'b1;
    layer2_outputs(3027) <= a and not b;
    layer2_outputs(3028) <= not b;
    layer2_outputs(3029) <= not a;
    layer2_outputs(3030) <= not b;
    layer2_outputs(3031) <= not a or b;
    layer2_outputs(3032) <= a xor b;
    layer2_outputs(3033) <= b and not a;
    layer2_outputs(3034) <= 1'b1;
    layer2_outputs(3035) <= a;
    layer2_outputs(3036) <= not b or a;
    layer2_outputs(3037) <= a;
    layer2_outputs(3038) <= a or b;
    layer2_outputs(3039) <= b;
    layer2_outputs(3040) <= not a;
    layer2_outputs(3041) <= not (a or b);
    layer2_outputs(3042) <= not (a or b);
    layer2_outputs(3043) <= a and b;
    layer2_outputs(3044) <= a;
    layer2_outputs(3045) <= not a or b;
    layer2_outputs(3046) <= 1'b1;
    layer2_outputs(3047) <= 1'b1;
    layer2_outputs(3048) <= b and not a;
    layer2_outputs(3049) <= not b or a;
    layer2_outputs(3050) <= a or b;
    layer2_outputs(3051) <= not a;
    layer2_outputs(3052) <= a and b;
    layer2_outputs(3053) <= a and b;
    layer2_outputs(3054) <= a and b;
    layer2_outputs(3055) <= a and b;
    layer2_outputs(3056) <= 1'b0;
    layer2_outputs(3057) <= not (a or b);
    layer2_outputs(3058) <= b;
    layer2_outputs(3059) <= not (a or b);
    layer2_outputs(3060) <= not b;
    layer2_outputs(3061) <= b;
    layer2_outputs(3062) <= b;
    layer2_outputs(3063) <= not a or b;
    layer2_outputs(3064) <= not (a or b);
    layer2_outputs(3065) <= a and b;
    layer2_outputs(3066) <= a;
    layer2_outputs(3067) <= not (a and b);
    layer2_outputs(3068) <= not a;
    layer2_outputs(3069) <= a;
    layer2_outputs(3070) <= a and not b;
    layer2_outputs(3071) <= a or b;
    layer2_outputs(3072) <= a and b;
    layer2_outputs(3073) <= a;
    layer2_outputs(3074) <= a and b;
    layer2_outputs(3075) <= b and not a;
    layer2_outputs(3076) <= not b;
    layer2_outputs(3077) <= a or b;
    layer2_outputs(3078) <= b;
    layer2_outputs(3079) <= a;
    layer2_outputs(3080) <= a and not b;
    layer2_outputs(3081) <= 1'b1;
    layer2_outputs(3082) <= not a;
    layer2_outputs(3083) <= 1'b1;
    layer2_outputs(3084) <= a xor b;
    layer2_outputs(3085) <= a;
    layer2_outputs(3086) <= b and not a;
    layer2_outputs(3087) <= not (a xor b);
    layer2_outputs(3088) <= a xor b;
    layer2_outputs(3089) <= not a;
    layer2_outputs(3090) <= not (a and b);
    layer2_outputs(3091) <= not (a and b);
    layer2_outputs(3092) <= not a;
    layer2_outputs(3093) <= a or b;
    layer2_outputs(3094) <= a;
    layer2_outputs(3095) <= not (a xor b);
    layer2_outputs(3096) <= not b or a;
    layer2_outputs(3097) <= b;
    layer2_outputs(3098) <= not b or a;
    layer2_outputs(3099) <= a xor b;
    layer2_outputs(3100) <= not (a xor b);
    layer2_outputs(3101) <= not a or b;
    layer2_outputs(3102) <= b;
    layer2_outputs(3103) <= a;
    layer2_outputs(3104) <= a and not b;
    layer2_outputs(3105) <= b and not a;
    layer2_outputs(3106) <= a and not b;
    layer2_outputs(3107) <= a;
    layer2_outputs(3108) <= b;
    layer2_outputs(3109) <= a or b;
    layer2_outputs(3110) <= not (a or b);
    layer2_outputs(3111) <= not b;
    layer2_outputs(3112) <= not b or a;
    layer2_outputs(3113) <= a xor b;
    layer2_outputs(3114) <= not a or b;
    layer2_outputs(3115) <= b and not a;
    layer2_outputs(3116) <= b;
    layer2_outputs(3117) <= a and b;
    layer2_outputs(3118) <= not (a or b);
    layer2_outputs(3119) <= b;
    layer2_outputs(3120) <= a;
    layer2_outputs(3121) <= not b;
    layer2_outputs(3122) <= a;
    layer2_outputs(3123) <= b and not a;
    layer2_outputs(3124) <= a;
    layer2_outputs(3125) <= b and not a;
    layer2_outputs(3126) <= a and b;
    layer2_outputs(3127) <= not b;
    layer2_outputs(3128) <= not (a xor b);
    layer2_outputs(3129) <= a and b;
    layer2_outputs(3130) <= not b;
    layer2_outputs(3131) <= not b;
    layer2_outputs(3132) <= not (a and b);
    layer2_outputs(3133) <= not a;
    layer2_outputs(3134) <= b and not a;
    layer2_outputs(3135) <= not b;
    layer2_outputs(3136) <= not b;
    layer2_outputs(3137) <= not (a and b);
    layer2_outputs(3138) <= a and not b;
    layer2_outputs(3139) <= not a or b;
    layer2_outputs(3140) <= a xor b;
    layer2_outputs(3141) <= a or b;
    layer2_outputs(3142) <= not a;
    layer2_outputs(3143) <= not a or b;
    layer2_outputs(3144) <= a or b;
    layer2_outputs(3145) <= b and not a;
    layer2_outputs(3146) <= not a;
    layer2_outputs(3147) <= b;
    layer2_outputs(3148) <= a and b;
    layer2_outputs(3149) <= not a or b;
    layer2_outputs(3150) <= b;
    layer2_outputs(3151) <= a or b;
    layer2_outputs(3152) <= not (a or b);
    layer2_outputs(3153) <= a xor b;
    layer2_outputs(3154) <= not (a xor b);
    layer2_outputs(3155) <= not a;
    layer2_outputs(3156) <= a or b;
    layer2_outputs(3157) <= a xor b;
    layer2_outputs(3158) <= b;
    layer2_outputs(3159) <= not (a xor b);
    layer2_outputs(3160) <= b and not a;
    layer2_outputs(3161) <= not b or a;
    layer2_outputs(3162) <= a or b;
    layer2_outputs(3163) <= not (a and b);
    layer2_outputs(3164) <= a or b;
    layer2_outputs(3165) <= a;
    layer2_outputs(3166) <= not b;
    layer2_outputs(3167) <= not (a or b);
    layer2_outputs(3168) <= 1'b0;
    layer2_outputs(3169) <= not b;
    layer2_outputs(3170) <= b and not a;
    layer2_outputs(3171) <= a xor b;
    layer2_outputs(3172) <= b;
    layer2_outputs(3173) <= not a or b;
    layer2_outputs(3174) <= a;
    layer2_outputs(3175) <= a;
    layer2_outputs(3176) <= a;
    layer2_outputs(3177) <= not a;
    layer2_outputs(3178) <= not (a and b);
    layer2_outputs(3179) <= not (a or b);
    layer2_outputs(3180) <= 1'b0;
    layer2_outputs(3181) <= a and b;
    layer2_outputs(3182) <= a and not b;
    layer2_outputs(3183) <= not a;
    layer2_outputs(3184) <= a or b;
    layer2_outputs(3185) <= a;
    layer2_outputs(3186) <= not (a xor b);
    layer2_outputs(3187) <= not (a xor b);
    layer2_outputs(3188) <= a and not b;
    layer2_outputs(3189) <= b and not a;
    layer2_outputs(3190) <= not b or a;
    layer2_outputs(3191) <= a xor b;
    layer2_outputs(3192) <= not a;
    layer2_outputs(3193) <= not a or b;
    layer2_outputs(3194) <= 1'b1;
    layer2_outputs(3195) <= not (a and b);
    layer2_outputs(3196) <= a and b;
    layer2_outputs(3197) <= not (a and b);
    layer2_outputs(3198) <= not b or a;
    layer2_outputs(3199) <= 1'b0;
    layer2_outputs(3200) <= not b or a;
    layer2_outputs(3201) <= b;
    layer2_outputs(3202) <= not (a and b);
    layer2_outputs(3203) <= a and not b;
    layer2_outputs(3204) <= b and not a;
    layer2_outputs(3205) <= b and not a;
    layer2_outputs(3206) <= not b or a;
    layer2_outputs(3207) <= not a;
    layer2_outputs(3208) <= not (a or b);
    layer2_outputs(3209) <= not b;
    layer2_outputs(3210) <= not a;
    layer2_outputs(3211) <= not (a or b);
    layer2_outputs(3212) <= not (a xor b);
    layer2_outputs(3213) <= a and b;
    layer2_outputs(3214) <= not a;
    layer2_outputs(3215) <= b;
    layer2_outputs(3216) <= not a or b;
    layer2_outputs(3217) <= not (a xor b);
    layer2_outputs(3218) <= a;
    layer2_outputs(3219) <= b;
    layer2_outputs(3220) <= a;
    layer2_outputs(3221) <= 1'b0;
    layer2_outputs(3222) <= not (a or b);
    layer2_outputs(3223) <= not b;
    layer2_outputs(3224) <= not b;
    layer2_outputs(3225) <= not (a xor b);
    layer2_outputs(3226) <= a and b;
    layer2_outputs(3227) <= b;
    layer2_outputs(3228) <= not b;
    layer2_outputs(3229) <= b;
    layer2_outputs(3230) <= b;
    layer2_outputs(3231) <= not b;
    layer2_outputs(3232) <= a;
    layer2_outputs(3233) <= not b or a;
    layer2_outputs(3234) <= not (a or b);
    layer2_outputs(3235) <= a and b;
    layer2_outputs(3236) <= a or b;
    layer2_outputs(3237) <= not (a or b);
    layer2_outputs(3238) <= a or b;
    layer2_outputs(3239) <= a;
    layer2_outputs(3240) <= a or b;
    layer2_outputs(3241) <= not a;
    layer2_outputs(3242) <= a or b;
    layer2_outputs(3243) <= a and b;
    layer2_outputs(3244) <= 1'b0;
    layer2_outputs(3245) <= not a;
    layer2_outputs(3246) <= not a or b;
    layer2_outputs(3247) <= not a;
    layer2_outputs(3248) <= a and b;
    layer2_outputs(3249) <= a xor b;
    layer2_outputs(3250) <= not b;
    layer2_outputs(3251) <= b and not a;
    layer2_outputs(3252) <= not b;
    layer2_outputs(3253) <= not b;
    layer2_outputs(3254) <= b;
    layer2_outputs(3255) <= b and not a;
    layer2_outputs(3256) <= not (a or b);
    layer2_outputs(3257) <= a and b;
    layer2_outputs(3258) <= not b;
    layer2_outputs(3259) <= b;
    layer2_outputs(3260) <= not a;
    layer2_outputs(3261) <= a and not b;
    layer2_outputs(3262) <= a xor b;
    layer2_outputs(3263) <= a xor b;
    layer2_outputs(3264) <= not (a xor b);
    layer2_outputs(3265) <= a or b;
    layer2_outputs(3266) <= not a;
    layer2_outputs(3267) <= b and not a;
    layer2_outputs(3268) <= not b;
    layer2_outputs(3269) <= not b;
    layer2_outputs(3270) <= not b;
    layer2_outputs(3271) <= not b;
    layer2_outputs(3272) <= not b;
    layer2_outputs(3273) <= not (a and b);
    layer2_outputs(3274) <= a;
    layer2_outputs(3275) <= not (a or b);
    layer2_outputs(3276) <= not a;
    layer2_outputs(3277) <= a;
    layer2_outputs(3278) <= a;
    layer2_outputs(3279) <= not a;
    layer2_outputs(3280) <= not a;
    layer2_outputs(3281) <= not (a and b);
    layer2_outputs(3282) <= a and b;
    layer2_outputs(3283) <= 1'b1;
    layer2_outputs(3284) <= b and not a;
    layer2_outputs(3285) <= a;
    layer2_outputs(3286) <= not a;
    layer2_outputs(3287) <= not b;
    layer2_outputs(3288) <= a and not b;
    layer2_outputs(3289) <= not (a and b);
    layer2_outputs(3290) <= not a;
    layer2_outputs(3291) <= b;
    layer2_outputs(3292) <= not (a and b);
    layer2_outputs(3293) <= not a or b;
    layer2_outputs(3294) <= 1'b0;
    layer2_outputs(3295) <= b;
    layer2_outputs(3296) <= a and b;
    layer2_outputs(3297) <= not (a and b);
    layer2_outputs(3298) <= not a;
    layer2_outputs(3299) <= a and not b;
    layer2_outputs(3300) <= not b;
    layer2_outputs(3301) <= 1'b1;
    layer2_outputs(3302) <= a or b;
    layer2_outputs(3303) <= 1'b1;
    layer2_outputs(3304) <= not (a xor b);
    layer2_outputs(3305) <= not (a xor b);
    layer2_outputs(3306) <= not a;
    layer2_outputs(3307) <= not b;
    layer2_outputs(3308) <= a and not b;
    layer2_outputs(3309) <= a and b;
    layer2_outputs(3310) <= not (a or b);
    layer2_outputs(3311) <= b;
    layer2_outputs(3312) <= a or b;
    layer2_outputs(3313) <= a or b;
    layer2_outputs(3314) <= 1'b1;
    layer2_outputs(3315) <= not b or a;
    layer2_outputs(3316) <= a or b;
    layer2_outputs(3317) <= b;
    layer2_outputs(3318) <= not (a and b);
    layer2_outputs(3319) <= not b;
    layer2_outputs(3320) <= not b;
    layer2_outputs(3321) <= not b;
    layer2_outputs(3322) <= b and not a;
    layer2_outputs(3323) <= not (a or b);
    layer2_outputs(3324) <= a or b;
    layer2_outputs(3325) <= not a or b;
    layer2_outputs(3326) <= not a;
    layer2_outputs(3327) <= not (a or b);
    layer2_outputs(3328) <= a;
    layer2_outputs(3329) <= not a or b;
    layer2_outputs(3330) <= a and not b;
    layer2_outputs(3331) <= b;
    layer2_outputs(3332) <= not b;
    layer2_outputs(3333) <= not (a or b);
    layer2_outputs(3334) <= a and not b;
    layer2_outputs(3335) <= not b;
    layer2_outputs(3336) <= a;
    layer2_outputs(3337) <= b;
    layer2_outputs(3338) <= not b;
    layer2_outputs(3339) <= not b;
    layer2_outputs(3340) <= 1'b1;
    layer2_outputs(3341) <= a and b;
    layer2_outputs(3342) <= not (a and b);
    layer2_outputs(3343) <= a and not b;
    layer2_outputs(3344) <= not (a or b);
    layer2_outputs(3345) <= a;
    layer2_outputs(3346) <= not b;
    layer2_outputs(3347) <= not b;
    layer2_outputs(3348) <= not (a or b);
    layer2_outputs(3349) <= b and not a;
    layer2_outputs(3350) <= b and not a;
    layer2_outputs(3351) <= a xor b;
    layer2_outputs(3352) <= b;
    layer2_outputs(3353) <= not (a and b);
    layer2_outputs(3354) <= not (a or b);
    layer2_outputs(3355) <= not (a xor b);
    layer2_outputs(3356) <= not (a and b);
    layer2_outputs(3357) <= a;
    layer2_outputs(3358) <= 1'b1;
    layer2_outputs(3359) <= a and b;
    layer2_outputs(3360) <= not a or b;
    layer2_outputs(3361) <= not a or b;
    layer2_outputs(3362) <= not a;
    layer2_outputs(3363) <= not a or b;
    layer2_outputs(3364) <= not b or a;
    layer2_outputs(3365) <= not (a and b);
    layer2_outputs(3366) <= a and not b;
    layer2_outputs(3367) <= b and not a;
    layer2_outputs(3368) <= a or b;
    layer2_outputs(3369) <= not a;
    layer2_outputs(3370) <= not a;
    layer2_outputs(3371) <= a and b;
    layer2_outputs(3372) <= a;
    layer2_outputs(3373) <= b and not a;
    layer2_outputs(3374) <= b;
    layer2_outputs(3375) <= a or b;
    layer2_outputs(3376) <= a and b;
    layer2_outputs(3377) <= not b;
    layer2_outputs(3378) <= not b;
    layer2_outputs(3379) <= a and not b;
    layer2_outputs(3380) <= not b;
    layer2_outputs(3381) <= not b or a;
    layer2_outputs(3382) <= not b or a;
    layer2_outputs(3383) <= b;
    layer2_outputs(3384) <= not (a or b);
    layer2_outputs(3385) <= a;
    layer2_outputs(3386) <= a xor b;
    layer2_outputs(3387) <= not a;
    layer2_outputs(3388) <= a or b;
    layer2_outputs(3389) <= a xor b;
    layer2_outputs(3390) <= not b;
    layer2_outputs(3391) <= b and not a;
    layer2_outputs(3392) <= 1'b0;
    layer2_outputs(3393) <= 1'b1;
    layer2_outputs(3394) <= 1'b1;
    layer2_outputs(3395) <= b and not a;
    layer2_outputs(3396) <= not a;
    layer2_outputs(3397) <= not a;
    layer2_outputs(3398) <= not b;
    layer2_outputs(3399) <= a and not b;
    layer2_outputs(3400) <= b;
    layer2_outputs(3401) <= a;
    layer2_outputs(3402) <= not a;
    layer2_outputs(3403) <= b and not a;
    layer2_outputs(3404) <= not b;
    layer2_outputs(3405) <= not b or a;
    layer2_outputs(3406) <= not a;
    layer2_outputs(3407) <= not b;
    layer2_outputs(3408) <= not (a or b);
    layer2_outputs(3409) <= not b or a;
    layer2_outputs(3410) <= not a;
    layer2_outputs(3411) <= not (a and b);
    layer2_outputs(3412) <= a;
    layer2_outputs(3413) <= not a or b;
    layer2_outputs(3414) <= not (a or b);
    layer2_outputs(3415) <= a and b;
    layer2_outputs(3416) <= not a or b;
    layer2_outputs(3417) <= b;
    layer2_outputs(3418) <= not (a and b);
    layer2_outputs(3419) <= a and not b;
    layer2_outputs(3420) <= not b;
    layer2_outputs(3421) <= a and not b;
    layer2_outputs(3422) <= not (a and b);
    layer2_outputs(3423) <= not a or b;
    layer2_outputs(3424) <= not b or a;
    layer2_outputs(3425) <= not b;
    layer2_outputs(3426) <= b;
    layer2_outputs(3427) <= not b;
    layer2_outputs(3428) <= not (a and b);
    layer2_outputs(3429) <= not a or b;
    layer2_outputs(3430) <= not b;
    layer2_outputs(3431) <= not a;
    layer2_outputs(3432) <= b;
    layer2_outputs(3433) <= not a;
    layer2_outputs(3434) <= a;
    layer2_outputs(3435) <= not (a and b);
    layer2_outputs(3436) <= not (a or b);
    layer2_outputs(3437) <= 1'b0;
    layer2_outputs(3438) <= not (a or b);
    layer2_outputs(3439) <= not a or b;
    layer2_outputs(3440) <= a and not b;
    layer2_outputs(3441) <= b;
    layer2_outputs(3442) <= a;
    layer2_outputs(3443) <= a;
    layer2_outputs(3444) <= a or b;
    layer2_outputs(3445) <= a and not b;
    layer2_outputs(3446) <= 1'b1;
    layer2_outputs(3447) <= not a or b;
    layer2_outputs(3448) <= 1'b1;
    layer2_outputs(3449) <= not b or a;
    layer2_outputs(3450) <= not a;
    layer2_outputs(3451) <= a xor b;
    layer2_outputs(3452) <= a and b;
    layer2_outputs(3453) <= b;
    layer2_outputs(3454) <= a or b;
    layer2_outputs(3455) <= not a;
    layer2_outputs(3456) <= a;
    layer2_outputs(3457) <= not (a and b);
    layer2_outputs(3458) <= not (a and b);
    layer2_outputs(3459) <= not a or b;
    layer2_outputs(3460) <= b;
    layer2_outputs(3461) <= b and not a;
    layer2_outputs(3462) <= not a or b;
    layer2_outputs(3463) <= a and b;
    layer2_outputs(3464) <= a;
    layer2_outputs(3465) <= not b;
    layer2_outputs(3466) <= a;
    layer2_outputs(3467) <= a;
    layer2_outputs(3468) <= not b;
    layer2_outputs(3469) <= a xor b;
    layer2_outputs(3470) <= a;
    layer2_outputs(3471) <= a;
    layer2_outputs(3472) <= b;
    layer2_outputs(3473) <= a;
    layer2_outputs(3474) <= not a;
    layer2_outputs(3475) <= a xor b;
    layer2_outputs(3476) <= a xor b;
    layer2_outputs(3477) <= a;
    layer2_outputs(3478) <= b and not a;
    layer2_outputs(3479) <= not b or a;
    layer2_outputs(3480) <= not (a and b);
    layer2_outputs(3481) <= a or b;
    layer2_outputs(3482) <= not b or a;
    layer2_outputs(3483) <= a;
    layer2_outputs(3484) <= b and not a;
    layer2_outputs(3485) <= a xor b;
    layer2_outputs(3486) <= not a;
    layer2_outputs(3487) <= not (a xor b);
    layer2_outputs(3488) <= not b or a;
    layer2_outputs(3489) <= b;
    layer2_outputs(3490) <= b and not a;
    layer2_outputs(3491) <= not a;
    layer2_outputs(3492) <= a and not b;
    layer2_outputs(3493) <= a or b;
    layer2_outputs(3494) <= a;
    layer2_outputs(3495) <= not (a xor b);
    layer2_outputs(3496) <= not (a xor b);
    layer2_outputs(3497) <= not a;
    layer2_outputs(3498) <= a or b;
    layer2_outputs(3499) <= not b or a;
    layer2_outputs(3500) <= not (a or b);
    layer2_outputs(3501) <= a and not b;
    layer2_outputs(3502) <= b and not a;
    layer2_outputs(3503) <= not b;
    layer2_outputs(3504) <= b;
    layer2_outputs(3505) <= not a or b;
    layer2_outputs(3506) <= not a or b;
    layer2_outputs(3507) <= not a;
    layer2_outputs(3508) <= a or b;
    layer2_outputs(3509) <= not b;
    layer2_outputs(3510) <= a or b;
    layer2_outputs(3511) <= not a;
    layer2_outputs(3512) <= 1'b0;
    layer2_outputs(3513) <= not (a and b);
    layer2_outputs(3514) <= a and b;
    layer2_outputs(3515) <= a;
    layer2_outputs(3516) <= b;
    layer2_outputs(3517) <= b and not a;
    layer2_outputs(3518) <= b and not a;
    layer2_outputs(3519) <= a;
    layer2_outputs(3520) <= a xor b;
    layer2_outputs(3521) <= not a;
    layer2_outputs(3522) <= not (a and b);
    layer2_outputs(3523) <= not (a or b);
    layer2_outputs(3524) <= b;
    layer2_outputs(3525) <= b and not a;
    layer2_outputs(3526) <= not (a or b);
    layer2_outputs(3527) <= not (a xor b);
    layer2_outputs(3528) <= b;
    layer2_outputs(3529) <= b;
    layer2_outputs(3530) <= not a;
    layer2_outputs(3531) <= a or b;
    layer2_outputs(3532) <= not a or b;
    layer2_outputs(3533) <= not a;
    layer2_outputs(3534) <= 1'b1;
    layer2_outputs(3535) <= a and b;
    layer2_outputs(3536) <= b and not a;
    layer2_outputs(3537) <= 1'b0;
    layer2_outputs(3538) <= not b or a;
    layer2_outputs(3539) <= not (a xor b);
    layer2_outputs(3540) <= a and not b;
    layer2_outputs(3541) <= not a or b;
    layer2_outputs(3542) <= b;
    layer2_outputs(3543) <= a;
    layer2_outputs(3544) <= b;
    layer2_outputs(3545) <= b and not a;
    layer2_outputs(3546) <= a and b;
    layer2_outputs(3547) <= b and not a;
    layer2_outputs(3548) <= not b;
    layer2_outputs(3549) <= a and b;
    layer2_outputs(3550) <= not b or a;
    layer2_outputs(3551) <= not (a and b);
    layer2_outputs(3552) <= not b;
    layer2_outputs(3553) <= not b or a;
    layer2_outputs(3554) <= 1'b1;
    layer2_outputs(3555) <= b;
    layer2_outputs(3556) <= a and not b;
    layer2_outputs(3557) <= a and not b;
    layer2_outputs(3558) <= not a;
    layer2_outputs(3559) <= a xor b;
    layer2_outputs(3560) <= not (a or b);
    layer2_outputs(3561) <= b;
    layer2_outputs(3562) <= a and not b;
    layer2_outputs(3563) <= not a or b;
    layer2_outputs(3564) <= not b;
    layer2_outputs(3565) <= a or b;
    layer2_outputs(3566) <= a and not b;
    layer2_outputs(3567) <= not (a xor b);
    layer2_outputs(3568) <= not a;
    layer2_outputs(3569) <= b;
    layer2_outputs(3570) <= not b;
    layer2_outputs(3571) <= a and not b;
    layer2_outputs(3572) <= not b or a;
    layer2_outputs(3573) <= not a or b;
    layer2_outputs(3574) <= not b;
    layer2_outputs(3575) <= a and not b;
    layer2_outputs(3576) <= not (a xor b);
    layer2_outputs(3577) <= not (a and b);
    layer2_outputs(3578) <= a and not b;
    layer2_outputs(3579) <= a and not b;
    layer2_outputs(3580) <= a;
    layer2_outputs(3581) <= not (a and b);
    layer2_outputs(3582) <= not (a and b);
    layer2_outputs(3583) <= a;
    layer2_outputs(3584) <= a and not b;
    layer2_outputs(3585) <= b and not a;
    layer2_outputs(3586) <= 1'b1;
    layer2_outputs(3587) <= b;
    layer2_outputs(3588) <= not a;
    layer2_outputs(3589) <= a and b;
    layer2_outputs(3590) <= not (a or b);
    layer2_outputs(3591) <= b;
    layer2_outputs(3592) <= not (a xor b);
    layer2_outputs(3593) <= a or b;
    layer2_outputs(3594) <= b;
    layer2_outputs(3595) <= a;
    layer2_outputs(3596) <= a and b;
    layer2_outputs(3597) <= not a or b;
    layer2_outputs(3598) <= not a;
    layer2_outputs(3599) <= not (a and b);
    layer2_outputs(3600) <= b and not a;
    layer2_outputs(3601) <= not a or b;
    layer2_outputs(3602) <= not b;
    layer2_outputs(3603) <= not b;
    layer2_outputs(3604) <= not b;
    layer2_outputs(3605) <= b;
    layer2_outputs(3606) <= a or b;
    layer2_outputs(3607) <= not a;
    layer2_outputs(3608) <= b and not a;
    layer2_outputs(3609) <= b;
    layer2_outputs(3610) <= a;
    layer2_outputs(3611) <= not (a or b);
    layer2_outputs(3612) <= not b;
    layer2_outputs(3613) <= a or b;
    layer2_outputs(3614) <= not (a and b);
    layer2_outputs(3615) <= not b;
    layer2_outputs(3616) <= not b or a;
    layer2_outputs(3617) <= not b;
    layer2_outputs(3618) <= a xor b;
    layer2_outputs(3619) <= b and not a;
    layer2_outputs(3620) <= a;
    layer2_outputs(3621) <= a;
    layer2_outputs(3622) <= a and not b;
    layer2_outputs(3623) <= not b;
    layer2_outputs(3624) <= a or b;
    layer2_outputs(3625) <= a;
    layer2_outputs(3626) <= not a or b;
    layer2_outputs(3627) <= not b or a;
    layer2_outputs(3628) <= b and not a;
    layer2_outputs(3629) <= not b;
    layer2_outputs(3630) <= a and b;
    layer2_outputs(3631) <= not (a or b);
    layer2_outputs(3632) <= not (a and b);
    layer2_outputs(3633) <= not b;
    layer2_outputs(3634) <= a and not b;
    layer2_outputs(3635) <= not b or a;
    layer2_outputs(3636) <= not a;
    layer2_outputs(3637) <= not a;
    layer2_outputs(3638) <= a;
    layer2_outputs(3639) <= a;
    layer2_outputs(3640) <= b;
    layer2_outputs(3641) <= not (a or b);
    layer2_outputs(3642) <= a and b;
    layer2_outputs(3643) <= a or b;
    layer2_outputs(3644) <= not a;
    layer2_outputs(3645) <= not (a or b);
    layer2_outputs(3646) <= a;
    layer2_outputs(3647) <= a or b;
    layer2_outputs(3648) <= 1'b0;
    layer2_outputs(3649) <= a and not b;
    layer2_outputs(3650) <= 1'b1;
    layer2_outputs(3651) <= not (a and b);
    layer2_outputs(3652) <= not (a and b);
    layer2_outputs(3653) <= b;
    layer2_outputs(3654) <= a or b;
    layer2_outputs(3655) <= a xor b;
    layer2_outputs(3656) <= not a or b;
    layer2_outputs(3657) <= b;
    layer2_outputs(3658) <= a and not b;
    layer2_outputs(3659) <= a and not b;
    layer2_outputs(3660) <= b;
    layer2_outputs(3661) <= b;
    layer2_outputs(3662) <= not (a and b);
    layer2_outputs(3663) <= not (a or b);
    layer2_outputs(3664) <= a and not b;
    layer2_outputs(3665) <= not b;
    layer2_outputs(3666) <= not b;
    layer2_outputs(3667) <= not b;
    layer2_outputs(3668) <= not a;
    layer2_outputs(3669) <= a or b;
    layer2_outputs(3670) <= not (a or b);
    layer2_outputs(3671) <= not b;
    layer2_outputs(3672) <= b;
    layer2_outputs(3673) <= not b;
    layer2_outputs(3674) <= not a or b;
    layer2_outputs(3675) <= a;
    layer2_outputs(3676) <= not (a or b);
    layer2_outputs(3677) <= not (a and b);
    layer2_outputs(3678) <= a and b;
    layer2_outputs(3679) <= not a or b;
    layer2_outputs(3680) <= not a;
    layer2_outputs(3681) <= b;
    layer2_outputs(3682) <= a or b;
    layer2_outputs(3683) <= a and b;
    layer2_outputs(3684) <= a and not b;
    layer2_outputs(3685) <= b;
    layer2_outputs(3686) <= not (a xor b);
    layer2_outputs(3687) <= a or b;
    layer2_outputs(3688) <= not a;
    layer2_outputs(3689) <= not (a or b);
    layer2_outputs(3690) <= a and b;
    layer2_outputs(3691) <= not a;
    layer2_outputs(3692) <= b;
    layer2_outputs(3693) <= a;
    layer2_outputs(3694) <= not b or a;
    layer2_outputs(3695) <= a or b;
    layer2_outputs(3696) <= not a or b;
    layer2_outputs(3697) <= not a;
    layer2_outputs(3698) <= not (a or b);
    layer2_outputs(3699) <= a and not b;
    layer2_outputs(3700) <= b and not a;
    layer2_outputs(3701) <= a and b;
    layer2_outputs(3702) <= not b;
    layer2_outputs(3703) <= a or b;
    layer2_outputs(3704) <= not a;
    layer2_outputs(3705) <= a;
    layer2_outputs(3706) <= not b or a;
    layer2_outputs(3707) <= not b;
    layer2_outputs(3708) <= not a or b;
    layer2_outputs(3709) <= not (a xor b);
    layer2_outputs(3710) <= a xor b;
    layer2_outputs(3711) <= a;
    layer2_outputs(3712) <= not a;
    layer2_outputs(3713) <= not b or a;
    layer2_outputs(3714) <= a;
    layer2_outputs(3715) <= a;
    layer2_outputs(3716) <= not b;
    layer2_outputs(3717) <= a or b;
    layer2_outputs(3718) <= not (a and b);
    layer2_outputs(3719) <= a;
    layer2_outputs(3720) <= not (a or b);
    layer2_outputs(3721) <= b;
    layer2_outputs(3722) <= a and not b;
    layer2_outputs(3723) <= b;
    layer2_outputs(3724) <= not a or b;
    layer2_outputs(3725) <= 1'b1;
    layer2_outputs(3726) <= not (a or b);
    layer2_outputs(3727) <= not b;
    layer2_outputs(3728) <= not (a xor b);
    layer2_outputs(3729) <= 1'b1;
    layer2_outputs(3730) <= b and not a;
    layer2_outputs(3731) <= a and not b;
    layer2_outputs(3732) <= not a or b;
    layer2_outputs(3733) <= not a;
    layer2_outputs(3734) <= 1'b0;
    layer2_outputs(3735) <= not b;
    layer2_outputs(3736) <= not b;
    layer2_outputs(3737) <= b;
    layer2_outputs(3738) <= b;
    layer2_outputs(3739) <= b;
    layer2_outputs(3740) <= not (a and b);
    layer2_outputs(3741) <= not a;
    layer2_outputs(3742) <= b;
    layer2_outputs(3743) <= a and b;
    layer2_outputs(3744) <= a and b;
    layer2_outputs(3745) <= not b;
    layer2_outputs(3746) <= not a;
    layer2_outputs(3747) <= a xor b;
    layer2_outputs(3748) <= not a;
    layer2_outputs(3749) <= a;
    layer2_outputs(3750) <= not a or b;
    layer2_outputs(3751) <= b;
    layer2_outputs(3752) <= a;
    layer2_outputs(3753) <= a and not b;
    layer2_outputs(3754) <= not (a xor b);
    layer2_outputs(3755) <= not b;
    layer2_outputs(3756) <= not (a xor b);
    layer2_outputs(3757) <= b;
    layer2_outputs(3758) <= not (a xor b);
    layer2_outputs(3759) <= not a;
    layer2_outputs(3760) <= not a;
    layer2_outputs(3761) <= a and not b;
    layer2_outputs(3762) <= a and b;
    layer2_outputs(3763) <= not a or b;
    layer2_outputs(3764) <= not (a or b);
    layer2_outputs(3765) <= a;
    layer2_outputs(3766) <= a or b;
    layer2_outputs(3767) <= b and not a;
    layer2_outputs(3768) <= a and b;
    layer2_outputs(3769) <= b;
    layer2_outputs(3770) <= not (a xor b);
    layer2_outputs(3771) <= a xor b;
    layer2_outputs(3772) <= a or b;
    layer2_outputs(3773) <= not a or b;
    layer2_outputs(3774) <= not a;
    layer2_outputs(3775) <= not b;
    layer2_outputs(3776) <= not (a or b);
    layer2_outputs(3777) <= a xor b;
    layer2_outputs(3778) <= not a or b;
    layer2_outputs(3779) <= not a or b;
    layer2_outputs(3780) <= not b or a;
    layer2_outputs(3781) <= a or b;
    layer2_outputs(3782) <= a and b;
    layer2_outputs(3783) <= not a or b;
    layer2_outputs(3784) <= b;
    layer2_outputs(3785) <= a;
    layer2_outputs(3786) <= a and b;
    layer2_outputs(3787) <= a or b;
    layer2_outputs(3788) <= a xor b;
    layer2_outputs(3789) <= b;
    layer2_outputs(3790) <= not a;
    layer2_outputs(3791) <= not (a or b);
    layer2_outputs(3792) <= not (a and b);
    layer2_outputs(3793) <= a and not b;
    layer2_outputs(3794) <= b and not a;
    layer2_outputs(3795) <= not b;
    layer2_outputs(3796) <= not b;
    layer2_outputs(3797) <= not (a or b);
    layer2_outputs(3798) <= not b or a;
    layer2_outputs(3799) <= a xor b;
    layer2_outputs(3800) <= not b;
    layer2_outputs(3801) <= a;
    layer2_outputs(3802) <= a;
    layer2_outputs(3803) <= a xor b;
    layer2_outputs(3804) <= a;
    layer2_outputs(3805) <= a;
    layer2_outputs(3806) <= b;
    layer2_outputs(3807) <= not (a or b);
    layer2_outputs(3808) <= not b;
    layer2_outputs(3809) <= a or b;
    layer2_outputs(3810) <= 1'b0;
    layer2_outputs(3811) <= not a or b;
    layer2_outputs(3812) <= b;
    layer2_outputs(3813) <= not (a and b);
    layer2_outputs(3814) <= a and b;
    layer2_outputs(3815) <= not a;
    layer2_outputs(3816) <= not a;
    layer2_outputs(3817) <= not b or a;
    layer2_outputs(3818) <= not b;
    layer2_outputs(3819) <= b and not a;
    layer2_outputs(3820) <= not a or b;
    layer2_outputs(3821) <= b;
    layer2_outputs(3822) <= a and not b;
    layer2_outputs(3823) <= a and not b;
    layer2_outputs(3824) <= not b or a;
    layer2_outputs(3825) <= not a or b;
    layer2_outputs(3826) <= not (a and b);
    layer2_outputs(3827) <= b;
    layer2_outputs(3828) <= not b or a;
    layer2_outputs(3829) <= a and b;
    layer2_outputs(3830) <= a;
    layer2_outputs(3831) <= a or b;
    layer2_outputs(3832) <= not a or b;
    layer2_outputs(3833) <= a;
    layer2_outputs(3834) <= a and b;
    layer2_outputs(3835) <= not a;
    layer2_outputs(3836) <= not a or b;
    layer2_outputs(3837) <= not b;
    layer2_outputs(3838) <= not b;
    layer2_outputs(3839) <= not a or b;
    layer2_outputs(3840) <= not b or a;
    layer2_outputs(3841) <= a and not b;
    layer2_outputs(3842) <= a and b;
    layer2_outputs(3843) <= not (a xor b);
    layer2_outputs(3844) <= not b or a;
    layer2_outputs(3845) <= a;
    layer2_outputs(3846) <= a;
    layer2_outputs(3847) <= a and b;
    layer2_outputs(3848) <= a and not b;
    layer2_outputs(3849) <= not a;
    layer2_outputs(3850) <= not (a and b);
    layer2_outputs(3851) <= not (a xor b);
    layer2_outputs(3852) <= b;
    layer2_outputs(3853) <= b and not a;
    layer2_outputs(3854) <= a and b;
    layer2_outputs(3855) <= not (a xor b);
    layer2_outputs(3856) <= not a or b;
    layer2_outputs(3857) <= not (a xor b);
    layer2_outputs(3858) <= not b;
    layer2_outputs(3859) <= not a or b;
    layer2_outputs(3860) <= b and not a;
    layer2_outputs(3861) <= not a or b;
    layer2_outputs(3862) <= not b;
    layer2_outputs(3863) <= a or b;
    layer2_outputs(3864) <= not (a or b);
    layer2_outputs(3865) <= not a;
    layer2_outputs(3866) <= b;
    layer2_outputs(3867) <= a and not b;
    layer2_outputs(3868) <= a and b;
    layer2_outputs(3869) <= a and b;
    layer2_outputs(3870) <= not b;
    layer2_outputs(3871) <= not (a and b);
    layer2_outputs(3872) <= b and not a;
    layer2_outputs(3873) <= a and b;
    layer2_outputs(3874) <= a or b;
    layer2_outputs(3875) <= not b or a;
    layer2_outputs(3876) <= not a or b;
    layer2_outputs(3877) <= a and not b;
    layer2_outputs(3878) <= b;
    layer2_outputs(3879) <= not (a xor b);
    layer2_outputs(3880) <= not b;
    layer2_outputs(3881) <= not a;
    layer2_outputs(3882) <= a and b;
    layer2_outputs(3883) <= a and not b;
    layer2_outputs(3884) <= not a or b;
    layer2_outputs(3885) <= a;
    layer2_outputs(3886) <= not b or a;
    layer2_outputs(3887) <= not a or b;
    layer2_outputs(3888) <= a;
    layer2_outputs(3889) <= not a;
    layer2_outputs(3890) <= a and b;
    layer2_outputs(3891) <= a;
    layer2_outputs(3892) <= a and not b;
    layer2_outputs(3893) <= not b;
    layer2_outputs(3894) <= not a;
    layer2_outputs(3895) <= not b;
    layer2_outputs(3896) <= a and not b;
    layer2_outputs(3897) <= not (a and b);
    layer2_outputs(3898) <= not (a xor b);
    layer2_outputs(3899) <= not (a and b);
    layer2_outputs(3900) <= not a;
    layer2_outputs(3901) <= not (a or b);
    layer2_outputs(3902) <= a;
    layer2_outputs(3903) <= not a or b;
    layer2_outputs(3904) <= a or b;
    layer2_outputs(3905) <= a xor b;
    layer2_outputs(3906) <= a xor b;
    layer2_outputs(3907) <= a xor b;
    layer2_outputs(3908) <= not a;
    layer2_outputs(3909) <= not a;
    layer2_outputs(3910) <= b and not a;
    layer2_outputs(3911) <= b;
    layer2_outputs(3912) <= not b;
    layer2_outputs(3913) <= a and not b;
    layer2_outputs(3914) <= not (a and b);
    layer2_outputs(3915) <= not b;
    layer2_outputs(3916) <= not a or b;
    layer2_outputs(3917) <= a;
    layer2_outputs(3918) <= not (a xor b);
    layer2_outputs(3919) <= 1'b0;
    layer2_outputs(3920) <= b and not a;
    layer2_outputs(3921) <= not a;
    layer2_outputs(3922) <= a;
    layer2_outputs(3923) <= not b;
    layer2_outputs(3924) <= not b or a;
    layer2_outputs(3925) <= b;
    layer2_outputs(3926) <= not (a and b);
    layer2_outputs(3927) <= b;
    layer2_outputs(3928) <= not (a or b);
    layer2_outputs(3929) <= not a;
    layer2_outputs(3930) <= b and not a;
    layer2_outputs(3931) <= not (a or b);
    layer2_outputs(3932) <= a;
    layer2_outputs(3933) <= a or b;
    layer2_outputs(3934) <= a;
    layer2_outputs(3935) <= a and b;
    layer2_outputs(3936) <= b;
    layer2_outputs(3937) <= not (a xor b);
    layer2_outputs(3938) <= not b or a;
    layer2_outputs(3939) <= not (a xor b);
    layer2_outputs(3940) <= a and not b;
    layer2_outputs(3941) <= not a or b;
    layer2_outputs(3942) <= not b or a;
    layer2_outputs(3943) <= not (a xor b);
    layer2_outputs(3944) <= a;
    layer2_outputs(3945) <= b;
    layer2_outputs(3946) <= a and not b;
    layer2_outputs(3947) <= not a;
    layer2_outputs(3948) <= not a or b;
    layer2_outputs(3949) <= a or b;
    layer2_outputs(3950) <= a and b;
    layer2_outputs(3951) <= b;
    layer2_outputs(3952) <= not a;
    layer2_outputs(3953) <= 1'b0;
    layer2_outputs(3954) <= not a or b;
    layer2_outputs(3955) <= not (a xor b);
    layer2_outputs(3956) <= b and not a;
    layer2_outputs(3957) <= a and not b;
    layer2_outputs(3958) <= not a;
    layer2_outputs(3959) <= not (a xor b);
    layer2_outputs(3960) <= not a;
    layer2_outputs(3961) <= b;
    layer2_outputs(3962) <= not a or b;
    layer2_outputs(3963) <= not (a and b);
    layer2_outputs(3964) <= not b;
    layer2_outputs(3965) <= a and b;
    layer2_outputs(3966) <= not b or a;
    layer2_outputs(3967) <= not b or a;
    layer2_outputs(3968) <= not (a xor b);
    layer2_outputs(3969) <= a;
    layer2_outputs(3970) <= a and b;
    layer2_outputs(3971) <= not (a xor b);
    layer2_outputs(3972) <= not (a xor b);
    layer2_outputs(3973) <= a and not b;
    layer2_outputs(3974) <= not b;
    layer2_outputs(3975) <= not a;
    layer2_outputs(3976) <= not a or b;
    layer2_outputs(3977) <= not a or b;
    layer2_outputs(3978) <= a or b;
    layer2_outputs(3979) <= not (a xor b);
    layer2_outputs(3980) <= a and not b;
    layer2_outputs(3981) <= a xor b;
    layer2_outputs(3982) <= not a;
    layer2_outputs(3983) <= a;
    layer2_outputs(3984) <= b;
    layer2_outputs(3985) <= not b or a;
    layer2_outputs(3986) <= b and not a;
    layer2_outputs(3987) <= not (a or b);
    layer2_outputs(3988) <= not b or a;
    layer2_outputs(3989) <= not a;
    layer2_outputs(3990) <= a xor b;
    layer2_outputs(3991) <= not (a or b);
    layer2_outputs(3992) <= not (a or b);
    layer2_outputs(3993) <= a and b;
    layer2_outputs(3994) <= not a or b;
    layer2_outputs(3995) <= a or b;
    layer2_outputs(3996) <= not b or a;
    layer2_outputs(3997) <= a xor b;
    layer2_outputs(3998) <= b and not a;
    layer2_outputs(3999) <= a and not b;
    layer2_outputs(4000) <= 1'b0;
    layer2_outputs(4001) <= not a;
    layer2_outputs(4002) <= a and b;
    layer2_outputs(4003) <= not (a xor b);
    layer2_outputs(4004) <= not (a and b);
    layer2_outputs(4005) <= a xor b;
    layer2_outputs(4006) <= b;
    layer2_outputs(4007) <= not a;
    layer2_outputs(4008) <= a and not b;
    layer2_outputs(4009) <= not b;
    layer2_outputs(4010) <= b and not a;
    layer2_outputs(4011) <= not a or b;
    layer2_outputs(4012) <= 1'b0;
    layer2_outputs(4013) <= a or b;
    layer2_outputs(4014) <= a and not b;
    layer2_outputs(4015) <= b;
    layer2_outputs(4016) <= a;
    layer2_outputs(4017) <= b and not a;
    layer2_outputs(4018) <= a and b;
    layer2_outputs(4019) <= b;
    layer2_outputs(4020) <= not a or b;
    layer2_outputs(4021) <= not b;
    layer2_outputs(4022) <= 1'b1;
    layer2_outputs(4023) <= not (a xor b);
    layer2_outputs(4024) <= not a;
    layer2_outputs(4025) <= not a;
    layer2_outputs(4026) <= a or b;
    layer2_outputs(4027) <= b;
    layer2_outputs(4028) <= b and not a;
    layer2_outputs(4029) <= not b or a;
    layer2_outputs(4030) <= not a;
    layer2_outputs(4031) <= a or b;
    layer2_outputs(4032) <= a;
    layer2_outputs(4033) <= b and not a;
    layer2_outputs(4034) <= b and not a;
    layer2_outputs(4035) <= not (a xor b);
    layer2_outputs(4036) <= not (a xor b);
    layer2_outputs(4037) <= not (a xor b);
    layer2_outputs(4038) <= not a;
    layer2_outputs(4039) <= not a or b;
    layer2_outputs(4040) <= not b;
    layer2_outputs(4041) <= b and not a;
    layer2_outputs(4042) <= a or b;
    layer2_outputs(4043) <= a and b;
    layer2_outputs(4044) <= not (a and b);
    layer2_outputs(4045) <= not (a or b);
    layer2_outputs(4046) <= b and not a;
    layer2_outputs(4047) <= not (a xor b);
    layer2_outputs(4048) <= not a or b;
    layer2_outputs(4049) <= b;
    layer2_outputs(4050) <= not (a xor b);
    layer2_outputs(4051) <= a xor b;
    layer2_outputs(4052) <= 1'b0;
    layer2_outputs(4053) <= a;
    layer2_outputs(4054) <= b;
    layer2_outputs(4055) <= not (a and b);
    layer2_outputs(4056) <= a;
    layer2_outputs(4057) <= a or b;
    layer2_outputs(4058) <= a xor b;
    layer2_outputs(4059) <= b and not a;
    layer2_outputs(4060) <= not b or a;
    layer2_outputs(4061) <= not (a or b);
    layer2_outputs(4062) <= not (a xor b);
    layer2_outputs(4063) <= 1'b1;
    layer2_outputs(4064) <= a;
    layer2_outputs(4065) <= not a or b;
    layer2_outputs(4066) <= not (a xor b);
    layer2_outputs(4067) <= a or b;
    layer2_outputs(4068) <= a;
    layer2_outputs(4069) <= not a;
    layer2_outputs(4070) <= not (a and b);
    layer2_outputs(4071) <= not a;
    layer2_outputs(4072) <= b;
    layer2_outputs(4073) <= not (a or b);
    layer2_outputs(4074) <= not a or b;
    layer2_outputs(4075) <= b;
    layer2_outputs(4076) <= b and not a;
    layer2_outputs(4077) <= a;
    layer2_outputs(4078) <= a and b;
    layer2_outputs(4079) <= a;
    layer2_outputs(4080) <= 1'b0;
    layer2_outputs(4081) <= not a;
    layer2_outputs(4082) <= not a;
    layer2_outputs(4083) <= not a or b;
    layer2_outputs(4084) <= not a;
    layer2_outputs(4085) <= not b;
    layer2_outputs(4086) <= a xor b;
    layer2_outputs(4087) <= not a;
    layer2_outputs(4088) <= not b or a;
    layer2_outputs(4089) <= b;
    layer2_outputs(4090) <= a and not b;
    layer2_outputs(4091) <= b and not a;
    layer2_outputs(4092) <= 1'b1;
    layer2_outputs(4093) <= a;
    layer2_outputs(4094) <= not (a or b);
    layer2_outputs(4095) <= not a or b;
    layer2_outputs(4096) <= not b;
    layer2_outputs(4097) <= a and b;
    layer2_outputs(4098) <= not a or b;
    layer2_outputs(4099) <= not (a xor b);
    layer2_outputs(4100) <= not b or a;
    layer2_outputs(4101) <= b;
    layer2_outputs(4102) <= b and not a;
    layer2_outputs(4103) <= b;
    layer2_outputs(4104) <= 1'b0;
    layer2_outputs(4105) <= b;
    layer2_outputs(4106) <= not b or a;
    layer2_outputs(4107) <= not b;
    layer2_outputs(4108) <= not a;
    layer2_outputs(4109) <= not (a xor b);
    layer2_outputs(4110) <= not (a xor b);
    layer2_outputs(4111) <= b;
    layer2_outputs(4112) <= not a or b;
    layer2_outputs(4113) <= a xor b;
    layer2_outputs(4114) <= not b;
    layer2_outputs(4115) <= b and not a;
    layer2_outputs(4116) <= not b or a;
    layer2_outputs(4117) <= not (a or b);
    layer2_outputs(4118) <= b and not a;
    layer2_outputs(4119) <= a and b;
    layer2_outputs(4120) <= not b or a;
    layer2_outputs(4121) <= not a;
    layer2_outputs(4122) <= not a;
    layer2_outputs(4123) <= not a or b;
    layer2_outputs(4124) <= a;
    layer2_outputs(4125) <= not a;
    layer2_outputs(4126) <= a;
    layer2_outputs(4127) <= a;
    layer2_outputs(4128) <= b and not a;
    layer2_outputs(4129) <= not a or b;
    layer2_outputs(4130) <= a and not b;
    layer2_outputs(4131) <= a and b;
    layer2_outputs(4132) <= not (a or b);
    layer2_outputs(4133) <= not a or b;
    layer2_outputs(4134) <= b;
    layer2_outputs(4135) <= a or b;
    layer2_outputs(4136) <= b;
    layer2_outputs(4137) <= not a;
    layer2_outputs(4138) <= not b;
    layer2_outputs(4139) <= not a;
    layer2_outputs(4140) <= b and not a;
    layer2_outputs(4141) <= a;
    layer2_outputs(4142) <= not b;
    layer2_outputs(4143) <= b and not a;
    layer2_outputs(4144) <= not b or a;
    layer2_outputs(4145) <= b;
    layer2_outputs(4146) <= not b;
    layer2_outputs(4147) <= a or b;
    layer2_outputs(4148) <= a and not b;
    layer2_outputs(4149) <= a and not b;
    layer2_outputs(4150) <= not (a and b);
    layer2_outputs(4151) <= not b or a;
    layer2_outputs(4152) <= not a or b;
    layer2_outputs(4153) <= not a;
    layer2_outputs(4154) <= a or b;
    layer2_outputs(4155) <= a and not b;
    layer2_outputs(4156) <= a;
    layer2_outputs(4157) <= a and b;
    layer2_outputs(4158) <= not a;
    layer2_outputs(4159) <= a;
    layer2_outputs(4160) <= not b;
    layer2_outputs(4161) <= a and not b;
    layer2_outputs(4162) <= not (a and b);
    layer2_outputs(4163) <= b and not a;
    layer2_outputs(4164) <= a and b;
    layer2_outputs(4165) <= not (a and b);
    layer2_outputs(4166) <= not a or b;
    layer2_outputs(4167) <= not a or b;
    layer2_outputs(4168) <= a xor b;
    layer2_outputs(4169) <= a xor b;
    layer2_outputs(4170) <= not b;
    layer2_outputs(4171) <= not b;
    layer2_outputs(4172) <= not b or a;
    layer2_outputs(4173) <= b and not a;
    layer2_outputs(4174) <= not a or b;
    layer2_outputs(4175) <= not a;
    layer2_outputs(4176) <= a;
    layer2_outputs(4177) <= a;
    layer2_outputs(4178) <= not (a or b);
    layer2_outputs(4179) <= a;
    layer2_outputs(4180) <= not b;
    layer2_outputs(4181) <= not a;
    layer2_outputs(4182) <= not (a and b);
    layer2_outputs(4183) <= not b or a;
    layer2_outputs(4184) <= not (a or b);
    layer2_outputs(4185) <= not b;
    layer2_outputs(4186) <= not (a xor b);
    layer2_outputs(4187) <= not b;
    layer2_outputs(4188) <= a and b;
    layer2_outputs(4189) <= a and b;
    layer2_outputs(4190) <= a or b;
    layer2_outputs(4191) <= b;
    layer2_outputs(4192) <= not (a and b);
    layer2_outputs(4193) <= b;
    layer2_outputs(4194) <= not (a or b);
    layer2_outputs(4195) <= a or b;
    layer2_outputs(4196) <= a xor b;
    layer2_outputs(4197) <= b and not a;
    layer2_outputs(4198) <= not b or a;
    layer2_outputs(4199) <= not b;
    layer2_outputs(4200) <= a and not b;
    layer2_outputs(4201) <= a xor b;
    layer2_outputs(4202) <= a xor b;
    layer2_outputs(4203) <= b;
    layer2_outputs(4204) <= a xor b;
    layer2_outputs(4205) <= not b or a;
    layer2_outputs(4206) <= a and not b;
    layer2_outputs(4207) <= b;
    layer2_outputs(4208) <= a and b;
    layer2_outputs(4209) <= a;
    layer2_outputs(4210) <= not (a or b);
    layer2_outputs(4211) <= not b or a;
    layer2_outputs(4212) <= a and b;
    layer2_outputs(4213) <= not (a or b);
    layer2_outputs(4214) <= not a;
    layer2_outputs(4215) <= not a or b;
    layer2_outputs(4216) <= a and b;
    layer2_outputs(4217) <= a and b;
    layer2_outputs(4218) <= not (a and b);
    layer2_outputs(4219) <= b and not a;
    layer2_outputs(4220) <= a or b;
    layer2_outputs(4221) <= not (a xor b);
    layer2_outputs(4222) <= not b or a;
    layer2_outputs(4223) <= not b or a;
    layer2_outputs(4224) <= b and not a;
    layer2_outputs(4225) <= 1'b1;
    layer2_outputs(4226) <= not b;
    layer2_outputs(4227) <= not b;
    layer2_outputs(4228) <= b;
    layer2_outputs(4229) <= not b or a;
    layer2_outputs(4230) <= a;
    layer2_outputs(4231) <= b and not a;
    layer2_outputs(4232) <= b;
    layer2_outputs(4233) <= not (a xor b);
    layer2_outputs(4234) <= not b or a;
    layer2_outputs(4235) <= a or b;
    layer2_outputs(4236) <= b and not a;
    layer2_outputs(4237) <= not a or b;
    layer2_outputs(4238) <= a xor b;
    layer2_outputs(4239) <= b and not a;
    layer2_outputs(4240) <= a;
    layer2_outputs(4241) <= a or b;
    layer2_outputs(4242) <= not a;
    layer2_outputs(4243) <= a;
    layer2_outputs(4244) <= not b;
    layer2_outputs(4245) <= a xor b;
    layer2_outputs(4246) <= a;
    layer2_outputs(4247) <= a or b;
    layer2_outputs(4248) <= not b or a;
    layer2_outputs(4249) <= a;
    layer2_outputs(4250) <= b and not a;
    layer2_outputs(4251) <= b;
    layer2_outputs(4252) <= b;
    layer2_outputs(4253) <= a;
    layer2_outputs(4254) <= a and not b;
    layer2_outputs(4255) <= not a or b;
    layer2_outputs(4256) <= not (a and b);
    layer2_outputs(4257) <= not (a and b);
    layer2_outputs(4258) <= not a or b;
    layer2_outputs(4259) <= a and not b;
    layer2_outputs(4260) <= a and b;
    layer2_outputs(4261) <= not a;
    layer2_outputs(4262) <= a or b;
    layer2_outputs(4263) <= not (a and b);
    layer2_outputs(4264) <= b;
    layer2_outputs(4265) <= not b or a;
    layer2_outputs(4266) <= not a;
    layer2_outputs(4267) <= not b or a;
    layer2_outputs(4268) <= not (a or b);
    layer2_outputs(4269) <= not (a xor b);
    layer2_outputs(4270) <= a and b;
    layer2_outputs(4271) <= b and not a;
    layer2_outputs(4272) <= b;
    layer2_outputs(4273) <= b;
    layer2_outputs(4274) <= b;
    layer2_outputs(4275) <= not b;
    layer2_outputs(4276) <= 1'b0;
    layer2_outputs(4277) <= not a;
    layer2_outputs(4278) <= not (a and b);
    layer2_outputs(4279) <= not b;
    layer2_outputs(4280) <= 1'b0;
    layer2_outputs(4281) <= not b;
    layer2_outputs(4282) <= a;
    layer2_outputs(4283) <= not a;
    layer2_outputs(4284) <= not b;
    layer2_outputs(4285) <= not b or a;
    layer2_outputs(4286) <= a and not b;
    layer2_outputs(4287) <= not b;
    layer2_outputs(4288) <= 1'b0;
    layer2_outputs(4289) <= not b;
    layer2_outputs(4290) <= not (a and b);
    layer2_outputs(4291) <= b;
    layer2_outputs(4292) <= b;
    layer2_outputs(4293) <= not a;
    layer2_outputs(4294) <= b and not a;
    layer2_outputs(4295) <= not b or a;
    layer2_outputs(4296) <= a;
    layer2_outputs(4297) <= a and not b;
    layer2_outputs(4298) <= not (a or b);
    layer2_outputs(4299) <= not b;
    layer2_outputs(4300) <= 1'b1;
    layer2_outputs(4301) <= not a;
    layer2_outputs(4302) <= b and not a;
    layer2_outputs(4303) <= a;
    layer2_outputs(4304) <= a or b;
    layer2_outputs(4305) <= a;
    layer2_outputs(4306) <= not a or b;
    layer2_outputs(4307) <= a and b;
    layer2_outputs(4308) <= not a;
    layer2_outputs(4309) <= not (a or b);
    layer2_outputs(4310) <= not a;
    layer2_outputs(4311) <= b;
    layer2_outputs(4312) <= 1'b1;
    layer2_outputs(4313) <= not (a or b);
    layer2_outputs(4314) <= not (a and b);
    layer2_outputs(4315) <= 1'b1;
    layer2_outputs(4316) <= b and not a;
    layer2_outputs(4317) <= a and b;
    layer2_outputs(4318) <= a and not b;
    layer2_outputs(4319) <= a and not b;
    layer2_outputs(4320) <= not a or b;
    layer2_outputs(4321) <= b and not a;
    layer2_outputs(4322) <= a xor b;
    layer2_outputs(4323) <= not (a and b);
    layer2_outputs(4324) <= not b or a;
    layer2_outputs(4325) <= a xor b;
    layer2_outputs(4326) <= not (a or b);
    layer2_outputs(4327) <= b and not a;
    layer2_outputs(4328) <= b;
    layer2_outputs(4329) <= 1'b1;
    layer2_outputs(4330) <= a and not b;
    layer2_outputs(4331) <= a or b;
    layer2_outputs(4332) <= a;
    layer2_outputs(4333) <= a or b;
    layer2_outputs(4334) <= a or b;
    layer2_outputs(4335) <= not (a or b);
    layer2_outputs(4336) <= not b;
    layer2_outputs(4337) <= not a;
    layer2_outputs(4338) <= a and b;
    layer2_outputs(4339) <= b and not a;
    layer2_outputs(4340) <= not a;
    layer2_outputs(4341) <= a and not b;
    layer2_outputs(4342) <= not (a and b);
    layer2_outputs(4343) <= not b;
    layer2_outputs(4344) <= a;
    layer2_outputs(4345) <= a;
    layer2_outputs(4346) <= not b;
    layer2_outputs(4347) <= not (a or b);
    layer2_outputs(4348) <= a or b;
    layer2_outputs(4349) <= not (a and b);
    layer2_outputs(4350) <= not (a and b);
    layer2_outputs(4351) <= a;
    layer2_outputs(4352) <= not a;
    layer2_outputs(4353) <= not a;
    layer2_outputs(4354) <= a;
    layer2_outputs(4355) <= 1'b1;
    layer2_outputs(4356) <= a and not b;
    layer2_outputs(4357) <= not (a xor b);
    layer2_outputs(4358) <= not a or b;
    layer2_outputs(4359) <= a and not b;
    layer2_outputs(4360) <= a;
    layer2_outputs(4361) <= a xor b;
    layer2_outputs(4362) <= not a or b;
    layer2_outputs(4363) <= a and not b;
    layer2_outputs(4364) <= a;
    layer2_outputs(4365) <= not a;
    layer2_outputs(4366) <= a or b;
    layer2_outputs(4367) <= b;
    layer2_outputs(4368) <= not a;
    layer2_outputs(4369) <= not a;
    layer2_outputs(4370) <= not b or a;
    layer2_outputs(4371) <= a xor b;
    layer2_outputs(4372) <= not (a or b);
    layer2_outputs(4373) <= not (a or b);
    layer2_outputs(4374) <= not (a and b);
    layer2_outputs(4375) <= not a;
    layer2_outputs(4376) <= b;
    layer2_outputs(4377) <= not a;
    layer2_outputs(4378) <= not b or a;
    layer2_outputs(4379) <= b;
    layer2_outputs(4380) <= not (a and b);
    layer2_outputs(4381) <= b and not a;
    layer2_outputs(4382) <= not (a and b);
    layer2_outputs(4383) <= a and not b;
    layer2_outputs(4384) <= a;
    layer2_outputs(4385) <= 1'b0;
    layer2_outputs(4386) <= b;
    layer2_outputs(4387) <= b;
    layer2_outputs(4388) <= a and not b;
    layer2_outputs(4389) <= b and not a;
    layer2_outputs(4390) <= not b;
    layer2_outputs(4391) <= not a or b;
    layer2_outputs(4392) <= not a or b;
    layer2_outputs(4393) <= not a;
    layer2_outputs(4394) <= not a or b;
    layer2_outputs(4395) <= a or b;
    layer2_outputs(4396) <= not b;
    layer2_outputs(4397) <= a or b;
    layer2_outputs(4398) <= not (a or b);
    layer2_outputs(4399) <= a or b;
    layer2_outputs(4400) <= not b;
    layer2_outputs(4401) <= 1'b1;
    layer2_outputs(4402) <= b;
    layer2_outputs(4403) <= not b or a;
    layer2_outputs(4404) <= a;
    layer2_outputs(4405) <= not a;
    layer2_outputs(4406) <= b and not a;
    layer2_outputs(4407) <= not a;
    layer2_outputs(4408) <= a or b;
    layer2_outputs(4409) <= a and b;
    layer2_outputs(4410) <= a or b;
    layer2_outputs(4411) <= not b;
    layer2_outputs(4412) <= a;
    layer2_outputs(4413) <= not a;
    layer2_outputs(4414) <= a or b;
    layer2_outputs(4415) <= a or b;
    layer2_outputs(4416) <= not b or a;
    layer2_outputs(4417) <= b and not a;
    layer2_outputs(4418) <= not b;
    layer2_outputs(4419) <= not a;
    layer2_outputs(4420) <= not a;
    layer2_outputs(4421) <= a or b;
    layer2_outputs(4422) <= not b or a;
    layer2_outputs(4423) <= not (a or b);
    layer2_outputs(4424) <= not (a xor b);
    layer2_outputs(4425) <= not b or a;
    layer2_outputs(4426) <= not a;
    layer2_outputs(4427) <= a;
    layer2_outputs(4428) <= not (a xor b);
    layer2_outputs(4429) <= a xor b;
    layer2_outputs(4430) <= a or b;
    layer2_outputs(4431) <= a;
    layer2_outputs(4432) <= b and not a;
    layer2_outputs(4433) <= b;
    layer2_outputs(4434) <= not (a and b);
    layer2_outputs(4435) <= a xor b;
    layer2_outputs(4436) <= a and b;
    layer2_outputs(4437) <= not a or b;
    layer2_outputs(4438) <= b;
    layer2_outputs(4439) <= a or b;
    layer2_outputs(4440) <= b and not a;
    layer2_outputs(4441) <= a;
    layer2_outputs(4442) <= not b;
    layer2_outputs(4443) <= b and not a;
    layer2_outputs(4444) <= a;
    layer2_outputs(4445) <= a and b;
    layer2_outputs(4446) <= b;
    layer2_outputs(4447) <= not b;
    layer2_outputs(4448) <= a and not b;
    layer2_outputs(4449) <= not (a and b);
    layer2_outputs(4450) <= not b;
    layer2_outputs(4451) <= not b or a;
    layer2_outputs(4452) <= b and not a;
    layer2_outputs(4453) <= not (a xor b);
    layer2_outputs(4454) <= not (a or b);
    layer2_outputs(4455) <= a or b;
    layer2_outputs(4456) <= a;
    layer2_outputs(4457) <= not b;
    layer2_outputs(4458) <= b and not a;
    layer2_outputs(4459) <= not (a or b);
    layer2_outputs(4460) <= not (a and b);
    layer2_outputs(4461) <= a and not b;
    layer2_outputs(4462) <= not (a or b);
    layer2_outputs(4463) <= a and not b;
    layer2_outputs(4464) <= b;
    layer2_outputs(4465) <= not (a or b);
    layer2_outputs(4466) <= not (a or b);
    layer2_outputs(4467) <= b;
    layer2_outputs(4468) <= a or b;
    layer2_outputs(4469) <= not (a and b);
    layer2_outputs(4470) <= not (a xor b);
    layer2_outputs(4471) <= a and b;
    layer2_outputs(4472) <= not a or b;
    layer2_outputs(4473) <= a xor b;
    layer2_outputs(4474) <= not (a xor b);
    layer2_outputs(4475) <= not b;
    layer2_outputs(4476) <= b and not a;
    layer2_outputs(4477) <= a or b;
    layer2_outputs(4478) <= a and not b;
    layer2_outputs(4479) <= a xor b;
    layer2_outputs(4480) <= not a;
    layer2_outputs(4481) <= b and not a;
    layer2_outputs(4482) <= not (a xor b);
    layer2_outputs(4483) <= a and b;
    layer2_outputs(4484) <= not a or b;
    layer2_outputs(4485) <= a;
    layer2_outputs(4486) <= a;
    layer2_outputs(4487) <= not (a or b);
    layer2_outputs(4488) <= not b;
    layer2_outputs(4489) <= a and not b;
    layer2_outputs(4490) <= 1'b1;
    layer2_outputs(4491) <= not b or a;
    layer2_outputs(4492) <= a xor b;
    layer2_outputs(4493) <= not (a or b);
    layer2_outputs(4494) <= not a;
    layer2_outputs(4495) <= not (a or b);
    layer2_outputs(4496) <= not (a xor b);
    layer2_outputs(4497) <= not (a or b);
    layer2_outputs(4498) <= not a;
    layer2_outputs(4499) <= a and not b;
    layer2_outputs(4500) <= a;
    layer2_outputs(4501) <= not (a and b);
    layer2_outputs(4502) <= b;
    layer2_outputs(4503) <= not a;
    layer2_outputs(4504) <= a;
    layer2_outputs(4505) <= not b;
    layer2_outputs(4506) <= not (a or b);
    layer2_outputs(4507) <= not b or a;
    layer2_outputs(4508) <= not b;
    layer2_outputs(4509) <= not (a xor b);
    layer2_outputs(4510) <= a;
    layer2_outputs(4511) <= a and not b;
    layer2_outputs(4512) <= not a;
    layer2_outputs(4513) <= not b or a;
    layer2_outputs(4514) <= a and not b;
    layer2_outputs(4515) <= not a or b;
    layer2_outputs(4516) <= b and not a;
    layer2_outputs(4517) <= not (a and b);
    layer2_outputs(4518) <= b;
    layer2_outputs(4519) <= a or b;
    layer2_outputs(4520) <= b and not a;
    layer2_outputs(4521) <= a and not b;
    layer2_outputs(4522) <= a and not b;
    layer2_outputs(4523) <= not b;
    layer2_outputs(4524) <= not b;
    layer2_outputs(4525) <= not b or a;
    layer2_outputs(4526) <= 1'b1;
    layer2_outputs(4527) <= not b or a;
    layer2_outputs(4528) <= a and not b;
    layer2_outputs(4529) <= a and b;
    layer2_outputs(4530) <= a or b;
    layer2_outputs(4531) <= not (a and b);
    layer2_outputs(4532) <= 1'b0;
    layer2_outputs(4533) <= b;
    layer2_outputs(4534) <= a and not b;
    layer2_outputs(4535) <= not (a or b);
    layer2_outputs(4536) <= a xor b;
    layer2_outputs(4537) <= 1'b0;
    layer2_outputs(4538) <= not a or b;
    layer2_outputs(4539) <= not (a and b);
    layer2_outputs(4540) <= b;
    layer2_outputs(4541) <= b;
    layer2_outputs(4542) <= b;
    layer2_outputs(4543) <= b;
    layer2_outputs(4544) <= b;
    layer2_outputs(4545) <= not b;
    layer2_outputs(4546) <= a xor b;
    layer2_outputs(4547) <= not a;
    layer2_outputs(4548) <= a;
    layer2_outputs(4549) <= a and not b;
    layer2_outputs(4550) <= not (a or b);
    layer2_outputs(4551) <= not (a xor b);
    layer2_outputs(4552) <= a and not b;
    layer2_outputs(4553) <= a;
    layer2_outputs(4554) <= not (a or b);
    layer2_outputs(4555) <= not b;
    layer2_outputs(4556) <= not b;
    layer2_outputs(4557) <= a or b;
    layer2_outputs(4558) <= not a;
    layer2_outputs(4559) <= a or b;
    layer2_outputs(4560) <= not b or a;
    layer2_outputs(4561) <= b and not a;
    layer2_outputs(4562) <= b;
    layer2_outputs(4563) <= not a or b;
    layer2_outputs(4564) <= b;
    layer2_outputs(4565) <= not a;
    layer2_outputs(4566) <= b and not a;
    layer2_outputs(4567) <= a and not b;
    layer2_outputs(4568) <= not (a xor b);
    layer2_outputs(4569) <= b;
    layer2_outputs(4570) <= b;
    layer2_outputs(4571) <= b;
    layer2_outputs(4572) <= not a;
    layer2_outputs(4573) <= a or b;
    layer2_outputs(4574) <= not a or b;
    layer2_outputs(4575) <= a or b;
    layer2_outputs(4576) <= not a;
    layer2_outputs(4577) <= not b or a;
    layer2_outputs(4578) <= a or b;
    layer2_outputs(4579) <= a;
    layer2_outputs(4580) <= a and b;
    layer2_outputs(4581) <= not (a and b);
    layer2_outputs(4582) <= not a or b;
    layer2_outputs(4583) <= a and not b;
    layer2_outputs(4584) <= not a;
    layer2_outputs(4585) <= a;
    layer2_outputs(4586) <= 1'b0;
    layer2_outputs(4587) <= not a;
    layer2_outputs(4588) <= b;
    layer2_outputs(4589) <= a and not b;
    layer2_outputs(4590) <= not a or b;
    layer2_outputs(4591) <= b;
    layer2_outputs(4592) <= b;
    layer2_outputs(4593) <= b;
    layer2_outputs(4594) <= a;
    layer2_outputs(4595) <= not b or a;
    layer2_outputs(4596) <= b;
    layer2_outputs(4597) <= not b;
    layer2_outputs(4598) <= not a;
    layer2_outputs(4599) <= a and b;
    layer2_outputs(4600) <= b and not a;
    layer2_outputs(4601) <= a;
    layer2_outputs(4602) <= b and not a;
    layer2_outputs(4603) <= a and not b;
    layer2_outputs(4604) <= a and not b;
    layer2_outputs(4605) <= not a;
    layer2_outputs(4606) <= a;
    layer2_outputs(4607) <= b;
    layer2_outputs(4608) <= not b or a;
    layer2_outputs(4609) <= a;
    layer2_outputs(4610) <= not a;
    layer2_outputs(4611) <= b;
    layer2_outputs(4612) <= not a or b;
    layer2_outputs(4613) <= not a;
    layer2_outputs(4614) <= 1'b1;
    layer2_outputs(4615) <= a xor b;
    layer2_outputs(4616) <= a and not b;
    layer2_outputs(4617) <= a xor b;
    layer2_outputs(4618) <= not (a xor b);
    layer2_outputs(4619) <= a xor b;
    layer2_outputs(4620) <= not (a or b);
    layer2_outputs(4621) <= a;
    layer2_outputs(4622) <= not a;
    layer2_outputs(4623) <= a or b;
    layer2_outputs(4624) <= not a;
    layer2_outputs(4625) <= b;
    layer2_outputs(4626) <= b;
    layer2_outputs(4627) <= not a or b;
    layer2_outputs(4628) <= b;
    layer2_outputs(4629) <= a;
    layer2_outputs(4630) <= b and not a;
    layer2_outputs(4631) <= not b;
    layer2_outputs(4632) <= not (a xor b);
    layer2_outputs(4633) <= not (a or b);
    layer2_outputs(4634) <= a and not b;
    layer2_outputs(4635) <= not a or b;
    layer2_outputs(4636) <= 1'b0;
    layer2_outputs(4637) <= b;
    layer2_outputs(4638) <= not (a xor b);
    layer2_outputs(4639) <= not b;
    layer2_outputs(4640) <= b;
    layer2_outputs(4641) <= not a or b;
    layer2_outputs(4642) <= b and not a;
    layer2_outputs(4643) <= a and b;
    layer2_outputs(4644) <= b;
    layer2_outputs(4645) <= b and not a;
    layer2_outputs(4646) <= not (a and b);
    layer2_outputs(4647) <= not (a or b);
    layer2_outputs(4648) <= a or b;
    layer2_outputs(4649) <= not b or a;
    layer2_outputs(4650) <= not (a and b);
    layer2_outputs(4651) <= not a;
    layer2_outputs(4652) <= not a or b;
    layer2_outputs(4653) <= not (a or b);
    layer2_outputs(4654) <= a and not b;
    layer2_outputs(4655) <= a xor b;
    layer2_outputs(4656) <= 1'b1;
    layer2_outputs(4657) <= a;
    layer2_outputs(4658) <= a and b;
    layer2_outputs(4659) <= not b;
    layer2_outputs(4660) <= not (a xor b);
    layer2_outputs(4661) <= b and not a;
    layer2_outputs(4662) <= a;
    layer2_outputs(4663) <= b;
    layer2_outputs(4664) <= b;
    layer2_outputs(4665) <= a and not b;
    layer2_outputs(4666) <= a;
    layer2_outputs(4667) <= not b or a;
    layer2_outputs(4668) <= not (a and b);
    layer2_outputs(4669) <= b and not a;
    layer2_outputs(4670) <= not (a and b);
    layer2_outputs(4671) <= not a or b;
    layer2_outputs(4672) <= not (a and b);
    layer2_outputs(4673) <= 1'b0;
    layer2_outputs(4674) <= not b;
    layer2_outputs(4675) <= not b or a;
    layer2_outputs(4676) <= not (a or b);
    layer2_outputs(4677) <= a and not b;
    layer2_outputs(4678) <= not (a or b);
    layer2_outputs(4679) <= not a;
    layer2_outputs(4680) <= a;
    layer2_outputs(4681) <= not b;
    layer2_outputs(4682) <= not a or b;
    layer2_outputs(4683) <= a and not b;
    layer2_outputs(4684) <= a and not b;
    layer2_outputs(4685) <= a and not b;
    layer2_outputs(4686) <= not a;
    layer2_outputs(4687) <= not b or a;
    layer2_outputs(4688) <= a and b;
    layer2_outputs(4689) <= not b;
    layer2_outputs(4690) <= a and not b;
    layer2_outputs(4691) <= a;
    layer2_outputs(4692) <= not a;
    layer2_outputs(4693) <= b;
    layer2_outputs(4694) <= not (a and b);
    layer2_outputs(4695) <= a;
    layer2_outputs(4696) <= not b;
    layer2_outputs(4697) <= a xor b;
    layer2_outputs(4698) <= not (a or b);
    layer2_outputs(4699) <= a xor b;
    layer2_outputs(4700) <= not b;
    layer2_outputs(4701) <= a xor b;
    layer2_outputs(4702) <= b;
    layer2_outputs(4703) <= not a;
    layer2_outputs(4704) <= a or b;
    layer2_outputs(4705) <= not a;
    layer2_outputs(4706) <= not b;
    layer2_outputs(4707) <= not a;
    layer2_outputs(4708) <= a or b;
    layer2_outputs(4709) <= b and not a;
    layer2_outputs(4710) <= not a or b;
    layer2_outputs(4711) <= b and not a;
    layer2_outputs(4712) <= a;
    layer2_outputs(4713) <= b;
    layer2_outputs(4714) <= not a;
    layer2_outputs(4715) <= b and not a;
    layer2_outputs(4716) <= a;
    layer2_outputs(4717) <= not b or a;
    layer2_outputs(4718) <= b;
    layer2_outputs(4719) <= not b;
    layer2_outputs(4720) <= not a;
    layer2_outputs(4721) <= not b;
    layer2_outputs(4722) <= b;
    layer2_outputs(4723) <= not a;
    layer2_outputs(4724) <= not a or b;
    layer2_outputs(4725) <= not b;
    layer2_outputs(4726) <= not b or a;
    layer2_outputs(4727) <= not b;
    layer2_outputs(4728) <= b and not a;
    layer2_outputs(4729) <= a;
    layer2_outputs(4730) <= a;
    layer2_outputs(4731) <= 1'b0;
    layer2_outputs(4732) <= not a;
    layer2_outputs(4733) <= a or b;
    layer2_outputs(4734) <= not b;
    layer2_outputs(4735) <= not a;
    layer2_outputs(4736) <= b;
    layer2_outputs(4737) <= not a or b;
    layer2_outputs(4738) <= not (a and b);
    layer2_outputs(4739) <= not b;
    layer2_outputs(4740) <= 1'b1;
    layer2_outputs(4741) <= b;
    layer2_outputs(4742) <= not a;
    layer2_outputs(4743) <= a or b;
    layer2_outputs(4744) <= a or b;
    layer2_outputs(4745) <= 1'b1;
    layer2_outputs(4746) <= a and not b;
    layer2_outputs(4747) <= not b;
    layer2_outputs(4748) <= b;
    layer2_outputs(4749) <= a xor b;
    layer2_outputs(4750) <= not b or a;
    layer2_outputs(4751) <= b;
    layer2_outputs(4752) <= not a;
    layer2_outputs(4753) <= not a;
    layer2_outputs(4754) <= a;
    layer2_outputs(4755) <= a or b;
    layer2_outputs(4756) <= not a or b;
    layer2_outputs(4757) <= a or b;
    layer2_outputs(4758) <= a xor b;
    layer2_outputs(4759) <= not (a xor b);
    layer2_outputs(4760) <= not (a and b);
    layer2_outputs(4761) <= not b or a;
    layer2_outputs(4762) <= not (a or b);
    layer2_outputs(4763) <= b;
    layer2_outputs(4764) <= not (a or b);
    layer2_outputs(4765) <= b;
    layer2_outputs(4766) <= 1'b0;
    layer2_outputs(4767) <= a and not b;
    layer2_outputs(4768) <= not (a or b);
    layer2_outputs(4769) <= a;
    layer2_outputs(4770) <= a and not b;
    layer2_outputs(4771) <= b;
    layer2_outputs(4772) <= b;
    layer2_outputs(4773) <= a;
    layer2_outputs(4774) <= not (a and b);
    layer2_outputs(4775) <= not b or a;
    layer2_outputs(4776) <= not (a or b);
    layer2_outputs(4777) <= a or b;
    layer2_outputs(4778) <= b;
    layer2_outputs(4779) <= not b or a;
    layer2_outputs(4780) <= not (a and b);
    layer2_outputs(4781) <= b;
    layer2_outputs(4782) <= a xor b;
    layer2_outputs(4783) <= a and not b;
    layer2_outputs(4784) <= a and b;
    layer2_outputs(4785) <= not (a or b);
    layer2_outputs(4786) <= b;
    layer2_outputs(4787) <= a or b;
    layer2_outputs(4788) <= not (a xor b);
    layer2_outputs(4789) <= b and not a;
    layer2_outputs(4790) <= not a or b;
    layer2_outputs(4791) <= not (a and b);
    layer2_outputs(4792) <= not (a or b);
    layer2_outputs(4793) <= not a or b;
    layer2_outputs(4794) <= not a or b;
    layer2_outputs(4795) <= 1'b1;
    layer2_outputs(4796) <= a;
    layer2_outputs(4797) <= 1'b0;
    layer2_outputs(4798) <= not (a xor b);
    layer2_outputs(4799) <= not (a xor b);
    layer2_outputs(4800) <= a;
    layer2_outputs(4801) <= a;
    layer2_outputs(4802) <= not (a xor b);
    layer2_outputs(4803) <= not b;
    layer2_outputs(4804) <= a;
    layer2_outputs(4805) <= b and not a;
    layer2_outputs(4806) <= a or b;
    layer2_outputs(4807) <= not (a and b);
    layer2_outputs(4808) <= a and b;
    layer2_outputs(4809) <= not b;
    layer2_outputs(4810) <= b;
    layer2_outputs(4811) <= not a;
    layer2_outputs(4812) <= a or b;
    layer2_outputs(4813) <= b;
    layer2_outputs(4814) <= b;
    layer2_outputs(4815) <= b and not a;
    layer2_outputs(4816) <= not b or a;
    layer2_outputs(4817) <= b;
    layer2_outputs(4818) <= a or b;
    layer2_outputs(4819) <= not a;
    layer2_outputs(4820) <= not a or b;
    layer2_outputs(4821) <= not (a xor b);
    layer2_outputs(4822) <= a;
    layer2_outputs(4823) <= not (a or b);
    layer2_outputs(4824) <= a;
    layer2_outputs(4825) <= b and not a;
    layer2_outputs(4826) <= not b;
    layer2_outputs(4827) <= not a or b;
    layer2_outputs(4828) <= not (a and b);
    layer2_outputs(4829) <= a;
    layer2_outputs(4830) <= a;
    layer2_outputs(4831) <= a and b;
    layer2_outputs(4832) <= not a;
    layer2_outputs(4833) <= not a or b;
    layer2_outputs(4834) <= a and b;
    layer2_outputs(4835) <= not a;
    layer2_outputs(4836) <= a and b;
    layer2_outputs(4837) <= a and not b;
    layer2_outputs(4838) <= not a or b;
    layer2_outputs(4839) <= not b;
    layer2_outputs(4840) <= a and b;
    layer2_outputs(4841) <= a or b;
    layer2_outputs(4842) <= a;
    layer2_outputs(4843) <= not a;
    layer2_outputs(4844) <= not b or a;
    layer2_outputs(4845) <= b;
    layer2_outputs(4846) <= b;
    layer2_outputs(4847) <= not a;
    layer2_outputs(4848) <= not b or a;
    layer2_outputs(4849) <= not (a and b);
    layer2_outputs(4850) <= b;
    layer2_outputs(4851) <= b;
    layer2_outputs(4852) <= not b;
    layer2_outputs(4853) <= not b;
    layer2_outputs(4854) <= not b or a;
    layer2_outputs(4855) <= a and not b;
    layer2_outputs(4856) <= not b or a;
    layer2_outputs(4857) <= not b;
    layer2_outputs(4858) <= not a;
    layer2_outputs(4859) <= a and not b;
    layer2_outputs(4860) <= not b;
    layer2_outputs(4861) <= b;
    layer2_outputs(4862) <= a and not b;
    layer2_outputs(4863) <= not a;
    layer2_outputs(4864) <= a and b;
    layer2_outputs(4865) <= a xor b;
    layer2_outputs(4866) <= not (a xor b);
    layer2_outputs(4867) <= not (a or b);
    layer2_outputs(4868) <= a and not b;
    layer2_outputs(4869) <= not (a xor b);
    layer2_outputs(4870) <= a;
    layer2_outputs(4871) <= not b;
    layer2_outputs(4872) <= not b or a;
    layer2_outputs(4873) <= a and not b;
    layer2_outputs(4874) <= not b;
    layer2_outputs(4875) <= not b;
    layer2_outputs(4876) <= not b;
    layer2_outputs(4877) <= not b;
    layer2_outputs(4878) <= a and b;
    layer2_outputs(4879) <= not (a or b);
    layer2_outputs(4880) <= a or b;
    layer2_outputs(4881) <= b;
    layer2_outputs(4882) <= not (a and b);
    layer2_outputs(4883) <= 1'b0;
    layer2_outputs(4884) <= a;
    layer2_outputs(4885) <= b;
    layer2_outputs(4886) <= not (a or b);
    layer2_outputs(4887) <= not b or a;
    layer2_outputs(4888) <= not a;
    layer2_outputs(4889) <= not a;
    layer2_outputs(4890) <= a xor b;
    layer2_outputs(4891) <= not a or b;
    layer2_outputs(4892) <= b and not a;
    layer2_outputs(4893) <= a and b;
    layer2_outputs(4894) <= a;
    layer2_outputs(4895) <= b and not a;
    layer2_outputs(4896) <= a and b;
    layer2_outputs(4897) <= b and not a;
    layer2_outputs(4898) <= not a;
    layer2_outputs(4899) <= not (a xor b);
    layer2_outputs(4900) <= not a;
    layer2_outputs(4901) <= not (a xor b);
    layer2_outputs(4902) <= a xor b;
    layer2_outputs(4903) <= not a or b;
    layer2_outputs(4904) <= b;
    layer2_outputs(4905) <= a and not b;
    layer2_outputs(4906) <= a or b;
    layer2_outputs(4907) <= b and not a;
    layer2_outputs(4908) <= a or b;
    layer2_outputs(4909) <= not (a and b);
    layer2_outputs(4910) <= 1'b0;
    layer2_outputs(4911) <= a and b;
    layer2_outputs(4912) <= not (a xor b);
    layer2_outputs(4913) <= b and not a;
    layer2_outputs(4914) <= not (a xor b);
    layer2_outputs(4915) <= a and not b;
    layer2_outputs(4916) <= a or b;
    layer2_outputs(4917) <= a xor b;
    layer2_outputs(4918) <= not b;
    layer2_outputs(4919) <= not a;
    layer2_outputs(4920) <= not (a or b);
    layer2_outputs(4921) <= a;
    layer2_outputs(4922) <= not a or b;
    layer2_outputs(4923) <= not b;
    layer2_outputs(4924) <= not b or a;
    layer2_outputs(4925) <= not a;
    layer2_outputs(4926) <= not (a xor b);
    layer2_outputs(4927) <= a or b;
    layer2_outputs(4928) <= not a;
    layer2_outputs(4929) <= b;
    layer2_outputs(4930) <= a;
    layer2_outputs(4931) <= not (a and b);
    layer2_outputs(4932) <= not a;
    layer2_outputs(4933) <= not (a or b);
    layer2_outputs(4934) <= b;
    layer2_outputs(4935) <= not a or b;
    layer2_outputs(4936) <= not (a and b);
    layer2_outputs(4937) <= a;
    layer2_outputs(4938) <= not b;
    layer2_outputs(4939) <= a and not b;
    layer2_outputs(4940) <= a and not b;
    layer2_outputs(4941) <= a;
    layer2_outputs(4942) <= not (a xor b);
    layer2_outputs(4943) <= a and not b;
    layer2_outputs(4944) <= not b or a;
    layer2_outputs(4945) <= a and b;
    layer2_outputs(4946) <= b;
    layer2_outputs(4947) <= not b or a;
    layer2_outputs(4948) <= not a or b;
    layer2_outputs(4949) <= b and not a;
    layer2_outputs(4950) <= b and not a;
    layer2_outputs(4951) <= not (a and b);
    layer2_outputs(4952) <= b;
    layer2_outputs(4953) <= a or b;
    layer2_outputs(4954) <= 1'b1;
    layer2_outputs(4955) <= a and not b;
    layer2_outputs(4956) <= not (a xor b);
    layer2_outputs(4957) <= a or b;
    layer2_outputs(4958) <= not a or b;
    layer2_outputs(4959) <= a and not b;
    layer2_outputs(4960) <= not a;
    layer2_outputs(4961) <= not a;
    layer2_outputs(4962) <= not (a or b);
    layer2_outputs(4963) <= not (a xor b);
    layer2_outputs(4964) <= not b;
    layer2_outputs(4965) <= not a;
    layer2_outputs(4966) <= b;
    layer2_outputs(4967) <= a and b;
    layer2_outputs(4968) <= not b;
    layer2_outputs(4969) <= not a;
    layer2_outputs(4970) <= not b;
    layer2_outputs(4971) <= not (a and b);
    layer2_outputs(4972) <= a;
    layer2_outputs(4973) <= not b or a;
    layer2_outputs(4974) <= b and not a;
    layer2_outputs(4975) <= 1'b0;
    layer2_outputs(4976) <= not b or a;
    layer2_outputs(4977) <= not (a xor b);
    layer2_outputs(4978) <= a and not b;
    layer2_outputs(4979) <= not b;
    layer2_outputs(4980) <= a and b;
    layer2_outputs(4981) <= not b;
    layer2_outputs(4982) <= 1'b0;
    layer2_outputs(4983) <= not (a or b);
    layer2_outputs(4984) <= a and b;
    layer2_outputs(4985) <= not a or b;
    layer2_outputs(4986) <= not (a and b);
    layer2_outputs(4987) <= b;
    layer2_outputs(4988) <= not a;
    layer2_outputs(4989) <= a or b;
    layer2_outputs(4990) <= 1'b0;
    layer2_outputs(4991) <= a and b;
    layer2_outputs(4992) <= not a or b;
    layer2_outputs(4993) <= not b;
    layer2_outputs(4994) <= not (a and b);
    layer2_outputs(4995) <= not (a and b);
    layer2_outputs(4996) <= not b;
    layer2_outputs(4997) <= a;
    layer2_outputs(4998) <= a;
    layer2_outputs(4999) <= b and not a;
    layer2_outputs(5000) <= not (a or b);
    layer2_outputs(5001) <= not a;
    layer2_outputs(5002) <= not a or b;
    layer2_outputs(5003) <= a and not b;
    layer2_outputs(5004) <= a;
    layer2_outputs(5005) <= b and not a;
    layer2_outputs(5006) <= not b;
    layer2_outputs(5007) <= a;
    layer2_outputs(5008) <= not b;
    layer2_outputs(5009) <= a and not b;
    layer2_outputs(5010) <= not a;
    layer2_outputs(5011) <= not a;
    layer2_outputs(5012) <= not b;
    layer2_outputs(5013) <= not b;
    layer2_outputs(5014) <= not a or b;
    layer2_outputs(5015) <= not (a or b);
    layer2_outputs(5016) <= b and not a;
    layer2_outputs(5017) <= b and not a;
    layer2_outputs(5018) <= not a;
    layer2_outputs(5019) <= not a or b;
    layer2_outputs(5020) <= a and not b;
    layer2_outputs(5021) <= a or b;
    layer2_outputs(5022) <= a and b;
    layer2_outputs(5023) <= not (a and b);
    layer2_outputs(5024) <= not b;
    layer2_outputs(5025) <= not b;
    layer2_outputs(5026) <= not a or b;
    layer2_outputs(5027) <= not b;
    layer2_outputs(5028) <= 1'b1;
    layer2_outputs(5029) <= not a;
    layer2_outputs(5030) <= b;
    layer2_outputs(5031) <= a and not b;
    layer2_outputs(5032) <= a and b;
    layer2_outputs(5033) <= not b;
    layer2_outputs(5034) <= a and b;
    layer2_outputs(5035) <= not (a or b);
    layer2_outputs(5036) <= not b;
    layer2_outputs(5037) <= b and not a;
    layer2_outputs(5038) <= not b or a;
    layer2_outputs(5039) <= a;
    layer2_outputs(5040) <= not (a or b);
    layer2_outputs(5041) <= 1'b0;
    layer2_outputs(5042) <= not (a xor b);
    layer2_outputs(5043) <= b and not a;
    layer2_outputs(5044) <= not a or b;
    layer2_outputs(5045) <= a and b;
    layer2_outputs(5046) <= a and not b;
    layer2_outputs(5047) <= b and not a;
    layer2_outputs(5048) <= not b or a;
    layer2_outputs(5049) <= not (a or b);
    layer2_outputs(5050) <= a and not b;
    layer2_outputs(5051) <= b and not a;
    layer2_outputs(5052) <= a;
    layer2_outputs(5053) <= not a or b;
    layer2_outputs(5054) <= not b or a;
    layer2_outputs(5055) <= not b or a;
    layer2_outputs(5056) <= a or b;
    layer2_outputs(5057) <= 1'b1;
    layer2_outputs(5058) <= a and b;
    layer2_outputs(5059) <= a;
    layer2_outputs(5060) <= not (a xor b);
    layer2_outputs(5061) <= not a or b;
    layer2_outputs(5062) <= not b;
    layer2_outputs(5063) <= not b;
    layer2_outputs(5064) <= a or b;
    layer2_outputs(5065) <= a xor b;
    layer2_outputs(5066) <= a xor b;
    layer2_outputs(5067) <= a;
    layer2_outputs(5068) <= not a;
    layer2_outputs(5069) <= not b;
    layer2_outputs(5070) <= a;
    layer2_outputs(5071) <= a xor b;
    layer2_outputs(5072) <= 1'b0;
    layer2_outputs(5073) <= 1'b0;
    layer2_outputs(5074) <= 1'b0;
    layer2_outputs(5075) <= a xor b;
    layer2_outputs(5076) <= a and b;
    layer2_outputs(5077) <= not a;
    layer2_outputs(5078) <= a;
    layer2_outputs(5079) <= not b or a;
    layer2_outputs(5080) <= a and b;
    layer2_outputs(5081) <= a and b;
    layer2_outputs(5082) <= not a;
    layer2_outputs(5083) <= not b or a;
    layer2_outputs(5084) <= b;
    layer2_outputs(5085) <= not a;
    layer2_outputs(5086) <= a;
    layer2_outputs(5087) <= a;
    layer2_outputs(5088) <= b;
    layer2_outputs(5089) <= not (a and b);
    layer2_outputs(5090) <= a xor b;
    layer2_outputs(5091) <= not (a xor b);
    layer2_outputs(5092) <= a;
    layer2_outputs(5093) <= not b or a;
    layer2_outputs(5094) <= a or b;
    layer2_outputs(5095) <= a or b;
    layer2_outputs(5096) <= a and not b;
    layer2_outputs(5097) <= a or b;
    layer2_outputs(5098) <= not b or a;
    layer2_outputs(5099) <= not a or b;
    layer2_outputs(5100) <= a;
    layer2_outputs(5101) <= a and b;
    layer2_outputs(5102) <= not b or a;
    layer2_outputs(5103) <= not a;
    layer2_outputs(5104) <= a xor b;
    layer2_outputs(5105) <= b;
    layer2_outputs(5106) <= not (a and b);
    layer2_outputs(5107) <= not (a and b);
    layer2_outputs(5108) <= 1'b0;
    layer2_outputs(5109) <= 1'b1;
    layer2_outputs(5110) <= not b;
    layer2_outputs(5111) <= not a;
    layer2_outputs(5112) <= b;
    layer2_outputs(5113) <= not a or b;
    layer2_outputs(5114) <= b;
    layer2_outputs(5115) <= not (a xor b);
    layer2_outputs(5116) <= a and not b;
    layer2_outputs(5117) <= not b;
    layer2_outputs(5118) <= b;
    layer2_outputs(5119) <= a;
    layer2_outputs(5120) <= b and not a;
    layer2_outputs(5121) <= not (a or b);
    layer2_outputs(5122) <= a and not b;
    layer2_outputs(5123) <= a;
    layer2_outputs(5124) <= not (a or b);
    layer2_outputs(5125) <= 1'b0;
    layer2_outputs(5126) <= not b;
    layer2_outputs(5127) <= not (a xor b);
    layer2_outputs(5128) <= not b or a;
    layer2_outputs(5129) <= a and b;
    layer2_outputs(5130) <= not b;
    layer2_outputs(5131) <= not a;
    layer2_outputs(5132) <= not a;
    layer2_outputs(5133) <= a and not b;
    layer2_outputs(5134) <= not b or a;
    layer2_outputs(5135) <= not b;
    layer2_outputs(5136) <= a or b;
    layer2_outputs(5137) <= a and b;
    layer2_outputs(5138) <= not a or b;
    layer2_outputs(5139) <= not (a xor b);
    layer2_outputs(5140) <= not a;
    layer2_outputs(5141) <= a and b;
    layer2_outputs(5142) <= not (a or b);
    layer2_outputs(5143) <= not b;
    layer2_outputs(5144) <= not (a and b);
    layer2_outputs(5145) <= a and b;
    layer2_outputs(5146) <= b;
    layer2_outputs(5147) <= a xor b;
    layer2_outputs(5148) <= a or b;
    layer2_outputs(5149) <= a;
    layer2_outputs(5150) <= a and not b;
    layer2_outputs(5151) <= a or b;
    layer2_outputs(5152) <= not (a and b);
    layer2_outputs(5153) <= a and not b;
    layer2_outputs(5154) <= not b;
    layer2_outputs(5155) <= a;
    layer2_outputs(5156) <= not (a or b);
    layer2_outputs(5157) <= not a;
    layer2_outputs(5158) <= not b;
    layer2_outputs(5159) <= b and not a;
    layer2_outputs(5160) <= b and not a;
    layer2_outputs(5161) <= not b;
    layer2_outputs(5162) <= a;
    layer2_outputs(5163) <= a;
    layer2_outputs(5164) <= not (a or b);
    layer2_outputs(5165) <= a and not b;
    layer2_outputs(5166) <= b and not a;
    layer2_outputs(5167) <= a;
    layer2_outputs(5168) <= not b or a;
    layer2_outputs(5169) <= not (a or b);
    layer2_outputs(5170) <= a;
    layer2_outputs(5171) <= not a;
    layer2_outputs(5172) <= b;
    layer2_outputs(5173) <= not b;
    layer2_outputs(5174) <= b and not a;
    layer2_outputs(5175) <= b;
    layer2_outputs(5176) <= a;
    layer2_outputs(5177) <= not b or a;
    layer2_outputs(5178) <= 1'b1;
    layer2_outputs(5179) <= not b;
    layer2_outputs(5180) <= not (a and b);
    layer2_outputs(5181) <= a xor b;
    layer2_outputs(5182) <= not b;
    layer2_outputs(5183) <= a or b;
    layer2_outputs(5184) <= a;
    layer2_outputs(5185) <= b;
    layer2_outputs(5186) <= 1'b1;
    layer2_outputs(5187) <= not b;
    layer2_outputs(5188) <= a;
    layer2_outputs(5189) <= not a;
    layer2_outputs(5190) <= a xor b;
    layer2_outputs(5191) <= b;
    layer2_outputs(5192) <= not (a and b);
    layer2_outputs(5193) <= a or b;
    layer2_outputs(5194) <= 1'b1;
    layer2_outputs(5195) <= 1'b1;
    layer2_outputs(5196) <= b;
    layer2_outputs(5197) <= b;
    layer2_outputs(5198) <= a;
    layer2_outputs(5199) <= not a or b;
    layer2_outputs(5200) <= b;
    layer2_outputs(5201) <= not b;
    layer2_outputs(5202) <= not (a xor b);
    layer2_outputs(5203) <= a or b;
    layer2_outputs(5204) <= b;
    layer2_outputs(5205) <= a;
    layer2_outputs(5206) <= 1'b0;
    layer2_outputs(5207) <= not a or b;
    layer2_outputs(5208) <= not a;
    layer2_outputs(5209) <= not b;
    layer2_outputs(5210) <= not (a xor b);
    layer2_outputs(5211) <= a;
    layer2_outputs(5212) <= not a;
    layer2_outputs(5213) <= 1'b1;
    layer2_outputs(5214) <= not a or b;
    layer2_outputs(5215) <= not b or a;
    layer2_outputs(5216) <= a and b;
    layer2_outputs(5217) <= not (a and b);
    layer2_outputs(5218) <= not b;
    layer2_outputs(5219) <= not (a xor b);
    layer2_outputs(5220) <= not a;
    layer2_outputs(5221) <= not a;
    layer2_outputs(5222) <= a or b;
    layer2_outputs(5223) <= not a or b;
    layer2_outputs(5224) <= not b;
    layer2_outputs(5225) <= b;
    layer2_outputs(5226) <= b;
    layer2_outputs(5227) <= b;
    layer2_outputs(5228) <= b;
    layer2_outputs(5229) <= not (a or b);
    layer2_outputs(5230) <= not b;
    layer2_outputs(5231) <= a;
    layer2_outputs(5232) <= not b or a;
    layer2_outputs(5233) <= not b or a;
    layer2_outputs(5234) <= b;
    layer2_outputs(5235) <= not (a xor b);
    layer2_outputs(5236) <= a and not b;
    layer2_outputs(5237) <= a or b;
    layer2_outputs(5238) <= not b;
    layer2_outputs(5239) <= not a or b;
    layer2_outputs(5240) <= not a or b;
    layer2_outputs(5241) <= b and not a;
    layer2_outputs(5242) <= not a;
    layer2_outputs(5243) <= not (a or b);
    layer2_outputs(5244) <= a;
    layer2_outputs(5245) <= a xor b;
    layer2_outputs(5246) <= 1'b1;
    layer2_outputs(5247) <= a;
    layer2_outputs(5248) <= a;
    layer2_outputs(5249) <= not b or a;
    layer2_outputs(5250) <= not (a or b);
    layer2_outputs(5251) <= a and not b;
    layer2_outputs(5252) <= not a;
    layer2_outputs(5253) <= a;
    layer2_outputs(5254) <= not a or b;
    layer2_outputs(5255) <= a xor b;
    layer2_outputs(5256) <= not a;
    layer2_outputs(5257) <= not (a or b);
    layer2_outputs(5258) <= 1'b1;
    layer2_outputs(5259) <= not b;
    layer2_outputs(5260) <= not a;
    layer2_outputs(5261) <= a and b;
    layer2_outputs(5262) <= not b;
    layer2_outputs(5263) <= a and not b;
    layer2_outputs(5264) <= not (a or b);
    layer2_outputs(5265) <= not b or a;
    layer2_outputs(5266) <= not a or b;
    layer2_outputs(5267) <= a xor b;
    layer2_outputs(5268) <= b and not a;
    layer2_outputs(5269) <= not b;
    layer2_outputs(5270) <= not (a or b);
    layer2_outputs(5271) <= not a;
    layer2_outputs(5272) <= not a;
    layer2_outputs(5273) <= a;
    layer2_outputs(5274) <= not b;
    layer2_outputs(5275) <= b and not a;
    layer2_outputs(5276) <= a and not b;
    layer2_outputs(5277) <= a;
    layer2_outputs(5278) <= a and b;
    layer2_outputs(5279) <= 1'b1;
    layer2_outputs(5280) <= a or b;
    layer2_outputs(5281) <= not a;
    layer2_outputs(5282) <= not b or a;
    layer2_outputs(5283) <= not (a xor b);
    layer2_outputs(5284) <= not b;
    layer2_outputs(5285) <= a or b;
    layer2_outputs(5286) <= a;
    layer2_outputs(5287) <= 1'b1;
    layer2_outputs(5288) <= not (a or b);
    layer2_outputs(5289) <= not b or a;
    layer2_outputs(5290) <= not b or a;
    layer2_outputs(5291) <= not b;
    layer2_outputs(5292) <= not b;
    layer2_outputs(5293) <= not (a and b);
    layer2_outputs(5294) <= not b;
    layer2_outputs(5295) <= 1'b1;
    layer2_outputs(5296) <= b;
    layer2_outputs(5297) <= b;
    layer2_outputs(5298) <= not a;
    layer2_outputs(5299) <= not b or a;
    layer2_outputs(5300) <= a;
    layer2_outputs(5301) <= not a or b;
    layer2_outputs(5302) <= not a or b;
    layer2_outputs(5303) <= a and b;
    layer2_outputs(5304) <= not (a and b);
    layer2_outputs(5305) <= a;
    layer2_outputs(5306) <= a and not b;
    layer2_outputs(5307) <= a or b;
    layer2_outputs(5308) <= not b or a;
    layer2_outputs(5309) <= not a;
    layer2_outputs(5310) <= a xor b;
    layer2_outputs(5311) <= not b or a;
    layer2_outputs(5312) <= not a;
    layer2_outputs(5313) <= not (a xor b);
    layer2_outputs(5314) <= a;
    layer2_outputs(5315) <= a and not b;
    layer2_outputs(5316) <= not (a or b);
    layer2_outputs(5317) <= b and not a;
    layer2_outputs(5318) <= not a or b;
    layer2_outputs(5319) <= a;
    layer2_outputs(5320) <= a and b;
    layer2_outputs(5321) <= b and not a;
    layer2_outputs(5322) <= a xor b;
    layer2_outputs(5323) <= b and not a;
    layer2_outputs(5324) <= not a;
    layer2_outputs(5325) <= not b;
    layer2_outputs(5326) <= not a;
    layer2_outputs(5327) <= a;
    layer2_outputs(5328) <= not b;
    layer2_outputs(5329) <= not a;
    layer2_outputs(5330) <= a and b;
    layer2_outputs(5331) <= not b;
    layer2_outputs(5332) <= a;
    layer2_outputs(5333) <= not b;
    layer2_outputs(5334) <= not a;
    layer2_outputs(5335) <= b;
    layer2_outputs(5336) <= b;
    layer2_outputs(5337) <= a xor b;
    layer2_outputs(5338) <= b;
    layer2_outputs(5339) <= not (a xor b);
    layer2_outputs(5340) <= not a;
    layer2_outputs(5341) <= not a;
    layer2_outputs(5342) <= not b or a;
    layer2_outputs(5343) <= b;
    layer2_outputs(5344) <= a or b;
    layer2_outputs(5345) <= b;
    layer2_outputs(5346) <= not a;
    layer2_outputs(5347) <= a or b;
    layer2_outputs(5348) <= not a;
    layer2_outputs(5349) <= a xor b;
    layer2_outputs(5350) <= not a;
    layer2_outputs(5351) <= b;
    layer2_outputs(5352) <= not a;
    layer2_outputs(5353) <= a and b;
    layer2_outputs(5354) <= not (a or b);
    layer2_outputs(5355) <= not b;
    layer2_outputs(5356) <= a;
    layer2_outputs(5357) <= a or b;
    layer2_outputs(5358) <= not a or b;
    layer2_outputs(5359) <= 1'b1;
    layer2_outputs(5360) <= not b or a;
    layer2_outputs(5361) <= not b or a;
    layer2_outputs(5362) <= b;
    layer2_outputs(5363) <= not (a xor b);
    layer2_outputs(5364) <= a and not b;
    layer2_outputs(5365) <= not a;
    layer2_outputs(5366) <= a;
    layer2_outputs(5367) <= a;
    layer2_outputs(5368) <= not a or b;
    layer2_outputs(5369) <= b;
    layer2_outputs(5370) <= b;
    layer2_outputs(5371) <= not a or b;
    layer2_outputs(5372) <= a;
    layer2_outputs(5373) <= not a;
    layer2_outputs(5374) <= not b;
    layer2_outputs(5375) <= not (a xor b);
    layer2_outputs(5376) <= not a;
    layer2_outputs(5377) <= not a;
    layer2_outputs(5378) <= not a;
    layer2_outputs(5379) <= a and not b;
    layer2_outputs(5380) <= a;
    layer2_outputs(5381) <= b;
    layer2_outputs(5382) <= not (a or b);
    layer2_outputs(5383) <= b;
    layer2_outputs(5384) <= a;
    layer2_outputs(5385) <= b;
    layer2_outputs(5386) <= not a;
    layer2_outputs(5387) <= not b;
    layer2_outputs(5388) <= a;
    layer2_outputs(5389) <= not (a xor b);
    layer2_outputs(5390) <= not a;
    layer2_outputs(5391) <= b;
    layer2_outputs(5392) <= not (a xor b);
    layer2_outputs(5393) <= not (a or b);
    layer2_outputs(5394) <= a and not b;
    layer2_outputs(5395) <= not (a xor b);
    layer2_outputs(5396) <= a;
    layer2_outputs(5397) <= not (a and b);
    layer2_outputs(5398) <= not a or b;
    layer2_outputs(5399) <= a and b;
    layer2_outputs(5400) <= a and not b;
    layer2_outputs(5401) <= not (a xor b);
    layer2_outputs(5402) <= b and not a;
    layer2_outputs(5403) <= a xor b;
    layer2_outputs(5404) <= b;
    layer2_outputs(5405) <= a;
    layer2_outputs(5406) <= a or b;
    layer2_outputs(5407) <= not a;
    layer2_outputs(5408) <= not a or b;
    layer2_outputs(5409) <= b and not a;
    layer2_outputs(5410) <= a;
    layer2_outputs(5411) <= not a;
    layer2_outputs(5412) <= a;
    layer2_outputs(5413) <= not (a or b);
    layer2_outputs(5414) <= not b;
    layer2_outputs(5415) <= not b;
    layer2_outputs(5416) <= not b or a;
    layer2_outputs(5417) <= a or b;
    layer2_outputs(5418) <= b;
    layer2_outputs(5419) <= not a;
    layer2_outputs(5420) <= 1'b1;
    layer2_outputs(5421) <= a or b;
    layer2_outputs(5422) <= a xor b;
    layer2_outputs(5423) <= not a or b;
    layer2_outputs(5424) <= a;
    layer2_outputs(5425) <= not (a or b);
    layer2_outputs(5426) <= not a;
    layer2_outputs(5427) <= b;
    layer2_outputs(5428) <= a;
    layer2_outputs(5429) <= not b;
    layer2_outputs(5430) <= a and not b;
    layer2_outputs(5431) <= not a or b;
    layer2_outputs(5432) <= a xor b;
    layer2_outputs(5433) <= not a;
    layer2_outputs(5434) <= not (a xor b);
    layer2_outputs(5435) <= b;
    layer2_outputs(5436) <= a and not b;
    layer2_outputs(5437) <= a or b;
    layer2_outputs(5438) <= b;
    layer2_outputs(5439) <= a xor b;
    layer2_outputs(5440) <= not b;
    layer2_outputs(5441) <= not (a xor b);
    layer2_outputs(5442) <= a xor b;
    layer2_outputs(5443) <= b and not a;
    layer2_outputs(5444) <= a;
    layer2_outputs(5445) <= a and not b;
    layer2_outputs(5446) <= a and not b;
    layer2_outputs(5447) <= a;
    layer2_outputs(5448) <= b;
    layer2_outputs(5449) <= 1'b1;
    layer2_outputs(5450) <= not a or b;
    layer2_outputs(5451) <= not (a and b);
    layer2_outputs(5452) <= not b;
    layer2_outputs(5453) <= b;
    layer2_outputs(5454) <= a and not b;
    layer2_outputs(5455) <= b;
    layer2_outputs(5456) <= not b;
    layer2_outputs(5457) <= not (a or b);
    layer2_outputs(5458) <= not (a and b);
    layer2_outputs(5459) <= a and not b;
    layer2_outputs(5460) <= not (a or b);
    layer2_outputs(5461) <= not b;
    layer2_outputs(5462) <= a and b;
    layer2_outputs(5463) <= not (a or b);
    layer2_outputs(5464) <= a;
    layer2_outputs(5465) <= a or b;
    layer2_outputs(5466) <= a and b;
    layer2_outputs(5467) <= not b;
    layer2_outputs(5468) <= not b;
    layer2_outputs(5469) <= not (a and b);
    layer2_outputs(5470) <= not b;
    layer2_outputs(5471) <= not a or b;
    layer2_outputs(5472) <= a and b;
    layer2_outputs(5473) <= a and b;
    layer2_outputs(5474) <= not (a xor b);
    layer2_outputs(5475) <= b;
    layer2_outputs(5476) <= not a;
    layer2_outputs(5477) <= not a;
    layer2_outputs(5478) <= a and b;
    layer2_outputs(5479) <= a;
    layer2_outputs(5480) <= not (a xor b);
    layer2_outputs(5481) <= b;
    layer2_outputs(5482) <= a or b;
    layer2_outputs(5483) <= not a;
    layer2_outputs(5484) <= not b;
    layer2_outputs(5485) <= a and not b;
    layer2_outputs(5486) <= not b or a;
    layer2_outputs(5487) <= a xor b;
    layer2_outputs(5488) <= not (a or b);
    layer2_outputs(5489) <= not (a and b);
    layer2_outputs(5490) <= not (a xor b);
    layer2_outputs(5491) <= b and not a;
    layer2_outputs(5492) <= not (a and b);
    layer2_outputs(5493) <= 1'b1;
    layer2_outputs(5494) <= a xor b;
    layer2_outputs(5495) <= not (a xor b);
    layer2_outputs(5496) <= a and b;
    layer2_outputs(5497) <= b;
    layer2_outputs(5498) <= a;
    layer2_outputs(5499) <= not a or b;
    layer2_outputs(5500) <= b and not a;
    layer2_outputs(5501) <= a and not b;
    layer2_outputs(5502) <= b;
    layer2_outputs(5503) <= not (a or b);
    layer2_outputs(5504) <= not a or b;
    layer2_outputs(5505) <= b;
    layer2_outputs(5506) <= a and b;
    layer2_outputs(5507) <= a and b;
    layer2_outputs(5508) <= a;
    layer2_outputs(5509) <= not (a xor b);
    layer2_outputs(5510) <= a;
    layer2_outputs(5511) <= a and b;
    layer2_outputs(5512) <= not b;
    layer2_outputs(5513) <= b;
    layer2_outputs(5514) <= b and not a;
    layer2_outputs(5515) <= b;
    layer2_outputs(5516) <= a and b;
    layer2_outputs(5517) <= 1'b0;
    layer2_outputs(5518) <= not (a or b);
    layer2_outputs(5519) <= not b;
    layer2_outputs(5520) <= a;
    layer2_outputs(5521) <= not a;
    layer2_outputs(5522) <= b;
    layer2_outputs(5523) <= not b;
    layer2_outputs(5524) <= not b;
    layer2_outputs(5525) <= a and b;
    layer2_outputs(5526) <= a or b;
    layer2_outputs(5527) <= not (a or b);
    layer2_outputs(5528) <= not (a or b);
    layer2_outputs(5529) <= a and not b;
    layer2_outputs(5530) <= not a;
    layer2_outputs(5531) <= a and not b;
    layer2_outputs(5532) <= a xor b;
    layer2_outputs(5533) <= not (a xor b);
    layer2_outputs(5534) <= not a;
    layer2_outputs(5535) <= 1'b1;
    layer2_outputs(5536) <= not (a xor b);
    layer2_outputs(5537) <= 1'b0;
    layer2_outputs(5538) <= not a or b;
    layer2_outputs(5539) <= 1'b0;
    layer2_outputs(5540) <= 1'b1;
    layer2_outputs(5541) <= not b or a;
    layer2_outputs(5542) <= a and not b;
    layer2_outputs(5543) <= a or b;
    layer2_outputs(5544) <= not a;
    layer2_outputs(5545) <= not (a and b);
    layer2_outputs(5546) <= a or b;
    layer2_outputs(5547) <= a and not b;
    layer2_outputs(5548) <= not (a or b);
    layer2_outputs(5549) <= not (a and b);
    layer2_outputs(5550) <= 1'b0;
    layer2_outputs(5551) <= not a or b;
    layer2_outputs(5552) <= not a or b;
    layer2_outputs(5553) <= a and b;
    layer2_outputs(5554) <= a and b;
    layer2_outputs(5555) <= a xor b;
    layer2_outputs(5556) <= not a or b;
    layer2_outputs(5557) <= not a;
    layer2_outputs(5558) <= not b;
    layer2_outputs(5559) <= not b;
    layer2_outputs(5560) <= not a;
    layer2_outputs(5561) <= b and not a;
    layer2_outputs(5562) <= not a;
    layer2_outputs(5563) <= not b or a;
    layer2_outputs(5564) <= not b or a;
    layer2_outputs(5565) <= a xor b;
    layer2_outputs(5566) <= not a;
    layer2_outputs(5567) <= a xor b;
    layer2_outputs(5568) <= not (a or b);
    layer2_outputs(5569) <= a;
    layer2_outputs(5570) <= a or b;
    layer2_outputs(5571) <= a and not b;
    layer2_outputs(5572) <= a and not b;
    layer2_outputs(5573) <= a or b;
    layer2_outputs(5574) <= not a;
    layer2_outputs(5575) <= a or b;
    layer2_outputs(5576) <= not (a or b);
    layer2_outputs(5577) <= b;
    layer2_outputs(5578) <= not b or a;
    layer2_outputs(5579) <= 1'b1;
    layer2_outputs(5580) <= not a or b;
    layer2_outputs(5581) <= a;
    layer2_outputs(5582) <= not (a and b);
    layer2_outputs(5583) <= 1'b0;
    layer2_outputs(5584) <= not b or a;
    layer2_outputs(5585) <= a;
    layer2_outputs(5586) <= not (a and b);
    layer2_outputs(5587) <= a;
    layer2_outputs(5588) <= not b or a;
    layer2_outputs(5589) <= not b;
    layer2_outputs(5590) <= not b;
    layer2_outputs(5591) <= 1'b0;
    layer2_outputs(5592) <= a;
    layer2_outputs(5593) <= a and not b;
    layer2_outputs(5594) <= not b;
    layer2_outputs(5595) <= a and not b;
    layer2_outputs(5596) <= not a;
    layer2_outputs(5597) <= a;
    layer2_outputs(5598) <= a xor b;
    layer2_outputs(5599) <= a and b;
    layer2_outputs(5600) <= a and not b;
    layer2_outputs(5601) <= b;
    layer2_outputs(5602) <= not b or a;
    layer2_outputs(5603) <= not b or a;
    layer2_outputs(5604) <= a and not b;
    layer2_outputs(5605) <= not a;
    layer2_outputs(5606) <= not b or a;
    layer2_outputs(5607) <= not (a or b);
    layer2_outputs(5608) <= not b or a;
    layer2_outputs(5609) <= a;
    layer2_outputs(5610) <= not b;
    layer2_outputs(5611) <= a;
    layer2_outputs(5612) <= a and b;
    layer2_outputs(5613) <= a;
    layer2_outputs(5614) <= not b;
    layer2_outputs(5615) <= not (a and b);
    layer2_outputs(5616) <= b;
    layer2_outputs(5617) <= 1'b0;
    layer2_outputs(5618) <= a and b;
    layer2_outputs(5619) <= a and not b;
    layer2_outputs(5620) <= a;
    layer2_outputs(5621) <= not a or b;
    layer2_outputs(5622) <= a;
    layer2_outputs(5623) <= a or b;
    layer2_outputs(5624) <= not (a xor b);
    layer2_outputs(5625) <= a xor b;
    layer2_outputs(5626) <= 1'b1;
    layer2_outputs(5627) <= a xor b;
    layer2_outputs(5628) <= not b;
    layer2_outputs(5629) <= b and not a;
    layer2_outputs(5630) <= not b or a;
    layer2_outputs(5631) <= b;
    layer2_outputs(5632) <= not (a and b);
    layer2_outputs(5633) <= not (a xor b);
    layer2_outputs(5634) <= 1'b0;
    layer2_outputs(5635) <= not a or b;
    layer2_outputs(5636) <= not b or a;
    layer2_outputs(5637) <= a and not b;
    layer2_outputs(5638) <= a xor b;
    layer2_outputs(5639) <= a xor b;
    layer2_outputs(5640) <= not b;
    layer2_outputs(5641) <= not a;
    layer2_outputs(5642) <= not a;
    layer2_outputs(5643) <= not (a or b);
    layer2_outputs(5644) <= not b or a;
    layer2_outputs(5645) <= not (a or b);
    layer2_outputs(5646) <= not b;
    layer2_outputs(5647) <= not b or a;
    layer2_outputs(5648) <= a;
    layer2_outputs(5649) <= a xor b;
    layer2_outputs(5650) <= a and not b;
    layer2_outputs(5651) <= b and not a;
    layer2_outputs(5652) <= not a;
    layer2_outputs(5653) <= not b or a;
    layer2_outputs(5654) <= not (a and b);
    layer2_outputs(5655) <= a and b;
    layer2_outputs(5656) <= not a;
    layer2_outputs(5657) <= not a;
    layer2_outputs(5658) <= not b or a;
    layer2_outputs(5659) <= b;
    layer2_outputs(5660) <= b;
    layer2_outputs(5661) <= not a or b;
    layer2_outputs(5662) <= a xor b;
    layer2_outputs(5663) <= b;
    layer2_outputs(5664) <= a;
    layer2_outputs(5665) <= not (a and b);
    layer2_outputs(5666) <= not a or b;
    layer2_outputs(5667) <= not a;
    layer2_outputs(5668) <= not (a or b);
    layer2_outputs(5669) <= not (a and b);
    layer2_outputs(5670) <= a and b;
    layer2_outputs(5671) <= a xor b;
    layer2_outputs(5672) <= b and not a;
    layer2_outputs(5673) <= not a;
    layer2_outputs(5674) <= not b or a;
    layer2_outputs(5675) <= b and not a;
    layer2_outputs(5676) <= not a;
    layer2_outputs(5677) <= a and not b;
    layer2_outputs(5678) <= not b;
    layer2_outputs(5679) <= not b;
    layer2_outputs(5680) <= not a or b;
    layer2_outputs(5681) <= not b or a;
    layer2_outputs(5682) <= not a or b;
    layer2_outputs(5683) <= not (a xor b);
    layer2_outputs(5684) <= not a;
    layer2_outputs(5685) <= b and not a;
    layer2_outputs(5686) <= a and not b;
    layer2_outputs(5687) <= a and b;
    layer2_outputs(5688) <= a;
    layer2_outputs(5689) <= 1'b0;
    layer2_outputs(5690) <= a xor b;
    layer2_outputs(5691) <= not (a or b);
    layer2_outputs(5692) <= a and b;
    layer2_outputs(5693) <= b;
    layer2_outputs(5694) <= a xor b;
    layer2_outputs(5695) <= a;
    layer2_outputs(5696) <= not a or b;
    layer2_outputs(5697) <= a;
    layer2_outputs(5698) <= b;
    layer2_outputs(5699) <= not (a or b);
    layer2_outputs(5700) <= not a;
    layer2_outputs(5701) <= not b;
    layer2_outputs(5702) <= not (a xor b);
    layer2_outputs(5703) <= not b or a;
    layer2_outputs(5704) <= not a;
    layer2_outputs(5705) <= not a or b;
    layer2_outputs(5706) <= not (a or b);
    layer2_outputs(5707) <= not a;
    layer2_outputs(5708) <= not a or b;
    layer2_outputs(5709) <= b and not a;
    layer2_outputs(5710) <= b;
    layer2_outputs(5711) <= not b or a;
    layer2_outputs(5712) <= a;
    layer2_outputs(5713) <= not (a xor b);
    layer2_outputs(5714) <= not a;
    layer2_outputs(5715) <= 1'b1;
    layer2_outputs(5716) <= not a;
    layer2_outputs(5717) <= not (a or b);
    layer2_outputs(5718) <= a xor b;
    layer2_outputs(5719) <= not a;
    layer2_outputs(5720) <= not b;
    layer2_outputs(5721) <= a;
    layer2_outputs(5722) <= not (a and b);
    layer2_outputs(5723) <= not a or b;
    layer2_outputs(5724) <= b;
    layer2_outputs(5725) <= a;
    layer2_outputs(5726) <= not a or b;
    layer2_outputs(5727) <= a or b;
    layer2_outputs(5728) <= not (a or b);
    layer2_outputs(5729) <= not b;
    layer2_outputs(5730) <= a xor b;
    layer2_outputs(5731) <= not (a or b);
    layer2_outputs(5732) <= a and b;
    layer2_outputs(5733) <= a and b;
    layer2_outputs(5734) <= b;
    layer2_outputs(5735) <= a xor b;
    layer2_outputs(5736) <= not b or a;
    layer2_outputs(5737) <= b;
    layer2_outputs(5738) <= b;
    layer2_outputs(5739) <= not b;
    layer2_outputs(5740) <= a and not b;
    layer2_outputs(5741) <= a or b;
    layer2_outputs(5742) <= not b;
    layer2_outputs(5743) <= b;
    layer2_outputs(5744) <= 1'b1;
    layer2_outputs(5745) <= not (a xor b);
    layer2_outputs(5746) <= b and not a;
    layer2_outputs(5747) <= b and not a;
    layer2_outputs(5748) <= not (a or b);
    layer2_outputs(5749) <= not a or b;
    layer2_outputs(5750) <= b and not a;
    layer2_outputs(5751) <= not (a and b);
    layer2_outputs(5752) <= b;
    layer2_outputs(5753) <= a and not b;
    layer2_outputs(5754) <= not b or a;
    layer2_outputs(5755) <= a and b;
    layer2_outputs(5756) <= a or b;
    layer2_outputs(5757) <= not a;
    layer2_outputs(5758) <= b;
    layer2_outputs(5759) <= not (a and b);
    layer2_outputs(5760) <= a xor b;
    layer2_outputs(5761) <= a xor b;
    layer2_outputs(5762) <= a or b;
    layer2_outputs(5763) <= a and b;
    layer2_outputs(5764) <= not b;
    layer2_outputs(5765) <= b;
    layer2_outputs(5766) <= a xor b;
    layer2_outputs(5767) <= a and b;
    layer2_outputs(5768) <= b;
    layer2_outputs(5769) <= a;
    layer2_outputs(5770) <= b and not a;
    layer2_outputs(5771) <= 1'b0;
    layer2_outputs(5772) <= a xor b;
    layer2_outputs(5773) <= a;
    layer2_outputs(5774) <= a;
    layer2_outputs(5775) <= not a or b;
    layer2_outputs(5776) <= b;
    layer2_outputs(5777) <= not b;
    layer2_outputs(5778) <= not b or a;
    layer2_outputs(5779) <= not b;
    layer2_outputs(5780) <= b;
    layer2_outputs(5781) <= not a;
    layer2_outputs(5782) <= not (a and b);
    layer2_outputs(5783) <= a;
    layer2_outputs(5784) <= not b or a;
    layer2_outputs(5785) <= b and not a;
    layer2_outputs(5786) <= not (a or b);
    layer2_outputs(5787) <= a and not b;
    layer2_outputs(5788) <= not b;
    layer2_outputs(5789) <= a and not b;
    layer2_outputs(5790) <= 1'b0;
    layer2_outputs(5791) <= a and b;
    layer2_outputs(5792) <= a;
    layer2_outputs(5793) <= not a;
    layer2_outputs(5794) <= a;
    layer2_outputs(5795) <= not b;
    layer2_outputs(5796) <= b;
    layer2_outputs(5797) <= not a;
    layer2_outputs(5798) <= not (a or b);
    layer2_outputs(5799) <= not b;
    layer2_outputs(5800) <= not (a and b);
    layer2_outputs(5801) <= not (a and b);
    layer2_outputs(5802) <= not a;
    layer2_outputs(5803) <= a and not b;
    layer2_outputs(5804) <= a;
    layer2_outputs(5805) <= not (a and b);
    layer2_outputs(5806) <= not (a and b);
    layer2_outputs(5807) <= a or b;
    layer2_outputs(5808) <= not (a and b);
    layer2_outputs(5809) <= b and not a;
    layer2_outputs(5810) <= not a;
    layer2_outputs(5811) <= a or b;
    layer2_outputs(5812) <= a and not b;
    layer2_outputs(5813) <= 1'b1;
    layer2_outputs(5814) <= not a or b;
    layer2_outputs(5815) <= b;
    layer2_outputs(5816) <= not a;
    layer2_outputs(5817) <= not (a and b);
    layer2_outputs(5818) <= a;
    layer2_outputs(5819) <= b;
    layer2_outputs(5820) <= not a;
    layer2_outputs(5821) <= not b;
    layer2_outputs(5822) <= b;
    layer2_outputs(5823) <= not (a and b);
    layer2_outputs(5824) <= not b;
    layer2_outputs(5825) <= not (a and b);
    layer2_outputs(5826) <= not (a or b);
    layer2_outputs(5827) <= not (a or b);
    layer2_outputs(5828) <= not b;
    layer2_outputs(5829) <= not b;
    layer2_outputs(5830) <= not a;
    layer2_outputs(5831) <= a and not b;
    layer2_outputs(5832) <= a or b;
    layer2_outputs(5833) <= a;
    layer2_outputs(5834) <= a and b;
    layer2_outputs(5835) <= not a or b;
    layer2_outputs(5836) <= a and not b;
    layer2_outputs(5837) <= a;
    layer2_outputs(5838) <= b and not a;
    layer2_outputs(5839) <= a xor b;
    layer2_outputs(5840) <= not a;
    layer2_outputs(5841) <= b and not a;
    layer2_outputs(5842) <= a and b;
    layer2_outputs(5843) <= not a or b;
    layer2_outputs(5844) <= b;
    layer2_outputs(5845) <= not (a or b);
    layer2_outputs(5846) <= not a or b;
    layer2_outputs(5847) <= b;
    layer2_outputs(5848) <= a xor b;
    layer2_outputs(5849) <= a;
    layer2_outputs(5850) <= b and not a;
    layer2_outputs(5851) <= a;
    layer2_outputs(5852) <= a or b;
    layer2_outputs(5853) <= a or b;
    layer2_outputs(5854) <= not (a xor b);
    layer2_outputs(5855) <= a;
    layer2_outputs(5856) <= b;
    layer2_outputs(5857) <= not b or a;
    layer2_outputs(5858) <= 1'b1;
    layer2_outputs(5859) <= not (a or b);
    layer2_outputs(5860) <= not b or a;
    layer2_outputs(5861) <= a xor b;
    layer2_outputs(5862) <= not (a xor b);
    layer2_outputs(5863) <= b and not a;
    layer2_outputs(5864) <= not a;
    layer2_outputs(5865) <= a;
    layer2_outputs(5866) <= not a;
    layer2_outputs(5867) <= not (a or b);
    layer2_outputs(5868) <= not (a xor b);
    layer2_outputs(5869) <= not b;
    layer2_outputs(5870) <= a or b;
    layer2_outputs(5871) <= not a;
    layer2_outputs(5872) <= a;
    layer2_outputs(5873) <= a and not b;
    layer2_outputs(5874) <= not a;
    layer2_outputs(5875) <= not b;
    layer2_outputs(5876) <= not a or b;
    layer2_outputs(5877) <= b;
    layer2_outputs(5878) <= b and not a;
    layer2_outputs(5879) <= a and b;
    layer2_outputs(5880) <= a and b;
    layer2_outputs(5881) <= b and not a;
    layer2_outputs(5882) <= 1'b0;
    layer2_outputs(5883) <= not b or a;
    layer2_outputs(5884) <= a and not b;
    layer2_outputs(5885) <= a and not b;
    layer2_outputs(5886) <= not a or b;
    layer2_outputs(5887) <= not b or a;
    layer2_outputs(5888) <= not (a or b);
    layer2_outputs(5889) <= b and not a;
    layer2_outputs(5890) <= a or b;
    layer2_outputs(5891) <= not a or b;
    layer2_outputs(5892) <= not b;
    layer2_outputs(5893) <= b and not a;
    layer2_outputs(5894) <= not a;
    layer2_outputs(5895) <= a and b;
    layer2_outputs(5896) <= not b;
    layer2_outputs(5897) <= not b;
    layer2_outputs(5898) <= not (a xor b);
    layer2_outputs(5899) <= not a;
    layer2_outputs(5900) <= a;
    layer2_outputs(5901) <= b;
    layer2_outputs(5902) <= a or b;
    layer2_outputs(5903) <= not (a and b);
    layer2_outputs(5904) <= a;
    layer2_outputs(5905) <= a;
    layer2_outputs(5906) <= a;
    layer2_outputs(5907) <= b;
    layer2_outputs(5908) <= not b or a;
    layer2_outputs(5909) <= a or b;
    layer2_outputs(5910) <= not (a xor b);
    layer2_outputs(5911) <= b;
    layer2_outputs(5912) <= not (a or b);
    layer2_outputs(5913) <= b;
    layer2_outputs(5914) <= not (a xor b);
    layer2_outputs(5915) <= a;
    layer2_outputs(5916) <= not b or a;
    layer2_outputs(5917) <= 1'b0;
    layer2_outputs(5918) <= b;
    layer2_outputs(5919) <= a or b;
    layer2_outputs(5920) <= not a;
    layer2_outputs(5921) <= a or b;
    layer2_outputs(5922) <= not (a and b);
    layer2_outputs(5923) <= a xor b;
    layer2_outputs(5924) <= a or b;
    layer2_outputs(5925) <= b and not a;
    layer2_outputs(5926) <= 1'b0;
    layer2_outputs(5927) <= a xor b;
    layer2_outputs(5928) <= a or b;
    layer2_outputs(5929) <= not b;
    layer2_outputs(5930) <= not (a xor b);
    layer2_outputs(5931) <= b and not a;
    layer2_outputs(5932) <= b;
    layer2_outputs(5933) <= not (a or b);
    layer2_outputs(5934) <= b;
    layer2_outputs(5935) <= not b;
    layer2_outputs(5936) <= a;
    layer2_outputs(5937) <= not b;
    layer2_outputs(5938) <= a and not b;
    layer2_outputs(5939) <= a;
    layer2_outputs(5940) <= not (a and b);
    layer2_outputs(5941) <= not b;
    layer2_outputs(5942) <= b;
    layer2_outputs(5943) <= a or b;
    layer2_outputs(5944) <= not b or a;
    layer2_outputs(5945) <= not (a or b);
    layer2_outputs(5946) <= a xor b;
    layer2_outputs(5947) <= a and b;
    layer2_outputs(5948) <= not b;
    layer2_outputs(5949) <= not a or b;
    layer2_outputs(5950) <= not (a or b);
    layer2_outputs(5951) <= not b or a;
    layer2_outputs(5952) <= not (a or b);
    layer2_outputs(5953) <= a and not b;
    layer2_outputs(5954) <= a xor b;
    layer2_outputs(5955) <= not (a xor b);
    layer2_outputs(5956) <= not b or a;
    layer2_outputs(5957) <= b;
    layer2_outputs(5958) <= a and not b;
    layer2_outputs(5959) <= not (a and b);
    layer2_outputs(5960) <= a;
    layer2_outputs(5961) <= not a;
    layer2_outputs(5962) <= not a;
    layer2_outputs(5963) <= not a or b;
    layer2_outputs(5964) <= not (a and b);
    layer2_outputs(5965) <= not b;
    layer2_outputs(5966) <= a and not b;
    layer2_outputs(5967) <= not b;
    layer2_outputs(5968) <= a or b;
    layer2_outputs(5969) <= b;
    layer2_outputs(5970) <= 1'b1;
    layer2_outputs(5971) <= 1'b0;
    layer2_outputs(5972) <= not b;
    layer2_outputs(5973) <= a and not b;
    layer2_outputs(5974) <= not b;
    layer2_outputs(5975) <= not b or a;
    layer2_outputs(5976) <= a or b;
    layer2_outputs(5977) <= a;
    layer2_outputs(5978) <= b;
    layer2_outputs(5979) <= a;
    layer2_outputs(5980) <= 1'b0;
    layer2_outputs(5981) <= not b or a;
    layer2_outputs(5982) <= not a;
    layer2_outputs(5983) <= a or b;
    layer2_outputs(5984) <= not b or a;
    layer2_outputs(5985) <= not a or b;
    layer2_outputs(5986) <= b;
    layer2_outputs(5987) <= a and not b;
    layer2_outputs(5988) <= not a;
    layer2_outputs(5989) <= not a or b;
    layer2_outputs(5990) <= not (a and b);
    layer2_outputs(5991) <= b;
    layer2_outputs(5992) <= b and not a;
    layer2_outputs(5993) <= not b;
    layer2_outputs(5994) <= not a;
    layer2_outputs(5995) <= b;
    layer2_outputs(5996) <= a or b;
    layer2_outputs(5997) <= a and b;
    layer2_outputs(5998) <= not (a and b);
    layer2_outputs(5999) <= not b;
    layer2_outputs(6000) <= not (a xor b);
    layer2_outputs(6001) <= not (a or b);
    layer2_outputs(6002) <= a or b;
    layer2_outputs(6003) <= b;
    layer2_outputs(6004) <= not (a and b);
    layer2_outputs(6005) <= b;
    layer2_outputs(6006) <= a and not b;
    layer2_outputs(6007) <= 1'b1;
    layer2_outputs(6008) <= b;
    layer2_outputs(6009) <= not b;
    layer2_outputs(6010) <= a;
    layer2_outputs(6011) <= a and not b;
    layer2_outputs(6012) <= not a;
    layer2_outputs(6013) <= b;
    layer2_outputs(6014) <= a;
    layer2_outputs(6015) <= b and not a;
    layer2_outputs(6016) <= a and b;
    layer2_outputs(6017) <= not b;
    layer2_outputs(6018) <= a;
    layer2_outputs(6019) <= a and not b;
    layer2_outputs(6020) <= not (a or b);
    layer2_outputs(6021) <= a or b;
    layer2_outputs(6022) <= a;
    layer2_outputs(6023) <= b and not a;
    layer2_outputs(6024) <= a and not b;
    layer2_outputs(6025) <= not (a and b);
    layer2_outputs(6026) <= a;
    layer2_outputs(6027) <= a;
    layer2_outputs(6028) <= not (a and b);
    layer2_outputs(6029) <= not b;
    layer2_outputs(6030) <= not b;
    layer2_outputs(6031) <= not a;
    layer2_outputs(6032) <= not b or a;
    layer2_outputs(6033) <= not (a or b);
    layer2_outputs(6034) <= not a;
    layer2_outputs(6035) <= not (a and b);
    layer2_outputs(6036) <= not (a or b);
    layer2_outputs(6037) <= a;
    layer2_outputs(6038) <= not b;
    layer2_outputs(6039) <= not b;
    layer2_outputs(6040) <= b;
    layer2_outputs(6041) <= not a or b;
    layer2_outputs(6042) <= not b or a;
    layer2_outputs(6043) <= b;
    layer2_outputs(6044) <= b and not a;
    layer2_outputs(6045) <= b;
    layer2_outputs(6046) <= a;
    layer2_outputs(6047) <= a;
    layer2_outputs(6048) <= a and b;
    layer2_outputs(6049) <= not a or b;
    layer2_outputs(6050) <= not b;
    layer2_outputs(6051) <= 1'b1;
    layer2_outputs(6052) <= b;
    layer2_outputs(6053) <= b;
    layer2_outputs(6054) <= not (a or b);
    layer2_outputs(6055) <= not (a xor b);
    layer2_outputs(6056) <= a or b;
    layer2_outputs(6057) <= not b or a;
    layer2_outputs(6058) <= b;
    layer2_outputs(6059) <= a and not b;
    layer2_outputs(6060) <= not a;
    layer2_outputs(6061) <= a or b;
    layer2_outputs(6062) <= a;
    layer2_outputs(6063) <= not a;
    layer2_outputs(6064) <= not (a xor b);
    layer2_outputs(6065) <= not b or a;
    layer2_outputs(6066) <= not (a and b);
    layer2_outputs(6067) <= not a or b;
    layer2_outputs(6068) <= not a;
    layer2_outputs(6069) <= a and not b;
    layer2_outputs(6070) <= not a;
    layer2_outputs(6071) <= not b;
    layer2_outputs(6072) <= a and not b;
    layer2_outputs(6073) <= a;
    layer2_outputs(6074) <= not b or a;
    layer2_outputs(6075) <= a and b;
    layer2_outputs(6076) <= not a or b;
    layer2_outputs(6077) <= a or b;
    layer2_outputs(6078) <= a and b;
    layer2_outputs(6079) <= not b;
    layer2_outputs(6080) <= b and not a;
    layer2_outputs(6081) <= not a;
    layer2_outputs(6082) <= not (a and b);
    layer2_outputs(6083) <= not (a and b);
    layer2_outputs(6084) <= not b or a;
    layer2_outputs(6085) <= not a;
    layer2_outputs(6086) <= not (a and b);
    layer2_outputs(6087) <= a xor b;
    layer2_outputs(6088) <= a;
    layer2_outputs(6089) <= not b or a;
    layer2_outputs(6090) <= not (a or b);
    layer2_outputs(6091) <= b;
    layer2_outputs(6092) <= a;
    layer2_outputs(6093) <= not a;
    layer2_outputs(6094) <= not (a xor b);
    layer2_outputs(6095) <= not a;
    layer2_outputs(6096) <= not (a and b);
    layer2_outputs(6097) <= b;
    layer2_outputs(6098) <= not a;
    layer2_outputs(6099) <= not (a xor b);
    layer2_outputs(6100) <= not b;
    layer2_outputs(6101) <= b;
    layer2_outputs(6102) <= a;
    layer2_outputs(6103) <= b and not a;
    layer2_outputs(6104) <= not a or b;
    layer2_outputs(6105) <= b;
    layer2_outputs(6106) <= 1'b0;
    layer2_outputs(6107) <= a;
    layer2_outputs(6108) <= not (a or b);
    layer2_outputs(6109) <= b and not a;
    layer2_outputs(6110) <= not b;
    layer2_outputs(6111) <= not (a or b);
    layer2_outputs(6112) <= a xor b;
    layer2_outputs(6113) <= a and b;
    layer2_outputs(6114) <= not b or a;
    layer2_outputs(6115) <= b;
    layer2_outputs(6116) <= not a;
    layer2_outputs(6117) <= not (a xor b);
    layer2_outputs(6118) <= a and not b;
    layer2_outputs(6119) <= a;
    layer2_outputs(6120) <= b;
    layer2_outputs(6121) <= not a or b;
    layer2_outputs(6122) <= not b;
    layer2_outputs(6123) <= not (a and b);
    layer2_outputs(6124) <= not b;
    layer2_outputs(6125) <= not b;
    layer2_outputs(6126) <= not b;
    layer2_outputs(6127) <= a xor b;
    layer2_outputs(6128) <= a;
    layer2_outputs(6129) <= not a;
    layer2_outputs(6130) <= not (a or b);
    layer2_outputs(6131) <= not b;
    layer2_outputs(6132) <= a;
    layer2_outputs(6133) <= not (a xor b);
    layer2_outputs(6134) <= a or b;
    layer2_outputs(6135) <= not a;
    layer2_outputs(6136) <= not a or b;
    layer2_outputs(6137) <= not b or a;
    layer2_outputs(6138) <= not a;
    layer2_outputs(6139) <= 1'b1;
    layer2_outputs(6140) <= b;
    layer2_outputs(6141) <= a;
    layer2_outputs(6142) <= not (a or b);
    layer2_outputs(6143) <= not a or b;
    layer2_outputs(6144) <= a and not b;
    layer2_outputs(6145) <= b and not a;
    layer2_outputs(6146) <= not b or a;
    layer2_outputs(6147) <= b;
    layer2_outputs(6148) <= not b or a;
    layer2_outputs(6149) <= a;
    layer2_outputs(6150) <= not a;
    layer2_outputs(6151) <= not a;
    layer2_outputs(6152) <= a or b;
    layer2_outputs(6153) <= not (a xor b);
    layer2_outputs(6154) <= not a;
    layer2_outputs(6155) <= not a;
    layer2_outputs(6156) <= a;
    layer2_outputs(6157) <= not a;
    layer2_outputs(6158) <= not (a or b);
    layer2_outputs(6159) <= 1'b0;
    layer2_outputs(6160) <= a or b;
    layer2_outputs(6161) <= b;
    layer2_outputs(6162) <= not a;
    layer2_outputs(6163) <= not a;
    layer2_outputs(6164) <= not b;
    layer2_outputs(6165) <= not b;
    layer2_outputs(6166) <= b and not a;
    layer2_outputs(6167) <= a;
    layer2_outputs(6168) <= not a or b;
    layer2_outputs(6169) <= not b or a;
    layer2_outputs(6170) <= b;
    layer2_outputs(6171) <= a or b;
    layer2_outputs(6172) <= not (a and b);
    layer2_outputs(6173) <= not b;
    layer2_outputs(6174) <= a and not b;
    layer2_outputs(6175) <= not a;
    layer2_outputs(6176) <= not (a and b);
    layer2_outputs(6177) <= not a or b;
    layer2_outputs(6178) <= a and not b;
    layer2_outputs(6179) <= a;
    layer2_outputs(6180) <= a and not b;
    layer2_outputs(6181) <= not (a or b);
    layer2_outputs(6182) <= not b or a;
    layer2_outputs(6183) <= not (a or b);
    layer2_outputs(6184) <= b;
    layer2_outputs(6185) <= not (a or b);
    layer2_outputs(6186) <= a xor b;
    layer2_outputs(6187) <= a and b;
    layer2_outputs(6188) <= not (a xor b);
    layer2_outputs(6189) <= not b or a;
    layer2_outputs(6190) <= b;
    layer2_outputs(6191) <= a and not b;
    layer2_outputs(6192) <= not a or b;
    layer2_outputs(6193) <= not b;
    layer2_outputs(6194) <= not (a or b);
    layer2_outputs(6195) <= not b or a;
    layer2_outputs(6196) <= not b;
    layer2_outputs(6197) <= b;
    layer2_outputs(6198) <= not a;
    layer2_outputs(6199) <= not a;
    layer2_outputs(6200) <= b;
    layer2_outputs(6201) <= b;
    layer2_outputs(6202) <= not (a and b);
    layer2_outputs(6203) <= b;
    layer2_outputs(6204) <= a and not b;
    layer2_outputs(6205) <= not b or a;
    layer2_outputs(6206) <= not a or b;
    layer2_outputs(6207) <= not (a or b);
    layer2_outputs(6208) <= not (a and b);
    layer2_outputs(6209) <= b;
    layer2_outputs(6210) <= b;
    layer2_outputs(6211) <= b;
    layer2_outputs(6212) <= a;
    layer2_outputs(6213) <= not (a or b);
    layer2_outputs(6214) <= not (a or b);
    layer2_outputs(6215) <= b;
    layer2_outputs(6216) <= not a;
    layer2_outputs(6217) <= not a;
    layer2_outputs(6218) <= not b or a;
    layer2_outputs(6219) <= b and not a;
    layer2_outputs(6220) <= not b or a;
    layer2_outputs(6221) <= not a;
    layer2_outputs(6222) <= a xor b;
    layer2_outputs(6223) <= not a;
    layer2_outputs(6224) <= 1'b1;
    layer2_outputs(6225) <= a;
    layer2_outputs(6226) <= not (a or b);
    layer2_outputs(6227) <= b and not a;
    layer2_outputs(6228) <= not b or a;
    layer2_outputs(6229) <= a xor b;
    layer2_outputs(6230) <= a;
    layer2_outputs(6231) <= not a;
    layer2_outputs(6232) <= b and not a;
    layer2_outputs(6233) <= a;
    layer2_outputs(6234) <= b and not a;
    layer2_outputs(6235) <= not a;
    layer2_outputs(6236) <= a;
    layer2_outputs(6237) <= a or b;
    layer2_outputs(6238) <= not b;
    layer2_outputs(6239) <= not b;
    layer2_outputs(6240) <= not a;
    layer2_outputs(6241) <= b and not a;
    layer2_outputs(6242) <= not b or a;
    layer2_outputs(6243) <= not (a xor b);
    layer2_outputs(6244) <= a xor b;
    layer2_outputs(6245) <= a;
    layer2_outputs(6246) <= a;
    layer2_outputs(6247) <= not (a xor b);
    layer2_outputs(6248) <= not a;
    layer2_outputs(6249) <= not b;
    layer2_outputs(6250) <= a and b;
    layer2_outputs(6251) <= not a or b;
    layer2_outputs(6252) <= b and not a;
    layer2_outputs(6253) <= 1'b1;
    layer2_outputs(6254) <= a and not b;
    layer2_outputs(6255) <= not (a xor b);
    layer2_outputs(6256) <= not (a xor b);
    layer2_outputs(6257) <= not a;
    layer2_outputs(6258) <= a xor b;
    layer2_outputs(6259) <= a or b;
    layer2_outputs(6260) <= not b;
    layer2_outputs(6261) <= a;
    layer2_outputs(6262) <= not (a and b);
    layer2_outputs(6263) <= not (a and b);
    layer2_outputs(6264) <= b;
    layer2_outputs(6265) <= a or b;
    layer2_outputs(6266) <= a xor b;
    layer2_outputs(6267) <= b and not a;
    layer2_outputs(6268) <= not (a xor b);
    layer2_outputs(6269) <= a and b;
    layer2_outputs(6270) <= not (a and b);
    layer2_outputs(6271) <= b;
    layer2_outputs(6272) <= not a;
    layer2_outputs(6273) <= b;
    layer2_outputs(6274) <= a or b;
    layer2_outputs(6275) <= b;
    layer2_outputs(6276) <= a or b;
    layer2_outputs(6277) <= not b;
    layer2_outputs(6278) <= a and b;
    layer2_outputs(6279) <= a and not b;
    layer2_outputs(6280) <= a and not b;
    layer2_outputs(6281) <= not b;
    layer2_outputs(6282) <= not (a xor b);
    layer2_outputs(6283) <= a;
    layer2_outputs(6284) <= not a;
    layer2_outputs(6285) <= not (a xor b);
    layer2_outputs(6286) <= b;
    layer2_outputs(6287) <= not a;
    layer2_outputs(6288) <= b;
    layer2_outputs(6289) <= not (a and b);
    layer2_outputs(6290) <= a;
    layer2_outputs(6291) <= b;
    layer2_outputs(6292) <= not b or a;
    layer2_outputs(6293) <= b;
    layer2_outputs(6294) <= a xor b;
    layer2_outputs(6295) <= not a or b;
    layer2_outputs(6296) <= not a;
    layer2_outputs(6297) <= not b;
    layer2_outputs(6298) <= not (a and b);
    layer2_outputs(6299) <= a and b;
    layer2_outputs(6300) <= a;
    layer2_outputs(6301) <= 1'b0;
    layer2_outputs(6302) <= a xor b;
    layer2_outputs(6303) <= a or b;
    layer2_outputs(6304) <= not (a and b);
    layer2_outputs(6305) <= 1'b1;
    layer2_outputs(6306) <= a;
    layer2_outputs(6307) <= not b or a;
    layer2_outputs(6308) <= not b;
    layer2_outputs(6309) <= 1'b1;
    layer2_outputs(6310) <= b and not a;
    layer2_outputs(6311) <= a xor b;
    layer2_outputs(6312) <= not b;
    layer2_outputs(6313) <= b;
    layer2_outputs(6314) <= not a or b;
    layer2_outputs(6315) <= not b;
    layer2_outputs(6316) <= a or b;
    layer2_outputs(6317) <= not a;
    layer2_outputs(6318) <= a and b;
    layer2_outputs(6319) <= a;
    layer2_outputs(6320) <= b and not a;
    layer2_outputs(6321) <= not b;
    layer2_outputs(6322) <= a and b;
    layer2_outputs(6323) <= b and not a;
    layer2_outputs(6324) <= not a;
    layer2_outputs(6325) <= a or b;
    layer2_outputs(6326) <= a xor b;
    layer2_outputs(6327) <= b;
    layer2_outputs(6328) <= a and not b;
    layer2_outputs(6329) <= a and not b;
    layer2_outputs(6330) <= b;
    layer2_outputs(6331) <= not b or a;
    layer2_outputs(6332) <= a and not b;
    layer2_outputs(6333) <= not (a and b);
    layer2_outputs(6334) <= a;
    layer2_outputs(6335) <= not (a or b);
    layer2_outputs(6336) <= not a;
    layer2_outputs(6337) <= not a or b;
    layer2_outputs(6338) <= not a or b;
    layer2_outputs(6339) <= not (a and b);
    layer2_outputs(6340) <= a;
    layer2_outputs(6341) <= not (a and b);
    layer2_outputs(6342) <= not b or a;
    layer2_outputs(6343) <= not (a xor b);
    layer2_outputs(6344) <= not b;
    layer2_outputs(6345) <= not b;
    layer2_outputs(6346) <= not (a xor b);
    layer2_outputs(6347) <= b;
    layer2_outputs(6348) <= not (a and b);
    layer2_outputs(6349) <= a xor b;
    layer2_outputs(6350) <= a;
    layer2_outputs(6351) <= not a;
    layer2_outputs(6352) <= not (a and b);
    layer2_outputs(6353) <= not b or a;
    layer2_outputs(6354) <= a and not b;
    layer2_outputs(6355) <= not (a or b);
    layer2_outputs(6356) <= not a;
    layer2_outputs(6357) <= not a;
    layer2_outputs(6358) <= a and b;
    layer2_outputs(6359) <= b;
    layer2_outputs(6360) <= not (a xor b);
    layer2_outputs(6361) <= a xor b;
    layer2_outputs(6362) <= not a or b;
    layer2_outputs(6363) <= b;
    layer2_outputs(6364) <= a and b;
    layer2_outputs(6365) <= a and b;
    layer2_outputs(6366) <= a or b;
    layer2_outputs(6367) <= not (a and b);
    layer2_outputs(6368) <= 1'b1;
    layer2_outputs(6369) <= not b;
    layer2_outputs(6370) <= not b or a;
    layer2_outputs(6371) <= a and not b;
    layer2_outputs(6372) <= b;
    layer2_outputs(6373) <= a or b;
    layer2_outputs(6374) <= a and b;
    layer2_outputs(6375) <= not b;
    layer2_outputs(6376) <= not b or a;
    layer2_outputs(6377) <= a;
    layer2_outputs(6378) <= a;
    layer2_outputs(6379) <= not (a or b);
    layer2_outputs(6380) <= not (a or b);
    layer2_outputs(6381) <= not b;
    layer2_outputs(6382) <= not b or a;
    layer2_outputs(6383) <= a and not b;
    layer2_outputs(6384) <= a;
    layer2_outputs(6385) <= b and not a;
    layer2_outputs(6386) <= not a;
    layer2_outputs(6387) <= not a or b;
    layer2_outputs(6388) <= b;
    layer2_outputs(6389) <= a or b;
    layer2_outputs(6390) <= not (a or b);
    layer2_outputs(6391) <= a or b;
    layer2_outputs(6392) <= not a or b;
    layer2_outputs(6393) <= 1'b1;
    layer2_outputs(6394) <= b;
    layer2_outputs(6395) <= a and b;
    layer2_outputs(6396) <= not b or a;
    layer2_outputs(6397) <= a;
    layer2_outputs(6398) <= not (a xor b);
    layer2_outputs(6399) <= not (a xor b);
    layer2_outputs(6400) <= not (a or b);
    layer2_outputs(6401) <= not a;
    layer2_outputs(6402) <= not (a xor b);
    layer2_outputs(6403) <= a and not b;
    layer2_outputs(6404) <= not (a xor b);
    layer2_outputs(6405) <= not a;
    layer2_outputs(6406) <= b and not a;
    layer2_outputs(6407) <= not (a and b);
    layer2_outputs(6408) <= not a;
    layer2_outputs(6409) <= b and not a;
    layer2_outputs(6410) <= a and b;
    layer2_outputs(6411) <= not b or a;
    layer2_outputs(6412) <= not b;
    layer2_outputs(6413) <= not a;
    layer2_outputs(6414) <= a and not b;
    layer2_outputs(6415) <= a;
    layer2_outputs(6416) <= not a or b;
    layer2_outputs(6417) <= a;
    layer2_outputs(6418) <= not (a or b);
    layer2_outputs(6419) <= a and b;
    layer2_outputs(6420) <= a;
    layer2_outputs(6421) <= a;
    layer2_outputs(6422) <= b;
    layer2_outputs(6423) <= not b;
    layer2_outputs(6424) <= a or b;
    layer2_outputs(6425) <= not (a and b);
    layer2_outputs(6426) <= b;
    layer2_outputs(6427) <= b;
    layer2_outputs(6428) <= not b;
    layer2_outputs(6429) <= not b;
    layer2_outputs(6430) <= not b;
    layer2_outputs(6431) <= not (a and b);
    layer2_outputs(6432) <= a and b;
    layer2_outputs(6433) <= not a;
    layer2_outputs(6434) <= a;
    layer2_outputs(6435) <= not (a or b);
    layer2_outputs(6436) <= not a;
    layer2_outputs(6437) <= a or b;
    layer2_outputs(6438) <= a or b;
    layer2_outputs(6439) <= b;
    layer2_outputs(6440) <= not a or b;
    layer2_outputs(6441) <= a and b;
    layer2_outputs(6442) <= not a or b;
    layer2_outputs(6443) <= b;
    layer2_outputs(6444) <= not a;
    layer2_outputs(6445) <= a and b;
    layer2_outputs(6446) <= 1'b0;
    layer2_outputs(6447) <= b;
    layer2_outputs(6448) <= not (a and b);
    layer2_outputs(6449) <= not b;
    layer2_outputs(6450) <= not a or b;
    layer2_outputs(6451) <= b;
    layer2_outputs(6452) <= a;
    layer2_outputs(6453) <= 1'b0;
    layer2_outputs(6454) <= not b or a;
    layer2_outputs(6455) <= a and b;
    layer2_outputs(6456) <= a and not b;
    layer2_outputs(6457) <= not (a or b);
    layer2_outputs(6458) <= not a;
    layer2_outputs(6459) <= a and not b;
    layer2_outputs(6460) <= a or b;
    layer2_outputs(6461) <= a or b;
    layer2_outputs(6462) <= a and b;
    layer2_outputs(6463) <= a and b;
    layer2_outputs(6464) <= not a or b;
    layer2_outputs(6465) <= not b or a;
    layer2_outputs(6466) <= not b;
    layer2_outputs(6467) <= 1'b0;
    layer2_outputs(6468) <= a xor b;
    layer2_outputs(6469) <= b and not a;
    layer2_outputs(6470) <= a and b;
    layer2_outputs(6471) <= not b or a;
    layer2_outputs(6472) <= a and not b;
    layer2_outputs(6473) <= not a;
    layer2_outputs(6474) <= a and not b;
    layer2_outputs(6475) <= b and not a;
    layer2_outputs(6476) <= not a;
    layer2_outputs(6477) <= 1'b0;
    layer2_outputs(6478) <= a;
    layer2_outputs(6479) <= not b;
    layer2_outputs(6480) <= not (a xor b);
    layer2_outputs(6481) <= not (a xor b);
    layer2_outputs(6482) <= a and not b;
    layer2_outputs(6483) <= b;
    layer2_outputs(6484) <= a or b;
    layer2_outputs(6485) <= b;
    layer2_outputs(6486) <= not b or a;
    layer2_outputs(6487) <= b and not a;
    layer2_outputs(6488) <= a and not b;
    layer2_outputs(6489) <= a;
    layer2_outputs(6490) <= not (a xor b);
    layer2_outputs(6491) <= not a or b;
    layer2_outputs(6492) <= a or b;
    layer2_outputs(6493) <= not (a or b);
    layer2_outputs(6494) <= not (a and b);
    layer2_outputs(6495) <= not b or a;
    layer2_outputs(6496) <= not a or b;
    layer2_outputs(6497) <= 1'b0;
    layer2_outputs(6498) <= a or b;
    layer2_outputs(6499) <= a;
    layer2_outputs(6500) <= 1'b0;
    layer2_outputs(6501) <= not a;
    layer2_outputs(6502) <= not b or a;
    layer2_outputs(6503) <= b;
    layer2_outputs(6504) <= a and b;
    layer2_outputs(6505) <= not a;
    layer2_outputs(6506) <= not a;
    layer2_outputs(6507) <= not a or b;
    layer2_outputs(6508) <= a;
    layer2_outputs(6509) <= not (a or b);
    layer2_outputs(6510) <= a and b;
    layer2_outputs(6511) <= a;
    layer2_outputs(6512) <= a and b;
    layer2_outputs(6513) <= not (a or b);
    layer2_outputs(6514) <= not (a xor b);
    layer2_outputs(6515) <= a xor b;
    layer2_outputs(6516) <= a xor b;
    layer2_outputs(6517) <= b;
    layer2_outputs(6518) <= a and b;
    layer2_outputs(6519) <= not a;
    layer2_outputs(6520) <= b;
    layer2_outputs(6521) <= not a or b;
    layer2_outputs(6522) <= not (a and b);
    layer2_outputs(6523) <= not b;
    layer2_outputs(6524) <= not a;
    layer2_outputs(6525) <= not b or a;
    layer2_outputs(6526) <= a;
    layer2_outputs(6527) <= 1'b1;
    layer2_outputs(6528) <= not a;
    layer2_outputs(6529) <= a xor b;
    layer2_outputs(6530) <= a or b;
    layer2_outputs(6531) <= b;
    layer2_outputs(6532) <= b and not a;
    layer2_outputs(6533) <= not a or b;
    layer2_outputs(6534) <= not b;
    layer2_outputs(6535) <= a and not b;
    layer2_outputs(6536) <= a xor b;
    layer2_outputs(6537) <= not b;
    layer2_outputs(6538) <= 1'b0;
    layer2_outputs(6539) <= not a or b;
    layer2_outputs(6540) <= a or b;
    layer2_outputs(6541) <= not (a and b);
    layer2_outputs(6542) <= not a;
    layer2_outputs(6543) <= not a;
    layer2_outputs(6544) <= a xor b;
    layer2_outputs(6545) <= a and b;
    layer2_outputs(6546) <= a or b;
    layer2_outputs(6547) <= not (a and b);
    layer2_outputs(6548) <= not (a and b);
    layer2_outputs(6549) <= not b;
    layer2_outputs(6550) <= a and not b;
    layer2_outputs(6551) <= a or b;
    layer2_outputs(6552) <= not b;
    layer2_outputs(6553) <= a and b;
    layer2_outputs(6554) <= not a or b;
    layer2_outputs(6555) <= not b;
    layer2_outputs(6556) <= 1'b1;
    layer2_outputs(6557) <= a and not b;
    layer2_outputs(6558) <= not (a xor b);
    layer2_outputs(6559) <= a;
    layer2_outputs(6560) <= b;
    layer2_outputs(6561) <= 1'b1;
    layer2_outputs(6562) <= not (a and b);
    layer2_outputs(6563) <= not b or a;
    layer2_outputs(6564) <= not b;
    layer2_outputs(6565) <= b and not a;
    layer2_outputs(6566) <= a and not b;
    layer2_outputs(6567) <= not a;
    layer2_outputs(6568) <= not (a xor b);
    layer2_outputs(6569) <= not (a and b);
    layer2_outputs(6570) <= a or b;
    layer2_outputs(6571) <= a and not b;
    layer2_outputs(6572) <= not a;
    layer2_outputs(6573) <= not a or b;
    layer2_outputs(6574) <= 1'b1;
    layer2_outputs(6575) <= not b or a;
    layer2_outputs(6576) <= b;
    layer2_outputs(6577) <= not a or b;
    layer2_outputs(6578) <= a and not b;
    layer2_outputs(6579) <= a xor b;
    layer2_outputs(6580) <= b;
    layer2_outputs(6581) <= a and b;
    layer2_outputs(6582) <= not (a or b);
    layer2_outputs(6583) <= not a;
    layer2_outputs(6584) <= not a;
    layer2_outputs(6585) <= not (a or b);
    layer2_outputs(6586) <= a;
    layer2_outputs(6587) <= not a;
    layer2_outputs(6588) <= not b;
    layer2_outputs(6589) <= a xor b;
    layer2_outputs(6590) <= 1'b0;
    layer2_outputs(6591) <= b;
    layer2_outputs(6592) <= a;
    layer2_outputs(6593) <= a or b;
    layer2_outputs(6594) <= not a;
    layer2_outputs(6595) <= b;
    layer2_outputs(6596) <= not b;
    layer2_outputs(6597) <= b;
    layer2_outputs(6598) <= a;
    layer2_outputs(6599) <= a and not b;
    layer2_outputs(6600) <= not b;
    layer2_outputs(6601) <= not a;
    layer2_outputs(6602) <= b;
    layer2_outputs(6603) <= a;
    layer2_outputs(6604) <= a and not b;
    layer2_outputs(6605) <= not a;
    layer2_outputs(6606) <= b and not a;
    layer2_outputs(6607) <= not (a xor b);
    layer2_outputs(6608) <= a and not b;
    layer2_outputs(6609) <= a xor b;
    layer2_outputs(6610) <= not (a or b);
    layer2_outputs(6611) <= a and b;
    layer2_outputs(6612) <= not b;
    layer2_outputs(6613) <= b;
    layer2_outputs(6614) <= a;
    layer2_outputs(6615) <= a;
    layer2_outputs(6616) <= not b;
    layer2_outputs(6617) <= a;
    layer2_outputs(6618) <= not b or a;
    layer2_outputs(6619) <= b;
    layer2_outputs(6620) <= a or b;
    layer2_outputs(6621) <= not (a and b);
    layer2_outputs(6622) <= b;
    layer2_outputs(6623) <= a or b;
    layer2_outputs(6624) <= not a or b;
    layer2_outputs(6625) <= not (a or b);
    layer2_outputs(6626) <= not (a or b);
    layer2_outputs(6627) <= b and not a;
    layer2_outputs(6628) <= not b;
    layer2_outputs(6629) <= a and b;
    layer2_outputs(6630) <= a and b;
    layer2_outputs(6631) <= not b or a;
    layer2_outputs(6632) <= a and b;
    layer2_outputs(6633) <= not b;
    layer2_outputs(6634) <= 1'b1;
    layer2_outputs(6635) <= not b;
    layer2_outputs(6636) <= not b;
    layer2_outputs(6637) <= not (a and b);
    layer2_outputs(6638) <= a or b;
    layer2_outputs(6639) <= 1'b1;
    layer2_outputs(6640) <= not (a xor b);
    layer2_outputs(6641) <= b;
    layer2_outputs(6642) <= not b or a;
    layer2_outputs(6643) <= a;
    layer2_outputs(6644) <= 1'b0;
    layer2_outputs(6645) <= a;
    layer2_outputs(6646) <= not (a or b);
    layer2_outputs(6647) <= a and not b;
    layer2_outputs(6648) <= a and not b;
    layer2_outputs(6649) <= not (a xor b);
    layer2_outputs(6650) <= not b or a;
    layer2_outputs(6651) <= a;
    layer2_outputs(6652) <= b;
    layer2_outputs(6653) <= not a;
    layer2_outputs(6654) <= a;
    layer2_outputs(6655) <= b;
    layer2_outputs(6656) <= not b or a;
    layer2_outputs(6657) <= b;
    layer2_outputs(6658) <= not (a and b);
    layer2_outputs(6659) <= not (a and b);
    layer2_outputs(6660) <= b and not a;
    layer2_outputs(6661) <= b;
    layer2_outputs(6662) <= a and b;
    layer2_outputs(6663) <= not (a xor b);
    layer2_outputs(6664) <= not b;
    layer2_outputs(6665) <= not a;
    layer2_outputs(6666) <= not b or a;
    layer2_outputs(6667) <= b and not a;
    layer2_outputs(6668) <= a;
    layer2_outputs(6669) <= a;
    layer2_outputs(6670) <= not (a and b);
    layer2_outputs(6671) <= a and b;
    layer2_outputs(6672) <= a xor b;
    layer2_outputs(6673) <= a and b;
    layer2_outputs(6674) <= not b;
    layer2_outputs(6675) <= not b;
    layer2_outputs(6676) <= b and not a;
    layer2_outputs(6677) <= not (a xor b);
    layer2_outputs(6678) <= b;
    layer2_outputs(6679) <= a or b;
    layer2_outputs(6680) <= not a;
    layer2_outputs(6681) <= a or b;
    layer2_outputs(6682) <= a;
    layer2_outputs(6683) <= b and not a;
    layer2_outputs(6684) <= b;
    layer2_outputs(6685) <= not b or a;
    layer2_outputs(6686) <= not b;
    layer2_outputs(6687) <= not b or a;
    layer2_outputs(6688) <= 1'b1;
    layer2_outputs(6689) <= 1'b1;
    layer2_outputs(6690) <= not b;
    layer2_outputs(6691) <= not b;
    layer2_outputs(6692) <= a and not b;
    layer2_outputs(6693) <= a xor b;
    layer2_outputs(6694) <= not b;
    layer2_outputs(6695) <= b;
    layer2_outputs(6696) <= a and not b;
    layer2_outputs(6697) <= a;
    layer2_outputs(6698) <= not b or a;
    layer2_outputs(6699) <= a;
    layer2_outputs(6700) <= not b or a;
    layer2_outputs(6701) <= a or b;
    layer2_outputs(6702) <= not b;
    layer2_outputs(6703) <= b;
    layer2_outputs(6704) <= not a or b;
    layer2_outputs(6705) <= not a;
    layer2_outputs(6706) <= b;
    layer2_outputs(6707) <= a;
    layer2_outputs(6708) <= a and not b;
    layer2_outputs(6709) <= a and not b;
    layer2_outputs(6710) <= not b;
    layer2_outputs(6711) <= not a or b;
    layer2_outputs(6712) <= not b;
    layer2_outputs(6713) <= not a;
    layer2_outputs(6714) <= b;
    layer2_outputs(6715) <= not (a or b);
    layer2_outputs(6716) <= not (a and b);
    layer2_outputs(6717) <= not (a or b);
    layer2_outputs(6718) <= a and b;
    layer2_outputs(6719) <= a;
    layer2_outputs(6720) <= b and not a;
    layer2_outputs(6721) <= not a;
    layer2_outputs(6722) <= not b;
    layer2_outputs(6723) <= not b or a;
    layer2_outputs(6724) <= not (a xor b);
    layer2_outputs(6725) <= not a;
    layer2_outputs(6726) <= b;
    layer2_outputs(6727) <= 1'b1;
    layer2_outputs(6728) <= not b;
    layer2_outputs(6729) <= not (a or b);
    layer2_outputs(6730) <= a and b;
    layer2_outputs(6731) <= not b;
    layer2_outputs(6732) <= a xor b;
    layer2_outputs(6733) <= not a or b;
    layer2_outputs(6734) <= b;
    layer2_outputs(6735) <= a xor b;
    layer2_outputs(6736) <= not a;
    layer2_outputs(6737) <= a;
    layer2_outputs(6738) <= not b or a;
    layer2_outputs(6739) <= a and not b;
    layer2_outputs(6740) <= not (a and b);
    layer2_outputs(6741) <= not a;
    layer2_outputs(6742) <= a or b;
    layer2_outputs(6743) <= b;
    layer2_outputs(6744) <= not a;
    layer2_outputs(6745) <= not a;
    layer2_outputs(6746) <= a and not b;
    layer2_outputs(6747) <= not a or b;
    layer2_outputs(6748) <= not (a and b);
    layer2_outputs(6749) <= a;
    layer2_outputs(6750) <= a and b;
    layer2_outputs(6751) <= a and b;
    layer2_outputs(6752) <= not a;
    layer2_outputs(6753) <= a and not b;
    layer2_outputs(6754) <= 1'b0;
    layer2_outputs(6755) <= a or b;
    layer2_outputs(6756) <= b and not a;
    layer2_outputs(6757) <= b and not a;
    layer2_outputs(6758) <= not a;
    layer2_outputs(6759) <= not a or b;
    layer2_outputs(6760) <= not b;
    layer2_outputs(6761) <= a or b;
    layer2_outputs(6762) <= not b or a;
    layer2_outputs(6763) <= not (a xor b);
    layer2_outputs(6764) <= a xor b;
    layer2_outputs(6765) <= not (a and b);
    layer2_outputs(6766) <= b and not a;
    layer2_outputs(6767) <= a;
    layer2_outputs(6768) <= a or b;
    layer2_outputs(6769) <= b and not a;
    layer2_outputs(6770) <= a or b;
    layer2_outputs(6771) <= a or b;
    layer2_outputs(6772) <= a;
    layer2_outputs(6773) <= not (a xor b);
    layer2_outputs(6774) <= not a or b;
    layer2_outputs(6775) <= 1'b0;
    layer2_outputs(6776) <= not b;
    layer2_outputs(6777) <= not (a and b);
    layer2_outputs(6778) <= a and b;
    layer2_outputs(6779) <= a and b;
    layer2_outputs(6780) <= b;
    layer2_outputs(6781) <= b and not a;
    layer2_outputs(6782) <= a;
    layer2_outputs(6783) <= b;
    layer2_outputs(6784) <= not b;
    layer2_outputs(6785) <= not b or a;
    layer2_outputs(6786) <= a;
    layer2_outputs(6787) <= not (a and b);
    layer2_outputs(6788) <= a;
    layer2_outputs(6789) <= not (a xor b);
    layer2_outputs(6790) <= not a or b;
    layer2_outputs(6791) <= a;
    layer2_outputs(6792) <= not b or a;
    layer2_outputs(6793) <= not (a or b);
    layer2_outputs(6794) <= not a or b;
    layer2_outputs(6795) <= b;
    layer2_outputs(6796) <= not a;
    layer2_outputs(6797) <= b;
    layer2_outputs(6798) <= a or b;
    layer2_outputs(6799) <= a;
    layer2_outputs(6800) <= not (a and b);
    layer2_outputs(6801) <= not b;
    layer2_outputs(6802) <= not (a and b);
    layer2_outputs(6803) <= a and b;
    layer2_outputs(6804) <= b;
    layer2_outputs(6805) <= a or b;
    layer2_outputs(6806) <= a and not b;
    layer2_outputs(6807) <= a or b;
    layer2_outputs(6808) <= a;
    layer2_outputs(6809) <= b;
    layer2_outputs(6810) <= b;
    layer2_outputs(6811) <= b;
    layer2_outputs(6812) <= b;
    layer2_outputs(6813) <= a;
    layer2_outputs(6814) <= not b;
    layer2_outputs(6815) <= b and not a;
    layer2_outputs(6816) <= b;
    layer2_outputs(6817) <= not a;
    layer2_outputs(6818) <= not b or a;
    layer2_outputs(6819) <= not a;
    layer2_outputs(6820) <= not (a and b);
    layer2_outputs(6821) <= b;
    layer2_outputs(6822) <= not a;
    layer2_outputs(6823) <= not a;
    layer2_outputs(6824) <= a xor b;
    layer2_outputs(6825) <= a;
    layer2_outputs(6826) <= a and b;
    layer2_outputs(6827) <= a and not b;
    layer2_outputs(6828) <= not b;
    layer2_outputs(6829) <= a and b;
    layer2_outputs(6830) <= not (a xor b);
    layer2_outputs(6831) <= not a or b;
    layer2_outputs(6832) <= a xor b;
    layer2_outputs(6833) <= a or b;
    layer2_outputs(6834) <= not (a xor b);
    layer2_outputs(6835) <= a and b;
    layer2_outputs(6836) <= not a or b;
    layer2_outputs(6837) <= not a;
    layer2_outputs(6838) <= 1'b0;
    layer2_outputs(6839) <= not (a or b);
    layer2_outputs(6840) <= not b;
    layer2_outputs(6841) <= a and b;
    layer2_outputs(6842) <= not (a and b);
    layer2_outputs(6843) <= b;
    layer2_outputs(6844) <= not b or a;
    layer2_outputs(6845) <= not (a and b);
    layer2_outputs(6846) <= a or b;
    layer2_outputs(6847) <= a and not b;
    layer2_outputs(6848) <= 1'b0;
    layer2_outputs(6849) <= not b or a;
    layer2_outputs(6850) <= b;
    layer2_outputs(6851) <= not b;
    layer2_outputs(6852) <= b;
    layer2_outputs(6853) <= a;
    layer2_outputs(6854) <= not a or b;
    layer2_outputs(6855) <= not a or b;
    layer2_outputs(6856) <= not a;
    layer2_outputs(6857) <= not (a and b);
    layer2_outputs(6858) <= a or b;
    layer2_outputs(6859) <= a;
    layer2_outputs(6860) <= b;
    layer2_outputs(6861) <= a and b;
    layer2_outputs(6862) <= b;
    layer2_outputs(6863) <= b and not a;
    layer2_outputs(6864) <= not (a and b);
    layer2_outputs(6865) <= not b;
    layer2_outputs(6866) <= not (a and b);
    layer2_outputs(6867) <= a;
    layer2_outputs(6868) <= not a;
    layer2_outputs(6869) <= not (a and b);
    layer2_outputs(6870) <= not b;
    layer2_outputs(6871) <= b;
    layer2_outputs(6872) <= a and not b;
    layer2_outputs(6873) <= not b;
    layer2_outputs(6874) <= b and not a;
    layer2_outputs(6875) <= a and not b;
    layer2_outputs(6876) <= b and not a;
    layer2_outputs(6877) <= 1'b1;
    layer2_outputs(6878) <= not a or b;
    layer2_outputs(6879) <= b;
    layer2_outputs(6880) <= b;
    layer2_outputs(6881) <= not (a or b);
    layer2_outputs(6882) <= not b or a;
    layer2_outputs(6883) <= b and not a;
    layer2_outputs(6884) <= not (a xor b);
    layer2_outputs(6885) <= a xor b;
    layer2_outputs(6886) <= a or b;
    layer2_outputs(6887) <= b;
    layer2_outputs(6888) <= a;
    layer2_outputs(6889) <= not a or b;
    layer2_outputs(6890) <= b;
    layer2_outputs(6891) <= not b or a;
    layer2_outputs(6892) <= not b;
    layer2_outputs(6893) <= 1'b0;
    layer2_outputs(6894) <= not b;
    layer2_outputs(6895) <= 1'b1;
    layer2_outputs(6896) <= a;
    layer2_outputs(6897) <= b;
    layer2_outputs(6898) <= a and not b;
    layer2_outputs(6899) <= 1'b1;
    layer2_outputs(6900) <= a or b;
    layer2_outputs(6901) <= not (a and b);
    layer2_outputs(6902) <= not a;
    layer2_outputs(6903) <= not a or b;
    layer2_outputs(6904) <= not (a and b);
    layer2_outputs(6905) <= a;
    layer2_outputs(6906) <= not b or a;
    layer2_outputs(6907) <= a;
    layer2_outputs(6908) <= b and not a;
    layer2_outputs(6909) <= not b;
    layer2_outputs(6910) <= a;
    layer2_outputs(6911) <= not (a or b);
    layer2_outputs(6912) <= not b;
    layer2_outputs(6913) <= b;
    layer2_outputs(6914) <= not a or b;
    layer2_outputs(6915) <= a or b;
    layer2_outputs(6916) <= a xor b;
    layer2_outputs(6917) <= a xor b;
    layer2_outputs(6918) <= not a;
    layer2_outputs(6919) <= a xor b;
    layer2_outputs(6920) <= not (a or b);
    layer2_outputs(6921) <= b and not a;
    layer2_outputs(6922) <= not (a or b);
    layer2_outputs(6923) <= b and not a;
    layer2_outputs(6924) <= not b;
    layer2_outputs(6925) <= not a or b;
    layer2_outputs(6926) <= not (a and b);
    layer2_outputs(6927) <= a;
    layer2_outputs(6928) <= not a or b;
    layer2_outputs(6929) <= 1'b0;
    layer2_outputs(6930) <= a;
    layer2_outputs(6931) <= b;
    layer2_outputs(6932) <= b;
    layer2_outputs(6933) <= b;
    layer2_outputs(6934) <= 1'b1;
    layer2_outputs(6935) <= not (a xor b);
    layer2_outputs(6936) <= 1'b0;
    layer2_outputs(6937) <= a xor b;
    layer2_outputs(6938) <= not (a or b);
    layer2_outputs(6939) <= a;
    layer2_outputs(6940) <= 1'b0;
    layer2_outputs(6941) <= 1'b0;
    layer2_outputs(6942) <= not (a and b);
    layer2_outputs(6943) <= 1'b1;
    layer2_outputs(6944) <= not a;
    layer2_outputs(6945) <= b;
    layer2_outputs(6946) <= a xor b;
    layer2_outputs(6947) <= b;
    layer2_outputs(6948) <= not a;
    layer2_outputs(6949) <= not (a xor b);
    layer2_outputs(6950) <= a and b;
    layer2_outputs(6951) <= 1'b1;
    layer2_outputs(6952) <= not (a and b);
    layer2_outputs(6953) <= not (a and b);
    layer2_outputs(6954) <= a and b;
    layer2_outputs(6955) <= not a;
    layer2_outputs(6956) <= a and not b;
    layer2_outputs(6957) <= a and b;
    layer2_outputs(6958) <= 1'b1;
    layer2_outputs(6959) <= a xor b;
    layer2_outputs(6960) <= not (a and b);
    layer2_outputs(6961) <= not b;
    layer2_outputs(6962) <= not b;
    layer2_outputs(6963) <= not b;
    layer2_outputs(6964) <= a and not b;
    layer2_outputs(6965) <= not b;
    layer2_outputs(6966) <= not (a or b);
    layer2_outputs(6967) <= not b or a;
    layer2_outputs(6968) <= b;
    layer2_outputs(6969) <= not b;
    layer2_outputs(6970) <= not (a or b);
    layer2_outputs(6971) <= not b or a;
    layer2_outputs(6972) <= a and not b;
    layer2_outputs(6973) <= b;
    layer2_outputs(6974) <= not a;
    layer2_outputs(6975) <= not b or a;
    layer2_outputs(6976) <= not (a and b);
    layer2_outputs(6977) <= a or b;
    layer2_outputs(6978) <= a or b;
    layer2_outputs(6979) <= not a;
    layer2_outputs(6980) <= not (a xor b);
    layer2_outputs(6981) <= b;
    layer2_outputs(6982) <= not b or a;
    layer2_outputs(6983) <= a;
    layer2_outputs(6984) <= a or b;
    layer2_outputs(6985) <= not a;
    layer2_outputs(6986) <= b and not a;
    layer2_outputs(6987) <= b and not a;
    layer2_outputs(6988) <= not a or b;
    layer2_outputs(6989) <= a or b;
    layer2_outputs(6990) <= not (a xor b);
    layer2_outputs(6991) <= a xor b;
    layer2_outputs(6992) <= not b;
    layer2_outputs(6993) <= b;
    layer2_outputs(6994) <= not b;
    layer2_outputs(6995) <= not a or b;
    layer2_outputs(6996) <= b;
    layer2_outputs(6997) <= not b or a;
    layer2_outputs(6998) <= not a;
    layer2_outputs(6999) <= a and b;
    layer2_outputs(7000) <= b and not a;
    layer2_outputs(7001) <= not a;
    layer2_outputs(7002) <= not a;
    layer2_outputs(7003) <= not b or a;
    layer2_outputs(7004) <= not b;
    layer2_outputs(7005) <= a and not b;
    layer2_outputs(7006) <= b and not a;
    layer2_outputs(7007) <= a and not b;
    layer2_outputs(7008) <= 1'b1;
    layer2_outputs(7009) <= a and not b;
    layer2_outputs(7010) <= not a;
    layer2_outputs(7011) <= 1'b0;
    layer2_outputs(7012) <= not a;
    layer2_outputs(7013) <= a xor b;
    layer2_outputs(7014) <= not (a and b);
    layer2_outputs(7015) <= a or b;
    layer2_outputs(7016) <= not a;
    layer2_outputs(7017) <= not (a xor b);
    layer2_outputs(7018) <= a or b;
    layer2_outputs(7019) <= b;
    layer2_outputs(7020) <= a and b;
    layer2_outputs(7021) <= a and not b;
    layer2_outputs(7022) <= a or b;
    layer2_outputs(7023) <= not b;
    layer2_outputs(7024) <= not b;
    layer2_outputs(7025) <= not b;
    layer2_outputs(7026) <= not a;
    layer2_outputs(7027) <= not b;
    layer2_outputs(7028) <= not b or a;
    layer2_outputs(7029) <= not b;
    layer2_outputs(7030) <= b;
    layer2_outputs(7031) <= a;
    layer2_outputs(7032) <= a;
    layer2_outputs(7033) <= not a;
    layer2_outputs(7034) <= a;
    layer2_outputs(7035) <= not b;
    layer2_outputs(7036) <= not (a xor b);
    layer2_outputs(7037) <= not a;
    layer2_outputs(7038) <= a;
    layer2_outputs(7039) <= not a or b;
    layer2_outputs(7040) <= a and not b;
    layer2_outputs(7041) <= a and b;
    layer2_outputs(7042) <= not a or b;
    layer2_outputs(7043) <= 1'b1;
    layer2_outputs(7044) <= 1'b0;
    layer2_outputs(7045) <= not (a xor b);
    layer2_outputs(7046) <= not a;
    layer2_outputs(7047) <= a and b;
    layer2_outputs(7048) <= not a;
    layer2_outputs(7049) <= a or b;
    layer2_outputs(7050) <= not b;
    layer2_outputs(7051) <= b;
    layer2_outputs(7052) <= not b;
    layer2_outputs(7053) <= not b or a;
    layer2_outputs(7054) <= b and not a;
    layer2_outputs(7055) <= not (a and b);
    layer2_outputs(7056) <= b;
    layer2_outputs(7057) <= not a;
    layer2_outputs(7058) <= not b;
    layer2_outputs(7059) <= b;
    layer2_outputs(7060) <= a and not b;
    layer2_outputs(7061) <= not (a xor b);
    layer2_outputs(7062) <= a and b;
    layer2_outputs(7063) <= not (a or b);
    layer2_outputs(7064) <= not (a or b);
    layer2_outputs(7065) <= a and b;
    layer2_outputs(7066) <= not (a and b);
    layer2_outputs(7067) <= a or b;
    layer2_outputs(7068) <= a xor b;
    layer2_outputs(7069) <= not (a xor b);
    layer2_outputs(7070) <= not b or a;
    layer2_outputs(7071) <= not (a and b);
    layer2_outputs(7072) <= not b;
    layer2_outputs(7073) <= a and b;
    layer2_outputs(7074) <= b;
    layer2_outputs(7075) <= a or b;
    layer2_outputs(7076) <= not b or a;
    layer2_outputs(7077) <= a xor b;
    layer2_outputs(7078) <= a;
    layer2_outputs(7079) <= not a or b;
    layer2_outputs(7080) <= a and not b;
    layer2_outputs(7081) <= a or b;
    layer2_outputs(7082) <= b and not a;
    layer2_outputs(7083) <= not (a xor b);
    layer2_outputs(7084) <= not a;
    layer2_outputs(7085) <= not a or b;
    layer2_outputs(7086) <= a xor b;
    layer2_outputs(7087) <= b and not a;
    layer2_outputs(7088) <= a and not b;
    layer2_outputs(7089) <= not (a or b);
    layer2_outputs(7090) <= not b;
    layer2_outputs(7091) <= not (a xor b);
    layer2_outputs(7092) <= not (a or b);
    layer2_outputs(7093) <= not b;
    layer2_outputs(7094) <= not (a and b);
    layer2_outputs(7095) <= not (a and b);
    layer2_outputs(7096) <= not b;
    layer2_outputs(7097) <= not a;
    layer2_outputs(7098) <= not a or b;
    layer2_outputs(7099) <= a xor b;
    layer2_outputs(7100) <= a or b;
    layer2_outputs(7101) <= a and b;
    layer2_outputs(7102) <= not a;
    layer2_outputs(7103) <= not a or b;
    layer2_outputs(7104) <= not b;
    layer2_outputs(7105) <= a;
    layer2_outputs(7106) <= 1'b1;
    layer2_outputs(7107) <= a or b;
    layer2_outputs(7108) <= not (a and b);
    layer2_outputs(7109) <= b;
    layer2_outputs(7110) <= a;
    layer2_outputs(7111) <= not b;
    layer2_outputs(7112) <= a xor b;
    layer2_outputs(7113) <= not a or b;
    layer2_outputs(7114) <= b;
    layer2_outputs(7115) <= a and b;
    layer2_outputs(7116) <= a and b;
    layer2_outputs(7117) <= not (a and b);
    layer2_outputs(7118) <= not (a or b);
    layer2_outputs(7119) <= a or b;
    layer2_outputs(7120) <= a and b;
    layer2_outputs(7121) <= a or b;
    layer2_outputs(7122) <= not b;
    layer2_outputs(7123) <= a xor b;
    layer2_outputs(7124) <= not b;
    layer2_outputs(7125) <= b;
    layer2_outputs(7126) <= a;
    layer2_outputs(7127) <= not (a and b);
    layer2_outputs(7128) <= b and not a;
    layer2_outputs(7129) <= 1'b0;
    layer2_outputs(7130) <= 1'b0;
    layer2_outputs(7131) <= b;
    layer2_outputs(7132) <= a;
    layer2_outputs(7133) <= b;
    layer2_outputs(7134) <= not (a or b);
    layer2_outputs(7135) <= not a;
    layer2_outputs(7136) <= not (a and b);
    layer2_outputs(7137) <= b;
    layer2_outputs(7138) <= a;
    layer2_outputs(7139) <= not b or a;
    layer2_outputs(7140) <= a;
    layer2_outputs(7141) <= not a or b;
    layer2_outputs(7142) <= a;
    layer2_outputs(7143) <= not b;
    layer2_outputs(7144) <= a xor b;
    layer2_outputs(7145) <= a and not b;
    layer2_outputs(7146) <= not a;
    layer2_outputs(7147) <= a;
    layer2_outputs(7148) <= b;
    layer2_outputs(7149) <= 1'b1;
    layer2_outputs(7150) <= a and b;
    layer2_outputs(7151) <= b and not a;
    layer2_outputs(7152) <= a or b;
    layer2_outputs(7153) <= 1'b1;
    layer2_outputs(7154) <= a and b;
    layer2_outputs(7155) <= not (a and b);
    layer2_outputs(7156) <= not a;
    layer2_outputs(7157) <= a and b;
    layer2_outputs(7158) <= not a;
    layer2_outputs(7159) <= not a or b;
    layer2_outputs(7160) <= not b;
    layer2_outputs(7161) <= a;
    layer2_outputs(7162) <= not a;
    layer2_outputs(7163) <= not (a or b);
    layer2_outputs(7164) <= a;
    layer2_outputs(7165) <= b and not a;
    layer2_outputs(7166) <= a or b;
    layer2_outputs(7167) <= a or b;
    layer2_outputs(7168) <= a;
    layer2_outputs(7169) <= a;
    layer2_outputs(7170) <= not a;
    layer2_outputs(7171) <= not (a or b);
    layer2_outputs(7172) <= not b;
    layer2_outputs(7173) <= 1'b1;
    layer2_outputs(7174) <= a;
    layer2_outputs(7175) <= not a or b;
    layer2_outputs(7176) <= not (a or b);
    layer2_outputs(7177) <= a;
    layer2_outputs(7178) <= a;
    layer2_outputs(7179) <= 1'b0;
    layer2_outputs(7180) <= not b or a;
    layer2_outputs(7181) <= not (a and b);
    layer2_outputs(7182) <= a and not b;
    layer2_outputs(7183) <= 1'b0;
    layer2_outputs(7184) <= a;
    layer2_outputs(7185) <= not b;
    layer2_outputs(7186) <= not b or a;
    layer2_outputs(7187) <= a and not b;
    layer2_outputs(7188) <= b;
    layer2_outputs(7189) <= b;
    layer2_outputs(7190) <= 1'b1;
    layer2_outputs(7191) <= a;
    layer2_outputs(7192) <= a and not b;
    layer2_outputs(7193) <= a and not b;
    layer2_outputs(7194) <= a xor b;
    layer2_outputs(7195) <= not (a xor b);
    layer2_outputs(7196) <= a and not b;
    layer2_outputs(7197) <= not b;
    layer2_outputs(7198) <= not b;
    layer2_outputs(7199) <= 1'b1;
    layer2_outputs(7200) <= not (a or b);
    layer2_outputs(7201) <= b and not a;
    layer2_outputs(7202) <= 1'b0;
    layer2_outputs(7203) <= not b;
    layer2_outputs(7204) <= a;
    layer2_outputs(7205) <= not a;
    layer2_outputs(7206) <= not b;
    layer2_outputs(7207) <= not a or b;
    layer2_outputs(7208) <= a;
    layer2_outputs(7209) <= not a;
    layer2_outputs(7210) <= not (a xor b);
    layer2_outputs(7211) <= not (a and b);
    layer2_outputs(7212) <= not b;
    layer2_outputs(7213) <= a and b;
    layer2_outputs(7214) <= not a or b;
    layer2_outputs(7215) <= not b;
    layer2_outputs(7216) <= a;
    layer2_outputs(7217) <= a and not b;
    layer2_outputs(7218) <= 1'b0;
    layer2_outputs(7219) <= b;
    layer2_outputs(7220) <= not b;
    layer2_outputs(7221) <= not (a and b);
    layer2_outputs(7222) <= a and b;
    layer2_outputs(7223) <= b;
    layer2_outputs(7224) <= not a or b;
    layer2_outputs(7225) <= not (a and b);
    layer2_outputs(7226) <= a;
    layer2_outputs(7227) <= b;
    layer2_outputs(7228) <= not (a or b);
    layer2_outputs(7229) <= b and not a;
    layer2_outputs(7230) <= a xor b;
    layer2_outputs(7231) <= not a or b;
    layer2_outputs(7232) <= a xor b;
    layer2_outputs(7233) <= a xor b;
    layer2_outputs(7234) <= not b or a;
    layer2_outputs(7235) <= not b;
    layer2_outputs(7236) <= not b or a;
    layer2_outputs(7237) <= a xor b;
    layer2_outputs(7238) <= a xor b;
    layer2_outputs(7239) <= not a;
    layer2_outputs(7240) <= b and not a;
    layer2_outputs(7241) <= not (a or b);
    layer2_outputs(7242) <= not b;
    layer2_outputs(7243) <= a or b;
    layer2_outputs(7244) <= not b;
    layer2_outputs(7245) <= not (a xor b);
    layer2_outputs(7246) <= b;
    layer2_outputs(7247) <= a or b;
    layer2_outputs(7248) <= not (a or b);
    layer2_outputs(7249) <= a xor b;
    layer2_outputs(7250) <= not a;
    layer2_outputs(7251) <= not a;
    layer2_outputs(7252) <= b and not a;
    layer2_outputs(7253) <= not a or b;
    layer2_outputs(7254) <= not a or b;
    layer2_outputs(7255) <= a and not b;
    layer2_outputs(7256) <= not a;
    layer2_outputs(7257) <= a and not b;
    layer2_outputs(7258) <= not b or a;
    layer2_outputs(7259) <= a;
    layer2_outputs(7260) <= a or b;
    layer2_outputs(7261) <= b and not a;
    layer2_outputs(7262) <= b and not a;
    layer2_outputs(7263) <= b and not a;
    layer2_outputs(7264) <= not b or a;
    layer2_outputs(7265) <= not (a and b);
    layer2_outputs(7266) <= a and b;
    layer2_outputs(7267) <= a;
    layer2_outputs(7268) <= not b;
    layer2_outputs(7269) <= not b;
    layer2_outputs(7270) <= a or b;
    layer2_outputs(7271) <= a xor b;
    layer2_outputs(7272) <= not a or b;
    layer2_outputs(7273) <= not b;
    layer2_outputs(7274) <= a and b;
    layer2_outputs(7275) <= not a or b;
    layer2_outputs(7276) <= not (a and b);
    layer2_outputs(7277) <= a;
    layer2_outputs(7278) <= a and b;
    layer2_outputs(7279) <= a or b;
    layer2_outputs(7280) <= not a;
    layer2_outputs(7281) <= a xor b;
    layer2_outputs(7282) <= a or b;
    layer2_outputs(7283) <= not b or a;
    layer2_outputs(7284) <= a;
    layer2_outputs(7285) <= not b;
    layer2_outputs(7286) <= not a;
    layer2_outputs(7287) <= a and not b;
    layer2_outputs(7288) <= not b or a;
    layer2_outputs(7289) <= not b;
    layer2_outputs(7290) <= not a;
    layer2_outputs(7291) <= not (a xor b);
    layer2_outputs(7292) <= not (a and b);
    layer2_outputs(7293) <= not a or b;
    layer2_outputs(7294) <= b;
    layer2_outputs(7295) <= not b or a;
    layer2_outputs(7296) <= not a;
    layer2_outputs(7297) <= not a;
    layer2_outputs(7298) <= not (a or b);
    layer2_outputs(7299) <= a;
    layer2_outputs(7300) <= not (a and b);
    layer2_outputs(7301) <= b;
    layer2_outputs(7302) <= not b;
    layer2_outputs(7303) <= a xor b;
    layer2_outputs(7304) <= b and not a;
    layer2_outputs(7305) <= not a or b;
    layer2_outputs(7306) <= a and b;
    layer2_outputs(7307) <= b;
    layer2_outputs(7308) <= a and not b;
    layer2_outputs(7309) <= not (a and b);
    layer2_outputs(7310) <= not a;
    layer2_outputs(7311) <= b;
    layer2_outputs(7312) <= a and b;
    layer2_outputs(7313) <= not (a and b);
    layer2_outputs(7314) <= a;
    layer2_outputs(7315) <= not b or a;
    layer2_outputs(7316) <= a;
    layer2_outputs(7317) <= not (a or b);
    layer2_outputs(7318) <= not b;
    layer2_outputs(7319) <= 1'b1;
    layer2_outputs(7320) <= a and b;
    layer2_outputs(7321) <= not (a or b);
    layer2_outputs(7322) <= b;
    layer2_outputs(7323) <= a;
    layer2_outputs(7324) <= not a;
    layer2_outputs(7325) <= not b or a;
    layer2_outputs(7326) <= not a or b;
    layer2_outputs(7327) <= a xor b;
    layer2_outputs(7328) <= not b;
    layer2_outputs(7329) <= b and not a;
    layer2_outputs(7330) <= not a or b;
    layer2_outputs(7331) <= not b or a;
    layer2_outputs(7332) <= not (a and b);
    layer2_outputs(7333) <= not (a xor b);
    layer2_outputs(7334) <= a;
    layer2_outputs(7335) <= not b;
    layer2_outputs(7336) <= b;
    layer2_outputs(7337) <= not b;
    layer2_outputs(7338) <= not b or a;
    layer2_outputs(7339) <= not (a xor b);
    layer2_outputs(7340) <= b;
    layer2_outputs(7341) <= not b;
    layer2_outputs(7342) <= a or b;
    layer2_outputs(7343) <= a and not b;
    layer2_outputs(7344) <= 1'b1;
    layer2_outputs(7345) <= a or b;
    layer2_outputs(7346) <= not a or b;
    layer2_outputs(7347) <= not a;
    layer2_outputs(7348) <= a;
    layer2_outputs(7349) <= not b;
    layer2_outputs(7350) <= a xor b;
    layer2_outputs(7351) <= not b;
    layer2_outputs(7352) <= a and b;
    layer2_outputs(7353) <= a or b;
    layer2_outputs(7354) <= a or b;
    layer2_outputs(7355) <= not b;
    layer2_outputs(7356) <= not b;
    layer2_outputs(7357) <= not (a xor b);
    layer2_outputs(7358) <= not a;
    layer2_outputs(7359) <= not a;
    layer2_outputs(7360) <= a;
    layer2_outputs(7361) <= not b;
    layer2_outputs(7362) <= not b;
    layer2_outputs(7363) <= not a or b;
    layer2_outputs(7364) <= a;
    layer2_outputs(7365) <= a and b;
    layer2_outputs(7366) <= b;
    layer2_outputs(7367) <= b;
    layer2_outputs(7368) <= b;
    layer2_outputs(7369) <= a;
    layer2_outputs(7370) <= not (a and b);
    layer2_outputs(7371) <= a;
    layer2_outputs(7372) <= not b or a;
    layer2_outputs(7373) <= not a;
    layer2_outputs(7374) <= not a or b;
    layer2_outputs(7375) <= a and not b;
    layer2_outputs(7376) <= a;
    layer2_outputs(7377) <= not (a xor b);
    layer2_outputs(7378) <= not (a xor b);
    layer2_outputs(7379) <= a and not b;
    layer2_outputs(7380) <= b;
    layer2_outputs(7381) <= not (a or b);
    layer2_outputs(7382) <= not a;
    layer2_outputs(7383) <= a;
    layer2_outputs(7384) <= not b or a;
    layer2_outputs(7385) <= a and not b;
    layer2_outputs(7386) <= b;
    layer2_outputs(7387) <= not b or a;
    layer2_outputs(7388) <= not (a xor b);
    layer2_outputs(7389) <= a;
    layer2_outputs(7390) <= not (a or b);
    layer2_outputs(7391) <= not a;
    layer2_outputs(7392) <= a or b;
    layer2_outputs(7393) <= b;
    layer2_outputs(7394) <= a and b;
    layer2_outputs(7395) <= not a;
    layer2_outputs(7396) <= not (a or b);
    layer2_outputs(7397) <= a xor b;
    layer2_outputs(7398) <= b;
    layer2_outputs(7399) <= not a;
    layer2_outputs(7400) <= a;
    layer2_outputs(7401) <= not (a or b);
    layer2_outputs(7402) <= b;
    layer2_outputs(7403) <= a and not b;
    layer2_outputs(7404) <= not a;
    layer2_outputs(7405) <= a or b;
    layer2_outputs(7406) <= not b or a;
    layer2_outputs(7407) <= not (a or b);
    layer2_outputs(7408) <= b;
    layer2_outputs(7409) <= a and b;
    layer2_outputs(7410) <= not b or a;
    layer2_outputs(7411) <= a and b;
    layer2_outputs(7412) <= not (a and b);
    layer2_outputs(7413) <= b;
    layer2_outputs(7414) <= a and not b;
    layer2_outputs(7415) <= b;
    layer2_outputs(7416) <= b and not a;
    layer2_outputs(7417) <= a or b;
    layer2_outputs(7418) <= not b;
    layer2_outputs(7419) <= not a;
    layer2_outputs(7420) <= not b;
    layer2_outputs(7421) <= a and not b;
    layer2_outputs(7422) <= a xor b;
    layer2_outputs(7423) <= not b or a;
    layer2_outputs(7424) <= a or b;
    layer2_outputs(7425) <= not a;
    layer2_outputs(7426) <= not b;
    layer2_outputs(7427) <= a and b;
    layer2_outputs(7428) <= not (a and b);
    layer2_outputs(7429) <= 1'b1;
    layer2_outputs(7430) <= a and not b;
    layer2_outputs(7431) <= not a or b;
    layer2_outputs(7432) <= a and not b;
    layer2_outputs(7433) <= not a or b;
    layer2_outputs(7434) <= a;
    layer2_outputs(7435) <= not (a or b);
    layer2_outputs(7436) <= not a or b;
    layer2_outputs(7437) <= not b or a;
    layer2_outputs(7438) <= not b or a;
    layer2_outputs(7439) <= not a or b;
    layer2_outputs(7440) <= b and not a;
    layer2_outputs(7441) <= a or b;
    layer2_outputs(7442) <= not (a and b);
    layer2_outputs(7443) <= not b;
    layer2_outputs(7444) <= 1'b0;
    layer2_outputs(7445) <= not (a xor b);
    layer2_outputs(7446) <= not (a or b);
    layer2_outputs(7447) <= a and b;
    layer2_outputs(7448) <= a or b;
    layer2_outputs(7449) <= a;
    layer2_outputs(7450) <= not a;
    layer2_outputs(7451) <= a and b;
    layer2_outputs(7452) <= not b;
    layer2_outputs(7453) <= not b;
    layer2_outputs(7454) <= not a;
    layer2_outputs(7455) <= not b or a;
    layer2_outputs(7456) <= a and b;
    layer2_outputs(7457) <= not (a and b);
    layer2_outputs(7458) <= not (a or b);
    layer2_outputs(7459) <= a and not b;
    layer2_outputs(7460) <= a xor b;
    layer2_outputs(7461) <= not b;
    layer2_outputs(7462) <= not a or b;
    layer2_outputs(7463) <= not a or b;
    layer2_outputs(7464) <= not (a or b);
    layer2_outputs(7465) <= b;
    layer2_outputs(7466) <= not (a and b);
    layer2_outputs(7467) <= not a;
    layer2_outputs(7468) <= not (a and b);
    layer2_outputs(7469) <= a or b;
    layer2_outputs(7470) <= a or b;
    layer2_outputs(7471) <= not b;
    layer2_outputs(7472) <= not b;
    layer2_outputs(7473) <= not (a xor b);
    layer2_outputs(7474) <= not a;
    layer2_outputs(7475) <= not a or b;
    layer2_outputs(7476) <= b;
    layer2_outputs(7477) <= a or b;
    layer2_outputs(7478) <= b;
    layer2_outputs(7479) <= not b or a;
    layer2_outputs(7480) <= not (a xor b);
    layer2_outputs(7481) <= not (a xor b);
    layer2_outputs(7482) <= b;
    layer2_outputs(7483) <= b;
    layer2_outputs(7484) <= a;
    layer2_outputs(7485) <= a and b;
    layer2_outputs(7486) <= not a or b;
    layer2_outputs(7487) <= b;
    layer2_outputs(7488) <= a;
    layer2_outputs(7489) <= a;
    layer2_outputs(7490) <= a and b;
    layer2_outputs(7491) <= not b;
    layer2_outputs(7492) <= a xor b;
    layer2_outputs(7493) <= not a;
    layer2_outputs(7494) <= 1'b0;
    layer2_outputs(7495) <= a and b;
    layer2_outputs(7496) <= not (a and b);
    layer2_outputs(7497) <= not (a and b);
    layer2_outputs(7498) <= not (a or b);
    layer2_outputs(7499) <= not (a and b);
    layer2_outputs(7500) <= not a;
    layer2_outputs(7501) <= not a;
    layer2_outputs(7502) <= not b;
    layer2_outputs(7503) <= b;
    layer2_outputs(7504) <= not b;
    layer2_outputs(7505) <= not b or a;
    layer2_outputs(7506) <= not b or a;
    layer2_outputs(7507) <= a and not b;
    layer2_outputs(7508) <= not a;
    layer2_outputs(7509) <= a;
    layer2_outputs(7510) <= not (a and b);
    layer2_outputs(7511) <= not a;
    layer2_outputs(7512) <= a or b;
    layer2_outputs(7513) <= a or b;
    layer2_outputs(7514) <= not a;
    layer2_outputs(7515) <= a and b;
    layer2_outputs(7516) <= a or b;
    layer2_outputs(7517) <= not b or a;
    layer2_outputs(7518) <= a;
    layer2_outputs(7519) <= not b or a;
    layer2_outputs(7520) <= not a;
    layer2_outputs(7521) <= b;
    layer2_outputs(7522) <= a or b;
    layer2_outputs(7523) <= a;
    layer2_outputs(7524) <= a;
    layer2_outputs(7525) <= b;
    layer2_outputs(7526) <= 1'b1;
    layer2_outputs(7527) <= not a;
    layer2_outputs(7528) <= b and not a;
    layer2_outputs(7529) <= b;
    layer2_outputs(7530) <= b and not a;
    layer2_outputs(7531) <= a;
    layer2_outputs(7532) <= b and not a;
    layer2_outputs(7533) <= a or b;
    layer2_outputs(7534) <= a or b;
    layer2_outputs(7535) <= not a;
    layer2_outputs(7536) <= a;
    layer2_outputs(7537) <= not a;
    layer2_outputs(7538) <= not a;
    layer2_outputs(7539) <= not b or a;
    layer2_outputs(7540) <= a xor b;
    layer2_outputs(7541) <= not a or b;
    layer2_outputs(7542) <= a or b;
    layer2_outputs(7543) <= not a;
    layer2_outputs(7544) <= not (a or b);
    layer2_outputs(7545) <= not (a or b);
    layer2_outputs(7546) <= b;
    layer2_outputs(7547) <= a or b;
    layer2_outputs(7548) <= not (a xor b);
    layer2_outputs(7549) <= 1'b0;
    layer2_outputs(7550) <= a;
    layer2_outputs(7551) <= b and not a;
    layer2_outputs(7552) <= a and not b;
    layer2_outputs(7553) <= 1'b1;
    layer2_outputs(7554) <= a;
    layer2_outputs(7555) <= a or b;
    layer2_outputs(7556) <= b;
    layer2_outputs(7557) <= a and not b;
    layer2_outputs(7558) <= a xor b;
    layer2_outputs(7559) <= not (a xor b);
    layer2_outputs(7560) <= not a;
    layer2_outputs(7561) <= b;
    layer2_outputs(7562) <= not a;
    layer2_outputs(7563) <= not b;
    layer2_outputs(7564) <= a xor b;
    layer2_outputs(7565) <= not b or a;
    layer2_outputs(7566) <= a;
    layer2_outputs(7567) <= a or b;
    layer2_outputs(7568) <= a xor b;
    layer2_outputs(7569) <= not (a or b);
    layer2_outputs(7570) <= not (a xor b);
    layer2_outputs(7571) <= not (a or b);
    layer2_outputs(7572) <= a;
    layer2_outputs(7573) <= b and not a;
    layer2_outputs(7574) <= a and not b;
    layer2_outputs(7575) <= a and b;
    layer2_outputs(7576) <= b;
    layer2_outputs(7577) <= b;
    layer2_outputs(7578) <= b;
    layer2_outputs(7579) <= a and not b;
    layer2_outputs(7580) <= not (a and b);
    layer2_outputs(7581) <= not b or a;
    layer2_outputs(7582) <= a and b;
    layer2_outputs(7583) <= b;
    layer2_outputs(7584) <= not a or b;
    layer2_outputs(7585) <= not b or a;
    layer2_outputs(7586) <= a xor b;
    layer2_outputs(7587) <= a or b;
    layer2_outputs(7588) <= b;
    layer2_outputs(7589) <= not b;
    layer2_outputs(7590) <= not b;
    layer2_outputs(7591) <= a and not b;
    layer2_outputs(7592) <= not a;
    layer2_outputs(7593) <= b and not a;
    layer2_outputs(7594) <= not a;
    layer2_outputs(7595) <= b and not a;
    layer2_outputs(7596) <= b;
    layer2_outputs(7597) <= b;
    layer2_outputs(7598) <= b;
    layer2_outputs(7599) <= a;
    layer2_outputs(7600) <= b and not a;
    layer2_outputs(7601) <= not (a and b);
    layer2_outputs(7602) <= a and not b;
    layer2_outputs(7603) <= a and b;
    layer2_outputs(7604) <= b;
    layer2_outputs(7605) <= not a;
    layer2_outputs(7606) <= not a or b;
    layer2_outputs(7607) <= a;
    layer2_outputs(7608) <= b;
    layer2_outputs(7609) <= a;
    layer2_outputs(7610) <= a xor b;
    layer2_outputs(7611) <= a;
    layer2_outputs(7612) <= not (a or b);
    layer2_outputs(7613) <= not (a or b);
    layer2_outputs(7614) <= b;
    layer2_outputs(7615) <= 1'b0;
    layer2_outputs(7616) <= not (a and b);
    layer2_outputs(7617) <= not b;
    layer2_outputs(7618) <= a xor b;
    layer2_outputs(7619) <= not a;
    layer2_outputs(7620) <= a xor b;
    layer2_outputs(7621) <= b;
    layer2_outputs(7622) <= a xor b;
    layer2_outputs(7623) <= not (a xor b);
    layer2_outputs(7624) <= a and b;
    layer2_outputs(7625) <= not a;
    layer2_outputs(7626) <= a;
    layer2_outputs(7627) <= not (a and b);
    layer2_outputs(7628) <= not b or a;
    layer2_outputs(7629) <= not a;
    layer2_outputs(7630) <= not b;
    layer2_outputs(7631) <= a or b;
    layer2_outputs(7632) <= 1'b0;
    layer2_outputs(7633) <= b;
    layer2_outputs(7634) <= a and not b;
    layer2_outputs(7635) <= a;
    layer2_outputs(7636) <= not (a and b);
    layer2_outputs(7637) <= not b or a;
    layer2_outputs(7638) <= a;
    layer2_outputs(7639) <= not a;
    layer2_outputs(7640) <= a and not b;
    layer2_outputs(7641) <= not a;
    layer2_outputs(7642) <= a or b;
    layer2_outputs(7643) <= a and not b;
    layer2_outputs(7644) <= a xor b;
    layer2_outputs(7645) <= a or b;
    layer2_outputs(7646) <= a or b;
    layer2_outputs(7647) <= not b;
    layer2_outputs(7648) <= a or b;
    layer2_outputs(7649) <= not (a and b);
    layer2_outputs(7650) <= a or b;
    layer2_outputs(7651) <= b;
    layer2_outputs(7652) <= b and not a;
    layer2_outputs(7653) <= a or b;
    layer2_outputs(7654) <= a and not b;
    layer2_outputs(7655) <= not (a and b);
    layer2_outputs(7656) <= a and b;
    layer2_outputs(7657) <= a and not b;
    layer2_outputs(7658) <= a and not b;
    layer2_outputs(7659) <= 1'b0;
    layer2_outputs(7660) <= not a or b;
    layer2_outputs(7661) <= not a;
    layer2_outputs(7662) <= a;
    layer2_outputs(7663) <= not a;
    layer2_outputs(7664) <= a or b;
    layer2_outputs(7665) <= a and not b;
    layer2_outputs(7666) <= not b;
    layer2_outputs(7667) <= b;
    layer2_outputs(7668) <= not a or b;
    layer2_outputs(7669) <= not a;
    layer2_outputs(7670) <= b and not a;
    layer2_outputs(7671) <= not (a or b);
    layer2_outputs(7672) <= not (a xor b);
    layer2_outputs(7673) <= a xor b;
    layer2_outputs(7674) <= a or b;
    layer2_outputs(7675) <= not b or a;
    layer2_outputs(7676) <= not (a and b);
    layer2_outputs(7677) <= not a or b;
    layer2_outputs(7678) <= a and not b;
    layer2_outputs(7679) <= not (a and b);
    layer2_outputs(7680) <= b and not a;
    layer2_outputs(7681) <= not b;
    layer2_outputs(7682) <= not b or a;
    layer2_outputs(7683) <= not b or a;
    layer2_outputs(7684) <= not b;
    layer2_outputs(7685) <= b;
    layer2_outputs(7686) <= b;
    layer2_outputs(7687) <= b;
    layer2_outputs(7688) <= not b;
    layer2_outputs(7689) <= not a or b;
    layer2_outputs(7690) <= not b;
    layer2_outputs(7691) <= a;
    layer2_outputs(7692) <= not a;
    layer2_outputs(7693) <= a and not b;
    layer2_outputs(7694) <= not b;
    layer2_outputs(7695) <= not (a and b);
    layer2_outputs(7696) <= not b or a;
    layer2_outputs(7697) <= b;
    layer2_outputs(7698) <= not b or a;
    layer2_outputs(7699) <= not b;
    layer2_outputs(7700) <= not b or a;
    layer2_outputs(7701) <= not (a and b);
    layer2_outputs(7702) <= a;
    layer2_outputs(7703) <= not b;
    layer2_outputs(7704) <= not a or b;
    layer2_outputs(7705) <= a xor b;
    layer2_outputs(7706) <= not (a and b);
    layer2_outputs(7707) <= not a or b;
    layer2_outputs(7708) <= a or b;
    layer2_outputs(7709) <= b;
    layer2_outputs(7710) <= not (a or b);
    layer2_outputs(7711) <= not b or a;
    layer2_outputs(7712) <= a or b;
    layer2_outputs(7713) <= not (a or b);
    layer2_outputs(7714) <= 1'b0;
    layer2_outputs(7715) <= a;
    layer2_outputs(7716) <= not a or b;
    layer2_outputs(7717) <= a or b;
    layer2_outputs(7718) <= a;
    layer2_outputs(7719) <= 1'b1;
    layer2_outputs(7720) <= b;
    layer2_outputs(7721) <= not b;
    layer2_outputs(7722) <= a;
    layer2_outputs(7723) <= b and not a;
    layer2_outputs(7724) <= a;
    layer2_outputs(7725) <= a;
    layer2_outputs(7726) <= not b or a;
    layer2_outputs(7727) <= a;
    layer2_outputs(7728) <= not (a and b);
    layer2_outputs(7729) <= not (a or b);
    layer2_outputs(7730) <= not (a xor b);
    layer2_outputs(7731) <= not a or b;
    layer2_outputs(7732) <= b;
    layer2_outputs(7733) <= a xor b;
    layer2_outputs(7734) <= a;
    layer2_outputs(7735) <= not a;
    layer2_outputs(7736) <= not b or a;
    layer2_outputs(7737) <= b;
    layer2_outputs(7738) <= not a or b;
    layer2_outputs(7739) <= not a or b;
    layer2_outputs(7740) <= not a;
    layer2_outputs(7741) <= b;
    layer2_outputs(7742) <= a and b;
    layer2_outputs(7743) <= a and not b;
    layer2_outputs(7744) <= not (a or b);
    layer2_outputs(7745) <= a;
    layer2_outputs(7746) <= b and not a;
    layer2_outputs(7747) <= b;
    layer2_outputs(7748) <= 1'b0;
    layer2_outputs(7749) <= not a;
    layer2_outputs(7750) <= not (a or b);
    layer2_outputs(7751) <= a and b;
    layer2_outputs(7752) <= a;
    layer2_outputs(7753) <= a and b;
    layer2_outputs(7754) <= a and not b;
    layer2_outputs(7755) <= a or b;
    layer2_outputs(7756) <= not a;
    layer2_outputs(7757) <= a;
    layer2_outputs(7758) <= a and b;
    layer2_outputs(7759) <= not (a and b);
    layer2_outputs(7760) <= not b;
    layer2_outputs(7761) <= b and not a;
    layer2_outputs(7762) <= not b;
    layer2_outputs(7763) <= a;
    layer2_outputs(7764) <= not (a xor b);
    layer2_outputs(7765) <= not b or a;
    layer2_outputs(7766) <= not a;
    layer2_outputs(7767) <= not (a xor b);
    layer2_outputs(7768) <= a and b;
    layer2_outputs(7769) <= a or b;
    layer2_outputs(7770) <= 1'b0;
    layer2_outputs(7771) <= not a;
    layer2_outputs(7772) <= not b or a;
    layer2_outputs(7773) <= not b or a;
    layer2_outputs(7774) <= not b or a;
    layer2_outputs(7775) <= a or b;
    layer2_outputs(7776) <= not b;
    layer2_outputs(7777) <= b and not a;
    layer2_outputs(7778) <= not (a xor b);
    layer2_outputs(7779) <= not (a or b);
    layer2_outputs(7780) <= not b or a;
    layer2_outputs(7781) <= b and not a;
    layer2_outputs(7782) <= not a or b;
    layer2_outputs(7783) <= not b;
    layer2_outputs(7784) <= a;
    layer2_outputs(7785) <= not a or b;
    layer2_outputs(7786) <= not (a or b);
    layer2_outputs(7787) <= not a;
    layer2_outputs(7788) <= a;
    layer2_outputs(7789) <= b;
    layer2_outputs(7790) <= b and not a;
    layer2_outputs(7791) <= a xor b;
    layer2_outputs(7792) <= not a;
    layer2_outputs(7793) <= not (a xor b);
    layer2_outputs(7794) <= a and not b;
    layer2_outputs(7795) <= a;
    layer2_outputs(7796) <= b;
    layer2_outputs(7797) <= not (a or b);
    layer2_outputs(7798) <= b and not a;
    layer2_outputs(7799) <= a xor b;
    layer2_outputs(7800) <= not a or b;
    layer2_outputs(7801) <= b;
    layer2_outputs(7802) <= not a or b;
    layer2_outputs(7803) <= a or b;
    layer2_outputs(7804) <= b;
    layer2_outputs(7805) <= not b or a;
    layer2_outputs(7806) <= 1'b1;
    layer2_outputs(7807) <= b and not a;
    layer2_outputs(7808) <= a and b;
    layer2_outputs(7809) <= a or b;
    layer2_outputs(7810) <= a or b;
    layer2_outputs(7811) <= a and not b;
    layer2_outputs(7812) <= 1'b1;
    layer2_outputs(7813) <= a xor b;
    layer2_outputs(7814) <= not (a or b);
    layer2_outputs(7815) <= a and b;
    layer2_outputs(7816) <= a and not b;
    layer2_outputs(7817) <= not a or b;
    layer2_outputs(7818) <= b and not a;
    layer2_outputs(7819) <= not a;
    layer2_outputs(7820) <= b and not a;
    layer2_outputs(7821) <= not a;
    layer2_outputs(7822) <= b;
    layer2_outputs(7823) <= a and b;
    layer2_outputs(7824) <= not a or b;
    layer2_outputs(7825) <= 1'b0;
    layer2_outputs(7826) <= a;
    layer2_outputs(7827) <= not a;
    layer2_outputs(7828) <= not a or b;
    layer2_outputs(7829) <= 1'b1;
    layer2_outputs(7830) <= 1'b0;
    layer2_outputs(7831) <= a xor b;
    layer2_outputs(7832) <= not (a xor b);
    layer2_outputs(7833) <= not b or a;
    layer2_outputs(7834) <= a and b;
    layer2_outputs(7835) <= not a;
    layer2_outputs(7836) <= a xor b;
    layer2_outputs(7837) <= a and b;
    layer2_outputs(7838) <= b;
    layer2_outputs(7839) <= b;
    layer2_outputs(7840) <= b;
    layer2_outputs(7841) <= not a;
    layer2_outputs(7842) <= not b or a;
    layer2_outputs(7843) <= a and b;
    layer2_outputs(7844) <= not b or a;
    layer2_outputs(7845) <= b;
    layer2_outputs(7846) <= a;
    layer2_outputs(7847) <= not b;
    layer2_outputs(7848) <= not (a or b);
    layer2_outputs(7849) <= not b;
    layer2_outputs(7850) <= not (a or b);
    layer2_outputs(7851) <= b and not a;
    layer2_outputs(7852) <= not b;
    layer2_outputs(7853) <= 1'b0;
    layer2_outputs(7854) <= not a;
    layer2_outputs(7855) <= not b;
    layer2_outputs(7856) <= b;
    layer2_outputs(7857) <= a and not b;
    layer2_outputs(7858) <= not (a or b);
    layer2_outputs(7859) <= not a or b;
    layer2_outputs(7860) <= not b;
    layer2_outputs(7861) <= not b or a;
    layer2_outputs(7862) <= not a;
    layer2_outputs(7863) <= a xor b;
    layer2_outputs(7864) <= not b or a;
    layer2_outputs(7865) <= a;
    layer2_outputs(7866) <= a or b;
    layer2_outputs(7867) <= b and not a;
    layer2_outputs(7868) <= not (a and b);
    layer2_outputs(7869) <= not (a xor b);
    layer2_outputs(7870) <= 1'b0;
    layer2_outputs(7871) <= 1'b1;
    layer2_outputs(7872) <= not b or a;
    layer2_outputs(7873) <= b and not a;
    layer2_outputs(7874) <= not b;
    layer2_outputs(7875) <= b and not a;
    layer2_outputs(7876) <= not b;
    layer2_outputs(7877) <= a;
    layer2_outputs(7878) <= not (a or b);
    layer2_outputs(7879) <= a xor b;
    layer2_outputs(7880) <= b;
    layer2_outputs(7881) <= not a or b;
    layer2_outputs(7882) <= a or b;
    layer2_outputs(7883) <= not b;
    layer2_outputs(7884) <= a xor b;
    layer2_outputs(7885) <= b and not a;
    layer2_outputs(7886) <= not b or a;
    layer2_outputs(7887) <= not b or a;
    layer2_outputs(7888) <= a and b;
    layer2_outputs(7889) <= a xor b;
    layer2_outputs(7890) <= a;
    layer2_outputs(7891) <= not (a and b);
    layer2_outputs(7892) <= not b;
    layer2_outputs(7893) <= not b or a;
    layer2_outputs(7894) <= a and b;
    layer2_outputs(7895) <= not (a and b);
    layer2_outputs(7896) <= a;
    layer2_outputs(7897) <= not a or b;
    layer2_outputs(7898) <= a;
    layer2_outputs(7899) <= b;
    layer2_outputs(7900) <= a or b;
    layer2_outputs(7901) <= a;
    layer2_outputs(7902) <= not a or b;
    layer2_outputs(7903) <= not a or b;
    layer2_outputs(7904) <= not b;
    layer2_outputs(7905) <= not (a xor b);
    layer2_outputs(7906) <= a or b;
    layer2_outputs(7907) <= b and not a;
    layer2_outputs(7908) <= b;
    layer2_outputs(7909) <= not a or b;
    layer2_outputs(7910) <= a;
    layer2_outputs(7911) <= not (a or b);
    layer2_outputs(7912) <= a and not b;
    layer2_outputs(7913) <= b;
    layer2_outputs(7914) <= not (a and b);
    layer2_outputs(7915) <= a and not b;
    layer2_outputs(7916) <= a and b;
    layer2_outputs(7917) <= not b or a;
    layer2_outputs(7918) <= not a;
    layer2_outputs(7919) <= b;
    layer2_outputs(7920) <= not (a and b);
    layer2_outputs(7921) <= not (a or b);
    layer2_outputs(7922) <= a or b;
    layer2_outputs(7923) <= a;
    layer2_outputs(7924) <= a;
    layer2_outputs(7925) <= a and b;
    layer2_outputs(7926) <= b and not a;
    layer2_outputs(7927) <= a and b;
    layer2_outputs(7928) <= not b;
    layer2_outputs(7929) <= a or b;
    layer2_outputs(7930) <= not b;
    layer2_outputs(7931) <= a or b;
    layer2_outputs(7932) <= b;
    layer2_outputs(7933) <= b;
    layer2_outputs(7934) <= not a;
    layer2_outputs(7935) <= a or b;
    layer2_outputs(7936) <= a or b;
    layer2_outputs(7937) <= not a;
    layer2_outputs(7938) <= a and not b;
    layer2_outputs(7939) <= 1'b0;
    layer2_outputs(7940) <= not (a and b);
    layer2_outputs(7941) <= not a or b;
    layer2_outputs(7942) <= a xor b;
    layer2_outputs(7943) <= not (a or b);
    layer2_outputs(7944) <= not (a and b);
    layer2_outputs(7945) <= not (a xor b);
    layer2_outputs(7946) <= a and b;
    layer2_outputs(7947) <= not (a xor b);
    layer2_outputs(7948) <= b;
    layer2_outputs(7949) <= 1'b0;
    layer2_outputs(7950) <= not (a and b);
    layer2_outputs(7951) <= a or b;
    layer2_outputs(7952) <= a and not b;
    layer2_outputs(7953) <= a;
    layer2_outputs(7954) <= b;
    layer2_outputs(7955) <= not a;
    layer2_outputs(7956) <= not (a and b);
    layer2_outputs(7957) <= not b;
    layer2_outputs(7958) <= not a;
    layer2_outputs(7959) <= not b;
    layer2_outputs(7960) <= b and not a;
    layer2_outputs(7961) <= a and b;
    layer2_outputs(7962) <= not b or a;
    layer2_outputs(7963) <= a;
    layer2_outputs(7964) <= not (a or b);
    layer2_outputs(7965) <= not (a xor b);
    layer2_outputs(7966) <= a;
    layer2_outputs(7967) <= not b;
    layer2_outputs(7968) <= a and b;
    layer2_outputs(7969) <= a;
    layer2_outputs(7970) <= a xor b;
    layer2_outputs(7971) <= a and b;
    layer2_outputs(7972) <= not a;
    layer2_outputs(7973) <= a;
    layer2_outputs(7974) <= not (a xor b);
    layer2_outputs(7975) <= b;
    layer2_outputs(7976) <= not b or a;
    layer2_outputs(7977) <= 1'b0;
    layer2_outputs(7978) <= a and not b;
    layer2_outputs(7979) <= 1'b0;
    layer2_outputs(7980) <= not b or a;
    layer2_outputs(7981) <= not (a and b);
    layer2_outputs(7982) <= not a;
    layer2_outputs(7983) <= not a;
    layer2_outputs(7984) <= not b;
    layer2_outputs(7985) <= not (a and b);
    layer2_outputs(7986) <= not (a and b);
    layer2_outputs(7987) <= 1'b0;
    layer2_outputs(7988) <= not (a and b);
    layer2_outputs(7989) <= b and not a;
    layer2_outputs(7990) <= not (a or b);
    layer2_outputs(7991) <= not (a or b);
    layer2_outputs(7992) <= not (a xor b);
    layer2_outputs(7993) <= not (a or b);
    layer2_outputs(7994) <= b;
    layer2_outputs(7995) <= a and not b;
    layer2_outputs(7996) <= a and not b;
    layer2_outputs(7997) <= a;
    layer2_outputs(7998) <= a and not b;
    layer2_outputs(7999) <= not (a or b);
    layer2_outputs(8000) <= not a or b;
    layer2_outputs(8001) <= a or b;
    layer2_outputs(8002) <= b and not a;
    layer2_outputs(8003) <= a and not b;
    layer2_outputs(8004) <= not b or a;
    layer2_outputs(8005) <= not (a xor b);
    layer2_outputs(8006) <= not a or b;
    layer2_outputs(8007) <= not b or a;
    layer2_outputs(8008) <= not a;
    layer2_outputs(8009) <= b;
    layer2_outputs(8010) <= 1'b1;
    layer2_outputs(8011) <= a;
    layer2_outputs(8012) <= not (a and b);
    layer2_outputs(8013) <= a and not b;
    layer2_outputs(8014) <= not (a or b);
    layer2_outputs(8015) <= a;
    layer2_outputs(8016) <= not a;
    layer2_outputs(8017) <= not a;
    layer2_outputs(8018) <= a xor b;
    layer2_outputs(8019) <= not a;
    layer2_outputs(8020) <= not b;
    layer2_outputs(8021) <= a;
    layer2_outputs(8022) <= not b;
    layer2_outputs(8023) <= a xor b;
    layer2_outputs(8024) <= b and not a;
    layer2_outputs(8025) <= b;
    layer2_outputs(8026) <= a;
    layer2_outputs(8027) <= a and b;
    layer2_outputs(8028) <= a and not b;
    layer2_outputs(8029) <= not (a or b);
    layer2_outputs(8030) <= not (a and b);
    layer2_outputs(8031) <= not a or b;
    layer2_outputs(8032) <= a or b;
    layer2_outputs(8033) <= not b or a;
    layer2_outputs(8034) <= not (a xor b);
    layer2_outputs(8035) <= not b or a;
    layer2_outputs(8036) <= a or b;
    layer2_outputs(8037) <= a;
    layer2_outputs(8038) <= b;
    layer2_outputs(8039) <= a and b;
    layer2_outputs(8040) <= a and not b;
    layer2_outputs(8041) <= not b;
    layer2_outputs(8042) <= a xor b;
    layer2_outputs(8043) <= not a;
    layer2_outputs(8044) <= not (a and b);
    layer2_outputs(8045) <= a and not b;
    layer2_outputs(8046) <= not b or a;
    layer2_outputs(8047) <= not a;
    layer2_outputs(8048) <= not b;
    layer2_outputs(8049) <= a and not b;
    layer2_outputs(8050) <= a or b;
    layer2_outputs(8051) <= a and not b;
    layer2_outputs(8052) <= not (a or b);
    layer2_outputs(8053) <= b;
    layer2_outputs(8054) <= b;
    layer2_outputs(8055) <= not b;
    layer2_outputs(8056) <= a;
    layer2_outputs(8057) <= a and not b;
    layer2_outputs(8058) <= a;
    layer2_outputs(8059) <= not a or b;
    layer2_outputs(8060) <= not b;
    layer2_outputs(8061) <= not b;
    layer2_outputs(8062) <= 1'b1;
    layer2_outputs(8063) <= 1'b0;
    layer2_outputs(8064) <= 1'b0;
    layer2_outputs(8065) <= a;
    layer2_outputs(8066) <= not b or a;
    layer2_outputs(8067) <= a;
    layer2_outputs(8068) <= 1'b1;
    layer2_outputs(8069) <= b and not a;
    layer2_outputs(8070) <= not b;
    layer2_outputs(8071) <= not b;
    layer2_outputs(8072) <= not (a xor b);
    layer2_outputs(8073) <= a and not b;
    layer2_outputs(8074) <= not b or a;
    layer2_outputs(8075) <= not a;
    layer2_outputs(8076) <= a;
    layer2_outputs(8077) <= a and not b;
    layer2_outputs(8078) <= not b or a;
    layer2_outputs(8079) <= not a;
    layer2_outputs(8080) <= b;
    layer2_outputs(8081) <= a;
    layer2_outputs(8082) <= not a;
    layer2_outputs(8083) <= a and b;
    layer2_outputs(8084) <= not b;
    layer2_outputs(8085) <= not b;
    layer2_outputs(8086) <= not b;
    layer2_outputs(8087) <= not a;
    layer2_outputs(8088) <= a and b;
    layer2_outputs(8089) <= not (a and b);
    layer2_outputs(8090) <= b and not a;
    layer2_outputs(8091) <= not a;
    layer2_outputs(8092) <= b;
    layer2_outputs(8093) <= b;
    layer2_outputs(8094) <= b;
    layer2_outputs(8095) <= not (a xor b);
    layer2_outputs(8096) <= a and b;
    layer2_outputs(8097) <= a and not b;
    layer2_outputs(8098) <= a and not b;
    layer2_outputs(8099) <= not b;
    layer2_outputs(8100) <= not a;
    layer2_outputs(8101) <= a;
    layer2_outputs(8102) <= not a;
    layer2_outputs(8103) <= not b;
    layer2_outputs(8104) <= 1'b1;
    layer2_outputs(8105) <= b;
    layer2_outputs(8106) <= b;
    layer2_outputs(8107) <= not a;
    layer2_outputs(8108) <= not a;
    layer2_outputs(8109) <= b and not a;
    layer2_outputs(8110) <= a and b;
    layer2_outputs(8111) <= not (a xor b);
    layer2_outputs(8112) <= not (a or b);
    layer2_outputs(8113) <= a and b;
    layer2_outputs(8114) <= not a;
    layer2_outputs(8115) <= not (a or b);
    layer2_outputs(8116) <= not b or a;
    layer2_outputs(8117) <= not b;
    layer2_outputs(8118) <= not b;
    layer2_outputs(8119) <= not (a and b);
    layer2_outputs(8120) <= not (a xor b);
    layer2_outputs(8121) <= not b or a;
    layer2_outputs(8122) <= a or b;
    layer2_outputs(8123) <= a or b;
    layer2_outputs(8124) <= a or b;
    layer2_outputs(8125) <= a and b;
    layer2_outputs(8126) <= not b;
    layer2_outputs(8127) <= a xor b;
    layer2_outputs(8128) <= b;
    layer2_outputs(8129) <= not a;
    layer2_outputs(8130) <= not a or b;
    layer2_outputs(8131) <= a;
    layer2_outputs(8132) <= b and not a;
    layer2_outputs(8133) <= not b or a;
    layer2_outputs(8134) <= a;
    layer2_outputs(8135) <= a;
    layer2_outputs(8136) <= not a;
    layer2_outputs(8137) <= not (a or b);
    layer2_outputs(8138) <= b;
    layer2_outputs(8139) <= b and not a;
    layer2_outputs(8140) <= b;
    layer2_outputs(8141) <= not b;
    layer2_outputs(8142) <= not b or a;
    layer2_outputs(8143) <= b;
    layer2_outputs(8144) <= not a or b;
    layer2_outputs(8145) <= a;
    layer2_outputs(8146) <= not b or a;
    layer2_outputs(8147) <= not a or b;
    layer2_outputs(8148) <= not a;
    layer2_outputs(8149) <= not (a or b);
    layer2_outputs(8150) <= not a;
    layer2_outputs(8151) <= a and not b;
    layer2_outputs(8152) <= b;
    layer2_outputs(8153) <= not (a and b);
    layer2_outputs(8154) <= b and not a;
    layer2_outputs(8155) <= a or b;
    layer2_outputs(8156) <= a xor b;
    layer2_outputs(8157) <= not a;
    layer2_outputs(8158) <= a and b;
    layer2_outputs(8159) <= not (a and b);
    layer2_outputs(8160) <= not b or a;
    layer2_outputs(8161) <= a xor b;
    layer2_outputs(8162) <= not b or a;
    layer2_outputs(8163) <= b;
    layer2_outputs(8164) <= 1'b0;
    layer2_outputs(8165) <= not a;
    layer2_outputs(8166) <= a or b;
    layer2_outputs(8167) <= a or b;
    layer2_outputs(8168) <= not b;
    layer2_outputs(8169) <= not (a xor b);
    layer2_outputs(8170) <= b and not a;
    layer2_outputs(8171) <= not (a and b);
    layer2_outputs(8172) <= not a;
    layer2_outputs(8173) <= 1'b0;
    layer2_outputs(8174) <= not (a xor b);
    layer2_outputs(8175) <= a and b;
    layer2_outputs(8176) <= not b or a;
    layer2_outputs(8177) <= not a;
    layer2_outputs(8178) <= a and b;
    layer2_outputs(8179) <= not b;
    layer2_outputs(8180) <= a;
    layer2_outputs(8181) <= a xor b;
    layer2_outputs(8182) <= a;
    layer2_outputs(8183) <= a and b;
    layer2_outputs(8184) <= not b;
    layer2_outputs(8185) <= not (a xor b);
    layer2_outputs(8186) <= not a;
    layer2_outputs(8187) <= b;
    layer2_outputs(8188) <= not (a and b);
    layer2_outputs(8189) <= not a;
    layer2_outputs(8190) <= a and b;
    layer2_outputs(8191) <= not a;
    layer2_outputs(8192) <= not a;
    layer2_outputs(8193) <= not (a or b);
    layer2_outputs(8194) <= a or b;
    layer2_outputs(8195) <= b and not a;
    layer2_outputs(8196) <= b;
    layer2_outputs(8197) <= a or b;
    layer2_outputs(8198) <= a or b;
    layer2_outputs(8199) <= a and not b;
    layer2_outputs(8200) <= not a;
    layer2_outputs(8201) <= b;
    layer2_outputs(8202) <= a;
    layer2_outputs(8203) <= a and b;
    layer2_outputs(8204) <= b;
    layer2_outputs(8205) <= not a;
    layer2_outputs(8206) <= not (a and b);
    layer2_outputs(8207) <= not a;
    layer2_outputs(8208) <= a or b;
    layer2_outputs(8209) <= not a;
    layer2_outputs(8210) <= a;
    layer2_outputs(8211) <= not b;
    layer2_outputs(8212) <= a;
    layer2_outputs(8213) <= a and b;
    layer2_outputs(8214) <= a and b;
    layer2_outputs(8215) <= a and not b;
    layer2_outputs(8216) <= a;
    layer2_outputs(8217) <= a or b;
    layer2_outputs(8218) <= a and not b;
    layer2_outputs(8219) <= not b;
    layer2_outputs(8220) <= b;
    layer2_outputs(8221) <= not b;
    layer2_outputs(8222) <= not b;
    layer2_outputs(8223) <= a and b;
    layer2_outputs(8224) <= not a;
    layer2_outputs(8225) <= a xor b;
    layer2_outputs(8226) <= a;
    layer2_outputs(8227) <= not b;
    layer2_outputs(8228) <= not a;
    layer2_outputs(8229) <= b and not a;
    layer2_outputs(8230) <= not (a or b);
    layer2_outputs(8231) <= a;
    layer2_outputs(8232) <= a;
    layer2_outputs(8233) <= not (a or b);
    layer2_outputs(8234) <= not b or a;
    layer2_outputs(8235) <= not (a xor b);
    layer2_outputs(8236) <= a;
    layer2_outputs(8237) <= a and not b;
    layer2_outputs(8238) <= b;
    layer2_outputs(8239) <= not a;
    layer2_outputs(8240) <= not a;
    layer2_outputs(8241) <= not b;
    layer2_outputs(8242) <= a and not b;
    layer2_outputs(8243) <= b;
    layer2_outputs(8244) <= not b;
    layer2_outputs(8245) <= a;
    layer2_outputs(8246) <= not a;
    layer2_outputs(8247) <= not a;
    layer2_outputs(8248) <= a or b;
    layer2_outputs(8249) <= a;
    layer2_outputs(8250) <= a;
    layer2_outputs(8251) <= a xor b;
    layer2_outputs(8252) <= not a or b;
    layer2_outputs(8253) <= a and b;
    layer2_outputs(8254) <= b and not a;
    layer2_outputs(8255) <= a xor b;
    layer2_outputs(8256) <= not (a xor b);
    layer2_outputs(8257) <= not a;
    layer2_outputs(8258) <= not a or b;
    layer2_outputs(8259) <= a;
    layer2_outputs(8260) <= a or b;
    layer2_outputs(8261) <= not b;
    layer2_outputs(8262) <= a xor b;
    layer2_outputs(8263) <= not (a xor b);
    layer2_outputs(8264) <= not b;
    layer2_outputs(8265) <= not a;
    layer2_outputs(8266) <= a and b;
    layer2_outputs(8267) <= not a or b;
    layer2_outputs(8268) <= a;
    layer2_outputs(8269) <= not (a or b);
    layer2_outputs(8270) <= a and b;
    layer2_outputs(8271) <= a or b;
    layer2_outputs(8272) <= b and not a;
    layer2_outputs(8273) <= not b or a;
    layer2_outputs(8274) <= not b or a;
    layer2_outputs(8275) <= not b;
    layer2_outputs(8276) <= b;
    layer2_outputs(8277) <= a;
    layer2_outputs(8278) <= a;
    layer2_outputs(8279) <= not (a and b);
    layer2_outputs(8280) <= not a;
    layer2_outputs(8281) <= not (a or b);
    layer2_outputs(8282) <= a xor b;
    layer2_outputs(8283) <= not b;
    layer2_outputs(8284) <= not (a xor b);
    layer2_outputs(8285) <= b and not a;
    layer2_outputs(8286) <= not b;
    layer2_outputs(8287) <= not a or b;
    layer2_outputs(8288) <= not b or a;
    layer2_outputs(8289) <= not b or a;
    layer2_outputs(8290) <= a or b;
    layer2_outputs(8291) <= a or b;
    layer2_outputs(8292) <= b;
    layer2_outputs(8293) <= b and not a;
    layer2_outputs(8294) <= b and not a;
    layer2_outputs(8295) <= not (a xor b);
    layer2_outputs(8296) <= not b;
    layer2_outputs(8297) <= not b;
    layer2_outputs(8298) <= a;
    layer2_outputs(8299) <= not (a or b);
    layer2_outputs(8300) <= not b or a;
    layer2_outputs(8301) <= not b or a;
    layer2_outputs(8302) <= b;
    layer2_outputs(8303) <= a xor b;
    layer2_outputs(8304) <= b;
    layer2_outputs(8305) <= not a;
    layer2_outputs(8306) <= 1'b1;
    layer2_outputs(8307) <= not a or b;
    layer2_outputs(8308) <= not a or b;
    layer2_outputs(8309) <= a and b;
    layer2_outputs(8310) <= a and b;
    layer2_outputs(8311) <= not (a xor b);
    layer2_outputs(8312) <= a and b;
    layer2_outputs(8313) <= 1'b0;
    layer2_outputs(8314) <= a;
    layer2_outputs(8315) <= not a or b;
    layer2_outputs(8316) <= not b;
    layer2_outputs(8317) <= not b or a;
    layer2_outputs(8318) <= a;
    layer2_outputs(8319) <= not (a and b);
    layer2_outputs(8320) <= not (a and b);
    layer2_outputs(8321) <= not (a and b);
    layer2_outputs(8322) <= not a;
    layer2_outputs(8323) <= not (a and b);
    layer2_outputs(8324) <= b and not a;
    layer2_outputs(8325) <= not (a and b);
    layer2_outputs(8326) <= not (a or b);
    layer2_outputs(8327) <= not (a or b);
    layer2_outputs(8328) <= not a;
    layer2_outputs(8329) <= a or b;
    layer2_outputs(8330) <= not b;
    layer2_outputs(8331) <= b;
    layer2_outputs(8332) <= not (a or b);
    layer2_outputs(8333) <= not b;
    layer2_outputs(8334) <= not (a or b);
    layer2_outputs(8335) <= b and not a;
    layer2_outputs(8336) <= not a or b;
    layer2_outputs(8337) <= not (a or b);
    layer2_outputs(8338) <= a;
    layer2_outputs(8339) <= not a;
    layer2_outputs(8340) <= a and b;
    layer2_outputs(8341) <= a;
    layer2_outputs(8342) <= not (a and b);
    layer2_outputs(8343) <= a;
    layer2_outputs(8344) <= a and b;
    layer2_outputs(8345) <= a or b;
    layer2_outputs(8346) <= not a or b;
    layer2_outputs(8347) <= a;
    layer2_outputs(8348) <= 1'b1;
    layer2_outputs(8349) <= not b;
    layer2_outputs(8350) <= a xor b;
    layer2_outputs(8351) <= a xor b;
    layer2_outputs(8352) <= a and b;
    layer2_outputs(8353) <= 1'b0;
    layer2_outputs(8354) <= not b;
    layer2_outputs(8355) <= not (a and b);
    layer2_outputs(8356) <= not b;
    layer2_outputs(8357) <= a;
    layer2_outputs(8358) <= 1'b0;
    layer2_outputs(8359) <= not (a and b);
    layer2_outputs(8360) <= b;
    layer2_outputs(8361) <= not a or b;
    layer2_outputs(8362) <= a;
    layer2_outputs(8363) <= not b;
    layer2_outputs(8364) <= a and not b;
    layer2_outputs(8365) <= not (a or b);
    layer2_outputs(8366) <= a;
    layer2_outputs(8367) <= a;
    layer2_outputs(8368) <= not (a and b);
    layer2_outputs(8369) <= not (a xor b);
    layer2_outputs(8370) <= not b or a;
    layer2_outputs(8371) <= b and not a;
    layer2_outputs(8372) <= a xor b;
    layer2_outputs(8373) <= a and not b;
    layer2_outputs(8374) <= not b;
    layer2_outputs(8375) <= not b or a;
    layer2_outputs(8376) <= not b;
    layer2_outputs(8377) <= a and not b;
    layer2_outputs(8378) <= a;
    layer2_outputs(8379) <= not (a xor b);
    layer2_outputs(8380) <= not b or a;
    layer2_outputs(8381) <= a and b;
    layer2_outputs(8382) <= not b;
    layer2_outputs(8383) <= not a;
    layer2_outputs(8384) <= not (a or b);
    layer2_outputs(8385) <= not (a and b);
    layer2_outputs(8386) <= not (a xor b);
    layer2_outputs(8387) <= a and not b;
    layer2_outputs(8388) <= a and b;
    layer2_outputs(8389) <= a xor b;
    layer2_outputs(8390) <= a;
    layer2_outputs(8391) <= not (a or b);
    layer2_outputs(8392) <= not (a and b);
    layer2_outputs(8393) <= b and not a;
    layer2_outputs(8394) <= b;
    layer2_outputs(8395) <= a and not b;
    layer2_outputs(8396) <= not (a xor b);
    layer2_outputs(8397) <= not a or b;
    layer2_outputs(8398) <= not (a or b);
    layer2_outputs(8399) <= not (a xor b);
    layer2_outputs(8400) <= b and not a;
    layer2_outputs(8401) <= 1'b1;
    layer2_outputs(8402) <= a or b;
    layer2_outputs(8403) <= a and not b;
    layer2_outputs(8404) <= a;
    layer2_outputs(8405) <= not a or b;
    layer2_outputs(8406) <= a;
    layer2_outputs(8407) <= a and not b;
    layer2_outputs(8408) <= a;
    layer2_outputs(8409) <= not b or a;
    layer2_outputs(8410) <= not (a or b);
    layer2_outputs(8411) <= not b;
    layer2_outputs(8412) <= not a;
    layer2_outputs(8413) <= not (a or b);
    layer2_outputs(8414) <= not a or b;
    layer2_outputs(8415) <= b;
    layer2_outputs(8416) <= a and b;
    layer2_outputs(8417) <= a and b;
    layer2_outputs(8418) <= a or b;
    layer2_outputs(8419) <= b;
    layer2_outputs(8420) <= not b;
    layer2_outputs(8421) <= not b or a;
    layer2_outputs(8422) <= not b;
    layer2_outputs(8423) <= not (a and b);
    layer2_outputs(8424) <= not a or b;
    layer2_outputs(8425) <= not a or b;
    layer2_outputs(8426) <= a or b;
    layer2_outputs(8427) <= a or b;
    layer2_outputs(8428) <= a;
    layer2_outputs(8429) <= a xor b;
    layer2_outputs(8430) <= b;
    layer2_outputs(8431) <= not a or b;
    layer2_outputs(8432) <= not a or b;
    layer2_outputs(8433) <= b;
    layer2_outputs(8434) <= not (a xor b);
    layer2_outputs(8435) <= not b;
    layer2_outputs(8436) <= not (a or b);
    layer2_outputs(8437) <= b;
    layer2_outputs(8438) <= not (a and b);
    layer2_outputs(8439) <= not a;
    layer2_outputs(8440) <= not b;
    layer2_outputs(8441) <= b and not a;
    layer2_outputs(8442) <= a and b;
    layer2_outputs(8443) <= not a;
    layer2_outputs(8444) <= a or b;
    layer2_outputs(8445) <= not (a xor b);
    layer2_outputs(8446) <= not a;
    layer2_outputs(8447) <= a;
    layer2_outputs(8448) <= not a;
    layer2_outputs(8449) <= not b;
    layer2_outputs(8450) <= not (a or b);
    layer2_outputs(8451) <= a;
    layer2_outputs(8452) <= not (a and b);
    layer2_outputs(8453) <= not (a and b);
    layer2_outputs(8454) <= not b;
    layer2_outputs(8455) <= a and b;
    layer2_outputs(8456) <= not (a and b);
    layer2_outputs(8457) <= not a;
    layer2_outputs(8458) <= not b;
    layer2_outputs(8459) <= not (a xor b);
    layer2_outputs(8460) <= b;
    layer2_outputs(8461) <= not (a xor b);
    layer2_outputs(8462) <= not b;
    layer2_outputs(8463) <= not b or a;
    layer2_outputs(8464) <= b and not a;
    layer2_outputs(8465) <= a;
    layer2_outputs(8466) <= a and not b;
    layer2_outputs(8467) <= 1'b0;
    layer2_outputs(8468) <= not b;
    layer2_outputs(8469) <= b;
    layer2_outputs(8470) <= a or b;
    layer2_outputs(8471) <= a;
    layer2_outputs(8472) <= not a or b;
    layer2_outputs(8473) <= not (a xor b);
    layer2_outputs(8474) <= not (a and b);
    layer2_outputs(8475) <= not b;
    layer2_outputs(8476) <= not (a and b);
    layer2_outputs(8477) <= a and not b;
    layer2_outputs(8478) <= not (a and b);
    layer2_outputs(8479) <= not (a xor b);
    layer2_outputs(8480) <= not (a or b);
    layer2_outputs(8481) <= not a or b;
    layer2_outputs(8482) <= a and b;
    layer2_outputs(8483) <= not b;
    layer2_outputs(8484) <= not a;
    layer2_outputs(8485) <= not a;
    layer2_outputs(8486) <= not (a and b);
    layer2_outputs(8487) <= not a;
    layer2_outputs(8488) <= a xor b;
    layer2_outputs(8489) <= a;
    layer2_outputs(8490) <= a xor b;
    layer2_outputs(8491) <= 1'b0;
    layer2_outputs(8492) <= a;
    layer2_outputs(8493) <= 1'b1;
    layer2_outputs(8494) <= b and not a;
    layer2_outputs(8495) <= b and not a;
    layer2_outputs(8496) <= b and not a;
    layer2_outputs(8497) <= b;
    layer2_outputs(8498) <= not a or b;
    layer2_outputs(8499) <= not (a or b);
    layer2_outputs(8500) <= a xor b;
    layer2_outputs(8501) <= b;
    layer2_outputs(8502) <= a and b;
    layer2_outputs(8503) <= not a;
    layer2_outputs(8504) <= a xor b;
    layer2_outputs(8505) <= not a;
    layer2_outputs(8506) <= b;
    layer2_outputs(8507) <= not a or b;
    layer2_outputs(8508) <= not (a or b);
    layer2_outputs(8509) <= not b;
    layer2_outputs(8510) <= b;
    layer2_outputs(8511) <= not (a and b);
    layer2_outputs(8512) <= a and not b;
    layer2_outputs(8513) <= a and b;
    layer2_outputs(8514) <= a;
    layer2_outputs(8515) <= a or b;
    layer2_outputs(8516) <= not a;
    layer2_outputs(8517) <= a and not b;
    layer2_outputs(8518) <= not a;
    layer2_outputs(8519) <= b;
    layer2_outputs(8520) <= not (a and b);
    layer2_outputs(8521) <= b;
    layer2_outputs(8522) <= a and b;
    layer2_outputs(8523) <= not a;
    layer2_outputs(8524) <= a xor b;
    layer2_outputs(8525) <= not b or a;
    layer2_outputs(8526) <= not a;
    layer2_outputs(8527) <= not a or b;
    layer2_outputs(8528) <= a and b;
    layer2_outputs(8529) <= a or b;
    layer2_outputs(8530) <= a;
    layer2_outputs(8531) <= a;
    layer2_outputs(8532) <= a and b;
    layer2_outputs(8533) <= not (a or b);
    layer2_outputs(8534) <= a;
    layer2_outputs(8535) <= a;
    layer2_outputs(8536) <= a and b;
    layer2_outputs(8537) <= a and not b;
    layer2_outputs(8538) <= b;
    layer2_outputs(8539) <= not a;
    layer2_outputs(8540) <= a and b;
    layer2_outputs(8541) <= a and not b;
    layer2_outputs(8542) <= not a;
    layer2_outputs(8543) <= not (a or b);
    layer2_outputs(8544) <= b;
    layer2_outputs(8545) <= not (a and b);
    layer2_outputs(8546) <= a or b;
    layer2_outputs(8547) <= b;
    layer2_outputs(8548) <= a;
    layer2_outputs(8549) <= 1'b0;
    layer2_outputs(8550) <= not b;
    layer2_outputs(8551) <= b and not a;
    layer2_outputs(8552) <= not a or b;
    layer2_outputs(8553) <= a and not b;
    layer2_outputs(8554) <= a;
    layer2_outputs(8555) <= not a;
    layer2_outputs(8556) <= a or b;
    layer2_outputs(8557) <= b;
    layer2_outputs(8558) <= not (a or b);
    layer2_outputs(8559) <= not b or a;
    layer2_outputs(8560) <= not b or a;
    layer2_outputs(8561) <= not a or b;
    layer2_outputs(8562) <= not a;
    layer2_outputs(8563) <= not a;
    layer2_outputs(8564) <= not (a or b);
    layer2_outputs(8565) <= not b;
    layer2_outputs(8566) <= b;
    layer2_outputs(8567) <= b;
    layer2_outputs(8568) <= a and not b;
    layer2_outputs(8569) <= a or b;
    layer2_outputs(8570) <= not (a or b);
    layer2_outputs(8571) <= not (a xor b);
    layer2_outputs(8572) <= not a;
    layer2_outputs(8573) <= b;
    layer2_outputs(8574) <= not b;
    layer2_outputs(8575) <= a xor b;
    layer2_outputs(8576) <= not b;
    layer2_outputs(8577) <= not (a or b);
    layer2_outputs(8578) <= b;
    layer2_outputs(8579) <= 1'b0;
    layer2_outputs(8580) <= not b;
    layer2_outputs(8581) <= not a or b;
    layer2_outputs(8582) <= b and not a;
    layer2_outputs(8583) <= b;
    layer2_outputs(8584) <= not (a and b);
    layer2_outputs(8585) <= not (a and b);
    layer2_outputs(8586) <= b and not a;
    layer2_outputs(8587) <= a and b;
    layer2_outputs(8588) <= not a;
    layer2_outputs(8589) <= not (a and b);
    layer2_outputs(8590) <= not b;
    layer2_outputs(8591) <= not b or a;
    layer2_outputs(8592) <= not a;
    layer2_outputs(8593) <= a and not b;
    layer2_outputs(8594) <= not (a xor b);
    layer2_outputs(8595) <= b;
    layer2_outputs(8596) <= a and b;
    layer2_outputs(8597) <= a;
    layer2_outputs(8598) <= a;
    layer2_outputs(8599) <= b;
    layer2_outputs(8600) <= not a or b;
    layer2_outputs(8601) <= a and not b;
    layer2_outputs(8602) <= a xor b;
    layer2_outputs(8603) <= not (a and b);
    layer2_outputs(8604) <= not a;
    layer2_outputs(8605) <= not a;
    layer2_outputs(8606) <= a and not b;
    layer2_outputs(8607) <= not a;
    layer2_outputs(8608) <= not a or b;
    layer2_outputs(8609) <= b and not a;
    layer2_outputs(8610) <= a xor b;
    layer2_outputs(8611) <= not b or a;
    layer2_outputs(8612) <= a and not b;
    layer2_outputs(8613) <= a and not b;
    layer2_outputs(8614) <= a and not b;
    layer2_outputs(8615) <= a;
    layer2_outputs(8616) <= not b;
    layer2_outputs(8617) <= not (a xor b);
    layer2_outputs(8618) <= not (a and b);
    layer2_outputs(8619) <= not a;
    layer2_outputs(8620) <= a;
    layer2_outputs(8621) <= a or b;
    layer2_outputs(8622) <= a xor b;
    layer2_outputs(8623) <= 1'b0;
    layer2_outputs(8624) <= 1'b0;
    layer2_outputs(8625) <= a and b;
    layer2_outputs(8626) <= not b;
    layer2_outputs(8627) <= not a or b;
    layer2_outputs(8628) <= b;
    layer2_outputs(8629) <= not (a or b);
    layer2_outputs(8630) <= not b;
    layer2_outputs(8631) <= a and not b;
    layer2_outputs(8632) <= not b;
    layer2_outputs(8633) <= 1'b0;
    layer2_outputs(8634) <= not b;
    layer2_outputs(8635) <= b;
    layer2_outputs(8636) <= a or b;
    layer2_outputs(8637) <= a and not b;
    layer2_outputs(8638) <= 1'b1;
    layer2_outputs(8639) <= b;
    layer2_outputs(8640) <= not (a and b);
    layer2_outputs(8641) <= a and b;
    layer2_outputs(8642) <= not b;
    layer2_outputs(8643) <= a xor b;
    layer2_outputs(8644) <= not (a xor b);
    layer2_outputs(8645) <= not b;
    layer2_outputs(8646) <= not b;
    layer2_outputs(8647) <= b;
    layer2_outputs(8648) <= b;
    layer2_outputs(8649) <= not a or b;
    layer2_outputs(8650) <= a or b;
    layer2_outputs(8651) <= not (a xor b);
    layer2_outputs(8652) <= a or b;
    layer2_outputs(8653) <= a and not b;
    layer2_outputs(8654) <= a and not b;
    layer2_outputs(8655) <= not b or a;
    layer2_outputs(8656) <= 1'b0;
    layer2_outputs(8657) <= not b;
    layer2_outputs(8658) <= a or b;
    layer2_outputs(8659) <= not a;
    layer2_outputs(8660) <= not (a or b);
    layer2_outputs(8661) <= not (a or b);
    layer2_outputs(8662) <= a or b;
    layer2_outputs(8663) <= a and not b;
    layer2_outputs(8664) <= a;
    layer2_outputs(8665) <= a;
    layer2_outputs(8666) <= a and not b;
    layer2_outputs(8667) <= a and not b;
    layer2_outputs(8668) <= not a;
    layer2_outputs(8669) <= not b;
    layer2_outputs(8670) <= not (a and b);
    layer2_outputs(8671) <= not a or b;
    layer2_outputs(8672) <= b;
    layer2_outputs(8673) <= a;
    layer2_outputs(8674) <= not b or a;
    layer2_outputs(8675) <= not (a or b);
    layer2_outputs(8676) <= not (a xor b);
    layer2_outputs(8677) <= not b or a;
    layer2_outputs(8678) <= a xor b;
    layer2_outputs(8679) <= not (a or b);
    layer2_outputs(8680) <= not (a xor b);
    layer2_outputs(8681) <= a;
    layer2_outputs(8682) <= not b;
    layer2_outputs(8683) <= a xor b;
    layer2_outputs(8684) <= a and b;
    layer2_outputs(8685) <= not b;
    layer2_outputs(8686) <= not (a or b);
    layer2_outputs(8687) <= a and b;
    layer2_outputs(8688) <= a or b;
    layer2_outputs(8689) <= b;
    layer2_outputs(8690) <= not a;
    layer2_outputs(8691) <= a or b;
    layer2_outputs(8692) <= b;
    layer2_outputs(8693) <= not a;
    layer2_outputs(8694) <= not (a or b);
    layer2_outputs(8695) <= not a or b;
    layer2_outputs(8696) <= a;
    layer2_outputs(8697) <= not b or a;
    layer2_outputs(8698) <= not a or b;
    layer2_outputs(8699) <= not b or a;
    layer2_outputs(8700) <= a and b;
    layer2_outputs(8701) <= not b;
    layer2_outputs(8702) <= a and b;
    layer2_outputs(8703) <= not a or b;
    layer2_outputs(8704) <= a;
    layer2_outputs(8705) <= a and b;
    layer2_outputs(8706) <= not a;
    layer2_outputs(8707) <= not (a and b);
    layer2_outputs(8708) <= b and not a;
    layer2_outputs(8709) <= not a;
    layer2_outputs(8710) <= a;
    layer2_outputs(8711) <= a or b;
    layer2_outputs(8712) <= not (a or b);
    layer2_outputs(8713) <= b and not a;
    layer2_outputs(8714) <= a and b;
    layer2_outputs(8715) <= a xor b;
    layer2_outputs(8716) <= not b;
    layer2_outputs(8717) <= a and not b;
    layer2_outputs(8718) <= not b or a;
    layer2_outputs(8719) <= not (a and b);
    layer2_outputs(8720) <= not (a xor b);
    layer2_outputs(8721) <= not b;
    layer2_outputs(8722) <= not (a or b);
    layer2_outputs(8723) <= not (a xor b);
    layer2_outputs(8724) <= a and b;
    layer2_outputs(8725) <= not (a or b);
    layer2_outputs(8726) <= not b;
    layer2_outputs(8727) <= a;
    layer2_outputs(8728) <= a xor b;
    layer2_outputs(8729) <= a and not b;
    layer2_outputs(8730) <= a and b;
    layer2_outputs(8731) <= a;
    layer2_outputs(8732) <= b;
    layer2_outputs(8733) <= a and not b;
    layer2_outputs(8734) <= not (a xor b);
    layer2_outputs(8735) <= not b;
    layer2_outputs(8736) <= not a;
    layer2_outputs(8737) <= not (a or b);
    layer2_outputs(8738) <= a and not b;
    layer2_outputs(8739) <= not a or b;
    layer2_outputs(8740) <= 1'b0;
    layer2_outputs(8741) <= not (a or b);
    layer2_outputs(8742) <= not b or a;
    layer2_outputs(8743) <= 1'b1;
    layer2_outputs(8744) <= 1'b0;
    layer2_outputs(8745) <= not (a xor b);
    layer2_outputs(8746) <= not b;
    layer2_outputs(8747) <= not b;
    layer2_outputs(8748) <= not (a and b);
    layer2_outputs(8749) <= not b;
    layer2_outputs(8750) <= b;
    layer2_outputs(8751) <= b and not a;
    layer2_outputs(8752) <= b and not a;
    layer2_outputs(8753) <= not b or a;
    layer2_outputs(8754) <= a xor b;
    layer2_outputs(8755) <= b;
    layer2_outputs(8756) <= a or b;
    layer2_outputs(8757) <= b;
    layer2_outputs(8758) <= not b;
    layer2_outputs(8759) <= not (a and b);
    layer2_outputs(8760) <= b;
    layer2_outputs(8761) <= not b;
    layer2_outputs(8762) <= not b;
    layer2_outputs(8763) <= a and not b;
    layer2_outputs(8764) <= a or b;
    layer2_outputs(8765) <= a or b;
    layer2_outputs(8766) <= not a;
    layer2_outputs(8767) <= b and not a;
    layer2_outputs(8768) <= b;
    layer2_outputs(8769) <= a or b;
    layer2_outputs(8770) <= 1'b1;
    layer2_outputs(8771) <= a or b;
    layer2_outputs(8772) <= not b or a;
    layer2_outputs(8773) <= a xor b;
    layer2_outputs(8774) <= b and not a;
    layer2_outputs(8775) <= not a or b;
    layer2_outputs(8776) <= not a;
    layer2_outputs(8777) <= 1'b0;
    layer2_outputs(8778) <= a or b;
    layer2_outputs(8779) <= not (a or b);
    layer2_outputs(8780) <= b;
    layer2_outputs(8781) <= a;
    layer2_outputs(8782) <= b and not a;
    layer2_outputs(8783) <= not (a or b);
    layer2_outputs(8784) <= not a;
    layer2_outputs(8785) <= not (a and b);
    layer2_outputs(8786) <= a;
    layer2_outputs(8787) <= b;
    layer2_outputs(8788) <= not (a xor b);
    layer2_outputs(8789) <= not (a and b);
    layer2_outputs(8790) <= a xor b;
    layer2_outputs(8791) <= not a;
    layer2_outputs(8792) <= a and not b;
    layer2_outputs(8793) <= not a or b;
    layer2_outputs(8794) <= not (a or b);
    layer2_outputs(8795) <= b;
    layer2_outputs(8796) <= a or b;
    layer2_outputs(8797) <= a xor b;
    layer2_outputs(8798) <= not (a and b);
    layer2_outputs(8799) <= a or b;
    layer2_outputs(8800) <= not a;
    layer2_outputs(8801) <= 1'b0;
    layer2_outputs(8802) <= a;
    layer2_outputs(8803) <= not a;
    layer2_outputs(8804) <= b and not a;
    layer2_outputs(8805) <= a xor b;
    layer2_outputs(8806) <= a and not b;
    layer2_outputs(8807) <= not (a and b);
    layer2_outputs(8808) <= not a;
    layer2_outputs(8809) <= a and not b;
    layer2_outputs(8810) <= a and not b;
    layer2_outputs(8811) <= not (a and b);
    layer2_outputs(8812) <= not b;
    layer2_outputs(8813) <= not b;
    layer2_outputs(8814) <= not a;
    layer2_outputs(8815) <= a xor b;
    layer2_outputs(8816) <= a and b;
    layer2_outputs(8817) <= not (a or b);
    layer2_outputs(8818) <= a;
    layer2_outputs(8819) <= a and not b;
    layer2_outputs(8820) <= a;
    layer2_outputs(8821) <= a xor b;
    layer2_outputs(8822) <= a or b;
    layer2_outputs(8823) <= not b;
    layer2_outputs(8824) <= a and not b;
    layer2_outputs(8825) <= a and not b;
    layer2_outputs(8826) <= b;
    layer2_outputs(8827) <= not b;
    layer2_outputs(8828) <= 1'b0;
    layer2_outputs(8829) <= not a or b;
    layer2_outputs(8830) <= a and not b;
    layer2_outputs(8831) <= 1'b0;
    layer2_outputs(8832) <= not a or b;
    layer2_outputs(8833) <= not (a xor b);
    layer2_outputs(8834) <= a or b;
    layer2_outputs(8835) <= not (a or b);
    layer2_outputs(8836) <= a xor b;
    layer2_outputs(8837) <= not (a and b);
    layer2_outputs(8838) <= 1'b0;
    layer2_outputs(8839) <= not a;
    layer2_outputs(8840) <= not b;
    layer2_outputs(8841) <= not (a xor b);
    layer2_outputs(8842) <= not a;
    layer2_outputs(8843) <= not (a and b);
    layer2_outputs(8844) <= b;
    layer2_outputs(8845) <= b;
    layer2_outputs(8846) <= not (a or b);
    layer2_outputs(8847) <= a or b;
    layer2_outputs(8848) <= 1'b0;
    layer2_outputs(8849) <= not (a xor b);
    layer2_outputs(8850) <= not (a or b);
    layer2_outputs(8851) <= a or b;
    layer2_outputs(8852) <= not (a or b);
    layer2_outputs(8853) <= not a;
    layer2_outputs(8854) <= a or b;
    layer2_outputs(8855) <= not (a or b);
    layer2_outputs(8856) <= not a;
    layer2_outputs(8857) <= not (a and b);
    layer2_outputs(8858) <= not b or a;
    layer2_outputs(8859) <= b;
    layer2_outputs(8860) <= not (a xor b);
    layer2_outputs(8861) <= b and not a;
    layer2_outputs(8862) <= not (a or b);
    layer2_outputs(8863) <= not a;
    layer2_outputs(8864) <= not b;
    layer2_outputs(8865) <= not a;
    layer2_outputs(8866) <= a and b;
    layer2_outputs(8867) <= a and not b;
    layer2_outputs(8868) <= a xor b;
    layer2_outputs(8869) <= a;
    layer2_outputs(8870) <= not (a xor b);
    layer2_outputs(8871) <= a xor b;
    layer2_outputs(8872) <= not (a or b);
    layer2_outputs(8873) <= b and not a;
    layer2_outputs(8874) <= not b;
    layer2_outputs(8875) <= a xor b;
    layer2_outputs(8876) <= a xor b;
    layer2_outputs(8877) <= not a;
    layer2_outputs(8878) <= a;
    layer2_outputs(8879) <= b;
    layer2_outputs(8880) <= a;
    layer2_outputs(8881) <= not (a and b);
    layer2_outputs(8882) <= a;
    layer2_outputs(8883) <= not (a or b);
    layer2_outputs(8884) <= a and not b;
    layer2_outputs(8885) <= not (a or b);
    layer2_outputs(8886) <= a and b;
    layer2_outputs(8887) <= not a;
    layer2_outputs(8888) <= not a or b;
    layer2_outputs(8889) <= not a or b;
    layer2_outputs(8890) <= a or b;
    layer2_outputs(8891) <= a or b;
    layer2_outputs(8892) <= b;
    layer2_outputs(8893) <= not b;
    layer2_outputs(8894) <= not (a xor b);
    layer2_outputs(8895) <= not (a xor b);
    layer2_outputs(8896) <= 1'b0;
    layer2_outputs(8897) <= b;
    layer2_outputs(8898) <= not b;
    layer2_outputs(8899) <= b;
    layer2_outputs(8900) <= b;
    layer2_outputs(8901) <= a and b;
    layer2_outputs(8902) <= b and not a;
    layer2_outputs(8903) <= not a;
    layer2_outputs(8904) <= b and not a;
    layer2_outputs(8905) <= not b;
    layer2_outputs(8906) <= not b;
    layer2_outputs(8907) <= not b;
    layer2_outputs(8908) <= not b;
    layer2_outputs(8909) <= 1'b0;
    layer2_outputs(8910) <= a and b;
    layer2_outputs(8911) <= not (a and b);
    layer2_outputs(8912) <= not b;
    layer2_outputs(8913) <= a and b;
    layer2_outputs(8914) <= a xor b;
    layer2_outputs(8915) <= a xor b;
    layer2_outputs(8916) <= a and b;
    layer2_outputs(8917) <= not (a or b);
    layer2_outputs(8918) <= not (a and b);
    layer2_outputs(8919) <= not b or a;
    layer2_outputs(8920) <= a and not b;
    layer2_outputs(8921) <= not a;
    layer2_outputs(8922) <= a or b;
    layer2_outputs(8923) <= not b;
    layer2_outputs(8924) <= not (a or b);
    layer2_outputs(8925) <= a and not b;
    layer2_outputs(8926) <= not (a and b);
    layer2_outputs(8927) <= 1'b1;
    layer2_outputs(8928) <= a or b;
    layer2_outputs(8929) <= a and b;
    layer2_outputs(8930) <= not (a or b);
    layer2_outputs(8931) <= a and b;
    layer2_outputs(8932) <= not (a xor b);
    layer2_outputs(8933) <= a or b;
    layer2_outputs(8934) <= a;
    layer2_outputs(8935) <= a;
    layer2_outputs(8936) <= not (a xor b);
    layer2_outputs(8937) <= b and not a;
    layer2_outputs(8938) <= not (a xor b);
    layer2_outputs(8939) <= not b or a;
    layer2_outputs(8940) <= a and not b;
    layer2_outputs(8941) <= a;
    layer2_outputs(8942) <= not a or b;
    layer2_outputs(8943) <= not b;
    layer2_outputs(8944) <= not b or a;
    layer2_outputs(8945) <= not (a or b);
    layer2_outputs(8946) <= a and b;
    layer2_outputs(8947) <= not a or b;
    layer2_outputs(8948) <= b;
    layer2_outputs(8949) <= b and not a;
    layer2_outputs(8950) <= not a;
    layer2_outputs(8951) <= not (a xor b);
    layer2_outputs(8952) <= not a;
    layer2_outputs(8953) <= not b;
    layer2_outputs(8954) <= not b or a;
    layer2_outputs(8955) <= b and not a;
    layer2_outputs(8956) <= b and not a;
    layer2_outputs(8957) <= a and b;
    layer2_outputs(8958) <= a;
    layer2_outputs(8959) <= b;
    layer2_outputs(8960) <= b;
    layer2_outputs(8961) <= not a;
    layer2_outputs(8962) <= not (a or b);
    layer2_outputs(8963) <= not a or b;
    layer2_outputs(8964) <= a or b;
    layer2_outputs(8965) <= a xor b;
    layer2_outputs(8966) <= a or b;
    layer2_outputs(8967) <= not b;
    layer2_outputs(8968) <= b and not a;
    layer2_outputs(8969) <= not a;
    layer2_outputs(8970) <= not b;
    layer2_outputs(8971) <= b and not a;
    layer2_outputs(8972) <= not (a and b);
    layer2_outputs(8973) <= not (a or b);
    layer2_outputs(8974) <= not (a or b);
    layer2_outputs(8975) <= not (a xor b);
    layer2_outputs(8976) <= b and not a;
    layer2_outputs(8977) <= a or b;
    layer2_outputs(8978) <= not b or a;
    layer2_outputs(8979) <= not (a or b);
    layer2_outputs(8980) <= not (a or b);
    layer2_outputs(8981) <= a and not b;
    layer2_outputs(8982) <= a;
    layer2_outputs(8983) <= a and b;
    layer2_outputs(8984) <= a and b;
    layer2_outputs(8985) <= not a;
    layer2_outputs(8986) <= a;
    layer2_outputs(8987) <= not a;
    layer2_outputs(8988) <= not (a or b);
    layer2_outputs(8989) <= a or b;
    layer2_outputs(8990) <= not (a or b);
    layer2_outputs(8991) <= 1'b0;
    layer2_outputs(8992) <= b and not a;
    layer2_outputs(8993) <= not b;
    layer2_outputs(8994) <= b;
    layer2_outputs(8995) <= not (a or b);
    layer2_outputs(8996) <= b;
    layer2_outputs(8997) <= a or b;
    layer2_outputs(8998) <= not b;
    layer2_outputs(8999) <= a and b;
    layer2_outputs(9000) <= a;
    layer2_outputs(9001) <= b and not a;
    layer2_outputs(9002) <= not a;
    layer2_outputs(9003) <= not (a xor b);
    layer2_outputs(9004) <= b;
    layer2_outputs(9005) <= not (a or b);
    layer2_outputs(9006) <= not a;
    layer2_outputs(9007) <= b;
    layer2_outputs(9008) <= not (a and b);
    layer2_outputs(9009) <= a and b;
    layer2_outputs(9010) <= not (a and b);
    layer2_outputs(9011) <= not a or b;
    layer2_outputs(9012) <= b and not a;
    layer2_outputs(9013) <= a and not b;
    layer2_outputs(9014) <= a and not b;
    layer2_outputs(9015) <= a and b;
    layer2_outputs(9016) <= not a or b;
    layer2_outputs(9017) <= b and not a;
    layer2_outputs(9018) <= 1'b1;
    layer2_outputs(9019) <= not (a or b);
    layer2_outputs(9020) <= a and not b;
    layer2_outputs(9021) <= a and b;
    layer2_outputs(9022) <= not a or b;
    layer2_outputs(9023) <= b and not a;
    layer2_outputs(9024) <= not b or a;
    layer2_outputs(9025) <= a;
    layer2_outputs(9026) <= not (a xor b);
    layer2_outputs(9027) <= a;
    layer2_outputs(9028) <= not a;
    layer2_outputs(9029) <= not b or a;
    layer2_outputs(9030) <= not (a and b);
    layer2_outputs(9031) <= a;
    layer2_outputs(9032) <= not a or b;
    layer2_outputs(9033) <= 1'b0;
    layer2_outputs(9034) <= not b;
    layer2_outputs(9035) <= not (a and b);
    layer2_outputs(9036) <= not (a or b);
    layer2_outputs(9037) <= a;
    layer2_outputs(9038) <= b and not a;
    layer2_outputs(9039) <= not (a or b);
    layer2_outputs(9040) <= not b;
    layer2_outputs(9041) <= not a;
    layer2_outputs(9042) <= 1'b0;
    layer2_outputs(9043) <= not b;
    layer2_outputs(9044) <= a and b;
    layer2_outputs(9045) <= a and not b;
    layer2_outputs(9046) <= 1'b0;
    layer2_outputs(9047) <= not (a and b);
    layer2_outputs(9048) <= a or b;
    layer2_outputs(9049) <= not a;
    layer2_outputs(9050) <= b;
    layer2_outputs(9051) <= not b or a;
    layer2_outputs(9052) <= b and not a;
    layer2_outputs(9053) <= not (a or b);
    layer2_outputs(9054) <= a or b;
    layer2_outputs(9055) <= a;
    layer2_outputs(9056) <= b;
    layer2_outputs(9057) <= a and not b;
    layer2_outputs(9058) <= a or b;
    layer2_outputs(9059) <= b;
    layer2_outputs(9060) <= b;
    layer2_outputs(9061) <= not a;
    layer2_outputs(9062) <= a or b;
    layer2_outputs(9063) <= not (a or b);
    layer2_outputs(9064) <= a;
    layer2_outputs(9065) <= not a;
    layer2_outputs(9066) <= 1'b1;
    layer2_outputs(9067) <= b and not a;
    layer2_outputs(9068) <= a and not b;
    layer2_outputs(9069) <= not b;
    layer2_outputs(9070) <= 1'b0;
    layer2_outputs(9071) <= not b or a;
    layer2_outputs(9072) <= a;
    layer2_outputs(9073) <= a;
    layer2_outputs(9074) <= not (a xor b);
    layer2_outputs(9075) <= b;
    layer2_outputs(9076) <= not (a and b);
    layer2_outputs(9077) <= not a;
    layer2_outputs(9078) <= b and not a;
    layer2_outputs(9079) <= b;
    layer2_outputs(9080) <= not a;
    layer2_outputs(9081) <= a and b;
    layer2_outputs(9082) <= not (a and b);
    layer2_outputs(9083) <= a;
    layer2_outputs(9084) <= a and not b;
    layer2_outputs(9085) <= 1'b0;
    layer2_outputs(9086) <= a and b;
    layer2_outputs(9087) <= not b or a;
    layer2_outputs(9088) <= not b;
    layer2_outputs(9089) <= not b;
    layer2_outputs(9090) <= a or b;
    layer2_outputs(9091) <= not (a and b);
    layer2_outputs(9092) <= not a;
    layer2_outputs(9093) <= a or b;
    layer2_outputs(9094) <= b;
    layer2_outputs(9095) <= a and not b;
    layer2_outputs(9096) <= not a or b;
    layer2_outputs(9097) <= b;
    layer2_outputs(9098) <= a;
    layer2_outputs(9099) <= b;
    layer2_outputs(9100) <= a;
    layer2_outputs(9101) <= a;
    layer2_outputs(9102) <= not a;
    layer2_outputs(9103) <= not b;
    layer2_outputs(9104) <= a xor b;
    layer2_outputs(9105) <= a or b;
    layer2_outputs(9106) <= not (a or b);
    layer2_outputs(9107) <= not (a and b);
    layer2_outputs(9108) <= b and not a;
    layer2_outputs(9109) <= not b or a;
    layer2_outputs(9110) <= b;
    layer2_outputs(9111) <= a or b;
    layer2_outputs(9112) <= a xor b;
    layer2_outputs(9113) <= not (a and b);
    layer2_outputs(9114) <= not b or a;
    layer2_outputs(9115) <= not a or b;
    layer2_outputs(9116) <= not b;
    layer2_outputs(9117) <= a and b;
    layer2_outputs(9118) <= not b;
    layer2_outputs(9119) <= a and not b;
    layer2_outputs(9120) <= 1'b1;
    layer2_outputs(9121) <= not (a xor b);
    layer2_outputs(9122) <= not b or a;
    layer2_outputs(9123) <= a or b;
    layer2_outputs(9124) <= not b or a;
    layer2_outputs(9125) <= not (a or b);
    layer2_outputs(9126) <= a or b;
    layer2_outputs(9127) <= b;
    layer2_outputs(9128) <= not b or a;
    layer2_outputs(9129) <= not a or b;
    layer2_outputs(9130) <= not (a and b);
    layer2_outputs(9131) <= a and not b;
    layer2_outputs(9132) <= 1'b1;
    layer2_outputs(9133) <= not b or a;
    layer2_outputs(9134) <= 1'b1;
    layer2_outputs(9135) <= a xor b;
    layer2_outputs(9136) <= not a;
    layer2_outputs(9137) <= a;
    layer2_outputs(9138) <= a and b;
    layer2_outputs(9139) <= a;
    layer2_outputs(9140) <= not (a and b);
    layer2_outputs(9141) <= b;
    layer2_outputs(9142) <= b;
    layer2_outputs(9143) <= not (a and b);
    layer2_outputs(9144) <= b;
    layer2_outputs(9145) <= not (a and b);
    layer2_outputs(9146) <= a and not b;
    layer2_outputs(9147) <= not (a or b);
    layer2_outputs(9148) <= not (a xor b);
    layer2_outputs(9149) <= a;
    layer2_outputs(9150) <= not (a or b);
    layer2_outputs(9151) <= a and not b;
    layer2_outputs(9152) <= a and not b;
    layer2_outputs(9153) <= not a;
    layer2_outputs(9154) <= a and not b;
    layer2_outputs(9155) <= b and not a;
    layer2_outputs(9156) <= not a;
    layer2_outputs(9157) <= not (a and b);
    layer2_outputs(9158) <= a and b;
    layer2_outputs(9159) <= a;
    layer2_outputs(9160) <= a or b;
    layer2_outputs(9161) <= b;
    layer2_outputs(9162) <= a or b;
    layer2_outputs(9163) <= not (a and b);
    layer2_outputs(9164) <= not a or b;
    layer2_outputs(9165) <= not b or a;
    layer2_outputs(9166) <= not (a or b);
    layer2_outputs(9167) <= not (a and b);
    layer2_outputs(9168) <= a xor b;
    layer2_outputs(9169) <= b;
    layer2_outputs(9170) <= not b;
    layer2_outputs(9171) <= not (a and b);
    layer2_outputs(9172) <= b;
    layer2_outputs(9173) <= a;
    layer2_outputs(9174) <= not a;
    layer2_outputs(9175) <= not (a xor b);
    layer2_outputs(9176) <= a or b;
    layer2_outputs(9177) <= a or b;
    layer2_outputs(9178) <= b;
    layer2_outputs(9179) <= not (a or b);
    layer2_outputs(9180) <= b and not a;
    layer2_outputs(9181) <= not b;
    layer2_outputs(9182) <= not (a or b);
    layer2_outputs(9183) <= a and not b;
    layer2_outputs(9184) <= a or b;
    layer2_outputs(9185) <= a;
    layer2_outputs(9186) <= 1'b1;
    layer2_outputs(9187) <= not a;
    layer2_outputs(9188) <= not (a or b);
    layer2_outputs(9189) <= not b;
    layer2_outputs(9190) <= a and not b;
    layer2_outputs(9191) <= a and not b;
    layer2_outputs(9192) <= not a or b;
    layer2_outputs(9193) <= b and not a;
    layer2_outputs(9194) <= not (a and b);
    layer2_outputs(9195) <= a and not b;
    layer2_outputs(9196) <= not a or b;
    layer2_outputs(9197) <= 1'b1;
    layer2_outputs(9198) <= not b or a;
    layer2_outputs(9199) <= b;
    layer2_outputs(9200) <= not b or a;
    layer2_outputs(9201) <= b and not a;
    layer2_outputs(9202) <= 1'b0;
    layer2_outputs(9203) <= b;
    layer2_outputs(9204) <= not b;
    layer2_outputs(9205) <= b;
    layer2_outputs(9206) <= not (a and b);
    layer2_outputs(9207) <= not (a and b);
    layer2_outputs(9208) <= b;
    layer2_outputs(9209) <= not (a xor b);
    layer2_outputs(9210) <= not b;
    layer2_outputs(9211) <= not b or a;
    layer2_outputs(9212) <= a or b;
    layer2_outputs(9213) <= not b;
    layer2_outputs(9214) <= not (a and b);
    layer2_outputs(9215) <= not (a and b);
    layer2_outputs(9216) <= not (a xor b);
    layer2_outputs(9217) <= a xor b;
    layer2_outputs(9218) <= b;
    layer2_outputs(9219) <= b;
    layer2_outputs(9220) <= b and not a;
    layer2_outputs(9221) <= b;
    layer2_outputs(9222) <= not (a or b);
    layer2_outputs(9223) <= not (a and b);
    layer2_outputs(9224) <= not (a or b);
    layer2_outputs(9225) <= a;
    layer2_outputs(9226) <= not (a xor b);
    layer2_outputs(9227) <= a xor b;
    layer2_outputs(9228) <= a and b;
    layer2_outputs(9229) <= b and not a;
    layer2_outputs(9230) <= a;
    layer2_outputs(9231) <= not (a xor b);
    layer2_outputs(9232) <= not b;
    layer2_outputs(9233) <= a or b;
    layer2_outputs(9234) <= not a or b;
    layer2_outputs(9235) <= b;
    layer2_outputs(9236) <= not (a and b);
    layer2_outputs(9237) <= not (a xor b);
    layer2_outputs(9238) <= a or b;
    layer2_outputs(9239) <= a and b;
    layer2_outputs(9240) <= b and not a;
    layer2_outputs(9241) <= b and not a;
    layer2_outputs(9242) <= not b or a;
    layer2_outputs(9243) <= a;
    layer2_outputs(9244) <= not (a and b);
    layer2_outputs(9245) <= not (a or b);
    layer2_outputs(9246) <= not (a xor b);
    layer2_outputs(9247) <= not (a or b);
    layer2_outputs(9248) <= b;
    layer2_outputs(9249) <= not a;
    layer2_outputs(9250) <= not b;
    layer2_outputs(9251) <= not (a and b);
    layer2_outputs(9252) <= a;
    layer2_outputs(9253) <= not (a xor b);
    layer2_outputs(9254) <= not (a xor b);
    layer2_outputs(9255) <= not b or a;
    layer2_outputs(9256) <= not (a or b);
    layer2_outputs(9257) <= b;
    layer2_outputs(9258) <= not b;
    layer2_outputs(9259) <= a and b;
    layer2_outputs(9260) <= not b;
    layer2_outputs(9261) <= a;
    layer2_outputs(9262) <= a and not b;
    layer2_outputs(9263) <= not a;
    layer2_outputs(9264) <= not a;
    layer2_outputs(9265) <= a xor b;
    layer2_outputs(9266) <= a;
    layer2_outputs(9267) <= not a;
    layer2_outputs(9268) <= not (a or b);
    layer2_outputs(9269) <= 1'b1;
    layer2_outputs(9270) <= b;
    layer2_outputs(9271) <= a;
    layer2_outputs(9272) <= not (a or b);
    layer2_outputs(9273) <= a and not b;
    layer2_outputs(9274) <= b;
    layer2_outputs(9275) <= not (a and b);
    layer2_outputs(9276) <= 1'b0;
    layer2_outputs(9277) <= not a or b;
    layer2_outputs(9278) <= a or b;
    layer2_outputs(9279) <= a or b;
    layer2_outputs(9280) <= 1'b1;
    layer2_outputs(9281) <= b and not a;
    layer2_outputs(9282) <= a or b;
    layer2_outputs(9283) <= not a or b;
    layer2_outputs(9284) <= a and b;
    layer2_outputs(9285) <= a;
    layer2_outputs(9286) <= not a;
    layer2_outputs(9287) <= a or b;
    layer2_outputs(9288) <= not b or a;
    layer2_outputs(9289) <= not a or b;
    layer2_outputs(9290) <= b;
    layer2_outputs(9291) <= b;
    layer2_outputs(9292) <= a xor b;
    layer2_outputs(9293) <= not a or b;
    layer2_outputs(9294) <= a or b;
    layer2_outputs(9295) <= not (a or b);
    layer2_outputs(9296) <= a or b;
    layer2_outputs(9297) <= a and not b;
    layer2_outputs(9298) <= not b or a;
    layer2_outputs(9299) <= a or b;
    layer2_outputs(9300) <= not b;
    layer2_outputs(9301) <= b and not a;
    layer2_outputs(9302) <= not (a and b);
    layer2_outputs(9303) <= a or b;
    layer2_outputs(9304) <= a and b;
    layer2_outputs(9305) <= a xor b;
    layer2_outputs(9306) <= b;
    layer2_outputs(9307) <= not a;
    layer2_outputs(9308) <= b;
    layer2_outputs(9309) <= not a;
    layer2_outputs(9310) <= a or b;
    layer2_outputs(9311) <= a and b;
    layer2_outputs(9312) <= a or b;
    layer2_outputs(9313) <= not (a and b);
    layer2_outputs(9314) <= b;
    layer2_outputs(9315) <= not b;
    layer2_outputs(9316) <= a and b;
    layer2_outputs(9317) <= not (a xor b);
    layer2_outputs(9318) <= a;
    layer2_outputs(9319) <= not a;
    layer2_outputs(9320) <= not a or b;
    layer2_outputs(9321) <= not b;
    layer2_outputs(9322) <= a and not b;
    layer2_outputs(9323) <= a;
    layer2_outputs(9324) <= a;
    layer2_outputs(9325) <= not a or b;
    layer2_outputs(9326) <= a;
    layer2_outputs(9327) <= not (a or b);
    layer2_outputs(9328) <= not b or a;
    layer2_outputs(9329) <= b and not a;
    layer2_outputs(9330) <= not (a xor b);
    layer2_outputs(9331) <= not b or a;
    layer2_outputs(9332) <= b;
    layer2_outputs(9333) <= 1'b0;
    layer2_outputs(9334) <= b;
    layer2_outputs(9335) <= a xor b;
    layer2_outputs(9336) <= a;
    layer2_outputs(9337) <= a;
    layer2_outputs(9338) <= b;
    layer2_outputs(9339) <= not b or a;
    layer2_outputs(9340) <= not b;
    layer2_outputs(9341) <= b and not a;
    layer2_outputs(9342) <= not b;
    layer2_outputs(9343) <= not b;
    layer2_outputs(9344) <= b;
    layer2_outputs(9345) <= 1'b0;
    layer2_outputs(9346) <= a and b;
    layer2_outputs(9347) <= b;
    layer2_outputs(9348) <= a and not b;
    layer2_outputs(9349) <= b and not a;
    layer2_outputs(9350) <= a and b;
    layer2_outputs(9351) <= not (a xor b);
    layer2_outputs(9352) <= not b;
    layer2_outputs(9353) <= a;
    layer2_outputs(9354) <= not (a xor b);
    layer2_outputs(9355) <= not (a or b);
    layer2_outputs(9356) <= a;
    layer2_outputs(9357) <= not a or b;
    layer2_outputs(9358) <= a;
    layer2_outputs(9359) <= b;
    layer2_outputs(9360) <= b;
    layer2_outputs(9361) <= not (a and b);
    layer2_outputs(9362) <= b;
    layer2_outputs(9363) <= not (a or b);
    layer2_outputs(9364) <= not (a and b);
    layer2_outputs(9365) <= not (a xor b);
    layer2_outputs(9366) <= a;
    layer2_outputs(9367) <= not b;
    layer2_outputs(9368) <= a xor b;
    layer2_outputs(9369) <= not b;
    layer2_outputs(9370) <= not a or b;
    layer2_outputs(9371) <= not b;
    layer2_outputs(9372) <= not (a or b);
    layer2_outputs(9373) <= not b;
    layer2_outputs(9374) <= not a;
    layer2_outputs(9375) <= not b;
    layer2_outputs(9376) <= not a;
    layer2_outputs(9377) <= not a;
    layer2_outputs(9378) <= not (a and b);
    layer2_outputs(9379) <= a and b;
    layer2_outputs(9380) <= a xor b;
    layer2_outputs(9381) <= 1'b1;
    layer2_outputs(9382) <= a;
    layer2_outputs(9383) <= b and not a;
    layer2_outputs(9384) <= a xor b;
    layer2_outputs(9385) <= a or b;
    layer2_outputs(9386) <= a or b;
    layer2_outputs(9387) <= 1'b1;
    layer2_outputs(9388) <= not (a and b);
    layer2_outputs(9389) <= b;
    layer2_outputs(9390) <= not b;
    layer2_outputs(9391) <= a xor b;
    layer2_outputs(9392) <= b;
    layer2_outputs(9393) <= not a;
    layer2_outputs(9394) <= not a;
    layer2_outputs(9395) <= not b or a;
    layer2_outputs(9396) <= not (a and b);
    layer2_outputs(9397) <= a;
    layer2_outputs(9398) <= not (a xor b);
    layer2_outputs(9399) <= not b;
    layer2_outputs(9400) <= not b;
    layer2_outputs(9401) <= not b;
    layer2_outputs(9402) <= not (a or b);
    layer2_outputs(9403) <= 1'b1;
    layer2_outputs(9404) <= not (a and b);
    layer2_outputs(9405) <= b;
    layer2_outputs(9406) <= a;
    layer2_outputs(9407) <= not b;
    layer2_outputs(9408) <= a xor b;
    layer2_outputs(9409) <= not (a or b);
    layer2_outputs(9410) <= a;
    layer2_outputs(9411) <= not a;
    layer2_outputs(9412) <= 1'b0;
    layer2_outputs(9413) <= b and not a;
    layer2_outputs(9414) <= a or b;
    layer2_outputs(9415) <= not (a and b);
    layer2_outputs(9416) <= b;
    layer2_outputs(9417) <= a;
    layer2_outputs(9418) <= 1'b0;
    layer2_outputs(9419) <= a and not b;
    layer2_outputs(9420) <= not a or b;
    layer2_outputs(9421) <= 1'b1;
    layer2_outputs(9422) <= a;
    layer2_outputs(9423) <= a and not b;
    layer2_outputs(9424) <= a xor b;
    layer2_outputs(9425) <= b and not a;
    layer2_outputs(9426) <= not b or a;
    layer2_outputs(9427) <= b and not a;
    layer2_outputs(9428) <= 1'b0;
    layer2_outputs(9429) <= 1'b0;
    layer2_outputs(9430) <= 1'b1;
    layer2_outputs(9431) <= not a or b;
    layer2_outputs(9432) <= a;
    layer2_outputs(9433) <= b;
    layer2_outputs(9434) <= not b;
    layer2_outputs(9435) <= not a;
    layer2_outputs(9436) <= not b;
    layer2_outputs(9437) <= a xor b;
    layer2_outputs(9438) <= not b or a;
    layer2_outputs(9439) <= 1'b0;
    layer2_outputs(9440) <= b;
    layer2_outputs(9441) <= a and b;
    layer2_outputs(9442) <= not b or a;
    layer2_outputs(9443) <= a;
    layer2_outputs(9444) <= not (a xor b);
    layer2_outputs(9445) <= not a or b;
    layer2_outputs(9446) <= b;
    layer2_outputs(9447) <= a and b;
    layer2_outputs(9448) <= a and b;
    layer2_outputs(9449) <= a or b;
    layer2_outputs(9450) <= not (a and b);
    layer2_outputs(9451) <= a xor b;
    layer2_outputs(9452) <= not (a and b);
    layer2_outputs(9453) <= b;
    layer2_outputs(9454) <= not a;
    layer2_outputs(9455) <= 1'b1;
    layer2_outputs(9456) <= a;
    layer2_outputs(9457) <= not a;
    layer2_outputs(9458) <= not (a xor b);
    layer2_outputs(9459) <= not (a or b);
    layer2_outputs(9460) <= not (a xor b);
    layer2_outputs(9461) <= a xor b;
    layer2_outputs(9462) <= a;
    layer2_outputs(9463) <= not a;
    layer2_outputs(9464) <= not a;
    layer2_outputs(9465) <= a and b;
    layer2_outputs(9466) <= not (a xor b);
    layer2_outputs(9467) <= not b or a;
    layer2_outputs(9468) <= a or b;
    layer2_outputs(9469) <= a;
    layer2_outputs(9470) <= not (a xor b);
    layer2_outputs(9471) <= not (a xor b);
    layer2_outputs(9472) <= b;
    layer2_outputs(9473) <= b and not a;
    layer2_outputs(9474) <= not (a xor b);
    layer2_outputs(9475) <= not a;
    layer2_outputs(9476) <= a and not b;
    layer2_outputs(9477) <= not a;
    layer2_outputs(9478) <= b;
    layer2_outputs(9479) <= not b;
    layer2_outputs(9480) <= 1'b1;
    layer2_outputs(9481) <= a and not b;
    layer2_outputs(9482) <= b and not a;
    layer2_outputs(9483) <= b;
    layer2_outputs(9484) <= a and not b;
    layer2_outputs(9485) <= not b;
    layer2_outputs(9486) <= not (a or b);
    layer2_outputs(9487) <= not a;
    layer2_outputs(9488) <= not (a or b);
    layer2_outputs(9489) <= a and b;
    layer2_outputs(9490) <= not a;
    layer2_outputs(9491) <= b;
    layer2_outputs(9492) <= not b;
    layer2_outputs(9493) <= not a or b;
    layer2_outputs(9494) <= not b;
    layer2_outputs(9495) <= a and not b;
    layer2_outputs(9496) <= not a;
    layer2_outputs(9497) <= not (a and b);
    layer2_outputs(9498) <= a or b;
    layer2_outputs(9499) <= not b;
    layer2_outputs(9500) <= not a;
    layer2_outputs(9501) <= a;
    layer2_outputs(9502) <= b and not a;
    layer2_outputs(9503) <= not a or b;
    layer2_outputs(9504) <= not (a or b);
    layer2_outputs(9505) <= a and not b;
    layer2_outputs(9506) <= not (a xor b);
    layer2_outputs(9507) <= not a or b;
    layer2_outputs(9508) <= not a;
    layer2_outputs(9509) <= not a or b;
    layer2_outputs(9510) <= not (a or b);
    layer2_outputs(9511) <= a and not b;
    layer2_outputs(9512) <= not b or a;
    layer2_outputs(9513) <= not a or b;
    layer2_outputs(9514) <= not b;
    layer2_outputs(9515) <= a and b;
    layer2_outputs(9516) <= not (a xor b);
    layer2_outputs(9517) <= not b;
    layer2_outputs(9518) <= b;
    layer2_outputs(9519) <= not a or b;
    layer2_outputs(9520) <= a;
    layer2_outputs(9521) <= not (a xor b);
    layer2_outputs(9522) <= b and not a;
    layer2_outputs(9523) <= not (a or b);
    layer2_outputs(9524) <= not a or b;
    layer2_outputs(9525) <= a xor b;
    layer2_outputs(9526) <= a xor b;
    layer2_outputs(9527) <= not b;
    layer2_outputs(9528) <= a;
    layer2_outputs(9529) <= not a;
    layer2_outputs(9530) <= not (a or b);
    layer2_outputs(9531) <= a xor b;
    layer2_outputs(9532) <= a and not b;
    layer2_outputs(9533) <= a;
    layer2_outputs(9534) <= a or b;
    layer2_outputs(9535) <= not (a xor b);
    layer2_outputs(9536) <= not b;
    layer2_outputs(9537) <= a;
    layer2_outputs(9538) <= a;
    layer2_outputs(9539) <= not (a xor b);
    layer2_outputs(9540) <= not b;
    layer2_outputs(9541) <= a and not b;
    layer2_outputs(9542) <= a or b;
    layer2_outputs(9543) <= b;
    layer2_outputs(9544) <= not (a or b);
    layer2_outputs(9545) <= not a;
    layer2_outputs(9546) <= not (a and b);
    layer2_outputs(9547) <= not a or b;
    layer2_outputs(9548) <= 1'b0;
    layer2_outputs(9549) <= a and b;
    layer2_outputs(9550) <= not a;
    layer2_outputs(9551) <= a and not b;
    layer2_outputs(9552) <= a;
    layer2_outputs(9553) <= not (a and b);
    layer2_outputs(9554) <= b and not a;
    layer2_outputs(9555) <= not b;
    layer2_outputs(9556) <= a or b;
    layer2_outputs(9557) <= not a;
    layer2_outputs(9558) <= a and b;
    layer2_outputs(9559) <= b and not a;
    layer2_outputs(9560) <= not a or b;
    layer2_outputs(9561) <= not b or a;
    layer2_outputs(9562) <= a or b;
    layer2_outputs(9563) <= not b or a;
    layer2_outputs(9564) <= not b;
    layer2_outputs(9565) <= not (a and b);
    layer2_outputs(9566) <= not a or b;
    layer2_outputs(9567) <= not a or b;
    layer2_outputs(9568) <= not b;
    layer2_outputs(9569) <= a or b;
    layer2_outputs(9570) <= b;
    layer2_outputs(9571) <= b;
    layer2_outputs(9572) <= a or b;
    layer2_outputs(9573) <= a;
    layer2_outputs(9574) <= a or b;
    layer2_outputs(9575) <= b;
    layer2_outputs(9576) <= not (a xor b);
    layer2_outputs(9577) <= not (a or b);
    layer2_outputs(9578) <= a and b;
    layer2_outputs(9579) <= not (a xor b);
    layer2_outputs(9580) <= not b;
    layer2_outputs(9581) <= a;
    layer2_outputs(9582) <= not b;
    layer2_outputs(9583) <= b and not a;
    layer2_outputs(9584) <= not a;
    layer2_outputs(9585) <= not b or a;
    layer2_outputs(9586) <= a and not b;
    layer2_outputs(9587) <= a and not b;
    layer2_outputs(9588) <= a;
    layer2_outputs(9589) <= not (a and b);
    layer2_outputs(9590) <= not b or a;
    layer2_outputs(9591) <= not a;
    layer2_outputs(9592) <= not b;
    layer2_outputs(9593) <= not (a or b);
    layer2_outputs(9594) <= a and not b;
    layer2_outputs(9595) <= a and not b;
    layer2_outputs(9596) <= a and b;
    layer2_outputs(9597) <= a or b;
    layer2_outputs(9598) <= a and b;
    layer2_outputs(9599) <= a;
    layer2_outputs(9600) <= not b;
    layer2_outputs(9601) <= a and not b;
    layer2_outputs(9602) <= b;
    layer2_outputs(9603) <= not (a xor b);
    layer2_outputs(9604) <= a xor b;
    layer2_outputs(9605) <= b;
    layer2_outputs(9606) <= not (a and b);
    layer2_outputs(9607) <= a xor b;
    layer2_outputs(9608) <= not b or a;
    layer2_outputs(9609) <= 1'b1;
    layer2_outputs(9610) <= not (a xor b);
    layer2_outputs(9611) <= a or b;
    layer2_outputs(9612) <= b and not a;
    layer2_outputs(9613) <= 1'b0;
    layer2_outputs(9614) <= b;
    layer2_outputs(9615) <= not b or a;
    layer2_outputs(9616) <= not b or a;
    layer2_outputs(9617) <= a;
    layer2_outputs(9618) <= not b or a;
    layer2_outputs(9619) <= a and not b;
    layer2_outputs(9620) <= a xor b;
    layer2_outputs(9621) <= a and not b;
    layer2_outputs(9622) <= not a;
    layer2_outputs(9623) <= a xor b;
    layer2_outputs(9624) <= not (a xor b);
    layer2_outputs(9625) <= not b or a;
    layer2_outputs(9626) <= not a;
    layer2_outputs(9627) <= not a or b;
    layer2_outputs(9628) <= a;
    layer2_outputs(9629) <= a or b;
    layer2_outputs(9630) <= not b;
    layer2_outputs(9631) <= not a;
    layer2_outputs(9632) <= not (a and b);
    layer2_outputs(9633) <= a or b;
    layer2_outputs(9634) <= b and not a;
    layer2_outputs(9635) <= not (a or b);
    layer2_outputs(9636) <= b;
    layer2_outputs(9637) <= not b;
    layer2_outputs(9638) <= b;
    layer2_outputs(9639) <= not b;
    layer2_outputs(9640) <= b and not a;
    layer2_outputs(9641) <= not (a and b);
    layer2_outputs(9642) <= a;
    layer2_outputs(9643) <= not a;
    layer2_outputs(9644) <= not a or b;
    layer2_outputs(9645) <= b;
    layer2_outputs(9646) <= not a;
    layer2_outputs(9647) <= a;
    layer2_outputs(9648) <= b and not a;
    layer2_outputs(9649) <= b and not a;
    layer2_outputs(9650) <= not b or a;
    layer2_outputs(9651) <= a xor b;
    layer2_outputs(9652) <= not b;
    layer2_outputs(9653) <= b;
    layer2_outputs(9654) <= not a;
    layer2_outputs(9655) <= not (a or b);
    layer2_outputs(9656) <= a and b;
    layer2_outputs(9657) <= not b;
    layer2_outputs(9658) <= not a;
    layer2_outputs(9659) <= a and b;
    layer2_outputs(9660) <= not (a and b);
    layer2_outputs(9661) <= a and b;
    layer2_outputs(9662) <= a xor b;
    layer2_outputs(9663) <= a and not b;
    layer2_outputs(9664) <= a and not b;
    layer2_outputs(9665) <= b;
    layer2_outputs(9666) <= not (a or b);
    layer2_outputs(9667) <= a xor b;
    layer2_outputs(9668) <= b;
    layer2_outputs(9669) <= not (a and b);
    layer2_outputs(9670) <= not (a xor b);
    layer2_outputs(9671) <= not b;
    layer2_outputs(9672) <= not b;
    layer2_outputs(9673) <= 1'b1;
    layer2_outputs(9674) <= b and not a;
    layer2_outputs(9675) <= b;
    layer2_outputs(9676) <= not (a and b);
    layer2_outputs(9677) <= not b or a;
    layer2_outputs(9678) <= not (a xor b);
    layer2_outputs(9679) <= b and not a;
    layer2_outputs(9680) <= a xor b;
    layer2_outputs(9681) <= a or b;
    layer2_outputs(9682) <= b;
    layer2_outputs(9683) <= not a;
    layer2_outputs(9684) <= a xor b;
    layer2_outputs(9685) <= b and not a;
    layer2_outputs(9686) <= not (a and b);
    layer2_outputs(9687) <= a or b;
    layer2_outputs(9688) <= b and not a;
    layer2_outputs(9689) <= b;
    layer2_outputs(9690) <= not b or a;
    layer2_outputs(9691) <= not (a and b);
    layer2_outputs(9692) <= not (a or b);
    layer2_outputs(9693) <= b;
    layer2_outputs(9694) <= b and not a;
    layer2_outputs(9695) <= b;
    layer2_outputs(9696) <= not b or a;
    layer2_outputs(9697) <= a and b;
    layer2_outputs(9698) <= not (a xor b);
    layer2_outputs(9699) <= not (a and b);
    layer2_outputs(9700) <= a and b;
    layer2_outputs(9701) <= a xor b;
    layer2_outputs(9702) <= not a;
    layer2_outputs(9703) <= not a;
    layer2_outputs(9704) <= a and not b;
    layer2_outputs(9705) <= not a or b;
    layer2_outputs(9706) <= not (a and b);
    layer2_outputs(9707) <= not a or b;
    layer2_outputs(9708) <= a and not b;
    layer2_outputs(9709) <= not b;
    layer2_outputs(9710) <= not b;
    layer2_outputs(9711) <= not (a or b);
    layer2_outputs(9712) <= not a or b;
    layer2_outputs(9713) <= not b;
    layer2_outputs(9714) <= not a or b;
    layer2_outputs(9715) <= b;
    layer2_outputs(9716) <= not (a xor b);
    layer2_outputs(9717) <= a and not b;
    layer2_outputs(9718) <= a and b;
    layer2_outputs(9719) <= b;
    layer2_outputs(9720) <= b;
    layer2_outputs(9721) <= not b or a;
    layer2_outputs(9722) <= not (a xor b);
    layer2_outputs(9723) <= not (a or b);
    layer2_outputs(9724) <= not a;
    layer2_outputs(9725) <= not (a xor b);
    layer2_outputs(9726) <= not b;
    layer2_outputs(9727) <= not b or a;
    layer2_outputs(9728) <= b and not a;
    layer2_outputs(9729) <= not b;
    layer2_outputs(9730) <= 1'b0;
    layer2_outputs(9731) <= b;
    layer2_outputs(9732) <= b;
    layer2_outputs(9733) <= a and b;
    layer2_outputs(9734) <= not a;
    layer2_outputs(9735) <= a or b;
    layer2_outputs(9736) <= not a or b;
    layer2_outputs(9737) <= not a;
    layer2_outputs(9738) <= not a;
    layer2_outputs(9739) <= not b or a;
    layer2_outputs(9740) <= a and not b;
    layer2_outputs(9741) <= a;
    layer2_outputs(9742) <= b;
    layer2_outputs(9743) <= not (a xor b);
    layer2_outputs(9744) <= not a;
    layer2_outputs(9745) <= a;
    layer2_outputs(9746) <= not a;
    layer2_outputs(9747) <= not a or b;
    layer2_outputs(9748) <= not b;
    layer2_outputs(9749) <= b and not a;
    layer2_outputs(9750) <= not b or a;
    layer2_outputs(9751) <= a xor b;
    layer2_outputs(9752) <= not a;
    layer2_outputs(9753) <= not (a xor b);
    layer2_outputs(9754) <= a;
    layer2_outputs(9755) <= a and not b;
    layer2_outputs(9756) <= a and not b;
    layer2_outputs(9757) <= a xor b;
    layer2_outputs(9758) <= a or b;
    layer2_outputs(9759) <= not (a or b);
    layer2_outputs(9760) <= not b;
    layer2_outputs(9761) <= a xor b;
    layer2_outputs(9762) <= a or b;
    layer2_outputs(9763) <= not a or b;
    layer2_outputs(9764) <= a xor b;
    layer2_outputs(9765) <= not b;
    layer2_outputs(9766) <= not (a and b);
    layer2_outputs(9767) <= not a;
    layer2_outputs(9768) <= not b;
    layer2_outputs(9769) <= b;
    layer2_outputs(9770) <= not (a and b);
    layer2_outputs(9771) <= not b or a;
    layer2_outputs(9772) <= not (a or b);
    layer2_outputs(9773) <= not b;
    layer2_outputs(9774) <= b;
    layer2_outputs(9775) <= a or b;
    layer2_outputs(9776) <= not (a and b);
    layer2_outputs(9777) <= a;
    layer2_outputs(9778) <= not b or a;
    layer2_outputs(9779) <= a and not b;
    layer2_outputs(9780) <= not (a or b);
    layer2_outputs(9781) <= not b;
    layer2_outputs(9782) <= not (a or b);
    layer2_outputs(9783) <= not b or a;
    layer2_outputs(9784) <= 1'b0;
    layer2_outputs(9785) <= not (a or b);
    layer2_outputs(9786) <= not a;
    layer2_outputs(9787) <= not (a or b);
    layer2_outputs(9788) <= 1'b0;
    layer2_outputs(9789) <= 1'b1;
    layer2_outputs(9790) <= a and b;
    layer2_outputs(9791) <= a and b;
    layer2_outputs(9792) <= a and not b;
    layer2_outputs(9793) <= not b or a;
    layer2_outputs(9794) <= b;
    layer2_outputs(9795) <= not (a and b);
    layer2_outputs(9796) <= a;
    layer2_outputs(9797) <= not a or b;
    layer2_outputs(9798) <= a and not b;
    layer2_outputs(9799) <= b and not a;
    layer2_outputs(9800) <= a xor b;
    layer2_outputs(9801) <= not b;
    layer2_outputs(9802) <= b;
    layer2_outputs(9803) <= not (a xor b);
    layer2_outputs(9804) <= not (a or b);
    layer2_outputs(9805) <= not (a or b);
    layer2_outputs(9806) <= b and not a;
    layer2_outputs(9807) <= a;
    layer2_outputs(9808) <= not a or b;
    layer2_outputs(9809) <= a;
    layer2_outputs(9810) <= b;
    layer2_outputs(9811) <= a;
    layer2_outputs(9812) <= b;
    layer2_outputs(9813) <= not a;
    layer2_outputs(9814) <= not b;
    layer2_outputs(9815) <= a and not b;
    layer2_outputs(9816) <= not a or b;
    layer2_outputs(9817) <= 1'b1;
    layer2_outputs(9818) <= b;
    layer2_outputs(9819) <= 1'b0;
    layer2_outputs(9820) <= a and b;
    layer2_outputs(9821) <= 1'b0;
    layer2_outputs(9822) <= a or b;
    layer2_outputs(9823) <= not (a and b);
    layer2_outputs(9824) <= not b or a;
    layer2_outputs(9825) <= not b;
    layer2_outputs(9826) <= a xor b;
    layer2_outputs(9827) <= a or b;
    layer2_outputs(9828) <= not a;
    layer2_outputs(9829) <= not (a or b);
    layer2_outputs(9830) <= not a;
    layer2_outputs(9831) <= a or b;
    layer2_outputs(9832) <= b;
    layer2_outputs(9833) <= not (a or b);
    layer2_outputs(9834) <= not (a xor b);
    layer2_outputs(9835) <= not a or b;
    layer2_outputs(9836) <= not (a or b);
    layer2_outputs(9837) <= b;
    layer2_outputs(9838) <= b and not a;
    layer2_outputs(9839) <= a xor b;
    layer2_outputs(9840) <= not b;
    layer2_outputs(9841) <= a;
    layer2_outputs(9842) <= not (a and b);
    layer2_outputs(9843) <= a xor b;
    layer2_outputs(9844) <= not b or a;
    layer2_outputs(9845) <= not (a and b);
    layer2_outputs(9846) <= not (a xor b);
    layer2_outputs(9847) <= b;
    layer2_outputs(9848) <= a and b;
    layer2_outputs(9849) <= not a;
    layer2_outputs(9850) <= a and not b;
    layer2_outputs(9851) <= a and not b;
    layer2_outputs(9852) <= not a;
    layer2_outputs(9853) <= b;
    layer2_outputs(9854) <= not (a or b);
    layer2_outputs(9855) <= 1'b1;
    layer2_outputs(9856) <= not b or a;
    layer2_outputs(9857) <= a xor b;
    layer2_outputs(9858) <= not a;
    layer2_outputs(9859) <= a;
    layer2_outputs(9860) <= b;
    layer2_outputs(9861) <= b;
    layer2_outputs(9862) <= a and b;
    layer2_outputs(9863) <= not a;
    layer2_outputs(9864) <= a and not b;
    layer2_outputs(9865) <= not (a or b);
    layer2_outputs(9866) <= 1'b1;
    layer2_outputs(9867) <= b and not a;
    layer2_outputs(9868) <= 1'b1;
    layer2_outputs(9869) <= a or b;
    layer2_outputs(9870) <= b;
    layer2_outputs(9871) <= b and not a;
    layer2_outputs(9872) <= a and not b;
    layer2_outputs(9873) <= not a;
    layer2_outputs(9874) <= a;
    layer2_outputs(9875) <= not (a and b);
    layer2_outputs(9876) <= 1'b1;
    layer2_outputs(9877) <= b;
    layer2_outputs(9878) <= not b;
    layer2_outputs(9879) <= not b;
    layer2_outputs(9880) <= a and not b;
    layer2_outputs(9881) <= a;
    layer2_outputs(9882) <= not a or b;
    layer2_outputs(9883) <= a and not b;
    layer2_outputs(9884) <= not (a xor b);
    layer2_outputs(9885) <= not a;
    layer2_outputs(9886) <= not a or b;
    layer2_outputs(9887) <= not a;
    layer2_outputs(9888) <= b;
    layer2_outputs(9889) <= not (a and b);
    layer2_outputs(9890) <= not a or b;
    layer2_outputs(9891) <= a;
    layer2_outputs(9892) <= not a;
    layer2_outputs(9893) <= 1'b1;
    layer2_outputs(9894) <= not a;
    layer2_outputs(9895) <= not b or a;
    layer2_outputs(9896) <= not b;
    layer2_outputs(9897) <= a;
    layer2_outputs(9898) <= not (a or b);
    layer2_outputs(9899) <= a and b;
    layer2_outputs(9900) <= a or b;
    layer2_outputs(9901) <= a and not b;
    layer2_outputs(9902) <= 1'b1;
    layer2_outputs(9903) <= not a;
    layer2_outputs(9904) <= a or b;
    layer2_outputs(9905) <= a or b;
    layer2_outputs(9906) <= b and not a;
    layer2_outputs(9907) <= b and not a;
    layer2_outputs(9908) <= a or b;
    layer2_outputs(9909) <= a xor b;
    layer2_outputs(9910) <= not b;
    layer2_outputs(9911) <= b;
    layer2_outputs(9912) <= not b;
    layer2_outputs(9913) <= not b;
    layer2_outputs(9914) <= a;
    layer2_outputs(9915) <= b;
    layer2_outputs(9916) <= a;
    layer2_outputs(9917) <= a;
    layer2_outputs(9918) <= a;
    layer2_outputs(9919) <= not a;
    layer2_outputs(9920) <= not b or a;
    layer2_outputs(9921) <= 1'b0;
    layer2_outputs(9922) <= not b or a;
    layer2_outputs(9923) <= b;
    layer2_outputs(9924) <= b;
    layer2_outputs(9925) <= b;
    layer2_outputs(9926) <= b;
    layer2_outputs(9927) <= a;
    layer2_outputs(9928) <= not (a xor b);
    layer2_outputs(9929) <= a xor b;
    layer2_outputs(9930) <= not a or b;
    layer2_outputs(9931) <= not b;
    layer2_outputs(9932) <= not b;
    layer2_outputs(9933) <= not (a or b);
    layer2_outputs(9934) <= not (a and b);
    layer2_outputs(9935) <= a and not b;
    layer2_outputs(9936) <= not a or b;
    layer2_outputs(9937) <= not b;
    layer2_outputs(9938) <= not b;
    layer2_outputs(9939) <= not a;
    layer2_outputs(9940) <= not a;
    layer2_outputs(9941) <= a and not b;
    layer2_outputs(9942) <= not (a xor b);
    layer2_outputs(9943) <= 1'b1;
    layer2_outputs(9944) <= not (a or b);
    layer2_outputs(9945) <= b;
    layer2_outputs(9946) <= a or b;
    layer2_outputs(9947) <= a or b;
    layer2_outputs(9948) <= b and not a;
    layer2_outputs(9949) <= b;
    layer2_outputs(9950) <= a;
    layer2_outputs(9951) <= a and b;
    layer2_outputs(9952) <= 1'b1;
    layer2_outputs(9953) <= not (a xor b);
    layer2_outputs(9954) <= a and not b;
    layer2_outputs(9955) <= not a;
    layer2_outputs(9956) <= 1'b0;
    layer2_outputs(9957) <= b;
    layer2_outputs(9958) <= not b;
    layer2_outputs(9959) <= b;
    layer2_outputs(9960) <= not b or a;
    layer2_outputs(9961) <= b;
    layer2_outputs(9962) <= b;
    layer2_outputs(9963) <= a;
    layer2_outputs(9964) <= 1'b1;
    layer2_outputs(9965) <= a and b;
    layer2_outputs(9966) <= a;
    layer2_outputs(9967) <= a and b;
    layer2_outputs(9968) <= a;
    layer2_outputs(9969) <= b;
    layer2_outputs(9970) <= b;
    layer2_outputs(9971) <= not b;
    layer2_outputs(9972) <= a and not b;
    layer2_outputs(9973) <= a;
    layer2_outputs(9974) <= not (a and b);
    layer2_outputs(9975) <= a and b;
    layer2_outputs(9976) <= a or b;
    layer2_outputs(9977) <= not (a xor b);
    layer2_outputs(9978) <= not (a and b);
    layer2_outputs(9979) <= not (a xor b);
    layer2_outputs(9980) <= a xor b;
    layer2_outputs(9981) <= not b or a;
    layer2_outputs(9982) <= not a;
    layer2_outputs(9983) <= a and b;
    layer2_outputs(9984) <= not (a xor b);
    layer2_outputs(9985) <= a;
    layer2_outputs(9986) <= a or b;
    layer2_outputs(9987) <= not (a xor b);
    layer2_outputs(9988) <= not b or a;
    layer2_outputs(9989) <= 1'b0;
    layer2_outputs(9990) <= a;
    layer2_outputs(9991) <= a;
    layer2_outputs(9992) <= b;
    layer2_outputs(9993) <= not (a and b);
    layer2_outputs(9994) <= not a;
    layer2_outputs(9995) <= not b or a;
    layer2_outputs(9996) <= not a or b;
    layer2_outputs(9997) <= b and not a;
    layer2_outputs(9998) <= b;
    layer2_outputs(9999) <= not (a and b);
    layer2_outputs(10000) <= a or b;
    layer2_outputs(10001) <= not (a and b);
    layer2_outputs(10002) <= a and not b;
    layer2_outputs(10003) <= b;
    layer2_outputs(10004) <= a;
    layer2_outputs(10005) <= b;
    layer2_outputs(10006) <= a or b;
    layer2_outputs(10007) <= not (a or b);
    layer2_outputs(10008) <= a;
    layer2_outputs(10009) <= a xor b;
    layer2_outputs(10010) <= a and not b;
    layer2_outputs(10011) <= 1'b0;
    layer2_outputs(10012) <= b;
    layer2_outputs(10013) <= b and not a;
    layer2_outputs(10014) <= b;
    layer2_outputs(10015) <= not (a xor b);
    layer2_outputs(10016) <= not a or b;
    layer2_outputs(10017) <= b and not a;
    layer2_outputs(10018) <= not b;
    layer2_outputs(10019) <= 1'b1;
    layer2_outputs(10020) <= not a;
    layer2_outputs(10021) <= a and b;
    layer2_outputs(10022) <= not a;
    layer2_outputs(10023) <= a or b;
    layer2_outputs(10024) <= a and not b;
    layer2_outputs(10025) <= a or b;
    layer2_outputs(10026) <= a;
    layer2_outputs(10027) <= a;
    layer2_outputs(10028) <= a and not b;
    layer2_outputs(10029) <= a xor b;
    layer2_outputs(10030) <= not (a or b);
    layer2_outputs(10031) <= a xor b;
    layer2_outputs(10032) <= a xor b;
    layer2_outputs(10033) <= not a;
    layer2_outputs(10034) <= a xor b;
    layer2_outputs(10035) <= b;
    layer2_outputs(10036) <= not (a or b);
    layer2_outputs(10037) <= not a;
    layer2_outputs(10038) <= b;
    layer2_outputs(10039) <= a xor b;
    layer2_outputs(10040) <= not (a and b);
    layer2_outputs(10041) <= 1'b0;
    layer2_outputs(10042) <= b and not a;
    layer2_outputs(10043) <= b and not a;
    layer2_outputs(10044) <= a or b;
    layer2_outputs(10045) <= not a or b;
    layer2_outputs(10046) <= not (a or b);
    layer2_outputs(10047) <= a and b;
    layer2_outputs(10048) <= not (a or b);
    layer2_outputs(10049) <= not a or b;
    layer2_outputs(10050) <= b;
    layer2_outputs(10051) <= a and not b;
    layer2_outputs(10052) <= not (a and b);
    layer2_outputs(10053) <= a;
    layer2_outputs(10054) <= a;
    layer2_outputs(10055) <= 1'b1;
    layer2_outputs(10056) <= a and not b;
    layer2_outputs(10057) <= not (a and b);
    layer2_outputs(10058) <= not a;
    layer2_outputs(10059) <= a and not b;
    layer2_outputs(10060) <= not (a xor b);
    layer2_outputs(10061) <= a or b;
    layer2_outputs(10062) <= a or b;
    layer2_outputs(10063) <= not a or b;
    layer2_outputs(10064) <= not b or a;
    layer2_outputs(10065) <= not a or b;
    layer2_outputs(10066) <= b and not a;
    layer2_outputs(10067) <= b;
    layer2_outputs(10068) <= a and not b;
    layer2_outputs(10069) <= b and not a;
    layer2_outputs(10070) <= a;
    layer2_outputs(10071) <= not b;
    layer2_outputs(10072) <= a;
    layer2_outputs(10073) <= 1'b0;
    layer2_outputs(10074) <= b;
    layer2_outputs(10075) <= a;
    layer2_outputs(10076) <= b and not a;
    layer2_outputs(10077) <= not b or a;
    layer2_outputs(10078) <= a or b;
    layer2_outputs(10079) <= a and not b;
    layer2_outputs(10080) <= not (a or b);
    layer2_outputs(10081) <= a and not b;
    layer2_outputs(10082) <= not a;
    layer2_outputs(10083) <= a;
    layer2_outputs(10084) <= b and not a;
    layer2_outputs(10085) <= a and b;
    layer2_outputs(10086) <= 1'b1;
    layer2_outputs(10087) <= not (a or b);
    layer2_outputs(10088) <= not b or a;
    layer2_outputs(10089) <= not b;
    layer2_outputs(10090) <= not a or b;
    layer2_outputs(10091) <= a or b;
    layer2_outputs(10092) <= a and b;
    layer2_outputs(10093) <= not (a or b);
    layer2_outputs(10094) <= a;
    layer2_outputs(10095) <= 1'b1;
    layer2_outputs(10096) <= a and b;
    layer2_outputs(10097) <= b;
    layer2_outputs(10098) <= a;
    layer2_outputs(10099) <= not (a and b);
    layer2_outputs(10100) <= not b;
    layer2_outputs(10101) <= not (a and b);
    layer2_outputs(10102) <= b;
    layer2_outputs(10103) <= not b or a;
    layer2_outputs(10104) <= not (a xor b);
    layer2_outputs(10105) <= not b;
    layer2_outputs(10106) <= not (a and b);
    layer2_outputs(10107) <= a and not b;
    layer2_outputs(10108) <= not a or b;
    layer2_outputs(10109) <= a;
    layer2_outputs(10110) <= a and b;
    layer2_outputs(10111) <= not a or b;
    layer2_outputs(10112) <= not b;
    layer2_outputs(10113) <= a and b;
    layer2_outputs(10114) <= 1'b1;
    layer2_outputs(10115) <= not a;
    layer2_outputs(10116) <= not a or b;
    layer2_outputs(10117) <= 1'b0;
    layer2_outputs(10118) <= not a or b;
    layer2_outputs(10119) <= a;
    layer2_outputs(10120) <= not a;
    layer2_outputs(10121) <= not (a or b);
    layer2_outputs(10122) <= a;
    layer2_outputs(10123) <= a or b;
    layer2_outputs(10124) <= a;
    layer2_outputs(10125) <= not a or b;
    layer2_outputs(10126) <= not a;
    layer2_outputs(10127) <= a or b;
    layer2_outputs(10128) <= a or b;
    layer2_outputs(10129) <= b;
    layer2_outputs(10130) <= not (a or b);
    layer2_outputs(10131) <= not a or b;
    layer2_outputs(10132) <= not (a or b);
    layer2_outputs(10133) <= 1'b1;
    layer2_outputs(10134) <= not a;
    layer2_outputs(10135) <= a xor b;
    layer2_outputs(10136) <= not b;
    layer2_outputs(10137) <= not a or b;
    layer2_outputs(10138) <= not (a or b);
    layer2_outputs(10139) <= not b or a;
    layer2_outputs(10140) <= a;
    layer2_outputs(10141) <= not a;
    layer2_outputs(10142) <= a and b;
    layer2_outputs(10143) <= not (a and b);
    layer2_outputs(10144) <= b;
    layer2_outputs(10145) <= not b or a;
    layer2_outputs(10146) <= a and b;
    layer2_outputs(10147) <= a and b;
    layer2_outputs(10148) <= not a or b;
    layer2_outputs(10149) <= a xor b;
    layer2_outputs(10150) <= not b;
    layer2_outputs(10151) <= 1'b1;
    layer2_outputs(10152) <= b;
    layer2_outputs(10153) <= b;
    layer2_outputs(10154) <= a or b;
    layer2_outputs(10155) <= not (a or b);
    layer2_outputs(10156) <= not (a or b);
    layer2_outputs(10157) <= not a;
    layer2_outputs(10158) <= a and not b;
    layer2_outputs(10159) <= a or b;
    layer2_outputs(10160) <= not a or b;
    layer2_outputs(10161) <= b and not a;
    layer2_outputs(10162) <= b and not a;
    layer2_outputs(10163) <= a and b;
    layer2_outputs(10164) <= a xor b;
    layer2_outputs(10165) <= a;
    layer2_outputs(10166) <= not a;
    layer2_outputs(10167) <= b;
    layer2_outputs(10168) <= 1'b0;
    layer2_outputs(10169) <= not b;
    layer2_outputs(10170) <= b and not a;
    layer2_outputs(10171) <= a and not b;
    layer2_outputs(10172) <= not a;
    layer2_outputs(10173) <= not a;
    layer2_outputs(10174) <= a and b;
    layer2_outputs(10175) <= a or b;
    layer2_outputs(10176) <= not a or b;
    layer2_outputs(10177) <= a;
    layer2_outputs(10178) <= not b;
    layer2_outputs(10179) <= not (a xor b);
    layer2_outputs(10180) <= not (a or b);
    layer2_outputs(10181) <= a or b;
    layer2_outputs(10182) <= not b;
    layer2_outputs(10183) <= a or b;
    layer2_outputs(10184) <= not (a or b);
    layer2_outputs(10185) <= not (a or b);
    layer2_outputs(10186) <= b;
    layer2_outputs(10187) <= not b;
    layer2_outputs(10188) <= not (a or b);
    layer2_outputs(10189) <= not b or a;
    layer2_outputs(10190) <= a and b;
    layer2_outputs(10191) <= not b;
    layer2_outputs(10192) <= b;
    layer2_outputs(10193) <= a xor b;
    layer2_outputs(10194) <= not (a xor b);
    layer2_outputs(10195) <= not a;
    layer2_outputs(10196) <= b and not a;
    layer2_outputs(10197) <= a and not b;
    layer2_outputs(10198) <= not a or b;
    layer2_outputs(10199) <= not (a or b);
    layer2_outputs(10200) <= b and not a;
    layer2_outputs(10201) <= not a or b;
    layer2_outputs(10202) <= not a;
    layer2_outputs(10203) <= a and not b;
    layer2_outputs(10204) <= not b;
    layer2_outputs(10205) <= a;
    layer2_outputs(10206) <= not (a and b);
    layer2_outputs(10207) <= a or b;
    layer2_outputs(10208) <= b;
    layer2_outputs(10209) <= not (a and b);
    layer2_outputs(10210) <= a and b;
    layer2_outputs(10211) <= not b;
    layer2_outputs(10212) <= 1'b1;
    layer2_outputs(10213) <= not (a xor b);
    layer2_outputs(10214) <= a or b;
    layer2_outputs(10215) <= a;
    layer2_outputs(10216) <= a and b;
    layer2_outputs(10217) <= a and b;
    layer2_outputs(10218) <= not a or b;
    layer2_outputs(10219) <= a xor b;
    layer2_outputs(10220) <= b;
    layer2_outputs(10221) <= not (a xor b);
    layer2_outputs(10222) <= a or b;
    layer2_outputs(10223) <= not b;
    layer2_outputs(10224) <= not (a or b);
    layer2_outputs(10225) <= a;
    layer2_outputs(10226) <= not a;
    layer2_outputs(10227) <= not a;
    layer2_outputs(10228) <= a and not b;
    layer2_outputs(10229) <= not a or b;
    layer2_outputs(10230) <= a xor b;
    layer2_outputs(10231) <= a or b;
    layer2_outputs(10232) <= a and b;
    layer2_outputs(10233) <= b;
    layer2_outputs(10234) <= not b;
    layer2_outputs(10235) <= not b or a;
    layer2_outputs(10236) <= not b or a;
    layer2_outputs(10237) <= b;
    layer2_outputs(10238) <= a xor b;
    layer2_outputs(10239) <= a;
    layer3_outputs(0) <= not (a xor b);
    layer3_outputs(1) <= a;
    layer3_outputs(2) <= 1'b1;
    layer3_outputs(3) <= a and not b;
    layer3_outputs(4) <= a xor b;
    layer3_outputs(5) <= b and not a;
    layer3_outputs(6) <= b;
    layer3_outputs(7) <= a and not b;
    layer3_outputs(8) <= not a;
    layer3_outputs(9) <= a and b;
    layer3_outputs(10) <= not a;
    layer3_outputs(11) <= a;
    layer3_outputs(12) <= not a;
    layer3_outputs(13) <= not a or b;
    layer3_outputs(14) <= b;
    layer3_outputs(15) <= not a;
    layer3_outputs(16) <= 1'b1;
    layer3_outputs(17) <= not a;
    layer3_outputs(18) <= a and b;
    layer3_outputs(19) <= b;
    layer3_outputs(20) <= not (a xor b);
    layer3_outputs(21) <= not a or b;
    layer3_outputs(22) <= not a;
    layer3_outputs(23) <= not (a or b);
    layer3_outputs(24) <= a or b;
    layer3_outputs(25) <= not (a and b);
    layer3_outputs(26) <= not a;
    layer3_outputs(27) <= a;
    layer3_outputs(28) <= not a;
    layer3_outputs(29) <= not a;
    layer3_outputs(30) <= b;
    layer3_outputs(31) <= not (a xor b);
    layer3_outputs(32) <= not b;
    layer3_outputs(33) <= a;
    layer3_outputs(34) <= not b;
    layer3_outputs(35) <= not (a and b);
    layer3_outputs(36) <= not a;
    layer3_outputs(37) <= not (a xor b);
    layer3_outputs(38) <= b and not a;
    layer3_outputs(39) <= a;
    layer3_outputs(40) <= not (a or b);
    layer3_outputs(41) <= not b;
    layer3_outputs(42) <= not b;
    layer3_outputs(43) <= b and not a;
    layer3_outputs(44) <= b and not a;
    layer3_outputs(45) <= b and not a;
    layer3_outputs(46) <= not (a xor b);
    layer3_outputs(47) <= a and b;
    layer3_outputs(48) <= b;
    layer3_outputs(49) <= not (a and b);
    layer3_outputs(50) <= not b;
    layer3_outputs(51) <= not (a or b);
    layer3_outputs(52) <= not b;
    layer3_outputs(53) <= a or b;
    layer3_outputs(54) <= not a;
    layer3_outputs(55) <= not b;
    layer3_outputs(56) <= not b or a;
    layer3_outputs(57) <= not a;
    layer3_outputs(58) <= not b;
    layer3_outputs(59) <= b;
    layer3_outputs(60) <= not b;
    layer3_outputs(61) <= not a or b;
    layer3_outputs(62) <= a;
    layer3_outputs(63) <= not b;
    layer3_outputs(64) <= a and b;
    layer3_outputs(65) <= a or b;
    layer3_outputs(66) <= not (a and b);
    layer3_outputs(67) <= b;
    layer3_outputs(68) <= not b or a;
    layer3_outputs(69) <= not (a and b);
    layer3_outputs(70) <= a and b;
    layer3_outputs(71) <= a and b;
    layer3_outputs(72) <= not a;
    layer3_outputs(73) <= b;
    layer3_outputs(74) <= not a;
    layer3_outputs(75) <= not b;
    layer3_outputs(76) <= a or b;
    layer3_outputs(77) <= not b;
    layer3_outputs(78) <= not (a and b);
    layer3_outputs(79) <= a and b;
    layer3_outputs(80) <= a and not b;
    layer3_outputs(81) <= a and not b;
    layer3_outputs(82) <= a;
    layer3_outputs(83) <= not b;
    layer3_outputs(84) <= not (a or b);
    layer3_outputs(85) <= not b or a;
    layer3_outputs(86) <= not (a or b);
    layer3_outputs(87) <= a;
    layer3_outputs(88) <= b;
    layer3_outputs(89) <= not (a or b);
    layer3_outputs(90) <= b;
    layer3_outputs(91) <= not (a and b);
    layer3_outputs(92) <= a;
    layer3_outputs(93) <= not b;
    layer3_outputs(94) <= b and not a;
    layer3_outputs(95) <= not (a and b);
    layer3_outputs(96) <= not a or b;
    layer3_outputs(97) <= a or b;
    layer3_outputs(98) <= b and not a;
    layer3_outputs(99) <= not b;
    layer3_outputs(100) <= not a or b;
    layer3_outputs(101) <= not b;
    layer3_outputs(102) <= a or b;
    layer3_outputs(103) <= a xor b;
    layer3_outputs(104) <= not (a and b);
    layer3_outputs(105) <= not (a and b);
    layer3_outputs(106) <= not (a or b);
    layer3_outputs(107) <= a or b;
    layer3_outputs(108) <= a xor b;
    layer3_outputs(109) <= not a or b;
    layer3_outputs(110) <= not a;
    layer3_outputs(111) <= not a or b;
    layer3_outputs(112) <= not a;
    layer3_outputs(113) <= not a;
    layer3_outputs(114) <= a xor b;
    layer3_outputs(115) <= not a or b;
    layer3_outputs(116) <= b;
    layer3_outputs(117) <= not b;
    layer3_outputs(118) <= not b;
    layer3_outputs(119) <= not b or a;
    layer3_outputs(120) <= a;
    layer3_outputs(121) <= not b or a;
    layer3_outputs(122) <= b and not a;
    layer3_outputs(123) <= not (a and b);
    layer3_outputs(124) <= b and not a;
    layer3_outputs(125) <= a xor b;
    layer3_outputs(126) <= a xor b;
    layer3_outputs(127) <= a xor b;
    layer3_outputs(128) <= b;
    layer3_outputs(129) <= not a;
    layer3_outputs(130) <= not b;
    layer3_outputs(131) <= a;
    layer3_outputs(132) <= a;
    layer3_outputs(133) <= b;
    layer3_outputs(134) <= not a;
    layer3_outputs(135) <= a xor b;
    layer3_outputs(136) <= not b;
    layer3_outputs(137) <= a xor b;
    layer3_outputs(138) <= a;
    layer3_outputs(139) <= a and not b;
    layer3_outputs(140) <= not (a or b);
    layer3_outputs(141) <= not (a xor b);
    layer3_outputs(142) <= 1'b1;
    layer3_outputs(143) <= a;
    layer3_outputs(144) <= a and b;
    layer3_outputs(145) <= a and b;
    layer3_outputs(146) <= a;
    layer3_outputs(147) <= not (a or b);
    layer3_outputs(148) <= not a;
    layer3_outputs(149) <= 1'b1;
    layer3_outputs(150) <= a or b;
    layer3_outputs(151) <= b;
    layer3_outputs(152) <= not (a and b);
    layer3_outputs(153) <= a or b;
    layer3_outputs(154) <= not a;
    layer3_outputs(155) <= a xor b;
    layer3_outputs(156) <= not (a xor b);
    layer3_outputs(157) <= not a or b;
    layer3_outputs(158) <= b;
    layer3_outputs(159) <= not b;
    layer3_outputs(160) <= a;
    layer3_outputs(161) <= not (a xor b);
    layer3_outputs(162) <= a and not b;
    layer3_outputs(163) <= not b or a;
    layer3_outputs(164) <= a xor b;
    layer3_outputs(165) <= not (a or b);
    layer3_outputs(166) <= a;
    layer3_outputs(167) <= not b;
    layer3_outputs(168) <= a or b;
    layer3_outputs(169) <= not b;
    layer3_outputs(170) <= not (a and b);
    layer3_outputs(171) <= not (a and b);
    layer3_outputs(172) <= a;
    layer3_outputs(173) <= not (a or b);
    layer3_outputs(174) <= not (a or b);
    layer3_outputs(175) <= b;
    layer3_outputs(176) <= not (a and b);
    layer3_outputs(177) <= not b or a;
    layer3_outputs(178) <= not (a and b);
    layer3_outputs(179) <= not a;
    layer3_outputs(180) <= b and not a;
    layer3_outputs(181) <= b;
    layer3_outputs(182) <= a and b;
    layer3_outputs(183) <= a and b;
    layer3_outputs(184) <= a and b;
    layer3_outputs(185) <= a and b;
    layer3_outputs(186) <= a and not b;
    layer3_outputs(187) <= a and b;
    layer3_outputs(188) <= b;
    layer3_outputs(189) <= not (a and b);
    layer3_outputs(190) <= a;
    layer3_outputs(191) <= not a;
    layer3_outputs(192) <= not a or b;
    layer3_outputs(193) <= not a;
    layer3_outputs(194) <= b and not a;
    layer3_outputs(195) <= not (a xor b);
    layer3_outputs(196) <= a and b;
    layer3_outputs(197) <= not b or a;
    layer3_outputs(198) <= not (a or b);
    layer3_outputs(199) <= a or b;
    layer3_outputs(200) <= not (a or b);
    layer3_outputs(201) <= not a;
    layer3_outputs(202) <= b;
    layer3_outputs(203) <= not b;
    layer3_outputs(204) <= a and b;
    layer3_outputs(205) <= 1'b0;
    layer3_outputs(206) <= not (a and b);
    layer3_outputs(207) <= not (a xor b);
    layer3_outputs(208) <= b;
    layer3_outputs(209) <= b;
    layer3_outputs(210) <= a;
    layer3_outputs(211) <= a;
    layer3_outputs(212) <= not (a and b);
    layer3_outputs(213) <= b;
    layer3_outputs(214) <= not (a or b);
    layer3_outputs(215) <= a;
    layer3_outputs(216) <= a and b;
    layer3_outputs(217) <= a and not b;
    layer3_outputs(218) <= not (a or b);
    layer3_outputs(219) <= not b;
    layer3_outputs(220) <= a;
    layer3_outputs(221) <= not (a and b);
    layer3_outputs(222) <= b and not a;
    layer3_outputs(223) <= b and not a;
    layer3_outputs(224) <= b;
    layer3_outputs(225) <= not (a or b);
    layer3_outputs(226) <= b;
    layer3_outputs(227) <= b and not a;
    layer3_outputs(228) <= not b or a;
    layer3_outputs(229) <= not a or b;
    layer3_outputs(230) <= a and b;
    layer3_outputs(231) <= not b;
    layer3_outputs(232) <= a;
    layer3_outputs(233) <= a or b;
    layer3_outputs(234) <= not (a xor b);
    layer3_outputs(235) <= not b;
    layer3_outputs(236) <= not (a xor b);
    layer3_outputs(237) <= b and not a;
    layer3_outputs(238) <= a;
    layer3_outputs(239) <= b;
    layer3_outputs(240) <= not (a or b);
    layer3_outputs(241) <= not (a and b);
    layer3_outputs(242) <= a or b;
    layer3_outputs(243) <= b;
    layer3_outputs(244) <= a;
    layer3_outputs(245) <= not a;
    layer3_outputs(246) <= b and not a;
    layer3_outputs(247) <= a and not b;
    layer3_outputs(248) <= a or b;
    layer3_outputs(249) <= a or b;
    layer3_outputs(250) <= not b;
    layer3_outputs(251) <= b;
    layer3_outputs(252) <= a xor b;
    layer3_outputs(253) <= b and not a;
    layer3_outputs(254) <= b;
    layer3_outputs(255) <= not a;
    layer3_outputs(256) <= not b or a;
    layer3_outputs(257) <= b;
    layer3_outputs(258) <= not b or a;
    layer3_outputs(259) <= not b;
    layer3_outputs(260) <= b and not a;
    layer3_outputs(261) <= a and b;
    layer3_outputs(262) <= a xor b;
    layer3_outputs(263) <= b;
    layer3_outputs(264) <= not b;
    layer3_outputs(265) <= not a;
    layer3_outputs(266) <= not a;
    layer3_outputs(267) <= not (a and b);
    layer3_outputs(268) <= a;
    layer3_outputs(269) <= a and b;
    layer3_outputs(270) <= not a or b;
    layer3_outputs(271) <= not a;
    layer3_outputs(272) <= not b or a;
    layer3_outputs(273) <= not (a and b);
    layer3_outputs(274) <= not a or b;
    layer3_outputs(275) <= not b;
    layer3_outputs(276) <= a and b;
    layer3_outputs(277) <= not (a xor b);
    layer3_outputs(278) <= not a;
    layer3_outputs(279) <= a and b;
    layer3_outputs(280) <= not a or b;
    layer3_outputs(281) <= not (a and b);
    layer3_outputs(282) <= not (a and b);
    layer3_outputs(283) <= a;
    layer3_outputs(284) <= not (a and b);
    layer3_outputs(285) <= not b;
    layer3_outputs(286) <= b and not a;
    layer3_outputs(287) <= b;
    layer3_outputs(288) <= a and b;
    layer3_outputs(289) <= not b or a;
    layer3_outputs(290) <= b and not a;
    layer3_outputs(291) <= not (a xor b);
    layer3_outputs(292) <= a or b;
    layer3_outputs(293) <= not b;
    layer3_outputs(294) <= a xor b;
    layer3_outputs(295) <= a or b;
    layer3_outputs(296) <= a and b;
    layer3_outputs(297) <= not (a or b);
    layer3_outputs(298) <= not b;
    layer3_outputs(299) <= not b;
    layer3_outputs(300) <= not a;
    layer3_outputs(301) <= not a or b;
    layer3_outputs(302) <= a xor b;
    layer3_outputs(303) <= not (a xor b);
    layer3_outputs(304) <= a;
    layer3_outputs(305) <= not a;
    layer3_outputs(306) <= a;
    layer3_outputs(307) <= not a;
    layer3_outputs(308) <= not (a and b);
    layer3_outputs(309) <= 1'b1;
    layer3_outputs(310) <= not a or b;
    layer3_outputs(311) <= b;
    layer3_outputs(312) <= not b or a;
    layer3_outputs(313) <= not a;
    layer3_outputs(314) <= a or b;
    layer3_outputs(315) <= a;
    layer3_outputs(316) <= not a;
    layer3_outputs(317) <= not a or b;
    layer3_outputs(318) <= a;
    layer3_outputs(319) <= b and not a;
    layer3_outputs(320) <= a or b;
    layer3_outputs(321) <= a;
    layer3_outputs(322) <= b;
    layer3_outputs(323) <= not b;
    layer3_outputs(324) <= a and b;
    layer3_outputs(325) <= a xor b;
    layer3_outputs(326) <= not b;
    layer3_outputs(327) <= not b;
    layer3_outputs(328) <= not a or b;
    layer3_outputs(329) <= not a or b;
    layer3_outputs(330) <= a;
    layer3_outputs(331) <= not a or b;
    layer3_outputs(332) <= not b;
    layer3_outputs(333) <= not (a and b);
    layer3_outputs(334) <= not a;
    layer3_outputs(335) <= a xor b;
    layer3_outputs(336) <= b and not a;
    layer3_outputs(337) <= a or b;
    layer3_outputs(338) <= b;
    layer3_outputs(339) <= not a;
    layer3_outputs(340) <= a and not b;
    layer3_outputs(341) <= not b or a;
    layer3_outputs(342) <= not (a xor b);
    layer3_outputs(343) <= a and not b;
    layer3_outputs(344) <= a;
    layer3_outputs(345) <= not b or a;
    layer3_outputs(346) <= a and b;
    layer3_outputs(347) <= not b or a;
    layer3_outputs(348) <= b and not a;
    layer3_outputs(349) <= not (a xor b);
    layer3_outputs(350) <= not b;
    layer3_outputs(351) <= a;
    layer3_outputs(352) <= a and not b;
    layer3_outputs(353) <= 1'b0;
    layer3_outputs(354) <= not a;
    layer3_outputs(355) <= a or b;
    layer3_outputs(356) <= not b;
    layer3_outputs(357) <= not (a xor b);
    layer3_outputs(358) <= b;
    layer3_outputs(359) <= not b;
    layer3_outputs(360) <= not b;
    layer3_outputs(361) <= not b or a;
    layer3_outputs(362) <= b;
    layer3_outputs(363) <= not (a and b);
    layer3_outputs(364) <= b;
    layer3_outputs(365) <= b and not a;
    layer3_outputs(366) <= not (a or b);
    layer3_outputs(367) <= not a;
    layer3_outputs(368) <= a xor b;
    layer3_outputs(369) <= 1'b0;
    layer3_outputs(370) <= not b;
    layer3_outputs(371) <= not (a xor b);
    layer3_outputs(372) <= a;
    layer3_outputs(373) <= not b;
    layer3_outputs(374) <= b;
    layer3_outputs(375) <= a and b;
    layer3_outputs(376) <= not (a xor b);
    layer3_outputs(377) <= not (a xor b);
    layer3_outputs(378) <= not (a and b);
    layer3_outputs(379) <= a;
    layer3_outputs(380) <= a and b;
    layer3_outputs(381) <= not (a and b);
    layer3_outputs(382) <= a and not b;
    layer3_outputs(383) <= not a;
    layer3_outputs(384) <= not (a or b);
    layer3_outputs(385) <= not (a and b);
    layer3_outputs(386) <= not (a xor b);
    layer3_outputs(387) <= not b or a;
    layer3_outputs(388) <= b;
    layer3_outputs(389) <= b;
    layer3_outputs(390) <= not b or a;
    layer3_outputs(391) <= a xor b;
    layer3_outputs(392) <= not (a and b);
    layer3_outputs(393) <= not a;
    layer3_outputs(394) <= 1'b0;
    layer3_outputs(395) <= a;
    layer3_outputs(396) <= b;
    layer3_outputs(397) <= a and not b;
    layer3_outputs(398) <= b and not a;
    layer3_outputs(399) <= a;
    layer3_outputs(400) <= a xor b;
    layer3_outputs(401) <= a and b;
    layer3_outputs(402) <= a and b;
    layer3_outputs(403) <= not a;
    layer3_outputs(404) <= b and not a;
    layer3_outputs(405) <= b;
    layer3_outputs(406) <= not a;
    layer3_outputs(407) <= a or b;
    layer3_outputs(408) <= a and not b;
    layer3_outputs(409) <= b;
    layer3_outputs(410) <= not a or b;
    layer3_outputs(411) <= not (a or b);
    layer3_outputs(412) <= a xor b;
    layer3_outputs(413) <= a;
    layer3_outputs(414) <= a and not b;
    layer3_outputs(415) <= not b;
    layer3_outputs(416) <= not a;
    layer3_outputs(417) <= a;
    layer3_outputs(418) <= b;
    layer3_outputs(419) <= a and not b;
    layer3_outputs(420) <= not b or a;
    layer3_outputs(421) <= a xor b;
    layer3_outputs(422) <= a or b;
    layer3_outputs(423) <= not b or a;
    layer3_outputs(424) <= not (a or b);
    layer3_outputs(425) <= not (a and b);
    layer3_outputs(426) <= b;
    layer3_outputs(427) <= not b or a;
    layer3_outputs(428) <= a;
    layer3_outputs(429) <= not b;
    layer3_outputs(430) <= not b or a;
    layer3_outputs(431) <= a or b;
    layer3_outputs(432) <= not b;
    layer3_outputs(433) <= a and not b;
    layer3_outputs(434) <= b;
    layer3_outputs(435) <= b;
    layer3_outputs(436) <= not b;
    layer3_outputs(437) <= b and not a;
    layer3_outputs(438) <= not a or b;
    layer3_outputs(439) <= not (a and b);
    layer3_outputs(440) <= not (a xor b);
    layer3_outputs(441) <= not a or b;
    layer3_outputs(442) <= b;
    layer3_outputs(443) <= not a;
    layer3_outputs(444) <= b;
    layer3_outputs(445) <= a xor b;
    layer3_outputs(446) <= a and not b;
    layer3_outputs(447) <= not (a or b);
    layer3_outputs(448) <= not (a xor b);
    layer3_outputs(449) <= a and not b;
    layer3_outputs(450) <= not (a xor b);
    layer3_outputs(451) <= a;
    layer3_outputs(452) <= not a;
    layer3_outputs(453) <= not a;
    layer3_outputs(454) <= not (a xor b);
    layer3_outputs(455) <= not b;
    layer3_outputs(456) <= not a or b;
    layer3_outputs(457) <= not a;
    layer3_outputs(458) <= a xor b;
    layer3_outputs(459) <= b and not a;
    layer3_outputs(460) <= not a;
    layer3_outputs(461) <= not (a and b);
    layer3_outputs(462) <= b;
    layer3_outputs(463) <= not (a xor b);
    layer3_outputs(464) <= not (a and b);
    layer3_outputs(465) <= b and not a;
    layer3_outputs(466) <= not b or a;
    layer3_outputs(467) <= a;
    layer3_outputs(468) <= a;
    layer3_outputs(469) <= not a;
    layer3_outputs(470) <= b;
    layer3_outputs(471) <= not b;
    layer3_outputs(472) <= not a;
    layer3_outputs(473) <= not a;
    layer3_outputs(474) <= not a;
    layer3_outputs(475) <= a;
    layer3_outputs(476) <= a xor b;
    layer3_outputs(477) <= not (a and b);
    layer3_outputs(478) <= a;
    layer3_outputs(479) <= b;
    layer3_outputs(480) <= a;
    layer3_outputs(481) <= not a or b;
    layer3_outputs(482) <= not a;
    layer3_outputs(483) <= b;
    layer3_outputs(484) <= a;
    layer3_outputs(485) <= b;
    layer3_outputs(486) <= not (a and b);
    layer3_outputs(487) <= not a;
    layer3_outputs(488) <= not (a xor b);
    layer3_outputs(489) <= a;
    layer3_outputs(490) <= a;
    layer3_outputs(491) <= not b or a;
    layer3_outputs(492) <= not b or a;
    layer3_outputs(493) <= not b;
    layer3_outputs(494) <= b;
    layer3_outputs(495) <= a xor b;
    layer3_outputs(496) <= b;
    layer3_outputs(497) <= a and b;
    layer3_outputs(498) <= not (a and b);
    layer3_outputs(499) <= a and not b;
    layer3_outputs(500) <= a and not b;
    layer3_outputs(501) <= a and not b;
    layer3_outputs(502) <= not (a or b);
    layer3_outputs(503) <= not a;
    layer3_outputs(504) <= not b or a;
    layer3_outputs(505) <= b and not a;
    layer3_outputs(506) <= not a;
    layer3_outputs(507) <= b;
    layer3_outputs(508) <= not a or b;
    layer3_outputs(509) <= not (a and b);
    layer3_outputs(510) <= a;
    layer3_outputs(511) <= 1'b0;
    layer3_outputs(512) <= not a or b;
    layer3_outputs(513) <= b;
    layer3_outputs(514) <= a;
    layer3_outputs(515) <= a and not b;
    layer3_outputs(516) <= not b;
    layer3_outputs(517) <= not (a and b);
    layer3_outputs(518) <= not a;
    layer3_outputs(519) <= not (a and b);
    layer3_outputs(520) <= a or b;
    layer3_outputs(521) <= a xor b;
    layer3_outputs(522) <= b and not a;
    layer3_outputs(523) <= b;
    layer3_outputs(524) <= b and not a;
    layer3_outputs(525) <= not (a and b);
    layer3_outputs(526) <= a;
    layer3_outputs(527) <= a xor b;
    layer3_outputs(528) <= b;
    layer3_outputs(529) <= a xor b;
    layer3_outputs(530) <= not (a or b);
    layer3_outputs(531) <= not a;
    layer3_outputs(532) <= a;
    layer3_outputs(533) <= not a;
    layer3_outputs(534) <= not b;
    layer3_outputs(535) <= a and b;
    layer3_outputs(536) <= b;
    layer3_outputs(537) <= not a;
    layer3_outputs(538) <= a;
    layer3_outputs(539) <= a and b;
    layer3_outputs(540) <= not b or a;
    layer3_outputs(541) <= b;
    layer3_outputs(542) <= not (a and b);
    layer3_outputs(543) <= a xor b;
    layer3_outputs(544) <= a and b;
    layer3_outputs(545) <= a xor b;
    layer3_outputs(546) <= a xor b;
    layer3_outputs(547) <= not (a xor b);
    layer3_outputs(548) <= b;
    layer3_outputs(549) <= not b or a;
    layer3_outputs(550) <= a or b;
    layer3_outputs(551) <= a;
    layer3_outputs(552) <= not b;
    layer3_outputs(553) <= not b;
    layer3_outputs(554) <= not a;
    layer3_outputs(555) <= not b;
    layer3_outputs(556) <= a;
    layer3_outputs(557) <= b and not a;
    layer3_outputs(558) <= not (a and b);
    layer3_outputs(559) <= a and b;
    layer3_outputs(560) <= not b;
    layer3_outputs(561) <= a and b;
    layer3_outputs(562) <= not b;
    layer3_outputs(563) <= not b;
    layer3_outputs(564) <= not (a or b);
    layer3_outputs(565) <= not (a or b);
    layer3_outputs(566) <= not (a and b);
    layer3_outputs(567) <= not b;
    layer3_outputs(568) <= a;
    layer3_outputs(569) <= not a or b;
    layer3_outputs(570) <= b;
    layer3_outputs(571) <= a;
    layer3_outputs(572) <= not (a xor b);
    layer3_outputs(573) <= not b or a;
    layer3_outputs(574) <= not b or a;
    layer3_outputs(575) <= not a;
    layer3_outputs(576) <= a or b;
    layer3_outputs(577) <= a xor b;
    layer3_outputs(578) <= not a;
    layer3_outputs(579) <= not a or b;
    layer3_outputs(580) <= not (a or b);
    layer3_outputs(581) <= a and not b;
    layer3_outputs(582) <= not a;
    layer3_outputs(583) <= not (a and b);
    layer3_outputs(584) <= not b;
    layer3_outputs(585) <= a and b;
    layer3_outputs(586) <= not a;
    layer3_outputs(587) <= not b;
    layer3_outputs(588) <= a;
    layer3_outputs(589) <= not (a xor b);
    layer3_outputs(590) <= b;
    layer3_outputs(591) <= a xor b;
    layer3_outputs(592) <= 1'b0;
    layer3_outputs(593) <= a and not b;
    layer3_outputs(594) <= b;
    layer3_outputs(595) <= not a or b;
    layer3_outputs(596) <= not a;
    layer3_outputs(597) <= b;
    layer3_outputs(598) <= not a;
    layer3_outputs(599) <= not b or a;
    layer3_outputs(600) <= not b;
    layer3_outputs(601) <= a and not b;
    layer3_outputs(602) <= not b;
    layer3_outputs(603) <= b and not a;
    layer3_outputs(604) <= a and not b;
    layer3_outputs(605) <= b and not a;
    layer3_outputs(606) <= a and b;
    layer3_outputs(607) <= b;
    layer3_outputs(608) <= not b;
    layer3_outputs(609) <= not (a and b);
    layer3_outputs(610) <= not a;
    layer3_outputs(611) <= a xor b;
    layer3_outputs(612) <= not b;
    layer3_outputs(613) <= not (a xor b);
    layer3_outputs(614) <= not (a or b);
    layer3_outputs(615) <= not b or a;
    layer3_outputs(616) <= not (a xor b);
    layer3_outputs(617) <= b;
    layer3_outputs(618) <= a xor b;
    layer3_outputs(619) <= a or b;
    layer3_outputs(620) <= not a;
    layer3_outputs(621) <= b;
    layer3_outputs(622) <= b;
    layer3_outputs(623) <= a and b;
    layer3_outputs(624) <= not a or b;
    layer3_outputs(625) <= a and not b;
    layer3_outputs(626) <= not (a and b);
    layer3_outputs(627) <= a;
    layer3_outputs(628) <= b;
    layer3_outputs(629) <= b;
    layer3_outputs(630) <= not (a xor b);
    layer3_outputs(631) <= not a;
    layer3_outputs(632) <= not b;
    layer3_outputs(633) <= a;
    layer3_outputs(634) <= a xor b;
    layer3_outputs(635) <= a and b;
    layer3_outputs(636) <= not a or b;
    layer3_outputs(637) <= a xor b;
    layer3_outputs(638) <= not b or a;
    layer3_outputs(639) <= a and not b;
    layer3_outputs(640) <= not a or b;
    layer3_outputs(641) <= a and b;
    layer3_outputs(642) <= not b or a;
    layer3_outputs(643) <= a;
    layer3_outputs(644) <= not (a xor b);
    layer3_outputs(645) <= not (a and b);
    layer3_outputs(646) <= 1'b0;
    layer3_outputs(647) <= a;
    layer3_outputs(648) <= 1'b1;
    layer3_outputs(649) <= a or b;
    layer3_outputs(650) <= not a;
    layer3_outputs(651) <= a;
    layer3_outputs(652) <= not (a and b);
    layer3_outputs(653) <= not (a xor b);
    layer3_outputs(654) <= a and b;
    layer3_outputs(655) <= not b or a;
    layer3_outputs(656) <= a and not b;
    layer3_outputs(657) <= not b;
    layer3_outputs(658) <= not b;
    layer3_outputs(659) <= not (a or b);
    layer3_outputs(660) <= b and not a;
    layer3_outputs(661) <= b;
    layer3_outputs(662) <= not b;
    layer3_outputs(663) <= a xor b;
    layer3_outputs(664) <= not b;
    layer3_outputs(665) <= not a or b;
    layer3_outputs(666) <= b;
    layer3_outputs(667) <= not b;
    layer3_outputs(668) <= b;
    layer3_outputs(669) <= a xor b;
    layer3_outputs(670) <= not a;
    layer3_outputs(671) <= b and not a;
    layer3_outputs(672) <= not (a xor b);
    layer3_outputs(673) <= not b;
    layer3_outputs(674) <= b;
    layer3_outputs(675) <= not a;
    layer3_outputs(676) <= a;
    layer3_outputs(677) <= b;
    layer3_outputs(678) <= not (a and b);
    layer3_outputs(679) <= b;
    layer3_outputs(680) <= 1'b1;
    layer3_outputs(681) <= not (a or b);
    layer3_outputs(682) <= a and b;
    layer3_outputs(683) <= b and not a;
    layer3_outputs(684) <= not a;
    layer3_outputs(685) <= a;
    layer3_outputs(686) <= b;
    layer3_outputs(687) <= b and not a;
    layer3_outputs(688) <= a;
    layer3_outputs(689) <= a;
    layer3_outputs(690) <= not b;
    layer3_outputs(691) <= a and not b;
    layer3_outputs(692) <= a;
    layer3_outputs(693) <= not b or a;
    layer3_outputs(694) <= not (a and b);
    layer3_outputs(695) <= not b or a;
    layer3_outputs(696) <= a xor b;
    layer3_outputs(697) <= a and b;
    layer3_outputs(698) <= not (a xor b);
    layer3_outputs(699) <= not b;
    layer3_outputs(700) <= not a;
    layer3_outputs(701) <= not b;
    layer3_outputs(702) <= not a;
    layer3_outputs(703) <= not b;
    layer3_outputs(704) <= not a;
    layer3_outputs(705) <= not (a xor b);
    layer3_outputs(706) <= not a;
    layer3_outputs(707) <= a or b;
    layer3_outputs(708) <= not a;
    layer3_outputs(709) <= not a;
    layer3_outputs(710) <= a and b;
    layer3_outputs(711) <= b and not a;
    layer3_outputs(712) <= b;
    layer3_outputs(713) <= a xor b;
    layer3_outputs(714) <= a or b;
    layer3_outputs(715) <= not a;
    layer3_outputs(716) <= a and b;
    layer3_outputs(717) <= not b;
    layer3_outputs(718) <= 1'b0;
    layer3_outputs(719) <= a and b;
    layer3_outputs(720) <= a and b;
    layer3_outputs(721) <= a or b;
    layer3_outputs(722) <= a or b;
    layer3_outputs(723) <= a and not b;
    layer3_outputs(724) <= b;
    layer3_outputs(725) <= a or b;
    layer3_outputs(726) <= b;
    layer3_outputs(727) <= a or b;
    layer3_outputs(728) <= not a;
    layer3_outputs(729) <= not b;
    layer3_outputs(730) <= not b;
    layer3_outputs(731) <= b;
    layer3_outputs(732) <= b and not a;
    layer3_outputs(733) <= not (a xor b);
    layer3_outputs(734) <= not (a or b);
    layer3_outputs(735) <= b;
    layer3_outputs(736) <= not a;
    layer3_outputs(737) <= not b or a;
    layer3_outputs(738) <= a;
    layer3_outputs(739) <= not b;
    layer3_outputs(740) <= not (a xor b);
    layer3_outputs(741) <= b;
    layer3_outputs(742) <= 1'b1;
    layer3_outputs(743) <= not a;
    layer3_outputs(744) <= not a or b;
    layer3_outputs(745) <= 1'b0;
    layer3_outputs(746) <= not (a xor b);
    layer3_outputs(747) <= a xor b;
    layer3_outputs(748) <= a;
    layer3_outputs(749) <= a or b;
    layer3_outputs(750) <= a;
    layer3_outputs(751) <= a and not b;
    layer3_outputs(752) <= b;
    layer3_outputs(753) <= a;
    layer3_outputs(754) <= a or b;
    layer3_outputs(755) <= not (a and b);
    layer3_outputs(756) <= a and b;
    layer3_outputs(757) <= not (a and b);
    layer3_outputs(758) <= b and not a;
    layer3_outputs(759) <= not b;
    layer3_outputs(760) <= not (a xor b);
    layer3_outputs(761) <= not (a xor b);
    layer3_outputs(762) <= a and not b;
    layer3_outputs(763) <= a xor b;
    layer3_outputs(764) <= b;
    layer3_outputs(765) <= b;
    layer3_outputs(766) <= 1'b1;
    layer3_outputs(767) <= not b;
    layer3_outputs(768) <= b and not a;
    layer3_outputs(769) <= a and b;
    layer3_outputs(770) <= a or b;
    layer3_outputs(771) <= b;
    layer3_outputs(772) <= a;
    layer3_outputs(773) <= b;
    layer3_outputs(774) <= not a;
    layer3_outputs(775) <= b and not a;
    layer3_outputs(776) <= a or b;
    layer3_outputs(777) <= b and not a;
    layer3_outputs(778) <= not a or b;
    layer3_outputs(779) <= a and not b;
    layer3_outputs(780) <= a or b;
    layer3_outputs(781) <= 1'b1;
    layer3_outputs(782) <= not (a xor b);
    layer3_outputs(783) <= a xor b;
    layer3_outputs(784) <= not (a xor b);
    layer3_outputs(785) <= a or b;
    layer3_outputs(786) <= not b;
    layer3_outputs(787) <= not (a xor b);
    layer3_outputs(788) <= a or b;
    layer3_outputs(789) <= not a or b;
    layer3_outputs(790) <= a and b;
    layer3_outputs(791) <= b;
    layer3_outputs(792) <= a;
    layer3_outputs(793) <= not a;
    layer3_outputs(794) <= not (a or b);
    layer3_outputs(795) <= not a;
    layer3_outputs(796) <= b;
    layer3_outputs(797) <= not (a xor b);
    layer3_outputs(798) <= b;
    layer3_outputs(799) <= a or b;
    layer3_outputs(800) <= a;
    layer3_outputs(801) <= not (a and b);
    layer3_outputs(802) <= a and not b;
    layer3_outputs(803) <= a and not b;
    layer3_outputs(804) <= not a;
    layer3_outputs(805) <= not (a xor b);
    layer3_outputs(806) <= a;
    layer3_outputs(807) <= not b;
    layer3_outputs(808) <= not a or b;
    layer3_outputs(809) <= b;
    layer3_outputs(810) <= not a;
    layer3_outputs(811) <= a or b;
    layer3_outputs(812) <= a or b;
    layer3_outputs(813) <= a and not b;
    layer3_outputs(814) <= a and b;
    layer3_outputs(815) <= not (a and b);
    layer3_outputs(816) <= a;
    layer3_outputs(817) <= not (a and b);
    layer3_outputs(818) <= b;
    layer3_outputs(819) <= b;
    layer3_outputs(820) <= b;
    layer3_outputs(821) <= not (a xor b);
    layer3_outputs(822) <= a or b;
    layer3_outputs(823) <= b;
    layer3_outputs(824) <= not a;
    layer3_outputs(825) <= a;
    layer3_outputs(826) <= not a;
    layer3_outputs(827) <= not a;
    layer3_outputs(828) <= not a or b;
    layer3_outputs(829) <= b;
    layer3_outputs(830) <= a;
    layer3_outputs(831) <= a xor b;
    layer3_outputs(832) <= a and not b;
    layer3_outputs(833) <= not b or a;
    layer3_outputs(834) <= b;
    layer3_outputs(835) <= not b or a;
    layer3_outputs(836) <= a or b;
    layer3_outputs(837) <= not a;
    layer3_outputs(838) <= not b or a;
    layer3_outputs(839) <= a and not b;
    layer3_outputs(840) <= not b or a;
    layer3_outputs(841) <= a or b;
    layer3_outputs(842) <= not b;
    layer3_outputs(843) <= not (a xor b);
    layer3_outputs(844) <= b;
    layer3_outputs(845) <= b;
    layer3_outputs(846) <= not b or a;
    layer3_outputs(847) <= a;
    layer3_outputs(848) <= not (a or b);
    layer3_outputs(849) <= not (a and b);
    layer3_outputs(850) <= a and b;
    layer3_outputs(851) <= not a;
    layer3_outputs(852) <= not b;
    layer3_outputs(853) <= not (a xor b);
    layer3_outputs(854) <= not (a xor b);
    layer3_outputs(855) <= a and b;
    layer3_outputs(856) <= a;
    layer3_outputs(857) <= a xor b;
    layer3_outputs(858) <= a and not b;
    layer3_outputs(859) <= not (a or b);
    layer3_outputs(860) <= a and not b;
    layer3_outputs(861) <= a and not b;
    layer3_outputs(862) <= not a;
    layer3_outputs(863) <= not (a xor b);
    layer3_outputs(864) <= b;
    layer3_outputs(865) <= not a;
    layer3_outputs(866) <= not (a or b);
    layer3_outputs(867) <= not (a and b);
    layer3_outputs(868) <= b;
    layer3_outputs(869) <= not b;
    layer3_outputs(870) <= b;
    layer3_outputs(871) <= not (a and b);
    layer3_outputs(872) <= b and not a;
    layer3_outputs(873) <= not b;
    layer3_outputs(874) <= b and not a;
    layer3_outputs(875) <= not b or a;
    layer3_outputs(876) <= not (a and b);
    layer3_outputs(877) <= b and not a;
    layer3_outputs(878) <= not b;
    layer3_outputs(879) <= a;
    layer3_outputs(880) <= a and b;
    layer3_outputs(881) <= not a;
    layer3_outputs(882) <= b;
    layer3_outputs(883) <= not b or a;
    layer3_outputs(884) <= a;
    layer3_outputs(885) <= b;
    layer3_outputs(886) <= not b;
    layer3_outputs(887) <= not (a and b);
    layer3_outputs(888) <= not (a and b);
    layer3_outputs(889) <= a or b;
    layer3_outputs(890) <= not a or b;
    layer3_outputs(891) <= a and not b;
    layer3_outputs(892) <= b;
    layer3_outputs(893) <= a;
    layer3_outputs(894) <= b;
    layer3_outputs(895) <= not b;
    layer3_outputs(896) <= not (a xor b);
    layer3_outputs(897) <= b;
    layer3_outputs(898) <= not a;
    layer3_outputs(899) <= not a;
    layer3_outputs(900) <= b;
    layer3_outputs(901) <= b and not a;
    layer3_outputs(902) <= not b;
    layer3_outputs(903) <= not b or a;
    layer3_outputs(904) <= not a or b;
    layer3_outputs(905) <= not b or a;
    layer3_outputs(906) <= a;
    layer3_outputs(907) <= not (a and b);
    layer3_outputs(908) <= a and b;
    layer3_outputs(909) <= not a;
    layer3_outputs(910) <= a;
    layer3_outputs(911) <= 1'b0;
    layer3_outputs(912) <= not a or b;
    layer3_outputs(913) <= a or b;
    layer3_outputs(914) <= not a;
    layer3_outputs(915) <= not b;
    layer3_outputs(916) <= a and b;
    layer3_outputs(917) <= not a;
    layer3_outputs(918) <= not a or b;
    layer3_outputs(919) <= a and not b;
    layer3_outputs(920) <= a xor b;
    layer3_outputs(921) <= a;
    layer3_outputs(922) <= not b;
    layer3_outputs(923) <= not a;
    layer3_outputs(924) <= a;
    layer3_outputs(925) <= not b;
    layer3_outputs(926) <= not (a xor b);
    layer3_outputs(927) <= not (a and b);
    layer3_outputs(928) <= not (a or b);
    layer3_outputs(929) <= a;
    layer3_outputs(930) <= not a;
    layer3_outputs(931) <= a or b;
    layer3_outputs(932) <= not b;
    layer3_outputs(933) <= a xor b;
    layer3_outputs(934) <= not b or a;
    layer3_outputs(935) <= not b or a;
    layer3_outputs(936) <= not (a xor b);
    layer3_outputs(937) <= not b;
    layer3_outputs(938) <= a;
    layer3_outputs(939) <= not b;
    layer3_outputs(940) <= a;
    layer3_outputs(941) <= not b or a;
    layer3_outputs(942) <= b;
    layer3_outputs(943) <= not a;
    layer3_outputs(944) <= not b;
    layer3_outputs(945) <= b and not a;
    layer3_outputs(946) <= b;
    layer3_outputs(947) <= not (a xor b);
    layer3_outputs(948) <= a;
    layer3_outputs(949) <= b and not a;
    layer3_outputs(950) <= not a or b;
    layer3_outputs(951) <= not (a or b);
    layer3_outputs(952) <= not b or a;
    layer3_outputs(953) <= b;
    layer3_outputs(954) <= a or b;
    layer3_outputs(955) <= not b;
    layer3_outputs(956) <= not a or b;
    layer3_outputs(957) <= not b or a;
    layer3_outputs(958) <= not (a or b);
    layer3_outputs(959) <= not (a xor b);
    layer3_outputs(960) <= not (a and b);
    layer3_outputs(961) <= a and not b;
    layer3_outputs(962) <= a and b;
    layer3_outputs(963) <= not (a xor b);
    layer3_outputs(964) <= a or b;
    layer3_outputs(965) <= not a or b;
    layer3_outputs(966) <= not (a and b);
    layer3_outputs(967) <= not (a or b);
    layer3_outputs(968) <= a and not b;
    layer3_outputs(969) <= a or b;
    layer3_outputs(970) <= a;
    layer3_outputs(971) <= not a;
    layer3_outputs(972) <= not a;
    layer3_outputs(973) <= not a or b;
    layer3_outputs(974) <= not a;
    layer3_outputs(975) <= not a;
    layer3_outputs(976) <= a and b;
    layer3_outputs(977) <= not (a or b);
    layer3_outputs(978) <= not a;
    layer3_outputs(979) <= a xor b;
    layer3_outputs(980) <= a;
    layer3_outputs(981) <= not a;
    layer3_outputs(982) <= b and not a;
    layer3_outputs(983) <= b;
    layer3_outputs(984) <= not a;
    layer3_outputs(985) <= not b or a;
    layer3_outputs(986) <= not a;
    layer3_outputs(987) <= not (a and b);
    layer3_outputs(988) <= a xor b;
    layer3_outputs(989) <= b;
    layer3_outputs(990) <= not (a or b);
    layer3_outputs(991) <= not a;
    layer3_outputs(992) <= a;
    layer3_outputs(993) <= b;
    layer3_outputs(994) <= a and not b;
    layer3_outputs(995) <= a;
    layer3_outputs(996) <= not a;
    layer3_outputs(997) <= b;
    layer3_outputs(998) <= not b;
    layer3_outputs(999) <= a;
    layer3_outputs(1000) <= not a;
    layer3_outputs(1001) <= not a;
    layer3_outputs(1002) <= a;
    layer3_outputs(1003) <= not (a and b);
    layer3_outputs(1004) <= not (a and b);
    layer3_outputs(1005) <= not a;
    layer3_outputs(1006) <= a or b;
    layer3_outputs(1007) <= not (a and b);
    layer3_outputs(1008) <= a xor b;
    layer3_outputs(1009) <= a and b;
    layer3_outputs(1010) <= b;
    layer3_outputs(1011) <= not a;
    layer3_outputs(1012) <= b;
    layer3_outputs(1013) <= not a or b;
    layer3_outputs(1014) <= a;
    layer3_outputs(1015) <= b;
    layer3_outputs(1016) <= not a;
    layer3_outputs(1017) <= not (a and b);
    layer3_outputs(1018) <= not (a and b);
    layer3_outputs(1019) <= b;
    layer3_outputs(1020) <= a or b;
    layer3_outputs(1021) <= a and not b;
    layer3_outputs(1022) <= not (a and b);
    layer3_outputs(1023) <= not (a xor b);
    layer3_outputs(1024) <= b and not a;
    layer3_outputs(1025) <= not (a or b);
    layer3_outputs(1026) <= a or b;
    layer3_outputs(1027) <= a;
    layer3_outputs(1028) <= b;
    layer3_outputs(1029) <= a;
    layer3_outputs(1030) <= not b or a;
    layer3_outputs(1031) <= not b or a;
    layer3_outputs(1032) <= not a or b;
    layer3_outputs(1033) <= a or b;
    layer3_outputs(1034) <= not a;
    layer3_outputs(1035) <= not b;
    layer3_outputs(1036) <= a;
    layer3_outputs(1037) <= b;
    layer3_outputs(1038) <= not (a and b);
    layer3_outputs(1039) <= b;
    layer3_outputs(1040) <= a;
    layer3_outputs(1041) <= a and b;
    layer3_outputs(1042) <= not a;
    layer3_outputs(1043) <= b;
    layer3_outputs(1044) <= a or b;
    layer3_outputs(1045) <= not b;
    layer3_outputs(1046) <= not (a or b);
    layer3_outputs(1047) <= not b;
    layer3_outputs(1048) <= a xor b;
    layer3_outputs(1049) <= a and b;
    layer3_outputs(1050) <= not a;
    layer3_outputs(1051) <= a or b;
    layer3_outputs(1052) <= not a;
    layer3_outputs(1053) <= not a or b;
    layer3_outputs(1054) <= not b;
    layer3_outputs(1055) <= not (a and b);
    layer3_outputs(1056) <= not (a xor b);
    layer3_outputs(1057) <= a xor b;
    layer3_outputs(1058) <= not (a xor b);
    layer3_outputs(1059) <= b;
    layer3_outputs(1060) <= not a or b;
    layer3_outputs(1061) <= a or b;
    layer3_outputs(1062) <= b;
    layer3_outputs(1063) <= a or b;
    layer3_outputs(1064) <= not (a or b);
    layer3_outputs(1065) <= not a or b;
    layer3_outputs(1066) <= not (a xor b);
    layer3_outputs(1067) <= not (a or b);
    layer3_outputs(1068) <= a;
    layer3_outputs(1069) <= not (a or b);
    layer3_outputs(1070) <= not (a or b);
    layer3_outputs(1071) <= not a;
    layer3_outputs(1072) <= a;
    layer3_outputs(1073) <= not a;
    layer3_outputs(1074) <= a;
    layer3_outputs(1075) <= a xor b;
    layer3_outputs(1076) <= not b;
    layer3_outputs(1077) <= not (a and b);
    layer3_outputs(1078) <= b and not a;
    layer3_outputs(1079) <= not b or a;
    layer3_outputs(1080) <= a;
    layer3_outputs(1081) <= 1'b0;
    layer3_outputs(1082) <= not a or b;
    layer3_outputs(1083) <= 1'b0;
    layer3_outputs(1084) <= a or b;
    layer3_outputs(1085) <= 1'b0;
    layer3_outputs(1086) <= a xor b;
    layer3_outputs(1087) <= a or b;
    layer3_outputs(1088) <= a and b;
    layer3_outputs(1089) <= not (a and b);
    layer3_outputs(1090) <= a and not b;
    layer3_outputs(1091) <= not (a or b);
    layer3_outputs(1092) <= not b;
    layer3_outputs(1093) <= not (a and b);
    layer3_outputs(1094) <= a or b;
    layer3_outputs(1095) <= b and not a;
    layer3_outputs(1096) <= not (a and b);
    layer3_outputs(1097) <= not a or b;
    layer3_outputs(1098) <= a xor b;
    layer3_outputs(1099) <= b;
    layer3_outputs(1100) <= a;
    layer3_outputs(1101) <= not b or a;
    layer3_outputs(1102) <= not (a or b);
    layer3_outputs(1103) <= not (a and b);
    layer3_outputs(1104) <= a;
    layer3_outputs(1105) <= not a;
    layer3_outputs(1106) <= not b;
    layer3_outputs(1107) <= a or b;
    layer3_outputs(1108) <= not a;
    layer3_outputs(1109) <= b and not a;
    layer3_outputs(1110) <= not a;
    layer3_outputs(1111) <= a and not b;
    layer3_outputs(1112) <= not a;
    layer3_outputs(1113) <= not a;
    layer3_outputs(1114) <= not b;
    layer3_outputs(1115) <= a;
    layer3_outputs(1116) <= not (a and b);
    layer3_outputs(1117) <= a;
    layer3_outputs(1118) <= not b;
    layer3_outputs(1119) <= a;
    layer3_outputs(1120) <= b;
    layer3_outputs(1121) <= not b;
    layer3_outputs(1122) <= b;
    layer3_outputs(1123) <= not (a or b);
    layer3_outputs(1124) <= a and b;
    layer3_outputs(1125) <= not a;
    layer3_outputs(1126) <= not (a xor b);
    layer3_outputs(1127) <= a and not b;
    layer3_outputs(1128) <= not (a xor b);
    layer3_outputs(1129) <= not (a or b);
    layer3_outputs(1130) <= not a;
    layer3_outputs(1131) <= not (a or b);
    layer3_outputs(1132) <= not a;
    layer3_outputs(1133) <= not b;
    layer3_outputs(1134) <= b;
    layer3_outputs(1135) <= a;
    layer3_outputs(1136) <= not b;
    layer3_outputs(1137) <= b;
    layer3_outputs(1138) <= not a;
    layer3_outputs(1139) <= b;
    layer3_outputs(1140) <= not a;
    layer3_outputs(1141) <= not a or b;
    layer3_outputs(1142) <= not a;
    layer3_outputs(1143) <= a and b;
    layer3_outputs(1144) <= a;
    layer3_outputs(1145) <= not b or a;
    layer3_outputs(1146) <= a xor b;
    layer3_outputs(1147) <= 1'b1;
    layer3_outputs(1148) <= a;
    layer3_outputs(1149) <= not a or b;
    layer3_outputs(1150) <= not a;
    layer3_outputs(1151) <= not (a and b);
    layer3_outputs(1152) <= a or b;
    layer3_outputs(1153) <= not (a or b);
    layer3_outputs(1154) <= a;
    layer3_outputs(1155) <= not (a and b);
    layer3_outputs(1156) <= b;
    layer3_outputs(1157) <= a and not b;
    layer3_outputs(1158) <= not a;
    layer3_outputs(1159) <= b and not a;
    layer3_outputs(1160) <= a or b;
    layer3_outputs(1161) <= b and not a;
    layer3_outputs(1162) <= not (a and b);
    layer3_outputs(1163) <= a xor b;
    layer3_outputs(1164) <= a or b;
    layer3_outputs(1165) <= b;
    layer3_outputs(1166) <= a and not b;
    layer3_outputs(1167) <= a;
    layer3_outputs(1168) <= a or b;
    layer3_outputs(1169) <= a or b;
    layer3_outputs(1170) <= a;
    layer3_outputs(1171) <= a;
    layer3_outputs(1172) <= a;
    layer3_outputs(1173) <= not b;
    layer3_outputs(1174) <= not (a xor b);
    layer3_outputs(1175) <= not a;
    layer3_outputs(1176) <= not a or b;
    layer3_outputs(1177) <= not a;
    layer3_outputs(1178) <= a and not b;
    layer3_outputs(1179) <= a and b;
    layer3_outputs(1180) <= not (a xor b);
    layer3_outputs(1181) <= not (a and b);
    layer3_outputs(1182) <= b;
    layer3_outputs(1183) <= not b or a;
    layer3_outputs(1184) <= a xor b;
    layer3_outputs(1185) <= a and not b;
    layer3_outputs(1186) <= b and not a;
    layer3_outputs(1187) <= not b;
    layer3_outputs(1188) <= a and not b;
    layer3_outputs(1189) <= not b or a;
    layer3_outputs(1190) <= not a;
    layer3_outputs(1191) <= b and not a;
    layer3_outputs(1192) <= not b;
    layer3_outputs(1193) <= not a;
    layer3_outputs(1194) <= a;
    layer3_outputs(1195) <= not a;
    layer3_outputs(1196) <= not (a xor b);
    layer3_outputs(1197) <= a and not b;
    layer3_outputs(1198) <= not b;
    layer3_outputs(1199) <= a;
    layer3_outputs(1200) <= not b or a;
    layer3_outputs(1201) <= a and b;
    layer3_outputs(1202) <= not b or a;
    layer3_outputs(1203) <= a;
    layer3_outputs(1204) <= not b;
    layer3_outputs(1205) <= not b;
    layer3_outputs(1206) <= b and not a;
    layer3_outputs(1207) <= b;
    layer3_outputs(1208) <= a;
    layer3_outputs(1209) <= a and not b;
    layer3_outputs(1210) <= not (a or b);
    layer3_outputs(1211) <= b;
    layer3_outputs(1212) <= not a;
    layer3_outputs(1213) <= not a;
    layer3_outputs(1214) <= a and not b;
    layer3_outputs(1215) <= a and not b;
    layer3_outputs(1216) <= not b;
    layer3_outputs(1217) <= a xor b;
    layer3_outputs(1218) <= a;
    layer3_outputs(1219) <= a;
    layer3_outputs(1220) <= not b or a;
    layer3_outputs(1221) <= b;
    layer3_outputs(1222) <= b and not a;
    layer3_outputs(1223) <= not (a xor b);
    layer3_outputs(1224) <= a or b;
    layer3_outputs(1225) <= not (a xor b);
    layer3_outputs(1226) <= b;
    layer3_outputs(1227) <= not b;
    layer3_outputs(1228) <= not (a xor b);
    layer3_outputs(1229) <= a and b;
    layer3_outputs(1230) <= not (a or b);
    layer3_outputs(1231) <= not b;
    layer3_outputs(1232) <= b and not a;
    layer3_outputs(1233) <= not a;
    layer3_outputs(1234) <= not (a xor b);
    layer3_outputs(1235) <= not a;
    layer3_outputs(1236) <= a;
    layer3_outputs(1237) <= not a;
    layer3_outputs(1238) <= not b;
    layer3_outputs(1239) <= not a;
    layer3_outputs(1240) <= not b;
    layer3_outputs(1241) <= a and b;
    layer3_outputs(1242) <= not a;
    layer3_outputs(1243) <= b;
    layer3_outputs(1244) <= a;
    layer3_outputs(1245) <= not b or a;
    layer3_outputs(1246) <= not a or b;
    layer3_outputs(1247) <= a and b;
    layer3_outputs(1248) <= not b or a;
    layer3_outputs(1249) <= not b;
    layer3_outputs(1250) <= not a or b;
    layer3_outputs(1251) <= a or b;
    layer3_outputs(1252) <= not (a or b);
    layer3_outputs(1253) <= not a;
    layer3_outputs(1254) <= not b or a;
    layer3_outputs(1255) <= a and b;
    layer3_outputs(1256) <= a and b;
    layer3_outputs(1257) <= not a or b;
    layer3_outputs(1258) <= not b or a;
    layer3_outputs(1259) <= not b or a;
    layer3_outputs(1260) <= not a;
    layer3_outputs(1261) <= a;
    layer3_outputs(1262) <= not a or b;
    layer3_outputs(1263) <= b;
    layer3_outputs(1264) <= b;
    layer3_outputs(1265) <= not b or a;
    layer3_outputs(1266) <= a and not b;
    layer3_outputs(1267) <= b and not a;
    layer3_outputs(1268) <= not b;
    layer3_outputs(1269) <= not (a and b);
    layer3_outputs(1270) <= not (a xor b);
    layer3_outputs(1271) <= not b or a;
    layer3_outputs(1272) <= a xor b;
    layer3_outputs(1273) <= a and not b;
    layer3_outputs(1274) <= 1'b1;
    layer3_outputs(1275) <= not a or b;
    layer3_outputs(1276) <= a;
    layer3_outputs(1277) <= not a or b;
    layer3_outputs(1278) <= b;
    layer3_outputs(1279) <= not a;
    layer3_outputs(1280) <= not b;
    layer3_outputs(1281) <= not a;
    layer3_outputs(1282) <= b;
    layer3_outputs(1283) <= not a or b;
    layer3_outputs(1284) <= not (a xor b);
    layer3_outputs(1285) <= not b or a;
    layer3_outputs(1286) <= a or b;
    layer3_outputs(1287) <= a xor b;
    layer3_outputs(1288) <= a;
    layer3_outputs(1289) <= a and b;
    layer3_outputs(1290) <= not (a xor b);
    layer3_outputs(1291) <= not (a xor b);
    layer3_outputs(1292) <= not a;
    layer3_outputs(1293) <= a;
    layer3_outputs(1294) <= not (a or b);
    layer3_outputs(1295) <= not b;
    layer3_outputs(1296) <= not (a or b);
    layer3_outputs(1297) <= a and not b;
    layer3_outputs(1298) <= not (a or b);
    layer3_outputs(1299) <= not a or b;
    layer3_outputs(1300) <= not b;
    layer3_outputs(1301) <= not (a or b);
    layer3_outputs(1302) <= not b;
    layer3_outputs(1303) <= a and b;
    layer3_outputs(1304) <= not a;
    layer3_outputs(1305) <= not (a xor b);
    layer3_outputs(1306) <= not a;
    layer3_outputs(1307) <= b;
    layer3_outputs(1308) <= not b;
    layer3_outputs(1309) <= not (a or b);
    layer3_outputs(1310) <= a;
    layer3_outputs(1311) <= not b;
    layer3_outputs(1312) <= not a;
    layer3_outputs(1313) <= not a;
    layer3_outputs(1314) <= b;
    layer3_outputs(1315) <= a xor b;
    layer3_outputs(1316) <= a xor b;
    layer3_outputs(1317) <= 1'b1;
    layer3_outputs(1318) <= not b or a;
    layer3_outputs(1319) <= a and b;
    layer3_outputs(1320) <= not a or b;
    layer3_outputs(1321) <= not a or b;
    layer3_outputs(1322) <= not b;
    layer3_outputs(1323) <= not b or a;
    layer3_outputs(1324) <= not a;
    layer3_outputs(1325) <= b and not a;
    layer3_outputs(1326) <= a;
    layer3_outputs(1327) <= a or b;
    layer3_outputs(1328) <= not b;
    layer3_outputs(1329) <= not a or b;
    layer3_outputs(1330) <= b and not a;
    layer3_outputs(1331) <= b;
    layer3_outputs(1332) <= a;
    layer3_outputs(1333) <= not a;
    layer3_outputs(1334) <= not b;
    layer3_outputs(1335) <= not b;
    layer3_outputs(1336) <= not b;
    layer3_outputs(1337) <= a and b;
    layer3_outputs(1338) <= b;
    layer3_outputs(1339) <= not a;
    layer3_outputs(1340) <= a and not b;
    layer3_outputs(1341) <= a or b;
    layer3_outputs(1342) <= not a;
    layer3_outputs(1343) <= not a;
    layer3_outputs(1344) <= not a or b;
    layer3_outputs(1345) <= not b;
    layer3_outputs(1346) <= a xor b;
    layer3_outputs(1347) <= not b;
    layer3_outputs(1348) <= a;
    layer3_outputs(1349) <= a;
    layer3_outputs(1350) <= not a;
    layer3_outputs(1351) <= a or b;
    layer3_outputs(1352) <= b;
    layer3_outputs(1353) <= a and not b;
    layer3_outputs(1354) <= a xor b;
    layer3_outputs(1355) <= a;
    layer3_outputs(1356) <= not a or b;
    layer3_outputs(1357) <= not a or b;
    layer3_outputs(1358) <= b;
    layer3_outputs(1359) <= not b or a;
    layer3_outputs(1360) <= a xor b;
    layer3_outputs(1361) <= a;
    layer3_outputs(1362) <= not (a xor b);
    layer3_outputs(1363) <= b;
    layer3_outputs(1364) <= a and not b;
    layer3_outputs(1365) <= not (a xor b);
    layer3_outputs(1366) <= b and not a;
    layer3_outputs(1367) <= a;
    layer3_outputs(1368) <= not (a xor b);
    layer3_outputs(1369) <= not b;
    layer3_outputs(1370) <= b;
    layer3_outputs(1371) <= b;
    layer3_outputs(1372) <= not a;
    layer3_outputs(1373) <= a or b;
    layer3_outputs(1374) <= not (a xor b);
    layer3_outputs(1375) <= not a or b;
    layer3_outputs(1376) <= not b or a;
    layer3_outputs(1377) <= b and not a;
    layer3_outputs(1378) <= a or b;
    layer3_outputs(1379) <= not b;
    layer3_outputs(1380) <= a;
    layer3_outputs(1381) <= not (a xor b);
    layer3_outputs(1382) <= 1'b1;
    layer3_outputs(1383) <= b and not a;
    layer3_outputs(1384) <= a and not b;
    layer3_outputs(1385) <= not (a or b);
    layer3_outputs(1386) <= not a or b;
    layer3_outputs(1387) <= not (a or b);
    layer3_outputs(1388) <= a xor b;
    layer3_outputs(1389) <= not b;
    layer3_outputs(1390) <= a and b;
    layer3_outputs(1391) <= not b;
    layer3_outputs(1392) <= not b;
    layer3_outputs(1393) <= not (a xor b);
    layer3_outputs(1394) <= not b or a;
    layer3_outputs(1395) <= not a or b;
    layer3_outputs(1396) <= not a;
    layer3_outputs(1397) <= b;
    layer3_outputs(1398) <= b;
    layer3_outputs(1399) <= 1'b0;
    layer3_outputs(1400) <= b;
    layer3_outputs(1401) <= not (a xor b);
    layer3_outputs(1402) <= a and b;
    layer3_outputs(1403) <= a xor b;
    layer3_outputs(1404) <= a xor b;
    layer3_outputs(1405) <= not b or a;
    layer3_outputs(1406) <= a xor b;
    layer3_outputs(1407) <= not (a and b);
    layer3_outputs(1408) <= not a or b;
    layer3_outputs(1409) <= a xor b;
    layer3_outputs(1410) <= a or b;
    layer3_outputs(1411) <= b;
    layer3_outputs(1412) <= a;
    layer3_outputs(1413) <= not a;
    layer3_outputs(1414) <= a;
    layer3_outputs(1415) <= not (a xor b);
    layer3_outputs(1416) <= not b or a;
    layer3_outputs(1417) <= not a;
    layer3_outputs(1418) <= not (a or b);
    layer3_outputs(1419) <= b and not a;
    layer3_outputs(1420) <= a and b;
    layer3_outputs(1421) <= a;
    layer3_outputs(1422) <= b;
    layer3_outputs(1423) <= not a or b;
    layer3_outputs(1424) <= a or b;
    layer3_outputs(1425) <= b;
    layer3_outputs(1426) <= 1'b1;
    layer3_outputs(1427) <= a;
    layer3_outputs(1428) <= a;
    layer3_outputs(1429) <= b;
    layer3_outputs(1430) <= a or b;
    layer3_outputs(1431) <= b;
    layer3_outputs(1432) <= a and not b;
    layer3_outputs(1433) <= not a or b;
    layer3_outputs(1434) <= a and not b;
    layer3_outputs(1435) <= not (a xor b);
    layer3_outputs(1436) <= b;
    layer3_outputs(1437) <= b;
    layer3_outputs(1438) <= a;
    layer3_outputs(1439) <= not b;
    layer3_outputs(1440) <= not (a xor b);
    layer3_outputs(1441) <= not (a xor b);
    layer3_outputs(1442) <= not b or a;
    layer3_outputs(1443) <= a and not b;
    layer3_outputs(1444) <= a;
    layer3_outputs(1445) <= not (a and b);
    layer3_outputs(1446) <= b and not a;
    layer3_outputs(1447) <= a;
    layer3_outputs(1448) <= not (a and b);
    layer3_outputs(1449) <= not b;
    layer3_outputs(1450) <= not b or a;
    layer3_outputs(1451) <= not a or b;
    layer3_outputs(1452) <= not (a or b);
    layer3_outputs(1453) <= not (a xor b);
    layer3_outputs(1454) <= not (a xor b);
    layer3_outputs(1455) <= not (a or b);
    layer3_outputs(1456) <= b and not a;
    layer3_outputs(1457) <= a and not b;
    layer3_outputs(1458) <= not (a or b);
    layer3_outputs(1459) <= not (a or b);
    layer3_outputs(1460) <= a and b;
    layer3_outputs(1461) <= a and not b;
    layer3_outputs(1462) <= b and not a;
    layer3_outputs(1463) <= a or b;
    layer3_outputs(1464) <= not (a or b);
    layer3_outputs(1465) <= b;
    layer3_outputs(1466) <= not a;
    layer3_outputs(1467) <= a and b;
    layer3_outputs(1468) <= not a or b;
    layer3_outputs(1469) <= a and not b;
    layer3_outputs(1470) <= a;
    layer3_outputs(1471) <= a or b;
    layer3_outputs(1472) <= a and b;
    layer3_outputs(1473) <= 1'b0;
    layer3_outputs(1474) <= a or b;
    layer3_outputs(1475) <= not a;
    layer3_outputs(1476) <= b and not a;
    layer3_outputs(1477) <= a;
    layer3_outputs(1478) <= a;
    layer3_outputs(1479) <= b and not a;
    layer3_outputs(1480) <= not b or a;
    layer3_outputs(1481) <= b;
    layer3_outputs(1482) <= not b;
    layer3_outputs(1483) <= b;
    layer3_outputs(1484) <= not b;
    layer3_outputs(1485) <= b and not a;
    layer3_outputs(1486) <= b;
    layer3_outputs(1487) <= not b;
    layer3_outputs(1488) <= not (a xor b);
    layer3_outputs(1489) <= not a or b;
    layer3_outputs(1490) <= b;
    layer3_outputs(1491) <= b;
    layer3_outputs(1492) <= a and b;
    layer3_outputs(1493) <= a and not b;
    layer3_outputs(1494) <= not (a and b);
    layer3_outputs(1495) <= not a or b;
    layer3_outputs(1496) <= not a;
    layer3_outputs(1497) <= a or b;
    layer3_outputs(1498) <= b;
    layer3_outputs(1499) <= b;
    layer3_outputs(1500) <= not (a and b);
    layer3_outputs(1501) <= not b;
    layer3_outputs(1502) <= b;
    layer3_outputs(1503) <= a;
    layer3_outputs(1504) <= not (a and b);
    layer3_outputs(1505) <= not (a or b);
    layer3_outputs(1506) <= not b or a;
    layer3_outputs(1507) <= not a or b;
    layer3_outputs(1508) <= b;
    layer3_outputs(1509) <= a;
    layer3_outputs(1510) <= a;
    layer3_outputs(1511) <= a and not b;
    layer3_outputs(1512) <= a and not b;
    layer3_outputs(1513) <= a and b;
    layer3_outputs(1514) <= not a or b;
    layer3_outputs(1515) <= not a;
    layer3_outputs(1516) <= not (a or b);
    layer3_outputs(1517) <= not (a xor b);
    layer3_outputs(1518) <= a or b;
    layer3_outputs(1519) <= a and not b;
    layer3_outputs(1520) <= not (a and b);
    layer3_outputs(1521) <= not a or b;
    layer3_outputs(1522) <= a xor b;
    layer3_outputs(1523) <= b and not a;
    layer3_outputs(1524) <= b and not a;
    layer3_outputs(1525) <= not a;
    layer3_outputs(1526) <= not (a and b);
    layer3_outputs(1527) <= a;
    layer3_outputs(1528) <= b and not a;
    layer3_outputs(1529) <= not (a or b);
    layer3_outputs(1530) <= not b;
    layer3_outputs(1531) <= not (a or b);
    layer3_outputs(1532) <= b;
    layer3_outputs(1533) <= b;
    layer3_outputs(1534) <= not (a xor b);
    layer3_outputs(1535) <= a and b;
    layer3_outputs(1536) <= not b;
    layer3_outputs(1537) <= not a or b;
    layer3_outputs(1538) <= b;
    layer3_outputs(1539) <= a or b;
    layer3_outputs(1540) <= not a or b;
    layer3_outputs(1541) <= 1'b0;
    layer3_outputs(1542) <= a xor b;
    layer3_outputs(1543) <= not b or a;
    layer3_outputs(1544) <= not b;
    layer3_outputs(1545) <= b;
    layer3_outputs(1546) <= b and not a;
    layer3_outputs(1547) <= not (a and b);
    layer3_outputs(1548) <= b;
    layer3_outputs(1549) <= a and b;
    layer3_outputs(1550) <= not a;
    layer3_outputs(1551) <= b;
    layer3_outputs(1552) <= not b or a;
    layer3_outputs(1553) <= a or b;
    layer3_outputs(1554) <= a xor b;
    layer3_outputs(1555) <= a and not b;
    layer3_outputs(1556) <= b;
    layer3_outputs(1557) <= b and not a;
    layer3_outputs(1558) <= b and not a;
    layer3_outputs(1559) <= not a;
    layer3_outputs(1560) <= not a;
    layer3_outputs(1561) <= not b;
    layer3_outputs(1562) <= b and not a;
    layer3_outputs(1563) <= not (a xor b);
    layer3_outputs(1564) <= b;
    layer3_outputs(1565) <= not b or a;
    layer3_outputs(1566) <= not a or b;
    layer3_outputs(1567) <= b and not a;
    layer3_outputs(1568) <= 1'b1;
    layer3_outputs(1569) <= not b;
    layer3_outputs(1570) <= not a;
    layer3_outputs(1571) <= not b or a;
    layer3_outputs(1572) <= a and not b;
    layer3_outputs(1573) <= a and b;
    layer3_outputs(1574) <= a or b;
    layer3_outputs(1575) <= not b;
    layer3_outputs(1576) <= b and not a;
    layer3_outputs(1577) <= a or b;
    layer3_outputs(1578) <= b;
    layer3_outputs(1579) <= not (a and b);
    layer3_outputs(1580) <= a xor b;
    layer3_outputs(1581) <= not a or b;
    layer3_outputs(1582) <= a and b;
    layer3_outputs(1583) <= not b;
    layer3_outputs(1584) <= b;
    layer3_outputs(1585) <= not a or b;
    layer3_outputs(1586) <= b;
    layer3_outputs(1587) <= b and not a;
    layer3_outputs(1588) <= not b;
    layer3_outputs(1589) <= b;
    layer3_outputs(1590) <= a or b;
    layer3_outputs(1591) <= a and b;
    layer3_outputs(1592) <= not a;
    layer3_outputs(1593) <= not a or b;
    layer3_outputs(1594) <= not b or a;
    layer3_outputs(1595) <= a;
    layer3_outputs(1596) <= b;
    layer3_outputs(1597) <= a xor b;
    layer3_outputs(1598) <= not a or b;
    layer3_outputs(1599) <= not a;
    layer3_outputs(1600) <= b and not a;
    layer3_outputs(1601) <= not (a xor b);
    layer3_outputs(1602) <= a xor b;
    layer3_outputs(1603) <= not b or a;
    layer3_outputs(1604) <= not a;
    layer3_outputs(1605) <= b;
    layer3_outputs(1606) <= not b;
    layer3_outputs(1607) <= b;
    layer3_outputs(1608) <= not b;
    layer3_outputs(1609) <= not (a or b);
    layer3_outputs(1610) <= a;
    layer3_outputs(1611) <= not (a and b);
    layer3_outputs(1612) <= not b;
    layer3_outputs(1613) <= a and b;
    layer3_outputs(1614) <= not a;
    layer3_outputs(1615) <= b;
    layer3_outputs(1616) <= not (a xor b);
    layer3_outputs(1617) <= not b or a;
    layer3_outputs(1618) <= not (a or b);
    layer3_outputs(1619) <= a and not b;
    layer3_outputs(1620) <= not b or a;
    layer3_outputs(1621) <= a;
    layer3_outputs(1622) <= b;
    layer3_outputs(1623) <= a;
    layer3_outputs(1624) <= not (a or b);
    layer3_outputs(1625) <= not (a xor b);
    layer3_outputs(1626) <= a and not b;
    layer3_outputs(1627) <= b;
    layer3_outputs(1628) <= not (a or b);
    layer3_outputs(1629) <= a xor b;
    layer3_outputs(1630) <= a;
    layer3_outputs(1631) <= b;
    layer3_outputs(1632) <= not a;
    layer3_outputs(1633) <= not b or a;
    layer3_outputs(1634) <= not (a and b);
    layer3_outputs(1635) <= b and not a;
    layer3_outputs(1636) <= a xor b;
    layer3_outputs(1637) <= b;
    layer3_outputs(1638) <= a;
    layer3_outputs(1639) <= b;
    layer3_outputs(1640) <= a and not b;
    layer3_outputs(1641) <= not b or a;
    layer3_outputs(1642) <= not a;
    layer3_outputs(1643) <= a;
    layer3_outputs(1644) <= not (a or b);
    layer3_outputs(1645) <= 1'b0;
    layer3_outputs(1646) <= not a;
    layer3_outputs(1647) <= not (a xor b);
    layer3_outputs(1648) <= not (a or b);
    layer3_outputs(1649) <= not (a and b);
    layer3_outputs(1650) <= a;
    layer3_outputs(1651) <= a;
    layer3_outputs(1652) <= not (a xor b);
    layer3_outputs(1653) <= a and b;
    layer3_outputs(1654) <= not a or b;
    layer3_outputs(1655) <= not (a and b);
    layer3_outputs(1656) <= b and not a;
    layer3_outputs(1657) <= not b or a;
    layer3_outputs(1658) <= not (a xor b);
    layer3_outputs(1659) <= b;
    layer3_outputs(1660) <= not a;
    layer3_outputs(1661) <= not b or a;
    layer3_outputs(1662) <= b and not a;
    layer3_outputs(1663) <= a or b;
    layer3_outputs(1664) <= not b;
    layer3_outputs(1665) <= b;
    layer3_outputs(1666) <= b;
    layer3_outputs(1667) <= a and b;
    layer3_outputs(1668) <= not (a and b);
    layer3_outputs(1669) <= not (a and b);
    layer3_outputs(1670) <= 1'b0;
    layer3_outputs(1671) <= not a;
    layer3_outputs(1672) <= a or b;
    layer3_outputs(1673) <= not a;
    layer3_outputs(1674) <= a;
    layer3_outputs(1675) <= not (a or b);
    layer3_outputs(1676) <= b;
    layer3_outputs(1677) <= a;
    layer3_outputs(1678) <= b;
    layer3_outputs(1679) <= not b;
    layer3_outputs(1680) <= not (a or b);
    layer3_outputs(1681) <= not b;
    layer3_outputs(1682) <= b and not a;
    layer3_outputs(1683) <= not a;
    layer3_outputs(1684) <= a and not b;
    layer3_outputs(1685) <= a or b;
    layer3_outputs(1686) <= not a;
    layer3_outputs(1687) <= b;
    layer3_outputs(1688) <= a and not b;
    layer3_outputs(1689) <= not (a and b);
    layer3_outputs(1690) <= not b or a;
    layer3_outputs(1691) <= not a;
    layer3_outputs(1692) <= not a;
    layer3_outputs(1693) <= not a;
    layer3_outputs(1694) <= not a;
    layer3_outputs(1695) <= not (a and b);
    layer3_outputs(1696) <= not (a and b);
    layer3_outputs(1697) <= b;
    layer3_outputs(1698) <= b;
    layer3_outputs(1699) <= not b or a;
    layer3_outputs(1700) <= not (a xor b);
    layer3_outputs(1701) <= not (a xor b);
    layer3_outputs(1702) <= b;
    layer3_outputs(1703) <= a or b;
    layer3_outputs(1704) <= a and not b;
    layer3_outputs(1705) <= a and b;
    layer3_outputs(1706) <= a xor b;
    layer3_outputs(1707) <= a xor b;
    layer3_outputs(1708) <= not a;
    layer3_outputs(1709) <= a;
    layer3_outputs(1710) <= b;
    layer3_outputs(1711) <= a and b;
    layer3_outputs(1712) <= b;
    layer3_outputs(1713) <= a or b;
    layer3_outputs(1714) <= b and not a;
    layer3_outputs(1715) <= not a;
    layer3_outputs(1716) <= not b;
    layer3_outputs(1717) <= not (a or b);
    layer3_outputs(1718) <= not b;
    layer3_outputs(1719) <= a;
    layer3_outputs(1720) <= not (a and b);
    layer3_outputs(1721) <= b and not a;
    layer3_outputs(1722) <= b;
    layer3_outputs(1723) <= a;
    layer3_outputs(1724) <= a and not b;
    layer3_outputs(1725) <= a;
    layer3_outputs(1726) <= not b;
    layer3_outputs(1727) <= b;
    layer3_outputs(1728) <= not a;
    layer3_outputs(1729) <= a;
    layer3_outputs(1730) <= not b or a;
    layer3_outputs(1731) <= 1'b1;
    layer3_outputs(1732) <= b and not a;
    layer3_outputs(1733) <= a;
    layer3_outputs(1734) <= not a or b;
    layer3_outputs(1735) <= b;
    layer3_outputs(1736) <= not a or b;
    layer3_outputs(1737) <= not b or a;
    layer3_outputs(1738) <= not (a xor b);
    layer3_outputs(1739) <= b;
    layer3_outputs(1740) <= not b or a;
    layer3_outputs(1741) <= 1'b0;
    layer3_outputs(1742) <= not (a and b);
    layer3_outputs(1743) <= 1'b1;
    layer3_outputs(1744) <= 1'b1;
    layer3_outputs(1745) <= not a or b;
    layer3_outputs(1746) <= a xor b;
    layer3_outputs(1747) <= not b;
    layer3_outputs(1748) <= a;
    layer3_outputs(1749) <= b;
    layer3_outputs(1750) <= not a or b;
    layer3_outputs(1751) <= b;
    layer3_outputs(1752) <= not (a xor b);
    layer3_outputs(1753) <= a and b;
    layer3_outputs(1754) <= not b;
    layer3_outputs(1755) <= not (a xor b);
    layer3_outputs(1756) <= not a;
    layer3_outputs(1757) <= not b;
    layer3_outputs(1758) <= a xor b;
    layer3_outputs(1759) <= not b;
    layer3_outputs(1760) <= 1'b0;
    layer3_outputs(1761) <= a;
    layer3_outputs(1762) <= a and not b;
    layer3_outputs(1763) <= not a or b;
    layer3_outputs(1764) <= not (a xor b);
    layer3_outputs(1765) <= not a;
    layer3_outputs(1766) <= a and not b;
    layer3_outputs(1767) <= not (a or b);
    layer3_outputs(1768) <= a and b;
    layer3_outputs(1769) <= b;
    layer3_outputs(1770) <= not (a xor b);
    layer3_outputs(1771) <= a or b;
    layer3_outputs(1772) <= not b or a;
    layer3_outputs(1773) <= a xor b;
    layer3_outputs(1774) <= not b or a;
    layer3_outputs(1775) <= not b;
    layer3_outputs(1776) <= not a;
    layer3_outputs(1777) <= a and b;
    layer3_outputs(1778) <= a and not b;
    layer3_outputs(1779) <= not b;
    layer3_outputs(1780) <= a and not b;
    layer3_outputs(1781) <= not (a or b);
    layer3_outputs(1782) <= b;
    layer3_outputs(1783) <= not (a xor b);
    layer3_outputs(1784) <= b and not a;
    layer3_outputs(1785) <= b and not a;
    layer3_outputs(1786) <= 1'b1;
    layer3_outputs(1787) <= not a;
    layer3_outputs(1788) <= b and not a;
    layer3_outputs(1789) <= a xor b;
    layer3_outputs(1790) <= b;
    layer3_outputs(1791) <= not (a and b);
    layer3_outputs(1792) <= not a or b;
    layer3_outputs(1793) <= not b;
    layer3_outputs(1794) <= not (a xor b);
    layer3_outputs(1795) <= a;
    layer3_outputs(1796) <= not b;
    layer3_outputs(1797) <= a xor b;
    layer3_outputs(1798) <= a and not b;
    layer3_outputs(1799) <= a or b;
    layer3_outputs(1800) <= not a;
    layer3_outputs(1801) <= a or b;
    layer3_outputs(1802) <= not a;
    layer3_outputs(1803) <= not b or a;
    layer3_outputs(1804) <= b and not a;
    layer3_outputs(1805) <= a and b;
    layer3_outputs(1806) <= not b;
    layer3_outputs(1807) <= a and b;
    layer3_outputs(1808) <= not (a xor b);
    layer3_outputs(1809) <= a;
    layer3_outputs(1810) <= b;
    layer3_outputs(1811) <= not b;
    layer3_outputs(1812) <= not b;
    layer3_outputs(1813) <= b and not a;
    layer3_outputs(1814) <= a xor b;
    layer3_outputs(1815) <= not (a xor b);
    layer3_outputs(1816) <= a and not b;
    layer3_outputs(1817) <= b and not a;
    layer3_outputs(1818) <= a xor b;
    layer3_outputs(1819) <= b;
    layer3_outputs(1820) <= not b;
    layer3_outputs(1821) <= a xor b;
    layer3_outputs(1822) <= a;
    layer3_outputs(1823) <= not b;
    layer3_outputs(1824) <= not a;
    layer3_outputs(1825) <= not a;
    layer3_outputs(1826) <= a and not b;
    layer3_outputs(1827) <= a;
    layer3_outputs(1828) <= not b or a;
    layer3_outputs(1829) <= b;
    layer3_outputs(1830) <= a and b;
    layer3_outputs(1831) <= a xor b;
    layer3_outputs(1832) <= not b or a;
    layer3_outputs(1833) <= not (a xor b);
    layer3_outputs(1834) <= not b or a;
    layer3_outputs(1835) <= a and not b;
    layer3_outputs(1836) <= not (a or b);
    layer3_outputs(1837) <= a and not b;
    layer3_outputs(1838) <= not (a xor b);
    layer3_outputs(1839) <= not b;
    layer3_outputs(1840) <= b;
    layer3_outputs(1841) <= a;
    layer3_outputs(1842) <= a and not b;
    layer3_outputs(1843) <= not (a and b);
    layer3_outputs(1844) <= b and not a;
    layer3_outputs(1845) <= not a or b;
    layer3_outputs(1846) <= not b;
    layer3_outputs(1847) <= b;
    layer3_outputs(1848) <= not a;
    layer3_outputs(1849) <= a and b;
    layer3_outputs(1850) <= a xor b;
    layer3_outputs(1851) <= a and not b;
    layer3_outputs(1852) <= b;
    layer3_outputs(1853) <= not b;
    layer3_outputs(1854) <= not (a xor b);
    layer3_outputs(1855) <= a xor b;
    layer3_outputs(1856) <= b and not a;
    layer3_outputs(1857) <= a xor b;
    layer3_outputs(1858) <= not (a or b);
    layer3_outputs(1859) <= not b or a;
    layer3_outputs(1860) <= not b or a;
    layer3_outputs(1861) <= b and not a;
    layer3_outputs(1862) <= a;
    layer3_outputs(1863) <= 1'b0;
    layer3_outputs(1864) <= not (a and b);
    layer3_outputs(1865) <= a;
    layer3_outputs(1866) <= not a;
    layer3_outputs(1867) <= a and b;
    layer3_outputs(1868) <= not (a and b);
    layer3_outputs(1869) <= a xor b;
    layer3_outputs(1870) <= not a or b;
    layer3_outputs(1871) <= b and not a;
    layer3_outputs(1872) <= not a;
    layer3_outputs(1873) <= not a;
    layer3_outputs(1874) <= a;
    layer3_outputs(1875) <= not a or b;
    layer3_outputs(1876) <= not a;
    layer3_outputs(1877) <= a;
    layer3_outputs(1878) <= a or b;
    layer3_outputs(1879) <= not b;
    layer3_outputs(1880) <= not (a and b);
    layer3_outputs(1881) <= not (a or b);
    layer3_outputs(1882) <= not a;
    layer3_outputs(1883) <= not b;
    layer3_outputs(1884) <= not b;
    layer3_outputs(1885) <= a xor b;
    layer3_outputs(1886) <= not (a and b);
    layer3_outputs(1887) <= a xor b;
    layer3_outputs(1888) <= a or b;
    layer3_outputs(1889) <= not (a and b);
    layer3_outputs(1890) <= a or b;
    layer3_outputs(1891) <= b and not a;
    layer3_outputs(1892) <= not (a and b);
    layer3_outputs(1893) <= not (a and b);
    layer3_outputs(1894) <= b and not a;
    layer3_outputs(1895) <= a;
    layer3_outputs(1896) <= not a or b;
    layer3_outputs(1897) <= a and not b;
    layer3_outputs(1898) <= not b or a;
    layer3_outputs(1899) <= not a or b;
    layer3_outputs(1900) <= not (a xor b);
    layer3_outputs(1901) <= b;
    layer3_outputs(1902) <= not b;
    layer3_outputs(1903) <= b and not a;
    layer3_outputs(1904) <= b;
    layer3_outputs(1905) <= not b;
    layer3_outputs(1906) <= not b;
    layer3_outputs(1907) <= a and not b;
    layer3_outputs(1908) <= b;
    layer3_outputs(1909) <= not a or b;
    layer3_outputs(1910) <= a and not b;
    layer3_outputs(1911) <= not (a and b);
    layer3_outputs(1912) <= a and b;
    layer3_outputs(1913) <= not (a or b);
    layer3_outputs(1914) <= not a or b;
    layer3_outputs(1915) <= not b;
    layer3_outputs(1916) <= a xor b;
    layer3_outputs(1917) <= not a or b;
    layer3_outputs(1918) <= not b or a;
    layer3_outputs(1919) <= a;
    layer3_outputs(1920) <= not a or b;
    layer3_outputs(1921) <= not a or b;
    layer3_outputs(1922) <= not (a and b);
    layer3_outputs(1923) <= not (a xor b);
    layer3_outputs(1924) <= a;
    layer3_outputs(1925) <= b and not a;
    layer3_outputs(1926) <= 1'b0;
    layer3_outputs(1927) <= a xor b;
    layer3_outputs(1928) <= not (a or b);
    layer3_outputs(1929) <= not b or a;
    layer3_outputs(1930) <= not b;
    layer3_outputs(1931) <= not (a xor b);
    layer3_outputs(1932) <= not b or a;
    layer3_outputs(1933) <= not (a or b);
    layer3_outputs(1934) <= not b;
    layer3_outputs(1935) <= not b;
    layer3_outputs(1936) <= not a;
    layer3_outputs(1937) <= not (a or b);
    layer3_outputs(1938) <= b;
    layer3_outputs(1939) <= not b;
    layer3_outputs(1940) <= a xor b;
    layer3_outputs(1941) <= not (a xor b);
    layer3_outputs(1942) <= b;
    layer3_outputs(1943) <= b and not a;
    layer3_outputs(1944) <= a and not b;
    layer3_outputs(1945) <= not a or b;
    layer3_outputs(1946) <= a or b;
    layer3_outputs(1947) <= not (a and b);
    layer3_outputs(1948) <= b;
    layer3_outputs(1949) <= a xor b;
    layer3_outputs(1950) <= not a;
    layer3_outputs(1951) <= a and not b;
    layer3_outputs(1952) <= a and not b;
    layer3_outputs(1953) <= not b;
    layer3_outputs(1954) <= not (a and b);
    layer3_outputs(1955) <= not b or a;
    layer3_outputs(1956) <= not a;
    layer3_outputs(1957) <= not (a xor b);
    layer3_outputs(1958) <= not b;
    layer3_outputs(1959) <= not b;
    layer3_outputs(1960) <= a or b;
    layer3_outputs(1961) <= a;
    layer3_outputs(1962) <= a xor b;
    layer3_outputs(1963) <= 1'b1;
    layer3_outputs(1964) <= not (a and b);
    layer3_outputs(1965) <= not a or b;
    layer3_outputs(1966) <= not b;
    layer3_outputs(1967) <= 1'b1;
    layer3_outputs(1968) <= not b;
    layer3_outputs(1969) <= not b;
    layer3_outputs(1970) <= a or b;
    layer3_outputs(1971) <= a and not b;
    layer3_outputs(1972) <= b;
    layer3_outputs(1973) <= not b;
    layer3_outputs(1974) <= not a;
    layer3_outputs(1975) <= b;
    layer3_outputs(1976) <= a;
    layer3_outputs(1977) <= not a or b;
    layer3_outputs(1978) <= not b;
    layer3_outputs(1979) <= a and not b;
    layer3_outputs(1980) <= a xor b;
    layer3_outputs(1981) <= not b;
    layer3_outputs(1982) <= 1'b0;
    layer3_outputs(1983) <= a and not b;
    layer3_outputs(1984) <= b;
    layer3_outputs(1985) <= a;
    layer3_outputs(1986) <= b;
    layer3_outputs(1987) <= not b;
    layer3_outputs(1988) <= a and b;
    layer3_outputs(1989) <= a;
    layer3_outputs(1990) <= not b;
    layer3_outputs(1991) <= b;
    layer3_outputs(1992) <= not a;
    layer3_outputs(1993) <= b;
    layer3_outputs(1994) <= not b;
    layer3_outputs(1995) <= b;
    layer3_outputs(1996) <= not (a xor b);
    layer3_outputs(1997) <= a xor b;
    layer3_outputs(1998) <= not (a and b);
    layer3_outputs(1999) <= a;
    layer3_outputs(2000) <= not a or b;
    layer3_outputs(2001) <= not b;
    layer3_outputs(2002) <= a;
    layer3_outputs(2003) <= not b or a;
    layer3_outputs(2004) <= not a;
    layer3_outputs(2005) <= a;
    layer3_outputs(2006) <= a and not b;
    layer3_outputs(2007) <= 1'b0;
    layer3_outputs(2008) <= not (a or b);
    layer3_outputs(2009) <= a;
    layer3_outputs(2010) <= not b or a;
    layer3_outputs(2011) <= not a or b;
    layer3_outputs(2012) <= b;
    layer3_outputs(2013) <= a xor b;
    layer3_outputs(2014) <= a;
    layer3_outputs(2015) <= a or b;
    layer3_outputs(2016) <= a and not b;
    layer3_outputs(2017) <= not b;
    layer3_outputs(2018) <= not a;
    layer3_outputs(2019) <= a and not b;
    layer3_outputs(2020) <= b;
    layer3_outputs(2021) <= a xor b;
    layer3_outputs(2022) <= b;
    layer3_outputs(2023) <= not b;
    layer3_outputs(2024) <= a;
    layer3_outputs(2025) <= a xor b;
    layer3_outputs(2026) <= b;
    layer3_outputs(2027) <= b and not a;
    layer3_outputs(2028) <= not (a or b);
    layer3_outputs(2029) <= 1'b0;
    layer3_outputs(2030) <= b and not a;
    layer3_outputs(2031) <= a and not b;
    layer3_outputs(2032) <= not (a or b);
    layer3_outputs(2033) <= a xor b;
    layer3_outputs(2034) <= a or b;
    layer3_outputs(2035) <= not b;
    layer3_outputs(2036) <= not b or a;
    layer3_outputs(2037) <= a;
    layer3_outputs(2038) <= a or b;
    layer3_outputs(2039) <= not (a xor b);
    layer3_outputs(2040) <= a or b;
    layer3_outputs(2041) <= b and not a;
    layer3_outputs(2042) <= not a;
    layer3_outputs(2043) <= 1'b1;
    layer3_outputs(2044) <= not b;
    layer3_outputs(2045) <= not b;
    layer3_outputs(2046) <= not b or a;
    layer3_outputs(2047) <= b;
    layer3_outputs(2048) <= 1'b0;
    layer3_outputs(2049) <= b and not a;
    layer3_outputs(2050) <= not a or b;
    layer3_outputs(2051) <= a and b;
    layer3_outputs(2052) <= b and not a;
    layer3_outputs(2053) <= a;
    layer3_outputs(2054) <= a and not b;
    layer3_outputs(2055) <= not (a xor b);
    layer3_outputs(2056) <= not a;
    layer3_outputs(2057) <= not a;
    layer3_outputs(2058) <= not (a and b);
    layer3_outputs(2059) <= b;
    layer3_outputs(2060) <= not a or b;
    layer3_outputs(2061) <= not a or b;
    layer3_outputs(2062) <= not b;
    layer3_outputs(2063) <= not b or a;
    layer3_outputs(2064) <= b;
    layer3_outputs(2065) <= not a;
    layer3_outputs(2066) <= not (a xor b);
    layer3_outputs(2067) <= b;
    layer3_outputs(2068) <= not b;
    layer3_outputs(2069) <= not a;
    layer3_outputs(2070) <= b and not a;
    layer3_outputs(2071) <= a xor b;
    layer3_outputs(2072) <= not (a xor b);
    layer3_outputs(2073) <= not (a and b);
    layer3_outputs(2074) <= not (a xor b);
    layer3_outputs(2075) <= a or b;
    layer3_outputs(2076) <= not (a or b);
    layer3_outputs(2077) <= not (a and b);
    layer3_outputs(2078) <= not (a xor b);
    layer3_outputs(2079) <= not a or b;
    layer3_outputs(2080) <= not (a xor b);
    layer3_outputs(2081) <= b;
    layer3_outputs(2082) <= not b;
    layer3_outputs(2083) <= not b;
    layer3_outputs(2084) <= a xor b;
    layer3_outputs(2085) <= 1'b0;
    layer3_outputs(2086) <= b;
    layer3_outputs(2087) <= a xor b;
    layer3_outputs(2088) <= a xor b;
    layer3_outputs(2089) <= a xor b;
    layer3_outputs(2090) <= not b;
    layer3_outputs(2091) <= not (a or b);
    layer3_outputs(2092) <= not a;
    layer3_outputs(2093) <= not b;
    layer3_outputs(2094) <= not b;
    layer3_outputs(2095) <= not b or a;
    layer3_outputs(2096) <= b;
    layer3_outputs(2097) <= a;
    layer3_outputs(2098) <= not b;
    layer3_outputs(2099) <= not (a or b);
    layer3_outputs(2100) <= not a;
    layer3_outputs(2101) <= a or b;
    layer3_outputs(2102) <= not a;
    layer3_outputs(2103) <= not (a or b);
    layer3_outputs(2104) <= not (a or b);
    layer3_outputs(2105) <= a and not b;
    layer3_outputs(2106) <= a and not b;
    layer3_outputs(2107) <= b;
    layer3_outputs(2108) <= a xor b;
    layer3_outputs(2109) <= b;
    layer3_outputs(2110) <= a and b;
    layer3_outputs(2111) <= not (a xor b);
    layer3_outputs(2112) <= a and not b;
    layer3_outputs(2113) <= a or b;
    layer3_outputs(2114) <= b;
    layer3_outputs(2115) <= a;
    layer3_outputs(2116) <= a or b;
    layer3_outputs(2117) <= a;
    layer3_outputs(2118) <= not b;
    layer3_outputs(2119) <= not b;
    layer3_outputs(2120) <= not a;
    layer3_outputs(2121) <= not b;
    layer3_outputs(2122) <= a xor b;
    layer3_outputs(2123) <= not (a or b);
    layer3_outputs(2124) <= a;
    layer3_outputs(2125) <= a or b;
    layer3_outputs(2126) <= not b;
    layer3_outputs(2127) <= not a;
    layer3_outputs(2128) <= not (a and b);
    layer3_outputs(2129) <= a;
    layer3_outputs(2130) <= not b or a;
    layer3_outputs(2131) <= not a;
    layer3_outputs(2132) <= a and b;
    layer3_outputs(2133) <= a or b;
    layer3_outputs(2134) <= not (a or b);
    layer3_outputs(2135) <= not (a or b);
    layer3_outputs(2136) <= a and not b;
    layer3_outputs(2137) <= b and not a;
    layer3_outputs(2138) <= not (a or b);
    layer3_outputs(2139) <= not a or b;
    layer3_outputs(2140) <= a;
    layer3_outputs(2141) <= a xor b;
    layer3_outputs(2142) <= not b;
    layer3_outputs(2143) <= not (a or b);
    layer3_outputs(2144) <= b;
    layer3_outputs(2145) <= not a or b;
    layer3_outputs(2146) <= not a;
    layer3_outputs(2147) <= a;
    layer3_outputs(2148) <= a and b;
    layer3_outputs(2149) <= not (a or b);
    layer3_outputs(2150) <= not (a xor b);
    layer3_outputs(2151) <= not a;
    layer3_outputs(2152) <= b;
    layer3_outputs(2153) <= not (a or b);
    layer3_outputs(2154) <= not (a or b);
    layer3_outputs(2155) <= not (a or b);
    layer3_outputs(2156) <= not b;
    layer3_outputs(2157) <= not (a xor b);
    layer3_outputs(2158) <= a;
    layer3_outputs(2159) <= 1'b1;
    layer3_outputs(2160) <= not a;
    layer3_outputs(2161) <= a and b;
    layer3_outputs(2162) <= a xor b;
    layer3_outputs(2163) <= not (a xor b);
    layer3_outputs(2164) <= not a;
    layer3_outputs(2165) <= a or b;
    layer3_outputs(2166) <= not b or a;
    layer3_outputs(2167) <= not (a or b);
    layer3_outputs(2168) <= a xor b;
    layer3_outputs(2169) <= b;
    layer3_outputs(2170) <= not (a or b);
    layer3_outputs(2171) <= not a;
    layer3_outputs(2172) <= a;
    layer3_outputs(2173) <= not a;
    layer3_outputs(2174) <= a xor b;
    layer3_outputs(2175) <= b;
    layer3_outputs(2176) <= not (a xor b);
    layer3_outputs(2177) <= 1'b0;
    layer3_outputs(2178) <= not b or a;
    layer3_outputs(2179) <= not a;
    layer3_outputs(2180) <= not b;
    layer3_outputs(2181) <= a and not b;
    layer3_outputs(2182) <= not (a or b);
    layer3_outputs(2183) <= a and b;
    layer3_outputs(2184) <= not a;
    layer3_outputs(2185) <= a or b;
    layer3_outputs(2186) <= not (a or b);
    layer3_outputs(2187) <= not b or a;
    layer3_outputs(2188) <= a or b;
    layer3_outputs(2189) <= not a or b;
    layer3_outputs(2190) <= a and b;
    layer3_outputs(2191) <= b;
    layer3_outputs(2192) <= a xor b;
    layer3_outputs(2193) <= a or b;
    layer3_outputs(2194) <= not a;
    layer3_outputs(2195) <= not b or a;
    layer3_outputs(2196) <= b and not a;
    layer3_outputs(2197) <= a and not b;
    layer3_outputs(2198) <= not (a and b);
    layer3_outputs(2199) <= a and b;
    layer3_outputs(2200) <= a and not b;
    layer3_outputs(2201) <= b;
    layer3_outputs(2202) <= a xor b;
    layer3_outputs(2203) <= a;
    layer3_outputs(2204) <= b;
    layer3_outputs(2205) <= a;
    layer3_outputs(2206) <= not (a xor b);
    layer3_outputs(2207) <= not b or a;
    layer3_outputs(2208) <= not b;
    layer3_outputs(2209) <= a xor b;
    layer3_outputs(2210) <= a xor b;
    layer3_outputs(2211) <= a;
    layer3_outputs(2212) <= b;
    layer3_outputs(2213) <= 1'b1;
    layer3_outputs(2214) <= not b;
    layer3_outputs(2215) <= b;
    layer3_outputs(2216) <= not a;
    layer3_outputs(2217) <= a;
    layer3_outputs(2218) <= not b;
    layer3_outputs(2219) <= 1'b0;
    layer3_outputs(2220) <= not a;
    layer3_outputs(2221) <= a;
    layer3_outputs(2222) <= not (a xor b);
    layer3_outputs(2223) <= not a;
    layer3_outputs(2224) <= b;
    layer3_outputs(2225) <= not a;
    layer3_outputs(2226) <= b;
    layer3_outputs(2227) <= b;
    layer3_outputs(2228) <= a xor b;
    layer3_outputs(2229) <= b and not a;
    layer3_outputs(2230) <= 1'b0;
    layer3_outputs(2231) <= not (a or b);
    layer3_outputs(2232) <= not b;
    layer3_outputs(2233) <= b;
    layer3_outputs(2234) <= not b;
    layer3_outputs(2235) <= a and not b;
    layer3_outputs(2236) <= a xor b;
    layer3_outputs(2237) <= a;
    layer3_outputs(2238) <= not b or a;
    layer3_outputs(2239) <= a or b;
    layer3_outputs(2240) <= a;
    layer3_outputs(2241) <= a;
    layer3_outputs(2242) <= not a;
    layer3_outputs(2243) <= b and not a;
    layer3_outputs(2244) <= a and not b;
    layer3_outputs(2245) <= not a;
    layer3_outputs(2246) <= not a;
    layer3_outputs(2247) <= not (a and b);
    layer3_outputs(2248) <= not (a xor b);
    layer3_outputs(2249) <= a;
    layer3_outputs(2250) <= not a;
    layer3_outputs(2251) <= a or b;
    layer3_outputs(2252) <= not a;
    layer3_outputs(2253) <= not (a and b);
    layer3_outputs(2254) <= not (a and b);
    layer3_outputs(2255) <= not a;
    layer3_outputs(2256) <= a and not b;
    layer3_outputs(2257) <= not b;
    layer3_outputs(2258) <= not (a xor b);
    layer3_outputs(2259) <= not b;
    layer3_outputs(2260) <= not a or b;
    layer3_outputs(2261) <= a and not b;
    layer3_outputs(2262) <= not b;
    layer3_outputs(2263) <= not b;
    layer3_outputs(2264) <= b;
    layer3_outputs(2265) <= b;
    layer3_outputs(2266) <= a and not b;
    layer3_outputs(2267) <= not b;
    layer3_outputs(2268) <= a and not b;
    layer3_outputs(2269) <= not (a xor b);
    layer3_outputs(2270) <= not (a xor b);
    layer3_outputs(2271) <= a xor b;
    layer3_outputs(2272) <= not b;
    layer3_outputs(2273) <= 1'b1;
    layer3_outputs(2274) <= a and not b;
    layer3_outputs(2275) <= not b or a;
    layer3_outputs(2276) <= not (a or b);
    layer3_outputs(2277) <= not b;
    layer3_outputs(2278) <= a and not b;
    layer3_outputs(2279) <= b;
    layer3_outputs(2280) <= b;
    layer3_outputs(2281) <= 1'b0;
    layer3_outputs(2282) <= not a;
    layer3_outputs(2283) <= b;
    layer3_outputs(2284) <= not a;
    layer3_outputs(2285) <= not (a or b);
    layer3_outputs(2286) <= not b;
    layer3_outputs(2287) <= a or b;
    layer3_outputs(2288) <= a and not b;
    layer3_outputs(2289) <= b;
    layer3_outputs(2290) <= not b;
    layer3_outputs(2291) <= not b or a;
    layer3_outputs(2292) <= a;
    layer3_outputs(2293) <= a and not b;
    layer3_outputs(2294) <= a and not b;
    layer3_outputs(2295) <= not a;
    layer3_outputs(2296) <= not (a xor b);
    layer3_outputs(2297) <= not (a xor b);
    layer3_outputs(2298) <= a and b;
    layer3_outputs(2299) <= a;
    layer3_outputs(2300) <= not b or a;
    layer3_outputs(2301) <= not a;
    layer3_outputs(2302) <= not a;
    layer3_outputs(2303) <= not b or a;
    layer3_outputs(2304) <= not b or a;
    layer3_outputs(2305) <= not b;
    layer3_outputs(2306) <= not (a xor b);
    layer3_outputs(2307) <= b and not a;
    layer3_outputs(2308) <= not (a xor b);
    layer3_outputs(2309) <= a;
    layer3_outputs(2310) <= not (a or b);
    layer3_outputs(2311) <= b and not a;
    layer3_outputs(2312) <= a or b;
    layer3_outputs(2313) <= a;
    layer3_outputs(2314) <= not (a and b);
    layer3_outputs(2315) <= a and b;
    layer3_outputs(2316) <= not (a xor b);
    layer3_outputs(2317) <= a;
    layer3_outputs(2318) <= not b or a;
    layer3_outputs(2319) <= not b;
    layer3_outputs(2320) <= not (a and b);
    layer3_outputs(2321) <= b;
    layer3_outputs(2322) <= b;
    layer3_outputs(2323) <= a or b;
    layer3_outputs(2324) <= a;
    layer3_outputs(2325) <= not (a and b);
    layer3_outputs(2326) <= not (a or b);
    layer3_outputs(2327) <= not b or a;
    layer3_outputs(2328) <= not (a xor b);
    layer3_outputs(2329) <= a and not b;
    layer3_outputs(2330) <= a;
    layer3_outputs(2331) <= not a;
    layer3_outputs(2332) <= not b or a;
    layer3_outputs(2333) <= b;
    layer3_outputs(2334) <= not (a or b);
    layer3_outputs(2335) <= a and not b;
    layer3_outputs(2336) <= b;
    layer3_outputs(2337) <= not (a xor b);
    layer3_outputs(2338) <= not a or b;
    layer3_outputs(2339) <= a;
    layer3_outputs(2340) <= a and b;
    layer3_outputs(2341) <= b and not a;
    layer3_outputs(2342) <= a and b;
    layer3_outputs(2343) <= a;
    layer3_outputs(2344) <= not (a and b);
    layer3_outputs(2345) <= not a or b;
    layer3_outputs(2346) <= not (a or b);
    layer3_outputs(2347) <= b;
    layer3_outputs(2348) <= not (a or b);
    layer3_outputs(2349) <= a and not b;
    layer3_outputs(2350) <= not (a xor b);
    layer3_outputs(2351) <= not a;
    layer3_outputs(2352) <= not a;
    layer3_outputs(2353) <= 1'b1;
    layer3_outputs(2354) <= a;
    layer3_outputs(2355) <= not a or b;
    layer3_outputs(2356) <= b;
    layer3_outputs(2357) <= a xor b;
    layer3_outputs(2358) <= a and b;
    layer3_outputs(2359) <= 1'b1;
    layer3_outputs(2360) <= not b or a;
    layer3_outputs(2361) <= b;
    layer3_outputs(2362) <= not b;
    layer3_outputs(2363) <= a and b;
    layer3_outputs(2364) <= not b;
    layer3_outputs(2365) <= not a;
    layer3_outputs(2366) <= not a;
    layer3_outputs(2367) <= a;
    layer3_outputs(2368) <= not b;
    layer3_outputs(2369) <= b;
    layer3_outputs(2370) <= not b;
    layer3_outputs(2371) <= a;
    layer3_outputs(2372) <= not b or a;
    layer3_outputs(2373) <= not b or a;
    layer3_outputs(2374) <= a and b;
    layer3_outputs(2375) <= a and not b;
    layer3_outputs(2376) <= a or b;
    layer3_outputs(2377) <= b;
    layer3_outputs(2378) <= not b;
    layer3_outputs(2379) <= not a;
    layer3_outputs(2380) <= not b;
    layer3_outputs(2381) <= 1'b0;
    layer3_outputs(2382) <= not (a and b);
    layer3_outputs(2383) <= not b;
    layer3_outputs(2384) <= a and b;
    layer3_outputs(2385) <= b;
    layer3_outputs(2386) <= b and not a;
    layer3_outputs(2387) <= a and b;
    layer3_outputs(2388) <= not a or b;
    layer3_outputs(2389) <= a and b;
    layer3_outputs(2390) <= a or b;
    layer3_outputs(2391) <= not a;
    layer3_outputs(2392) <= b and not a;
    layer3_outputs(2393) <= not b;
    layer3_outputs(2394) <= not a;
    layer3_outputs(2395) <= a;
    layer3_outputs(2396) <= a and not b;
    layer3_outputs(2397) <= a and not b;
    layer3_outputs(2398) <= a xor b;
    layer3_outputs(2399) <= a and not b;
    layer3_outputs(2400) <= not a;
    layer3_outputs(2401) <= a and not b;
    layer3_outputs(2402) <= not (a or b);
    layer3_outputs(2403) <= a;
    layer3_outputs(2404) <= not b or a;
    layer3_outputs(2405) <= not (a or b);
    layer3_outputs(2406) <= not a;
    layer3_outputs(2407) <= a;
    layer3_outputs(2408) <= b;
    layer3_outputs(2409) <= not (a and b);
    layer3_outputs(2410) <= not a or b;
    layer3_outputs(2411) <= not b or a;
    layer3_outputs(2412) <= a and not b;
    layer3_outputs(2413) <= a and not b;
    layer3_outputs(2414) <= not a or b;
    layer3_outputs(2415) <= a and b;
    layer3_outputs(2416) <= not (a xor b);
    layer3_outputs(2417) <= not (a and b);
    layer3_outputs(2418) <= not (a xor b);
    layer3_outputs(2419) <= a and b;
    layer3_outputs(2420) <= a;
    layer3_outputs(2421) <= not a;
    layer3_outputs(2422) <= not b;
    layer3_outputs(2423) <= not (a and b);
    layer3_outputs(2424) <= not a or b;
    layer3_outputs(2425) <= b;
    layer3_outputs(2426) <= a and not b;
    layer3_outputs(2427) <= not b or a;
    layer3_outputs(2428) <= not a;
    layer3_outputs(2429) <= 1'b0;
    layer3_outputs(2430) <= not (a xor b);
    layer3_outputs(2431) <= a or b;
    layer3_outputs(2432) <= b and not a;
    layer3_outputs(2433) <= not (a xor b);
    layer3_outputs(2434) <= b and not a;
    layer3_outputs(2435) <= a and b;
    layer3_outputs(2436) <= not (a and b);
    layer3_outputs(2437) <= not (a and b);
    layer3_outputs(2438) <= not (a or b);
    layer3_outputs(2439) <= a and b;
    layer3_outputs(2440) <= b and not a;
    layer3_outputs(2441) <= not b;
    layer3_outputs(2442) <= a or b;
    layer3_outputs(2443) <= a xor b;
    layer3_outputs(2444) <= b and not a;
    layer3_outputs(2445) <= a;
    layer3_outputs(2446) <= not (a xor b);
    layer3_outputs(2447) <= not b;
    layer3_outputs(2448) <= a xor b;
    layer3_outputs(2449) <= b and not a;
    layer3_outputs(2450) <= a xor b;
    layer3_outputs(2451) <= not a;
    layer3_outputs(2452) <= b;
    layer3_outputs(2453) <= not a or b;
    layer3_outputs(2454) <= 1'b1;
    layer3_outputs(2455) <= b;
    layer3_outputs(2456) <= not (a xor b);
    layer3_outputs(2457) <= not b;
    layer3_outputs(2458) <= not a;
    layer3_outputs(2459) <= not (a xor b);
    layer3_outputs(2460) <= a;
    layer3_outputs(2461) <= not a;
    layer3_outputs(2462) <= a and b;
    layer3_outputs(2463) <= not a or b;
    layer3_outputs(2464) <= not b or a;
    layer3_outputs(2465) <= a;
    layer3_outputs(2466) <= a xor b;
    layer3_outputs(2467) <= b and not a;
    layer3_outputs(2468) <= a;
    layer3_outputs(2469) <= a;
    layer3_outputs(2470) <= a and b;
    layer3_outputs(2471) <= not b;
    layer3_outputs(2472) <= not (a and b);
    layer3_outputs(2473) <= not b or a;
    layer3_outputs(2474) <= a;
    layer3_outputs(2475) <= a;
    layer3_outputs(2476) <= 1'b1;
    layer3_outputs(2477) <= not b or a;
    layer3_outputs(2478) <= not b or a;
    layer3_outputs(2479) <= a;
    layer3_outputs(2480) <= not a;
    layer3_outputs(2481) <= a;
    layer3_outputs(2482) <= not (a and b);
    layer3_outputs(2483) <= b;
    layer3_outputs(2484) <= not (a or b);
    layer3_outputs(2485) <= not (a or b);
    layer3_outputs(2486) <= a;
    layer3_outputs(2487) <= a;
    layer3_outputs(2488) <= not a;
    layer3_outputs(2489) <= not b or a;
    layer3_outputs(2490) <= a xor b;
    layer3_outputs(2491) <= not a or b;
    layer3_outputs(2492) <= not (a xor b);
    layer3_outputs(2493) <= b;
    layer3_outputs(2494) <= not (a xor b);
    layer3_outputs(2495) <= b;
    layer3_outputs(2496) <= b;
    layer3_outputs(2497) <= a or b;
    layer3_outputs(2498) <= b;
    layer3_outputs(2499) <= b;
    layer3_outputs(2500) <= not b;
    layer3_outputs(2501) <= not b;
    layer3_outputs(2502) <= b;
    layer3_outputs(2503) <= not b or a;
    layer3_outputs(2504) <= not (a and b);
    layer3_outputs(2505) <= not b or a;
    layer3_outputs(2506) <= not (a and b);
    layer3_outputs(2507) <= a;
    layer3_outputs(2508) <= b;
    layer3_outputs(2509) <= a and b;
    layer3_outputs(2510) <= a xor b;
    layer3_outputs(2511) <= a or b;
    layer3_outputs(2512) <= a or b;
    layer3_outputs(2513) <= not a;
    layer3_outputs(2514) <= not b;
    layer3_outputs(2515) <= b and not a;
    layer3_outputs(2516) <= not b;
    layer3_outputs(2517) <= a and b;
    layer3_outputs(2518) <= b;
    layer3_outputs(2519) <= not b;
    layer3_outputs(2520) <= a;
    layer3_outputs(2521) <= a;
    layer3_outputs(2522) <= not (a and b);
    layer3_outputs(2523) <= a xor b;
    layer3_outputs(2524) <= not b or a;
    layer3_outputs(2525) <= not b or a;
    layer3_outputs(2526) <= not b;
    layer3_outputs(2527) <= not b or a;
    layer3_outputs(2528) <= not a or b;
    layer3_outputs(2529) <= not (a and b);
    layer3_outputs(2530) <= not (a xor b);
    layer3_outputs(2531) <= a or b;
    layer3_outputs(2532) <= not a;
    layer3_outputs(2533) <= not a;
    layer3_outputs(2534) <= a xor b;
    layer3_outputs(2535) <= not b;
    layer3_outputs(2536) <= not (a xor b);
    layer3_outputs(2537) <= not (a xor b);
    layer3_outputs(2538) <= a;
    layer3_outputs(2539) <= not a;
    layer3_outputs(2540) <= a xor b;
    layer3_outputs(2541) <= b;
    layer3_outputs(2542) <= b;
    layer3_outputs(2543) <= a and not b;
    layer3_outputs(2544) <= not b;
    layer3_outputs(2545) <= not b;
    layer3_outputs(2546) <= not a or b;
    layer3_outputs(2547) <= not a or b;
    layer3_outputs(2548) <= a and b;
    layer3_outputs(2549) <= not (a and b);
    layer3_outputs(2550) <= a xor b;
    layer3_outputs(2551) <= not a;
    layer3_outputs(2552) <= a xor b;
    layer3_outputs(2553) <= b;
    layer3_outputs(2554) <= not a;
    layer3_outputs(2555) <= b and not a;
    layer3_outputs(2556) <= not a or b;
    layer3_outputs(2557) <= not b;
    layer3_outputs(2558) <= not (a xor b);
    layer3_outputs(2559) <= a xor b;
    layer3_outputs(2560) <= a;
    layer3_outputs(2561) <= a;
    layer3_outputs(2562) <= a;
    layer3_outputs(2563) <= a;
    layer3_outputs(2564) <= a and b;
    layer3_outputs(2565) <= not b;
    layer3_outputs(2566) <= not b;
    layer3_outputs(2567) <= not a or b;
    layer3_outputs(2568) <= a and not b;
    layer3_outputs(2569) <= not (a and b);
    layer3_outputs(2570) <= not b or a;
    layer3_outputs(2571) <= b;
    layer3_outputs(2572) <= b;
    layer3_outputs(2573) <= a or b;
    layer3_outputs(2574) <= b;
    layer3_outputs(2575) <= not b;
    layer3_outputs(2576) <= not b;
    layer3_outputs(2577) <= b and not a;
    layer3_outputs(2578) <= b;
    layer3_outputs(2579) <= not a or b;
    layer3_outputs(2580) <= not a;
    layer3_outputs(2581) <= b;
    layer3_outputs(2582) <= a;
    layer3_outputs(2583) <= b;
    layer3_outputs(2584) <= b;
    layer3_outputs(2585) <= b and not a;
    layer3_outputs(2586) <= not b;
    layer3_outputs(2587) <= a or b;
    layer3_outputs(2588) <= not b or a;
    layer3_outputs(2589) <= not b;
    layer3_outputs(2590) <= not b or a;
    layer3_outputs(2591) <= a xor b;
    layer3_outputs(2592) <= b;
    layer3_outputs(2593) <= not (a xor b);
    layer3_outputs(2594) <= a and b;
    layer3_outputs(2595) <= a or b;
    layer3_outputs(2596) <= b;
    layer3_outputs(2597) <= not b;
    layer3_outputs(2598) <= b and not a;
    layer3_outputs(2599) <= b and not a;
    layer3_outputs(2600) <= b and not a;
    layer3_outputs(2601) <= a;
    layer3_outputs(2602) <= not (a and b);
    layer3_outputs(2603) <= a;
    layer3_outputs(2604) <= a;
    layer3_outputs(2605) <= not b;
    layer3_outputs(2606) <= 1'b1;
    layer3_outputs(2607) <= a and b;
    layer3_outputs(2608) <= not a;
    layer3_outputs(2609) <= not a;
    layer3_outputs(2610) <= not b;
    layer3_outputs(2611) <= not (a and b);
    layer3_outputs(2612) <= not (a and b);
    layer3_outputs(2613) <= not (a or b);
    layer3_outputs(2614) <= not a or b;
    layer3_outputs(2615) <= b;
    layer3_outputs(2616) <= not b;
    layer3_outputs(2617) <= a;
    layer3_outputs(2618) <= b;
    layer3_outputs(2619) <= 1'b0;
    layer3_outputs(2620) <= not a;
    layer3_outputs(2621) <= b;
    layer3_outputs(2622) <= a or b;
    layer3_outputs(2623) <= b;
    layer3_outputs(2624) <= a;
    layer3_outputs(2625) <= a xor b;
    layer3_outputs(2626) <= not (a and b);
    layer3_outputs(2627) <= not b or a;
    layer3_outputs(2628) <= not (a and b);
    layer3_outputs(2629) <= not a;
    layer3_outputs(2630) <= a;
    layer3_outputs(2631) <= b;
    layer3_outputs(2632) <= a;
    layer3_outputs(2633) <= not (a xor b);
    layer3_outputs(2634) <= not (a and b);
    layer3_outputs(2635) <= a;
    layer3_outputs(2636) <= not b;
    layer3_outputs(2637) <= b;
    layer3_outputs(2638) <= not a or b;
    layer3_outputs(2639) <= not b or a;
    layer3_outputs(2640) <= not (a and b);
    layer3_outputs(2641) <= a and b;
    layer3_outputs(2642) <= b;
    layer3_outputs(2643) <= not (a or b);
    layer3_outputs(2644) <= a;
    layer3_outputs(2645) <= a and b;
    layer3_outputs(2646) <= b;
    layer3_outputs(2647) <= a and b;
    layer3_outputs(2648) <= not a or b;
    layer3_outputs(2649) <= b and not a;
    layer3_outputs(2650) <= a and not b;
    layer3_outputs(2651) <= b;
    layer3_outputs(2652) <= a and b;
    layer3_outputs(2653) <= a;
    layer3_outputs(2654) <= not b;
    layer3_outputs(2655) <= a;
    layer3_outputs(2656) <= b;
    layer3_outputs(2657) <= not (a and b);
    layer3_outputs(2658) <= not a or b;
    layer3_outputs(2659) <= a;
    layer3_outputs(2660) <= not a or b;
    layer3_outputs(2661) <= not (a xor b);
    layer3_outputs(2662) <= b;
    layer3_outputs(2663) <= a and b;
    layer3_outputs(2664) <= a;
    layer3_outputs(2665) <= b;
    layer3_outputs(2666) <= a and b;
    layer3_outputs(2667) <= a xor b;
    layer3_outputs(2668) <= a and not b;
    layer3_outputs(2669) <= not a;
    layer3_outputs(2670) <= not (a or b);
    layer3_outputs(2671) <= not (a or b);
    layer3_outputs(2672) <= not a;
    layer3_outputs(2673) <= b;
    layer3_outputs(2674) <= a;
    layer3_outputs(2675) <= b and not a;
    layer3_outputs(2676) <= b;
    layer3_outputs(2677) <= not b or a;
    layer3_outputs(2678) <= not (a and b);
    layer3_outputs(2679) <= a and b;
    layer3_outputs(2680) <= a and not b;
    layer3_outputs(2681) <= not b or a;
    layer3_outputs(2682) <= not b;
    layer3_outputs(2683) <= not (a and b);
    layer3_outputs(2684) <= b;
    layer3_outputs(2685) <= b;
    layer3_outputs(2686) <= a;
    layer3_outputs(2687) <= not b;
    layer3_outputs(2688) <= a xor b;
    layer3_outputs(2689) <= a;
    layer3_outputs(2690) <= a or b;
    layer3_outputs(2691) <= not (a xor b);
    layer3_outputs(2692) <= b;
    layer3_outputs(2693) <= b;
    layer3_outputs(2694) <= not (a and b);
    layer3_outputs(2695) <= a and not b;
    layer3_outputs(2696) <= not (a or b);
    layer3_outputs(2697) <= a xor b;
    layer3_outputs(2698) <= 1'b0;
    layer3_outputs(2699) <= a xor b;
    layer3_outputs(2700) <= a or b;
    layer3_outputs(2701) <= b;
    layer3_outputs(2702) <= a;
    layer3_outputs(2703) <= a;
    layer3_outputs(2704) <= not (a or b);
    layer3_outputs(2705) <= not (a xor b);
    layer3_outputs(2706) <= a xor b;
    layer3_outputs(2707) <= a;
    layer3_outputs(2708) <= a;
    layer3_outputs(2709) <= a;
    layer3_outputs(2710) <= b;
    layer3_outputs(2711) <= a or b;
    layer3_outputs(2712) <= not b or a;
    layer3_outputs(2713) <= not a or b;
    layer3_outputs(2714) <= not b or a;
    layer3_outputs(2715) <= b;
    layer3_outputs(2716) <= a and not b;
    layer3_outputs(2717) <= b;
    layer3_outputs(2718) <= not (a xor b);
    layer3_outputs(2719) <= not (a or b);
    layer3_outputs(2720) <= a;
    layer3_outputs(2721) <= not (a xor b);
    layer3_outputs(2722) <= a and not b;
    layer3_outputs(2723) <= not b or a;
    layer3_outputs(2724) <= not a or b;
    layer3_outputs(2725) <= a xor b;
    layer3_outputs(2726) <= not (a xor b);
    layer3_outputs(2727) <= a and b;
    layer3_outputs(2728) <= not a;
    layer3_outputs(2729) <= a xor b;
    layer3_outputs(2730) <= a or b;
    layer3_outputs(2731) <= not (a xor b);
    layer3_outputs(2732) <= not b;
    layer3_outputs(2733) <= a and b;
    layer3_outputs(2734) <= not (a and b);
    layer3_outputs(2735) <= b;
    layer3_outputs(2736) <= not b;
    layer3_outputs(2737) <= a and not b;
    layer3_outputs(2738) <= not (a or b);
    layer3_outputs(2739) <= b;
    layer3_outputs(2740) <= b;
    layer3_outputs(2741) <= not b;
    layer3_outputs(2742) <= a;
    layer3_outputs(2743) <= not (a xor b);
    layer3_outputs(2744) <= not (a or b);
    layer3_outputs(2745) <= a and b;
    layer3_outputs(2746) <= a;
    layer3_outputs(2747) <= b;
    layer3_outputs(2748) <= b;
    layer3_outputs(2749) <= a or b;
    layer3_outputs(2750) <= not (a or b);
    layer3_outputs(2751) <= not b;
    layer3_outputs(2752) <= not (a or b);
    layer3_outputs(2753) <= not (a xor b);
    layer3_outputs(2754) <= b and not a;
    layer3_outputs(2755) <= a and b;
    layer3_outputs(2756) <= a and not b;
    layer3_outputs(2757) <= a;
    layer3_outputs(2758) <= a;
    layer3_outputs(2759) <= a;
    layer3_outputs(2760) <= not (a xor b);
    layer3_outputs(2761) <= 1'b1;
    layer3_outputs(2762) <= a xor b;
    layer3_outputs(2763) <= not a;
    layer3_outputs(2764) <= not a;
    layer3_outputs(2765) <= not a or b;
    layer3_outputs(2766) <= b;
    layer3_outputs(2767) <= not (a and b);
    layer3_outputs(2768) <= b;
    layer3_outputs(2769) <= not b;
    layer3_outputs(2770) <= a;
    layer3_outputs(2771) <= not a;
    layer3_outputs(2772) <= a xor b;
    layer3_outputs(2773) <= a and not b;
    layer3_outputs(2774) <= a xor b;
    layer3_outputs(2775) <= not (a xor b);
    layer3_outputs(2776) <= not b;
    layer3_outputs(2777) <= not a or b;
    layer3_outputs(2778) <= not a;
    layer3_outputs(2779) <= b;
    layer3_outputs(2780) <= not (a or b);
    layer3_outputs(2781) <= not b;
    layer3_outputs(2782) <= not b or a;
    layer3_outputs(2783) <= a xor b;
    layer3_outputs(2784) <= a;
    layer3_outputs(2785) <= 1'b1;
    layer3_outputs(2786) <= not (a xor b);
    layer3_outputs(2787) <= a and b;
    layer3_outputs(2788) <= not (a xor b);
    layer3_outputs(2789) <= 1'b0;
    layer3_outputs(2790) <= b;
    layer3_outputs(2791) <= not a or b;
    layer3_outputs(2792) <= a;
    layer3_outputs(2793) <= not b or a;
    layer3_outputs(2794) <= a and not b;
    layer3_outputs(2795) <= not b;
    layer3_outputs(2796) <= b;
    layer3_outputs(2797) <= a or b;
    layer3_outputs(2798) <= a and b;
    layer3_outputs(2799) <= not b or a;
    layer3_outputs(2800) <= not (a and b);
    layer3_outputs(2801) <= a;
    layer3_outputs(2802) <= a xor b;
    layer3_outputs(2803) <= a or b;
    layer3_outputs(2804) <= b and not a;
    layer3_outputs(2805) <= not (a xor b);
    layer3_outputs(2806) <= not a;
    layer3_outputs(2807) <= not a;
    layer3_outputs(2808) <= 1'b0;
    layer3_outputs(2809) <= a xor b;
    layer3_outputs(2810) <= a and not b;
    layer3_outputs(2811) <= a and b;
    layer3_outputs(2812) <= not b or a;
    layer3_outputs(2813) <= not b;
    layer3_outputs(2814) <= not a;
    layer3_outputs(2815) <= not a;
    layer3_outputs(2816) <= a or b;
    layer3_outputs(2817) <= not b or a;
    layer3_outputs(2818) <= not (a and b);
    layer3_outputs(2819) <= not (a or b);
    layer3_outputs(2820) <= not b;
    layer3_outputs(2821) <= a and b;
    layer3_outputs(2822) <= b;
    layer3_outputs(2823) <= a;
    layer3_outputs(2824) <= not b;
    layer3_outputs(2825) <= not b or a;
    layer3_outputs(2826) <= not (a or b);
    layer3_outputs(2827) <= a xor b;
    layer3_outputs(2828) <= not a;
    layer3_outputs(2829) <= not a;
    layer3_outputs(2830) <= a and b;
    layer3_outputs(2831) <= a xor b;
    layer3_outputs(2832) <= b and not a;
    layer3_outputs(2833) <= not b;
    layer3_outputs(2834) <= not b or a;
    layer3_outputs(2835) <= not b;
    layer3_outputs(2836) <= not a or b;
    layer3_outputs(2837) <= b;
    layer3_outputs(2838) <= b;
    layer3_outputs(2839) <= not (a and b);
    layer3_outputs(2840) <= not b or a;
    layer3_outputs(2841) <= not a;
    layer3_outputs(2842) <= not a;
    layer3_outputs(2843) <= a;
    layer3_outputs(2844) <= a xor b;
    layer3_outputs(2845) <= a;
    layer3_outputs(2846) <= a xor b;
    layer3_outputs(2847) <= b;
    layer3_outputs(2848) <= a xor b;
    layer3_outputs(2849) <= not (a or b);
    layer3_outputs(2850) <= a;
    layer3_outputs(2851) <= a and not b;
    layer3_outputs(2852) <= not a;
    layer3_outputs(2853) <= not a;
    layer3_outputs(2854) <= not (a or b);
    layer3_outputs(2855) <= b;
    layer3_outputs(2856) <= not (a xor b);
    layer3_outputs(2857) <= not (a or b);
    layer3_outputs(2858) <= a or b;
    layer3_outputs(2859) <= not b;
    layer3_outputs(2860) <= a or b;
    layer3_outputs(2861) <= b and not a;
    layer3_outputs(2862) <= a and not b;
    layer3_outputs(2863) <= a or b;
    layer3_outputs(2864) <= not a;
    layer3_outputs(2865) <= not (a or b);
    layer3_outputs(2866) <= not b;
    layer3_outputs(2867) <= not b or a;
    layer3_outputs(2868) <= b;
    layer3_outputs(2869) <= not (a xor b);
    layer3_outputs(2870) <= not (a or b);
    layer3_outputs(2871) <= b;
    layer3_outputs(2872) <= not (a xor b);
    layer3_outputs(2873) <= a and not b;
    layer3_outputs(2874) <= a;
    layer3_outputs(2875) <= not (a or b);
    layer3_outputs(2876) <= not b or a;
    layer3_outputs(2877) <= not b;
    layer3_outputs(2878) <= not a or b;
    layer3_outputs(2879) <= not (a xor b);
    layer3_outputs(2880) <= b;
    layer3_outputs(2881) <= not (a and b);
    layer3_outputs(2882) <= b;
    layer3_outputs(2883) <= b and not a;
    layer3_outputs(2884) <= a and not b;
    layer3_outputs(2885) <= a;
    layer3_outputs(2886) <= not a;
    layer3_outputs(2887) <= a and b;
    layer3_outputs(2888) <= a xor b;
    layer3_outputs(2889) <= a;
    layer3_outputs(2890) <= b and not a;
    layer3_outputs(2891) <= b;
    layer3_outputs(2892) <= not a or b;
    layer3_outputs(2893) <= not (a and b);
    layer3_outputs(2894) <= b;
    layer3_outputs(2895) <= not a;
    layer3_outputs(2896) <= not (a and b);
    layer3_outputs(2897) <= not b or a;
    layer3_outputs(2898) <= b;
    layer3_outputs(2899) <= a and not b;
    layer3_outputs(2900) <= not a;
    layer3_outputs(2901) <= not b;
    layer3_outputs(2902) <= a xor b;
    layer3_outputs(2903) <= a and b;
    layer3_outputs(2904) <= not b;
    layer3_outputs(2905) <= not a;
    layer3_outputs(2906) <= not a;
    layer3_outputs(2907) <= not (a and b);
    layer3_outputs(2908) <= not a;
    layer3_outputs(2909) <= 1'b1;
    layer3_outputs(2910) <= not a;
    layer3_outputs(2911) <= b and not a;
    layer3_outputs(2912) <= not a or b;
    layer3_outputs(2913) <= a;
    layer3_outputs(2914) <= not a;
    layer3_outputs(2915) <= b and not a;
    layer3_outputs(2916) <= not (a and b);
    layer3_outputs(2917) <= a and not b;
    layer3_outputs(2918) <= not a or b;
    layer3_outputs(2919) <= a or b;
    layer3_outputs(2920) <= not (a xor b);
    layer3_outputs(2921) <= a;
    layer3_outputs(2922) <= not a;
    layer3_outputs(2923) <= not a or b;
    layer3_outputs(2924) <= not (a xor b);
    layer3_outputs(2925) <= 1'b1;
    layer3_outputs(2926) <= not b;
    layer3_outputs(2927) <= not (a and b);
    layer3_outputs(2928) <= a;
    layer3_outputs(2929) <= not a or b;
    layer3_outputs(2930) <= a xor b;
    layer3_outputs(2931) <= not a or b;
    layer3_outputs(2932) <= not a or b;
    layer3_outputs(2933) <= b;
    layer3_outputs(2934) <= 1'b0;
    layer3_outputs(2935) <= a xor b;
    layer3_outputs(2936) <= not a or b;
    layer3_outputs(2937) <= not a or b;
    layer3_outputs(2938) <= 1'b1;
    layer3_outputs(2939) <= not a or b;
    layer3_outputs(2940) <= b;
    layer3_outputs(2941) <= not (a or b);
    layer3_outputs(2942) <= a;
    layer3_outputs(2943) <= a or b;
    layer3_outputs(2944) <= not (a or b);
    layer3_outputs(2945) <= a;
    layer3_outputs(2946) <= not (a and b);
    layer3_outputs(2947) <= a;
    layer3_outputs(2948) <= a;
    layer3_outputs(2949) <= a;
    layer3_outputs(2950) <= not a;
    layer3_outputs(2951) <= not (a xor b);
    layer3_outputs(2952) <= not b or a;
    layer3_outputs(2953) <= not b;
    layer3_outputs(2954) <= not b;
    layer3_outputs(2955) <= not a;
    layer3_outputs(2956) <= not b;
    layer3_outputs(2957) <= a xor b;
    layer3_outputs(2958) <= a and b;
    layer3_outputs(2959) <= a and not b;
    layer3_outputs(2960) <= a and not b;
    layer3_outputs(2961) <= a;
    layer3_outputs(2962) <= not a;
    layer3_outputs(2963) <= not b;
    layer3_outputs(2964) <= not (a and b);
    layer3_outputs(2965) <= not (a or b);
    layer3_outputs(2966) <= a or b;
    layer3_outputs(2967) <= not b;
    layer3_outputs(2968) <= not b;
    layer3_outputs(2969) <= b;
    layer3_outputs(2970) <= not b or a;
    layer3_outputs(2971) <= a;
    layer3_outputs(2972) <= a;
    layer3_outputs(2973) <= a and b;
    layer3_outputs(2974) <= b;
    layer3_outputs(2975) <= a or b;
    layer3_outputs(2976) <= a and b;
    layer3_outputs(2977) <= b;
    layer3_outputs(2978) <= b and not a;
    layer3_outputs(2979) <= not (a and b);
    layer3_outputs(2980) <= a and b;
    layer3_outputs(2981) <= a xor b;
    layer3_outputs(2982) <= not a;
    layer3_outputs(2983) <= not (a xor b);
    layer3_outputs(2984) <= a;
    layer3_outputs(2985) <= not (a or b);
    layer3_outputs(2986) <= a and b;
    layer3_outputs(2987) <= a and not b;
    layer3_outputs(2988) <= not a;
    layer3_outputs(2989) <= b and not a;
    layer3_outputs(2990) <= b and not a;
    layer3_outputs(2991) <= a;
    layer3_outputs(2992) <= a and not b;
    layer3_outputs(2993) <= a;
    layer3_outputs(2994) <= not b or a;
    layer3_outputs(2995) <= a or b;
    layer3_outputs(2996) <= not (a xor b);
    layer3_outputs(2997) <= a xor b;
    layer3_outputs(2998) <= not (a or b);
    layer3_outputs(2999) <= a and not b;
    layer3_outputs(3000) <= not b or a;
    layer3_outputs(3001) <= not (a and b);
    layer3_outputs(3002) <= a;
    layer3_outputs(3003) <= a;
    layer3_outputs(3004) <= a and not b;
    layer3_outputs(3005) <= b;
    layer3_outputs(3006) <= a and b;
    layer3_outputs(3007) <= a and b;
    layer3_outputs(3008) <= a xor b;
    layer3_outputs(3009) <= not b;
    layer3_outputs(3010) <= a and b;
    layer3_outputs(3011) <= a and b;
    layer3_outputs(3012) <= a;
    layer3_outputs(3013) <= not (a xor b);
    layer3_outputs(3014) <= a or b;
    layer3_outputs(3015) <= a;
    layer3_outputs(3016) <= a xor b;
    layer3_outputs(3017) <= b and not a;
    layer3_outputs(3018) <= b and not a;
    layer3_outputs(3019) <= b and not a;
    layer3_outputs(3020) <= not (a or b);
    layer3_outputs(3021) <= a xor b;
    layer3_outputs(3022) <= a and not b;
    layer3_outputs(3023) <= not b;
    layer3_outputs(3024) <= a;
    layer3_outputs(3025) <= b;
    layer3_outputs(3026) <= b;
    layer3_outputs(3027) <= not (a xor b);
    layer3_outputs(3028) <= not b or a;
    layer3_outputs(3029) <= b and not a;
    layer3_outputs(3030) <= a or b;
    layer3_outputs(3031) <= not (a and b);
    layer3_outputs(3032) <= a xor b;
    layer3_outputs(3033) <= not a or b;
    layer3_outputs(3034) <= a;
    layer3_outputs(3035) <= a;
    layer3_outputs(3036) <= not a;
    layer3_outputs(3037) <= a and b;
    layer3_outputs(3038) <= a and not b;
    layer3_outputs(3039) <= b;
    layer3_outputs(3040) <= 1'b1;
    layer3_outputs(3041) <= not a or b;
    layer3_outputs(3042) <= a;
    layer3_outputs(3043) <= not b or a;
    layer3_outputs(3044) <= b;
    layer3_outputs(3045) <= not (a and b);
    layer3_outputs(3046) <= not (a and b);
    layer3_outputs(3047) <= not b;
    layer3_outputs(3048) <= b;
    layer3_outputs(3049) <= a xor b;
    layer3_outputs(3050) <= not (a xor b);
    layer3_outputs(3051) <= not b;
    layer3_outputs(3052) <= not (a and b);
    layer3_outputs(3053) <= not b;
    layer3_outputs(3054) <= a or b;
    layer3_outputs(3055) <= not a or b;
    layer3_outputs(3056) <= not a;
    layer3_outputs(3057) <= not a;
    layer3_outputs(3058) <= not a or b;
    layer3_outputs(3059) <= not a or b;
    layer3_outputs(3060) <= not a;
    layer3_outputs(3061) <= not a;
    layer3_outputs(3062) <= b;
    layer3_outputs(3063) <= not a or b;
    layer3_outputs(3064) <= b;
    layer3_outputs(3065) <= a and not b;
    layer3_outputs(3066) <= not a or b;
    layer3_outputs(3067) <= not (a and b);
    layer3_outputs(3068) <= b;
    layer3_outputs(3069) <= a;
    layer3_outputs(3070) <= a and not b;
    layer3_outputs(3071) <= not (a and b);
    layer3_outputs(3072) <= not b;
    layer3_outputs(3073) <= a or b;
    layer3_outputs(3074) <= not (a or b);
    layer3_outputs(3075) <= not a;
    layer3_outputs(3076) <= b;
    layer3_outputs(3077) <= 1'b0;
    layer3_outputs(3078) <= not a;
    layer3_outputs(3079) <= not (a xor b);
    layer3_outputs(3080) <= not b;
    layer3_outputs(3081) <= b and not a;
    layer3_outputs(3082) <= not a or b;
    layer3_outputs(3083) <= b and not a;
    layer3_outputs(3084) <= b and not a;
    layer3_outputs(3085) <= not (a or b);
    layer3_outputs(3086) <= a and not b;
    layer3_outputs(3087) <= not (a and b);
    layer3_outputs(3088) <= not a or b;
    layer3_outputs(3089) <= a xor b;
    layer3_outputs(3090) <= a;
    layer3_outputs(3091) <= a and b;
    layer3_outputs(3092) <= not b or a;
    layer3_outputs(3093) <= not b or a;
    layer3_outputs(3094) <= a or b;
    layer3_outputs(3095) <= a or b;
    layer3_outputs(3096) <= not a;
    layer3_outputs(3097) <= a and b;
    layer3_outputs(3098) <= a;
    layer3_outputs(3099) <= not b;
    layer3_outputs(3100) <= not b or a;
    layer3_outputs(3101) <= a and b;
    layer3_outputs(3102) <= not a;
    layer3_outputs(3103) <= not (a and b);
    layer3_outputs(3104) <= b;
    layer3_outputs(3105) <= a and b;
    layer3_outputs(3106) <= not a;
    layer3_outputs(3107) <= not b;
    layer3_outputs(3108) <= a;
    layer3_outputs(3109) <= not (a xor b);
    layer3_outputs(3110) <= b;
    layer3_outputs(3111) <= not b;
    layer3_outputs(3112) <= not b;
    layer3_outputs(3113) <= not a;
    layer3_outputs(3114) <= b and not a;
    layer3_outputs(3115) <= not b;
    layer3_outputs(3116) <= b;
    layer3_outputs(3117) <= b and not a;
    layer3_outputs(3118) <= not (a or b);
    layer3_outputs(3119) <= a and b;
    layer3_outputs(3120) <= not a;
    layer3_outputs(3121) <= not (a xor b);
    layer3_outputs(3122) <= a;
    layer3_outputs(3123) <= not a;
    layer3_outputs(3124) <= a;
    layer3_outputs(3125) <= not b;
    layer3_outputs(3126) <= not b;
    layer3_outputs(3127) <= b;
    layer3_outputs(3128) <= not (a xor b);
    layer3_outputs(3129) <= a and not b;
    layer3_outputs(3130) <= a;
    layer3_outputs(3131) <= not b or a;
    layer3_outputs(3132) <= a xor b;
    layer3_outputs(3133) <= a;
    layer3_outputs(3134) <= not a;
    layer3_outputs(3135) <= not a or b;
    layer3_outputs(3136) <= not b or a;
    layer3_outputs(3137) <= b;
    layer3_outputs(3138) <= 1'b1;
    layer3_outputs(3139) <= not (a or b);
    layer3_outputs(3140) <= not b or a;
    layer3_outputs(3141) <= a;
    layer3_outputs(3142) <= a or b;
    layer3_outputs(3143) <= not (a or b);
    layer3_outputs(3144) <= a and not b;
    layer3_outputs(3145) <= b;
    layer3_outputs(3146) <= not (a and b);
    layer3_outputs(3147) <= a xor b;
    layer3_outputs(3148) <= not (a and b);
    layer3_outputs(3149) <= a;
    layer3_outputs(3150) <= b;
    layer3_outputs(3151) <= not b or a;
    layer3_outputs(3152) <= not (a or b);
    layer3_outputs(3153) <= not b or a;
    layer3_outputs(3154) <= not (a xor b);
    layer3_outputs(3155) <= a;
    layer3_outputs(3156) <= a;
    layer3_outputs(3157) <= not (a and b);
    layer3_outputs(3158) <= a;
    layer3_outputs(3159) <= a xor b;
    layer3_outputs(3160) <= a or b;
    layer3_outputs(3161) <= not b;
    layer3_outputs(3162) <= a;
    layer3_outputs(3163) <= not b;
    layer3_outputs(3164) <= b;
    layer3_outputs(3165) <= not (a and b);
    layer3_outputs(3166) <= b and not a;
    layer3_outputs(3167) <= a and b;
    layer3_outputs(3168) <= a and b;
    layer3_outputs(3169) <= b;
    layer3_outputs(3170) <= not a or b;
    layer3_outputs(3171) <= not a;
    layer3_outputs(3172) <= not b;
    layer3_outputs(3173) <= not (a and b);
    layer3_outputs(3174) <= a or b;
    layer3_outputs(3175) <= not a;
    layer3_outputs(3176) <= not b;
    layer3_outputs(3177) <= b and not a;
    layer3_outputs(3178) <= not b or a;
    layer3_outputs(3179) <= not (a or b);
    layer3_outputs(3180) <= a;
    layer3_outputs(3181) <= not b;
    layer3_outputs(3182) <= a xor b;
    layer3_outputs(3183) <= not b;
    layer3_outputs(3184) <= not b;
    layer3_outputs(3185) <= a and not b;
    layer3_outputs(3186) <= a and not b;
    layer3_outputs(3187) <= 1'b0;
    layer3_outputs(3188) <= a;
    layer3_outputs(3189) <= not (a and b);
    layer3_outputs(3190) <= not (a or b);
    layer3_outputs(3191) <= a and not b;
    layer3_outputs(3192) <= not b or a;
    layer3_outputs(3193) <= b;
    layer3_outputs(3194) <= a xor b;
    layer3_outputs(3195) <= not b;
    layer3_outputs(3196) <= b;
    layer3_outputs(3197) <= a xor b;
    layer3_outputs(3198) <= a or b;
    layer3_outputs(3199) <= a or b;
    layer3_outputs(3200) <= not b or a;
    layer3_outputs(3201) <= not (a xor b);
    layer3_outputs(3202) <= not b or a;
    layer3_outputs(3203) <= b;
    layer3_outputs(3204) <= not a or b;
    layer3_outputs(3205) <= not (a or b);
    layer3_outputs(3206) <= not a or b;
    layer3_outputs(3207) <= a xor b;
    layer3_outputs(3208) <= not a;
    layer3_outputs(3209) <= not a;
    layer3_outputs(3210) <= not a or b;
    layer3_outputs(3211) <= not (a xor b);
    layer3_outputs(3212) <= a;
    layer3_outputs(3213) <= a;
    layer3_outputs(3214) <= not a;
    layer3_outputs(3215) <= not (a and b);
    layer3_outputs(3216) <= not b or a;
    layer3_outputs(3217) <= not a or b;
    layer3_outputs(3218) <= not a;
    layer3_outputs(3219) <= not a or b;
    layer3_outputs(3220) <= not (a and b);
    layer3_outputs(3221) <= not b or a;
    layer3_outputs(3222) <= b;
    layer3_outputs(3223) <= not a or b;
    layer3_outputs(3224) <= b and not a;
    layer3_outputs(3225) <= not (a and b);
    layer3_outputs(3226) <= a;
    layer3_outputs(3227) <= b and not a;
    layer3_outputs(3228) <= not (a and b);
    layer3_outputs(3229) <= a and not b;
    layer3_outputs(3230) <= not a or b;
    layer3_outputs(3231) <= b;
    layer3_outputs(3232) <= not (a or b);
    layer3_outputs(3233) <= a or b;
    layer3_outputs(3234) <= not b;
    layer3_outputs(3235) <= not (a and b);
    layer3_outputs(3236) <= not b or a;
    layer3_outputs(3237) <= a and not b;
    layer3_outputs(3238) <= a;
    layer3_outputs(3239) <= b;
    layer3_outputs(3240) <= not (a or b);
    layer3_outputs(3241) <= not (a xor b);
    layer3_outputs(3242) <= not a;
    layer3_outputs(3243) <= not a or b;
    layer3_outputs(3244) <= a;
    layer3_outputs(3245) <= a or b;
    layer3_outputs(3246) <= b and not a;
    layer3_outputs(3247) <= b and not a;
    layer3_outputs(3248) <= 1'b1;
    layer3_outputs(3249) <= a;
    layer3_outputs(3250) <= not a;
    layer3_outputs(3251) <= not b or a;
    layer3_outputs(3252) <= a and not b;
    layer3_outputs(3253) <= b;
    layer3_outputs(3254) <= not b;
    layer3_outputs(3255) <= not (a and b);
    layer3_outputs(3256) <= not b;
    layer3_outputs(3257) <= a xor b;
    layer3_outputs(3258) <= b;
    layer3_outputs(3259) <= a;
    layer3_outputs(3260) <= not a or b;
    layer3_outputs(3261) <= a or b;
    layer3_outputs(3262) <= not a;
    layer3_outputs(3263) <= a xor b;
    layer3_outputs(3264) <= not (a xor b);
    layer3_outputs(3265) <= not b or a;
    layer3_outputs(3266) <= b and not a;
    layer3_outputs(3267) <= a;
    layer3_outputs(3268) <= not (a xor b);
    layer3_outputs(3269) <= b;
    layer3_outputs(3270) <= not b;
    layer3_outputs(3271) <= not (a and b);
    layer3_outputs(3272) <= b;
    layer3_outputs(3273) <= not (a xor b);
    layer3_outputs(3274) <= not (a and b);
    layer3_outputs(3275) <= not (a xor b);
    layer3_outputs(3276) <= b;
    layer3_outputs(3277) <= not (a or b);
    layer3_outputs(3278) <= not (a and b);
    layer3_outputs(3279) <= not (a and b);
    layer3_outputs(3280) <= not b;
    layer3_outputs(3281) <= b;
    layer3_outputs(3282) <= not a;
    layer3_outputs(3283) <= a;
    layer3_outputs(3284) <= not b;
    layer3_outputs(3285) <= b;
    layer3_outputs(3286) <= not (a xor b);
    layer3_outputs(3287) <= a;
    layer3_outputs(3288) <= b and not a;
    layer3_outputs(3289) <= not b;
    layer3_outputs(3290) <= b and not a;
    layer3_outputs(3291) <= a and b;
    layer3_outputs(3292) <= not b;
    layer3_outputs(3293) <= not (a xor b);
    layer3_outputs(3294) <= b and not a;
    layer3_outputs(3295) <= b;
    layer3_outputs(3296) <= not a;
    layer3_outputs(3297) <= b;
    layer3_outputs(3298) <= a xor b;
    layer3_outputs(3299) <= b;
    layer3_outputs(3300) <= a and not b;
    layer3_outputs(3301) <= not a;
    layer3_outputs(3302) <= a and b;
    layer3_outputs(3303) <= not a;
    layer3_outputs(3304) <= b;
    layer3_outputs(3305) <= b;
    layer3_outputs(3306) <= not a;
    layer3_outputs(3307) <= a;
    layer3_outputs(3308) <= b;
    layer3_outputs(3309) <= not b;
    layer3_outputs(3310) <= a xor b;
    layer3_outputs(3311) <= not a or b;
    layer3_outputs(3312) <= 1'b0;
    layer3_outputs(3313) <= a;
    layer3_outputs(3314) <= a;
    layer3_outputs(3315) <= a and not b;
    layer3_outputs(3316) <= not (a and b);
    layer3_outputs(3317) <= a;
    layer3_outputs(3318) <= not a or b;
    layer3_outputs(3319) <= a or b;
    layer3_outputs(3320) <= b;
    layer3_outputs(3321) <= a and not b;
    layer3_outputs(3322) <= not b or a;
    layer3_outputs(3323) <= not (a or b);
    layer3_outputs(3324) <= b;
    layer3_outputs(3325) <= not (a and b);
    layer3_outputs(3326) <= a or b;
    layer3_outputs(3327) <= not b;
    layer3_outputs(3328) <= a xor b;
    layer3_outputs(3329) <= not b;
    layer3_outputs(3330) <= a or b;
    layer3_outputs(3331) <= not b;
    layer3_outputs(3332) <= not a;
    layer3_outputs(3333) <= b and not a;
    layer3_outputs(3334) <= a xor b;
    layer3_outputs(3335) <= not (a and b);
    layer3_outputs(3336) <= a or b;
    layer3_outputs(3337) <= a and not b;
    layer3_outputs(3338) <= a;
    layer3_outputs(3339) <= a xor b;
    layer3_outputs(3340) <= not (a or b);
    layer3_outputs(3341) <= a and b;
    layer3_outputs(3342) <= not b;
    layer3_outputs(3343) <= not b;
    layer3_outputs(3344) <= not a;
    layer3_outputs(3345) <= b;
    layer3_outputs(3346) <= not a;
    layer3_outputs(3347) <= a and not b;
    layer3_outputs(3348) <= not a or b;
    layer3_outputs(3349) <= not b;
    layer3_outputs(3350) <= not a;
    layer3_outputs(3351) <= not b or a;
    layer3_outputs(3352) <= b;
    layer3_outputs(3353) <= not b;
    layer3_outputs(3354) <= b;
    layer3_outputs(3355) <= b;
    layer3_outputs(3356) <= not (a and b);
    layer3_outputs(3357) <= not b;
    layer3_outputs(3358) <= a xor b;
    layer3_outputs(3359) <= not b;
    layer3_outputs(3360) <= not a or b;
    layer3_outputs(3361) <= a and b;
    layer3_outputs(3362) <= not b;
    layer3_outputs(3363) <= a;
    layer3_outputs(3364) <= a;
    layer3_outputs(3365) <= a;
    layer3_outputs(3366) <= not (a xor b);
    layer3_outputs(3367) <= not b or a;
    layer3_outputs(3368) <= not (a xor b);
    layer3_outputs(3369) <= a and not b;
    layer3_outputs(3370) <= a and b;
    layer3_outputs(3371) <= a and not b;
    layer3_outputs(3372) <= b;
    layer3_outputs(3373) <= not b or a;
    layer3_outputs(3374) <= 1'b0;
    layer3_outputs(3375) <= a xor b;
    layer3_outputs(3376) <= a;
    layer3_outputs(3377) <= a and b;
    layer3_outputs(3378) <= not b;
    layer3_outputs(3379) <= not (a or b);
    layer3_outputs(3380) <= not b;
    layer3_outputs(3381) <= not b or a;
    layer3_outputs(3382) <= not a;
    layer3_outputs(3383) <= not a;
    layer3_outputs(3384) <= a;
    layer3_outputs(3385) <= b and not a;
    layer3_outputs(3386) <= not (a and b);
    layer3_outputs(3387) <= not (a xor b);
    layer3_outputs(3388) <= b and not a;
    layer3_outputs(3389) <= a and not b;
    layer3_outputs(3390) <= b;
    layer3_outputs(3391) <= b;
    layer3_outputs(3392) <= not a;
    layer3_outputs(3393) <= a and b;
    layer3_outputs(3394) <= not (a or b);
    layer3_outputs(3395) <= not b or a;
    layer3_outputs(3396) <= b and not a;
    layer3_outputs(3397) <= a and b;
    layer3_outputs(3398) <= a or b;
    layer3_outputs(3399) <= 1'b0;
    layer3_outputs(3400) <= a;
    layer3_outputs(3401) <= a and not b;
    layer3_outputs(3402) <= not a or b;
    layer3_outputs(3403) <= not a;
    layer3_outputs(3404) <= not b or a;
    layer3_outputs(3405) <= a;
    layer3_outputs(3406) <= b;
    layer3_outputs(3407) <= a and b;
    layer3_outputs(3408) <= b and not a;
    layer3_outputs(3409) <= a;
    layer3_outputs(3410) <= a or b;
    layer3_outputs(3411) <= a and b;
    layer3_outputs(3412) <= not (a or b);
    layer3_outputs(3413) <= not (a or b);
    layer3_outputs(3414) <= not (a or b);
    layer3_outputs(3415) <= not b;
    layer3_outputs(3416) <= a;
    layer3_outputs(3417) <= not a;
    layer3_outputs(3418) <= a and not b;
    layer3_outputs(3419) <= a and b;
    layer3_outputs(3420) <= a or b;
    layer3_outputs(3421) <= a and b;
    layer3_outputs(3422) <= not (a and b);
    layer3_outputs(3423) <= a xor b;
    layer3_outputs(3424) <= a and not b;
    layer3_outputs(3425) <= not (a and b);
    layer3_outputs(3426) <= not (a and b);
    layer3_outputs(3427) <= a and b;
    layer3_outputs(3428) <= not b;
    layer3_outputs(3429) <= b and not a;
    layer3_outputs(3430) <= b;
    layer3_outputs(3431) <= a;
    layer3_outputs(3432) <= not b or a;
    layer3_outputs(3433) <= not (a or b);
    layer3_outputs(3434) <= not (a and b);
    layer3_outputs(3435) <= 1'b1;
    layer3_outputs(3436) <= not (a or b);
    layer3_outputs(3437) <= a or b;
    layer3_outputs(3438) <= not b or a;
    layer3_outputs(3439) <= not (a and b);
    layer3_outputs(3440) <= 1'b0;
    layer3_outputs(3441) <= a xor b;
    layer3_outputs(3442) <= not b;
    layer3_outputs(3443) <= b and not a;
    layer3_outputs(3444) <= a and not b;
    layer3_outputs(3445) <= not b;
    layer3_outputs(3446) <= b;
    layer3_outputs(3447) <= a xor b;
    layer3_outputs(3448) <= not (a xor b);
    layer3_outputs(3449) <= not a;
    layer3_outputs(3450) <= not (a xor b);
    layer3_outputs(3451) <= a and b;
    layer3_outputs(3452) <= not b;
    layer3_outputs(3453) <= not (a or b);
    layer3_outputs(3454) <= not a;
    layer3_outputs(3455) <= a and not b;
    layer3_outputs(3456) <= a xor b;
    layer3_outputs(3457) <= not (a or b);
    layer3_outputs(3458) <= not a or b;
    layer3_outputs(3459) <= not b;
    layer3_outputs(3460) <= b;
    layer3_outputs(3461) <= a xor b;
    layer3_outputs(3462) <= not (a xor b);
    layer3_outputs(3463) <= not (a and b);
    layer3_outputs(3464) <= not (a or b);
    layer3_outputs(3465) <= not a;
    layer3_outputs(3466) <= a and not b;
    layer3_outputs(3467) <= not b;
    layer3_outputs(3468) <= a;
    layer3_outputs(3469) <= not b or a;
    layer3_outputs(3470) <= not b or a;
    layer3_outputs(3471) <= not a;
    layer3_outputs(3472) <= a or b;
    layer3_outputs(3473) <= not (a xor b);
    layer3_outputs(3474) <= not (a and b);
    layer3_outputs(3475) <= not (a xor b);
    layer3_outputs(3476) <= a and b;
    layer3_outputs(3477) <= a and b;
    layer3_outputs(3478) <= a and not b;
    layer3_outputs(3479) <= not a;
    layer3_outputs(3480) <= not a or b;
    layer3_outputs(3481) <= not b or a;
    layer3_outputs(3482) <= b;
    layer3_outputs(3483) <= not b;
    layer3_outputs(3484) <= a or b;
    layer3_outputs(3485) <= not (a or b);
    layer3_outputs(3486) <= 1'b0;
    layer3_outputs(3487) <= b and not a;
    layer3_outputs(3488) <= b;
    layer3_outputs(3489) <= not b or a;
    layer3_outputs(3490) <= not b or a;
    layer3_outputs(3491) <= b;
    layer3_outputs(3492) <= b;
    layer3_outputs(3493) <= not (a or b);
    layer3_outputs(3494) <= a xor b;
    layer3_outputs(3495) <= not (a and b);
    layer3_outputs(3496) <= not b;
    layer3_outputs(3497) <= a or b;
    layer3_outputs(3498) <= not (a or b);
    layer3_outputs(3499) <= not b;
    layer3_outputs(3500) <= not b;
    layer3_outputs(3501) <= a and not b;
    layer3_outputs(3502) <= not b or a;
    layer3_outputs(3503) <= a and b;
    layer3_outputs(3504) <= a;
    layer3_outputs(3505) <= not a;
    layer3_outputs(3506) <= not b;
    layer3_outputs(3507) <= a and b;
    layer3_outputs(3508) <= a;
    layer3_outputs(3509) <= b;
    layer3_outputs(3510) <= not b;
    layer3_outputs(3511) <= not a;
    layer3_outputs(3512) <= not (a and b);
    layer3_outputs(3513) <= not (a or b);
    layer3_outputs(3514) <= a or b;
    layer3_outputs(3515) <= not a or b;
    layer3_outputs(3516) <= not a;
    layer3_outputs(3517) <= not a or b;
    layer3_outputs(3518) <= a;
    layer3_outputs(3519) <= b;
    layer3_outputs(3520) <= a and not b;
    layer3_outputs(3521) <= not (a or b);
    layer3_outputs(3522) <= a;
    layer3_outputs(3523) <= a;
    layer3_outputs(3524) <= not a;
    layer3_outputs(3525) <= not (a or b);
    layer3_outputs(3526) <= b;
    layer3_outputs(3527) <= not a;
    layer3_outputs(3528) <= a and b;
    layer3_outputs(3529) <= not (a and b);
    layer3_outputs(3530) <= a xor b;
    layer3_outputs(3531) <= not (a and b);
    layer3_outputs(3532) <= not (a and b);
    layer3_outputs(3533) <= a;
    layer3_outputs(3534) <= a xor b;
    layer3_outputs(3535) <= a and b;
    layer3_outputs(3536) <= b;
    layer3_outputs(3537) <= a or b;
    layer3_outputs(3538) <= not a;
    layer3_outputs(3539) <= not b;
    layer3_outputs(3540) <= a and b;
    layer3_outputs(3541) <= not (a xor b);
    layer3_outputs(3542) <= not a;
    layer3_outputs(3543) <= not a or b;
    layer3_outputs(3544) <= not b or a;
    layer3_outputs(3545) <= a or b;
    layer3_outputs(3546) <= not b;
    layer3_outputs(3547) <= a;
    layer3_outputs(3548) <= not b;
    layer3_outputs(3549) <= a or b;
    layer3_outputs(3550) <= a and b;
    layer3_outputs(3551) <= a xor b;
    layer3_outputs(3552) <= b;
    layer3_outputs(3553) <= a;
    layer3_outputs(3554) <= not b;
    layer3_outputs(3555) <= not b or a;
    layer3_outputs(3556) <= a;
    layer3_outputs(3557) <= b and not a;
    layer3_outputs(3558) <= not a or b;
    layer3_outputs(3559) <= not (a xor b);
    layer3_outputs(3560) <= not (a xor b);
    layer3_outputs(3561) <= not b;
    layer3_outputs(3562) <= not (a or b);
    layer3_outputs(3563) <= not a or b;
    layer3_outputs(3564) <= b and not a;
    layer3_outputs(3565) <= a;
    layer3_outputs(3566) <= a;
    layer3_outputs(3567) <= b and not a;
    layer3_outputs(3568) <= not b;
    layer3_outputs(3569) <= not b;
    layer3_outputs(3570) <= b;
    layer3_outputs(3571) <= b and not a;
    layer3_outputs(3572) <= a and not b;
    layer3_outputs(3573) <= a;
    layer3_outputs(3574) <= b and not a;
    layer3_outputs(3575) <= a and not b;
    layer3_outputs(3576) <= b;
    layer3_outputs(3577) <= a;
    layer3_outputs(3578) <= 1'b0;
    layer3_outputs(3579) <= not a;
    layer3_outputs(3580) <= a and not b;
    layer3_outputs(3581) <= not (a xor b);
    layer3_outputs(3582) <= a;
    layer3_outputs(3583) <= a or b;
    layer3_outputs(3584) <= b;
    layer3_outputs(3585) <= a;
    layer3_outputs(3586) <= not b;
    layer3_outputs(3587) <= not a;
    layer3_outputs(3588) <= b and not a;
    layer3_outputs(3589) <= a and not b;
    layer3_outputs(3590) <= a xor b;
    layer3_outputs(3591) <= a and not b;
    layer3_outputs(3592) <= not a;
    layer3_outputs(3593) <= a xor b;
    layer3_outputs(3594) <= a;
    layer3_outputs(3595) <= a;
    layer3_outputs(3596) <= not b or a;
    layer3_outputs(3597) <= a or b;
    layer3_outputs(3598) <= b and not a;
    layer3_outputs(3599) <= a or b;
    layer3_outputs(3600) <= b;
    layer3_outputs(3601) <= not (a or b);
    layer3_outputs(3602) <= a and not b;
    layer3_outputs(3603) <= not a or b;
    layer3_outputs(3604) <= b;
    layer3_outputs(3605) <= b;
    layer3_outputs(3606) <= a or b;
    layer3_outputs(3607) <= a and not b;
    layer3_outputs(3608) <= not (a or b);
    layer3_outputs(3609) <= not b or a;
    layer3_outputs(3610) <= not a or b;
    layer3_outputs(3611) <= not a;
    layer3_outputs(3612) <= a or b;
    layer3_outputs(3613) <= not a;
    layer3_outputs(3614) <= not b;
    layer3_outputs(3615) <= not (a or b);
    layer3_outputs(3616) <= not (a xor b);
    layer3_outputs(3617) <= not b;
    layer3_outputs(3618) <= not b or a;
    layer3_outputs(3619) <= a or b;
    layer3_outputs(3620) <= a and not b;
    layer3_outputs(3621) <= b;
    layer3_outputs(3622) <= a;
    layer3_outputs(3623) <= b;
    layer3_outputs(3624) <= not a or b;
    layer3_outputs(3625) <= not a;
    layer3_outputs(3626) <= a;
    layer3_outputs(3627) <= a;
    layer3_outputs(3628) <= not (a or b);
    layer3_outputs(3629) <= a or b;
    layer3_outputs(3630) <= not a;
    layer3_outputs(3631) <= not (a xor b);
    layer3_outputs(3632) <= b and not a;
    layer3_outputs(3633) <= a;
    layer3_outputs(3634) <= a and not b;
    layer3_outputs(3635) <= a;
    layer3_outputs(3636) <= a and not b;
    layer3_outputs(3637) <= not (a xor b);
    layer3_outputs(3638) <= not a;
    layer3_outputs(3639) <= not (a xor b);
    layer3_outputs(3640) <= a or b;
    layer3_outputs(3641) <= b;
    layer3_outputs(3642) <= b;
    layer3_outputs(3643) <= not b;
    layer3_outputs(3644) <= b;
    layer3_outputs(3645) <= not (a or b);
    layer3_outputs(3646) <= not b or a;
    layer3_outputs(3647) <= a xor b;
    layer3_outputs(3648) <= b;
    layer3_outputs(3649) <= a or b;
    layer3_outputs(3650) <= 1'b1;
    layer3_outputs(3651) <= a and not b;
    layer3_outputs(3652) <= not a or b;
    layer3_outputs(3653) <= a;
    layer3_outputs(3654) <= b;
    layer3_outputs(3655) <= b;
    layer3_outputs(3656) <= a;
    layer3_outputs(3657) <= not (a or b);
    layer3_outputs(3658) <= a xor b;
    layer3_outputs(3659) <= not a;
    layer3_outputs(3660) <= b;
    layer3_outputs(3661) <= not a;
    layer3_outputs(3662) <= not (a xor b);
    layer3_outputs(3663) <= b;
    layer3_outputs(3664) <= not (a and b);
    layer3_outputs(3665) <= b;
    layer3_outputs(3666) <= a xor b;
    layer3_outputs(3667) <= a;
    layer3_outputs(3668) <= not (a xor b);
    layer3_outputs(3669) <= not (a xor b);
    layer3_outputs(3670) <= not b;
    layer3_outputs(3671) <= a xor b;
    layer3_outputs(3672) <= not b;
    layer3_outputs(3673) <= not (a and b);
    layer3_outputs(3674) <= a;
    layer3_outputs(3675) <= not (a xor b);
    layer3_outputs(3676) <= b and not a;
    layer3_outputs(3677) <= not (a and b);
    layer3_outputs(3678) <= not b;
    layer3_outputs(3679) <= a or b;
    layer3_outputs(3680) <= not (a and b);
    layer3_outputs(3681) <= b;
    layer3_outputs(3682) <= a;
    layer3_outputs(3683) <= not b or a;
    layer3_outputs(3684) <= not b or a;
    layer3_outputs(3685) <= b and not a;
    layer3_outputs(3686) <= not b;
    layer3_outputs(3687) <= not (a or b);
    layer3_outputs(3688) <= 1'b1;
    layer3_outputs(3689) <= not a or b;
    layer3_outputs(3690) <= not a;
    layer3_outputs(3691) <= not a;
    layer3_outputs(3692) <= not a or b;
    layer3_outputs(3693) <= not b;
    layer3_outputs(3694) <= not b;
    layer3_outputs(3695) <= b;
    layer3_outputs(3696) <= b;
    layer3_outputs(3697) <= not a;
    layer3_outputs(3698) <= 1'b0;
    layer3_outputs(3699) <= b;
    layer3_outputs(3700) <= a and b;
    layer3_outputs(3701) <= not a;
    layer3_outputs(3702) <= not a;
    layer3_outputs(3703) <= not (a xor b);
    layer3_outputs(3704) <= not (a and b);
    layer3_outputs(3705) <= not b;
    layer3_outputs(3706) <= not b;
    layer3_outputs(3707) <= b and not a;
    layer3_outputs(3708) <= a;
    layer3_outputs(3709) <= a and not b;
    layer3_outputs(3710) <= not a;
    layer3_outputs(3711) <= b;
    layer3_outputs(3712) <= not a;
    layer3_outputs(3713) <= a;
    layer3_outputs(3714) <= a xor b;
    layer3_outputs(3715) <= a;
    layer3_outputs(3716) <= b and not a;
    layer3_outputs(3717) <= a and not b;
    layer3_outputs(3718) <= not b;
    layer3_outputs(3719) <= b and not a;
    layer3_outputs(3720) <= a xor b;
    layer3_outputs(3721) <= a and not b;
    layer3_outputs(3722) <= not (a or b);
    layer3_outputs(3723) <= a xor b;
    layer3_outputs(3724) <= 1'b0;
    layer3_outputs(3725) <= a;
    layer3_outputs(3726) <= not (a xor b);
    layer3_outputs(3727) <= not (a xor b);
    layer3_outputs(3728) <= a or b;
    layer3_outputs(3729) <= not (a or b);
    layer3_outputs(3730) <= a xor b;
    layer3_outputs(3731) <= not (a or b);
    layer3_outputs(3732) <= a or b;
    layer3_outputs(3733) <= b;
    layer3_outputs(3734) <= not (a or b);
    layer3_outputs(3735) <= a and not b;
    layer3_outputs(3736) <= a;
    layer3_outputs(3737) <= a and b;
    layer3_outputs(3738) <= a and not b;
    layer3_outputs(3739) <= not (a or b);
    layer3_outputs(3740) <= a xor b;
    layer3_outputs(3741) <= not (a xor b);
    layer3_outputs(3742) <= not a;
    layer3_outputs(3743) <= a xor b;
    layer3_outputs(3744) <= not (a and b);
    layer3_outputs(3745) <= a or b;
    layer3_outputs(3746) <= a and b;
    layer3_outputs(3747) <= b;
    layer3_outputs(3748) <= not b or a;
    layer3_outputs(3749) <= a and not b;
    layer3_outputs(3750) <= not (a or b);
    layer3_outputs(3751) <= b and not a;
    layer3_outputs(3752) <= a and b;
    layer3_outputs(3753) <= b;
    layer3_outputs(3754) <= not (a and b);
    layer3_outputs(3755) <= not b;
    layer3_outputs(3756) <= a xor b;
    layer3_outputs(3757) <= a xor b;
    layer3_outputs(3758) <= b;
    layer3_outputs(3759) <= b and not a;
    layer3_outputs(3760) <= not (a and b);
    layer3_outputs(3761) <= not (a and b);
    layer3_outputs(3762) <= not (a xor b);
    layer3_outputs(3763) <= not a or b;
    layer3_outputs(3764) <= a;
    layer3_outputs(3765) <= a xor b;
    layer3_outputs(3766) <= b;
    layer3_outputs(3767) <= a;
    layer3_outputs(3768) <= a xor b;
    layer3_outputs(3769) <= a;
    layer3_outputs(3770) <= not b;
    layer3_outputs(3771) <= not b;
    layer3_outputs(3772) <= a and b;
    layer3_outputs(3773) <= not b or a;
    layer3_outputs(3774) <= a;
    layer3_outputs(3775) <= not (a xor b);
    layer3_outputs(3776) <= b;
    layer3_outputs(3777) <= not a or b;
    layer3_outputs(3778) <= a xor b;
    layer3_outputs(3779) <= not b or a;
    layer3_outputs(3780) <= a or b;
    layer3_outputs(3781) <= not a;
    layer3_outputs(3782) <= not a;
    layer3_outputs(3783) <= not b or a;
    layer3_outputs(3784) <= not a;
    layer3_outputs(3785) <= a;
    layer3_outputs(3786) <= a;
    layer3_outputs(3787) <= not (a xor b);
    layer3_outputs(3788) <= a or b;
    layer3_outputs(3789) <= not a;
    layer3_outputs(3790) <= b and not a;
    layer3_outputs(3791) <= 1'b0;
    layer3_outputs(3792) <= b;
    layer3_outputs(3793) <= b and not a;
    layer3_outputs(3794) <= not b;
    layer3_outputs(3795) <= not b;
    layer3_outputs(3796) <= b and not a;
    layer3_outputs(3797) <= a;
    layer3_outputs(3798) <= not a;
    layer3_outputs(3799) <= not (a xor b);
    layer3_outputs(3800) <= a;
    layer3_outputs(3801) <= b;
    layer3_outputs(3802) <= a;
    layer3_outputs(3803) <= not b or a;
    layer3_outputs(3804) <= not b;
    layer3_outputs(3805) <= not a;
    layer3_outputs(3806) <= not b or a;
    layer3_outputs(3807) <= not (a or b);
    layer3_outputs(3808) <= a;
    layer3_outputs(3809) <= not a or b;
    layer3_outputs(3810) <= a xor b;
    layer3_outputs(3811) <= a and not b;
    layer3_outputs(3812) <= b and not a;
    layer3_outputs(3813) <= not b;
    layer3_outputs(3814) <= not b;
    layer3_outputs(3815) <= b;
    layer3_outputs(3816) <= not (a and b);
    layer3_outputs(3817) <= b;
    layer3_outputs(3818) <= not a or b;
    layer3_outputs(3819) <= a or b;
    layer3_outputs(3820) <= b and not a;
    layer3_outputs(3821) <= not a;
    layer3_outputs(3822) <= b;
    layer3_outputs(3823) <= not b;
    layer3_outputs(3824) <= b;
    layer3_outputs(3825) <= not b;
    layer3_outputs(3826) <= not a;
    layer3_outputs(3827) <= b;
    layer3_outputs(3828) <= not a or b;
    layer3_outputs(3829) <= b and not a;
    layer3_outputs(3830) <= a;
    layer3_outputs(3831) <= b;
    layer3_outputs(3832) <= a or b;
    layer3_outputs(3833) <= b and not a;
    layer3_outputs(3834) <= not b or a;
    layer3_outputs(3835) <= not (a or b);
    layer3_outputs(3836) <= not (a xor b);
    layer3_outputs(3837) <= not (a xor b);
    layer3_outputs(3838) <= a;
    layer3_outputs(3839) <= not b;
    layer3_outputs(3840) <= not b;
    layer3_outputs(3841) <= not b;
    layer3_outputs(3842) <= b;
    layer3_outputs(3843) <= a;
    layer3_outputs(3844) <= a and not b;
    layer3_outputs(3845) <= not b or a;
    layer3_outputs(3846) <= a;
    layer3_outputs(3847) <= not (a or b);
    layer3_outputs(3848) <= a xor b;
    layer3_outputs(3849) <= b;
    layer3_outputs(3850) <= not b;
    layer3_outputs(3851) <= b;
    layer3_outputs(3852) <= a or b;
    layer3_outputs(3853) <= a and b;
    layer3_outputs(3854) <= not b;
    layer3_outputs(3855) <= not a;
    layer3_outputs(3856) <= not a or b;
    layer3_outputs(3857) <= not b or a;
    layer3_outputs(3858) <= b and not a;
    layer3_outputs(3859) <= not a;
    layer3_outputs(3860) <= a or b;
    layer3_outputs(3861) <= not (a xor b);
    layer3_outputs(3862) <= not a;
    layer3_outputs(3863) <= a or b;
    layer3_outputs(3864) <= not a;
    layer3_outputs(3865) <= not (a or b);
    layer3_outputs(3866) <= a and not b;
    layer3_outputs(3867) <= a and b;
    layer3_outputs(3868) <= b;
    layer3_outputs(3869) <= not (a xor b);
    layer3_outputs(3870) <= a;
    layer3_outputs(3871) <= a or b;
    layer3_outputs(3872) <= a or b;
    layer3_outputs(3873) <= a xor b;
    layer3_outputs(3874) <= b;
    layer3_outputs(3875) <= not b;
    layer3_outputs(3876) <= not b;
    layer3_outputs(3877) <= not a;
    layer3_outputs(3878) <= b;
    layer3_outputs(3879) <= not b or a;
    layer3_outputs(3880) <= not b or a;
    layer3_outputs(3881) <= not b;
    layer3_outputs(3882) <= b;
    layer3_outputs(3883) <= b;
    layer3_outputs(3884) <= not b or a;
    layer3_outputs(3885) <= a;
    layer3_outputs(3886) <= a;
    layer3_outputs(3887) <= not b;
    layer3_outputs(3888) <= 1'b1;
    layer3_outputs(3889) <= b;
    layer3_outputs(3890) <= a or b;
    layer3_outputs(3891) <= a and not b;
    layer3_outputs(3892) <= a and not b;
    layer3_outputs(3893) <= b;
    layer3_outputs(3894) <= not b;
    layer3_outputs(3895) <= not (a or b);
    layer3_outputs(3896) <= a xor b;
    layer3_outputs(3897) <= a or b;
    layer3_outputs(3898) <= not b or a;
    layer3_outputs(3899) <= b and not a;
    layer3_outputs(3900) <= a;
    layer3_outputs(3901) <= a xor b;
    layer3_outputs(3902) <= a xor b;
    layer3_outputs(3903) <= not a;
    layer3_outputs(3904) <= not a;
    layer3_outputs(3905) <= a;
    layer3_outputs(3906) <= a and not b;
    layer3_outputs(3907) <= not b;
    layer3_outputs(3908) <= not b;
    layer3_outputs(3909) <= not a or b;
    layer3_outputs(3910) <= not (a xor b);
    layer3_outputs(3911) <= not (a or b);
    layer3_outputs(3912) <= b;
    layer3_outputs(3913) <= a xor b;
    layer3_outputs(3914) <= not b;
    layer3_outputs(3915) <= b and not a;
    layer3_outputs(3916) <= a xor b;
    layer3_outputs(3917) <= not a;
    layer3_outputs(3918) <= not (a or b);
    layer3_outputs(3919) <= not (a or b);
    layer3_outputs(3920) <= b and not a;
    layer3_outputs(3921) <= not b or a;
    layer3_outputs(3922) <= not b;
    layer3_outputs(3923) <= not b;
    layer3_outputs(3924) <= a and not b;
    layer3_outputs(3925) <= not b or a;
    layer3_outputs(3926) <= not a;
    layer3_outputs(3927) <= b and not a;
    layer3_outputs(3928) <= 1'b0;
    layer3_outputs(3929) <= a;
    layer3_outputs(3930) <= a;
    layer3_outputs(3931) <= a or b;
    layer3_outputs(3932) <= a and not b;
    layer3_outputs(3933) <= not (a or b);
    layer3_outputs(3934) <= a xor b;
    layer3_outputs(3935) <= not (a xor b);
    layer3_outputs(3936) <= a;
    layer3_outputs(3937) <= a;
    layer3_outputs(3938) <= a or b;
    layer3_outputs(3939) <= not a;
    layer3_outputs(3940) <= b;
    layer3_outputs(3941) <= a;
    layer3_outputs(3942) <= b and not a;
    layer3_outputs(3943) <= not (a and b);
    layer3_outputs(3944) <= b and not a;
    layer3_outputs(3945) <= a xor b;
    layer3_outputs(3946) <= a or b;
    layer3_outputs(3947) <= not (a or b);
    layer3_outputs(3948) <= a;
    layer3_outputs(3949) <= not (a and b);
    layer3_outputs(3950) <= not b;
    layer3_outputs(3951) <= a;
    layer3_outputs(3952) <= not a or b;
    layer3_outputs(3953) <= a;
    layer3_outputs(3954) <= not b;
    layer3_outputs(3955) <= b and not a;
    layer3_outputs(3956) <= not a;
    layer3_outputs(3957) <= not a;
    layer3_outputs(3958) <= not (a and b);
    layer3_outputs(3959) <= b;
    layer3_outputs(3960) <= b;
    layer3_outputs(3961) <= a;
    layer3_outputs(3962) <= not b;
    layer3_outputs(3963) <= a xor b;
    layer3_outputs(3964) <= not b or a;
    layer3_outputs(3965) <= a or b;
    layer3_outputs(3966) <= a and not b;
    layer3_outputs(3967) <= a or b;
    layer3_outputs(3968) <= not (a xor b);
    layer3_outputs(3969) <= a;
    layer3_outputs(3970) <= not b or a;
    layer3_outputs(3971) <= b and not a;
    layer3_outputs(3972) <= not b;
    layer3_outputs(3973) <= b;
    layer3_outputs(3974) <= b and not a;
    layer3_outputs(3975) <= a and not b;
    layer3_outputs(3976) <= not (a xor b);
    layer3_outputs(3977) <= not a;
    layer3_outputs(3978) <= a or b;
    layer3_outputs(3979) <= a;
    layer3_outputs(3980) <= not (a or b);
    layer3_outputs(3981) <= not a or b;
    layer3_outputs(3982) <= not b or a;
    layer3_outputs(3983) <= a or b;
    layer3_outputs(3984) <= a and not b;
    layer3_outputs(3985) <= not a or b;
    layer3_outputs(3986) <= b and not a;
    layer3_outputs(3987) <= a;
    layer3_outputs(3988) <= not (a or b);
    layer3_outputs(3989) <= not (a xor b);
    layer3_outputs(3990) <= not (a or b);
    layer3_outputs(3991) <= not b;
    layer3_outputs(3992) <= a or b;
    layer3_outputs(3993) <= 1'b1;
    layer3_outputs(3994) <= not b;
    layer3_outputs(3995) <= b and not a;
    layer3_outputs(3996) <= not b or a;
    layer3_outputs(3997) <= not a;
    layer3_outputs(3998) <= not b;
    layer3_outputs(3999) <= not (a xor b);
    layer3_outputs(4000) <= not a or b;
    layer3_outputs(4001) <= not (a and b);
    layer3_outputs(4002) <= not b or a;
    layer3_outputs(4003) <= a xor b;
    layer3_outputs(4004) <= not a;
    layer3_outputs(4005) <= a and b;
    layer3_outputs(4006) <= not (a and b);
    layer3_outputs(4007) <= not b;
    layer3_outputs(4008) <= not a;
    layer3_outputs(4009) <= not a;
    layer3_outputs(4010) <= not a;
    layer3_outputs(4011) <= not b or a;
    layer3_outputs(4012) <= a;
    layer3_outputs(4013) <= not (a or b);
    layer3_outputs(4014) <= not (a or b);
    layer3_outputs(4015) <= not b;
    layer3_outputs(4016) <= not (a and b);
    layer3_outputs(4017) <= not b or a;
    layer3_outputs(4018) <= not (a xor b);
    layer3_outputs(4019) <= not (a or b);
    layer3_outputs(4020) <= not b;
    layer3_outputs(4021) <= not (a and b);
    layer3_outputs(4022) <= a;
    layer3_outputs(4023) <= not b;
    layer3_outputs(4024) <= not b;
    layer3_outputs(4025) <= not (a xor b);
    layer3_outputs(4026) <= b;
    layer3_outputs(4027) <= not b;
    layer3_outputs(4028) <= a xor b;
    layer3_outputs(4029) <= a and b;
    layer3_outputs(4030) <= 1'b0;
    layer3_outputs(4031) <= a and b;
    layer3_outputs(4032) <= not (a or b);
    layer3_outputs(4033) <= not (a or b);
    layer3_outputs(4034) <= not a;
    layer3_outputs(4035) <= not (a or b);
    layer3_outputs(4036) <= a or b;
    layer3_outputs(4037) <= a xor b;
    layer3_outputs(4038) <= a and not b;
    layer3_outputs(4039) <= a or b;
    layer3_outputs(4040) <= b and not a;
    layer3_outputs(4041) <= b and not a;
    layer3_outputs(4042) <= a and not b;
    layer3_outputs(4043) <= a;
    layer3_outputs(4044) <= not (a or b);
    layer3_outputs(4045) <= a;
    layer3_outputs(4046) <= b and not a;
    layer3_outputs(4047) <= not b;
    layer3_outputs(4048) <= a xor b;
    layer3_outputs(4049) <= a and b;
    layer3_outputs(4050) <= not b;
    layer3_outputs(4051) <= not b;
    layer3_outputs(4052) <= a or b;
    layer3_outputs(4053) <= a;
    layer3_outputs(4054) <= not b;
    layer3_outputs(4055) <= b and not a;
    layer3_outputs(4056) <= b;
    layer3_outputs(4057) <= not b or a;
    layer3_outputs(4058) <= not (a xor b);
    layer3_outputs(4059) <= b;
    layer3_outputs(4060) <= a or b;
    layer3_outputs(4061) <= not (a xor b);
    layer3_outputs(4062) <= b;
    layer3_outputs(4063) <= not a;
    layer3_outputs(4064) <= not (a xor b);
    layer3_outputs(4065) <= not b or a;
    layer3_outputs(4066) <= a;
    layer3_outputs(4067) <= a and b;
    layer3_outputs(4068) <= a xor b;
    layer3_outputs(4069) <= not (a or b);
    layer3_outputs(4070) <= b;
    layer3_outputs(4071) <= not a or b;
    layer3_outputs(4072) <= not b;
    layer3_outputs(4073) <= not a;
    layer3_outputs(4074) <= a or b;
    layer3_outputs(4075) <= not a;
    layer3_outputs(4076) <= a and b;
    layer3_outputs(4077) <= not b;
    layer3_outputs(4078) <= not (a and b);
    layer3_outputs(4079) <= b;
    layer3_outputs(4080) <= a or b;
    layer3_outputs(4081) <= not (a or b);
    layer3_outputs(4082) <= b;
    layer3_outputs(4083) <= not a or b;
    layer3_outputs(4084) <= a xor b;
    layer3_outputs(4085) <= b;
    layer3_outputs(4086) <= not (a xor b);
    layer3_outputs(4087) <= not (a or b);
    layer3_outputs(4088) <= a xor b;
    layer3_outputs(4089) <= not b;
    layer3_outputs(4090) <= b;
    layer3_outputs(4091) <= b and not a;
    layer3_outputs(4092) <= not a;
    layer3_outputs(4093) <= b and not a;
    layer3_outputs(4094) <= not a;
    layer3_outputs(4095) <= not (a xor b);
    layer3_outputs(4096) <= a and b;
    layer3_outputs(4097) <= b;
    layer3_outputs(4098) <= not (a and b);
    layer3_outputs(4099) <= not b;
    layer3_outputs(4100) <= not b or a;
    layer3_outputs(4101) <= a xor b;
    layer3_outputs(4102) <= a xor b;
    layer3_outputs(4103) <= a and not b;
    layer3_outputs(4104) <= not b;
    layer3_outputs(4105) <= not b or a;
    layer3_outputs(4106) <= not b;
    layer3_outputs(4107) <= not a;
    layer3_outputs(4108) <= b and not a;
    layer3_outputs(4109) <= not b;
    layer3_outputs(4110) <= a or b;
    layer3_outputs(4111) <= b;
    layer3_outputs(4112) <= a and b;
    layer3_outputs(4113) <= not (a and b);
    layer3_outputs(4114) <= not b;
    layer3_outputs(4115) <= b and not a;
    layer3_outputs(4116) <= not (a xor b);
    layer3_outputs(4117) <= not b;
    layer3_outputs(4118) <= not (a xor b);
    layer3_outputs(4119) <= a and b;
    layer3_outputs(4120) <= b;
    layer3_outputs(4121) <= a xor b;
    layer3_outputs(4122) <= not (a and b);
    layer3_outputs(4123) <= not (a or b);
    layer3_outputs(4124) <= not b;
    layer3_outputs(4125) <= b;
    layer3_outputs(4126) <= a xor b;
    layer3_outputs(4127) <= a xor b;
    layer3_outputs(4128) <= a or b;
    layer3_outputs(4129) <= 1'b0;
    layer3_outputs(4130) <= a;
    layer3_outputs(4131) <= a and not b;
    layer3_outputs(4132) <= not (a and b);
    layer3_outputs(4133) <= not b or a;
    layer3_outputs(4134) <= not (a or b);
    layer3_outputs(4135) <= not b;
    layer3_outputs(4136) <= not a or b;
    layer3_outputs(4137) <= not b;
    layer3_outputs(4138) <= not b;
    layer3_outputs(4139) <= a;
    layer3_outputs(4140) <= not (a or b);
    layer3_outputs(4141) <= b and not a;
    layer3_outputs(4142) <= not (a and b);
    layer3_outputs(4143) <= not (a and b);
    layer3_outputs(4144) <= a;
    layer3_outputs(4145) <= not a;
    layer3_outputs(4146) <= b;
    layer3_outputs(4147) <= not (a xor b);
    layer3_outputs(4148) <= not b or a;
    layer3_outputs(4149) <= not b or a;
    layer3_outputs(4150) <= a and not b;
    layer3_outputs(4151) <= not b;
    layer3_outputs(4152) <= not b;
    layer3_outputs(4153) <= not a or b;
    layer3_outputs(4154) <= not (a or b);
    layer3_outputs(4155) <= not a;
    layer3_outputs(4156) <= not b;
    layer3_outputs(4157) <= b;
    layer3_outputs(4158) <= 1'b0;
    layer3_outputs(4159) <= not (a xor b);
    layer3_outputs(4160) <= not a;
    layer3_outputs(4161) <= not a or b;
    layer3_outputs(4162) <= a xor b;
    layer3_outputs(4163) <= a;
    layer3_outputs(4164) <= a;
    layer3_outputs(4165) <= b;
    layer3_outputs(4166) <= not (a xor b);
    layer3_outputs(4167) <= a and b;
    layer3_outputs(4168) <= b;
    layer3_outputs(4169) <= b;
    layer3_outputs(4170) <= not a or b;
    layer3_outputs(4171) <= not b or a;
    layer3_outputs(4172) <= a and b;
    layer3_outputs(4173) <= b;
    layer3_outputs(4174) <= not (a and b);
    layer3_outputs(4175) <= not b or a;
    layer3_outputs(4176) <= not b;
    layer3_outputs(4177) <= a or b;
    layer3_outputs(4178) <= b and not a;
    layer3_outputs(4179) <= a xor b;
    layer3_outputs(4180) <= a;
    layer3_outputs(4181) <= b and not a;
    layer3_outputs(4182) <= not (a or b);
    layer3_outputs(4183) <= not (a and b);
    layer3_outputs(4184) <= not b;
    layer3_outputs(4185) <= not a;
    layer3_outputs(4186) <= not b or a;
    layer3_outputs(4187) <= not (a and b);
    layer3_outputs(4188) <= not b or a;
    layer3_outputs(4189) <= not (a or b);
    layer3_outputs(4190) <= a;
    layer3_outputs(4191) <= not b;
    layer3_outputs(4192) <= a;
    layer3_outputs(4193) <= b;
    layer3_outputs(4194) <= not a or b;
    layer3_outputs(4195) <= a;
    layer3_outputs(4196) <= not b;
    layer3_outputs(4197) <= a and b;
    layer3_outputs(4198) <= a;
    layer3_outputs(4199) <= not a;
    layer3_outputs(4200) <= a;
    layer3_outputs(4201) <= a and b;
    layer3_outputs(4202) <= 1'b1;
    layer3_outputs(4203) <= a and b;
    layer3_outputs(4204) <= not a or b;
    layer3_outputs(4205) <= not (a and b);
    layer3_outputs(4206) <= a;
    layer3_outputs(4207) <= not b;
    layer3_outputs(4208) <= a and b;
    layer3_outputs(4209) <= not (a and b);
    layer3_outputs(4210) <= b;
    layer3_outputs(4211) <= not a;
    layer3_outputs(4212) <= not a;
    layer3_outputs(4213) <= a;
    layer3_outputs(4214) <= not a;
    layer3_outputs(4215) <= not b or a;
    layer3_outputs(4216) <= not (a and b);
    layer3_outputs(4217) <= not (a and b);
    layer3_outputs(4218) <= a and not b;
    layer3_outputs(4219) <= not (a and b);
    layer3_outputs(4220) <= not a;
    layer3_outputs(4221) <= a or b;
    layer3_outputs(4222) <= not (a xor b);
    layer3_outputs(4223) <= a xor b;
    layer3_outputs(4224) <= not b;
    layer3_outputs(4225) <= not a;
    layer3_outputs(4226) <= b;
    layer3_outputs(4227) <= not a;
    layer3_outputs(4228) <= a and not b;
    layer3_outputs(4229) <= not b;
    layer3_outputs(4230) <= not a;
    layer3_outputs(4231) <= not (a and b);
    layer3_outputs(4232) <= a xor b;
    layer3_outputs(4233) <= not a;
    layer3_outputs(4234) <= not b;
    layer3_outputs(4235) <= not (a xor b);
    layer3_outputs(4236) <= b;
    layer3_outputs(4237) <= a or b;
    layer3_outputs(4238) <= not b;
    layer3_outputs(4239) <= not b;
    layer3_outputs(4240) <= not (a and b);
    layer3_outputs(4241) <= a and b;
    layer3_outputs(4242) <= not b or a;
    layer3_outputs(4243) <= not b or a;
    layer3_outputs(4244) <= not b;
    layer3_outputs(4245) <= a or b;
    layer3_outputs(4246) <= a or b;
    layer3_outputs(4247) <= a;
    layer3_outputs(4248) <= a or b;
    layer3_outputs(4249) <= b;
    layer3_outputs(4250) <= b and not a;
    layer3_outputs(4251) <= not a;
    layer3_outputs(4252) <= a and not b;
    layer3_outputs(4253) <= b;
    layer3_outputs(4254) <= not (a and b);
    layer3_outputs(4255) <= not a or b;
    layer3_outputs(4256) <= b and not a;
    layer3_outputs(4257) <= b;
    layer3_outputs(4258) <= a xor b;
    layer3_outputs(4259) <= not (a xor b);
    layer3_outputs(4260) <= not b;
    layer3_outputs(4261) <= not (a and b);
    layer3_outputs(4262) <= not (a or b);
    layer3_outputs(4263) <= a and not b;
    layer3_outputs(4264) <= a and b;
    layer3_outputs(4265) <= not b;
    layer3_outputs(4266) <= a and not b;
    layer3_outputs(4267) <= not (a or b);
    layer3_outputs(4268) <= not (a and b);
    layer3_outputs(4269) <= a and b;
    layer3_outputs(4270) <= not b;
    layer3_outputs(4271) <= a and b;
    layer3_outputs(4272) <= b;
    layer3_outputs(4273) <= a and b;
    layer3_outputs(4274) <= not (a and b);
    layer3_outputs(4275) <= a and b;
    layer3_outputs(4276) <= a and b;
    layer3_outputs(4277) <= not (a xor b);
    layer3_outputs(4278) <= a;
    layer3_outputs(4279) <= not (a or b);
    layer3_outputs(4280) <= not b;
    layer3_outputs(4281) <= not (a or b);
    layer3_outputs(4282) <= b;
    layer3_outputs(4283) <= a or b;
    layer3_outputs(4284) <= b;
    layer3_outputs(4285) <= b and not a;
    layer3_outputs(4286) <= not a;
    layer3_outputs(4287) <= not b or a;
    layer3_outputs(4288) <= 1'b1;
    layer3_outputs(4289) <= not a;
    layer3_outputs(4290) <= a and not b;
    layer3_outputs(4291) <= a or b;
    layer3_outputs(4292) <= not a;
    layer3_outputs(4293) <= a and b;
    layer3_outputs(4294) <= a and not b;
    layer3_outputs(4295) <= not b or a;
    layer3_outputs(4296) <= a and not b;
    layer3_outputs(4297) <= not a;
    layer3_outputs(4298) <= b;
    layer3_outputs(4299) <= not a;
    layer3_outputs(4300) <= not a;
    layer3_outputs(4301) <= a xor b;
    layer3_outputs(4302) <= not b or a;
    layer3_outputs(4303) <= not b or a;
    layer3_outputs(4304) <= a;
    layer3_outputs(4305) <= not b or a;
    layer3_outputs(4306) <= a;
    layer3_outputs(4307) <= 1'b1;
    layer3_outputs(4308) <= a;
    layer3_outputs(4309) <= b;
    layer3_outputs(4310) <= not (a xor b);
    layer3_outputs(4311) <= a xor b;
    layer3_outputs(4312) <= not (a and b);
    layer3_outputs(4313) <= a;
    layer3_outputs(4314) <= not (a or b);
    layer3_outputs(4315) <= b;
    layer3_outputs(4316) <= not (a xor b);
    layer3_outputs(4317) <= a and not b;
    layer3_outputs(4318) <= a;
    layer3_outputs(4319) <= not a;
    layer3_outputs(4320) <= a and b;
    layer3_outputs(4321) <= not (a xor b);
    layer3_outputs(4322) <= not b or a;
    layer3_outputs(4323) <= not b;
    layer3_outputs(4324) <= a;
    layer3_outputs(4325) <= a xor b;
    layer3_outputs(4326) <= not b or a;
    layer3_outputs(4327) <= not a;
    layer3_outputs(4328) <= not (a or b);
    layer3_outputs(4329) <= a and b;
    layer3_outputs(4330) <= not a;
    layer3_outputs(4331) <= a and not b;
    layer3_outputs(4332) <= a and b;
    layer3_outputs(4333) <= a xor b;
    layer3_outputs(4334) <= not (a or b);
    layer3_outputs(4335) <= b;
    layer3_outputs(4336) <= a;
    layer3_outputs(4337) <= b and not a;
    layer3_outputs(4338) <= not b;
    layer3_outputs(4339) <= a and b;
    layer3_outputs(4340) <= not a or b;
    layer3_outputs(4341) <= not (a xor b);
    layer3_outputs(4342) <= 1'b1;
    layer3_outputs(4343) <= a xor b;
    layer3_outputs(4344) <= b;
    layer3_outputs(4345) <= not (a or b);
    layer3_outputs(4346) <= a and not b;
    layer3_outputs(4347) <= not b or a;
    layer3_outputs(4348) <= a;
    layer3_outputs(4349) <= not (a and b);
    layer3_outputs(4350) <= not (a or b);
    layer3_outputs(4351) <= a;
    layer3_outputs(4352) <= not (a or b);
    layer3_outputs(4353) <= a and not b;
    layer3_outputs(4354) <= not a or b;
    layer3_outputs(4355) <= a;
    layer3_outputs(4356) <= not (a xor b);
    layer3_outputs(4357) <= a and b;
    layer3_outputs(4358) <= a xor b;
    layer3_outputs(4359) <= not b or a;
    layer3_outputs(4360) <= b;
    layer3_outputs(4361) <= not a or b;
    layer3_outputs(4362) <= a xor b;
    layer3_outputs(4363) <= b and not a;
    layer3_outputs(4364) <= a;
    layer3_outputs(4365) <= b;
    layer3_outputs(4366) <= a and b;
    layer3_outputs(4367) <= b;
    layer3_outputs(4368) <= not b;
    layer3_outputs(4369) <= not (a and b);
    layer3_outputs(4370) <= not a or b;
    layer3_outputs(4371) <= not b or a;
    layer3_outputs(4372) <= not b;
    layer3_outputs(4373) <= a and not b;
    layer3_outputs(4374) <= not b;
    layer3_outputs(4375) <= not a;
    layer3_outputs(4376) <= a xor b;
    layer3_outputs(4377) <= not b;
    layer3_outputs(4378) <= a or b;
    layer3_outputs(4379) <= not b or a;
    layer3_outputs(4380) <= not (a xor b);
    layer3_outputs(4381) <= not (a or b);
    layer3_outputs(4382) <= a or b;
    layer3_outputs(4383) <= not a;
    layer3_outputs(4384) <= not (a xor b);
    layer3_outputs(4385) <= not (a and b);
    layer3_outputs(4386) <= b;
    layer3_outputs(4387) <= not b;
    layer3_outputs(4388) <= a and b;
    layer3_outputs(4389) <= a and not b;
    layer3_outputs(4390) <= b;
    layer3_outputs(4391) <= b;
    layer3_outputs(4392) <= not (a and b);
    layer3_outputs(4393) <= a xor b;
    layer3_outputs(4394) <= not a;
    layer3_outputs(4395) <= a;
    layer3_outputs(4396) <= b;
    layer3_outputs(4397) <= not b;
    layer3_outputs(4398) <= not (a or b);
    layer3_outputs(4399) <= not a;
    layer3_outputs(4400) <= not b or a;
    layer3_outputs(4401) <= b;
    layer3_outputs(4402) <= 1'b0;
    layer3_outputs(4403) <= not (a and b);
    layer3_outputs(4404) <= a and b;
    layer3_outputs(4405) <= b and not a;
    layer3_outputs(4406) <= not (a xor b);
    layer3_outputs(4407) <= a and not b;
    layer3_outputs(4408) <= not b;
    layer3_outputs(4409) <= not (a and b);
    layer3_outputs(4410) <= not (a xor b);
    layer3_outputs(4411) <= not b;
    layer3_outputs(4412) <= not b;
    layer3_outputs(4413) <= not (a xor b);
    layer3_outputs(4414) <= b;
    layer3_outputs(4415) <= not a;
    layer3_outputs(4416) <= not b;
    layer3_outputs(4417) <= a xor b;
    layer3_outputs(4418) <= b and not a;
    layer3_outputs(4419) <= not (a and b);
    layer3_outputs(4420) <= b and not a;
    layer3_outputs(4421) <= a;
    layer3_outputs(4422) <= not b;
    layer3_outputs(4423) <= not a;
    layer3_outputs(4424) <= not (a and b);
    layer3_outputs(4425) <= not a or b;
    layer3_outputs(4426) <= not (a and b);
    layer3_outputs(4427) <= not (a or b);
    layer3_outputs(4428) <= a and not b;
    layer3_outputs(4429) <= b and not a;
    layer3_outputs(4430) <= a;
    layer3_outputs(4431) <= not b;
    layer3_outputs(4432) <= a and b;
    layer3_outputs(4433) <= not b;
    layer3_outputs(4434) <= not b;
    layer3_outputs(4435) <= b and not a;
    layer3_outputs(4436) <= not a;
    layer3_outputs(4437) <= b;
    layer3_outputs(4438) <= a and not b;
    layer3_outputs(4439) <= a;
    layer3_outputs(4440) <= a and not b;
    layer3_outputs(4441) <= not (a and b);
    layer3_outputs(4442) <= not (a and b);
    layer3_outputs(4443) <= not b;
    layer3_outputs(4444) <= a and b;
    layer3_outputs(4445) <= not b;
    layer3_outputs(4446) <= not (a xor b);
    layer3_outputs(4447) <= not (a xor b);
    layer3_outputs(4448) <= not a;
    layer3_outputs(4449) <= not a or b;
    layer3_outputs(4450) <= a;
    layer3_outputs(4451) <= a and not b;
    layer3_outputs(4452) <= not b or a;
    layer3_outputs(4453) <= not a or b;
    layer3_outputs(4454) <= not a;
    layer3_outputs(4455) <= a;
    layer3_outputs(4456) <= a and b;
    layer3_outputs(4457) <= a;
    layer3_outputs(4458) <= not (a xor b);
    layer3_outputs(4459) <= not (a xor b);
    layer3_outputs(4460) <= not a or b;
    layer3_outputs(4461) <= not (a xor b);
    layer3_outputs(4462) <= not a;
    layer3_outputs(4463) <= not b or a;
    layer3_outputs(4464) <= a and not b;
    layer3_outputs(4465) <= not b;
    layer3_outputs(4466) <= not b or a;
    layer3_outputs(4467) <= 1'b0;
    layer3_outputs(4468) <= not (a or b);
    layer3_outputs(4469) <= not a;
    layer3_outputs(4470) <= a and not b;
    layer3_outputs(4471) <= b;
    layer3_outputs(4472) <= not (a or b);
    layer3_outputs(4473) <= a;
    layer3_outputs(4474) <= not b or a;
    layer3_outputs(4475) <= a and b;
    layer3_outputs(4476) <= not b;
    layer3_outputs(4477) <= b;
    layer3_outputs(4478) <= not (a or b);
    layer3_outputs(4479) <= not a;
    layer3_outputs(4480) <= a or b;
    layer3_outputs(4481) <= not (a xor b);
    layer3_outputs(4482) <= a;
    layer3_outputs(4483) <= a;
    layer3_outputs(4484) <= not b or a;
    layer3_outputs(4485) <= a;
    layer3_outputs(4486) <= not a;
    layer3_outputs(4487) <= not b or a;
    layer3_outputs(4488) <= a;
    layer3_outputs(4489) <= a and not b;
    layer3_outputs(4490) <= not (a or b);
    layer3_outputs(4491) <= not (a or b);
    layer3_outputs(4492) <= not a;
    layer3_outputs(4493) <= a xor b;
    layer3_outputs(4494) <= a or b;
    layer3_outputs(4495) <= a xor b;
    layer3_outputs(4496) <= a;
    layer3_outputs(4497) <= not (a xor b);
    layer3_outputs(4498) <= a;
    layer3_outputs(4499) <= b;
    layer3_outputs(4500) <= not a or b;
    layer3_outputs(4501) <= not (a or b);
    layer3_outputs(4502) <= a;
    layer3_outputs(4503) <= b;
    layer3_outputs(4504) <= a;
    layer3_outputs(4505) <= not (a and b);
    layer3_outputs(4506) <= not a;
    layer3_outputs(4507) <= not b;
    layer3_outputs(4508) <= not a;
    layer3_outputs(4509) <= a or b;
    layer3_outputs(4510) <= a or b;
    layer3_outputs(4511) <= a and b;
    layer3_outputs(4512) <= not (a and b);
    layer3_outputs(4513) <= a or b;
    layer3_outputs(4514) <= not a;
    layer3_outputs(4515) <= not b;
    layer3_outputs(4516) <= a and not b;
    layer3_outputs(4517) <= not b;
    layer3_outputs(4518) <= a and not b;
    layer3_outputs(4519) <= not a;
    layer3_outputs(4520) <= a and not b;
    layer3_outputs(4521) <= not b;
    layer3_outputs(4522) <= not a;
    layer3_outputs(4523) <= b;
    layer3_outputs(4524) <= b;
    layer3_outputs(4525) <= not a or b;
    layer3_outputs(4526) <= b and not a;
    layer3_outputs(4527) <= a;
    layer3_outputs(4528) <= b;
    layer3_outputs(4529) <= a and b;
    layer3_outputs(4530) <= a or b;
    layer3_outputs(4531) <= a;
    layer3_outputs(4532) <= not b;
    layer3_outputs(4533) <= not a or b;
    layer3_outputs(4534) <= b and not a;
    layer3_outputs(4535) <= 1'b1;
    layer3_outputs(4536) <= not (a xor b);
    layer3_outputs(4537) <= not a;
    layer3_outputs(4538) <= a and b;
    layer3_outputs(4539) <= b;
    layer3_outputs(4540) <= not b;
    layer3_outputs(4541) <= a xor b;
    layer3_outputs(4542) <= a xor b;
    layer3_outputs(4543) <= b and not a;
    layer3_outputs(4544) <= not (a and b);
    layer3_outputs(4545) <= not a;
    layer3_outputs(4546) <= 1'b1;
    layer3_outputs(4547) <= a and b;
    layer3_outputs(4548) <= not b;
    layer3_outputs(4549) <= a and b;
    layer3_outputs(4550) <= a;
    layer3_outputs(4551) <= a xor b;
    layer3_outputs(4552) <= a xor b;
    layer3_outputs(4553) <= not b;
    layer3_outputs(4554) <= b and not a;
    layer3_outputs(4555) <= not (a or b);
    layer3_outputs(4556) <= b;
    layer3_outputs(4557) <= not b or a;
    layer3_outputs(4558) <= a and b;
    layer3_outputs(4559) <= not b or a;
    layer3_outputs(4560) <= b;
    layer3_outputs(4561) <= not b or a;
    layer3_outputs(4562) <= not a;
    layer3_outputs(4563) <= not b;
    layer3_outputs(4564) <= a;
    layer3_outputs(4565) <= a xor b;
    layer3_outputs(4566) <= a and not b;
    layer3_outputs(4567) <= a and not b;
    layer3_outputs(4568) <= not a or b;
    layer3_outputs(4569) <= b;
    layer3_outputs(4570) <= not a or b;
    layer3_outputs(4571) <= b;
    layer3_outputs(4572) <= a and b;
    layer3_outputs(4573) <= 1'b1;
    layer3_outputs(4574) <= not b or a;
    layer3_outputs(4575) <= not b or a;
    layer3_outputs(4576) <= b;
    layer3_outputs(4577) <= not b or a;
    layer3_outputs(4578) <= not b or a;
    layer3_outputs(4579) <= not b or a;
    layer3_outputs(4580) <= b;
    layer3_outputs(4581) <= not b or a;
    layer3_outputs(4582) <= b;
    layer3_outputs(4583) <= b;
    layer3_outputs(4584) <= not (a and b);
    layer3_outputs(4585) <= not b;
    layer3_outputs(4586) <= b and not a;
    layer3_outputs(4587) <= not b;
    layer3_outputs(4588) <= not (a or b);
    layer3_outputs(4589) <= not a or b;
    layer3_outputs(4590) <= b;
    layer3_outputs(4591) <= not b;
    layer3_outputs(4592) <= not b;
    layer3_outputs(4593) <= a and not b;
    layer3_outputs(4594) <= b;
    layer3_outputs(4595) <= not (a or b);
    layer3_outputs(4596) <= not (a and b);
    layer3_outputs(4597) <= not a;
    layer3_outputs(4598) <= a or b;
    layer3_outputs(4599) <= a and not b;
    layer3_outputs(4600) <= not (a and b);
    layer3_outputs(4601) <= b and not a;
    layer3_outputs(4602) <= not a;
    layer3_outputs(4603) <= not (a xor b);
    layer3_outputs(4604) <= not a;
    layer3_outputs(4605) <= a xor b;
    layer3_outputs(4606) <= 1'b0;
    layer3_outputs(4607) <= a and b;
    layer3_outputs(4608) <= a;
    layer3_outputs(4609) <= not b or a;
    layer3_outputs(4610) <= not a or b;
    layer3_outputs(4611) <= a and b;
    layer3_outputs(4612) <= not a;
    layer3_outputs(4613) <= not (a or b);
    layer3_outputs(4614) <= a;
    layer3_outputs(4615) <= not (a and b);
    layer3_outputs(4616) <= a xor b;
    layer3_outputs(4617) <= not a or b;
    layer3_outputs(4618) <= not a;
    layer3_outputs(4619) <= a or b;
    layer3_outputs(4620) <= not a;
    layer3_outputs(4621) <= a;
    layer3_outputs(4622) <= b;
    layer3_outputs(4623) <= not a or b;
    layer3_outputs(4624) <= a;
    layer3_outputs(4625) <= not (a and b);
    layer3_outputs(4626) <= not b;
    layer3_outputs(4627) <= 1'b0;
    layer3_outputs(4628) <= not (a or b);
    layer3_outputs(4629) <= a or b;
    layer3_outputs(4630) <= not (a xor b);
    layer3_outputs(4631) <= a and b;
    layer3_outputs(4632) <= not a;
    layer3_outputs(4633) <= not b;
    layer3_outputs(4634) <= b;
    layer3_outputs(4635) <= not (a and b);
    layer3_outputs(4636) <= not (a xor b);
    layer3_outputs(4637) <= not b or a;
    layer3_outputs(4638) <= b;
    layer3_outputs(4639) <= not a;
    layer3_outputs(4640) <= a and b;
    layer3_outputs(4641) <= b;
    layer3_outputs(4642) <= a;
    layer3_outputs(4643) <= a;
    layer3_outputs(4644) <= b;
    layer3_outputs(4645) <= not a;
    layer3_outputs(4646) <= b and not a;
    layer3_outputs(4647) <= b;
    layer3_outputs(4648) <= a xor b;
    layer3_outputs(4649) <= not (a or b);
    layer3_outputs(4650) <= a;
    layer3_outputs(4651) <= a xor b;
    layer3_outputs(4652) <= b;
    layer3_outputs(4653) <= b;
    layer3_outputs(4654) <= not (a or b);
    layer3_outputs(4655) <= a and not b;
    layer3_outputs(4656) <= a;
    layer3_outputs(4657) <= a and b;
    layer3_outputs(4658) <= not (a and b);
    layer3_outputs(4659) <= a xor b;
    layer3_outputs(4660) <= not a;
    layer3_outputs(4661) <= not (a and b);
    layer3_outputs(4662) <= b;
    layer3_outputs(4663) <= not b or a;
    layer3_outputs(4664) <= a or b;
    layer3_outputs(4665) <= a or b;
    layer3_outputs(4666) <= a and b;
    layer3_outputs(4667) <= b;
    layer3_outputs(4668) <= not b;
    layer3_outputs(4669) <= not b;
    layer3_outputs(4670) <= not a;
    layer3_outputs(4671) <= a xor b;
    layer3_outputs(4672) <= a xor b;
    layer3_outputs(4673) <= a;
    layer3_outputs(4674) <= a or b;
    layer3_outputs(4675) <= b;
    layer3_outputs(4676) <= a or b;
    layer3_outputs(4677) <= a and not b;
    layer3_outputs(4678) <= not (a xor b);
    layer3_outputs(4679) <= b;
    layer3_outputs(4680) <= a xor b;
    layer3_outputs(4681) <= not b;
    layer3_outputs(4682) <= b;
    layer3_outputs(4683) <= not a;
    layer3_outputs(4684) <= a or b;
    layer3_outputs(4685) <= 1'b1;
    layer3_outputs(4686) <= not b or a;
    layer3_outputs(4687) <= a and b;
    layer3_outputs(4688) <= a and not b;
    layer3_outputs(4689) <= not (a or b);
    layer3_outputs(4690) <= b;
    layer3_outputs(4691) <= not b;
    layer3_outputs(4692) <= not a;
    layer3_outputs(4693) <= a and b;
    layer3_outputs(4694) <= a;
    layer3_outputs(4695) <= a;
    layer3_outputs(4696) <= not (a or b);
    layer3_outputs(4697) <= a xor b;
    layer3_outputs(4698) <= not b or a;
    layer3_outputs(4699) <= b and not a;
    layer3_outputs(4700) <= not b or a;
    layer3_outputs(4701) <= a;
    layer3_outputs(4702) <= not (a and b);
    layer3_outputs(4703) <= b;
    layer3_outputs(4704) <= not (a xor b);
    layer3_outputs(4705) <= not (a and b);
    layer3_outputs(4706) <= not a or b;
    layer3_outputs(4707) <= not a;
    layer3_outputs(4708) <= not a or b;
    layer3_outputs(4709) <= a;
    layer3_outputs(4710) <= a;
    layer3_outputs(4711) <= not (a and b);
    layer3_outputs(4712) <= a;
    layer3_outputs(4713) <= a;
    layer3_outputs(4714) <= a;
    layer3_outputs(4715) <= not b or a;
    layer3_outputs(4716) <= a and not b;
    layer3_outputs(4717) <= not a;
    layer3_outputs(4718) <= b;
    layer3_outputs(4719) <= not (a and b);
    layer3_outputs(4720) <= a and b;
    layer3_outputs(4721) <= a;
    layer3_outputs(4722) <= a;
    layer3_outputs(4723) <= a;
    layer3_outputs(4724) <= not (a and b);
    layer3_outputs(4725) <= a;
    layer3_outputs(4726) <= not a or b;
    layer3_outputs(4727) <= a and b;
    layer3_outputs(4728) <= b and not a;
    layer3_outputs(4729) <= a;
    layer3_outputs(4730) <= not (a and b);
    layer3_outputs(4731) <= b;
    layer3_outputs(4732) <= not b or a;
    layer3_outputs(4733) <= not b;
    layer3_outputs(4734) <= b;
    layer3_outputs(4735) <= a or b;
    layer3_outputs(4736) <= a or b;
    layer3_outputs(4737) <= not (a and b);
    layer3_outputs(4738) <= not (a and b);
    layer3_outputs(4739) <= a or b;
    layer3_outputs(4740) <= a;
    layer3_outputs(4741) <= a and b;
    layer3_outputs(4742) <= not (a or b);
    layer3_outputs(4743) <= not a;
    layer3_outputs(4744) <= not (a and b);
    layer3_outputs(4745) <= not b;
    layer3_outputs(4746) <= a;
    layer3_outputs(4747) <= b;
    layer3_outputs(4748) <= a and not b;
    layer3_outputs(4749) <= b and not a;
    layer3_outputs(4750) <= not b or a;
    layer3_outputs(4751) <= b and not a;
    layer3_outputs(4752) <= not (a and b);
    layer3_outputs(4753) <= not (a xor b);
    layer3_outputs(4754) <= a or b;
    layer3_outputs(4755) <= not b;
    layer3_outputs(4756) <= b;
    layer3_outputs(4757) <= not (a and b);
    layer3_outputs(4758) <= not b;
    layer3_outputs(4759) <= not b or a;
    layer3_outputs(4760) <= a;
    layer3_outputs(4761) <= not a;
    layer3_outputs(4762) <= a and not b;
    layer3_outputs(4763) <= a;
    layer3_outputs(4764) <= not b or a;
    layer3_outputs(4765) <= not (a and b);
    layer3_outputs(4766) <= not a;
    layer3_outputs(4767) <= a and not b;
    layer3_outputs(4768) <= not (a xor b);
    layer3_outputs(4769) <= a and not b;
    layer3_outputs(4770) <= a and b;
    layer3_outputs(4771) <= not b;
    layer3_outputs(4772) <= b;
    layer3_outputs(4773) <= a and not b;
    layer3_outputs(4774) <= not (a or b);
    layer3_outputs(4775) <= a xor b;
    layer3_outputs(4776) <= not a or b;
    layer3_outputs(4777) <= a xor b;
    layer3_outputs(4778) <= a and b;
    layer3_outputs(4779) <= not (a xor b);
    layer3_outputs(4780) <= b;
    layer3_outputs(4781) <= not b;
    layer3_outputs(4782) <= a xor b;
    layer3_outputs(4783) <= a;
    layer3_outputs(4784) <= not (a xor b);
    layer3_outputs(4785) <= a;
    layer3_outputs(4786) <= a;
    layer3_outputs(4787) <= not a;
    layer3_outputs(4788) <= b;
    layer3_outputs(4789) <= not (a or b);
    layer3_outputs(4790) <= not b;
    layer3_outputs(4791) <= a and b;
    layer3_outputs(4792) <= a or b;
    layer3_outputs(4793) <= a and not b;
    layer3_outputs(4794) <= not (a or b);
    layer3_outputs(4795) <= b and not a;
    layer3_outputs(4796) <= a xor b;
    layer3_outputs(4797) <= a and b;
    layer3_outputs(4798) <= not b;
    layer3_outputs(4799) <= not (a and b);
    layer3_outputs(4800) <= not (a or b);
    layer3_outputs(4801) <= not b;
    layer3_outputs(4802) <= not (a xor b);
    layer3_outputs(4803) <= not a;
    layer3_outputs(4804) <= a;
    layer3_outputs(4805) <= not a;
    layer3_outputs(4806) <= not (a or b);
    layer3_outputs(4807) <= a xor b;
    layer3_outputs(4808) <= b;
    layer3_outputs(4809) <= a;
    layer3_outputs(4810) <= not a or b;
    layer3_outputs(4811) <= not a;
    layer3_outputs(4812) <= b and not a;
    layer3_outputs(4813) <= not b;
    layer3_outputs(4814) <= b;
    layer3_outputs(4815) <= not (a or b);
    layer3_outputs(4816) <= not (a and b);
    layer3_outputs(4817) <= a;
    layer3_outputs(4818) <= b and not a;
    layer3_outputs(4819) <= b;
    layer3_outputs(4820) <= a;
    layer3_outputs(4821) <= a;
    layer3_outputs(4822) <= a and b;
    layer3_outputs(4823) <= not a;
    layer3_outputs(4824) <= not b or a;
    layer3_outputs(4825) <= not a;
    layer3_outputs(4826) <= not a or b;
    layer3_outputs(4827) <= a and not b;
    layer3_outputs(4828) <= not b;
    layer3_outputs(4829) <= not b;
    layer3_outputs(4830) <= not b or a;
    layer3_outputs(4831) <= a;
    layer3_outputs(4832) <= a xor b;
    layer3_outputs(4833) <= not (a xor b);
    layer3_outputs(4834) <= not b;
    layer3_outputs(4835) <= a and b;
    layer3_outputs(4836) <= not (a xor b);
    layer3_outputs(4837) <= a;
    layer3_outputs(4838) <= not a;
    layer3_outputs(4839) <= a;
    layer3_outputs(4840) <= not b or a;
    layer3_outputs(4841) <= b;
    layer3_outputs(4842) <= not a or b;
    layer3_outputs(4843) <= not b;
    layer3_outputs(4844) <= a;
    layer3_outputs(4845) <= b;
    layer3_outputs(4846) <= not (a or b);
    layer3_outputs(4847) <= a or b;
    layer3_outputs(4848) <= not (a and b);
    layer3_outputs(4849) <= a or b;
    layer3_outputs(4850) <= a or b;
    layer3_outputs(4851) <= not (a or b);
    layer3_outputs(4852) <= not b or a;
    layer3_outputs(4853) <= not (a or b);
    layer3_outputs(4854) <= a xor b;
    layer3_outputs(4855) <= b and not a;
    layer3_outputs(4856) <= not a or b;
    layer3_outputs(4857) <= b;
    layer3_outputs(4858) <= a;
    layer3_outputs(4859) <= b and not a;
    layer3_outputs(4860) <= 1'b0;
    layer3_outputs(4861) <= a;
    layer3_outputs(4862) <= not (a and b);
    layer3_outputs(4863) <= a;
    layer3_outputs(4864) <= not (a xor b);
    layer3_outputs(4865) <= not a;
    layer3_outputs(4866) <= a and b;
    layer3_outputs(4867) <= not b or a;
    layer3_outputs(4868) <= not b;
    layer3_outputs(4869) <= not a or b;
    layer3_outputs(4870) <= not (a or b);
    layer3_outputs(4871) <= a and not b;
    layer3_outputs(4872) <= b;
    layer3_outputs(4873) <= b;
    layer3_outputs(4874) <= not a or b;
    layer3_outputs(4875) <= b;
    layer3_outputs(4876) <= a;
    layer3_outputs(4877) <= b;
    layer3_outputs(4878) <= a and not b;
    layer3_outputs(4879) <= b and not a;
    layer3_outputs(4880) <= not (a or b);
    layer3_outputs(4881) <= 1'b1;
    layer3_outputs(4882) <= not b or a;
    layer3_outputs(4883) <= not (a and b);
    layer3_outputs(4884) <= not a or b;
    layer3_outputs(4885) <= not a or b;
    layer3_outputs(4886) <= a or b;
    layer3_outputs(4887) <= a or b;
    layer3_outputs(4888) <= 1'b0;
    layer3_outputs(4889) <= a and not b;
    layer3_outputs(4890) <= not (a or b);
    layer3_outputs(4891) <= b;
    layer3_outputs(4892) <= not a or b;
    layer3_outputs(4893) <= not (a and b);
    layer3_outputs(4894) <= a and b;
    layer3_outputs(4895) <= not b;
    layer3_outputs(4896) <= not b;
    layer3_outputs(4897) <= not (a and b);
    layer3_outputs(4898) <= a and not b;
    layer3_outputs(4899) <= a or b;
    layer3_outputs(4900) <= not b;
    layer3_outputs(4901) <= a;
    layer3_outputs(4902) <= a or b;
    layer3_outputs(4903) <= not (a and b);
    layer3_outputs(4904) <= not (a and b);
    layer3_outputs(4905) <= 1'b1;
    layer3_outputs(4906) <= b;
    layer3_outputs(4907) <= a xor b;
    layer3_outputs(4908) <= not b;
    layer3_outputs(4909) <= b;
    layer3_outputs(4910) <= not (a and b);
    layer3_outputs(4911) <= a;
    layer3_outputs(4912) <= not b;
    layer3_outputs(4913) <= not a;
    layer3_outputs(4914) <= not b;
    layer3_outputs(4915) <= not b or a;
    layer3_outputs(4916) <= not a;
    layer3_outputs(4917) <= not b;
    layer3_outputs(4918) <= not a or b;
    layer3_outputs(4919) <= 1'b1;
    layer3_outputs(4920) <= not b;
    layer3_outputs(4921) <= not (a xor b);
    layer3_outputs(4922) <= b;
    layer3_outputs(4923) <= a and b;
    layer3_outputs(4924) <= not b;
    layer3_outputs(4925) <= not a;
    layer3_outputs(4926) <= not b;
    layer3_outputs(4927) <= not a;
    layer3_outputs(4928) <= not b;
    layer3_outputs(4929) <= a xor b;
    layer3_outputs(4930) <= b;
    layer3_outputs(4931) <= not b or a;
    layer3_outputs(4932) <= not a;
    layer3_outputs(4933) <= a and b;
    layer3_outputs(4934) <= a and not b;
    layer3_outputs(4935) <= b;
    layer3_outputs(4936) <= not b;
    layer3_outputs(4937) <= a;
    layer3_outputs(4938) <= not (a and b);
    layer3_outputs(4939) <= a;
    layer3_outputs(4940) <= not b;
    layer3_outputs(4941) <= not b or a;
    layer3_outputs(4942) <= a or b;
    layer3_outputs(4943) <= not a or b;
    layer3_outputs(4944) <= 1'b1;
    layer3_outputs(4945) <= a and not b;
    layer3_outputs(4946) <= not a or b;
    layer3_outputs(4947) <= not (a and b);
    layer3_outputs(4948) <= not a or b;
    layer3_outputs(4949) <= b;
    layer3_outputs(4950) <= a or b;
    layer3_outputs(4951) <= not a or b;
    layer3_outputs(4952) <= b;
    layer3_outputs(4953) <= not b;
    layer3_outputs(4954) <= a xor b;
    layer3_outputs(4955) <= a or b;
    layer3_outputs(4956) <= a;
    layer3_outputs(4957) <= b;
    layer3_outputs(4958) <= not (a and b);
    layer3_outputs(4959) <= not a or b;
    layer3_outputs(4960) <= a or b;
    layer3_outputs(4961) <= not b;
    layer3_outputs(4962) <= not (a and b);
    layer3_outputs(4963) <= b;
    layer3_outputs(4964) <= not (a or b);
    layer3_outputs(4965) <= a and b;
    layer3_outputs(4966) <= not a;
    layer3_outputs(4967) <= not a or b;
    layer3_outputs(4968) <= not b or a;
    layer3_outputs(4969) <= b;
    layer3_outputs(4970) <= not (a or b);
    layer3_outputs(4971) <= not (a and b);
    layer3_outputs(4972) <= not b;
    layer3_outputs(4973) <= b;
    layer3_outputs(4974) <= not b;
    layer3_outputs(4975) <= not (a or b);
    layer3_outputs(4976) <= not b or a;
    layer3_outputs(4977) <= not (a xor b);
    layer3_outputs(4978) <= not b or a;
    layer3_outputs(4979) <= not b or a;
    layer3_outputs(4980) <= not (a or b);
    layer3_outputs(4981) <= not a;
    layer3_outputs(4982) <= b and not a;
    layer3_outputs(4983) <= not a or b;
    layer3_outputs(4984) <= not a or b;
    layer3_outputs(4985) <= not a or b;
    layer3_outputs(4986) <= not (a or b);
    layer3_outputs(4987) <= not (a and b);
    layer3_outputs(4988) <= b and not a;
    layer3_outputs(4989) <= a and not b;
    layer3_outputs(4990) <= not (a xor b);
    layer3_outputs(4991) <= not (a xor b);
    layer3_outputs(4992) <= not (a and b);
    layer3_outputs(4993) <= not a or b;
    layer3_outputs(4994) <= b;
    layer3_outputs(4995) <= not b;
    layer3_outputs(4996) <= not (a and b);
    layer3_outputs(4997) <= a and not b;
    layer3_outputs(4998) <= not (a and b);
    layer3_outputs(4999) <= not (a or b);
    layer3_outputs(5000) <= b;
    layer3_outputs(5001) <= not (a and b);
    layer3_outputs(5002) <= not (a or b);
    layer3_outputs(5003) <= not b;
    layer3_outputs(5004) <= a xor b;
    layer3_outputs(5005) <= a and not b;
    layer3_outputs(5006) <= not a;
    layer3_outputs(5007) <= a;
    layer3_outputs(5008) <= not a;
    layer3_outputs(5009) <= a and not b;
    layer3_outputs(5010) <= a and not b;
    layer3_outputs(5011) <= not (a and b);
    layer3_outputs(5012) <= not (a and b);
    layer3_outputs(5013) <= a;
    layer3_outputs(5014) <= not (a and b);
    layer3_outputs(5015) <= a;
    layer3_outputs(5016) <= b;
    layer3_outputs(5017) <= 1'b1;
    layer3_outputs(5018) <= b;
    layer3_outputs(5019) <= a xor b;
    layer3_outputs(5020) <= b;
    layer3_outputs(5021) <= not a or b;
    layer3_outputs(5022) <= not b or a;
    layer3_outputs(5023) <= not a;
    layer3_outputs(5024) <= a xor b;
    layer3_outputs(5025) <= b;
    layer3_outputs(5026) <= a and not b;
    layer3_outputs(5027) <= b;
    layer3_outputs(5028) <= not b or a;
    layer3_outputs(5029) <= not b;
    layer3_outputs(5030) <= a;
    layer3_outputs(5031) <= b;
    layer3_outputs(5032) <= a or b;
    layer3_outputs(5033) <= b;
    layer3_outputs(5034) <= a and b;
    layer3_outputs(5035) <= a;
    layer3_outputs(5036) <= b;
    layer3_outputs(5037) <= not b;
    layer3_outputs(5038) <= a or b;
    layer3_outputs(5039) <= b;
    layer3_outputs(5040) <= b;
    layer3_outputs(5041) <= not (a xor b);
    layer3_outputs(5042) <= not (a xor b);
    layer3_outputs(5043) <= a xor b;
    layer3_outputs(5044) <= not a;
    layer3_outputs(5045) <= not (a and b);
    layer3_outputs(5046) <= a;
    layer3_outputs(5047) <= not a;
    layer3_outputs(5048) <= not b or a;
    layer3_outputs(5049) <= not (a or b);
    layer3_outputs(5050) <= not b or a;
    layer3_outputs(5051) <= not b;
    layer3_outputs(5052) <= not (a or b);
    layer3_outputs(5053) <= b;
    layer3_outputs(5054) <= not (a xor b);
    layer3_outputs(5055) <= a and not b;
    layer3_outputs(5056) <= not a;
    layer3_outputs(5057) <= a or b;
    layer3_outputs(5058) <= a xor b;
    layer3_outputs(5059) <= a xor b;
    layer3_outputs(5060) <= not (a xor b);
    layer3_outputs(5061) <= not a or b;
    layer3_outputs(5062) <= a xor b;
    layer3_outputs(5063) <= not b;
    layer3_outputs(5064) <= not a;
    layer3_outputs(5065) <= b;
    layer3_outputs(5066) <= a or b;
    layer3_outputs(5067) <= 1'b0;
    layer3_outputs(5068) <= not b or a;
    layer3_outputs(5069) <= a;
    layer3_outputs(5070) <= a;
    layer3_outputs(5071) <= a;
    layer3_outputs(5072) <= a;
    layer3_outputs(5073) <= a or b;
    layer3_outputs(5074) <= a;
    layer3_outputs(5075) <= not a;
    layer3_outputs(5076) <= 1'b1;
    layer3_outputs(5077) <= not (a and b);
    layer3_outputs(5078) <= a and not b;
    layer3_outputs(5079) <= b;
    layer3_outputs(5080) <= not a;
    layer3_outputs(5081) <= not (a or b);
    layer3_outputs(5082) <= a xor b;
    layer3_outputs(5083) <= not (a or b);
    layer3_outputs(5084) <= not b;
    layer3_outputs(5085) <= a or b;
    layer3_outputs(5086) <= not a or b;
    layer3_outputs(5087) <= a and not b;
    layer3_outputs(5088) <= a xor b;
    layer3_outputs(5089) <= a and b;
    layer3_outputs(5090) <= a;
    layer3_outputs(5091) <= a xor b;
    layer3_outputs(5092) <= not a or b;
    layer3_outputs(5093) <= a xor b;
    layer3_outputs(5094) <= a or b;
    layer3_outputs(5095) <= a and b;
    layer3_outputs(5096) <= a or b;
    layer3_outputs(5097) <= not b;
    layer3_outputs(5098) <= not (a and b);
    layer3_outputs(5099) <= a or b;
    layer3_outputs(5100) <= not a;
    layer3_outputs(5101) <= not a;
    layer3_outputs(5102) <= a;
    layer3_outputs(5103) <= a;
    layer3_outputs(5104) <= b;
    layer3_outputs(5105) <= not (a or b);
    layer3_outputs(5106) <= not a or b;
    layer3_outputs(5107) <= b and not a;
    layer3_outputs(5108) <= not b;
    layer3_outputs(5109) <= a and not b;
    layer3_outputs(5110) <= a and not b;
    layer3_outputs(5111) <= a;
    layer3_outputs(5112) <= a and not b;
    layer3_outputs(5113) <= a and not b;
    layer3_outputs(5114) <= not b;
    layer3_outputs(5115) <= b;
    layer3_outputs(5116) <= not b;
    layer3_outputs(5117) <= a xor b;
    layer3_outputs(5118) <= not b;
    layer3_outputs(5119) <= b;
    layer3_outputs(5120) <= not b;
    layer3_outputs(5121) <= a or b;
    layer3_outputs(5122) <= a;
    layer3_outputs(5123) <= not a;
    layer3_outputs(5124) <= not a;
    layer3_outputs(5125) <= not b;
    layer3_outputs(5126) <= not a;
    layer3_outputs(5127) <= not b or a;
    layer3_outputs(5128) <= a xor b;
    layer3_outputs(5129) <= a;
    layer3_outputs(5130) <= a or b;
    layer3_outputs(5131) <= a or b;
    layer3_outputs(5132) <= not (a xor b);
    layer3_outputs(5133) <= a;
    layer3_outputs(5134) <= not (a xor b);
    layer3_outputs(5135) <= not b;
    layer3_outputs(5136) <= not a;
    layer3_outputs(5137) <= not a;
    layer3_outputs(5138) <= not a;
    layer3_outputs(5139) <= b;
    layer3_outputs(5140) <= a and b;
    layer3_outputs(5141) <= not (a and b);
    layer3_outputs(5142) <= not a or b;
    layer3_outputs(5143) <= not a;
    layer3_outputs(5144) <= b and not a;
    layer3_outputs(5145) <= a;
    layer3_outputs(5146) <= not (a xor b);
    layer3_outputs(5147) <= not b;
    layer3_outputs(5148) <= 1'b1;
    layer3_outputs(5149) <= not a;
    layer3_outputs(5150) <= not (a and b);
    layer3_outputs(5151) <= not a or b;
    layer3_outputs(5152) <= not b;
    layer3_outputs(5153) <= b and not a;
    layer3_outputs(5154) <= a;
    layer3_outputs(5155) <= a and not b;
    layer3_outputs(5156) <= not (a or b);
    layer3_outputs(5157) <= not b;
    layer3_outputs(5158) <= b and not a;
    layer3_outputs(5159) <= not a;
    layer3_outputs(5160) <= a and b;
    layer3_outputs(5161) <= not (a xor b);
    layer3_outputs(5162) <= a;
    layer3_outputs(5163) <= b;
    layer3_outputs(5164) <= a xor b;
    layer3_outputs(5165) <= not a;
    layer3_outputs(5166) <= not b or a;
    layer3_outputs(5167) <= a and b;
    layer3_outputs(5168) <= not (a and b);
    layer3_outputs(5169) <= a xor b;
    layer3_outputs(5170) <= not a;
    layer3_outputs(5171) <= b;
    layer3_outputs(5172) <= a;
    layer3_outputs(5173) <= b;
    layer3_outputs(5174) <= a and b;
    layer3_outputs(5175) <= not b or a;
    layer3_outputs(5176) <= a and b;
    layer3_outputs(5177) <= not b;
    layer3_outputs(5178) <= a xor b;
    layer3_outputs(5179) <= not (a or b);
    layer3_outputs(5180) <= b and not a;
    layer3_outputs(5181) <= not b;
    layer3_outputs(5182) <= not b;
    layer3_outputs(5183) <= not (a or b);
    layer3_outputs(5184) <= b and not a;
    layer3_outputs(5185) <= not b;
    layer3_outputs(5186) <= not a or b;
    layer3_outputs(5187) <= not b;
    layer3_outputs(5188) <= a and b;
    layer3_outputs(5189) <= not b;
    layer3_outputs(5190) <= a;
    layer3_outputs(5191) <= a;
    layer3_outputs(5192) <= 1'b1;
    layer3_outputs(5193) <= not (a xor b);
    layer3_outputs(5194) <= not b;
    layer3_outputs(5195) <= a and b;
    layer3_outputs(5196) <= not a;
    layer3_outputs(5197) <= not a or b;
    layer3_outputs(5198) <= not a or b;
    layer3_outputs(5199) <= b;
    layer3_outputs(5200) <= a;
    layer3_outputs(5201) <= not (a or b);
    layer3_outputs(5202) <= a and b;
    layer3_outputs(5203) <= a or b;
    layer3_outputs(5204) <= not (a or b);
    layer3_outputs(5205) <= not b or a;
    layer3_outputs(5206) <= not b or a;
    layer3_outputs(5207) <= b;
    layer3_outputs(5208) <= not b;
    layer3_outputs(5209) <= b;
    layer3_outputs(5210) <= not b;
    layer3_outputs(5211) <= not b;
    layer3_outputs(5212) <= not (a xor b);
    layer3_outputs(5213) <= b and not a;
    layer3_outputs(5214) <= b and not a;
    layer3_outputs(5215) <= not b or a;
    layer3_outputs(5216) <= a;
    layer3_outputs(5217) <= not a;
    layer3_outputs(5218) <= b and not a;
    layer3_outputs(5219) <= a and not b;
    layer3_outputs(5220) <= not b;
    layer3_outputs(5221) <= a or b;
    layer3_outputs(5222) <= b;
    layer3_outputs(5223) <= not (a xor b);
    layer3_outputs(5224) <= a and not b;
    layer3_outputs(5225) <= a and not b;
    layer3_outputs(5226) <= not a;
    layer3_outputs(5227) <= not (a or b);
    layer3_outputs(5228) <= not b or a;
    layer3_outputs(5229) <= not b or a;
    layer3_outputs(5230) <= a;
    layer3_outputs(5231) <= not b;
    layer3_outputs(5232) <= a;
    layer3_outputs(5233) <= a and b;
    layer3_outputs(5234) <= not b or a;
    layer3_outputs(5235) <= not b;
    layer3_outputs(5236) <= not a or b;
    layer3_outputs(5237) <= a;
    layer3_outputs(5238) <= not a;
    layer3_outputs(5239) <= a xor b;
    layer3_outputs(5240) <= b;
    layer3_outputs(5241) <= a;
    layer3_outputs(5242) <= 1'b0;
    layer3_outputs(5243) <= b and not a;
    layer3_outputs(5244) <= not a or b;
    layer3_outputs(5245) <= not (a or b);
    layer3_outputs(5246) <= not (a or b);
    layer3_outputs(5247) <= b;
    layer3_outputs(5248) <= b;
    layer3_outputs(5249) <= a and not b;
    layer3_outputs(5250) <= a or b;
    layer3_outputs(5251) <= not a;
    layer3_outputs(5252) <= b and not a;
    layer3_outputs(5253) <= not a;
    layer3_outputs(5254) <= not (a and b);
    layer3_outputs(5255) <= b;
    layer3_outputs(5256) <= not b;
    layer3_outputs(5257) <= a;
    layer3_outputs(5258) <= a and not b;
    layer3_outputs(5259) <= b;
    layer3_outputs(5260) <= not (a xor b);
    layer3_outputs(5261) <= b;
    layer3_outputs(5262) <= not (a or b);
    layer3_outputs(5263) <= a;
    layer3_outputs(5264) <= a;
    layer3_outputs(5265) <= a;
    layer3_outputs(5266) <= not (a and b);
    layer3_outputs(5267) <= a and b;
    layer3_outputs(5268) <= a;
    layer3_outputs(5269) <= b;
    layer3_outputs(5270) <= not a or b;
    layer3_outputs(5271) <= b;
    layer3_outputs(5272) <= 1'b1;
    layer3_outputs(5273) <= not (a or b);
    layer3_outputs(5274) <= not b;
    layer3_outputs(5275) <= a xor b;
    layer3_outputs(5276) <= b;
    layer3_outputs(5277) <= b;
    layer3_outputs(5278) <= not b;
    layer3_outputs(5279) <= a xor b;
    layer3_outputs(5280) <= not a;
    layer3_outputs(5281) <= a xor b;
    layer3_outputs(5282) <= b and not a;
    layer3_outputs(5283) <= b;
    layer3_outputs(5284) <= b;
    layer3_outputs(5285) <= a;
    layer3_outputs(5286) <= b and not a;
    layer3_outputs(5287) <= a and b;
    layer3_outputs(5288) <= a;
    layer3_outputs(5289) <= not (a or b);
    layer3_outputs(5290) <= not (a xor b);
    layer3_outputs(5291) <= not b;
    layer3_outputs(5292) <= not (a or b);
    layer3_outputs(5293) <= not a;
    layer3_outputs(5294) <= not (a and b);
    layer3_outputs(5295) <= a or b;
    layer3_outputs(5296) <= b;
    layer3_outputs(5297) <= a;
    layer3_outputs(5298) <= not b;
    layer3_outputs(5299) <= not b;
    layer3_outputs(5300) <= a and not b;
    layer3_outputs(5301) <= b;
    layer3_outputs(5302) <= not a or b;
    layer3_outputs(5303) <= a xor b;
    layer3_outputs(5304) <= not a;
    layer3_outputs(5305) <= not b;
    layer3_outputs(5306) <= not b;
    layer3_outputs(5307) <= a and b;
    layer3_outputs(5308) <= a xor b;
    layer3_outputs(5309) <= a and b;
    layer3_outputs(5310) <= not (a xor b);
    layer3_outputs(5311) <= not a or b;
    layer3_outputs(5312) <= a and not b;
    layer3_outputs(5313) <= a;
    layer3_outputs(5314) <= not (a or b);
    layer3_outputs(5315) <= not a or b;
    layer3_outputs(5316) <= a;
    layer3_outputs(5317) <= not a;
    layer3_outputs(5318) <= a;
    layer3_outputs(5319) <= a or b;
    layer3_outputs(5320) <= b;
    layer3_outputs(5321) <= not b or a;
    layer3_outputs(5322) <= not a or b;
    layer3_outputs(5323) <= not b;
    layer3_outputs(5324) <= a;
    layer3_outputs(5325) <= not a;
    layer3_outputs(5326) <= a xor b;
    layer3_outputs(5327) <= b and not a;
    layer3_outputs(5328) <= not (a and b);
    layer3_outputs(5329) <= a;
    layer3_outputs(5330) <= b;
    layer3_outputs(5331) <= a xor b;
    layer3_outputs(5332) <= not (a and b);
    layer3_outputs(5333) <= not a or b;
    layer3_outputs(5334) <= not b or a;
    layer3_outputs(5335) <= not b;
    layer3_outputs(5336) <= a and not b;
    layer3_outputs(5337) <= a and b;
    layer3_outputs(5338) <= not a;
    layer3_outputs(5339) <= a;
    layer3_outputs(5340) <= not a;
    layer3_outputs(5341) <= a and b;
    layer3_outputs(5342) <= a and not b;
    layer3_outputs(5343) <= a;
    layer3_outputs(5344) <= a xor b;
    layer3_outputs(5345) <= not b or a;
    layer3_outputs(5346) <= b;
    layer3_outputs(5347) <= a and not b;
    layer3_outputs(5348) <= a xor b;
    layer3_outputs(5349) <= a and b;
    layer3_outputs(5350) <= not b;
    layer3_outputs(5351) <= not (a and b);
    layer3_outputs(5352) <= a or b;
    layer3_outputs(5353) <= b;
    layer3_outputs(5354) <= not a;
    layer3_outputs(5355) <= not b or a;
    layer3_outputs(5356) <= not (a or b);
    layer3_outputs(5357) <= a and not b;
    layer3_outputs(5358) <= a and b;
    layer3_outputs(5359) <= not (a and b);
    layer3_outputs(5360) <= a or b;
    layer3_outputs(5361) <= not a or b;
    layer3_outputs(5362) <= not (a or b);
    layer3_outputs(5363) <= b;
    layer3_outputs(5364) <= b;
    layer3_outputs(5365) <= not b;
    layer3_outputs(5366) <= b;
    layer3_outputs(5367) <= b;
    layer3_outputs(5368) <= not (a or b);
    layer3_outputs(5369) <= not (a xor b);
    layer3_outputs(5370) <= a or b;
    layer3_outputs(5371) <= not (a or b);
    layer3_outputs(5372) <= not b;
    layer3_outputs(5373) <= b and not a;
    layer3_outputs(5374) <= a;
    layer3_outputs(5375) <= not a;
    layer3_outputs(5376) <= not a or b;
    layer3_outputs(5377) <= not (a xor b);
    layer3_outputs(5378) <= a;
    layer3_outputs(5379) <= not b or a;
    layer3_outputs(5380) <= a and b;
    layer3_outputs(5381) <= not a or b;
    layer3_outputs(5382) <= a;
    layer3_outputs(5383) <= not (a and b);
    layer3_outputs(5384) <= a and b;
    layer3_outputs(5385) <= not a;
    layer3_outputs(5386) <= a;
    layer3_outputs(5387) <= not b;
    layer3_outputs(5388) <= not a or b;
    layer3_outputs(5389) <= a or b;
    layer3_outputs(5390) <= not a or b;
    layer3_outputs(5391) <= not (a or b);
    layer3_outputs(5392) <= a xor b;
    layer3_outputs(5393) <= not a;
    layer3_outputs(5394) <= not b;
    layer3_outputs(5395) <= 1'b0;
    layer3_outputs(5396) <= not a;
    layer3_outputs(5397) <= not a;
    layer3_outputs(5398) <= not b;
    layer3_outputs(5399) <= a xor b;
    layer3_outputs(5400) <= 1'b0;
    layer3_outputs(5401) <= b;
    layer3_outputs(5402) <= b and not a;
    layer3_outputs(5403) <= b;
    layer3_outputs(5404) <= not a or b;
    layer3_outputs(5405) <= not (a or b);
    layer3_outputs(5406) <= not a;
    layer3_outputs(5407) <= not b;
    layer3_outputs(5408) <= not b or a;
    layer3_outputs(5409) <= a and not b;
    layer3_outputs(5410) <= b;
    layer3_outputs(5411) <= b;
    layer3_outputs(5412) <= a;
    layer3_outputs(5413) <= a and b;
    layer3_outputs(5414) <= not b or a;
    layer3_outputs(5415) <= not b;
    layer3_outputs(5416) <= not (a xor b);
    layer3_outputs(5417) <= not a;
    layer3_outputs(5418) <= a and not b;
    layer3_outputs(5419) <= a xor b;
    layer3_outputs(5420) <= 1'b1;
    layer3_outputs(5421) <= not b or a;
    layer3_outputs(5422) <= not b;
    layer3_outputs(5423) <= not b or a;
    layer3_outputs(5424) <= b;
    layer3_outputs(5425) <= b;
    layer3_outputs(5426) <= b;
    layer3_outputs(5427) <= a or b;
    layer3_outputs(5428) <= a and b;
    layer3_outputs(5429) <= not a;
    layer3_outputs(5430) <= not b;
    layer3_outputs(5431) <= not a;
    layer3_outputs(5432) <= not a or b;
    layer3_outputs(5433) <= not a or b;
    layer3_outputs(5434) <= b and not a;
    layer3_outputs(5435) <= not (a xor b);
    layer3_outputs(5436) <= a and b;
    layer3_outputs(5437) <= a;
    layer3_outputs(5438) <= a or b;
    layer3_outputs(5439) <= not b;
    layer3_outputs(5440) <= not (a xor b);
    layer3_outputs(5441) <= not (a and b);
    layer3_outputs(5442) <= not b;
    layer3_outputs(5443) <= not (a or b);
    layer3_outputs(5444) <= b;
    layer3_outputs(5445) <= a;
    layer3_outputs(5446) <= 1'b1;
    layer3_outputs(5447) <= not a;
    layer3_outputs(5448) <= b;
    layer3_outputs(5449) <= not b;
    layer3_outputs(5450) <= a;
    layer3_outputs(5451) <= not (a and b);
    layer3_outputs(5452) <= a;
    layer3_outputs(5453) <= a and b;
    layer3_outputs(5454) <= a xor b;
    layer3_outputs(5455) <= not b or a;
    layer3_outputs(5456) <= not (a xor b);
    layer3_outputs(5457) <= not b;
    layer3_outputs(5458) <= a xor b;
    layer3_outputs(5459) <= a;
    layer3_outputs(5460) <= a and b;
    layer3_outputs(5461) <= not b or a;
    layer3_outputs(5462) <= a and b;
    layer3_outputs(5463) <= not (a and b);
    layer3_outputs(5464) <= a or b;
    layer3_outputs(5465) <= 1'b0;
    layer3_outputs(5466) <= a;
    layer3_outputs(5467) <= not a;
    layer3_outputs(5468) <= a or b;
    layer3_outputs(5469) <= not a;
    layer3_outputs(5470) <= a and not b;
    layer3_outputs(5471) <= a and b;
    layer3_outputs(5472) <= b and not a;
    layer3_outputs(5473) <= a xor b;
    layer3_outputs(5474) <= a or b;
    layer3_outputs(5475) <= a xor b;
    layer3_outputs(5476) <= a and b;
    layer3_outputs(5477) <= not b or a;
    layer3_outputs(5478) <= not a;
    layer3_outputs(5479) <= b;
    layer3_outputs(5480) <= b;
    layer3_outputs(5481) <= b;
    layer3_outputs(5482) <= a and not b;
    layer3_outputs(5483) <= a;
    layer3_outputs(5484) <= a and not b;
    layer3_outputs(5485) <= b and not a;
    layer3_outputs(5486) <= not a;
    layer3_outputs(5487) <= not (a xor b);
    layer3_outputs(5488) <= b;
    layer3_outputs(5489) <= a xor b;
    layer3_outputs(5490) <= not a or b;
    layer3_outputs(5491) <= a and not b;
    layer3_outputs(5492) <= b;
    layer3_outputs(5493) <= a xor b;
    layer3_outputs(5494) <= b;
    layer3_outputs(5495) <= a xor b;
    layer3_outputs(5496) <= not b;
    layer3_outputs(5497) <= not (a xor b);
    layer3_outputs(5498) <= 1'b0;
    layer3_outputs(5499) <= a;
    layer3_outputs(5500) <= not a or b;
    layer3_outputs(5501) <= not a or b;
    layer3_outputs(5502) <= not a;
    layer3_outputs(5503) <= b;
    layer3_outputs(5504) <= a or b;
    layer3_outputs(5505) <= not b;
    layer3_outputs(5506) <= not (a xor b);
    layer3_outputs(5507) <= a and b;
    layer3_outputs(5508) <= not a;
    layer3_outputs(5509) <= not b;
    layer3_outputs(5510) <= not b;
    layer3_outputs(5511) <= not a;
    layer3_outputs(5512) <= a xor b;
    layer3_outputs(5513) <= 1'b0;
    layer3_outputs(5514) <= a;
    layer3_outputs(5515) <= b;
    layer3_outputs(5516) <= not (a and b);
    layer3_outputs(5517) <= not b or a;
    layer3_outputs(5518) <= not a;
    layer3_outputs(5519) <= not (a or b);
    layer3_outputs(5520) <= not (a or b);
    layer3_outputs(5521) <= not b;
    layer3_outputs(5522) <= not b;
    layer3_outputs(5523) <= a;
    layer3_outputs(5524) <= a;
    layer3_outputs(5525) <= a;
    layer3_outputs(5526) <= not (a and b);
    layer3_outputs(5527) <= a and not b;
    layer3_outputs(5528) <= not b;
    layer3_outputs(5529) <= a;
    layer3_outputs(5530) <= not a;
    layer3_outputs(5531) <= not a;
    layer3_outputs(5532) <= not b or a;
    layer3_outputs(5533) <= a or b;
    layer3_outputs(5534) <= not a or b;
    layer3_outputs(5535) <= a xor b;
    layer3_outputs(5536) <= not (a or b);
    layer3_outputs(5537) <= a and not b;
    layer3_outputs(5538) <= a or b;
    layer3_outputs(5539) <= b;
    layer3_outputs(5540) <= not (a or b);
    layer3_outputs(5541) <= b;
    layer3_outputs(5542) <= not a;
    layer3_outputs(5543) <= a;
    layer3_outputs(5544) <= not b or a;
    layer3_outputs(5545) <= b;
    layer3_outputs(5546) <= b and not a;
    layer3_outputs(5547) <= not (a and b);
    layer3_outputs(5548) <= a or b;
    layer3_outputs(5549) <= a xor b;
    layer3_outputs(5550) <= not a or b;
    layer3_outputs(5551) <= a;
    layer3_outputs(5552) <= not b;
    layer3_outputs(5553) <= not a;
    layer3_outputs(5554) <= a and b;
    layer3_outputs(5555) <= not a;
    layer3_outputs(5556) <= not a or b;
    layer3_outputs(5557) <= not a or b;
    layer3_outputs(5558) <= not a;
    layer3_outputs(5559) <= a;
    layer3_outputs(5560) <= a xor b;
    layer3_outputs(5561) <= not a;
    layer3_outputs(5562) <= not b;
    layer3_outputs(5563) <= not (a xor b);
    layer3_outputs(5564) <= not (a xor b);
    layer3_outputs(5565) <= not (a and b);
    layer3_outputs(5566) <= not a;
    layer3_outputs(5567) <= b;
    layer3_outputs(5568) <= not b;
    layer3_outputs(5569) <= a xor b;
    layer3_outputs(5570) <= not b;
    layer3_outputs(5571) <= not a or b;
    layer3_outputs(5572) <= b;
    layer3_outputs(5573) <= not a;
    layer3_outputs(5574) <= a and not b;
    layer3_outputs(5575) <= not a;
    layer3_outputs(5576) <= not b or a;
    layer3_outputs(5577) <= not (a and b);
    layer3_outputs(5578) <= not a;
    layer3_outputs(5579) <= not b or a;
    layer3_outputs(5580) <= not b;
    layer3_outputs(5581) <= a;
    layer3_outputs(5582) <= b and not a;
    layer3_outputs(5583) <= not b;
    layer3_outputs(5584) <= 1'b0;
    layer3_outputs(5585) <= not a or b;
    layer3_outputs(5586) <= b;
    layer3_outputs(5587) <= a xor b;
    layer3_outputs(5588) <= not b or a;
    layer3_outputs(5589) <= 1'b1;
    layer3_outputs(5590) <= a and b;
    layer3_outputs(5591) <= not b;
    layer3_outputs(5592) <= not b;
    layer3_outputs(5593) <= a;
    layer3_outputs(5594) <= a xor b;
    layer3_outputs(5595) <= a xor b;
    layer3_outputs(5596) <= b;
    layer3_outputs(5597) <= b and not a;
    layer3_outputs(5598) <= a;
    layer3_outputs(5599) <= not (a or b);
    layer3_outputs(5600) <= not b;
    layer3_outputs(5601) <= a;
    layer3_outputs(5602) <= a xor b;
    layer3_outputs(5603) <= a or b;
    layer3_outputs(5604) <= a and not b;
    layer3_outputs(5605) <= a xor b;
    layer3_outputs(5606) <= a xor b;
    layer3_outputs(5607) <= not b;
    layer3_outputs(5608) <= 1'b1;
    layer3_outputs(5609) <= not b or a;
    layer3_outputs(5610) <= a or b;
    layer3_outputs(5611) <= not (a xor b);
    layer3_outputs(5612) <= b;
    layer3_outputs(5613) <= not b or a;
    layer3_outputs(5614) <= not a or b;
    layer3_outputs(5615) <= b;
    layer3_outputs(5616) <= a and b;
    layer3_outputs(5617) <= a;
    layer3_outputs(5618) <= not a;
    layer3_outputs(5619) <= a and b;
    layer3_outputs(5620) <= b;
    layer3_outputs(5621) <= a or b;
    layer3_outputs(5622) <= 1'b0;
    layer3_outputs(5623) <= not a or b;
    layer3_outputs(5624) <= not a;
    layer3_outputs(5625) <= a;
    layer3_outputs(5626) <= 1'b1;
    layer3_outputs(5627) <= b and not a;
    layer3_outputs(5628) <= not (a and b);
    layer3_outputs(5629) <= not a;
    layer3_outputs(5630) <= not (a xor b);
    layer3_outputs(5631) <= not a;
    layer3_outputs(5632) <= b and not a;
    layer3_outputs(5633) <= not b;
    layer3_outputs(5634) <= b;
    layer3_outputs(5635) <= not a;
    layer3_outputs(5636) <= a and b;
    layer3_outputs(5637) <= a and not b;
    layer3_outputs(5638) <= not a;
    layer3_outputs(5639) <= not (a and b);
    layer3_outputs(5640) <= not b or a;
    layer3_outputs(5641) <= not a;
    layer3_outputs(5642) <= not a or b;
    layer3_outputs(5643) <= b;
    layer3_outputs(5644) <= not b;
    layer3_outputs(5645) <= not (a xor b);
    layer3_outputs(5646) <= a or b;
    layer3_outputs(5647) <= not (a xor b);
    layer3_outputs(5648) <= a or b;
    layer3_outputs(5649) <= not b;
    layer3_outputs(5650) <= not (a xor b);
    layer3_outputs(5651) <= not (a xor b);
    layer3_outputs(5652) <= not (a xor b);
    layer3_outputs(5653) <= not a or b;
    layer3_outputs(5654) <= 1'b1;
    layer3_outputs(5655) <= not a;
    layer3_outputs(5656) <= b and not a;
    layer3_outputs(5657) <= a or b;
    layer3_outputs(5658) <= not (a xor b);
    layer3_outputs(5659) <= not b;
    layer3_outputs(5660) <= not b;
    layer3_outputs(5661) <= b;
    layer3_outputs(5662) <= not (a or b);
    layer3_outputs(5663) <= not (a xor b);
    layer3_outputs(5664) <= a xor b;
    layer3_outputs(5665) <= b;
    layer3_outputs(5666) <= not (a and b);
    layer3_outputs(5667) <= not a or b;
    layer3_outputs(5668) <= not (a or b);
    layer3_outputs(5669) <= a;
    layer3_outputs(5670) <= a;
    layer3_outputs(5671) <= not (a and b);
    layer3_outputs(5672) <= not a;
    layer3_outputs(5673) <= b;
    layer3_outputs(5674) <= not a;
    layer3_outputs(5675) <= not a;
    layer3_outputs(5676) <= not a or b;
    layer3_outputs(5677) <= not (a xor b);
    layer3_outputs(5678) <= not b;
    layer3_outputs(5679) <= a and not b;
    layer3_outputs(5680) <= not (a or b);
    layer3_outputs(5681) <= a;
    layer3_outputs(5682) <= 1'b1;
    layer3_outputs(5683) <= a xor b;
    layer3_outputs(5684) <= b;
    layer3_outputs(5685) <= a;
    layer3_outputs(5686) <= a;
    layer3_outputs(5687) <= not b;
    layer3_outputs(5688) <= b;
    layer3_outputs(5689) <= b;
    layer3_outputs(5690) <= not b or a;
    layer3_outputs(5691) <= not (a or b);
    layer3_outputs(5692) <= not (a or b);
    layer3_outputs(5693) <= not (a and b);
    layer3_outputs(5694) <= b;
    layer3_outputs(5695) <= 1'b0;
    layer3_outputs(5696) <= not (a and b);
    layer3_outputs(5697) <= not b or a;
    layer3_outputs(5698) <= a and b;
    layer3_outputs(5699) <= a;
    layer3_outputs(5700) <= a;
    layer3_outputs(5701) <= not a;
    layer3_outputs(5702) <= a;
    layer3_outputs(5703) <= a and b;
    layer3_outputs(5704) <= not (a and b);
    layer3_outputs(5705) <= not (a or b);
    layer3_outputs(5706) <= a and b;
    layer3_outputs(5707) <= a;
    layer3_outputs(5708) <= b and not a;
    layer3_outputs(5709) <= a xor b;
    layer3_outputs(5710) <= a and not b;
    layer3_outputs(5711) <= a and b;
    layer3_outputs(5712) <= not b;
    layer3_outputs(5713) <= a or b;
    layer3_outputs(5714) <= a;
    layer3_outputs(5715) <= a xor b;
    layer3_outputs(5716) <= a or b;
    layer3_outputs(5717) <= not b;
    layer3_outputs(5718) <= not b;
    layer3_outputs(5719) <= a xor b;
    layer3_outputs(5720) <= b and not a;
    layer3_outputs(5721) <= a or b;
    layer3_outputs(5722) <= not a or b;
    layer3_outputs(5723) <= b;
    layer3_outputs(5724) <= not a;
    layer3_outputs(5725) <= not b;
    layer3_outputs(5726) <= a xor b;
    layer3_outputs(5727) <= b and not a;
    layer3_outputs(5728) <= a and not b;
    layer3_outputs(5729) <= a or b;
    layer3_outputs(5730) <= not a;
    layer3_outputs(5731) <= not (a xor b);
    layer3_outputs(5732) <= 1'b1;
    layer3_outputs(5733) <= not a;
    layer3_outputs(5734) <= b and not a;
    layer3_outputs(5735) <= a;
    layer3_outputs(5736) <= not b or a;
    layer3_outputs(5737) <= a;
    layer3_outputs(5738) <= a and not b;
    layer3_outputs(5739) <= not (a xor b);
    layer3_outputs(5740) <= not a or b;
    layer3_outputs(5741) <= not b;
    layer3_outputs(5742) <= not (a and b);
    layer3_outputs(5743) <= not (a or b);
    layer3_outputs(5744) <= b;
    layer3_outputs(5745) <= not (a xor b);
    layer3_outputs(5746) <= a and b;
    layer3_outputs(5747) <= b and not a;
    layer3_outputs(5748) <= not a or b;
    layer3_outputs(5749) <= not (a xor b);
    layer3_outputs(5750) <= not (a xor b);
    layer3_outputs(5751) <= not b or a;
    layer3_outputs(5752) <= not (a and b);
    layer3_outputs(5753) <= b and not a;
    layer3_outputs(5754) <= b;
    layer3_outputs(5755) <= not b;
    layer3_outputs(5756) <= a and b;
    layer3_outputs(5757) <= not b;
    layer3_outputs(5758) <= a and not b;
    layer3_outputs(5759) <= not b;
    layer3_outputs(5760) <= not a or b;
    layer3_outputs(5761) <= a and not b;
    layer3_outputs(5762) <= a xor b;
    layer3_outputs(5763) <= not a;
    layer3_outputs(5764) <= a;
    layer3_outputs(5765) <= b;
    layer3_outputs(5766) <= not (a or b);
    layer3_outputs(5767) <= 1'b1;
    layer3_outputs(5768) <= a;
    layer3_outputs(5769) <= a;
    layer3_outputs(5770) <= not a or b;
    layer3_outputs(5771) <= a;
    layer3_outputs(5772) <= a;
    layer3_outputs(5773) <= b;
    layer3_outputs(5774) <= b;
    layer3_outputs(5775) <= not a;
    layer3_outputs(5776) <= a and not b;
    layer3_outputs(5777) <= a and not b;
    layer3_outputs(5778) <= b and not a;
    layer3_outputs(5779) <= b;
    layer3_outputs(5780) <= not b;
    layer3_outputs(5781) <= not (a or b);
    layer3_outputs(5782) <= a and not b;
    layer3_outputs(5783) <= a and b;
    layer3_outputs(5784) <= a and not b;
    layer3_outputs(5785) <= a and b;
    layer3_outputs(5786) <= a xor b;
    layer3_outputs(5787) <= not b;
    layer3_outputs(5788) <= a;
    layer3_outputs(5789) <= not (a or b);
    layer3_outputs(5790) <= b;
    layer3_outputs(5791) <= a;
    layer3_outputs(5792) <= b;
    layer3_outputs(5793) <= not (a or b);
    layer3_outputs(5794) <= b;
    layer3_outputs(5795) <= not (a or b);
    layer3_outputs(5796) <= a;
    layer3_outputs(5797) <= a and not b;
    layer3_outputs(5798) <= a and b;
    layer3_outputs(5799) <= not (a and b);
    layer3_outputs(5800) <= not a;
    layer3_outputs(5801) <= not b or a;
    layer3_outputs(5802) <= a;
    layer3_outputs(5803) <= not a;
    layer3_outputs(5804) <= not (a or b);
    layer3_outputs(5805) <= not b or a;
    layer3_outputs(5806) <= not a or b;
    layer3_outputs(5807) <= not b;
    layer3_outputs(5808) <= not a or b;
    layer3_outputs(5809) <= b;
    layer3_outputs(5810) <= a and b;
    layer3_outputs(5811) <= not (a and b);
    layer3_outputs(5812) <= not (a and b);
    layer3_outputs(5813) <= not (a and b);
    layer3_outputs(5814) <= a;
    layer3_outputs(5815) <= b;
    layer3_outputs(5816) <= not b or a;
    layer3_outputs(5817) <= a;
    layer3_outputs(5818) <= not (a or b);
    layer3_outputs(5819) <= not b or a;
    layer3_outputs(5820) <= a and not b;
    layer3_outputs(5821) <= a or b;
    layer3_outputs(5822) <= a and b;
    layer3_outputs(5823) <= not a or b;
    layer3_outputs(5824) <= not b;
    layer3_outputs(5825) <= not (a xor b);
    layer3_outputs(5826) <= not (a and b);
    layer3_outputs(5827) <= a;
    layer3_outputs(5828) <= not b;
    layer3_outputs(5829) <= a xor b;
    layer3_outputs(5830) <= not (a or b);
    layer3_outputs(5831) <= a;
    layer3_outputs(5832) <= a;
    layer3_outputs(5833) <= not b;
    layer3_outputs(5834) <= not a;
    layer3_outputs(5835) <= 1'b0;
    layer3_outputs(5836) <= 1'b1;
    layer3_outputs(5837) <= a xor b;
    layer3_outputs(5838) <= not a;
    layer3_outputs(5839) <= a and b;
    layer3_outputs(5840) <= a and not b;
    layer3_outputs(5841) <= not a;
    layer3_outputs(5842) <= not b or a;
    layer3_outputs(5843) <= 1'b1;
    layer3_outputs(5844) <= not b;
    layer3_outputs(5845) <= not b;
    layer3_outputs(5846) <= b and not a;
    layer3_outputs(5847) <= a and b;
    layer3_outputs(5848) <= a;
    layer3_outputs(5849) <= not (a or b);
    layer3_outputs(5850) <= a xor b;
    layer3_outputs(5851) <= not (a or b);
    layer3_outputs(5852) <= not a;
    layer3_outputs(5853) <= b;
    layer3_outputs(5854) <= not (a xor b);
    layer3_outputs(5855) <= a and not b;
    layer3_outputs(5856) <= not b;
    layer3_outputs(5857) <= not a;
    layer3_outputs(5858) <= a and b;
    layer3_outputs(5859) <= a or b;
    layer3_outputs(5860) <= not b;
    layer3_outputs(5861) <= a xor b;
    layer3_outputs(5862) <= a and not b;
    layer3_outputs(5863) <= not b;
    layer3_outputs(5864) <= a and not b;
    layer3_outputs(5865) <= not b;
    layer3_outputs(5866) <= not b;
    layer3_outputs(5867) <= not b or a;
    layer3_outputs(5868) <= not (a and b);
    layer3_outputs(5869) <= b;
    layer3_outputs(5870) <= a xor b;
    layer3_outputs(5871) <= b;
    layer3_outputs(5872) <= a or b;
    layer3_outputs(5873) <= a xor b;
    layer3_outputs(5874) <= not (a xor b);
    layer3_outputs(5875) <= not a;
    layer3_outputs(5876) <= not b;
    layer3_outputs(5877) <= b;
    layer3_outputs(5878) <= not b or a;
    layer3_outputs(5879) <= a;
    layer3_outputs(5880) <= a;
    layer3_outputs(5881) <= not a or b;
    layer3_outputs(5882) <= a and not b;
    layer3_outputs(5883) <= b;
    layer3_outputs(5884) <= b;
    layer3_outputs(5885) <= a xor b;
    layer3_outputs(5886) <= not b;
    layer3_outputs(5887) <= a xor b;
    layer3_outputs(5888) <= not a;
    layer3_outputs(5889) <= b;
    layer3_outputs(5890) <= a or b;
    layer3_outputs(5891) <= not a or b;
    layer3_outputs(5892) <= not b or a;
    layer3_outputs(5893) <= b;
    layer3_outputs(5894) <= not b;
    layer3_outputs(5895) <= a and not b;
    layer3_outputs(5896) <= not b;
    layer3_outputs(5897) <= a and b;
    layer3_outputs(5898) <= a or b;
    layer3_outputs(5899) <= a;
    layer3_outputs(5900) <= not b or a;
    layer3_outputs(5901) <= a and b;
    layer3_outputs(5902) <= a or b;
    layer3_outputs(5903) <= not b;
    layer3_outputs(5904) <= a;
    layer3_outputs(5905) <= a;
    layer3_outputs(5906) <= a or b;
    layer3_outputs(5907) <= not (a or b);
    layer3_outputs(5908) <= not b or a;
    layer3_outputs(5909) <= a and not b;
    layer3_outputs(5910) <= not (a or b);
    layer3_outputs(5911) <= not b;
    layer3_outputs(5912) <= not a or b;
    layer3_outputs(5913) <= not (a or b);
    layer3_outputs(5914) <= not a;
    layer3_outputs(5915) <= not a or b;
    layer3_outputs(5916) <= not a or b;
    layer3_outputs(5917) <= not b;
    layer3_outputs(5918) <= not (a xor b);
    layer3_outputs(5919) <= not b;
    layer3_outputs(5920) <= a or b;
    layer3_outputs(5921) <= a xor b;
    layer3_outputs(5922) <= not b or a;
    layer3_outputs(5923) <= not a;
    layer3_outputs(5924) <= a and not b;
    layer3_outputs(5925) <= a xor b;
    layer3_outputs(5926) <= not (a and b);
    layer3_outputs(5927) <= b and not a;
    layer3_outputs(5928) <= not (a xor b);
    layer3_outputs(5929) <= not a;
    layer3_outputs(5930) <= not (a and b);
    layer3_outputs(5931) <= a xor b;
    layer3_outputs(5932) <= not (a and b);
    layer3_outputs(5933) <= a and not b;
    layer3_outputs(5934) <= b;
    layer3_outputs(5935) <= a xor b;
    layer3_outputs(5936) <= not b;
    layer3_outputs(5937) <= a;
    layer3_outputs(5938) <= not (a or b);
    layer3_outputs(5939) <= b;
    layer3_outputs(5940) <= b;
    layer3_outputs(5941) <= b;
    layer3_outputs(5942) <= a;
    layer3_outputs(5943) <= not a;
    layer3_outputs(5944) <= not b;
    layer3_outputs(5945) <= not a or b;
    layer3_outputs(5946) <= a;
    layer3_outputs(5947) <= a and not b;
    layer3_outputs(5948) <= a xor b;
    layer3_outputs(5949) <= 1'b1;
    layer3_outputs(5950) <= a or b;
    layer3_outputs(5951) <= a and not b;
    layer3_outputs(5952) <= a xor b;
    layer3_outputs(5953) <= a or b;
    layer3_outputs(5954) <= b;
    layer3_outputs(5955) <= a;
    layer3_outputs(5956) <= not b;
    layer3_outputs(5957) <= not a;
    layer3_outputs(5958) <= not b or a;
    layer3_outputs(5959) <= a;
    layer3_outputs(5960) <= not b;
    layer3_outputs(5961) <= a xor b;
    layer3_outputs(5962) <= not a;
    layer3_outputs(5963) <= b;
    layer3_outputs(5964) <= not (a xor b);
    layer3_outputs(5965) <= not b;
    layer3_outputs(5966) <= not b;
    layer3_outputs(5967) <= not b;
    layer3_outputs(5968) <= not b;
    layer3_outputs(5969) <= not (a xor b);
    layer3_outputs(5970) <= b;
    layer3_outputs(5971) <= b and not a;
    layer3_outputs(5972) <= a and not b;
    layer3_outputs(5973) <= a and b;
    layer3_outputs(5974) <= a or b;
    layer3_outputs(5975) <= b and not a;
    layer3_outputs(5976) <= not b;
    layer3_outputs(5977) <= a xor b;
    layer3_outputs(5978) <= b;
    layer3_outputs(5979) <= not b or a;
    layer3_outputs(5980) <= not b or a;
    layer3_outputs(5981) <= not b;
    layer3_outputs(5982) <= not b;
    layer3_outputs(5983) <= not a or b;
    layer3_outputs(5984) <= not b or a;
    layer3_outputs(5985) <= not b or a;
    layer3_outputs(5986) <= not (a xor b);
    layer3_outputs(5987) <= a;
    layer3_outputs(5988) <= not (a and b);
    layer3_outputs(5989) <= not b or a;
    layer3_outputs(5990) <= not (a xor b);
    layer3_outputs(5991) <= not a;
    layer3_outputs(5992) <= not b or a;
    layer3_outputs(5993) <= not b or a;
    layer3_outputs(5994) <= b;
    layer3_outputs(5995) <= a;
    layer3_outputs(5996) <= a and not b;
    layer3_outputs(5997) <= a and not b;
    layer3_outputs(5998) <= not (a or b);
    layer3_outputs(5999) <= not b or a;
    layer3_outputs(6000) <= b;
    layer3_outputs(6001) <= not a;
    layer3_outputs(6002) <= b and not a;
    layer3_outputs(6003) <= a xor b;
    layer3_outputs(6004) <= b and not a;
    layer3_outputs(6005) <= a and b;
    layer3_outputs(6006) <= a;
    layer3_outputs(6007) <= a and not b;
    layer3_outputs(6008) <= not a;
    layer3_outputs(6009) <= not b;
    layer3_outputs(6010) <= a or b;
    layer3_outputs(6011) <= not (a and b);
    layer3_outputs(6012) <= not (a or b);
    layer3_outputs(6013) <= not b;
    layer3_outputs(6014) <= b;
    layer3_outputs(6015) <= b and not a;
    layer3_outputs(6016) <= a;
    layer3_outputs(6017) <= not a;
    layer3_outputs(6018) <= not a;
    layer3_outputs(6019) <= not b or a;
    layer3_outputs(6020) <= not a;
    layer3_outputs(6021) <= a;
    layer3_outputs(6022) <= a and b;
    layer3_outputs(6023) <= a xor b;
    layer3_outputs(6024) <= not (a xor b);
    layer3_outputs(6025) <= a or b;
    layer3_outputs(6026) <= b and not a;
    layer3_outputs(6027) <= not a;
    layer3_outputs(6028) <= b;
    layer3_outputs(6029) <= a and b;
    layer3_outputs(6030) <= a;
    layer3_outputs(6031) <= b;
    layer3_outputs(6032) <= not b;
    layer3_outputs(6033) <= a xor b;
    layer3_outputs(6034) <= a xor b;
    layer3_outputs(6035) <= b;
    layer3_outputs(6036) <= not a;
    layer3_outputs(6037) <= a and b;
    layer3_outputs(6038) <= 1'b0;
    layer3_outputs(6039) <= a and not b;
    layer3_outputs(6040) <= a and not b;
    layer3_outputs(6041) <= not (a xor b);
    layer3_outputs(6042) <= not a;
    layer3_outputs(6043) <= not a;
    layer3_outputs(6044) <= 1'b0;
    layer3_outputs(6045) <= not a;
    layer3_outputs(6046) <= b;
    layer3_outputs(6047) <= not a;
    layer3_outputs(6048) <= a;
    layer3_outputs(6049) <= not (a xor b);
    layer3_outputs(6050) <= a xor b;
    layer3_outputs(6051) <= b;
    layer3_outputs(6052) <= not a;
    layer3_outputs(6053) <= not b;
    layer3_outputs(6054) <= not a;
    layer3_outputs(6055) <= a;
    layer3_outputs(6056) <= not a or b;
    layer3_outputs(6057) <= not (a or b);
    layer3_outputs(6058) <= a;
    layer3_outputs(6059) <= b;
    layer3_outputs(6060) <= a or b;
    layer3_outputs(6061) <= 1'b1;
    layer3_outputs(6062) <= not a;
    layer3_outputs(6063) <= a or b;
    layer3_outputs(6064) <= not (a or b);
    layer3_outputs(6065) <= a xor b;
    layer3_outputs(6066) <= a;
    layer3_outputs(6067) <= not b or a;
    layer3_outputs(6068) <= not (a or b);
    layer3_outputs(6069) <= not b or a;
    layer3_outputs(6070) <= not a;
    layer3_outputs(6071) <= a and not b;
    layer3_outputs(6072) <= a and not b;
    layer3_outputs(6073) <= b;
    layer3_outputs(6074) <= a and b;
    layer3_outputs(6075) <= not (a xor b);
    layer3_outputs(6076) <= b and not a;
    layer3_outputs(6077) <= b;
    layer3_outputs(6078) <= not a;
    layer3_outputs(6079) <= a xor b;
    layer3_outputs(6080) <= a xor b;
    layer3_outputs(6081) <= 1'b1;
    layer3_outputs(6082) <= not b;
    layer3_outputs(6083) <= a or b;
    layer3_outputs(6084) <= not a;
    layer3_outputs(6085) <= not (a and b);
    layer3_outputs(6086) <= not b;
    layer3_outputs(6087) <= not a;
    layer3_outputs(6088) <= not (a or b);
    layer3_outputs(6089) <= not a;
    layer3_outputs(6090) <= not a or b;
    layer3_outputs(6091) <= not (a xor b);
    layer3_outputs(6092) <= a or b;
    layer3_outputs(6093) <= a or b;
    layer3_outputs(6094) <= not b or a;
    layer3_outputs(6095) <= b;
    layer3_outputs(6096) <= not b or a;
    layer3_outputs(6097) <= not (a and b);
    layer3_outputs(6098) <= b and not a;
    layer3_outputs(6099) <= a;
    layer3_outputs(6100) <= b;
    layer3_outputs(6101) <= a;
    layer3_outputs(6102) <= b;
    layer3_outputs(6103) <= not a;
    layer3_outputs(6104) <= not b or a;
    layer3_outputs(6105) <= a;
    layer3_outputs(6106) <= a and b;
    layer3_outputs(6107) <= b and not a;
    layer3_outputs(6108) <= a or b;
    layer3_outputs(6109) <= not b;
    layer3_outputs(6110) <= a xor b;
    layer3_outputs(6111) <= a;
    layer3_outputs(6112) <= not a;
    layer3_outputs(6113) <= a and b;
    layer3_outputs(6114) <= a;
    layer3_outputs(6115) <= not a or b;
    layer3_outputs(6116) <= a or b;
    layer3_outputs(6117) <= a xor b;
    layer3_outputs(6118) <= not (a and b);
    layer3_outputs(6119) <= a and not b;
    layer3_outputs(6120) <= a and not b;
    layer3_outputs(6121) <= a xor b;
    layer3_outputs(6122) <= a;
    layer3_outputs(6123) <= b;
    layer3_outputs(6124) <= a;
    layer3_outputs(6125) <= not b;
    layer3_outputs(6126) <= not b or a;
    layer3_outputs(6127) <= not a;
    layer3_outputs(6128) <= not (a or b);
    layer3_outputs(6129) <= a or b;
    layer3_outputs(6130) <= not a;
    layer3_outputs(6131) <= not (a and b);
    layer3_outputs(6132) <= b;
    layer3_outputs(6133) <= a and b;
    layer3_outputs(6134) <= not a or b;
    layer3_outputs(6135) <= not (a or b);
    layer3_outputs(6136) <= a and not b;
    layer3_outputs(6137) <= a or b;
    layer3_outputs(6138) <= a;
    layer3_outputs(6139) <= a;
    layer3_outputs(6140) <= b;
    layer3_outputs(6141) <= not a or b;
    layer3_outputs(6142) <= not a or b;
    layer3_outputs(6143) <= a and not b;
    layer3_outputs(6144) <= a;
    layer3_outputs(6145) <= a xor b;
    layer3_outputs(6146) <= not a;
    layer3_outputs(6147) <= not b or a;
    layer3_outputs(6148) <= not b or a;
    layer3_outputs(6149) <= not (a or b);
    layer3_outputs(6150) <= not b;
    layer3_outputs(6151) <= not b or a;
    layer3_outputs(6152) <= not (a or b);
    layer3_outputs(6153) <= b;
    layer3_outputs(6154) <= not b or a;
    layer3_outputs(6155) <= a;
    layer3_outputs(6156) <= not b;
    layer3_outputs(6157) <= a or b;
    layer3_outputs(6158) <= not b or a;
    layer3_outputs(6159) <= 1'b0;
    layer3_outputs(6160) <= not (a or b);
    layer3_outputs(6161) <= b and not a;
    layer3_outputs(6162) <= not b;
    layer3_outputs(6163) <= not (a or b);
    layer3_outputs(6164) <= 1'b1;
    layer3_outputs(6165) <= b;
    layer3_outputs(6166) <= a xor b;
    layer3_outputs(6167) <= not b;
    layer3_outputs(6168) <= not b or a;
    layer3_outputs(6169) <= not b;
    layer3_outputs(6170) <= not a;
    layer3_outputs(6171) <= not (a and b);
    layer3_outputs(6172) <= not b;
    layer3_outputs(6173) <= a xor b;
    layer3_outputs(6174) <= 1'b0;
    layer3_outputs(6175) <= b;
    layer3_outputs(6176) <= not b or a;
    layer3_outputs(6177) <= b and not a;
    layer3_outputs(6178) <= not a or b;
    layer3_outputs(6179) <= a;
    layer3_outputs(6180) <= a and b;
    layer3_outputs(6181) <= b and not a;
    layer3_outputs(6182) <= not b;
    layer3_outputs(6183) <= a;
    layer3_outputs(6184) <= a;
    layer3_outputs(6185) <= b and not a;
    layer3_outputs(6186) <= not a;
    layer3_outputs(6187) <= b;
    layer3_outputs(6188) <= not (a or b);
    layer3_outputs(6189) <= a;
    layer3_outputs(6190) <= not a;
    layer3_outputs(6191) <= a xor b;
    layer3_outputs(6192) <= not (a xor b);
    layer3_outputs(6193) <= not (a xor b);
    layer3_outputs(6194) <= not (a or b);
    layer3_outputs(6195) <= b and not a;
    layer3_outputs(6196) <= not a;
    layer3_outputs(6197) <= b;
    layer3_outputs(6198) <= a;
    layer3_outputs(6199) <= a;
    layer3_outputs(6200) <= not a or b;
    layer3_outputs(6201) <= a xor b;
    layer3_outputs(6202) <= b and not a;
    layer3_outputs(6203) <= a;
    layer3_outputs(6204) <= b and not a;
    layer3_outputs(6205) <= not (a xor b);
    layer3_outputs(6206) <= a and not b;
    layer3_outputs(6207) <= b;
    layer3_outputs(6208) <= not b;
    layer3_outputs(6209) <= not a or b;
    layer3_outputs(6210) <= a and b;
    layer3_outputs(6211) <= not a;
    layer3_outputs(6212) <= not a;
    layer3_outputs(6213) <= not a;
    layer3_outputs(6214) <= not a;
    layer3_outputs(6215) <= a xor b;
    layer3_outputs(6216) <= a;
    layer3_outputs(6217) <= 1'b0;
    layer3_outputs(6218) <= not b or a;
    layer3_outputs(6219) <= b;
    layer3_outputs(6220) <= not a;
    layer3_outputs(6221) <= a and not b;
    layer3_outputs(6222) <= b;
    layer3_outputs(6223) <= not a or b;
    layer3_outputs(6224) <= not a or b;
    layer3_outputs(6225) <= a xor b;
    layer3_outputs(6226) <= b;
    layer3_outputs(6227) <= 1'b1;
    layer3_outputs(6228) <= b;
    layer3_outputs(6229) <= b and not a;
    layer3_outputs(6230) <= not a;
    layer3_outputs(6231) <= not b;
    layer3_outputs(6232) <= a and not b;
    layer3_outputs(6233) <= b;
    layer3_outputs(6234) <= a;
    layer3_outputs(6235) <= not b;
    layer3_outputs(6236) <= a xor b;
    layer3_outputs(6237) <= b and not a;
    layer3_outputs(6238) <= not a or b;
    layer3_outputs(6239) <= not (a xor b);
    layer3_outputs(6240) <= not a or b;
    layer3_outputs(6241) <= b;
    layer3_outputs(6242) <= not (a or b);
    layer3_outputs(6243) <= a and not b;
    layer3_outputs(6244) <= not a;
    layer3_outputs(6245) <= not b;
    layer3_outputs(6246) <= b;
    layer3_outputs(6247) <= not b;
    layer3_outputs(6248) <= not (a or b);
    layer3_outputs(6249) <= a;
    layer3_outputs(6250) <= b and not a;
    layer3_outputs(6251) <= not b;
    layer3_outputs(6252) <= 1'b1;
    layer3_outputs(6253) <= not (a xor b);
    layer3_outputs(6254) <= not a;
    layer3_outputs(6255) <= 1'b0;
    layer3_outputs(6256) <= not a;
    layer3_outputs(6257) <= not a;
    layer3_outputs(6258) <= a xor b;
    layer3_outputs(6259) <= not (a and b);
    layer3_outputs(6260) <= a;
    layer3_outputs(6261) <= not b or a;
    layer3_outputs(6262) <= b;
    layer3_outputs(6263) <= a;
    layer3_outputs(6264) <= not (a and b);
    layer3_outputs(6265) <= a;
    layer3_outputs(6266) <= a and b;
    layer3_outputs(6267) <= a or b;
    layer3_outputs(6268) <= not a;
    layer3_outputs(6269) <= b;
    layer3_outputs(6270) <= not b;
    layer3_outputs(6271) <= not b;
    layer3_outputs(6272) <= a;
    layer3_outputs(6273) <= not b;
    layer3_outputs(6274) <= a and not b;
    layer3_outputs(6275) <= not b;
    layer3_outputs(6276) <= not a;
    layer3_outputs(6277) <= a or b;
    layer3_outputs(6278) <= a;
    layer3_outputs(6279) <= b;
    layer3_outputs(6280) <= b and not a;
    layer3_outputs(6281) <= not a;
    layer3_outputs(6282) <= a and not b;
    layer3_outputs(6283) <= not b;
    layer3_outputs(6284) <= a xor b;
    layer3_outputs(6285) <= not a;
    layer3_outputs(6286) <= not b;
    layer3_outputs(6287) <= not a;
    layer3_outputs(6288) <= a;
    layer3_outputs(6289) <= a xor b;
    layer3_outputs(6290) <= b and not a;
    layer3_outputs(6291) <= a xor b;
    layer3_outputs(6292) <= a and b;
    layer3_outputs(6293) <= a or b;
    layer3_outputs(6294) <= a or b;
    layer3_outputs(6295) <= not a;
    layer3_outputs(6296) <= not b or a;
    layer3_outputs(6297) <= not (a xor b);
    layer3_outputs(6298) <= not b;
    layer3_outputs(6299) <= not (a xor b);
    layer3_outputs(6300) <= a;
    layer3_outputs(6301) <= a xor b;
    layer3_outputs(6302) <= a and not b;
    layer3_outputs(6303) <= b;
    layer3_outputs(6304) <= not a;
    layer3_outputs(6305) <= b;
    layer3_outputs(6306) <= b and not a;
    layer3_outputs(6307) <= a and b;
    layer3_outputs(6308) <= not (a or b);
    layer3_outputs(6309) <= not b or a;
    layer3_outputs(6310) <= a xor b;
    layer3_outputs(6311) <= 1'b0;
    layer3_outputs(6312) <= a;
    layer3_outputs(6313) <= not a;
    layer3_outputs(6314) <= a xor b;
    layer3_outputs(6315) <= a and not b;
    layer3_outputs(6316) <= b;
    layer3_outputs(6317) <= not b;
    layer3_outputs(6318) <= not a or b;
    layer3_outputs(6319) <= a;
    layer3_outputs(6320) <= a and b;
    layer3_outputs(6321) <= not b or a;
    layer3_outputs(6322) <= a and not b;
    layer3_outputs(6323) <= not (a and b);
    layer3_outputs(6324) <= not a;
    layer3_outputs(6325) <= a;
    layer3_outputs(6326) <= not a;
    layer3_outputs(6327) <= a;
    layer3_outputs(6328) <= a and not b;
    layer3_outputs(6329) <= not (a or b);
    layer3_outputs(6330) <= a or b;
    layer3_outputs(6331) <= a and not b;
    layer3_outputs(6332) <= 1'b0;
    layer3_outputs(6333) <= not a or b;
    layer3_outputs(6334) <= b and not a;
    layer3_outputs(6335) <= not (a xor b);
    layer3_outputs(6336) <= b and not a;
    layer3_outputs(6337) <= not b;
    layer3_outputs(6338) <= not a or b;
    layer3_outputs(6339) <= not a or b;
    layer3_outputs(6340) <= a;
    layer3_outputs(6341) <= not b;
    layer3_outputs(6342) <= not a or b;
    layer3_outputs(6343) <= not b or a;
    layer3_outputs(6344) <= b and not a;
    layer3_outputs(6345) <= a and not b;
    layer3_outputs(6346) <= a and b;
    layer3_outputs(6347) <= not b;
    layer3_outputs(6348) <= not (a and b);
    layer3_outputs(6349) <= not (a and b);
    layer3_outputs(6350) <= not a;
    layer3_outputs(6351) <= b;
    layer3_outputs(6352) <= a;
    layer3_outputs(6353) <= 1'b1;
    layer3_outputs(6354) <= not b;
    layer3_outputs(6355) <= not a or b;
    layer3_outputs(6356) <= not a;
    layer3_outputs(6357) <= a and b;
    layer3_outputs(6358) <= a;
    layer3_outputs(6359) <= b;
    layer3_outputs(6360) <= not (a and b);
    layer3_outputs(6361) <= not b;
    layer3_outputs(6362) <= a and b;
    layer3_outputs(6363) <= not (a and b);
    layer3_outputs(6364) <= not a or b;
    layer3_outputs(6365) <= b;
    layer3_outputs(6366) <= a;
    layer3_outputs(6367) <= b;
    layer3_outputs(6368) <= not a;
    layer3_outputs(6369) <= not (a or b);
    layer3_outputs(6370) <= a and b;
    layer3_outputs(6371) <= not a;
    layer3_outputs(6372) <= not a;
    layer3_outputs(6373) <= not a or b;
    layer3_outputs(6374) <= a;
    layer3_outputs(6375) <= a;
    layer3_outputs(6376) <= not (a xor b);
    layer3_outputs(6377) <= a;
    layer3_outputs(6378) <= b and not a;
    layer3_outputs(6379) <= not a;
    layer3_outputs(6380) <= not a;
    layer3_outputs(6381) <= a or b;
    layer3_outputs(6382) <= a and b;
    layer3_outputs(6383) <= a or b;
    layer3_outputs(6384) <= not b;
    layer3_outputs(6385) <= not (a or b);
    layer3_outputs(6386) <= not b or a;
    layer3_outputs(6387) <= a;
    layer3_outputs(6388) <= not (a xor b);
    layer3_outputs(6389) <= a and not b;
    layer3_outputs(6390) <= not (a xor b);
    layer3_outputs(6391) <= not b or a;
    layer3_outputs(6392) <= not (a or b);
    layer3_outputs(6393) <= a or b;
    layer3_outputs(6394) <= not b or a;
    layer3_outputs(6395) <= not a or b;
    layer3_outputs(6396) <= not (a or b);
    layer3_outputs(6397) <= b and not a;
    layer3_outputs(6398) <= not (a xor b);
    layer3_outputs(6399) <= a;
    layer3_outputs(6400) <= a and not b;
    layer3_outputs(6401) <= b;
    layer3_outputs(6402) <= not (a xor b);
    layer3_outputs(6403) <= not a;
    layer3_outputs(6404) <= a or b;
    layer3_outputs(6405) <= a;
    layer3_outputs(6406) <= b;
    layer3_outputs(6407) <= a or b;
    layer3_outputs(6408) <= 1'b0;
    layer3_outputs(6409) <= a;
    layer3_outputs(6410) <= not (a xor b);
    layer3_outputs(6411) <= not (a xor b);
    layer3_outputs(6412) <= not b;
    layer3_outputs(6413) <= b;
    layer3_outputs(6414) <= a;
    layer3_outputs(6415) <= not b;
    layer3_outputs(6416) <= not a;
    layer3_outputs(6417) <= a or b;
    layer3_outputs(6418) <= 1'b1;
    layer3_outputs(6419) <= a and b;
    layer3_outputs(6420) <= b;
    layer3_outputs(6421) <= not (a and b);
    layer3_outputs(6422) <= not b or a;
    layer3_outputs(6423) <= not b or a;
    layer3_outputs(6424) <= a and b;
    layer3_outputs(6425) <= a or b;
    layer3_outputs(6426) <= not a or b;
    layer3_outputs(6427) <= a xor b;
    layer3_outputs(6428) <= not b or a;
    layer3_outputs(6429) <= not a or b;
    layer3_outputs(6430) <= not a;
    layer3_outputs(6431) <= a;
    layer3_outputs(6432) <= a xor b;
    layer3_outputs(6433) <= not b;
    layer3_outputs(6434) <= a and b;
    layer3_outputs(6435) <= b;
    layer3_outputs(6436) <= a and b;
    layer3_outputs(6437) <= not b;
    layer3_outputs(6438) <= a;
    layer3_outputs(6439) <= not a;
    layer3_outputs(6440) <= a and b;
    layer3_outputs(6441) <= not a;
    layer3_outputs(6442) <= not (a or b);
    layer3_outputs(6443) <= not a or b;
    layer3_outputs(6444) <= not b or a;
    layer3_outputs(6445) <= b;
    layer3_outputs(6446) <= not (a xor b);
    layer3_outputs(6447) <= a;
    layer3_outputs(6448) <= b;
    layer3_outputs(6449) <= not b;
    layer3_outputs(6450) <= a or b;
    layer3_outputs(6451) <= not (a and b);
    layer3_outputs(6452) <= a;
    layer3_outputs(6453) <= a or b;
    layer3_outputs(6454) <= a and not b;
    layer3_outputs(6455) <= a;
    layer3_outputs(6456) <= not a;
    layer3_outputs(6457) <= not a or b;
    layer3_outputs(6458) <= a and not b;
    layer3_outputs(6459) <= not a;
    layer3_outputs(6460) <= not b;
    layer3_outputs(6461) <= a and b;
    layer3_outputs(6462) <= not b;
    layer3_outputs(6463) <= a and b;
    layer3_outputs(6464) <= a;
    layer3_outputs(6465) <= not a or b;
    layer3_outputs(6466) <= a xor b;
    layer3_outputs(6467) <= a xor b;
    layer3_outputs(6468) <= a xor b;
    layer3_outputs(6469) <= a xor b;
    layer3_outputs(6470) <= a or b;
    layer3_outputs(6471) <= b;
    layer3_outputs(6472) <= a;
    layer3_outputs(6473) <= a;
    layer3_outputs(6474) <= not (a xor b);
    layer3_outputs(6475) <= a or b;
    layer3_outputs(6476) <= b;
    layer3_outputs(6477) <= a and not b;
    layer3_outputs(6478) <= a or b;
    layer3_outputs(6479) <= not (a or b);
    layer3_outputs(6480) <= not b;
    layer3_outputs(6481) <= a and not b;
    layer3_outputs(6482) <= not (a xor b);
    layer3_outputs(6483) <= not a;
    layer3_outputs(6484) <= 1'b0;
    layer3_outputs(6485) <= a and b;
    layer3_outputs(6486) <= a or b;
    layer3_outputs(6487) <= not (a and b);
    layer3_outputs(6488) <= not b;
    layer3_outputs(6489) <= b;
    layer3_outputs(6490) <= a;
    layer3_outputs(6491) <= b and not a;
    layer3_outputs(6492) <= a xor b;
    layer3_outputs(6493) <= not b or a;
    layer3_outputs(6494) <= not (a and b);
    layer3_outputs(6495) <= not a;
    layer3_outputs(6496) <= not a;
    layer3_outputs(6497) <= a and b;
    layer3_outputs(6498) <= not b;
    layer3_outputs(6499) <= not (a or b);
    layer3_outputs(6500) <= b;
    layer3_outputs(6501) <= b and not a;
    layer3_outputs(6502) <= a and b;
    layer3_outputs(6503) <= not b;
    layer3_outputs(6504) <= not (a or b);
    layer3_outputs(6505) <= not (a and b);
    layer3_outputs(6506) <= not (a and b);
    layer3_outputs(6507) <= a and b;
    layer3_outputs(6508) <= not (a xor b);
    layer3_outputs(6509) <= a or b;
    layer3_outputs(6510) <= a;
    layer3_outputs(6511) <= not b or a;
    layer3_outputs(6512) <= not b or a;
    layer3_outputs(6513) <= a or b;
    layer3_outputs(6514) <= b;
    layer3_outputs(6515) <= a xor b;
    layer3_outputs(6516) <= not a;
    layer3_outputs(6517) <= not b;
    layer3_outputs(6518) <= b;
    layer3_outputs(6519) <= a and b;
    layer3_outputs(6520) <= not a;
    layer3_outputs(6521) <= b and not a;
    layer3_outputs(6522) <= a and b;
    layer3_outputs(6523) <= not b or a;
    layer3_outputs(6524) <= not a;
    layer3_outputs(6525) <= not (a xor b);
    layer3_outputs(6526) <= not (a and b);
    layer3_outputs(6527) <= a or b;
    layer3_outputs(6528) <= not (a and b);
    layer3_outputs(6529) <= a;
    layer3_outputs(6530) <= b;
    layer3_outputs(6531) <= not a;
    layer3_outputs(6532) <= 1'b1;
    layer3_outputs(6533) <= not a;
    layer3_outputs(6534) <= a xor b;
    layer3_outputs(6535) <= not a;
    layer3_outputs(6536) <= a xor b;
    layer3_outputs(6537) <= not b;
    layer3_outputs(6538) <= a;
    layer3_outputs(6539) <= not b;
    layer3_outputs(6540) <= a xor b;
    layer3_outputs(6541) <= a;
    layer3_outputs(6542) <= not a;
    layer3_outputs(6543) <= b;
    layer3_outputs(6544) <= a and b;
    layer3_outputs(6545) <= 1'b0;
    layer3_outputs(6546) <= not a;
    layer3_outputs(6547) <= a and not b;
    layer3_outputs(6548) <= b;
    layer3_outputs(6549) <= a or b;
    layer3_outputs(6550) <= a;
    layer3_outputs(6551) <= a;
    layer3_outputs(6552) <= not a;
    layer3_outputs(6553) <= a and not b;
    layer3_outputs(6554) <= b;
    layer3_outputs(6555) <= a and b;
    layer3_outputs(6556) <= not a;
    layer3_outputs(6557) <= a and not b;
    layer3_outputs(6558) <= a or b;
    layer3_outputs(6559) <= not (a and b);
    layer3_outputs(6560) <= a and not b;
    layer3_outputs(6561) <= not a;
    layer3_outputs(6562) <= a;
    layer3_outputs(6563) <= not a;
    layer3_outputs(6564) <= b and not a;
    layer3_outputs(6565) <= b;
    layer3_outputs(6566) <= b;
    layer3_outputs(6567) <= not a;
    layer3_outputs(6568) <= a and b;
    layer3_outputs(6569) <= not a;
    layer3_outputs(6570) <= not b;
    layer3_outputs(6571) <= not b;
    layer3_outputs(6572) <= a and not b;
    layer3_outputs(6573) <= not (a or b);
    layer3_outputs(6574) <= a and b;
    layer3_outputs(6575) <= not (a xor b);
    layer3_outputs(6576) <= a;
    layer3_outputs(6577) <= not b or a;
    layer3_outputs(6578) <= not b;
    layer3_outputs(6579) <= b;
    layer3_outputs(6580) <= a or b;
    layer3_outputs(6581) <= not a;
    layer3_outputs(6582) <= a;
    layer3_outputs(6583) <= a and not b;
    layer3_outputs(6584) <= not a;
    layer3_outputs(6585) <= not b or a;
    layer3_outputs(6586) <= not (a or b);
    layer3_outputs(6587) <= not (a or b);
    layer3_outputs(6588) <= a;
    layer3_outputs(6589) <= b;
    layer3_outputs(6590) <= a xor b;
    layer3_outputs(6591) <= b and not a;
    layer3_outputs(6592) <= not a;
    layer3_outputs(6593) <= not (a and b);
    layer3_outputs(6594) <= not a;
    layer3_outputs(6595) <= b and not a;
    layer3_outputs(6596) <= not (a xor b);
    layer3_outputs(6597) <= b;
    layer3_outputs(6598) <= b;
    layer3_outputs(6599) <= b;
    layer3_outputs(6600) <= b;
    layer3_outputs(6601) <= not a or b;
    layer3_outputs(6602) <= not b;
    layer3_outputs(6603) <= not (a and b);
    layer3_outputs(6604) <= a;
    layer3_outputs(6605) <= b and not a;
    layer3_outputs(6606) <= not b or a;
    layer3_outputs(6607) <= not a or b;
    layer3_outputs(6608) <= not b;
    layer3_outputs(6609) <= 1'b1;
    layer3_outputs(6610) <= not b;
    layer3_outputs(6611) <= not a;
    layer3_outputs(6612) <= b;
    layer3_outputs(6613) <= not (a and b);
    layer3_outputs(6614) <= not a;
    layer3_outputs(6615) <= not b;
    layer3_outputs(6616) <= b;
    layer3_outputs(6617) <= not a or b;
    layer3_outputs(6618) <= not b;
    layer3_outputs(6619) <= a;
    layer3_outputs(6620) <= a and b;
    layer3_outputs(6621) <= a;
    layer3_outputs(6622) <= a and b;
    layer3_outputs(6623) <= not (a or b);
    layer3_outputs(6624) <= not (a xor b);
    layer3_outputs(6625) <= not a;
    layer3_outputs(6626) <= b;
    layer3_outputs(6627) <= a;
    layer3_outputs(6628) <= not a;
    layer3_outputs(6629) <= not (a xor b);
    layer3_outputs(6630) <= a;
    layer3_outputs(6631) <= a;
    layer3_outputs(6632) <= not (a and b);
    layer3_outputs(6633) <= a;
    layer3_outputs(6634) <= a and not b;
    layer3_outputs(6635) <= a;
    layer3_outputs(6636) <= a or b;
    layer3_outputs(6637) <= not a;
    layer3_outputs(6638) <= b;
    layer3_outputs(6639) <= a xor b;
    layer3_outputs(6640) <= not (a xor b);
    layer3_outputs(6641) <= a;
    layer3_outputs(6642) <= a;
    layer3_outputs(6643) <= a xor b;
    layer3_outputs(6644) <= b and not a;
    layer3_outputs(6645) <= not b;
    layer3_outputs(6646) <= not (a or b);
    layer3_outputs(6647) <= a xor b;
    layer3_outputs(6648) <= a;
    layer3_outputs(6649) <= not a;
    layer3_outputs(6650) <= not b;
    layer3_outputs(6651) <= not (a xor b);
    layer3_outputs(6652) <= not (a xor b);
    layer3_outputs(6653) <= not a or b;
    layer3_outputs(6654) <= a or b;
    layer3_outputs(6655) <= not (a xor b);
    layer3_outputs(6656) <= a and b;
    layer3_outputs(6657) <= not (a xor b);
    layer3_outputs(6658) <= not b;
    layer3_outputs(6659) <= not (a or b);
    layer3_outputs(6660) <= b;
    layer3_outputs(6661) <= not a;
    layer3_outputs(6662) <= not a or b;
    layer3_outputs(6663) <= not a;
    layer3_outputs(6664) <= not a;
    layer3_outputs(6665) <= a;
    layer3_outputs(6666) <= not b;
    layer3_outputs(6667) <= not (a or b);
    layer3_outputs(6668) <= not b;
    layer3_outputs(6669) <= not a or b;
    layer3_outputs(6670) <= not a;
    layer3_outputs(6671) <= 1'b1;
    layer3_outputs(6672) <= a and b;
    layer3_outputs(6673) <= a and b;
    layer3_outputs(6674) <= a or b;
    layer3_outputs(6675) <= b and not a;
    layer3_outputs(6676) <= b;
    layer3_outputs(6677) <= a;
    layer3_outputs(6678) <= not (a or b);
    layer3_outputs(6679) <= not b or a;
    layer3_outputs(6680) <= not a;
    layer3_outputs(6681) <= not (a and b);
    layer3_outputs(6682) <= b and not a;
    layer3_outputs(6683) <= a and b;
    layer3_outputs(6684) <= not (a xor b);
    layer3_outputs(6685) <= not b or a;
    layer3_outputs(6686) <= a and b;
    layer3_outputs(6687) <= not (a xor b);
    layer3_outputs(6688) <= a or b;
    layer3_outputs(6689) <= a xor b;
    layer3_outputs(6690) <= not (a or b);
    layer3_outputs(6691) <= not a;
    layer3_outputs(6692) <= not b;
    layer3_outputs(6693) <= not (a xor b);
    layer3_outputs(6694) <= not a;
    layer3_outputs(6695) <= b;
    layer3_outputs(6696) <= not b or a;
    layer3_outputs(6697) <= not a;
    layer3_outputs(6698) <= a;
    layer3_outputs(6699) <= not (a xor b);
    layer3_outputs(6700) <= not (a xor b);
    layer3_outputs(6701) <= b;
    layer3_outputs(6702) <= not b or a;
    layer3_outputs(6703) <= 1'b0;
    layer3_outputs(6704) <= not (a xor b);
    layer3_outputs(6705) <= not b;
    layer3_outputs(6706) <= a or b;
    layer3_outputs(6707) <= b and not a;
    layer3_outputs(6708) <= not a;
    layer3_outputs(6709) <= not b;
    layer3_outputs(6710) <= b and not a;
    layer3_outputs(6711) <= not (a or b);
    layer3_outputs(6712) <= a and b;
    layer3_outputs(6713) <= not (a xor b);
    layer3_outputs(6714) <= b;
    layer3_outputs(6715) <= a or b;
    layer3_outputs(6716) <= a and not b;
    layer3_outputs(6717) <= not a;
    layer3_outputs(6718) <= a xor b;
    layer3_outputs(6719) <= a and b;
    layer3_outputs(6720) <= not a;
    layer3_outputs(6721) <= a or b;
    layer3_outputs(6722) <= b;
    layer3_outputs(6723) <= not b or a;
    layer3_outputs(6724) <= a or b;
    layer3_outputs(6725) <= not (a or b);
    layer3_outputs(6726) <= b and not a;
    layer3_outputs(6727) <= b;
    layer3_outputs(6728) <= a;
    layer3_outputs(6729) <= a and b;
    layer3_outputs(6730) <= not b;
    layer3_outputs(6731) <= a and b;
    layer3_outputs(6732) <= a or b;
    layer3_outputs(6733) <= a xor b;
    layer3_outputs(6734) <= a;
    layer3_outputs(6735) <= b;
    layer3_outputs(6736) <= not b;
    layer3_outputs(6737) <= not a or b;
    layer3_outputs(6738) <= a and b;
    layer3_outputs(6739) <= b;
    layer3_outputs(6740) <= not a or b;
    layer3_outputs(6741) <= b and not a;
    layer3_outputs(6742) <= not (a xor b);
    layer3_outputs(6743) <= not b;
    layer3_outputs(6744) <= a xor b;
    layer3_outputs(6745) <= a xor b;
    layer3_outputs(6746) <= not a;
    layer3_outputs(6747) <= a and b;
    layer3_outputs(6748) <= a and b;
    layer3_outputs(6749) <= not b;
    layer3_outputs(6750) <= not (a xor b);
    layer3_outputs(6751) <= b and not a;
    layer3_outputs(6752) <= not b;
    layer3_outputs(6753) <= b and not a;
    layer3_outputs(6754) <= not b;
    layer3_outputs(6755) <= a xor b;
    layer3_outputs(6756) <= not (a and b);
    layer3_outputs(6757) <= not (a xor b);
    layer3_outputs(6758) <= a xor b;
    layer3_outputs(6759) <= not b or a;
    layer3_outputs(6760) <= b;
    layer3_outputs(6761) <= a;
    layer3_outputs(6762) <= a xor b;
    layer3_outputs(6763) <= a and not b;
    layer3_outputs(6764) <= not a;
    layer3_outputs(6765) <= not (a and b);
    layer3_outputs(6766) <= not b or a;
    layer3_outputs(6767) <= a or b;
    layer3_outputs(6768) <= b and not a;
    layer3_outputs(6769) <= a and b;
    layer3_outputs(6770) <= b;
    layer3_outputs(6771) <= not (a and b);
    layer3_outputs(6772) <= not (a or b);
    layer3_outputs(6773) <= a or b;
    layer3_outputs(6774) <= b;
    layer3_outputs(6775) <= b;
    layer3_outputs(6776) <= not (a or b);
    layer3_outputs(6777) <= not (a or b);
    layer3_outputs(6778) <= b and not a;
    layer3_outputs(6779) <= b;
    layer3_outputs(6780) <= not a;
    layer3_outputs(6781) <= not a or b;
    layer3_outputs(6782) <= a and not b;
    layer3_outputs(6783) <= a xor b;
    layer3_outputs(6784) <= not a;
    layer3_outputs(6785) <= not (a or b);
    layer3_outputs(6786) <= not b;
    layer3_outputs(6787) <= a or b;
    layer3_outputs(6788) <= a;
    layer3_outputs(6789) <= not a or b;
    layer3_outputs(6790) <= b and not a;
    layer3_outputs(6791) <= b;
    layer3_outputs(6792) <= a and not b;
    layer3_outputs(6793) <= not b;
    layer3_outputs(6794) <= not b or a;
    layer3_outputs(6795) <= a;
    layer3_outputs(6796) <= not (a or b);
    layer3_outputs(6797) <= a or b;
    layer3_outputs(6798) <= a;
    layer3_outputs(6799) <= a;
    layer3_outputs(6800) <= not b or a;
    layer3_outputs(6801) <= 1'b0;
    layer3_outputs(6802) <= a;
    layer3_outputs(6803) <= a;
    layer3_outputs(6804) <= b and not a;
    layer3_outputs(6805) <= a and not b;
    layer3_outputs(6806) <= not (a and b);
    layer3_outputs(6807) <= not b;
    layer3_outputs(6808) <= a xor b;
    layer3_outputs(6809) <= a;
    layer3_outputs(6810) <= b;
    layer3_outputs(6811) <= a xor b;
    layer3_outputs(6812) <= not (a xor b);
    layer3_outputs(6813) <= not (a xor b);
    layer3_outputs(6814) <= not b or a;
    layer3_outputs(6815) <= not b or a;
    layer3_outputs(6816) <= a and not b;
    layer3_outputs(6817) <= 1'b0;
    layer3_outputs(6818) <= a or b;
    layer3_outputs(6819) <= not b;
    layer3_outputs(6820) <= a and b;
    layer3_outputs(6821) <= b;
    layer3_outputs(6822) <= not a or b;
    layer3_outputs(6823) <= b;
    layer3_outputs(6824) <= b and not a;
    layer3_outputs(6825) <= not a;
    layer3_outputs(6826) <= a and b;
    layer3_outputs(6827) <= not (a or b);
    layer3_outputs(6828) <= a and b;
    layer3_outputs(6829) <= not a;
    layer3_outputs(6830) <= not b;
    layer3_outputs(6831) <= not a or b;
    layer3_outputs(6832) <= not b or a;
    layer3_outputs(6833) <= not a;
    layer3_outputs(6834) <= a;
    layer3_outputs(6835) <= a xor b;
    layer3_outputs(6836) <= b and not a;
    layer3_outputs(6837) <= a;
    layer3_outputs(6838) <= not (a and b);
    layer3_outputs(6839) <= a and b;
    layer3_outputs(6840) <= not a;
    layer3_outputs(6841) <= not (a xor b);
    layer3_outputs(6842) <= not (a and b);
    layer3_outputs(6843) <= not a or b;
    layer3_outputs(6844) <= not a or b;
    layer3_outputs(6845) <= not b;
    layer3_outputs(6846) <= a and not b;
    layer3_outputs(6847) <= not (a xor b);
    layer3_outputs(6848) <= not a or b;
    layer3_outputs(6849) <= a xor b;
    layer3_outputs(6850) <= a and b;
    layer3_outputs(6851) <= not a;
    layer3_outputs(6852) <= a and not b;
    layer3_outputs(6853) <= not a or b;
    layer3_outputs(6854) <= b;
    layer3_outputs(6855) <= not b;
    layer3_outputs(6856) <= not (a xor b);
    layer3_outputs(6857) <= not b;
    layer3_outputs(6858) <= not b;
    layer3_outputs(6859) <= a and b;
    layer3_outputs(6860) <= not b;
    layer3_outputs(6861) <= not b;
    layer3_outputs(6862) <= a and not b;
    layer3_outputs(6863) <= a;
    layer3_outputs(6864) <= b and not a;
    layer3_outputs(6865) <= not b;
    layer3_outputs(6866) <= a and not b;
    layer3_outputs(6867) <= not (a or b);
    layer3_outputs(6868) <= not a;
    layer3_outputs(6869) <= not b;
    layer3_outputs(6870) <= not a or b;
    layer3_outputs(6871) <= not b;
    layer3_outputs(6872) <= a and b;
    layer3_outputs(6873) <= b;
    layer3_outputs(6874) <= not a;
    layer3_outputs(6875) <= not (a and b);
    layer3_outputs(6876) <= not a;
    layer3_outputs(6877) <= not b or a;
    layer3_outputs(6878) <= not a or b;
    layer3_outputs(6879) <= not (a or b);
    layer3_outputs(6880) <= not b;
    layer3_outputs(6881) <= not (a xor b);
    layer3_outputs(6882) <= a and not b;
    layer3_outputs(6883) <= 1'b0;
    layer3_outputs(6884) <= not b;
    layer3_outputs(6885) <= not b;
    layer3_outputs(6886) <= not (a and b);
    layer3_outputs(6887) <= not a;
    layer3_outputs(6888) <= a;
    layer3_outputs(6889) <= a xor b;
    layer3_outputs(6890) <= not (a xor b);
    layer3_outputs(6891) <= not (a or b);
    layer3_outputs(6892) <= not b or a;
    layer3_outputs(6893) <= a;
    layer3_outputs(6894) <= a and b;
    layer3_outputs(6895) <= not a;
    layer3_outputs(6896) <= a;
    layer3_outputs(6897) <= b;
    layer3_outputs(6898) <= not b;
    layer3_outputs(6899) <= not a;
    layer3_outputs(6900) <= a;
    layer3_outputs(6901) <= a or b;
    layer3_outputs(6902) <= a and b;
    layer3_outputs(6903) <= not (a xor b);
    layer3_outputs(6904) <= a;
    layer3_outputs(6905) <= b;
    layer3_outputs(6906) <= a xor b;
    layer3_outputs(6907) <= not b;
    layer3_outputs(6908) <= not b or a;
    layer3_outputs(6909) <= b;
    layer3_outputs(6910) <= 1'b0;
    layer3_outputs(6911) <= a;
    layer3_outputs(6912) <= b;
    layer3_outputs(6913) <= b;
    layer3_outputs(6914) <= a xor b;
    layer3_outputs(6915) <= a xor b;
    layer3_outputs(6916) <= a or b;
    layer3_outputs(6917) <= not a or b;
    layer3_outputs(6918) <= not a;
    layer3_outputs(6919) <= b;
    layer3_outputs(6920) <= 1'b0;
    layer3_outputs(6921) <= not a;
    layer3_outputs(6922) <= b and not a;
    layer3_outputs(6923) <= not b or a;
    layer3_outputs(6924) <= not b;
    layer3_outputs(6925) <= a;
    layer3_outputs(6926) <= a xor b;
    layer3_outputs(6927) <= b and not a;
    layer3_outputs(6928) <= not b or a;
    layer3_outputs(6929) <= b and not a;
    layer3_outputs(6930) <= a or b;
    layer3_outputs(6931) <= not (a or b);
    layer3_outputs(6932) <= not a;
    layer3_outputs(6933) <= not a;
    layer3_outputs(6934) <= b;
    layer3_outputs(6935) <= not (a and b);
    layer3_outputs(6936) <= a or b;
    layer3_outputs(6937) <= not b or a;
    layer3_outputs(6938) <= 1'b1;
    layer3_outputs(6939) <= not a or b;
    layer3_outputs(6940) <= not (a or b);
    layer3_outputs(6941) <= not a or b;
    layer3_outputs(6942) <= a;
    layer3_outputs(6943) <= b;
    layer3_outputs(6944) <= b;
    layer3_outputs(6945) <= a and b;
    layer3_outputs(6946) <= not (a and b);
    layer3_outputs(6947) <= not a;
    layer3_outputs(6948) <= b and not a;
    layer3_outputs(6949) <= b;
    layer3_outputs(6950) <= not b;
    layer3_outputs(6951) <= not (a xor b);
    layer3_outputs(6952) <= a and b;
    layer3_outputs(6953) <= not b;
    layer3_outputs(6954) <= not (a and b);
    layer3_outputs(6955) <= a and not b;
    layer3_outputs(6956) <= a;
    layer3_outputs(6957) <= not (a and b);
    layer3_outputs(6958) <= not (a xor b);
    layer3_outputs(6959) <= a xor b;
    layer3_outputs(6960) <= b;
    layer3_outputs(6961) <= a xor b;
    layer3_outputs(6962) <= a;
    layer3_outputs(6963) <= not b;
    layer3_outputs(6964) <= a and b;
    layer3_outputs(6965) <= a;
    layer3_outputs(6966) <= a;
    layer3_outputs(6967) <= a or b;
    layer3_outputs(6968) <= b;
    layer3_outputs(6969) <= not (a and b);
    layer3_outputs(6970) <= 1'b0;
    layer3_outputs(6971) <= a and not b;
    layer3_outputs(6972) <= b and not a;
    layer3_outputs(6973) <= a xor b;
    layer3_outputs(6974) <= not (a and b);
    layer3_outputs(6975) <= a and not b;
    layer3_outputs(6976) <= b;
    layer3_outputs(6977) <= a and not b;
    layer3_outputs(6978) <= not b;
    layer3_outputs(6979) <= not (a and b);
    layer3_outputs(6980) <= not b;
    layer3_outputs(6981) <= a and not b;
    layer3_outputs(6982) <= a xor b;
    layer3_outputs(6983) <= 1'b1;
    layer3_outputs(6984) <= a xor b;
    layer3_outputs(6985) <= b;
    layer3_outputs(6986) <= a;
    layer3_outputs(6987) <= b;
    layer3_outputs(6988) <= not b;
    layer3_outputs(6989) <= not a or b;
    layer3_outputs(6990) <= a;
    layer3_outputs(6991) <= not b;
    layer3_outputs(6992) <= a or b;
    layer3_outputs(6993) <= not b;
    layer3_outputs(6994) <= a xor b;
    layer3_outputs(6995) <= a and b;
    layer3_outputs(6996) <= not b;
    layer3_outputs(6997) <= not b or a;
    layer3_outputs(6998) <= a and b;
    layer3_outputs(6999) <= b;
    layer3_outputs(7000) <= a;
    layer3_outputs(7001) <= b and not a;
    layer3_outputs(7002) <= a or b;
    layer3_outputs(7003) <= b;
    layer3_outputs(7004) <= not a;
    layer3_outputs(7005) <= not b;
    layer3_outputs(7006) <= not (a and b);
    layer3_outputs(7007) <= not (a or b);
    layer3_outputs(7008) <= a;
    layer3_outputs(7009) <= not b;
    layer3_outputs(7010) <= not (a and b);
    layer3_outputs(7011) <= not (a xor b);
    layer3_outputs(7012) <= not b;
    layer3_outputs(7013) <= a;
    layer3_outputs(7014) <= not b;
    layer3_outputs(7015) <= not a;
    layer3_outputs(7016) <= b;
    layer3_outputs(7017) <= a or b;
    layer3_outputs(7018) <= a xor b;
    layer3_outputs(7019) <= not (a xor b);
    layer3_outputs(7020) <= not (a or b);
    layer3_outputs(7021) <= a and b;
    layer3_outputs(7022) <= not (a xor b);
    layer3_outputs(7023) <= not (a xor b);
    layer3_outputs(7024) <= a xor b;
    layer3_outputs(7025) <= 1'b1;
    layer3_outputs(7026) <= not b;
    layer3_outputs(7027) <= not (a or b);
    layer3_outputs(7028) <= not b;
    layer3_outputs(7029) <= a;
    layer3_outputs(7030) <= not a or b;
    layer3_outputs(7031) <= not a or b;
    layer3_outputs(7032) <= a;
    layer3_outputs(7033) <= b;
    layer3_outputs(7034) <= a;
    layer3_outputs(7035) <= a;
    layer3_outputs(7036) <= not a;
    layer3_outputs(7037) <= not (a or b);
    layer3_outputs(7038) <= not a or b;
    layer3_outputs(7039) <= not (a xor b);
    layer3_outputs(7040) <= not b or a;
    layer3_outputs(7041) <= 1'b1;
    layer3_outputs(7042) <= a xor b;
    layer3_outputs(7043) <= not a;
    layer3_outputs(7044) <= a and not b;
    layer3_outputs(7045) <= not a or b;
    layer3_outputs(7046) <= not a or b;
    layer3_outputs(7047) <= not (a or b);
    layer3_outputs(7048) <= a;
    layer3_outputs(7049) <= a and b;
    layer3_outputs(7050) <= not (a and b);
    layer3_outputs(7051) <= b;
    layer3_outputs(7052) <= a and b;
    layer3_outputs(7053) <= b;
    layer3_outputs(7054) <= not (a xor b);
    layer3_outputs(7055) <= not a or b;
    layer3_outputs(7056) <= b and not a;
    layer3_outputs(7057) <= a and b;
    layer3_outputs(7058) <= b and not a;
    layer3_outputs(7059) <= not (a or b);
    layer3_outputs(7060) <= b and not a;
    layer3_outputs(7061) <= a;
    layer3_outputs(7062) <= not b;
    layer3_outputs(7063) <= not b or a;
    layer3_outputs(7064) <= not a;
    layer3_outputs(7065) <= not b;
    layer3_outputs(7066) <= a xor b;
    layer3_outputs(7067) <= b;
    layer3_outputs(7068) <= a;
    layer3_outputs(7069) <= not a or b;
    layer3_outputs(7070) <= not a or b;
    layer3_outputs(7071) <= not b;
    layer3_outputs(7072) <= b and not a;
    layer3_outputs(7073) <= a xor b;
    layer3_outputs(7074) <= a and b;
    layer3_outputs(7075) <= not (a or b);
    layer3_outputs(7076) <= b;
    layer3_outputs(7077) <= not (a xor b);
    layer3_outputs(7078) <= not b;
    layer3_outputs(7079) <= b and not a;
    layer3_outputs(7080) <= b;
    layer3_outputs(7081) <= 1'b1;
    layer3_outputs(7082) <= not (a and b);
    layer3_outputs(7083) <= a and not b;
    layer3_outputs(7084) <= not b or a;
    layer3_outputs(7085) <= a or b;
    layer3_outputs(7086) <= b;
    layer3_outputs(7087) <= not (a and b);
    layer3_outputs(7088) <= not a;
    layer3_outputs(7089) <= a xor b;
    layer3_outputs(7090) <= b;
    layer3_outputs(7091) <= a and not b;
    layer3_outputs(7092) <= not (a and b);
    layer3_outputs(7093) <= a;
    layer3_outputs(7094) <= not (a or b);
    layer3_outputs(7095) <= not a;
    layer3_outputs(7096) <= not (a xor b);
    layer3_outputs(7097) <= a or b;
    layer3_outputs(7098) <= b and not a;
    layer3_outputs(7099) <= not b;
    layer3_outputs(7100) <= not (a and b);
    layer3_outputs(7101) <= b;
    layer3_outputs(7102) <= b;
    layer3_outputs(7103) <= a and b;
    layer3_outputs(7104) <= not b;
    layer3_outputs(7105) <= not a;
    layer3_outputs(7106) <= b;
    layer3_outputs(7107) <= not a;
    layer3_outputs(7108) <= a and b;
    layer3_outputs(7109) <= b;
    layer3_outputs(7110) <= not b;
    layer3_outputs(7111) <= a and not b;
    layer3_outputs(7112) <= not a;
    layer3_outputs(7113) <= not a;
    layer3_outputs(7114) <= 1'b1;
    layer3_outputs(7115) <= not (a or b);
    layer3_outputs(7116) <= a or b;
    layer3_outputs(7117) <= a;
    layer3_outputs(7118) <= not (a xor b);
    layer3_outputs(7119) <= a or b;
    layer3_outputs(7120) <= a and b;
    layer3_outputs(7121) <= a and not b;
    layer3_outputs(7122) <= a or b;
    layer3_outputs(7123) <= not a;
    layer3_outputs(7124) <= not b;
    layer3_outputs(7125) <= not (a xor b);
    layer3_outputs(7126) <= 1'b0;
    layer3_outputs(7127) <= not b;
    layer3_outputs(7128) <= a xor b;
    layer3_outputs(7129) <= not (a xor b);
    layer3_outputs(7130) <= not b;
    layer3_outputs(7131) <= b;
    layer3_outputs(7132) <= a xor b;
    layer3_outputs(7133) <= a;
    layer3_outputs(7134) <= a and not b;
    layer3_outputs(7135) <= b;
    layer3_outputs(7136) <= b;
    layer3_outputs(7137) <= a and not b;
    layer3_outputs(7138) <= 1'b1;
    layer3_outputs(7139) <= not a;
    layer3_outputs(7140) <= not (a or b);
    layer3_outputs(7141) <= not (a and b);
    layer3_outputs(7142) <= not a;
    layer3_outputs(7143) <= b;
    layer3_outputs(7144) <= a xor b;
    layer3_outputs(7145) <= b;
    layer3_outputs(7146) <= a and not b;
    layer3_outputs(7147) <= not (a xor b);
    layer3_outputs(7148) <= a;
    layer3_outputs(7149) <= not a;
    layer3_outputs(7150) <= b;
    layer3_outputs(7151) <= a and b;
    layer3_outputs(7152) <= not a or b;
    layer3_outputs(7153) <= a and b;
    layer3_outputs(7154) <= not (a xor b);
    layer3_outputs(7155) <= a xor b;
    layer3_outputs(7156) <= a;
    layer3_outputs(7157) <= not (a xor b);
    layer3_outputs(7158) <= not (a and b);
    layer3_outputs(7159) <= b and not a;
    layer3_outputs(7160) <= a and b;
    layer3_outputs(7161) <= not (a xor b);
    layer3_outputs(7162) <= not (a xor b);
    layer3_outputs(7163) <= b;
    layer3_outputs(7164) <= b;
    layer3_outputs(7165) <= b;
    layer3_outputs(7166) <= not a;
    layer3_outputs(7167) <= not b;
    layer3_outputs(7168) <= not (a and b);
    layer3_outputs(7169) <= a or b;
    layer3_outputs(7170) <= a;
    layer3_outputs(7171) <= b;
    layer3_outputs(7172) <= b;
    layer3_outputs(7173) <= a xor b;
    layer3_outputs(7174) <= not a;
    layer3_outputs(7175) <= not b;
    layer3_outputs(7176) <= not b;
    layer3_outputs(7177) <= not a;
    layer3_outputs(7178) <= not (a and b);
    layer3_outputs(7179) <= not b;
    layer3_outputs(7180) <= not a;
    layer3_outputs(7181) <= not (a xor b);
    layer3_outputs(7182) <= not b or a;
    layer3_outputs(7183) <= a;
    layer3_outputs(7184) <= not b;
    layer3_outputs(7185) <= not b or a;
    layer3_outputs(7186) <= a xor b;
    layer3_outputs(7187) <= not (a xor b);
    layer3_outputs(7188) <= not (a or b);
    layer3_outputs(7189) <= not (a and b);
    layer3_outputs(7190) <= a;
    layer3_outputs(7191) <= a or b;
    layer3_outputs(7192) <= not (a xor b);
    layer3_outputs(7193) <= a;
    layer3_outputs(7194) <= not a;
    layer3_outputs(7195) <= not (a xor b);
    layer3_outputs(7196) <= a;
    layer3_outputs(7197) <= not (a and b);
    layer3_outputs(7198) <= not (a xor b);
    layer3_outputs(7199) <= not (a and b);
    layer3_outputs(7200) <= a and not b;
    layer3_outputs(7201) <= a;
    layer3_outputs(7202) <= a and not b;
    layer3_outputs(7203) <= b and not a;
    layer3_outputs(7204) <= not (a xor b);
    layer3_outputs(7205) <= a;
    layer3_outputs(7206) <= not (a or b);
    layer3_outputs(7207) <= b and not a;
    layer3_outputs(7208) <= not (a or b);
    layer3_outputs(7209) <= not b;
    layer3_outputs(7210) <= not b;
    layer3_outputs(7211) <= 1'b0;
    layer3_outputs(7212) <= a xor b;
    layer3_outputs(7213) <= a and not b;
    layer3_outputs(7214) <= not b or a;
    layer3_outputs(7215) <= not b;
    layer3_outputs(7216) <= b and not a;
    layer3_outputs(7217) <= a and not b;
    layer3_outputs(7218) <= a xor b;
    layer3_outputs(7219) <= not a;
    layer3_outputs(7220) <= a;
    layer3_outputs(7221) <= a and not b;
    layer3_outputs(7222) <= a or b;
    layer3_outputs(7223) <= a and not b;
    layer3_outputs(7224) <= not b;
    layer3_outputs(7225) <= not (a or b);
    layer3_outputs(7226) <= not (a or b);
    layer3_outputs(7227) <= a and b;
    layer3_outputs(7228) <= b and not a;
    layer3_outputs(7229) <= not b;
    layer3_outputs(7230) <= a xor b;
    layer3_outputs(7231) <= a or b;
    layer3_outputs(7232) <= a;
    layer3_outputs(7233) <= not (a or b);
    layer3_outputs(7234) <= a and not b;
    layer3_outputs(7235) <= a or b;
    layer3_outputs(7236) <= not b;
    layer3_outputs(7237) <= b;
    layer3_outputs(7238) <= not a;
    layer3_outputs(7239) <= not b or a;
    layer3_outputs(7240) <= not a;
    layer3_outputs(7241) <= a or b;
    layer3_outputs(7242) <= b;
    layer3_outputs(7243) <= a xor b;
    layer3_outputs(7244) <= b;
    layer3_outputs(7245) <= a;
    layer3_outputs(7246) <= not b;
    layer3_outputs(7247) <= not a;
    layer3_outputs(7248) <= not a;
    layer3_outputs(7249) <= not (a xor b);
    layer3_outputs(7250) <= b;
    layer3_outputs(7251) <= a and b;
    layer3_outputs(7252) <= not (a or b);
    layer3_outputs(7253) <= a and b;
    layer3_outputs(7254) <= a or b;
    layer3_outputs(7255) <= b;
    layer3_outputs(7256) <= not (a xor b);
    layer3_outputs(7257) <= a;
    layer3_outputs(7258) <= not (a or b);
    layer3_outputs(7259) <= not a;
    layer3_outputs(7260) <= not a;
    layer3_outputs(7261) <= not b;
    layer3_outputs(7262) <= not b;
    layer3_outputs(7263) <= a;
    layer3_outputs(7264) <= a and not b;
    layer3_outputs(7265) <= 1'b0;
    layer3_outputs(7266) <= a;
    layer3_outputs(7267) <= a;
    layer3_outputs(7268) <= not b or a;
    layer3_outputs(7269) <= a and b;
    layer3_outputs(7270) <= not (a and b);
    layer3_outputs(7271) <= b;
    layer3_outputs(7272) <= not a;
    layer3_outputs(7273) <= a;
    layer3_outputs(7274) <= not a;
    layer3_outputs(7275) <= a xor b;
    layer3_outputs(7276) <= not b;
    layer3_outputs(7277) <= not (a or b);
    layer3_outputs(7278) <= not a;
    layer3_outputs(7279) <= a;
    layer3_outputs(7280) <= not (a xor b);
    layer3_outputs(7281) <= not b;
    layer3_outputs(7282) <= not (a and b);
    layer3_outputs(7283) <= b;
    layer3_outputs(7284) <= a;
    layer3_outputs(7285) <= a and not b;
    layer3_outputs(7286) <= not a;
    layer3_outputs(7287) <= a and b;
    layer3_outputs(7288) <= not a;
    layer3_outputs(7289) <= a and b;
    layer3_outputs(7290) <= a;
    layer3_outputs(7291) <= 1'b0;
    layer3_outputs(7292) <= not b;
    layer3_outputs(7293) <= not a;
    layer3_outputs(7294) <= a and b;
    layer3_outputs(7295) <= a and b;
    layer3_outputs(7296) <= a xor b;
    layer3_outputs(7297) <= not a or b;
    layer3_outputs(7298) <= not (a or b);
    layer3_outputs(7299) <= b;
    layer3_outputs(7300) <= b;
    layer3_outputs(7301) <= not b;
    layer3_outputs(7302) <= b;
    layer3_outputs(7303) <= not (a or b);
    layer3_outputs(7304) <= not b;
    layer3_outputs(7305) <= a or b;
    layer3_outputs(7306) <= not a;
    layer3_outputs(7307) <= not a or b;
    layer3_outputs(7308) <= not a or b;
    layer3_outputs(7309) <= a or b;
    layer3_outputs(7310) <= not (a and b);
    layer3_outputs(7311) <= not b;
    layer3_outputs(7312) <= a and b;
    layer3_outputs(7313) <= not a;
    layer3_outputs(7314) <= not (a xor b);
    layer3_outputs(7315) <= b and not a;
    layer3_outputs(7316) <= a and b;
    layer3_outputs(7317) <= not (a xor b);
    layer3_outputs(7318) <= b;
    layer3_outputs(7319) <= not b;
    layer3_outputs(7320) <= not (a and b);
    layer3_outputs(7321) <= b and not a;
    layer3_outputs(7322) <= a and not b;
    layer3_outputs(7323) <= not (a and b);
    layer3_outputs(7324) <= not a;
    layer3_outputs(7325) <= not (a or b);
    layer3_outputs(7326) <= not (a xor b);
    layer3_outputs(7327) <= a or b;
    layer3_outputs(7328) <= not a;
    layer3_outputs(7329) <= not a;
    layer3_outputs(7330) <= a;
    layer3_outputs(7331) <= not b or a;
    layer3_outputs(7332) <= a and b;
    layer3_outputs(7333) <= not a;
    layer3_outputs(7334) <= not b;
    layer3_outputs(7335) <= a xor b;
    layer3_outputs(7336) <= a xor b;
    layer3_outputs(7337) <= not (a xor b);
    layer3_outputs(7338) <= not (a xor b);
    layer3_outputs(7339) <= b;
    layer3_outputs(7340) <= not (a or b);
    layer3_outputs(7341) <= not (a and b);
    layer3_outputs(7342) <= a and not b;
    layer3_outputs(7343) <= a and b;
    layer3_outputs(7344) <= not (a xor b);
    layer3_outputs(7345) <= a and not b;
    layer3_outputs(7346) <= 1'b0;
    layer3_outputs(7347) <= a and not b;
    layer3_outputs(7348) <= a;
    layer3_outputs(7349) <= a;
    layer3_outputs(7350) <= a;
    layer3_outputs(7351) <= not (a and b);
    layer3_outputs(7352) <= not a or b;
    layer3_outputs(7353) <= not a;
    layer3_outputs(7354) <= 1'b0;
    layer3_outputs(7355) <= not (a xor b);
    layer3_outputs(7356) <= not b;
    layer3_outputs(7357) <= a or b;
    layer3_outputs(7358) <= b;
    layer3_outputs(7359) <= b;
    layer3_outputs(7360) <= b;
    layer3_outputs(7361) <= a;
    layer3_outputs(7362) <= a and b;
    layer3_outputs(7363) <= a;
    layer3_outputs(7364) <= not (a xor b);
    layer3_outputs(7365) <= not a;
    layer3_outputs(7366) <= a;
    layer3_outputs(7367) <= not b;
    layer3_outputs(7368) <= not a;
    layer3_outputs(7369) <= not b;
    layer3_outputs(7370) <= a xor b;
    layer3_outputs(7371) <= b and not a;
    layer3_outputs(7372) <= not b;
    layer3_outputs(7373) <= b;
    layer3_outputs(7374) <= b and not a;
    layer3_outputs(7375) <= not a or b;
    layer3_outputs(7376) <= a and b;
    layer3_outputs(7377) <= a and not b;
    layer3_outputs(7378) <= not (a or b);
    layer3_outputs(7379) <= a or b;
    layer3_outputs(7380) <= not (a and b);
    layer3_outputs(7381) <= a or b;
    layer3_outputs(7382) <= not b;
    layer3_outputs(7383) <= not a;
    layer3_outputs(7384) <= b;
    layer3_outputs(7385) <= not b;
    layer3_outputs(7386) <= not a;
    layer3_outputs(7387) <= 1'b0;
    layer3_outputs(7388) <= a xor b;
    layer3_outputs(7389) <= a or b;
    layer3_outputs(7390) <= not a or b;
    layer3_outputs(7391) <= not a or b;
    layer3_outputs(7392) <= not a or b;
    layer3_outputs(7393) <= b;
    layer3_outputs(7394) <= not (a xor b);
    layer3_outputs(7395) <= not a;
    layer3_outputs(7396) <= not b or a;
    layer3_outputs(7397) <= not a;
    layer3_outputs(7398) <= a and not b;
    layer3_outputs(7399) <= not a or b;
    layer3_outputs(7400) <= a xor b;
    layer3_outputs(7401) <= a;
    layer3_outputs(7402) <= a and b;
    layer3_outputs(7403) <= not b;
    layer3_outputs(7404) <= a;
    layer3_outputs(7405) <= not (a xor b);
    layer3_outputs(7406) <= a or b;
    layer3_outputs(7407) <= a xor b;
    layer3_outputs(7408) <= not (a xor b);
    layer3_outputs(7409) <= a;
    layer3_outputs(7410) <= a or b;
    layer3_outputs(7411) <= b and not a;
    layer3_outputs(7412) <= not a or b;
    layer3_outputs(7413) <= not a;
    layer3_outputs(7414) <= not (a xor b);
    layer3_outputs(7415) <= a or b;
    layer3_outputs(7416) <= not (a xor b);
    layer3_outputs(7417) <= 1'b1;
    layer3_outputs(7418) <= not b or a;
    layer3_outputs(7419) <= a;
    layer3_outputs(7420) <= a or b;
    layer3_outputs(7421) <= not (a and b);
    layer3_outputs(7422) <= b and not a;
    layer3_outputs(7423) <= not b or a;
    layer3_outputs(7424) <= not (a xor b);
    layer3_outputs(7425) <= a xor b;
    layer3_outputs(7426) <= not a;
    layer3_outputs(7427) <= a;
    layer3_outputs(7428) <= not b or a;
    layer3_outputs(7429) <= b and not a;
    layer3_outputs(7430) <= a;
    layer3_outputs(7431) <= a and not b;
    layer3_outputs(7432) <= b;
    layer3_outputs(7433) <= not a;
    layer3_outputs(7434) <= not a;
    layer3_outputs(7435) <= b and not a;
    layer3_outputs(7436) <= a;
    layer3_outputs(7437) <= a;
    layer3_outputs(7438) <= b;
    layer3_outputs(7439) <= b and not a;
    layer3_outputs(7440) <= not (a xor b);
    layer3_outputs(7441) <= a;
    layer3_outputs(7442) <= b;
    layer3_outputs(7443) <= b;
    layer3_outputs(7444) <= not b;
    layer3_outputs(7445) <= b and not a;
    layer3_outputs(7446) <= a;
    layer3_outputs(7447) <= not (a or b);
    layer3_outputs(7448) <= a;
    layer3_outputs(7449) <= not b;
    layer3_outputs(7450) <= a xor b;
    layer3_outputs(7451) <= a;
    layer3_outputs(7452) <= not b;
    layer3_outputs(7453) <= not (a and b);
    layer3_outputs(7454) <= a;
    layer3_outputs(7455) <= a;
    layer3_outputs(7456) <= b;
    layer3_outputs(7457) <= not a;
    layer3_outputs(7458) <= not a;
    layer3_outputs(7459) <= not b or a;
    layer3_outputs(7460) <= 1'b0;
    layer3_outputs(7461) <= not a;
    layer3_outputs(7462) <= not (a xor b);
    layer3_outputs(7463) <= a;
    layer3_outputs(7464) <= not (a xor b);
    layer3_outputs(7465) <= not a;
    layer3_outputs(7466) <= not b;
    layer3_outputs(7467) <= b;
    layer3_outputs(7468) <= b;
    layer3_outputs(7469) <= not (a xor b);
    layer3_outputs(7470) <= not a;
    layer3_outputs(7471) <= b and not a;
    layer3_outputs(7472) <= a;
    layer3_outputs(7473) <= b;
    layer3_outputs(7474) <= a and b;
    layer3_outputs(7475) <= not (a xor b);
    layer3_outputs(7476) <= not b or a;
    layer3_outputs(7477) <= a xor b;
    layer3_outputs(7478) <= not b;
    layer3_outputs(7479) <= a or b;
    layer3_outputs(7480) <= not a;
    layer3_outputs(7481) <= b;
    layer3_outputs(7482) <= a or b;
    layer3_outputs(7483) <= b;
    layer3_outputs(7484) <= a;
    layer3_outputs(7485) <= a and not b;
    layer3_outputs(7486) <= a and b;
    layer3_outputs(7487) <= b;
    layer3_outputs(7488) <= a xor b;
    layer3_outputs(7489) <= a xor b;
    layer3_outputs(7490) <= not (a and b);
    layer3_outputs(7491) <= not (a or b);
    layer3_outputs(7492) <= b and not a;
    layer3_outputs(7493) <= not (a and b);
    layer3_outputs(7494) <= not (a xor b);
    layer3_outputs(7495) <= not (a and b);
    layer3_outputs(7496) <= a and b;
    layer3_outputs(7497) <= a;
    layer3_outputs(7498) <= b and not a;
    layer3_outputs(7499) <= not (a xor b);
    layer3_outputs(7500) <= b;
    layer3_outputs(7501) <= not b or a;
    layer3_outputs(7502) <= a and b;
    layer3_outputs(7503) <= not a;
    layer3_outputs(7504) <= a or b;
    layer3_outputs(7505) <= not b or a;
    layer3_outputs(7506) <= not b;
    layer3_outputs(7507) <= a or b;
    layer3_outputs(7508) <= a and not b;
    layer3_outputs(7509) <= not b or a;
    layer3_outputs(7510) <= b;
    layer3_outputs(7511) <= a or b;
    layer3_outputs(7512) <= not b or a;
    layer3_outputs(7513) <= b;
    layer3_outputs(7514) <= not b;
    layer3_outputs(7515) <= a;
    layer3_outputs(7516) <= not (a xor b);
    layer3_outputs(7517) <= not (a and b);
    layer3_outputs(7518) <= a and not b;
    layer3_outputs(7519) <= not (a and b);
    layer3_outputs(7520) <= a or b;
    layer3_outputs(7521) <= a;
    layer3_outputs(7522) <= a xor b;
    layer3_outputs(7523) <= b and not a;
    layer3_outputs(7524) <= a and b;
    layer3_outputs(7525) <= a;
    layer3_outputs(7526) <= b;
    layer3_outputs(7527) <= a;
    layer3_outputs(7528) <= not (a and b);
    layer3_outputs(7529) <= a and b;
    layer3_outputs(7530) <= a and b;
    layer3_outputs(7531) <= not (a xor b);
    layer3_outputs(7532) <= not a;
    layer3_outputs(7533) <= not b or a;
    layer3_outputs(7534) <= not a or b;
    layer3_outputs(7535) <= not (a and b);
    layer3_outputs(7536) <= not a or b;
    layer3_outputs(7537) <= b;
    layer3_outputs(7538) <= not b;
    layer3_outputs(7539) <= a xor b;
    layer3_outputs(7540) <= not b or a;
    layer3_outputs(7541) <= a;
    layer3_outputs(7542) <= not b;
    layer3_outputs(7543) <= not b;
    layer3_outputs(7544) <= a;
    layer3_outputs(7545) <= b;
    layer3_outputs(7546) <= not b;
    layer3_outputs(7547) <= b and not a;
    layer3_outputs(7548) <= a;
    layer3_outputs(7549) <= a xor b;
    layer3_outputs(7550) <= not (a or b);
    layer3_outputs(7551) <= a;
    layer3_outputs(7552) <= not b or a;
    layer3_outputs(7553) <= b;
    layer3_outputs(7554) <= b;
    layer3_outputs(7555) <= b;
    layer3_outputs(7556) <= not a;
    layer3_outputs(7557) <= not (a or b);
    layer3_outputs(7558) <= 1'b0;
    layer3_outputs(7559) <= a and not b;
    layer3_outputs(7560) <= not (a and b);
    layer3_outputs(7561) <= not a;
    layer3_outputs(7562) <= not (a and b);
    layer3_outputs(7563) <= not a or b;
    layer3_outputs(7564) <= not a;
    layer3_outputs(7565) <= b and not a;
    layer3_outputs(7566) <= b;
    layer3_outputs(7567) <= not (a or b);
    layer3_outputs(7568) <= a and not b;
    layer3_outputs(7569) <= b;
    layer3_outputs(7570) <= not a;
    layer3_outputs(7571) <= not (a xor b);
    layer3_outputs(7572) <= a;
    layer3_outputs(7573) <= not (a xor b);
    layer3_outputs(7574) <= a xor b;
    layer3_outputs(7575) <= b and not a;
    layer3_outputs(7576) <= b and not a;
    layer3_outputs(7577) <= not (a or b);
    layer3_outputs(7578) <= b and not a;
    layer3_outputs(7579) <= not (a and b);
    layer3_outputs(7580) <= b and not a;
    layer3_outputs(7581) <= not b;
    layer3_outputs(7582) <= b and not a;
    layer3_outputs(7583) <= a or b;
    layer3_outputs(7584) <= a;
    layer3_outputs(7585) <= b and not a;
    layer3_outputs(7586) <= a and b;
    layer3_outputs(7587) <= b;
    layer3_outputs(7588) <= b;
    layer3_outputs(7589) <= not b or a;
    layer3_outputs(7590) <= a;
    layer3_outputs(7591) <= not (a xor b);
    layer3_outputs(7592) <= b and not a;
    layer3_outputs(7593) <= not b or a;
    layer3_outputs(7594) <= b and not a;
    layer3_outputs(7595) <= not b or a;
    layer3_outputs(7596) <= not (a or b);
    layer3_outputs(7597) <= a xor b;
    layer3_outputs(7598) <= a and b;
    layer3_outputs(7599) <= a and not b;
    layer3_outputs(7600) <= a xor b;
    layer3_outputs(7601) <= not b;
    layer3_outputs(7602) <= not a or b;
    layer3_outputs(7603) <= b;
    layer3_outputs(7604) <= not (a or b);
    layer3_outputs(7605) <= a;
    layer3_outputs(7606) <= a xor b;
    layer3_outputs(7607) <= not b;
    layer3_outputs(7608) <= b and not a;
    layer3_outputs(7609) <= not (a or b);
    layer3_outputs(7610) <= not a;
    layer3_outputs(7611) <= not a or b;
    layer3_outputs(7612) <= a or b;
    layer3_outputs(7613) <= not b;
    layer3_outputs(7614) <= a;
    layer3_outputs(7615) <= b;
    layer3_outputs(7616) <= not b or a;
    layer3_outputs(7617) <= not a or b;
    layer3_outputs(7618) <= b;
    layer3_outputs(7619) <= a or b;
    layer3_outputs(7620) <= not (a or b);
    layer3_outputs(7621) <= not (a xor b);
    layer3_outputs(7622) <= a and b;
    layer3_outputs(7623) <= a and b;
    layer3_outputs(7624) <= not b;
    layer3_outputs(7625) <= not b;
    layer3_outputs(7626) <= a;
    layer3_outputs(7627) <= a and b;
    layer3_outputs(7628) <= 1'b0;
    layer3_outputs(7629) <= a and b;
    layer3_outputs(7630) <= not b;
    layer3_outputs(7631) <= not b;
    layer3_outputs(7632) <= a or b;
    layer3_outputs(7633) <= a or b;
    layer3_outputs(7634) <= a;
    layer3_outputs(7635) <= a or b;
    layer3_outputs(7636) <= not a;
    layer3_outputs(7637) <= not b;
    layer3_outputs(7638) <= not (a xor b);
    layer3_outputs(7639) <= not b;
    layer3_outputs(7640) <= a or b;
    layer3_outputs(7641) <= not b;
    layer3_outputs(7642) <= not b;
    layer3_outputs(7643) <= a and b;
    layer3_outputs(7644) <= not (a and b);
    layer3_outputs(7645) <= not a;
    layer3_outputs(7646) <= a xor b;
    layer3_outputs(7647) <= b and not a;
    layer3_outputs(7648) <= b;
    layer3_outputs(7649) <= a;
    layer3_outputs(7650) <= not b;
    layer3_outputs(7651) <= a;
    layer3_outputs(7652) <= a xor b;
    layer3_outputs(7653) <= not b;
    layer3_outputs(7654) <= not a;
    layer3_outputs(7655) <= a and b;
    layer3_outputs(7656) <= a and b;
    layer3_outputs(7657) <= a xor b;
    layer3_outputs(7658) <= not (a or b);
    layer3_outputs(7659) <= not a;
    layer3_outputs(7660) <= a;
    layer3_outputs(7661) <= a and not b;
    layer3_outputs(7662) <= not (a xor b);
    layer3_outputs(7663) <= b and not a;
    layer3_outputs(7664) <= not (a xor b);
    layer3_outputs(7665) <= not (a and b);
    layer3_outputs(7666) <= not (a xor b);
    layer3_outputs(7667) <= a or b;
    layer3_outputs(7668) <= not a;
    layer3_outputs(7669) <= a and not b;
    layer3_outputs(7670) <= not a or b;
    layer3_outputs(7671) <= not b;
    layer3_outputs(7672) <= b and not a;
    layer3_outputs(7673) <= a and not b;
    layer3_outputs(7674) <= b;
    layer3_outputs(7675) <= a and b;
    layer3_outputs(7676) <= not (a or b);
    layer3_outputs(7677) <= a;
    layer3_outputs(7678) <= not (a xor b);
    layer3_outputs(7679) <= not b or a;
    layer3_outputs(7680) <= b;
    layer3_outputs(7681) <= a and not b;
    layer3_outputs(7682) <= a;
    layer3_outputs(7683) <= not (a and b);
    layer3_outputs(7684) <= b;
    layer3_outputs(7685) <= not a or b;
    layer3_outputs(7686) <= not a or b;
    layer3_outputs(7687) <= a;
    layer3_outputs(7688) <= a xor b;
    layer3_outputs(7689) <= b;
    layer3_outputs(7690) <= b;
    layer3_outputs(7691) <= not b or a;
    layer3_outputs(7692) <= a xor b;
    layer3_outputs(7693) <= not a;
    layer3_outputs(7694) <= not (a or b);
    layer3_outputs(7695) <= not b or a;
    layer3_outputs(7696) <= not b;
    layer3_outputs(7697) <= a and not b;
    layer3_outputs(7698) <= not a or b;
    layer3_outputs(7699) <= not a;
    layer3_outputs(7700) <= not b;
    layer3_outputs(7701) <= a;
    layer3_outputs(7702) <= not (a or b);
    layer3_outputs(7703) <= a and not b;
    layer3_outputs(7704) <= not b or a;
    layer3_outputs(7705) <= a and not b;
    layer3_outputs(7706) <= not (a or b);
    layer3_outputs(7707) <= not b;
    layer3_outputs(7708) <= a xor b;
    layer3_outputs(7709) <= not (a or b);
    layer3_outputs(7710) <= b;
    layer3_outputs(7711) <= not b;
    layer3_outputs(7712) <= not a or b;
    layer3_outputs(7713) <= not (a xor b);
    layer3_outputs(7714) <= not (a xor b);
    layer3_outputs(7715) <= 1'b0;
    layer3_outputs(7716) <= not (a or b);
    layer3_outputs(7717) <= a;
    layer3_outputs(7718) <= not a;
    layer3_outputs(7719) <= a or b;
    layer3_outputs(7720) <= b;
    layer3_outputs(7721) <= b;
    layer3_outputs(7722) <= b and not a;
    layer3_outputs(7723) <= 1'b1;
    layer3_outputs(7724) <= a and not b;
    layer3_outputs(7725) <= a;
    layer3_outputs(7726) <= not (a xor b);
    layer3_outputs(7727) <= not a;
    layer3_outputs(7728) <= not b;
    layer3_outputs(7729) <= not (a xor b);
    layer3_outputs(7730) <= a;
    layer3_outputs(7731) <= not a;
    layer3_outputs(7732) <= b;
    layer3_outputs(7733) <= b;
    layer3_outputs(7734) <= b;
    layer3_outputs(7735) <= not a or b;
    layer3_outputs(7736) <= a xor b;
    layer3_outputs(7737) <= b;
    layer3_outputs(7738) <= b;
    layer3_outputs(7739) <= a xor b;
    layer3_outputs(7740) <= not (a xor b);
    layer3_outputs(7741) <= a;
    layer3_outputs(7742) <= b;
    layer3_outputs(7743) <= b;
    layer3_outputs(7744) <= not b;
    layer3_outputs(7745) <= a or b;
    layer3_outputs(7746) <= not a or b;
    layer3_outputs(7747) <= a and b;
    layer3_outputs(7748) <= not a;
    layer3_outputs(7749) <= a;
    layer3_outputs(7750) <= not a;
    layer3_outputs(7751) <= not b;
    layer3_outputs(7752) <= not a or b;
    layer3_outputs(7753) <= not b or a;
    layer3_outputs(7754) <= a;
    layer3_outputs(7755) <= not a;
    layer3_outputs(7756) <= not (a and b);
    layer3_outputs(7757) <= not b or a;
    layer3_outputs(7758) <= not a;
    layer3_outputs(7759) <= a;
    layer3_outputs(7760) <= a or b;
    layer3_outputs(7761) <= not b or a;
    layer3_outputs(7762) <= b;
    layer3_outputs(7763) <= not (a xor b);
    layer3_outputs(7764) <= b;
    layer3_outputs(7765) <= not b;
    layer3_outputs(7766) <= a or b;
    layer3_outputs(7767) <= not (a xor b);
    layer3_outputs(7768) <= not (a xor b);
    layer3_outputs(7769) <= a or b;
    layer3_outputs(7770) <= not (a or b);
    layer3_outputs(7771) <= b;
    layer3_outputs(7772) <= b;
    layer3_outputs(7773) <= a and b;
    layer3_outputs(7774) <= a or b;
    layer3_outputs(7775) <= not a or b;
    layer3_outputs(7776) <= not b;
    layer3_outputs(7777) <= a;
    layer3_outputs(7778) <= a and b;
    layer3_outputs(7779) <= not (a or b);
    layer3_outputs(7780) <= not (a xor b);
    layer3_outputs(7781) <= a or b;
    layer3_outputs(7782) <= a;
    layer3_outputs(7783) <= a and not b;
    layer3_outputs(7784) <= a;
    layer3_outputs(7785) <= not (a and b);
    layer3_outputs(7786) <= a xor b;
    layer3_outputs(7787) <= not (a and b);
    layer3_outputs(7788) <= not a;
    layer3_outputs(7789) <= a;
    layer3_outputs(7790) <= not (a or b);
    layer3_outputs(7791) <= not b or a;
    layer3_outputs(7792) <= not a or b;
    layer3_outputs(7793) <= a or b;
    layer3_outputs(7794) <= not (a and b);
    layer3_outputs(7795) <= a and b;
    layer3_outputs(7796) <= not a or b;
    layer3_outputs(7797) <= a and b;
    layer3_outputs(7798) <= not b;
    layer3_outputs(7799) <= b;
    layer3_outputs(7800) <= not a;
    layer3_outputs(7801) <= b;
    layer3_outputs(7802) <= b;
    layer3_outputs(7803) <= not b or a;
    layer3_outputs(7804) <= b;
    layer3_outputs(7805) <= not a or b;
    layer3_outputs(7806) <= a;
    layer3_outputs(7807) <= a and b;
    layer3_outputs(7808) <= b;
    layer3_outputs(7809) <= not a or b;
    layer3_outputs(7810) <= b;
    layer3_outputs(7811) <= a and b;
    layer3_outputs(7812) <= not (a and b);
    layer3_outputs(7813) <= not b or a;
    layer3_outputs(7814) <= not a;
    layer3_outputs(7815) <= not a or b;
    layer3_outputs(7816) <= not b or a;
    layer3_outputs(7817) <= b;
    layer3_outputs(7818) <= not a;
    layer3_outputs(7819) <= not a;
    layer3_outputs(7820) <= a and not b;
    layer3_outputs(7821) <= a;
    layer3_outputs(7822) <= b and not a;
    layer3_outputs(7823) <= a or b;
    layer3_outputs(7824) <= not b;
    layer3_outputs(7825) <= b;
    layer3_outputs(7826) <= b;
    layer3_outputs(7827) <= not b;
    layer3_outputs(7828) <= b and not a;
    layer3_outputs(7829) <= not a;
    layer3_outputs(7830) <= not b;
    layer3_outputs(7831) <= a and b;
    layer3_outputs(7832) <= not (a or b);
    layer3_outputs(7833) <= b and not a;
    layer3_outputs(7834) <= not a;
    layer3_outputs(7835) <= a;
    layer3_outputs(7836) <= a or b;
    layer3_outputs(7837) <= a and b;
    layer3_outputs(7838) <= not a;
    layer3_outputs(7839) <= a;
    layer3_outputs(7840) <= not a;
    layer3_outputs(7841) <= not a;
    layer3_outputs(7842) <= not (a or b);
    layer3_outputs(7843) <= not b or a;
    layer3_outputs(7844) <= a;
    layer3_outputs(7845) <= b;
    layer3_outputs(7846) <= not a;
    layer3_outputs(7847) <= b and not a;
    layer3_outputs(7848) <= not b;
    layer3_outputs(7849) <= not (a or b);
    layer3_outputs(7850) <= b and not a;
    layer3_outputs(7851) <= not a;
    layer3_outputs(7852) <= a;
    layer3_outputs(7853) <= b;
    layer3_outputs(7854) <= not a;
    layer3_outputs(7855) <= a xor b;
    layer3_outputs(7856) <= not (a xor b);
    layer3_outputs(7857) <= a;
    layer3_outputs(7858) <= not a;
    layer3_outputs(7859) <= not b or a;
    layer3_outputs(7860) <= not b;
    layer3_outputs(7861) <= a or b;
    layer3_outputs(7862) <= b and not a;
    layer3_outputs(7863) <= a and b;
    layer3_outputs(7864) <= not b;
    layer3_outputs(7865) <= a or b;
    layer3_outputs(7866) <= a xor b;
    layer3_outputs(7867) <= b;
    layer3_outputs(7868) <= 1'b1;
    layer3_outputs(7869) <= not b or a;
    layer3_outputs(7870) <= a;
    layer3_outputs(7871) <= a and b;
    layer3_outputs(7872) <= a and not b;
    layer3_outputs(7873) <= a or b;
    layer3_outputs(7874) <= not a or b;
    layer3_outputs(7875) <= not b;
    layer3_outputs(7876) <= b;
    layer3_outputs(7877) <= b;
    layer3_outputs(7878) <= b;
    layer3_outputs(7879) <= not b or a;
    layer3_outputs(7880) <= b;
    layer3_outputs(7881) <= b and not a;
    layer3_outputs(7882) <= a;
    layer3_outputs(7883) <= not a or b;
    layer3_outputs(7884) <= not (a and b);
    layer3_outputs(7885) <= a and not b;
    layer3_outputs(7886) <= a and b;
    layer3_outputs(7887) <= b;
    layer3_outputs(7888) <= not b;
    layer3_outputs(7889) <= not b;
    layer3_outputs(7890) <= not a;
    layer3_outputs(7891) <= a and not b;
    layer3_outputs(7892) <= a and not b;
    layer3_outputs(7893) <= a and b;
    layer3_outputs(7894) <= a;
    layer3_outputs(7895) <= a or b;
    layer3_outputs(7896) <= a;
    layer3_outputs(7897) <= b;
    layer3_outputs(7898) <= not (a and b);
    layer3_outputs(7899) <= not b;
    layer3_outputs(7900) <= not (a and b);
    layer3_outputs(7901) <= b;
    layer3_outputs(7902) <= 1'b1;
    layer3_outputs(7903) <= not a;
    layer3_outputs(7904) <= b;
    layer3_outputs(7905) <= not a;
    layer3_outputs(7906) <= b;
    layer3_outputs(7907) <= not b;
    layer3_outputs(7908) <= not a;
    layer3_outputs(7909) <= b and not a;
    layer3_outputs(7910) <= b and not a;
    layer3_outputs(7911) <= a;
    layer3_outputs(7912) <= a and b;
    layer3_outputs(7913) <= a and b;
    layer3_outputs(7914) <= a xor b;
    layer3_outputs(7915) <= b;
    layer3_outputs(7916) <= not (a and b);
    layer3_outputs(7917) <= b and not a;
    layer3_outputs(7918) <= a;
    layer3_outputs(7919) <= a and b;
    layer3_outputs(7920) <= b;
    layer3_outputs(7921) <= b;
    layer3_outputs(7922) <= 1'b0;
    layer3_outputs(7923) <= not b;
    layer3_outputs(7924) <= a;
    layer3_outputs(7925) <= a and not b;
    layer3_outputs(7926) <= not a;
    layer3_outputs(7927) <= not b or a;
    layer3_outputs(7928) <= b and not a;
    layer3_outputs(7929) <= a and b;
    layer3_outputs(7930) <= not (a and b);
    layer3_outputs(7931) <= b;
    layer3_outputs(7932) <= a and not b;
    layer3_outputs(7933) <= not (a xor b);
    layer3_outputs(7934) <= not b;
    layer3_outputs(7935) <= 1'b0;
    layer3_outputs(7936) <= not b or a;
    layer3_outputs(7937) <= a and not b;
    layer3_outputs(7938) <= a and b;
    layer3_outputs(7939) <= b;
    layer3_outputs(7940) <= not (a or b);
    layer3_outputs(7941) <= b;
    layer3_outputs(7942) <= not b;
    layer3_outputs(7943) <= a and b;
    layer3_outputs(7944) <= not (a or b);
    layer3_outputs(7945) <= not b;
    layer3_outputs(7946) <= a;
    layer3_outputs(7947) <= not (a xor b);
    layer3_outputs(7948) <= not (a and b);
    layer3_outputs(7949) <= a and b;
    layer3_outputs(7950) <= a and not b;
    layer3_outputs(7951) <= not b;
    layer3_outputs(7952) <= not b;
    layer3_outputs(7953) <= a and not b;
    layer3_outputs(7954) <= b;
    layer3_outputs(7955) <= b and not a;
    layer3_outputs(7956) <= a or b;
    layer3_outputs(7957) <= not (a or b);
    layer3_outputs(7958) <= b;
    layer3_outputs(7959) <= b;
    layer3_outputs(7960) <= a or b;
    layer3_outputs(7961) <= not a;
    layer3_outputs(7962) <= not b;
    layer3_outputs(7963) <= not b;
    layer3_outputs(7964) <= a and not b;
    layer3_outputs(7965) <= not a or b;
    layer3_outputs(7966) <= a;
    layer3_outputs(7967) <= a xor b;
    layer3_outputs(7968) <= b;
    layer3_outputs(7969) <= not b;
    layer3_outputs(7970) <= 1'b1;
    layer3_outputs(7971) <= not a or b;
    layer3_outputs(7972) <= not a;
    layer3_outputs(7973) <= not b or a;
    layer3_outputs(7974) <= b;
    layer3_outputs(7975) <= not (a xor b);
    layer3_outputs(7976) <= not b or a;
    layer3_outputs(7977) <= a and not b;
    layer3_outputs(7978) <= not (a xor b);
    layer3_outputs(7979) <= not b or a;
    layer3_outputs(7980) <= not b;
    layer3_outputs(7981) <= not a;
    layer3_outputs(7982) <= b;
    layer3_outputs(7983) <= a and b;
    layer3_outputs(7984) <= a or b;
    layer3_outputs(7985) <= 1'b1;
    layer3_outputs(7986) <= not (a xor b);
    layer3_outputs(7987) <= not a;
    layer3_outputs(7988) <= not b;
    layer3_outputs(7989) <= a or b;
    layer3_outputs(7990) <= not (a or b);
    layer3_outputs(7991) <= a and not b;
    layer3_outputs(7992) <= not b;
    layer3_outputs(7993) <= a;
    layer3_outputs(7994) <= a or b;
    layer3_outputs(7995) <= a and b;
    layer3_outputs(7996) <= a or b;
    layer3_outputs(7997) <= a and not b;
    layer3_outputs(7998) <= a and not b;
    layer3_outputs(7999) <= not b;
    layer3_outputs(8000) <= b and not a;
    layer3_outputs(8001) <= not a;
    layer3_outputs(8002) <= not (a xor b);
    layer3_outputs(8003) <= a;
    layer3_outputs(8004) <= b;
    layer3_outputs(8005) <= not (a or b);
    layer3_outputs(8006) <= a and b;
    layer3_outputs(8007) <= b and not a;
    layer3_outputs(8008) <= not a or b;
    layer3_outputs(8009) <= b and not a;
    layer3_outputs(8010) <= a or b;
    layer3_outputs(8011) <= 1'b0;
    layer3_outputs(8012) <= a and b;
    layer3_outputs(8013) <= not (a or b);
    layer3_outputs(8014) <= a xor b;
    layer3_outputs(8015) <= not a;
    layer3_outputs(8016) <= b and not a;
    layer3_outputs(8017) <= not a;
    layer3_outputs(8018) <= a;
    layer3_outputs(8019) <= a xor b;
    layer3_outputs(8020) <= a or b;
    layer3_outputs(8021) <= a xor b;
    layer3_outputs(8022) <= b and not a;
    layer3_outputs(8023) <= 1'b0;
    layer3_outputs(8024) <= not a;
    layer3_outputs(8025) <= a and b;
    layer3_outputs(8026) <= not b;
    layer3_outputs(8027) <= a and not b;
    layer3_outputs(8028) <= a or b;
    layer3_outputs(8029) <= not b;
    layer3_outputs(8030) <= b and not a;
    layer3_outputs(8031) <= not b or a;
    layer3_outputs(8032) <= not a;
    layer3_outputs(8033) <= not (a xor b);
    layer3_outputs(8034) <= not a or b;
    layer3_outputs(8035) <= a;
    layer3_outputs(8036) <= 1'b0;
    layer3_outputs(8037) <= a or b;
    layer3_outputs(8038) <= not (a and b);
    layer3_outputs(8039) <= b and not a;
    layer3_outputs(8040) <= not a;
    layer3_outputs(8041) <= not a or b;
    layer3_outputs(8042) <= a or b;
    layer3_outputs(8043) <= b and not a;
    layer3_outputs(8044) <= not (a xor b);
    layer3_outputs(8045) <= not a or b;
    layer3_outputs(8046) <= not (a and b);
    layer3_outputs(8047) <= a;
    layer3_outputs(8048) <= a and not b;
    layer3_outputs(8049) <= a xor b;
    layer3_outputs(8050) <= b;
    layer3_outputs(8051) <= not (a or b);
    layer3_outputs(8052) <= not b;
    layer3_outputs(8053) <= a or b;
    layer3_outputs(8054) <= not b;
    layer3_outputs(8055) <= not (a xor b);
    layer3_outputs(8056) <= b;
    layer3_outputs(8057) <= not b or a;
    layer3_outputs(8058) <= b;
    layer3_outputs(8059) <= not a or b;
    layer3_outputs(8060) <= not (a xor b);
    layer3_outputs(8061) <= not a;
    layer3_outputs(8062) <= b;
    layer3_outputs(8063) <= a;
    layer3_outputs(8064) <= a xor b;
    layer3_outputs(8065) <= b and not a;
    layer3_outputs(8066) <= a;
    layer3_outputs(8067) <= not a;
    layer3_outputs(8068) <= not a;
    layer3_outputs(8069) <= not (a and b);
    layer3_outputs(8070) <= not (a xor b);
    layer3_outputs(8071) <= 1'b1;
    layer3_outputs(8072) <= not b;
    layer3_outputs(8073) <= 1'b0;
    layer3_outputs(8074) <= a and not b;
    layer3_outputs(8075) <= not b;
    layer3_outputs(8076) <= a and b;
    layer3_outputs(8077) <= not b;
    layer3_outputs(8078) <= not (a xor b);
    layer3_outputs(8079) <= not (a and b);
    layer3_outputs(8080) <= not a;
    layer3_outputs(8081) <= not a;
    layer3_outputs(8082) <= a and not b;
    layer3_outputs(8083) <= a or b;
    layer3_outputs(8084) <= b;
    layer3_outputs(8085) <= b;
    layer3_outputs(8086) <= not b or a;
    layer3_outputs(8087) <= not b or a;
    layer3_outputs(8088) <= b and not a;
    layer3_outputs(8089) <= a and not b;
    layer3_outputs(8090) <= a or b;
    layer3_outputs(8091) <= not a or b;
    layer3_outputs(8092) <= b;
    layer3_outputs(8093) <= not (a and b);
    layer3_outputs(8094) <= b and not a;
    layer3_outputs(8095) <= a;
    layer3_outputs(8096) <= 1'b1;
    layer3_outputs(8097) <= not a or b;
    layer3_outputs(8098) <= not (a or b);
    layer3_outputs(8099) <= not a or b;
    layer3_outputs(8100) <= a and not b;
    layer3_outputs(8101) <= not a;
    layer3_outputs(8102) <= not b;
    layer3_outputs(8103) <= not b or a;
    layer3_outputs(8104) <= not a;
    layer3_outputs(8105) <= b;
    layer3_outputs(8106) <= a xor b;
    layer3_outputs(8107) <= b;
    layer3_outputs(8108) <= a xor b;
    layer3_outputs(8109) <= b and not a;
    layer3_outputs(8110) <= not b;
    layer3_outputs(8111) <= a and b;
    layer3_outputs(8112) <= not (a and b);
    layer3_outputs(8113) <= not a;
    layer3_outputs(8114) <= a xor b;
    layer3_outputs(8115) <= a or b;
    layer3_outputs(8116) <= a or b;
    layer3_outputs(8117) <= a;
    layer3_outputs(8118) <= not b or a;
    layer3_outputs(8119) <= a and b;
    layer3_outputs(8120) <= a and b;
    layer3_outputs(8121) <= not a or b;
    layer3_outputs(8122) <= a and b;
    layer3_outputs(8123) <= not (a xor b);
    layer3_outputs(8124) <= a and b;
    layer3_outputs(8125) <= not a;
    layer3_outputs(8126) <= a and b;
    layer3_outputs(8127) <= a;
    layer3_outputs(8128) <= not a or b;
    layer3_outputs(8129) <= not b or a;
    layer3_outputs(8130) <= not (a xor b);
    layer3_outputs(8131) <= a or b;
    layer3_outputs(8132) <= not b;
    layer3_outputs(8133) <= not b;
    layer3_outputs(8134) <= a and not b;
    layer3_outputs(8135) <= b;
    layer3_outputs(8136) <= not b;
    layer3_outputs(8137) <= not (a and b);
    layer3_outputs(8138) <= a;
    layer3_outputs(8139) <= b and not a;
    layer3_outputs(8140) <= a;
    layer3_outputs(8141) <= not a;
    layer3_outputs(8142) <= a and not b;
    layer3_outputs(8143) <= a xor b;
    layer3_outputs(8144) <= not b or a;
    layer3_outputs(8145) <= not a or b;
    layer3_outputs(8146) <= a;
    layer3_outputs(8147) <= not a or b;
    layer3_outputs(8148) <= not b or a;
    layer3_outputs(8149) <= not a;
    layer3_outputs(8150) <= a;
    layer3_outputs(8151) <= not b;
    layer3_outputs(8152) <= a;
    layer3_outputs(8153) <= not b;
    layer3_outputs(8154) <= not (a or b);
    layer3_outputs(8155) <= not (a and b);
    layer3_outputs(8156) <= b;
    layer3_outputs(8157) <= not b;
    layer3_outputs(8158) <= not b or a;
    layer3_outputs(8159) <= a;
    layer3_outputs(8160) <= not b;
    layer3_outputs(8161) <= not (a and b);
    layer3_outputs(8162) <= b;
    layer3_outputs(8163) <= 1'b0;
    layer3_outputs(8164) <= b;
    layer3_outputs(8165) <= not (a and b);
    layer3_outputs(8166) <= a or b;
    layer3_outputs(8167) <= a;
    layer3_outputs(8168) <= not a;
    layer3_outputs(8169) <= not (a or b);
    layer3_outputs(8170) <= b;
    layer3_outputs(8171) <= not b;
    layer3_outputs(8172) <= b and not a;
    layer3_outputs(8173) <= a and b;
    layer3_outputs(8174) <= 1'b0;
    layer3_outputs(8175) <= not (a xor b);
    layer3_outputs(8176) <= a xor b;
    layer3_outputs(8177) <= b;
    layer3_outputs(8178) <= b;
    layer3_outputs(8179) <= a or b;
    layer3_outputs(8180) <= not (a or b);
    layer3_outputs(8181) <= not (a or b);
    layer3_outputs(8182) <= not a;
    layer3_outputs(8183) <= not (a or b);
    layer3_outputs(8184) <= not b;
    layer3_outputs(8185) <= not (a and b);
    layer3_outputs(8186) <= b;
    layer3_outputs(8187) <= not a;
    layer3_outputs(8188) <= a;
    layer3_outputs(8189) <= a xor b;
    layer3_outputs(8190) <= not a;
    layer3_outputs(8191) <= b;
    layer3_outputs(8192) <= not a or b;
    layer3_outputs(8193) <= not b;
    layer3_outputs(8194) <= not b;
    layer3_outputs(8195) <= b and not a;
    layer3_outputs(8196) <= not a;
    layer3_outputs(8197) <= b and not a;
    layer3_outputs(8198) <= a xor b;
    layer3_outputs(8199) <= not (a xor b);
    layer3_outputs(8200) <= not a;
    layer3_outputs(8201) <= not (a or b);
    layer3_outputs(8202) <= not (a and b);
    layer3_outputs(8203) <= not a;
    layer3_outputs(8204) <= not (a and b);
    layer3_outputs(8205) <= not (a xor b);
    layer3_outputs(8206) <= b and not a;
    layer3_outputs(8207) <= a and not b;
    layer3_outputs(8208) <= a or b;
    layer3_outputs(8209) <= not a;
    layer3_outputs(8210) <= a;
    layer3_outputs(8211) <= b;
    layer3_outputs(8212) <= a;
    layer3_outputs(8213) <= not (a or b);
    layer3_outputs(8214) <= a xor b;
    layer3_outputs(8215) <= not a;
    layer3_outputs(8216) <= a xor b;
    layer3_outputs(8217) <= a and b;
    layer3_outputs(8218) <= not a;
    layer3_outputs(8219) <= not (a xor b);
    layer3_outputs(8220) <= a;
    layer3_outputs(8221) <= not a or b;
    layer3_outputs(8222) <= not a;
    layer3_outputs(8223) <= not (a and b);
    layer3_outputs(8224) <= not b;
    layer3_outputs(8225) <= not a;
    layer3_outputs(8226) <= a;
    layer3_outputs(8227) <= not a or b;
    layer3_outputs(8228) <= a or b;
    layer3_outputs(8229) <= 1'b0;
    layer3_outputs(8230) <= not (a and b);
    layer3_outputs(8231) <= a;
    layer3_outputs(8232) <= not a;
    layer3_outputs(8233) <= not (a and b);
    layer3_outputs(8234) <= not (a xor b);
    layer3_outputs(8235) <= not b;
    layer3_outputs(8236) <= not a or b;
    layer3_outputs(8237) <= b;
    layer3_outputs(8238) <= not (a or b);
    layer3_outputs(8239) <= a and not b;
    layer3_outputs(8240) <= not (a and b);
    layer3_outputs(8241) <= b and not a;
    layer3_outputs(8242) <= not b or a;
    layer3_outputs(8243) <= not a;
    layer3_outputs(8244) <= not b;
    layer3_outputs(8245) <= a;
    layer3_outputs(8246) <= not (a xor b);
    layer3_outputs(8247) <= a or b;
    layer3_outputs(8248) <= not (a or b);
    layer3_outputs(8249) <= a or b;
    layer3_outputs(8250) <= not b;
    layer3_outputs(8251) <= not (a xor b);
    layer3_outputs(8252) <= not a;
    layer3_outputs(8253) <= not (a and b);
    layer3_outputs(8254) <= a or b;
    layer3_outputs(8255) <= not b;
    layer3_outputs(8256) <= not a or b;
    layer3_outputs(8257) <= not b;
    layer3_outputs(8258) <= b;
    layer3_outputs(8259) <= not a;
    layer3_outputs(8260) <= not a;
    layer3_outputs(8261) <= b;
    layer3_outputs(8262) <= b;
    layer3_outputs(8263) <= not a or b;
    layer3_outputs(8264) <= not b;
    layer3_outputs(8265) <= not (a and b);
    layer3_outputs(8266) <= b;
    layer3_outputs(8267) <= not (a or b);
    layer3_outputs(8268) <= a;
    layer3_outputs(8269) <= a and not b;
    layer3_outputs(8270) <= not a;
    layer3_outputs(8271) <= not (a or b);
    layer3_outputs(8272) <= 1'b0;
    layer3_outputs(8273) <= not b;
    layer3_outputs(8274) <= not b;
    layer3_outputs(8275) <= not (a and b);
    layer3_outputs(8276) <= not (a xor b);
    layer3_outputs(8277) <= not b;
    layer3_outputs(8278) <= not b;
    layer3_outputs(8279) <= not a;
    layer3_outputs(8280) <= not b;
    layer3_outputs(8281) <= a or b;
    layer3_outputs(8282) <= a or b;
    layer3_outputs(8283) <= not (a xor b);
    layer3_outputs(8284) <= not b;
    layer3_outputs(8285) <= b;
    layer3_outputs(8286) <= not b;
    layer3_outputs(8287) <= not (a or b);
    layer3_outputs(8288) <= not (a or b);
    layer3_outputs(8289) <= a xor b;
    layer3_outputs(8290) <= not b;
    layer3_outputs(8291) <= not a or b;
    layer3_outputs(8292) <= a;
    layer3_outputs(8293) <= not a;
    layer3_outputs(8294) <= not (a xor b);
    layer3_outputs(8295) <= not (a and b);
    layer3_outputs(8296) <= not (a or b);
    layer3_outputs(8297) <= a and b;
    layer3_outputs(8298) <= not b or a;
    layer3_outputs(8299) <= a;
    layer3_outputs(8300) <= a or b;
    layer3_outputs(8301) <= not a;
    layer3_outputs(8302) <= a and not b;
    layer3_outputs(8303) <= not b or a;
    layer3_outputs(8304) <= a or b;
    layer3_outputs(8305) <= not (a or b);
    layer3_outputs(8306) <= b;
    layer3_outputs(8307) <= not (a or b);
    layer3_outputs(8308) <= not b or a;
    layer3_outputs(8309) <= a xor b;
    layer3_outputs(8310) <= a or b;
    layer3_outputs(8311) <= not a;
    layer3_outputs(8312) <= not (a xor b);
    layer3_outputs(8313) <= not (a or b);
    layer3_outputs(8314) <= a;
    layer3_outputs(8315) <= not a;
    layer3_outputs(8316) <= b;
    layer3_outputs(8317) <= a and b;
    layer3_outputs(8318) <= not b;
    layer3_outputs(8319) <= b;
    layer3_outputs(8320) <= not (a xor b);
    layer3_outputs(8321) <= a;
    layer3_outputs(8322) <= not (a and b);
    layer3_outputs(8323) <= not a;
    layer3_outputs(8324) <= not (a and b);
    layer3_outputs(8325) <= b and not a;
    layer3_outputs(8326) <= a and b;
    layer3_outputs(8327) <= not a;
    layer3_outputs(8328) <= not (a xor b);
    layer3_outputs(8329) <= not b;
    layer3_outputs(8330) <= not (a xor b);
    layer3_outputs(8331) <= a;
    layer3_outputs(8332) <= not a;
    layer3_outputs(8333) <= not a;
    layer3_outputs(8334) <= a;
    layer3_outputs(8335) <= a;
    layer3_outputs(8336) <= not b;
    layer3_outputs(8337) <= a and b;
    layer3_outputs(8338) <= a xor b;
    layer3_outputs(8339) <= not (a xor b);
    layer3_outputs(8340) <= not b;
    layer3_outputs(8341) <= not a;
    layer3_outputs(8342) <= not b;
    layer3_outputs(8343) <= a and not b;
    layer3_outputs(8344) <= not a;
    layer3_outputs(8345) <= a and b;
    layer3_outputs(8346) <= a xor b;
    layer3_outputs(8347) <= b;
    layer3_outputs(8348) <= not (a and b);
    layer3_outputs(8349) <= a;
    layer3_outputs(8350) <= a and not b;
    layer3_outputs(8351) <= a;
    layer3_outputs(8352) <= a;
    layer3_outputs(8353) <= not b;
    layer3_outputs(8354) <= not a;
    layer3_outputs(8355) <= not b;
    layer3_outputs(8356) <= b;
    layer3_outputs(8357) <= a and not b;
    layer3_outputs(8358) <= not b;
    layer3_outputs(8359) <= a xor b;
    layer3_outputs(8360) <= not b;
    layer3_outputs(8361) <= not b;
    layer3_outputs(8362) <= not (a or b);
    layer3_outputs(8363) <= not a or b;
    layer3_outputs(8364) <= not (a xor b);
    layer3_outputs(8365) <= a and b;
    layer3_outputs(8366) <= a xor b;
    layer3_outputs(8367) <= a;
    layer3_outputs(8368) <= not a;
    layer3_outputs(8369) <= not a;
    layer3_outputs(8370) <= a xor b;
    layer3_outputs(8371) <= b;
    layer3_outputs(8372) <= a and b;
    layer3_outputs(8373) <= b and not a;
    layer3_outputs(8374) <= a;
    layer3_outputs(8375) <= b and not a;
    layer3_outputs(8376) <= not (a or b);
    layer3_outputs(8377) <= b;
    layer3_outputs(8378) <= a;
    layer3_outputs(8379) <= b and not a;
    layer3_outputs(8380) <= b and not a;
    layer3_outputs(8381) <= not a;
    layer3_outputs(8382) <= b;
    layer3_outputs(8383) <= b;
    layer3_outputs(8384) <= not b;
    layer3_outputs(8385) <= a and b;
    layer3_outputs(8386) <= a;
    layer3_outputs(8387) <= not b or a;
    layer3_outputs(8388) <= not a or b;
    layer3_outputs(8389) <= a;
    layer3_outputs(8390) <= a and not b;
    layer3_outputs(8391) <= not b or a;
    layer3_outputs(8392) <= a or b;
    layer3_outputs(8393) <= not b;
    layer3_outputs(8394) <= 1'b1;
    layer3_outputs(8395) <= not a or b;
    layer3_outputs(8396) <= not a;
    layer3_outputs(8397) <= a;
    layer3_outputs(8398) <= b;
    layer3_outputs(8399) <= b;
    layer3_outputs(8400) <= a;
    layer3_outputs(8401) <= b;
    layer3_outputs(8402) <= a xor b;
    layer3_outputs(8403) <= b;
    layer3_outputs(8404) <= b and not a;
    layer3_outputs(8405) <= not a;
    layer3_outputs(8406) <= a;
    layer3_outputs(8407) <= not a;
    layer3_outputs(8408) <= not (a or b);
    layer3_outputs(8409) <= not a or b;
    layer3_outputs(8410) <= not (a or b);
    layer3_outputs(8411) <= a and not b;
    layer3_outputs(8412) <= b and not a;
    layer3_outputs(8413) <= not b;
    layer3_outputs(8414) <= not a;
    layer3_outputs(8415) <= b and not a;
    layer3_outputs(8416) <= not a;
    layer3_outputs(8417) <= b and not a;
    layer3_outputs(8418) <= b and not a;
    layer3_outputs(8419) <= b;
    layer3_outputs(8420) <= a;
    layer3_outputs(8421) <= a xor b;
    layer3_outputs(8422) <= not (a or b);
    layer3_outputs(8423) <= b;
    layer3_outputs(8424) <= b;
    layer3_outputs(8425) <= b;
    layer3_outputs(8426) <= not (a and b);
    layer3_outputs(8427) <= not a or b;
    layer3_outputs(8428) <= b;
    layer3_outputs(8429) <= not a;
    layer3_outputs(8430) <= not b;
    layer3_outputs(8431) <= a or b;
    layer3_outputs(8432) <= a;
    layer3_outputs(8433) <= a;
    layer3_outputs(8434) <= not (a xor b);
    layer3_outputs(8435) <= not b;
    layer3_outputs(8436) <= a and b;
    layer3_outputs(8437) <= not a;
    layer3_outputs(8438) <= not a or b;
    layer3_outputs(8439) <= not a;
    layer3_outputs(8440) <= not (a xor b);
    layer3_outputs(8441) <= b;
    layer3_outputs(8442) <= a xor b;
    layer3_outputs(8443) <= not b;
    layer3_outputs(8444) <= a or b;
    layer3_outputs(8445) <= b and not a;
    layer3_outputs(8446) <= b;
    layer3_outputs(8447) <= not (a or b);
    layer3_outputs(8448) <= a;
    layer3_outputs(8449) <= not a;
    layer3_outputs(8450) <= 1'b0;
    layer3_outputs(8451) <= a;
    layer3_outputs(8452) <= not b or a;
    layer3_outputs(8453) <= not b;
    layer3_outputs(8454) <= 1'b0;
    layer3_outputs(8455) <= b;
    layer3_outputs(8456) <= b;
    layer3_outputs(8457) <= not (a and b);
    layer3_outputs(8458) <= not b or a;
    layer3_outputs(8459) <= a and not b;
    layer3_outputs(8460) <= not (a xor b);
    layer3_outputs(8461) <= a or b;
    layer3_outputs(8462) <= not a or b;
    layer3_outputs(8463) <= not b;
    layer3_outputs(8464) <= a;
    layer3_outputs(8465) <= a or b;
    layer3_outputs(8466) <= b;
    layer3_outputs(8467) <= a and b;
    layer3_outputs(8468) <= not b;
    layer3_outputs(8469) <= not b;
    layer3_outputs(8470) <= a and b;
    layer3_outputs(8471) <= not (a xor b);
    layer3_outputs(8472) <= a xor b;
    layer3_outputs(8473) <= not (a or b);
    layer3_outputs(8474) <= a xor b;
    layer3_outputs(8475) <= b;
    layer3_outputs(8476) <= not b or a;
    layer3_outputs(8477) <= not b;
    layer3_outputs(8478) <= a;
    layer3_outputs(8479) <= not (a and b);
    layer3_outputs(8480) <= a;
    layer3_outputs(8481) <= not b;
    layer3_outputs(8482) <= not (a xor b);
    layer3_outputs(8483) <= a;
    layer3_outputs(8484) <= a;
    layer3_outputs(8485) <= b and not a;
    layer3_outputs(8486) <= a and b;
    layer3_outputs(8487) <= not b;
    layer3_outputs(8488) <= not a or b;
    layer3_outputs(8489) <= a;
    layer3_outputs(8490) <= not (a or b);
    layer3_outputs(8491) <= not a;
    layer3_outputs(8492) <= not (a and b);
    layer3_outputs(8493) <= a or b;
    layer3_outputs(8494) <= a or b;
    layer3_outputs(8495) <= not a;
    layer3_outputs(8496) <= not (a and b);
    layer3_outputs(8497) <= a xor b;
    layer3_outputs(8498) <= a;
    layer3_outputs(8499) <= not a;
    layer3_outputs(8500) <= not (a or b);
    layer3_outputs(8501) <= not a;
    layer3_outputs(8502) <= a;
    layer3_outputs(8503) <= a xor b;
    layer3_outputs(8504) <= not b;
    layer3_outputs(8505) <= a xor b;
    layer3_outputs(8506) <= not a;
    layer3_outputs(8507) <= b;
    layer3_outputs(8508) <= a and b;
    layer3_outputs(8509) <= not b;
    layer3_outputs(8510) <= not b or a;
    layer3_outputs(8511) <= a or b;
    layer3_outputs(8512) <= a or b;
    layer3_outputs(8513) <= a and b;
    layer3_outputs(8514) <= not b or a;
    layer3_outputs(8515) <= a;
    layer3_outputs(8516) <= b and not a;
    layer3_outputs(8517) <= not (a xor b);
    layer3_outputs(8518) <= a;
    layer3_outputs(8519) <= b;
    layer3_outputs(8520) <= b;
    layer3_outputs(8521) <= not b;
    layer3_outputs(8522) <= not a;
    layer3_outputs(8523) <= a xor b;
    layer3_outputs(8524) <= not a;
    layer3_outputs(8525) <= a and b;
    layer3_outputs(8526) <= not b;
    layer3_outputs(8527) <= a;
    layer3_outputs(8528) <= b and not a;
    layer3_outputs(8529) <= a xor b;
    layer3_outputs(8530) <= b;
    layer3_outputs(8531) <= a and not b;
    layer3_outputs(8532) <= not (a or b);
    layer3_outputs(8533) <= a;
    layer3_outputs(8534) <= not (a or b);
    layer3_outputs(8535) <= a;
    layer3_outputs(8536) <= not a or b;
    layer3_outputs(8537) <= b and not a;
    layer3_outputs(8538) <= a xor b;
    layer3_outputs(8539) <= not a or b;
    layer3_outputs(8540) <= a or b;
    layer3_outputs(8541) <= not b;
    layer3_outputs(8542) <= not (a and b);
    layer3_outputs(8543) <= not a;
    layer3_outputs(8544) <= not (a or b);
    layer3_outputs(8545) <= b and not a;
    layer3_outputs(8546) <= a or b;
    layer3_outputs(8547) <= b and not a;
    layer3_outputs(8548) <= b and not a;
    layer3_outputs(8549) <= a;
    layer3_outputs(8550) <= a and not b;
    layer3_outputs(8551) <= not a or b;
    layer3_outputs(8552) <= a or b;
    layer3_outputs(8553) <= not a;
    layer3_outputs(8554) <= not a;
    layer3_outputs(8555) <= a and not b;
    layer3_outputs(8556) <= 1'b0;
    layer3_outputs(8557) <= not b;
    layer3_outputs(8558) <= b;
    layer3_outputs(8559) <= b;
    layer3_outputs(8560) <= not b;
    layer3_outputs(8561) <= 1'b1;
    layer3_outputs(8562) <= a xor b;
    layer3_outputs(8563) <= not (a or b);
    layer3_outputs(8564) <= a or b;
    layer3_outputs(8565) <= not (a xor b);
    layer3_outputs(8566) <= b;
    layer3_outputs(8567) <= b and not a;
    layer3_outputs(8568) <= b and not a;
    layer3_outputs(8569) <= b;
    layer3_outputs(8570) <= b;
    layer3_outputs(8571) <= not b;
    layer3_outputs(8572) <= not b;
    layer3_outputs(8573) <= a and not b;
    layer3_outputs(8574) <= b and not a;
    layer3_outputs(8575) <= not a;
    layer3_outputs(8576) <= a or b;
    layer3_outputs(8577) <= a and not b;
    layer3_outputs(8578) <= not a;
    layer3_outputs(8579) <= a or b;
    layer3_outputs(8580) <= not b;
    layer3_outputs(8581) <= a;
    layer3_outputs(8582) <= not (a and b);
    layer3_outputs(8583) <= a xor b;
    layer3_outputs(8584) <= b and not a;
    layer3_outputs(8585) <= not a;
    layer3_outputs(8586) <= not a or b;
    layer3_outputs(8587) <= not a;
    layer3_outputs(8588) <= not b or a;
    layer3_outputs(8589) <= a;
    layer3_outputs(8590) <= b and not a;
    layer3_outputs(8591) <= not a or b;
    layer3_outputs(8592) <= not a;
    layer3_outputs(8593) <= a;
    layer3_outputs(8594) <= b;
    layer3_outputs(8595) <= not (a and b);
    layer3_outputs(8596) <= a or b;
    layer3_outputs(8597) <= b and not a;
    layer3_outputs(8598) <= a xor b;
    layer3_outputs(8599) <= a;
    layer3_outputs(8600) <= a;
    layer3_outputs(8601) <= a;
    layer3_outputs(8602) <= a;
    layer3_outputs(8603) <= b;
    layer3_outputs(8604) <= not (a xor b);
    layer3_outputs(8605) <= not b or a;
    layer3_outputs(8606) <= a;
    layer3_outputs(8607) <= a or b;
    layer3_outputs(8608) <= not (a or b);
    layer3_outputs(8609) <= b;
    layer3_outputs(8610) <= not (a or b);
    layer3_outputs(8611) <= not a;
    layer3_outputs(8612) <= a;
    layer3_outputs(8613) <= b;
    layer3_outputs(8614) <= not (a xor b);
    layer3_outputs(8615) <= not (a or b);
    layer3_outputs(8616) <= a or b;
    layer3_outputs(8617) <= a and b;
    layer3_outputs(8618) <= not (a xor b);
    layer3_outputs(8619) <= b;
    layer3_outputs(8620) <= not (a xor b);
    layer3_outputs(8621) <= not a or b;
    layer3_outputs(8622) <= b;
    layer3_outputs(8623) <= not (a or b);
    layer3_outputs(8624) <= 1'b1;
    layer3_outputs(8625) <= not a;
    layer3_outputs(8626) <= not a;
    layer3_outputs(8627) <= a;
    layer3_outputs(8628) <= not b;
    layer3_outputs(8629) <= a and b;
    layer3_outputs(8630) <= not (a xor b);
    layer3_outputs(8631) <= not b;
    layer3_outputs(8632) <= b and not a;
    layer3_outputs(8633) <= not (a and b);
    layer3_outputs(8634) <= not a;
    layer3_outputs(8635) <= b;
    layer3_outputs(8636) <= a xor b;
    layer3_outputs(8637) <= not (a and b);
    layer3_outputs(8638) <= a and not b;
    layer3_outputs(8639) <= a or b;
    layer3_outputs(8640) <= not a;
    layer3_outputs(8641) <= b;
    layer3_outputs(8642) <= b;
    layer3_outputs(8643) <= not (a or b);
    layer3_outputs(8644) <= not (a xor b);
    layer3_outputs(8645) <= b and not a;
    layer3_outputs(8646) <= b;
    layer3_outputs(8647) <= not (a or b);
    layer3_outputs(8648) <= b and not a;
    layer3_outputs(8649) <= a and not b;
    layer3_outputs(8650) <= a and b;
    layer3_outputs(8651) <= not (a xor b);
    layer3_outputs(8652) <= not a;
    layer3_outputs(8653) <= not b or a;
    layer3_outputs(8654) <= not (a and b);
    layer3_outputs(8655) <= not (a or b);
    layer3_outputs(8656) <= b;
    layer3_outputs(8657) <= a xor b;
    layer3_outputs(8658) <= b and not a;
    layer3_outputs(8659) <= not (a xor b);
    layer3_outputs(8660) <= a;
    layer3_outputs(8661) <= not (a xor b);
    layer3_outputs(8662) <= a and b;
    layer3_outputs(8663) <= not b;
    layer3_outputs(8664) <= b;
    layer3_outputs(8665) <= a;
    layer3_outputs(8666) <= not a;
    layer3_outputs(8667) <= a;
    layer3_outputs(8668) <= a and not b;
    layer3_outputs(8669) <= not b;
    layer3_outputs(8670) <= a or b;
    layer3_outputs(8671) <= b;
    layer3_outputs(8672) <= a or b;
    layer3_outputs(8673) <= not (a and b);
    layer3_outputs(8674) <= a and b;
    layer3_outputs(8675) <= not b;
    layer3_outputs(8676) <= not b;
    layer3_outputs(8677) <= a;
    layer3_outputs(8678) <= not (a and b);
    layer3_outputs(8679) <= b;
    layer3_outputs(8680) <= a xor b;
    layer3_outputs(8681) <= b and not a;
    layer3_outputs(8682) <= not (a and b);
    layer3_outputs(8683) <= not a;
    layer3_outputs(8684) <= b;
    layer3_outputs(8685) <= a;
    layer3_outputs(8686) <= not (a and b);
    layer3_outputs(8687) <= 1'b0;
    layer3_outputs(8688) <= a xor b;
    layer3_outputs(8689) <= b;
    layer3_outputs(8690) <= a and b;
    layer3_outputs(8691) <= b;
    layer3_outputs(8692) <= not a or b;
    layer3_outputs(8693) <= not (a xor b);
    layer3_outputs(8694) <= a xor b;
    layer3_outputs(8695) <= not a;
    layer3_outputs(8696) <= a and b;
    layer3_outputs(8697) <= not a;
    layer3_outputs(8698) <= not (a or b);
    layer3_outputs(8699) <= not b or a;
    layer3_outputs(8700) <= b;
    layer3_outputs(8701) <= not a;
    layer3_outputs(8702) <= a;
    layer3_outputs(8703) <= not a;
    layer3_outputs(8704) <= a;
    layer3_outputs(8705) <= a and b;
    layer3_outputs(8706) <= a;
    layer3_outputs(8707) <= a;
    layer3_outputs(8708) <= b;
    layer3_outputs(8709) <= not a or b;
    layer3_outputs(8710) <= not (a or b);
    layer3_outputs(8711) <= 1'b1;
    layer3_outputs(8712) <= b;
    layer3_outputs(8713) <= not (a and b);
    layer3_outputs(8714) <= b;
    layer3_outputs(8715) <= not a;
    layer3_outputs(8716) <= not a;
    layer3_outputs(8717) <= a or b;
    layer3_outputs(8718) <= b;
    layer3_outputs(8719) <= a or b;
    layer3_outputs(8720) <= b;
    layer3_outputs(8721) <= not (a xor b);
    layer3_outputs(8722) <= not b;
    layer3_outputs(8723) <= not a or b;
    layer3_outputs(8724) <= a;
    layer3_outputs(8725) <= a or b;
    layer3_outputs(8726) <= not a;
    layer3_outputs(8727) <= not b;
    layer3_outputs(8728) <= not a;
    layer3_outputs(8729) <= not a;
    layer3_outputs(8730) <= not b;
    layer3_outputs(8731) <= a and not b;
    layer3_outputs(8732) <= b;
    layer3_outputs(8733) <= not a or b;
    layer3_outputs(8734) <= not (a and b);
    layer3_outputs(8735) <= a;
    layer3_outputs(8736) <= not a or b;
    layer3_outputs(8737) <= b;
    layer3_outputs(8738) <= b;
    layer3_outputs(8739) <= b and not a;
    layer3_outputs(8740) <= b;
    layer3_outputs(8741) <= b and not a;
    layer3_outputs(8742) <= not b;
    layer3_outputs(8743) <= not a or b;
    layer3_outputs(8744) <= not (a or b);
    layer3_outputs(8745) <= a;
    layer3_outputs(8746) <= not b or a;
    layer3_outputs(8747) <= not a;
    layer3_outputs(8748) <= b;
    layer3_outputs(8749) <= not b;
    layer3_outputs(8750) <= b and not a;
    layer3_outputs(8751) <= not (a xor b);
    layer3_outputs(8752) <= a and b;
    layer3_outputs(8753) <= a;
    layer3_outputs(8754) <= not a;
    layer3_outputs(8755) <= not b;
    layer3_outputs(8756) <= not (a or b);
    layer3_outputs(8757) <= not (a or b);
    layer3_outputs(8758) <= not a;
    layer3_outputs(8759) <= not b or a;
    layer3_outputs(8760) <= not a;
    layer3_outputs(8761) <= a xor b;
    layer3_outputs(8762) <= a;
    layer3_outputs(8763) <= not a or b;
    layer3_outputs(8764) <= not a;
    layer3_outputs(8765) <= a;
    layer3_outputs(8766) <= not a or b;
    layer3_outputs(8767) <= 1'b1;
    layer3_outputs(8768) <= b and not a;
    layer3_outputs(8769) <= not a;
    layer3_outputs(8770) <= not b or a;
    layer3_outputs(8771) <= a;
    layer3_outputs(8772) <= not b or a;
    layer3_outputs(8773) <= a or b;
    layer3_outputs(8774) <= not a;
    layer3_outputs(8775) <= a and b;
    layer3_outputs(8776) <= not b;
    layer3_outputs(8777) <= not (a xor b);
    layer3_outputs(8778) <= not (a xor b);
    layer3_outputs(8779) <= not (a and b);
    layer3_outputs(8780) <= not a;
    layer3_outputs(8781) <= a or b;
    layer3_outputs(8782) <= not a;
    layer3_outputs(8783) <= not (a or b);
    layer3_outputs(8784) <= not (a or b);
    layer3_outputs(8785) <= not a;
    layer3_outputs(8786) <= a and not b;
    layer3_outputs(8787) <= a xor b;
    layer3_outputs(8788) <= a;
    layer3_outputs(8789) <= not a;
    layer3_outputs(8790) <= a and b;
    layer3_outputs(8791) <= a;
    layer3_outputs(8792) <= not b;
    layer3_outputs(8793) <= not b;
    layer3_outputs(8794) <= not (a xor b);
    layer3_outputs(8795) <= a or b;
    layer3_outputs(8796) <= a or b;
    layer3_outputs(8797) <= not (a xor b);
    layer3_outputs(8798) <= a and not b;
    layer3_outputs(8799) <= a;
    layer3_outputs(8800) <= a;
    layer3_outputs(8801) <= a;
    layer3_outputs(8802) <= b;
    layer3_outputs(8803) <= not (a xor b);
    layer3_outputs(8804) <= a xor b;
    layer3_outputs(8805) <= not (a xor b);
    layer3_outputs(8806) <= not a;
    layer3_outputs(8807) <= not b;
    layer3_outputs(8808) <= a xor b;
    layer3_outputs(8809) <= a and b;
    layer3_outputs(8810) <= 1'b1;
    layer3_outputs(8811) <= not a;
    layer3_outputs(8812) <= not (a xor b);
    layer3_outputs(8813) <= b;
    layer3_outputs(8814) <= not b or a;
    layer3_outputs(8815) <= not b;
    layer3_outputs(8816) <= b;
    layer3_outputs(8817) <= not b;
    layer3_outputs(8818) <= a;
    layer3_outputs(8819) <= b;
    layer3_outputs(8820) <= not (a and b);
    layer3_outputs(8821) <= b and not a;
    layer3_outputs(8822) <= not b;
    layer3_outputs(8823) <= a;
    layer3_outputs(8824) <= a;
    layer3_outputs(8825) <= not b or a;
    layer3_outputs(8826) <= not b;
    layer3_outputs(8827) <= a;
    layer3_outputs(8828) <= a and not b;
    layer3_outputs(8829) <= not a or b;
    layer3_outputs(8830) <= not a;
    layer3_outputs(8831) <= a xor b;
    layer3_outputs(8832) <= a;
    layer3_outputs(8833) <= not b;
    layer3_outputs(8834) <= a;
    layer3_outputs(8835) <= not a or b;
    layer3_outputs(8836) <= not b;
    layer3_outputs(8837) <= not b;
    layer3_outputs(8838) <= a or b;
    layer3_outputs(8839) <= a;
    layer3_outputs(8840) <= b;
    layer3_outputs(8841) <= not (a xor b);
    layer3_outputs(8842) <= not a or b;
    layer3_outputs(8843) <= a;
    layer3_outputs(8844) <= not b or a;
    layer3_outputs(8845) <= not (a and b);
    layer3_outputs(8846) <= not (a xor b);
    layer3_outputs(8847) <= b;
    layer3_outputs(8848) <= not a or b;
    layer3_outputs(8849) <= 1'b1;
    layer3_outputs(8850) <= b and not a;
    layer3_outputs(8851) <= a or b;
    layer3_outputs(8852) <= not a;
    layer3_outputs(8853) <= a xor b;
    layer3_outputs(8854) <= not a;
    layer3_outputs(8855) <= not (a or b);
    layer3_outputs(8856) <= not a;
    layer3_outputs(8857) <= b and not a;
    layer3_outputs(8858) <= a and b;
    layer3_outputs(8859) <= b;
    layer3_outputs(8860) <= not a;
    layer3_outputs(8861) <= a;
    layer3_outputs(8862) <= 1'b0;
    layer3_outputs(8863) <= not b or a;
    layer3_outputs(8864) <= not b;
    layer3_outputs(8865) <= a;
    layer3_outputs(8866) <= a;
    layer3_outputs(8867) <= b;
    layer3_outputs(8868) <= not b or a;
    layer3_outputs(8869) <= b and not a;
    layer3_outputs(8870) <= not (a xor b);
    layer3_outputs(8871) <= not a;
    layer3_outputs(8872) <= a;
    layer3_outputs(8873) <= b and not a;
    layer3_outputs(8874) <= not b;
    layer3_outputs(8875) <= a and not b;
    layer3_outputs(8876) <= a or b;
    layer3_outputs(8877) <= b;
    layer3_outputs(8878) <= a xor b;
    layer3_outputs(8879) <= a xor b;
    layer3_outputs(8880) <= a;
    layer3_outputs(8881) <= b;
    layer3_outputs(8882) <= not (a and b);
    layer3_outputs(8883) <= not (a and b);
    layer3_outputs(8884) <= not a;
    layer3_outputs(8885) <= a xor b;
    layer3_outputs(8886) <= not b;
    layer3_outputs(8887) <= not (a and b);
    layer3_outputs(8888) <= not (a and b);
    layer3_outputs(8889) <= b;
    layer3_outputs(8890) <= not a;
    layer3_outputs(8891) <= not (a and b);
    layer3_outputs(8892) <= 1'b1;
    layer3_outputs(8893) <= not b;
    layer3_outputs(8894) <= not a;
    layer3_outputs(8895) <= a and not b;
    layer3_outputs(8896) <= a and b;
    layer3_outputs(8897) <= not a;
    layer3_outputs(8898) <= not b;
    layer3_outputs(8899) <= a and b;
    layer3_outputs(8900) <= not (a xor b);
    layer3_outputs(8901) <= not b or a;
    layer3_outputs(8902) <= not a or b;
    layer3_outputs(8903) <= a xor b;
    layer3_outputs(8904) <= a;
    layer3_outputs(8905) <= not (a and b);
    layer3_outputs(8906) <= a xor b;
    layer3_outputs(8907) <= b;
    layer3_outputs(8908) <= a xor b;
    layer3_outputs(8909) <= not (a or b);
    layer3_outputs(8910) <= not a;
    layer3_outputs(8911) <= not (a xor b);
    layer3_outputs(8912) <= a xor b;
    layer3_outputs(8913) <= b and not a;
    layer3_outputs(8914) <= not b or a;
    layer3_outputs(8915) <= a;
    layer3_outputs(8916) <= a;
    layer3_outputs(8917) <= not a;
    layer3_outputs(8918) <= b and not a;
    layer3_outputs(8919) <= not b;
    layer3_outputs(8920) <= a xor b;
    layer3_outputs(8921) <= not b or a;
    layer3_outputs(8922) <= not a;
    layer3_outputs(8923) <= not (a xor b);
    layer3_outputs(8924) <= a xor b;
    layer3_outputs(8925) <= a;
    layer3_outputs(8926) <= a and not b;
    layer3_outputs(8927) <= b and not a;
    layer3_outputs(8928) <= a and not b;
    layer3_outputs(8929) <= not (a xor b);
    layer3_outputs(8930) <= a and not b;
    layer3_outputs(8931) <= a;
    layer3_outputs(8932) <= not (a xor b);
    layer3_outputs(8933) <= not a;
    layer3_outputs(8934) <= not (a and b);
    layer3_outputs(8935) <= not b or a;
    layer3_outputs(8936) <= not a;
    layer3_outputs(8937) <= a xor b;
    layer3_outputs(8938) <= b;
    layer3_outputs(8939) <= not b or a;
    layer3_outputs(8940) <= not b or a;
    layer3_outputs(8941) <= not a or b;
    layer3_outputs(8942) <= a;
    layer3_outputs(8943) <= not (a xor b);
    layer3_outputs(8944) <= not (a and b);
    layer3_outputs(8945) <= b and not a;
    layer3_outputs(8946) <= b;
    layer3_outputs(8947) <= not (a xor b);
    layer3_outputs(8948) <= not b;
    layer3_outputs(8949) <= b and not a;
    layer3_outputs(8950) <= not (a xor b);
    layer3_outputs(8951) <= not b;
    layer3_outputs(8952) <= not b;
    layer3_outputs(8953) <= b;
    layer3_outputs(8954) <= a;
    layer3_outputs(8955) <= a;
    layer3_outputs(8956) <= not (a and b);
    layer3_outputs(8957) <= a;
    layer3_outputs(8958) <= not a;
    layer3_outputs(8959) <= not b;
    layer3_outputs(8960) <= not a or b;
    layer3_outputs(8961) <= b;
    layer3_outputs(8962) <= not b;
    layer3_outputs(8963) <= not a;
    layer3_outputs(8964) <= not (a or b);
    layer3_outputs(8965) <= not a;
    layer3_outputs(8966) <= not b;
    layer3_outputs(8967) <= b;
    layer3_outputs(8968) <= b;
    layer3_outputs(8969) <= a;
    layer3_outputs(8970) <= not a;
    layer3_outputs(8971) <= not b or a;
    layer3_outputs(8972) <= a;
    layer3_outputs(8973) <= a and b;
    layer3_outputs(8974) <= not (a xor b);
    layer3_outputs(8975) <= a and b;
    layer3_outputs(8976) <= not a;
    layer3_outputs(8977) <= a or b;
    layer3_outputs(8978) <= a or b;
    layer3_outputs(8979) <= not a;
    layer3_outputs(8980) <= not a;
    layer3_outputs(8981) <= a and b;
    layer3_outputs(8982) <= not b;
    layer3_outputs(8983) <= not (a xor b);
    layer3_outputs(8984) <= a and b;
    layer3_outputs(8985) <= not b;
    layer3_outputs(8986) <= not a;
    layer3_outputs(8987) <= not (a or b);
    layer3_outputs(8988) <= a and not b;
    layer3_outputs(8989) <= not (a and b);
    layer3_outputs(8990) <= not b;
    layer3_outputs(8991) <= a;
    layer3_outputs(8992) <= not b or a;
    layer3_outputs(8993) <= a and b;
    layer3_outputs(8994) <= a and b;
    layer3_outputs(8995) <= not b or a;
    layer3_outputs(8996) <= 1'b1;
    layer3_outputs(8997) <= a or b;
    layer3_outputs(8998) <= not (a or b);
    layer3_outputs(8999) <= not (a and b);
    layer3_outputs(9000) <= not a;
    layer3_outputs(9001) <= b;
    layer3_outputs(9002) <= a;
    layer3_outputs(9003) <= a xor b;
    layer3_outputs(9004) <= not a;
    layer3_outputs(9005) <= a or b;
    layer3_outputs(9006) <= a or b;
    layer3_outputs(9007) <= not (a or b);
    layer3_outputs(9008) <= not a or b;
    layer3_outputs(9009) <= not (a xor b);
    layer3_outputs(9010) <= not (a xor b);
    layer3_outputs(9011) <= a xor b;
    layer3_outputs(9012) <= not (a or b);
    layer3_outputs(9013) <= a and not b;
    layer3_outputs(9014) <= not b;
    layer3_outputs(9015) <= not b or a;
    layer3_outputs(9016) <= a xor b;
    layer3_outputs(9017) <= not a;
    layer3_outputs(9018) <= b;
    layer3_outputs(9019) <= not (a or b);
    layer3_outputs(9020) <= a or b;
    layer3_outputs(9021) <= a;
    layer3_outputs(9022) <= not a;
    layer3_outputs(9023) <= not b;
    layer3_outputs(9024) <= not b;
    layer3_outputs(9025) <= b;
    layer3_outputs(9026) <= not (a xor b);
    layer3_outputs(9027) <= not (a xor b);
    layer3_outputs(9028) <= not b;
    layer3_outputs(9029) <= a or b;
    layer3_outputs(9030) <= b;
    layer3_outputs(9031) <= a and not b;
    layer3_outputs(9032) <= not b;
    layer3_outputs(9033) <= a;
    layer3_outputs(9034) <= a and b;
    layer3_outputs(9035) <= 1'b1;
    layer3_outputs(9036) <= a and b;
    layer3_outputs(9037) <= a;
    layer3_outputs(9038) <= not (a and b);
    layer3_outputs(9039) <= a and not b;
    layer3_outputs(9040) <= a or b;
    layer3_outputs(9041) <= not a or b;
    layer3_outputs(9042) <= not a;
    layer3_outputs(9043) <= a and b;
    layer3_outputs(9044) <= not (a or b);
    layer3_outputs(9045) <= not (a and b);
    layer3_outputs(9046) <= not b;
    layer3_outputs(9047) <= not b;
    layer3_outputs(9048) <= not a or b;
    layer3_outputs(9049) <= b;
    layer3_outputs(9050) <= not (a xor b);
    layer3_outputs(9051) <= a or b;
    layer3_outputs(9052) <= not b;
    layer3_outputs(9053) <= not b;
    layer3_outputs(9054) <= a and b;
    layer3_outputs(9055) <= a xor b;
    layer3_outputs(9056) <= 1'b0;
    layer3_outputs(9057) <= a and not b;
    layer3_outputs(9058) <= not b;
    layer3_outputs(9059) <= not (a or b);
    layer3_outputs(9060) <= not (a and b);
    layer3_outputs(9061) <= b;
    layer3_outputs(9062) <= a and b;
    layer3_outputs(9063) <= not b or a;
    layer3_outputs(9064) <= a and b;
    layer3_outputs(9065) <= a;
    layer3_outputs(9066) <= a and b;
    layer3_outputs(9067) <= a;
    layer3_outputs(9068) <= a or b;
    layer3_outputs(9069) <= a;
    layer3_outputs(9070) <= not b;
    layer3_outputs(9071) <= not b or a;
    layer3_outputs(9072) <= a and b;
    layer3_outputs(9073) <= not (a and b);
    layer3_outputs(9074) <= b and not a;
    layer3_outputs(9075) <= b;
    layer3_outputs(9076) <= a;
    layer3_outputs(9077) <= not b or a;
    layer3_outputs(9078) <= not a;
    layer3_outputs(9079) <= a;
    layer3_outputs(9080) <= a or b;
    layer3_outputs(9081) <= not a;
    layer3_outputs(9082) <= not b;
    layer3_outputs(9083) <= a and not b;
    layer3_outputs(9084) <= a and b;
    layer3_outputs(9085) <= a xor b;
    layer3_outputs(9086) <= not b or a;
    layer3_outputs(9087) <= not (a and b);
    layer3_outputs(9088) <= a;
    layer3_outputs(9089) <= a;
    layer3_outputs(9090) <= b and not a;
    layer3_outputs(9091) <= not (a and b);
    layer3_outputs(9092) <= b and not a;
    layer3_outputs(9093) <= b;
    layer3_outputs(9094) <= not a;
    layer3_outputs(9095) <= a;
    layer3_outputs(9096) <= a xor b;
    layer3_outputs(9097) <= not (a and b);
    layer3_outputs(9098) <= not a;
    layer3_outputs(9099) <= not (a and b);
    layer3_outputs(9100) <= not (a xor b);
    layer3_outputs(9101) <= not a or b;
    layer3_outputs(9102) <= not (a or b);
    layer3_outputs(9103) <= not a;
    layer3_outputs(9104) <= b;
    layer3_outputs(9105) <= a;
    layer3_outputs(9106) <= not (a or b);
    layer3_outputs(9107) <= b;
    layer3_outputs(9108) <= a and b;
    layer3_outputs(9109) <= not (a xor b);
    layer3_outputs(9110) <= a xor b;
    layer3_outputs(9111) <= a xor b;
    layer3_outputs(9112) <= not b or a;
    layer3_outputs(9113) <= not a or b;
    layer3_outputs(9114) <= not a or b;
    layer3_outputs(9115) <= not a;
    layer3_outputs(9116) <= not a;
    layer3_outputs(9117) <= a;
    layer3_outputs(9118) <= not (a and b);
    layer3_outputs(9119) <= not b;
    layer3_outputs(9120) <= not b or a;
    layer3_outputs(9121) <= 1'b1;
    layer3_outputs(9122) <= not b or a;
    layer3_outputs(9123) <= not (a xor b);
    layer3_outputs(9124) <= a;
    layer3_outputs(9125) <= not a;
    layer3_outputs(9126) <= a and b;
    layer3_outputs(9127) <= not a or b;
    layer3_outputs(9128) <= a;
    layer3_outputs(9129) <= b;
    layer3_outputs(9130) <= a xor b;
    layer3_outputs(9131) <= not b;
    layer3_outputs(9132) <= b;
    layer3_outputs(9133) <= a xor b;
    layer3_outputs(9134) <= a;
    layer3_outputs(9135) <= not a;
    layer3_outputs(9136) <= a and not b;
    layer3_outputs(9137) <= not a or b;
    layer3_outputs(9138) <= not a;
    layer3_outputs(9139) <= not b;
    layer3_outputs(9140) <= a or b;
    layer3_outputs(9141) <= not b or a;
    layer3_outputs(9142) <= b;
    layer3_outputs(9143) <= a;
    layer3_outputs(9144) <= b;
    layer3_outputs(9145) <= b;
    layer3_outputs(9146) <= not (a and b);
    layer3_outputs(9147) <= b and not a;
    layer3_outputs(9148) <= a;
    layer3_outputs(9149) <= not a;
    layer3_outputs(9150) <= b;
    layer3_outputs(9151) <= b;
    layer3_outputs(9152) <= b;
    layer3_outputs(9153) <= a xor b;
    layer3_outputs(9154) <= a xor b;
    layer3_outputs(9155) <= not b or a;
    layer3_outputs(9156) <= not b or a;
    layer3_outputs(9157) <= a or b;
    layer3_outputs(9158) <= a or b;
    layer3_outputs(9159) <= a and not b;
    layer3_outputs(9160) <= a;
    layer3_outputs(9161) <= not (a and b);
    layer3_outputs(9162) <= not a or b;
    layer3_outputs(9163) <= not a;
    layer3_outputs(9164) <= not a;
    layer3_outputs(9165) <= not b;
    layer3_outputs(9166) <= 1'b0;
    layer3_outputs(9167) <= 1'b0;
    layer3_outputs(9168) <= b;
    layer3_outputs(9169) <= b;
    layer3_outputs(9170) <= a xor b;
    layer3_outputs(9171) <= a;
    layer3_outputs(9172) <= not (a xor b);
    layer3_outputs(9173) <= a and b;
    layer3_outputs(9174) <= not b;
    layer3_outputs(9175) <= not a;
    layer3_outputs(9176) <= a and b;
    layer3_outputs(9177) <= b;
    layer3_outputs(9178) <= not b;
    layer3_outputs(9179) <= not b;
    layer3_outputs(9180) <= b and not a;
    layer3_outputs(9181) <= a;
    layer3_outputs(9182) <= not b or a;
    layer3_outputs(9183) <= not (a or b);
    layer3_outputs(9184) <= a and not b;
    layer3_outputs(9185) <= not b;
    layer3_outputs(9186) <= not a;
    layer3_outputs(9187) <= a and b;
    layer3_outputs(9188) <= a xor b;
    layer3_outputs(9189) <= a and b;
    layer3_outputs(9190) <= b and not a;
    layer3_outputs(9191) <= not (a and b);
    layer3_outputs(9192) <= a and b;
    layer3_outputs(9193) <= a or b;
    layer3_outputs(9194) <= a;
    layer3_outputs(9195) <= not b or a;
    layer3_outputs(9196) <= a and b;
    layer3_outputs(9197) <= a;
    layer3_outputs(9198) <= b;
    layer3_outputs(9199) <= not a;
    layer3_outputs(9200) <= a and not b;
    layer3_outputs(9201) <= not (a or b);
    layer3_outputs(9202) <= not a;
    layer3_outputs(9203) <= not b or a;
    layer3_outputs(9204) <= not b;
    layer3_outputs(9205) <= a and b;
    layer3_outputs(9206) <= not b;
    layer3_outputs(9207) <= not (a xor b);
    layer3_outputs(9208) <= not a or b;
    layer3_outputs(9209) <= not a;
    layer3_outputs(9210) <= not a;
    layer3_outputs(9211) <= not (a or b);
    layer3_outputs(9212) <= b;
    layer3_outputs(9213) <= a;
    layer3_outputs(9214) <= a or b;
    layer3_outputs(9215) <= a;
    layer3_outputs(9216) <= not b;
    layer3_outputs(9217) <= not a;
    layer3_outputs(9218) <= not b;
    layer3_outputs(9219) <= not b or a;
    layer3_outputs(9220) <= b;
    layer3_outputs(9221) <= not (a or b);
    layer3_outputs(9222) <= a;
    layer3_outputs(9223) <= not (a xor b);
    layer3_outputs(9224) <= b;
    layer3_outputs(9225) <= b;
    layer3_outputs(9226) <= a xor b;
    layer3_outputs(9227) <= not b or a;
    layer3_outputs(9228) <= a;
    layer3_outputs(9229) <= not a;
    layer3_outputs(9230) <= not b;
    layer3_outputs(9231) <= a and not b;
    layer3_outputs(9232) <= not (a or b);
    layer3_outputs(9233) <= not a;
    layer3_outputs(9234) <= 1'b1;
    layer3_outputs(9235) <= not (a and b);
    layer3_outputs(9236) <= not a;
    layer3_outputs(9237) <= not b;
    layer3_outputs(9238) <= b and not a;
    layer3_outputs(9239) <= a xor b;
    layer3_outputs(9240) <= a and b;
    layer3_outputs(9241) <= not b;
    layer3_outputs(9242) <= not (a or b);
    layer3_outputs(9243) <= 1'b0;
    layer3_outputs(9244) <= not b;
    layer3_outputs(9245) <= a or b;
    layer3_outputs(9246) <= not (a xor b);
    layer3_outputs(9247) <= a xor b;
    layer3_outputs(9248) <= not (a xor b);
    layer3_outputs(9249) <= a or b;
    layer3_outputs(9250) <= 1'b0;
    layer3_outputs(9251) <= a and not b;
    layer3_outputs(9252) <= not b;
    layer3_outputs(9253) <= not b;
    layer3_outputs(9254) <= b;
    layer3_outputs(9255) <= a;
    layer3_outputs(9256) <= not (a or b);
    layer3_outputs(9257) <= a and not b;
    layer3_outputs(9258) <= a;
    layer3_outputs(9259) <= a;
    layer3_outputs(9260) <= not b or a;
    layer3_outputs(9261) <= b;
    layer3_outputs(9262) <= a;
    layer3_outputs(9263) <= not a or b;
    layer3_outputs(9264) <= not a;
    layer3_outputs(9265) <= not b;
    layer3_outputs(9266) <= a or b;
    layer3_outputs(9267) <= a;
    layer3_outputs(9268) <= not b or a;
    layer3_outputs(9269) <= a;
    layer3_outputs(9270) <= not (a xor b);
    layer3_outputs(9271) <= not (a or b);
    layer3_outputs(9272) <= a or b;
    layer3_outputs(9273) <= not b;
    layer3_outputs(9274) <= a or b;
    layer3_outputs(9275) <= a xor b;
    layer3_outputs(9276) <= not (a or b);
    layer3_outputs(9277) <= b;
    layer3_outputs(9278) <= not a;
    layer3_outputs(9279) <= not b;
    layer3_outputs(9280) <= not (a xor b);
    layer3_outputs(9281) <= a and b;
    layer3_outputs(9282) <= not a;
    layer3_outputs(9283) <= a xor b;
    layer3_outputs(9284) <= not (a xor b);
    layer3_outputs(9285) <= b;
    layer3_outputs(9286) <= not (a xor b);
    layer3_outputs(9287) <= a or b;
    layer3_outputs(9288) <= a;
    layer3_outputs(9289) <= 1'b1;
    layer3_outputs(9290) <= not (a or b);
    layer3_outputs(9291) <= not (a and b);
    layer3_outputs(9292) <= 1'b1;
    layer3_outputs(9293) <= not (a xor b);
    layer3_outputs(9294) <= not a or b;
    layer3_outputs(9295) <= b;
    layer3_outputs(9296) <= not b or a;
    layer3_outputs(9297) <= not a;
    layer3_outputs(9298) <= b;
    layer3_outputs(9299) <= not b or a;
    layer3_outputs(9300) <= not (a xor b);
    layer3_outputs(9301) <= not (a and b);
    layer3_outputs(9302) <= a;
    layer3_outputs(9303) <= a or b;
    layer3_outputs(9304) <= not (a xor b);
    layer3_outputs(9305) <= not (a or b);
    layer3_outputs(9306) <= b;
    layer3_outputs(9307) <= not a;
    layer3_outputs(9308) <= not a or b;
    layer3_outputs(9309) <= a xor b;
    layer3_outputs(9310) <= a xor b;
    layer3_outputs(9311) <= b and not a;
    layer3_outputs(9312) <= not (a and b);
    layer3_outputs(9313) <= not (a or b);
    layer3_outputs(9314) <= b and not a;
    layer3_outputs(9315) <= b;
    layer3_outputs(9316) <= not (a xor b);
    layer3_outputs(9317) <= b;
    layer3_outputs(9318) <= a;
    layer3_outputs(9319) <= a and b;
    layer3_outputs(9320) <= not b or a;
    layer3_outputs(9321) <= a and not b;
    layer3_outputs(9322) <= not (a and b);
    layer3_outputs(9323) <= not a or b;
    layer3_outputs(9324) <= not (a xor b);
    layer3_outputs(9325) <= not b or a;
    layer3_outputs(9326) <= not b;
    layer3_outputs(9327) <= not (a xor b);
    layer3_outputs(9328) <= not b;
    layer3_outputs(9329) <= a and not b;
    layer3_outputs(9330) <= not (a xor b);
    layer3_outputs(9331) <= not (a and b);
    layer3_outputs(9332) <= a;
    layer3_outputs(9333) <= a and b;
    layer3_outputs(9334) <= b;
    layer3_outputs(9335) <= not b;
    layer3_outputs(9336) <= b;
    layer3_outputs(9337) <= a and not b;
    layer3_outputs(9338) <= b;
    layer3_outputs(9339) <= a xor b;
    layer3_outputs(9340) <= 1'b1;
    layer3_outputs(9341) <= not (a or b);
    layer3_outputs(9342) <= not b;
    layer3_outputs(9343) <= not a or b;
    layer3_outputs(9344) <= not a;
    layer3_outputs(9345) <= a or b;
    layer3_outputs(9346) <= not (a and b);
    layer3_outputs(9347) <= b;
    layer3_outputs(9348) <= not a;
    layer3_outputs(9349) <= not b;
    layer3_outputs(9350) <= b;
    layer3_outputs(9351) <= a;
    layer3_outputs(9352) <= a and b;
    layer3_outputs(9353) <= not (a or b);
    layer3_outputs(9354) <= b;
    layer3_outputs(9355) <= b and not a;
    layer3_outputs(9356) <= a and b;
    layer3_outputs(9357) <= a;
    layer3_outputs(9358) <= not b or a;
    layer3_outputs(9359) <= not a or b;
    layer3_outputs(9360) <= not b;
    layer3_outputs(9361) <= a or b;
    layer3_outputs(9362) <= not (a or b);
    layer3_outputs(9363) <= 1'b0;
    layer3_outputs(9364) <= b and not a;
    layer3_outputs(9365) <= a and not b;
    layer3_outputs(9366) <= not b;
    layer3_outputs(9367) <= a or b;
    layer3_outputs(9368) <= not b or a;
    layer3_outputs(9369) <= not a;
    layer3_outputs(9370) <= b;
    layer3_outputs(9371) <= not (a or b);
    layer3_outputs(9372) <= not (a and b);
    layer3_outputs(9373) <= a and b;
    layer3_outputs(9374) <= b and not a;
    layer3_outputs(9375) <= b;
    layer3_outputs(9376) <= a and not b;
    layer3_outputs(9377) <= a and not b;
    layer3_outputs(9378) <= b;
    layer3_outputs(9379) <= not a or b;
    layer3_outputs(9380) <= not a or b;
    layer3_outputs(9381) <= not b;
    layer3_outputs(9382) <= not b;
    layer3_outputs(9383) <= b;
    layer3_outputs(9384) <= not a or b;
    layer3_outputs(9385) <= a;
    layer3_outputs(9386) <= 1'b0;
    layer3_outputs(9387) <= a and b;
    layer3_outputs(9388) <= b;
    layer3_outputs(9389) <= a;
    layer3_outputs(9390) <= a or b;
    layer3_outputs(9391) <= not a or b;
    layer3_outputs(9392) <= not b;
    layer3_outputs(9393) <= a and not b;
    layer3_outputs(9394) <= not (a or b);
    layer3_outputs(9395) <= not (a xor b);
    layer3_outputs(9396) <= not (a xor b);
    layer3_outputs(9397) <= not b or a;
    layer3_outputs(9398) <= a;
    layer3_outputs(9399) <= not (a and b);
    layer3_outputs(9400) <= not a;
    layer3_outputs(9401) <= not (a xor b);
    layer3_outputs(9402) <= not b or a;
    layer3_outputs(9403) <= not a;
    layer3_outputs(9404) <= not b or a;
    layer3_outputs(9405) <= b;
    layer3_outputs(9406) <= a;
    layer3_outputs(9407) <= a and b;
    layer3_outputs(9408) <= not b or a;
    layer3_outputs(9409) <= a xor b;
    layer3_outputs(9410) <= not b;
    layer3_outputs(9411) <= a and b;
    layer3_outputs(9412) <= not a or b;
    layer3_outputs(9413) <= not (a and b);
    layer3_outputs(9414) <= b and not a;
    layer3_outputs(9415) <= not (a xor b);
    layer3_outputs(9416) <= not a;
    layer3_outputs(9417) <= not a;
    layer3_outputs(9418) <= a and not b;
    layer3_outputs(9419) <= a;
    layer3_outputs(9420) <= not a or b;
    layer3_outputs(9421) <= a;
    layer3_outputs(9422) <= a;
    layer3_outputs(9423) <= not a;
    layer3_outputs(9424) <= not (a and b);
    layer3_outputs(9425) <= b;
    layer3_outputs(9426) <= a or b;
    layer3_outputs(9427) <= not (a xor b);
    layer3_outputs(9428) <= 1'b0;
    layer3_outputs(9429) <= b;
    layer3_outputs(9430) <= a;
    layer3_outputs(9431) <= not (a or b);
    layer3_outputs(9432) <= b and not a;
    layer3_outputs(9433) <= not (a xor b);
    layer3_outputs(9434) <= b and not a;
    layer3_outputs(9435) <= a or b;
    layer3_outputs(9436) <= not a;
    layer3_outputs(9437) <= b;
    layer3_outputs(9438) <= a or b;
    layer3_outputs(9439) <= not a;
    layer3_outputs(9440) <= not a;
    layer3_outputs(9441) <= not (a xor b);
    layer3_outputs(9442) <= not (a xor b);
    layer3_outputs(9443) <= a;
    layer3_outputs(9444) <= not a;
    layer3_outputs(9445) <= b and not a;
    layer3_outputs(9446) <= not b;
    layer3_outputs(9447) <= not b or a;
    layer3_outputs(9448) <= a;
    layer3_outputs(9449) <= not b;
    layer3_outputs(9450) <= not (a or b);
    layer3_outputs(9451) <= not (a xor b);
    layer3_outputs(9452) <= not (a or b);
    layer3_outputs(9453) <= a;
    layer3_outputs(9454) <= b;
    layer3_outputs(9455) <= b;
    layer3_outputs(9456) <= a and b;
    layer3_outputs(9457) <= a or b;
    layer3_outputs(9458) <= not b;
    layer3_outputs(9459) <= not b;
    layer3_outputs(9460) <= a;
    layer3_outputs(9461) <= not (a and b);
    layer3_outputs(9462) <= a xor b;
    layer3_outputs(9463) <= 1'b1;
    layer3_outputs(9464) <= a and not b;
    layer3_outputs(9465) <= not (a or b);
    layer3_outputs(9466) <= a and b;
    layer3_outputs(9467) <= not (a or b);
    layer3_outputs(9468) <= a;
    layer3_outputs(9469) <= a xor b;
    layer3_outputs(9470) <= b;
    layer3_outputs(9471) <= a;
    layer3_outputs(9472) <= not a or b;
    layer3_outputs(9473) <= a;
    layer3_outputs(9474) <= not b;
    layer3_outputs(9475) <= not (a xor b);
    layer3_outputs(9476) <= not a;
    layer3_outputs(9477) <= b and not a;
    layer3_outputs(9478) <= a;
    layer3_outputs(9479) <= not b;
    layer3_outputs(9480) <= a and not b;
    layer3_outputs(9481) <= a;
    layer3_outputs(9482) <= not b;
    layer3_outputs(9483) <= a;
    layer3_outputs(9484) <= a or b;
    layer3_outputs(9485) <= not (a or b);
    layer3_outputs(9486) <= a;
    layer3_outputs(9487) <= a or b;
    layer3_outputs(9488) <= not (a xor b);
    layer3_outputs(9489) <= a or b;
    layer3_outputs(9490) <= a or b;
    layer3_outputs(9491) <= a and b;
    layer3_outputs(9492) <= not a;
    layer3_outputs(9493) <= a and not b;
    layer3_outputs(9494) <= not a or b;
    layer3_outputs(9495) <= a;
    layer3_outputs(9496) <= a or b;
    layer3_outputs(9497) <= 1'b0;
    layer3_outputs(9498) <= not a or b;
    layer3_outputs(9499) <= b and not a;
    layer3_outputs(9500) <= b;
    layer3_outputs(9501) <= 1'b0;
    layer3_outputs(9502) <= a and b;
    layer3_outputs(9503) <= not (a or b);
    layer3_outputs(9504) <= a;
    layer3_outputs(9505) <= b;
    layer3_outputs(9506) <= b and not a;
    layer3_outputs(9507) <= not a;
    layer3_outputs(9508) <= a or b;
    layer3_outputs(9509) <= a or b;
    layer3_outputs(9510) <= a and not b;
    layer3_outputs(9511) <= b and not a;
    layer3_outputs(9512) <= not a;
    layer3_outputs(9513) <= a;
    layer3_outputs(9514) <= a and b;
    layer3_outputs(9515) <= not (a or b);
    layer3_outputs(9516) <= a;
    layer3_outputs(9517) <= not (a xor b);
    layer3_outputs(9518) <= b;
    layer3_outputs(9519) <= not a;
    layer3_outputs(9520) <= a xor b;
    layer3_outputs(9521) <= not b or a;
    layer3_outputs(9522) <= a;
    layer3_outputs(9523) <= not a;
    layer3_outputs(9524) <= a;
    layer3_outputs(9525) <= b;
    layer3_outputs(9526) <= not (a xor b);
    layer3_outputs(9527) <= a or b;
    layer3_outputs(9528) <= b and not a;
    layer3_outputs(9529) <= a or b;
    layer3_outputs(9530) <= not (a and b);
    layer3_outputs(9531) <= not a;
    layer3_outputs(9532) <= a or b;
    layer3_outputs(9533) <= not a;
    layer3_outputs(9534) <= a and not b;
    layer3_outputs(9535) <= not (a xor b);
    layer3_outputs(9536) <= b;
    layer3_outputs(9537) <= not b;
    layer3_outputs(9538) <= not b or a;
    layer3_outputs(9539) <= a;
    layer3_outputs(9540) <= b and not a;
    layer3_outputs(9541) <= not (a xor b);
    layer3_outputs(9542) <= a;
    layer3_outputs(9543) <= not b;
    layer3_outputs(9544) <= a;
    layer3_outputs(9545) <= not b or a;
    layer3_outputs(9546) <= not a;
    layer3_outputs(9547) <= a or b;
    layer3_outputs(9548) <= b and not a;
    layer3_outputs(9549) <= not (a or b);
    layer3_outputs(9550) <= not b;
    layer3_outputs(9551) <= not a;
    layer3_outputs(9552) <= a and b;
    layer3_outputs(9553) <= not b;
    layer3_outputs(9554) <= not b;
    layer3_outputs(9555) <= not (a xor b);
    layer3_outputs(9556) <= not a;
    layer3_outputs(9557) <= not a;
    layer3_outputs(9558) <= b;
    layer3_outputs(9559) <= a;
    layer3_outputs(9560) <= a;
    layer3_outputs(9561) <= a;
    layer3_outputs(9562) <= not b;
    layer3_outputs(9563) <= b;
    layer3_outputs(9564) <= not (a xor b);
    layer3_outputs(9565) <= a and not b;
    layer3_outputs(9566) <= b;
    layer3_outputs(9567) <= not (a xor b);
    layer3_outputs(9568) <= not a or b;
    layer3_outputs(9569) <= not (a and b);
    layer3_outputs(9570) <= not (a and b);
    layer3_outputs(9571) <= a or b;
    layer3_outputs(9572) <= not (a or b);
    layer3_outputs(9573) <= a and not b;
    layer3_outputs(9574) <= a;
    layer3_outputs(9575) <= not (a or b);
    layer3_outputs(9576) <= a;
    layer3_outputs(9577) <= not a;
    layer3_outputs(9578) <= not a;
    layer3_outputs(9579) <= a or b;
    layer3_outputs(9580) <= a xor b;
    layer3_outputs(9581) <= a and b;
    layer3_outputs(9582) <= b;
    layer3_outputs(9583) <= not (a and b);
    layer3_outputs(9584) <= a xor b;
    layer3_outputs(9585) <= a;
    layer3_outputs(9586) <= not (a and b);
    layer3_outputs(9587) <= not a;
    layer3_outputs(9588) <= not a;
    layer3_outputs(9589) <= b and not a;
    layer3_outputs(9590) <= not a or b;
    layer3_outputs(9591) <= not a;
    layer3_outputs(9592) <= not a;
    layer3_outputs(9593) <= a;
    layer3_outputs(9594) <= a;
    layer3_outputs(9595) <= not b;
    layer3_outputs(9596) <= not b or a;
    layer3_outputs(9597) <= not (a or b);
    layer3_outputs(9598) <= a or b;
    layer3_outputs(9599) <= b;
    layer3_outputs(9600) <= b;
    layer3_outputs(9601) <= a;
    layer3_outputs(9602) <= b;
    layer3_outputs(9603) <= b;
    layer3_outputs(9604) <= b;
    layer3_outputs(9605) <= not (a or b);
    layer3_outputs(9606) <= b and not a;
    layer3_outputs(9607) <= not (a or b);
    layer3_outputs(9608) <= not b or a;
    layer3_outputs(9609) <= a and not b;
    layer3_outputs(9610) <= a xor b;
    layer3_outputs(9611) <= not (a or b);
    layer3_outputs(9612) <= a and b;
    layer3_outputs(9613) <= a or b;
    layer3_outputs(9614) <= not a;
    layer3_outputs(9615) <= a and not b;
    layer3_outputs(9616) <= b;
    layer3_outputs(9617) <= not b or a;
    layer3_outputs(9618) <= a and b;
    layer3_outputs(9619) <= a xor b;
    layer3_outputs(9620) <= not b or a;
    layer3_outputs(9621) <= a;
    layer3_outputs(9622) <= not (a xor b);
    layer3_outputs(9623) <= not a or b;
    layer3_outputs(9624) <= a;
    layer3_outputs(9625) <= a and not b;
    layer3_outputs(9626) <= not a or b;
    layer3_outputs(9627) <= a;
    layer3_outputs(9628) <= not b;
    layer3_outputs(9629) <= b;
    layer3_outputs(9630) <= not (a xor b);
    layer3_outputs(9631) <= not (a or b);
    layer3_outputs(9632) <= b;
    layer3_outputs(9633) <= not b;
    layer3_outputs(9634) <= a or b;
    layer3_outputs(9635) <= a xor b;
    layer3_outputs(9636) <= not a;
    layer3_outputs(9637) <= a xor b;
    layer3_outputs(9638) <= not b or a;
    layer3_outputs(9639) <= not a;
    layer3_outputs(9640) <= not (a xor b);
    layer3_outputs(9641) <= a;
    layer3_outputs(9642) <= a and b;
    layer3_outputs(9643) <= a and b;
    layer3_outputs(9644) <= a and not b;
    layer3_outputs(9645) <= a or b;
    layer3_outputs(9646) <= a or b;
    layer3_outputs(9647) <= not a;
    layer3_outputs(9648) <= not b;
    layer3_outputs(9649) <= not a;
    layer3_outputs(9650) <= a and b;
    layer3_outputs(9651) <= not b;
    layer3_outputs(9652) <= b;
    layer3_outputs(9653) <= a xor b;
    layer3_outputs(9654) <= b;
    layer3_outputs(9655) <= a and b;
    layer3_outputs(9656) <= not a or b;
    layer3_outputs(9657) <= not b;
    layer3_outputs(9658) <= a;
    layer3_outputs(9659) <= b;
    layer3_outputs(9660) <= not (a and b);
    layer3_outputs(9661) <= not a;
    layer3_outputs(9662) <= a;
    layer3_outputs(9663) <= a and not b;
    layer3_outputs(9664) <= a;
    layer3_outputs(9665) <= not (a or b);
    layer3_outputs(9666) <= b;
    layer3_outputs(9667) <= not (a and b);
    layer3_outputs(9668) <= a xor b;
    layer3_outputs(9669) <= 1'b1;
    layer3_outputs(9670) <= a and b;
    layer3_outputs(9671) <= a and b;
    layer3_outputs(9672) <= a xor b;
    layer3_outputs(9673) <= not a;
    layer3_outputs(9674) <= a and not b;
    layer3_outputs(9675) <= a;
    layer3_outputs(9676) <= a;
    layer3_outputs(9677) <= not b or a;
    layer3_outputs(9678) <= a;
    layer3_outputs(9679) <= not b;
    layer3_outputs(9680) <= not b;
    layer3_outputs(9681) <= not b or a;
    layer3_outputs(9682) <= not b;
    layer3_outputs(9683) <= not b;
    layer3_outputs(9684) <= a and not b;
    layer3_outputs(9685) <= 1'b1;
    layer3_outputs(9686) <= not (a and b);
    layer3_outputs(9687) <= b;
    layer3_outputs(9688) <= a and b;
    layer3_outputs(9689) <= not (a xor b);
    layer3_outputs(9690) <= a;
    layer3_outputs(9691) <= not (a and b);
    layer3_outputs(9692) <= not b;
    layer3_outputs(9693) <= not a;
    layer3_outputs(9694) <= a;
    layer3_outputs(9695) <= 1'b0;
    layer3_outputs(9696) <= not (a and b);
    layer3_outputs(9697) <= a;
    layer3_outputs(9698) <= a and b;
    layer3_outputs(9699) <= a xor b;
    layer3_outputs(9700) <= b;
    layer3_outputs(9701) <= not a;
    layer3_outputs(9702) <= not b;
    layer3_outputs(9703) <= not a or b;
    layer3_outputs(9704) <= not b;
    layer3_outputs(9705) <= not (a xor b);
    layer3_outputs(9706) <= not (a xor b);
    layer3_outputs(9707) <= a xor b;
    layer3_outputs(9708) <= b and not a;
    layer3_outputs(9709) <= not b;
    layer3_outputs(9710) <= not b or a;
    layer3_outputs(9711) <= a and b;
    layer3_outputs(9712) <= b;
    layer3_outputs(9713) <= a xor b;
    layer3_outputs(9714) <= b;
    layer3_outputs(9715) <= a and not b;
    layer3_outputs(9716) <= not b or a;
    layer3_outputs(9717) <= not (a xor b);
    layer3_outputs(9718) <= not (a xor b);
    layer3_outputs(9719) <= b and not a;
    layer3_outputs(9720) <= not b or a;
    layer3_outputs(9721) <= a;
    layer3_outputs(9722) <= a or b;
    layer3_outputs(9723) <= a and b;
    layer3_outputs(9724) <= not (a xor b);
    layer3_outputs(9725) <= not b;
    layer3_outputs(9726) <= a and b;
    layer3_outputs(9727) <= a and b;
    layer3_outputs(9728) <= not b;
    layer3_outputs(9729) <= a and b;
    layer3_outputs(9730) <= not a;
    layer3_outputs(9731) <= a;
    layer3_outputs(9732) <= not (a xor b);
    layer3_outputs(9733) <= a xor b;
    layer3_outputs(9734) <= a and not b;
    layer3_outputs(9735) <= a or b;
    layer3_outputs(9736) <= not (a and b);
    layer3_outputs(9737) <= a or b;
    layer3_outputs(9738) <= not a;
    layer3_outputs(9739) <= not b or a;
    layer3_outputs(9740) <= not (a xor b);
    layer3_outputs(9741) <= not a;
    layer3_outputs(9742) <= not (a and b);
    layer3_outputs(9743) <= 1'b1;
    layer3_outputs(9744) <= b and not a;
    layer3_outputs(9745) <= b and not a;
    layer3_outputs(9746) <= not (a and b);
    layer3_outputs(9747) <= a or b;
    layer3_outputs(9748) <= not b or a;
    layer3_outputs(9749) <= b;
    layer3_outputs(9750) <= not b;
    layer3_outputs(9751) <= not (a and b);
    layer3_outputs(9752) <= not b;
    layer3_outputs(9753) <= a xor b;
    layer3_outputs(9754) <= not (a xor b);
    layer3_outputs(9755) <= a;
    layer3_outputs(9756) <= b;
    layer3_outputs(9757) <= 1'b0;
    layer3_outputs(9758) <= not a;
    layer3_outputs(9759) <= b;
    layer3_outputs(9760) <= not b;
    layer3_outputs(9761) <= a and b;
    layer3_outputs(9762) <= a and not b;
    layer3_outputs(9763) <= a;
    layer3_outputs(9764) <= b and not a;
    layer3_outputs(9765) <= a and not b;
    layer3_outputs(9766) <= a;
    layer3_outputs(9767) <= not b;
    layer3_outputs(9768) <= not (a or b);
    layer3_outputs(9769) <= a and b;
    layer3_outputs(9770) <= not a;
    layer3_outputs(9771) <= not (a or b);
    layer3_outputs(9772) <= not b or a;
    layer3_outputs(9773) <= not a;
    layer3_outputs(9774) <= b;
    layer3_outputs(9775) <= not b;
    layer3_outputs(9776) <= not b;
    layer3_outputs(9777) <= not a or b;
    layer3_outputs(9778) <= not b;
    layer3_outputs(9779) <= a or b;
    layer3_outputs(9780) <= not b;
    layer3_outputs(9781) <= not b;
    layer3_outputs(9782) <= a;
    layer3_outputs(9783) <= a and not b;
    layer3_outputs(9784) <= a and b;
    layer3_outputs(9785) <= not (a xor b);
    layer3_outputs(9786) <= not (a or b);
    layer3_outputs(9787) <= not b;
    layer3_outputs(9788) <= a and b;
    layer3_outputs(9789) <= a;
    layer3_outputs(9790) <= b;
    layer3_outputs(9791) <= not b or a;
    layer3_outputs(9792) <= b;
    layer3_outputs(9793) <= a xor b;
    layer3_outputs(9794) <= a and b;
    layer3_outputs(9795) <= not (a and b);
    layer3_outputs(9796) <= a xor b;
    layer3_outputs(9797) <= a xor b;
    layer3_outputs(9798) <= not (a or b);
    layer3_outputs(9799) <= not b or a;
    layer3_outputs(9800) <= a xor b;
    layer3_outputs(9801) <= not b;
    layer3_outputs(9802) <= b;
    layer3_outputs(9803) <= not b;
    layer3_outputs(9804) <= b and not a;
    layer3_outputs(9805) <= not a or b;
    layer3_outputs(9806) <= not b;
    layer3_outputs(9807) <= b;
    layer3_outputs(9808) <= a or b;
    layer3_outputs(9809) <= not (a or b);
    layer3_outputs(9810) <= a;
    layer3_outputs(9811) <= not b or a;
    layer3_outputs(9812) <= not a;
    layer3_outputs(9813) <= a and b;
    layer3_outputs(9814) <= b;
    layer3_outputs(9815) <= b;
    layer3_outputs(9816) <= a and not b;
    layer3_outputs(9817) <= a and not b;
    layer3_outputs(9818) <= a;
    layer3_outputs(9819) <= b;
    layer3_outputs(9820) <= a xor b;
    layer3_outputs(9821) <= not a or b;
    layer3_outputs(9822) <= not (a and b);
    layer3_outputs(9823) <= a xor b;
    layer3_outputs(9824) <= a or b;
    layer3_outputs(9825) <= not b;
    layer3_outputs(9826) <= b and not a;
    layer3_outputs(9827) <= not b or a;
    layer3_outputs(9828) <= not (a or b);
    layer3_outputs(9829) <= b and not a;
    layer3_outputs(9830) <= a and b;
    layer3_outputs(9831) <= a xor b;
    layer3_outputs(9832) <= b;
    layer3_outputs(9833) <= b;
    layer3_outputs(9834) <= not a;
    layer3_outputs(9835) <= a or b;
    layer3_outputs(9836) <= not b;
    layer3_outputs(9837) <= not b;
    layer3_outputs(9838) <= not (a or b);
    layer3_outputs(9839) <= a;
    layer3_outputs(9840) <= b;
    layer3_outputs(9841) <= a or b;
    layer3_outputs(9842) <= not b or a;
    layer3_outputs(9843) <= b and not a;
    layer3_outputs(9844) <= b;
    layer3_outputs(9845) <= a;
    layer3_outputs(9846) <= a and b;
    layer3_outputs(9847) <= not (a or b);
    layer3_outputs(9848) <= not a;
    layer3_outputs(9849) <= a;
    layer3_outputs(9850) <= a and not b;
    layer3_outputs(9851) <= a and not b;
    layer3_outputs(9852) <= not (a and b);
    layer3_outputs(9853) <= a and not b;
    layer3_outputs(9854) <= not (a and b);
    layer3_outputs(9855) <= a and b;
    layer3_outputs(9856) <= not b;
    layer3_outputs(9857) <= not (a xor b);
    layer3_outputs(9858) <= a;
    layer3_outputs(9859) <= not (a and b);
    layer3_outputs(9860) <= b and not a;
    layer3_outputs(9861) <= not a or b;
    layer3_outputs(9862) <= a;
    layer3_outputs(9863) <= a;
    layer3_outputs(9864) <= not b;
    layer3_outputs(9865) <= a;
    layer3_outputs(9866) <= a and not b;
    layer3_outputs(9867) <= not a or b;
    layer3_outputs(9868) <= not b or a;
    layer3_outputs(9869) <= a and not b;
    layer3_outputs(9870) <= not a;
    layer3_outputs(9871) <= not a;
    layer3_outputs(9872) <= b;
    layer3_outputs(9873) <= a and b;
    layer3_outputs(9874) <= a and b;
    layer3_outputs(9875) <= not (a xor b);
    layer3_outputs(9876) <= a;
    layer3_outputs(9877) <= a xor b;
    layer3_outputs(9878) <= a and not b;
    layer3_outputs(9879) <= b;
    layer3_outputs(9880) <= not b;
    layer3_outputs(9881) <= not b or a;
    layer3_outputs(9882) <= a and b;
    layer3_outputs(9883) <= not (a and b);
    layer3_outputs(9884) <= not b or a;
    layer3_outputs(9885) <= a or b;
    layer3_outputs(9886) <= a;
    layer3_outputs(9887) <= a;
    layer3_outputs(9888) <= not b;
    layer3_outputs(9889) <= b;
    layer3_outputs(9890) <= not b;
    layer3_outputs(9891) <= not a or b;
    layer3_outputs(9892) <= b and not a;
    layer3_outputs(9893) <= not b or a;
    layer3_outputs(9894) <= a or b;
    layer3_outputs(9895) <= not b;
    layer3_outputs(9896) <= a xor b;
    layer3_outputs(9897) <= a and b;
    layer3_outputs(9898) <= not a;
    layer3_outputs(9899) <= a xor b;
    layer3_outputs(9900) <= not b or a;
    layer3_outputs(9901) <= not b or a;
    layer3_outputs(9902) <= b;
    layer3_outputs(9903) <= not (a and b);
    layer3_outputs(9904) <= not a;
    layer3_outputs(9905) <= a xor b;
    layer3_outputs(9906) <= a;
    layer3_outputs(9907) <= not b;
    layer3_outputs(9908) <= a or b;
    layer3_outputs(9909) <= b;
    layer3_outputs(9910) <= 1'b1;
    layer3_outputs(9911) <= not b;
    layer3_outputs(9912) <= a xor b;
    layer3_outputs(9913) <= a or b;
    layer3_outputs(9914) <= a and not b;
    layer3_outputs(9915) <= not b or a;
    layer3_outputs(9916) <= a xor b;
    layer3_outputs(9917) <= a;
    layer3_outputs(9918) <= 1'b0;
    layer3_outputs(9919) <= not b;
    layer3_outputs(9920) <= 1'b0;
    layer3_outputs(9921) <= not a;
    layer3_outputs(9922) <= not (a xor b);
    layer3_outputs(9923) <= a;
    layer3_outputs(9924) <= a or b;
    layer3_outputs(9925) <= a and b;
    layer3_outputs(9926) <= not a or b;
    layer3_outputs(9927) <= not (a and b);
    layer3_outputs(9928) <= not a or b;
    layer3_outputs(9929) <= not b;
    layer3_outputs(9930) <= a and b;
    layer3_outputs(9931) <= not a;
    layer3_outputs(9932) <= a;
    layer3_outputs(9933) <= a;
    layer3_outputs(9934) <= not b or a;
    layer3_outputs(9935) <= a xor b;
    layer3_outputs(9936) <= not a;
    layer3_outputs(9937) <= b and not a;
    layer3_outputs(9938) <= a xor b;
    layer3_outputs(9939) <= b and not a;
    layer3_outputs(9940) <= a and not b;
    layer3_outputs(9941) <= a;
    layer3_outputs(9942) <= a xor b;
    layer3_outputs(9943) <= not a;
    layer3_outputs(9944) <= not a or b;
    layer3_outputs(9945) <= a or b;
    layer3_outputs(9946) <= not b;
    layer3_outputs(9947) <= a;
    layer3_outputs(9948) <= not b;
    layer3_outputs(9949) <= b and not a;
    layer3_outputs(9950) <= not (a xor b);
    layer3_outputs(9951) <= a;
    layer3_outputs(9952) <= not (a and b);
    layer3_outputs(9953) <= not (a xor b);
    layer3_outputs(9954) <= a and not b;
    layer3_outputs(9955) <= not (a xor b);
    layer3_outputs(9956) <= a xor b;
    layer3_outputs(9957) <= not a;
    layer3_outputs(9958) <= not a;
    layer3_outputs(9959) <= not a;
    layer3_outputs(9960) <= b and not a;
    layer3_outputs(9961) <= not (a or b);
    layer3_outputs(9962) <= not b or a;
    layer3_outputs(9963) <= a and not b;
    layer3_outputs(9964) <= a or b;
    layer3_outputs(9965) <= not a or b;
    layer3_outputs(9966) <= a or b;
    layer3_outputs(9967) <= a or b;
    layer3_outputs(9968) <= not a or b;
    layer3_outputs(9969) <= not a or b;
    layer3_outputs(9970) <= 1'b0;
    layer3_outputs(9971) <= not a or b;
    layer3_outputs(9972) <= a and b;
    layer3_outputs(9973) <= not a;
    layer3_outputs(9974) <= not a;
    layer3_outputs(9975) <= a;
    layer3_outputs(9976) <= a;
    layer3_outputs(9977) <= not b or a;
    layer3_outputs(9978) <= a and b;
    layer3_outputs(9979) <= not (a and b);
    layer3_outputs(9980) <= not b;
    layer3_outputs(9981) <= not a or b;
    layer3_outputs(9982) <= not b;
    layer3_outputs(9983) <= not (a and b);
    layer3_outputs(9984) <= b and not a;
    layer3_outputs(9985) <= not a;
    layer3_outputs(9986) <= a and b;
    layer3_outputs(9987) <= not (a xor b);
    layer3_outputs(9988) <= b;
    layer3_outputs(9989) <= a xor b;
    layer3_outputs(9990) <= not a or b;
    layer3_outputs(9991) <= b and not a;
    layer3_outputs(9992) <= 1'b1;
    layer3_outputs(9993) <= not (a and b);
    layer3_outputs(9994) <= not a;
    layer3_outputs(9995) <= not (a and b);
    layer3_outputs(9996) <= not b;
    layer3_outputs(9997) <= not (a xor b);
    layer3_outputs(9998) <= a;
    layer3_outputs(9999) <= b;
    layer3_outputs(10000) <= not (a xor b);
    layer3_outputs(10001) <= not b or a;
    layer3_outputs(10002) <= not b;
    layer3_outputs(10003) <= a;
    layer3_outputs(10004) <= b and not a;
    layer3_outputs(10005) <= not (a and b);
    layer3_outputs(10006) <= not a;
    layer3_outputs(10007) <= a and not b;
    layer3_outputs(10008) <= not a;
    layer3_outputs(10009) <= not (a xor b);
    layer3_outputs(10010) <= b and not a;
    layer3_outputs(10011) <= not b;
    layer3_outputs(10012) <= not a or b;
    layer3_outputs(10013) <= not b;
    layer3_outputs(10014) <= b;
    layer3_outputs(10015) <= not a;
    layer3_outputs(10016) <= b;
    layer3_outputs(10017) <= a and b;
    layer3_outputs(10018) <= a;
    layer3_outputs(10019) <= not (a and b);
    layer3_outputs(10020) <= 1'b0;
    layer3_outputs(10021) <= a or b;
    layer3_outputs(10022) <= not (a or b);
    layer3_outputs(10023) <= b;
    layer3_outputs(10024) <= b and not a;
    layer3_outputs(10025) <= a or b;
    layer3_outputs(10026) <= a and not b;
    layer3_outputs(10027) <= not (a and b);
    layer3_outputs(10028) <= not b;
    layer3_outputs(10029) <= a and b;
    layer3_outputs(10030) <= not (a xor b);
    layer3_outputs(10031) <= a;
    layer3_outputs(10032) <= b and not a;
    layer3_outputs(10033) <= b;
    layer3_outputs(10034) <= a or b;
    layer3_outputs(10035) <= not b or a;
    layer3_outputs(10036) <= a or b;
    layer3_outputs(10037) <= not b;
    layer3_outputs(10038) <= not b or a;
    layer3_outputs(10039) <= not b;
    layer3_outputs(10040) <= not a;
    layer3_outputs(10041) <= not a;
    layer3_outputs(10042) <= not (a or b);
    layer3_outputs(10043) <= a and b;
    layer3_outputs(10044) <= not (a and b);
    layer3_outputs(10045) <= not (a and b);
    layer3_outputs(10046) <= not b;
    layer3_outputs(10047) <= not a or b;
    layer3_outputs(10048) <= a xor b;
    layer3_outputs(10049) <= 1'b0;
    layer3_outputs(10050) <= a xor b;
    layer3_outputs(10051) <= a and not b;
    layer3_outputs(10052) <= a and not b;
    layer3_outputs(10053) <= 1'b0;
    layer3_outputs(10054) <= b;
    layer3_outputs(10055) <= b;
    layer3_outputs(10056) <= a;
    layer3_outputs(10057) <= b and not a;
    layer3_outputs(10058) <= not a;
    layer3_outputs(10059) <= not (a or b);
    layer3_outputs(10060) <= not a;
    layer3_outputs(10061) <= not a or b;
    layer3_outputs(10062) <= b;
    layer3_outputs(10063) <= not (a xor b);
    layer3_outputs(10064) <= a and b;
    layer3_outputs(10065) <= not a;
    layer3_outputs(10066) <= not b;
    layer3_outputs(10067) <= not (a xor b);
    layer3_outputs(10068) <= b;
    layer3_outputs(10069) <= a and b;
    layer3_outputs(10070) <= b and not a;
    layer3_outputs(10071) <= a and b;
    layer3_outputs(10072) <= a or b;
    layer3_outputs(10073) <= not (a or b);
    layer3_outputs(10074) <= not a;
    layer3_outputs(10075) <= not b;
    layer3_outputs(10076) <= 1'b0;
    layer3_outputs(10077) <= a and not b;
    layer3_outputs(10078) <= not b;
    layer3_outputs(10079) <= not b or a;
    layer3_outputs(10080) <= not b or a;
    layer3_outputs(10081) <= a and not b;
    layer3_outputs(10082) <= b;
    layer3_outputs(10083) <= not a;
    layer3_outputs(10084) <= not (a and b);
    layer3_outputs(10085) <= b;
    layer3_outputs(10086) <= a and not b;
    layer3_outputs(10087) <= a xor b;
    layer3_outputs(10088) <= a xor b;
    layer3_outputs(10089) <= not (a and b);
    layer3_outputs(10090) <= a xor b;
    layer3_outputs(10091) <= b;
    layer3_outputs(10092) <= b;
    layer3_outputs(10093) <= not a or b;
    layer3_outputs(10094) <= not a;
    layer3_outputs(10095) <= not (a or b);
    layer3_outputs(10096) <= a xor b;
    layer3_outputs(10097) <= a xor b;
    layer3_outputs(10098) <= not a;
    layer3_outputs(10099) <= not a;
    layer3_outputs(10100) <= not b or a;
    layer3_outputs(10101) <= not a;
    layer3_outputs(10102) <= a and not b;
    layer3_outputs(10103) <= a;
    layer3_outputs(10104) <= a xor b;
    layer3_outputs(10105) <= not (a xor b);
    layer3_outputs(10106) <= 1'b0;
    layer3_outputs(10107) <= b and not a;
    layer3_outputs(10108) <= not b or a;
    layer3_outputs(10109) <= a xor b;
    layer3_outputs(10110) <= not (a xor b);
    layer3_outputs(10111) <= a and b;
    layer3_outputs(10112) <= a;
    layer3_outputs(10113) <= b and not a;
    layer3_outputs(10114) <= a or b;
    layer3_outputs(10115) <= not a;
    layer3_outputs(10116) <= not (a and b);
    layer3_outputs(10117) <= not b;
    layer3_outputs(10118) <= not (a and b);
    layer3_outputs(10119) <= not b;
    layer3_outputs(10120) <= b;
    layer3_outputs(10121) <= not a;
    layer3_outputs(10122) <= a and not b;
    layer3_outputs(10123) <= a;
    layer3_outputs(10124) <= not (a or b);
    layer3_outputs(10125) <= a;
    layer3_outputs(10126) <= b and not a;
    layer3_outputs(10127) <= not b or a;
    layer3_outputs(10128) <= not a or b;
    layer3_outputs(10129) <= a and b;
    layer3_outputs(10130) <= not (a or b);
    layer3_outputs(10131) <= 1'b0;
    layer3_outputs(10132) <= b and not a;
    layer3_outputs(10133) <= a;
    layer3_outputs(10134) <= a or b;
    layer3_outputs(10135) <= not a;
    layer3_outputs(10136) <= b;
    layer3_outputs(10137) <= not b or a;
    layer3_outputs(10138) <= not (a and b);
    layer3_outputs(10139) <= not (a xor b);
    layer3_outputs(10140) <= a and b;
    layer3_outputs(10141) <= a;
    layer3_outputs(10142) <= a and not b;
    layer3_outputs(10143) <= b and not a;
    layer3_outputs(10144) <= a xor b;
    layer3_outputs(10145) <= not (a and b);
    layer3_outputs(10146) <= not b;
    layer3_outputs(10147) <= not a;
    layer3_outputs(10148) <= a;
    layer3_outputs(10149) <= a or b;
    layer3_outputs(10150) <= not (a and b);
    layer3_outputs(10151) <= not a;
    layer3_outputs(10152) <= a and b;
    layer3_outputs(10153) <= not a;
    layer3_outputs(10154) <= b and not a;
    layer3_outputs(10155) <= a;
    layer3_outputs(10156) <= not b;
    layer3_outputs(10157) <= a;
    layer3_outputs(10158) <= not (a xor b);
    layer3_outputs(10159) <= a and b;
    layer3_outputs(10160) <= not a;
    layer3_outputs(10161) <= not a;
    layer3_outputs(10162) <= 1'b1;
    layer3_outputs(10163) <= not b or a;
    layer3_outputs(10164) <= not (a xor b);
    layer3_outputs(10165) <= not (a or b);
    layer3_outputs(10166) <= b;
    layer3_outputs(10167) <= a xor b;
    layer3_outputs(10168) <= not b;
    layer3_outputs(10169) <= a;
    layer3_outputs(10170) <= not (a and b);
    layer3_outputs(10171) <= not a or b;
    layer3_outputs(10172) <= not a or b;
    layer3_outputs(10173) <= not a;
    layer3_outputs(10174) <= b;
    layer3_outputs(10175) <= not a;
    layer3_outputs(10176) <= a;
    layer3_outputs(10177) <= not b or a;
    layer3_outputs(10178) <= b and not a;
    layer3_outputs(10179) <= a and b;
    layer3_outputs(10180) <= b;
    layer3_outputs(10181) <= a xor b;
    layer3_outputs(10182) <= a;
    layer3_outputs(10183) <= not (a or b);
    layer3_outputs(10184) <= not a;
    layer3_outputs(10185) <= not (a xor b);
    layer3_outputs(10186) <= not a;
    layer3_outputs(10187) <= a;
    layer3_outputs(10188) <= not a;
    layer3_outputs(10189) <= not b;
    layer3_outputs(10190) <= not b;
    layer3_outputs(10191) <= b;
    layer3_outputs(10192) <= a;
    layer3_outputs(10193) <= a and not b;
    layer3_outputs(10194) <= not a;
    layer3_outputs(10195) <= b;
    layer3_outputs(10196) <= not b;
    layer3_outputs(10197) <= b;
    layer3_outputs(10198) <= a xor b;
    layer3_outputs(10199) <= b and not a;
    layer3_outputs(10200) <= a or b;
    layer3_outputs(10201) <= a or b;
    layer3_outputs(10202) <= not a;
    layer3_outputs(10203) <= not (a or b);
    layer3_outputs(10204) <= a and not b;
    layer3_outputs(10205) <= not a;
    layer3_outputs(10206) <= not a or b;
    layer3_outputs(10207) <= b and not a;
    layer3_outputs(10208) <= not (a and b);
    layer3_outputs(10209) <= a;
    layer3_outputs(10210) <= 1'b1;
    layer3_outputs(10211) <= a and not b;
    layer3_outputs(10212) <= not (a or b);
    layer3_outputs(10213) <= 1'b1;
    layer3_outputs(10214) <= a or b;
    layer3_outputs(10215) <= not b;
    layer3_outputs(10216) <= a and not b;
    layer3_outputs(10217) <= b and not a;
    layer3_outputs(10218) <= not (a xor b);
    layer3_outputs(10219) <= a or b;
    layer3_outputs(10220) <= a or b;
    layer3_outputs(10221) <= a;
    layer3_outputs(10222) <= not a;
    layer3_outputs(10223) <= not a or b;
    layer3_outputs(10224) <= not b or a;
    layer3_outputs(10225) <= a xor b;
    layer3_outputs(10226) <= a and b;
    layer3_outputs(10227) <= a xor b;
    layer3_outputs(10228) <= a;
    layer3_outputs(10229) <= a;
    layer3_outputs(10230) <= a or b;
    layer3_outputs(10231) <= a;
    layer3_outputs(10232) <= a;
    layer3_outputs(10233) <= not b;
    layer3_outputs(10234) <= b and not a;
    layer3_outputs(10235) <= not b;
    layer3_outputs(10236) <= a and not b;
    layer3_outputs(10237) <= not a;
    layer3_outputs(10238) <= a and b;
    layer3_outputs(10239) <= a;
    layer4_outputs(0) <= b;
    layer4_outputs(1) <= a;
    layer4_outputs(2) <= not b;
    layer4_outputs(3) <= a xor b;
    layer4_outputs(4) <= not a;
    layer4_outputs(5) <= b;
    layer4_outputs(6) <= a;
    layer4_outputs(7) <= b;
    layer4_outputs(8) <= not b;
    layer4_outputs(9) <= b;
    layer4_outputs(10) <= a xor b;
    layer4_outputs(11) <= not a or b;
    layer4_outputs(12) <= not a;
    layer4_outputs(13) <= not b;
    layer4_outputs(14) <= not b;
    layer4_outputs(15) <= not a or b;
    layer4_outputs(16) <= not (a or b);
    layer4_outputs(17) <= a;
    layer4_outputs(18) <= a or b;
    layer4_outputs(19) <= b;
    layer4_outputs(20) <= a and b;
    layer4_outputs(21) <= a;
    layer4_outputs(22) <= not (a xor b);
    layer4_outputs(23) <= not a;
    layer4_outputs(24) <= a;
    layer4_outputs(25) <= not b;
    layer4_outputs(26) <= not b;
    layer4_outputs(27) <= a;
    layer4_outputs(28) <= not (a and b);
    layer4_outputs(29) <= b;
    layer4_outputs(30) <= not b or a;
    layer4_outputs(31) <= not b;
    layer4_outputs(32) <= b;
    layer4_outputs(33) <= not b or a;
    layer4_outputs(34) <= not b;
    layer4_outputs(35) <= not a;
    layer4_outputs(36) <= not (a xor b);
    layer4_outputs(37) <= not a;
    layer4_outputs(38) <= b;
    layer4_outputs(39) <= not (a and b);
    layer4_outputs(40) <= not (a xor b);
    layer4_outputs(41) <= a;
    layer4_outputs(42) <= not a or b;
    layer4_outputs(43) <= a xor b;
    layer4_outputs(44) <= not a;
    layer4_outputs(45) <= not b or a;
    layer4_outputs(46) <= a;
    layer4_outputs(47) <= a;
    layer4_outputs(48) <= a and not b;
    layer4_outputs(49) <= not (a xor b);
    layer4_outputs(50) <= a or b;
    layer4_outputs(51) <= not (a xor b);
    layer4_outputs(52) <= not b;
    layer4_outputs(53) <= not b;
    layer4_outputs(54) <= not (a xor b);
    layer4_outputs(55) <= a and not b;
    layer4_outputs(56) <= b;
    layer4_outputs(57) <= a xor b;
    layer4_outputs(58) <= a xor b;
    layer4_outputs(59) <= not (a or b);
    layer4_outputs(60) <= a and not b;
    layer4_outputs(61) <= not a;
    layer4_outputs(62) <= a xor b;
    layer4_outputs(63) <= a;
    layer4_outputs(64) <= not a;
    layer4_outputs(65) <= not b;
    layer4_outputs(66) <= not b;
    layer4_outputs(67) <= a xor b;
    layer4_outputs(68) <= a;
    layer4_outputs(69) <= b;
    layer4_outputs(70) <= not (a or b);
    layer4_outputs(71) <= not b or a;
    layer4_outputs(72) <= not b;
    layer4_outputs(73) <= a;
    layer4_outputs(74) <= not (a xor b);
    layer4_outputs(75) <= not (a xor b);
    layer4_outputs(76) <= not a;
    layer4_outputs(77) <= not (a and b);
    layer4_outputs(78) <= not a;
    layer4_outputs(79) <= b;
    layer4_outputs(80) <= not (a or b);
    layer4_outputs(81) <= a xor b;
    layer4_outputs(82) <= not (a and b);
    layer4_outputs(83) <= a;
    layer4_outputs(84) <= a;
    layer4_outputs(85) <= not b;
    layer4_outputs(86) <= not b or a;
    layer4_outputs(87) <= not (a xor b);
    layer4_outputs(88) <= not a;
    layer4_outputs(89) <= not (a xor b);
    layer4_outputs(90) <= a and b;
    layer4_outputs(91) <= not b;
    layer4_outputs(92) <= not (a or b);
    layer4_outputs(93) <= a;
    layer4_outputs(94) <= not b;
    layer4_outputs(95) <= not b;
    layer4_outputs(96) <= b;
    layer4_outputs(97) <= a and b;
    layer4_outputs(98) <= not b;
    layer4_outputs(99) <= a and not b;
    layer4_outputs(100) <= b and not a;
    layer4_outputs(101) <= not (a and b);
    layer4_outputs(102) <= not b;
    layer4_outputs(103) <= not b;
    layer4_outputs(104) <= not (a xor b);
    layer4_outputs(105) <= not (a xor b);
    layer4_outputs(106) <= not a;
    layer4_outputs(107) <= a or b;
    layer4_outputs(108) <= not b;
    layer4_outputs(109) <= b;
    layer4_outputs(110) <= a and not b;
    layer4_outputs(111) <= not b;
    layer4_outputs(112) <= not b;
    layer4_outputs(113) <= not (a and b);
    layer4_outputs(114) <= a;
    layer4_outputs(115) <= not a;
    layer4_outputs(116) <= a;
    layer4_outputs(117) <= a;
    layer4_outputs(118) <= not b;
    layer4_outputs(119) <= not b;
    layer4_outputs(120) <= b;
    layer4_outputs(121) <= a xor b;
    layer4_outputs(122) <= b and not a;
    layer4_outputs(123) <= a or b;
    layer4_outputs(124) <= a or b;
    layer4_outputs(125) <= not a or b;
    layer4_outputs(126) <= b;
    layer4_outputs(127) <= a xor b;
    layer4_outputs(128) <= a;
    layer4_outputs(129) <= a and b;
    layer4_outputs(130) <= a and b;
    layer4_outputs(131) <= b;
    layer4_outputs(132) <= a;
    layer4_outputs(133) <= not b;
    layer4_outputs(134) <= not (a xor b);
    layer4_outputs(135) <= a;
    layer4_outputs(136) <= b and not a;
    layer4_outputs(137) <= b;
    layer4_outputs(138) <= b and not a;
    layer4_outputs(139) <= b;
    layer4_outputs(140) <= a and not b;
    layer4_outputs(141) <= not (a and b);
    layer4_outputs(142) <= not (a and b);
    layer4_outputs(143) <= not (a or b);
    layer4_outputs(144) <= b;
    layer4_outputs(145) <= a;
    layer4_outputs(146) <= a;
    layer4_outputs(147) <= a and b;
    layer4_outputs(148) <= b and not a;
    layer4_outputs(149) <= not b;
    layer4_outputs(150) <= a and b;
    layer4_outputs(151) <= not a;
    layer4_outputs(152) <= not (a and b);
    layer4_outputs(153) <= not (a xor b);
    layer4_outputs(154) <= not (a or b);
    layer4_outputs(155) <= a and not b;
    layer4_outputs(156) <= b;
    layer4_outputs(157) <= not (a and b);
    layer4_outputs(158) <= b and not a;
    layer4_outputs(159) <= not (a xor b);
    layer4_outputs(160) <= a;
    layer4_outputs(161) <= not a or b;
    layer4_outputs(162) <= a xor b;
    layer4_outputs(163) <= not b;
    layer4_outputs(164) <= not b;
    layer4_outputs(165) <= not b;
    layer4_outputs(166) <= not a;
    layer4_outputs(167) <= a or b;
    layer4_outputs(168) <= not b;
    layer4_outputs(169) <= a and b;
    layer4_outputs(170) <= not (a and b);
    layer4_outputs(171) <= not a or b;
    layer4_outputs(172) <= a;
    layer4_outputs(173) <= a or b;
    layer4_outputs(174) <= a xor b;
    layer4_outputs(175) <= a;
    layer4_outputs(176) <= not (a and b);
    layer4_outputs(177) <= b and not a;
    layer4_outputs(178) <= not b;
    layer4_outputs(179) <= a xor b;
    layer4_outputs(180) <= b;
    layer4_outputs(181) <= a and not b;
    layer4_outputs(182) <= a;
    layer4_outputs(183) <= b and not a;
    layer4_outputs(184) <= not (a or b);
    layer4_outputs(185) <= not (a xor b);
    layer4_outputs(186) <= a xor b;
    layer4_outputs(187) <= b;
    layer4_outputs(188) <= b;
    layer4_outputs(189) <= not b;
    layer4_outputs(190) <= b and not a;
    layer4_outputs(191) <= not a;
    layer4_outputs(192) <= a and not b;
    layer4_outputs(193) <= not (a xor b);
    layer4_outputs(194) <= not (a or b);
    layer4_outputs(195) <= not (a xor b);
    layer4_outputs(196) <= a or b;
    layer4_outputs(197) <= not b;
    layer4_outputs(198) <= 1'b1;
    layer4_outputs(199) <= not b;
    layer4_outputs(200) <= not (a xor b);
    layer4_outputs(201) <= not b;
    layer4_outputs(202) <= not b;
    layer4_outputs(203) <= not a;
    layer4_outputs(204) <= not b;
    layer4_outputs(205) <= a xor b;
    layer4_outputs(206) <= a and b;
    layer4_outputs(207) <= b;
    layer4_outputs(208) <= b;
    layer4_outputs(209) <= not a;
    layer4_outputs(210) <= not a or b;
    layer4_outputs(211) <= a xor b;
    layer4_outputs(212) <= not b or a;
    layer4_outputs(213) <= not b;
    layer4_outputs(214) <= not (a or b);
    layer4_outputs(215) <= a;
    layer4_outputs(216) <= a;
    layer4_outputs(217) <= not a;
    layer4_outputs(218) <= a;
    layer4_outputs(219) <= a xor b;
    layer4_outputs(220) <= not (a xor b);
    layer4_outputs(221) <= not b;
    layer4_outputs(222) <= not a;
    layer4_outputs(223) <= a;
    layer4_outputs(224) <= not a;
    layer4_outputs(225) <= not b;
    layer4_outputs(226) <= not (a xor b);
    layer4_outputs(227) <= a;
    layer4_outputs(228) <= not b;
    layer4_outputs(229) <= not (a xor b);
    layer4_outputs(230) <= 1'b0;
    layer4_outputs(231) <= a xor b;
    layer4_outputs(232) <= not (a and b);
    layer4_outputs(233) <= a;
    layer4_outputs(234) <= not (a or b);
    layer4_outputs(235) <= b;
    layer4_outputs(236) <= a;
    layer4_outputs(237) <= not a;
    layer4_outputs(238) <= not (a and b);
    layer4_outputs(239) <= b;
    layer4_outputs(240) <= not b or a;
    layer4_outputs(241) <= a xor b;
    layer4_outputs(242) <= not a or b;
    layer4_outputs(243) <= b and not a;
    layer4_outputs(244) <= not (a and b);
    layer4_outputs(245) <= not a;
    layer4_outputs(246) <= b;
    layer4_outputs(247) <= not a or b;
    layer4_outputs(248) <= not a or b;
    layer4_outputs(249) <= a and b;
    layer4_outputs(250) <= not b;
    layer4_outputs(251) <= a;
    layer4_outputs(252) <= 1'b0;
    layer4_outputs(253) <= not b;
    layer4_outputs(254) <= not (a or b);
    layer4_outputs(255) <= a;
    layer4_outputs(256) <= not a;
    layer4_outputs(257) <= a;
    layer4_outputs(258) <= not b;
    layer4_outputs(259) <= a and b;
    layer4_outputs(260) <= not b;
    layer4_outputs(261) <= not b;
    layer4_outputs(262) <= not b;
    layer4_outputs(263) <= not (a xor b);
    layer4_outputs(264) <= a;
    layer4_outputs(265) <= a xor b;
    layer4_outputs(266) <= b;
    layer4_outputs(267) <= not (a xor b);
    layer4_outputs(268) <= a;
    layer4_outputs(269) <= a;
    layer4_outputs(270) <= a and not b;
    layer4_outputs(271) <= b;
    layer4_outputs(272) <= b;
    layer4_outputs(273) <= not (a or b);
    layer4_outputs(274) <= not (a or b);
    layer4_outputs(275) <= a;
    layer4_outputs(276) <= not (a and b);
    layer4_outputs(277) <= not (a or b);
    layer4_outputs(278) <= not a;
    layer4_outputs(279) <= b and not a;
    layer4_outputs(280) <= a and not b;
    layer4_outputs(281) <= b;
    layer4_outputs(282) <= a and not b;
    layer4_outputs(283) <= a and b;
    layer4_outputs(284) <= not (a and b);
    layer4_outputs(285) <= a and not b;
    layer4_outputs(286) <= not b;
    layer4_outputs(287) <= a;
    layer4_outputs(288) <= b and not a;
    layer4_outputs(289) <= not a or b;
    layer4_outputs(290) <= not (a and b);
    layer4_outputs(291) <= not a or b;
    layer4_outputs(292) <= not (a and b);
    layer4_outputs(293) <= a and not b;
    layer4_outputs(294) <= not b;
    layer4_outputs(295) <= a and b;
    layer4_outputs(296) <= not b;
    layer4_outputs(297) <= not (a xor b);
    layer4_outputs(298) <= b;
    layer4_outputs(299) <= a;
    layer4_outputs(300) <= not b or a;
    layer4_outputs(301) <= not b;
    layer4_outputs(302) <= a and b;
    layer4_outputs(303) <= b;
    layer4_outputs(304) <= not (a xor b);
    layer4_outputs(305) <= not a or b;
    layer4_outputs(306) <= b and not a;
    layer4_outputs(307) <= b;
    layer4_outputs(308) <= a and b;
    layer4_outputs(309) <= a;
    layer4_outputs(310) <= a or b;
    layer4_outputs(311) <= a and b;
    layer4_outputs(312) <= a and b;
    layer4_outputs(313) <= a;
    layer4_outputs(314) <= not a;
    layer4_outputs(315) <= a or b;
    layer4_outputs(316) <= not (a xor b);
    layer4_outputs(317) <= not (a and b);
    layer4_outputs(318) <= not b;
    layer4_outputs(319) <= b;
    layer4_outputs(320) <= not b or a;
    layer4_outputs(321) <= not (a xor b);
    layer4_outputs(322) <= not a or b;
    layer4_outputs(323) <= b and not a;
    layer4_outputs(324) <= a;
    layer4_outputs(325) <= not b;
    layer4_outputs(326) <= not a or b;
    layer4_outputs(327) <= not a or b;
    layer4_outputs(328) <= a xor b;
    layer4_outputs(329) <= not (a or b);
    layer4_outputs(330) <= b;
    layer4_outputs(331) <= not (a or b);
    layer4_outputs(332) <= not b;
    layer4_outputs(333) <= b;
    layer4_outputs(334) <= not a;
    layer4_outputs(335) <= b;
    layer4_outputs(336) <= not (a xor b);
    layer4_outputs(337) <= a and b;
    layer4_outputs(338) <= b and not a;
    layer4_outputs(339) <= not b;
    layer4_outputs(340) <= not a;
    layer4_outputs(341) <= a;
    layer4_outputs(342) <= a and not b;
    layer4_outputs(343) <= not (a xor b);
    layer4_outputs(344) <= not a;
    layer4_outputs(345) <= not b or a;
    layer4_outputs(346) <= not (a xor b);
    layer4_outputs(347) <= not (a and b);
    layer4_outputs(348) <= not b or a;
    layer4_outputs(349) <= not a;
    layer4_outputs(350) <= a;
    layer4_outputs(351) <= not b;
    layer4_outputs(352) <= a or b;
    layer4_outputs(353) <= a or b;
    layer4_outputs(354) <= not (a xor b);
    layer4_outputs(355) <= not a;
    layer4_outputs(356) <= not (a xor b);
    layer4_outputs(357) <= a and not b;
    layer4_outputs(358) <= b;
    layer4_outputs(359) <= not b;
    layer4_outputs(360) <= b;
    layer4_outputs(361) <= not a;
    layer4_outputs(362) <= a;
    layer4_outputs(363) <= not a;
    layer4_outputs(364) <= 1'b1;
    layer4_outputs(365) <= a;
    layer4_outputs(366) <= a and not b;
    layer4_outputs(367) <= not a;
    layer4_outputs(368) <= not a or b;
    layer4_outputs(369) <= b and not a;
    layer4_outputs(370) <= a;
    layer4_outputs(371) <= a and not b;
    layer4_outputs(372) <= a and b;
    layer4_outputs(373) <= not a;
    layer4_outputs(374) <= not (a and b);
    layer4_outputs(375) <= a xor b;
    layer4_outputs(376) <= not (a xor b);
    layer4_outputs(377) <= a;
    layer4_outputs(378) <= b and not a;
    layer4_outputs(379) <= not a;
    layer4_outputs(380) <= not a;
    layer4_outputs(381) <= b and not a;
    layer4_outputs(382) <= not (a xor b);
    layer4_outputs(383) <= not (a and b);
    layer4_outputs(384) <= not b or a;
    layer4_outputs(385) <= not (a and b);
    layer4_outputs(386) <= a;
    layer4_outputs(387) <= a;
    layer4_outputs(388) <= not (a xor b);
    layer4_outputs(389) <= b;
    layer4_outputs(390) <= not b or a;
    layer4_outputs(391) <= not (a xor b);
    layer4_outputs(392) <= b and not a;
    layer4_outputs(393) <= a xor b;
    layer4_outputs(394) <= a and not b;
    layer4_outputs(395) <= a and b;
    layer4_outputs(396) <= b;
    layer4_outputs(397) <= not a;
    layer4_outputs(398) <= not a or b;
    layer4_outputs(399) <= not a or b;
    layer4_outputs(400) <= a;
    layer4_outputs(401) <= not a or b;
    layer4_outputs(402) <= not b;
    layer4_outputs(403) <= a and not b;
    layer4_outputs(404) <= not a or b;
    layer4_outputs(405) <= not a or b;
    layer4_outputs(406) <= not b;
    layer4_outputs(407) <= b and not a;
    layer4_outputs(408) <= 1'b1;
    layer4_outputs(409) <= a;
    layer4_outputs(410) <= a or b;
    layer4_outputs(411) <= not a or b;
    layer4_outputs(412) <= not b;
    layer4_outputs(413) <= not (a xor b);
    layer4_outputs(414) <= not a;
    layer4_outputs(415) <= b and not a;
    layer4_outputs(416) <= a or b;
    layer4_outputs(417) <= a xor b;
    layer4_outputs(418) <= not b;
    layer4_outputs(419) <= not b;
    layer4_outputs(420) <= a or b;
    layer4_outputs(421) <= not a;
    layer4_outputs(422) <= not a;
    layer4_outputs(423) <= not b or a;
    layer4_outputs(424) <= b;
    layer4_outputs(425) <= not a;
    layer4_outputs(426) <= a;
    layer4_outputs(427) <= a xor b;
    layer4_outputs(428) <= a xor b;
    layer4_outputs(429) <= b and not a;
    layer4_outputs(430) <= a;
    layer4_outputs(431) <= a;
    layer4_outputs(432) <= not b or a;
    layer4_outputs(433) <= not (a xor b);
    layer4_outputs(434) <= a;
    layer4_outputs(435) <= not (a xor b);
    layer4_outputs(436) <= not b;
    layer4_outputs(437) <= not a or b;
    layer4_outputs(438) <= a or b;
    layer4_outputs(439) <= not (a or b);
    layer4_outputs(440) <= b and not a;
    layer4_outputs(441) <= a and not b;
    layer4_outputs(442) <= a and b;
    layer4_outputs(443) <= a or b;
    layer4_outputs(444) <= not (a xor b);
    layer4_outputs(445) <= a;
    layer4_outputs(446) <= a or b;
    layer4_outputs(447) <= not (a and b);
    layer4_outputs(448) <= a xor b;
    layer4_outputs(449) <= not (a or b);
    layer4_outputs(450) <= not b;
    layer4_outputs(451) <= b and not a;
    layer4_outputs(452) <= b;
    layer4_outputs(453) <= not (a xor b);
    layer4_outputs(454) <= not (a or b);
    layer4_outputs(455) <= not b;
    layer4_outputs(456) <= b and not a;
    layer4_outputs(457) <= not (a or b);
    layer4_outputs(458) <= b and not a;
    layer4_outputs(459) <= not (a or b);
    layer4_outputs(460) <= a;
    layer4_outputs(461) <= b and not a;
    layer4_outputs(462) <= not b or a;
    layer4_outputs(463) <= a or b;
    layer4_outputs(464) <= not (a or b);
    layer4_outputs(465) <= not b;
    layer4_outputs(466) <= not a;
    layer4_outputs(467) <= a xor b;
    layer4_outputs(468) <= not (a or b);
    layer4_outputs(469) <= not a;
    layer4_outputs(470) <= not a;
    layer4_outputs(471) <= not b;
    layer4_outputs(472) <= not (a and b);
    layer4_outputs(473) <= not (a xor b);
    layer4_outputs(474) <= not (a xor b);
    layer4_outputs(475) <= not a;
    layer4_outputs(476) <= a and not b;
    layer4_outputs(477) <= not (a and b);
    layer4_outputs(478) <= a;
    layer4_outputs(479) <= b;
    layer4_outputs(480) <= not (a xor b);
    layer4_outputs(481) <= not a;
    layer4_outputs(482) <= a and b;
    layer4_outputs(483) <= not b or a;
    layer4_outputs(484) <= not b;
    layer4_outputs(485) <= not (a xor b);
    layer4_outputs(486) <= a;
    layer4_outputs(487) <= not a;
    layer4_outputs(488) <= not a;
    layer4_outputs(489) <= b;
    layer4_outputs(490) <= not (a xor b);
    layer4_outputs(491) <= b;
    layer4_outputs(492) <= b;
    layer4_outputs(493) <= not (a xor b);
    layer4_outputs(494) <= not a or b;
    layer4_outputs(495) <= a;
    layer4_outputs(496) <= a;
    layer4_outputs(497) <= not (a and b);
    layer4_outputs(498) <= not b;
    layer4_outputs(499) <= not a;
    layer4_outputs(500) <= b;
    layer4_outputs(501) <= a xor b;
    layer4_outputs(502) <= not b;
    layer4_outputs(503) <= not b or a;
    layer4_outputs(504) <= b;
    layer4_outputs(505) <= b;
    layer4_outputs(506) <= not a;
    layer4_outputs(507) <= b;
    layer4_outputs(508) <= b;
    layer4_outputs(509) <= not a or b;
    layer4_outputs(510) <= a;
    layer4_outputs(511) <= not b or a;
    layer4_outputs(512) <= not b;
    layer4_outputs(513) <= not b or a;
    layer4_outputs(514) <= not (a xor b);
    layer4_outputs(515) <= b and not a;
    layer4_outputs(516) <= 1'b1;
    layer4_outputs(517) <= b and not a;
    layer4_outputs(518) <= a and b;
    layer4_outputs(519) <= a and not b;
    layer4_outputs(520) <= not (a xor b);
    layer4_outputs(521) <= not (a xor b);
    layer4_outputs(522) <= a xor b;
    layer4_outputs(523) <= not (a and b);
    layer4_outputs(524) <= a;
    layer4_outputs(525) <= not (a or b);
    layer4_outputs(526) <= a or b;
    layer4_outputs(527) <= not (a or b);
    layer4_outputs(528) <= a or b;
    layer4_outputs(529) <= a and b;
    layer4_outputs(530) <= not b or a;
    layer4_outputs(531) <= not (a or b);
    layer4_outputs(532) <= a and not b;
    layer4_outputs(533) <= not b;
    layer4_outputs(534) <= a or b;
    layer4_outputs(535) <= a;
    layer4_outputs(536) <= not b;
    layer4_outputs(537) <= not b;
    layer4_outputs(538) <= not (a xor b);
    layer4_outputs(539) <= not (a xor b);
    layer4_outputs(540) <= not a;
    layer4_outputs(541) <= a;
    layer4_outputs(542) <= not (a xor b);
    layer4_outputs(543) <= b and not a;
    layer4_outputs(544) <= not a or b;
    layer4_outputs(545) <= a;
    layer4_outputs(546) <= not b or a;
    layer4_outputs(547) <= a;
    layer4_outputs(548) <= b;
    layer4_outputs(549) <= not b;
    layer4_outputs(550) <= not b or a;
    layer4_outputs(551) <= a;
    layer4_outputs(552) <= not a or b;
    layer4_outputs(553) <= 1'b0;
    layer4_outputs(554) <= a or b;
    layer4_outputs(555) <= not (a and b);
    layer4_outputs(556) <= a and not b;
    layer4_outputs(557) <= a xor b;
    layer4_outputs(558) <= not (a or b);
    layer4_outputs(559) <= not b;
    layer4_outputs(560) <= not b;
    layer4_outputs(561) <= a;
    layer4_outputs(562) <= not a;
    layer4_outputs(563) <= a;
    layer4_outputs(564) <= not a;
    layer4_outputs(565) <= b;
    layer4_outputs(566) <= b;
    layer4_outputs(567) <= not (a or b);
    layer4_outputs(568) <= not b;
    layer4_outputs(569) <= not a;
    layer4_outputs(570) <= not (a or b);
    layer4_outputs(571) <= a or b;
    layer4_outputs(572) <= a and not b;
    layer4_outputs(573) <= not b;
    layer4_outputs(574) <= not b or a;
    layer4_outputs(575) <= not a;
    layer4_outputs(576) <= a xor b;
    layer4_outputs(577) <= not a;
    layer4_outputs(578) <= not (a xor b);
    layer4_outputs(579) <= not (a and b);
    layer4_outputs(580) <= b;
    layer4_outputs(581) <= not b;
    layer4_outputs(582) <= not b or a;
    layer4_outputs(583) <= not b;
    layer4_outputs(584) <= a and not b;
    layer4_outputs(585) <= b;
    layer4_outputs(586) <= b;
    layer4_outputs(587) <= 1'b0;
    layer4_outputs(588) <= a;
    layer4_outputs(589) <= a xor b;
    layer4_outputs(590) <= not (a or b);
    layer4_outputs(591) <= b;
    layer4_outputs(592) <= a;
    layer4_outputs(593) <= not (a and b);
    layer4_outputs(594) <= a;
    layer4_outputs(595) <= a;
    layer4_outputs(596) <= not b;
    layer4_outputs(597) <= b;
    layer4_outputs(598) <= a xor b;
    layer4_outputs(599) <= not (a or b);
    layer4_outputs(600) <= not (a xor b);
    layer4_outputs(601) <= a and b;
    layer4_outputs(602) <= not b;
    layer4_outputs(603) <= a;
    layer4_outputs(604) <= not (a and b);
    layer4_outputs(605) <= not (a xor b);
    layer4_outputs(606) <= a and b;
    layer4_outputs(607) <= b and not a;
    layer4_outputs(608) <= b and not a;
    layer4_outputs(609) <= b;
    layer4_outputs(610) <= b;
    layer4_outputs(611) <= not b;
    layer4_outputs(612) <= not a or b;
    layer4_outputs(613) <= not (a or b);
    layer4_outputs(614) <= a;
    layer4_outputs(615) <= a xor b;
    layer4_outputs(616) <= a and b;
    layer4_outputs(617) <= not b;
    layer4_outputs(618) <= b;
    layer4_outputs(619) <= a;
    layer4_outputs(620) <= a;
    layer4_outputs(621) <= b and not a;
    layer4_outputs(622) <= a and not b;
    layer4_outputs(623) <= not a or b;
    layer4_outputs(624) <= not a;
    layer4_outputs(625) <= a or b;
    layer4_outputs(626) <= not a;
    layer4_outputs(627) <= a and b;
    layer4_outputs(628) <= b;
    layer4_outputs(629) <= not a;
    layer4_outputs(630) <= not b;
    layer4_outputs(631) <= b and not a;
    layer4_outputs(632) <= not a;
    layer4_outputs(633) <= a and b;
    layer4_outputs(634) <= not (a and b);
    layer4_outputs(635) <= a and b;
    layer4_outputs(636) <= a or b;
    layer4_outputs(637) <= a;
    layer4_outputs(638) <= a and not b;
    layer4_outputs(639) <= b;
    layer4_outputs(640) <= not a;
    layer4_outputs(641) <= not b;
    layer4_outputs(642) <= b;
    layer4_outputs(643) <= a and b;
    layer4_outputs(644) <= not (a or b);
    layer4_outputs(645) <= not b;
    layer4_outputs(646) <= b;
    layer4_outputs(647) <= not a;
    layer4_outputs(648) <= a and b;
    layer4_outputs(649) <= not b;
    layer4_outputs(650) <= b;
    layer4_outputs(651) <= not a;
    layer4_outputs(652) <= a and not b;
    layer4_outputs(653) <= not b;
    layer4_outputs(654) <= a xor b;
    layer4_outputs(655) <= a;
    layer4_outputs(656) <= b;
    layer4_outputs(657) <= a xor b;
    layer4_outputs(658) <= not (a and b);
    layer4_outputs(659) <= not (a xor b);
    layer4_outputs(660) <= not (a xor b);
    layer4_outputs(661) <= a xor b;
    layer4_outputs(662) <= not a or b;
    layer4_outputs(663) <= not (a or b);
    layer4_outputs(664) <= not (a xor b);
    layer4_outputs(665) <= not (a and b);
    layer4_outputs(666) <= a;
    layer4_outputs(667) <= not b;
    layer4_outputs(668) <= b and not a;
    layer4_outputs(669) <= b;
    layer4_outputs(670) <= 1'b0;
    layer4_outputs(671) <= a xor b;
    layer4_outputs(672) <= not (a or b);
    layer4_outputs(673) <= a;
    layer4_outputs(674) <= not a;
    layer4_outputs(675) <= not b;
    layer4_outputs(676) <= not (a xor b);
    layer4_outputs(677) <= not b;
    layer4_outputs(678) <= a or b;
    layer4_outputs(679) <= not b;
    layer4_outputs(680) <= not (a or b);
    layer4_outputs(681) <= b;
    layer4_outputs(682) <= not a or b;
    layer4_outputs(683) <= b and not a;
    layer4_outputs(684) <= a and b;
    layer4_outputs(685) <= not b;
    layer4_outputs(686) <= a;
    layer4_outputs(687) <= not b or a;
    layer4_outputs(688) <= not (a or b);
    layer4_outputs(689) <= a or b;
    layer4_outputs(690) <= a and not b;
    layer4_outputs(691) <= a and b;
    layer4_outputs(692) <= a;
    layer4_outputs(693) <= b;
    layer4_outputs(694) <= not a or b;
    layer4_outputs(695) <= not a;
    layer4_outputs(696) <= a xor b;
    layer4_outputs(697) <= not b or a;
    layer4_outputs(698) <= b;
    layer4_outputs(699) <= not (a or b);
    layer4_outputs(700) <= a;
    layer4_outputs(701) <= not (a xor b);
    layer4_outputs(702) <= a or b;
    layer4_outputs(703) <= not (a and b);
    layer4_outputs(704) <= not (a xor b);
    layer4_outputs(705) <= not b;
    layer4_outputs(706) <= a xor b;
    layer4_outputs(707) <= not b or a;
    layer4_outputs(708) <= b;
    layer4_outputs(709) <= not a or b;
    layer4_outputs(710) <= b;
    layer4_outputs(711) <= not b;
    layer4_outputs(712) <= a xor b;
    layer4_outputs(713) <= not a or b;
    layer4_outputs(714) <= not (a xor b);
    layer4_outputs(715) <= a;
    layer4_outputs(716) <= a xor b;
    layer4_outputs(717) <= not (a or b);
    layer4_outputs(718) <= not a or b;
    layer4_outputs(719) <= a or b;
    layer4_outputs(720) <= a xor b;
    layer4_outputs(721) <= b and not a;
    layer4_outputs(722) <= not (a xor b);
    layer4_outputs(723) <= b;
    layer4_outputs(724) <= not (a xor b);
    layer4_outputs(725) <= not (a and b);
    layer4_outputs(726) <= b;
    layer4_outputs(727) <= not b;
    layer4_outputs(728) <= not (a and b);
    layer4_outputs(729) <= not b;
    layer4_outputs(730) <= a and not b;
    layer4_outputs(731) <= a xor b;
    layer4_outputs(732) <= a and not b;
    layer4_outputs(733) <= not (a xor b);
    layer4_outputs(734) <= b;
    layer4_outputs(735) <= a xor b;
    layer4_outputs(736) <= a xor b;
    layer4_outputs(737) <= not a;
    layer4_outputs(738) <= b and not a;
    layer4_outputs(739) <= a and b;
    layer4_outputs(740) <= a xor b;
    layer4_outputs(741) <= a and not b;
    layer4_outputs(742) <= not b;
    layer4_outputs(743) <= not b;
    layer4_outputs(744) <= a and b;
    layer4_outputs(745) <= a and b;
    layer4_outputs(746) <= not (a xor b);
    layer4_outputs(747) <= not (a xor b);
    layer4_outputs(748) <= not b or a;
    layer4_outputs(749) <= b;
    layer4_outputs(750) <= a or b;
    layer4_outputs(751) <= b;
    layer4_outputs(752) <= not (a or b);
    layer4_outputs(753) <= not b;
    layer4_outputs(754) <= not (a and b);
    layer4_outputs(755) <= b;
    layer4_outputs(756) <= not (a or b);
    layer4_outputs(757) <= a;
    layer4_outputs(758) <= not b or a;
    layer4_outputs(759) <= b;
    layer4_outputs(760) <= a xor b;
    layer4_outputs(761) <= b;
    layer4_outputs(762) <= a;
    layer4_outputs(763) <= not b;
    layer4_outputs(764) <= not a;
    layer4_outputs(765) <= not b;
    layer4_outputs(766) <= b;
    layer4_outputs(767) <= a xor b;
    layer4_outputs(768) <= a and b;
    layer4_outputs(769) <= b;
    layer4_outputs(770) <= not b or a;
    layer4_outputs(771) <= a and not b;
    layer4_outputs(772) <= not a or b;
    layer4_outputs(773) <= not b;
    layer4_outputs(774) <= a and b;
    layer4_outputs(775) <= not (a and b);
    layer4_outputs(776) <= not a;
    layer4_outputs(777) <= a xor b;
    layer4_outputs(778) <= a xor b;
    layer4_outputs(779) <= not a;
    layer4_outputs(780) <= not (a xor b);
    layer4_outputs(781) <= a or b;
    layer4_outputs(782) <= a or b;
    layer4_outputs(783) <= not b;
    layer4_outputs(784) <= a and not b;
    layer4_outputs(785) <= not (a xor b);
    layer4_outputs(786) <= not b;
    layer4_outputs(787) <= a;
    layer4_outputs(788) <= not (a xor b);
    layer4_outputs(789) <= a xor b;
    layer4_outputs(790) <= not b or a;
    layer4_outputs(791) <= not b or a;
    layer4_outputs(792) <= a;
    layer4_outputs(793) <= not a;
    layer4_outputs(794) <= b;
    layer4_outputs(795) <= not (a xor b);
    layer4_outputs(796) <= a xor b;
    layer4_outputs(797) <= a;
    layer4_outputs(798) <= a and not b;
    layer4_outputs(799) <= not (a xor b);
    layer4_outputs(800) <= not b;
    layer4_outputs(801) <= a and b;
    layer4_outputs(802) <= not a or b;
    layer4_outputs(803) <= not (a xor b);
    layer4_outputs(804) <= not a;
    layer4_outputs(805) <= not (a xor b);
    layer4_outputs(806) <= not a or b;
    layer4_outputs(807) <= b;
    layer4_outputs(808) <= b;
    layer4_outputs(809) <= a xor b;
    layer4_outputs(810) <= b;
    layer4_outputs(811) <= b;
    layer4_outputs(812) <= a xor b;
    layer4_outputs(813) <= not (a xor b);
    layer4_outputs(814) <= not a;
    layer4_outputs(815) <= a;
    layer4_outputs(816) <= not (a xor b);
    layer4_outputs(817) <= b;
    layer4_outputs(818) <= a and not b;
    layer4_outputs(819) <= not (a xor b);
    layer4_outputs(820) <= a xor b;
    layer4_outputs(821) <= b;
    layer4_outputs(822) <= not (a and b);
    layer4_outputs(823) <= a;
    layer4_outputs(824) <= not a;
    layer4_outputs(825) <= not b;
    layer4_outputs(826) <= a xor b;
    layer4_outputs(827) <= a and b;
    layer4_outputs(828) <= a;
    layer4_outputs(829) <= not a;
    layer4_outputs(830) <= not b;
    layer4_outputs(831) <= b;
    layer4_outputs(832) <= not (a or b);
    layer4_outputs(833) <= not a or b;
    layer4_outputs(834) <= b;
    layer4_outputs(835) <= a or b;
    layer4_outputs(836) <= b;
    layer4_outputs(837) <= a and not b;
    layer4_outputs(838) <= not (a xor b);
    layer4_outputs(839) <= a or b;
    layer4_outputs(840) <= not a;
    layer4_outputs(841) <= b;
    layer4_outputs(842) <= a;
    layer4_outputs(843) <= b and not a;
    layer4_outputs(844) <= not b;
    layer4_outputs(845) <= not (a or b);
    layer4_outputs(846) <= a xor b;
    layer4_outputs(847) <= a and not b;
    layer4_outputs(848) <= not a or b;
    layer4_outputs(849) <= not a;
    layer4_outputs(850) <= not (a or b);
    layer4_outputs(851) <= a or b;
    layer4_outputs(852) <= not b or a;
    layer4_outputs(853) <= not (a xor b);
    layer4_outputs(854) <= not (a and b);
    layer4_outputs(855) <= not b or a;
    layer4_outputs(856) <= b;
    layer4_outputs(857) <= a xor b;
    layer4_outputs(858) <= a;
    layer4_outputs(859) <= a;
    layer4_outputs(860) <= not a;
    layer4_outputs(861) <= a or b;
    layer4_outputs(862) <= a and not b;
    layer4_outputs(863) <= not a;
    layer4_outputs(864) <= not b;
    layer4_outputs(865) <= a and b;
    layer4_outputs(866) <= not (a and b);
    layer4_outputs(867) <= not a;
    layer4_outputs(868) <= not b;
    layer4_outputs(869) <= a and not b;
    layer4_outputs(870) <= not (a or b);
    layer4_outputs(871) <= not b or a;
    layer4_outputs(872) <= b;
    layer4_outputs(873) <= b and not a;
    layer4_outputs(874) <= b;
    layer4_outputs(875) <= a or b;
    layer4_outputs(876) <= a xor b;
    layer4_outputs(877) <= a;
    layer4_outputs(878) <= not a or b;
    layer4_outputs(879) <= a and b;
    layer4_outputs(880) <= not (a and b);
    layer4_outputs(881) <= not (a xor b);
    layer4_outputs(882) <= a and b;
    layer4_outputs(883) <= not (a or b);
    layer4_outputs(884) <= not b;
    layer4_outputs(885) <= a;
    layer4_outputs(886) <= a and b;
    layer4_outputs(887) <= not b;
    layer4_outputs(888) <= not b;
    layer4_outputs(889) <= a xor b;
    layer4_outputs(890) <= not b;
    layer4_outputs(891) <= b and not a;
    layer4_outputs(892) <= not (a xor b);
    layer4_outputs(893) <= not b or a;
    layer4_outputs(894) <= not a;
    layer4_outputs(895) <= a or b;
    layer4_outputs(896) <= not (a or b);
    layer4_outputs(897) <= b;
    layer4_outputs(898) <= a and b;
    layer4_outputs(899) <= a;
    layer4_outputs(900) <= not (a or b);
    layer4_outputs(901) <= a;
    layer4_outputs(902) <= a and not b;
    layer4_outputs(903) <= not b;
    layer4_outputs(904) <= b;
    layer4_outputs(905) <= not (a and b);
    layer4_outputs(906) <= b;
    layer4_outputs(907) <= a and b;
    layer4_outputs(908) <= a xor b;
    layer4_outputs(909) <= b;
    layer4_outputs(910) <= a;
    layer4_outputs(911) <= not a or b;
    layer4_outputs(912) <= a or b;
    layer4_outputs(913) <= b;
    layer4_outputs(914) <= not b;
    layer4_outputs(915) <= b;
    layer4_outputs(916) <= not b;
    layer4_outputs(917) <= not a;
    layer4_outputs(918) <= a xor b;
    layer4_outputs(919) <= not b;
    layer4_outputs(920) <= not a or b;
    layer4_outputs(921) <= a and b;
    layer4_outputs(922) <= b;
    layer4_outputs(923) <= a;
    layer4_outputs(924) <= a xor b;
    layer4_outputs(925) <= not (a or b);
    layer4_outputs(926) <= not a;
    layer4_outputs(927) <= not (a and b);
    layer4_outputs(928) <= b and not a;
    layer4_outputs(929) <= a;
    layer4_outputs(930) <= b;
    layer4_outputs(931) <= not (a xor b);
    layer4_outputs(932) <= a or b;
    layer4_outputs(933) <= a xor b;
    layer4_outputs(934) <= a xor b;
    layer4_outputs(935) <= b;
    layer4_outputs(936) <= b;
    layer4_outputs(937) <= a xor b;
    layer4_outputs(938) <= a;
    layer4_outputs(939) <= not (a or b);
    layer4_outputs(940) <= not b;
    layer4_outputs(941) <= a and not b;
    layer4_outputs(942) <= a;
    layer4_outputs(943) <= not b or a;
    layer4_outputs(944) <= not (a or b);
    layer4_outputs(945) <= a and not b;
    layer4_outputs(946) <= not b or a;
    layer4_outputs(947) <= not b or a;
    layer4_outputs(948) <= not (a xor b);
    layer4_outputs(949) <= a xor b;
    layer4_outputs(950) <= b and not a;
    layer4_outputs(951) <= not a or b;
    layer4_outputs(952) <= not (a and b);
    layer4_outputs(953) <= b;
    layer4_outputs(954) <= not (a xor b);
    layer4_outputs(955) <= not a;
    layer4_outputs(956) <= b;
    layer4_outputs(957) <= a;
    layer4_outputs(958) <= not (a xor b);
    layer4_outputs(959) <= a and not b;
    layer4_outputs(960) <= b and not a;
    layer4_outputs(961) <= b and not a;
    layer4_outputs(962) <= not a or b;
    layer4_outputs(963) <= not b;
    layer4_outputs(964) <= not (a xor b);
    layer4_outputs(965) <= b and not a;
    layer4_outputs(966) <= a and not b;
    layer4_outputs(967) <= not b;
    layer4_outputs(968) <= not a;
    layer4_outputs(969) <= not (a xor b);
    layer4_outputs(970) <= not a or b;
    layer4_outputs(971) <= not (a xor b);
    layer4_outputs(972) <= b;
    layer4_outputs(973) <= a;
    layer4_outputs(974) <= not a or b;
    layer4_outputs(975) <= a;
    layer4_outputs(976) <= b and not a;
    layer4_outputs(977) <= not (a and b);
    layer4_outputs(978) <= not b or a;
    layer4_outputs(979) <= not b;
    layer4_outputs(980) <= a xor b;
    layer4_outputs(981) <= a;
    layer4_outputs(982) <= b;
    layer4_outputs(983) <= a;
    layer4_outputs(984) <= b;
    layer4_outputs(985) <= a;
    layer4_outputs(986) <= a and not b;
    layer4_outputs(987) <= not b;
    layer4_outputs(988) <= b;
    layer4_outputs(989) <= not b or a;
    layer4_outputs(990) <= a or b;
    layer4_outputs(991) <= not (a xor b);
    layer4_outputs(992) <= a xor b;
    layer4_outputs(993) <= a xor b;
    layer4_outputs(994) <= a and b;
    layer4_outputs(995) <= a or b;
    layer4_outputs(996) <= a;
    layer4_outputs(997) <= a or b;
    layer4_outputs(998) <= not (a xor b);
    layer4_outputs(999) <= not (a xor b);
    layer4_outputs(1000) <= b and not a;
    layer4_outputs(1001) <= a xor b;
    layer4_outputs(1002) <= not (a or b);
    layer4_outputs(1003) <= not b or a;
    layer4_outputs(1004) <= not a;
    layer4_outputs(1005) <= a;
    layer4_outputs(1006) <= a and not b;
    layer4_outputs(1007) <= a and not b;
    layer4_outputs(1008) <= not (a xor b);
    layer4_outputs(1009) <= not b or a;
    layer4_outputs(1010) <= a xor b;
    layer4_outputs(1011) <= not b or a;
    layer4_outputs(1012) <= not (a and b);
    layer4_outputs(1013) <= not (a xor b);
    layer4_outputs(1014) <= a xor b;
    layer4_outputs(1015) <= a and not b;
    layer4_outputs(1016) <= a xor b;
    layer4_outputs(1017) <= a xor b;
    layer4_outputs(1018) <= 1'b1;
    layer4_outputs(1019) <= not (a and b);
    layer4_outputs(1020) <= a and b;
    layer4_outputs(1021) <= not (a xor b);
    layer4_outputs(1022) <= a;
    layer4_outputs(1023) <= not (a and b);
    layer4_outputs(1024) <= a;
    layer4_outputs(1025) <= a or b;
    layer4_outputs(1026) <= not a;
    layer4_outputs(1027) <= a;
    layer4_outputs(1028) <= not (a xor b);
    layer4_outputs(1029) <= a and not b;
    layer4_outputs(1030) <= not a or b;
    layer4_outputs(1031) <= b;
    layer4_outputs(1032) <= not b;
    layer4_outputs(1033) <= b and not a;
    layer4_outputs(1034) <= not b or a;
    layer4_outputs(1035) <= not a;
    layer4_outputs(1036) <= not (a or b);
    layer4_outputs(1037) <= b and not a;
    layer4_outputs(1038) <= not (a or b);
    layer4_outputs(1039) <= a;
    layer4_outputs(1040) <= not (a and b);
    layer4_outputs(1041) <= a xor b;
    layer4_outputs(1042) <= b and not a;
    layer4_outputs(1043) <= a;
    layer4_outputs(1044) <= not a;
    layer4_outputs(1045) <= not (a xor b);
    layer4_outputs(1046) <= not b or a;
    layer4_outputs(1047) <= a or b;
    layer4_outputs(1048) <= not b or a;
    layer4_outputs(1049) <= a and not b;
    layer4_outputs(1050) <= not (a xor b);
    layer4_outputs(1051) <= not (a xor b);
    layer4_outputs(1052) <= not b or a;
    layer4_outputs(1053) <= not (a and b);
    layer4_outputs(1054) <= a and not b;
    layer4_outputs(1055) <= a or b;
    layer4_outputs(1056) <= a;
    layer4_outputs(1057) <= not (a and b);
    layer4_outputs(1058) <= b;
    layer4_outputs(1059) <= not a;
    layer4_outputs(1060) <= b;
    layer4_outputs(1061) <= b and not a;
    layer4_outputs(1062) <= not a;
    layer4_outputs(1063) <= b;
    layer4_outputs(1064) <= a xor b;
    layer4_outputs(1065) <= a xor b;
    layer4_outputs(1066) <= b;
    layer4_outputs(1067) <= a xor b;
    layer4_outputs(1068) <= b;
    layer4_outputs(1069) <= a xor b;
    layer4_outputs(1070) <= not b;
    layer4_outputs(1071) <= 1'b0;
    layer4_outputs(1072) <= not b;
    layer4_outputs(1073) <= b;
    layer4_outputs(1074) <= not (a or b);
    layer4_outputs(1075) <= not b;
    layer4_outputs(1076) <= a;
    layer4_outputs(1077) <= a;
    layer4_outputs(1078) <= a or b;
    layer4_outputs(1079) <= b and not a;
    layer4_outputs(1080) <= b and not a;
    layer4_outputs(1081) <= b;
    layer4_outputs(1082) <= a or b;
    layer4_outputs(1083) <= not a;
    layer4_outputs(1084) <= a or b;
    layer4_outputs(1085) <= a or b;
    layer4_outputs(1086) <= not b;
    layer4_outputs(1087) <= b;
    layer4_outputs(1088) <= not b;
    layer4_outputs(1089) <= b;
    layer4_outputs(1090) <= a xor b;
    layer4_outputs(1091) <= not b;
    layer4_outputs(1092) <= b;
    layer4_outputs(1093) <= b;
    layer4_outputs(1094) <= a and not b;
    layer4_outputs(1095) <= a xor b;
    layer4_outputs(1096) <= not (a xor b);
    layer4_outputs(1097) <= not b;
    layer4_outputs(1098) <= a and not b;
    layer4_outputs(1099) <= b;
    layer4_outputs(1100) <= b and not a;
    layer4_outputs(1101) <= a and b;
    layer4_outputs(1102) <= b;
    layer4_outputs(1103) <= a and b;
    layer4_outputs(1104) <= b;
    layer4_outputs(1105) <= a;
    layer4_outputs(1106) <= a and b;
    layer4_outputs(1107) <= b and not a;
    layer4_outputs(1108) <= a xor b;
    layer4_outputs(1109) <= a and not b;
    layer4_outputs(1110) <= not a;
    layer4_outputs(1111) <= a xor b;
    layer4_outputs(1112) <= not b;
    layer4_outputs(1113) <= not a or b;
    layer4_outputs(1114) <= a and not b;
    layer4_outputs(1115) <= not a;
    layer4_outputs(1116) <= not (a or b);
    layer4_outputs(1117) <= b and not a;
    layer4_outputs(1118) <= a;
    layer4_outputs(1119) <= not a;
    layer4_outputs(1120) <= a;
    layer4_outputs(1121) <= a xor b;
    layer4_outputs(1122) <= not (a xor b);
    layer4_outputs(1123) <= not b;
    layer4_outputs(1124) <= a xor b;
    layer4_outputs(1125) <= not (a xor b);
    layer4_outputs(1126) <= 1'b0;
    layer4_outputs(1127) <= not a or b;
    layer4_outputs(1128) <= a;
    layer4_outputs(1129) <= not b;
    layer4_outputs(1130) <= a and b;
    layer4_outputs(1131) <= a xor b;
    layer4_outputs(1132) <= a and not b;
    layer4_outputs(1133) <= not (a and b);
    layer4_outputs(1134) <= not a;
    layer4_outputs(1135) <= a;
    layer4_outputs(1136) <= not (a and b);
    layer4_outputs(1137) <= b and not a;
    layer4_outputs(1138) <= not a or b;
    layer4_outputs(1139) <= a and not b;
    layer4_outputs(1140) <= a and b;
    layer4_outputs(1141) <= not (a or b);
    layer4_outputs(1142) <= b;
    layer4_outputs(1143) <= b and not a;
    layer4_outputs(1144) <= not (a xor b);
    layer4_outputs(1145) <= a or b;
    layer4_outputs(1146) <= a xor b;
    layer4_outputs(1147) <= a;
    layer4_outputs(1148) <= b;
    layer4_outputs(1149) <= not (a or b);
    layer4_outputs(1150) <= not b or a;
    layer4_outputs(1151) <= b;
    layer4_outputs(1152) <= a;
    layer4_outputs(1153) <= not (a xor b);
    layer4_outputs(1154) <= not a;
    layer4_outputs(1155) <= not (a and b);
    layer4_outputs(1156) <= a;
    layer4_outputs(1157) <= not b or a;
    layer4_outputs(1158) <= a;
    layer4_outputs(1159) <= not a;
    layer4_outputs(1160) <= b;
    layer4_outputs(1161) <= not b;
    layer4_outputs(1162) <= b;
    layer4_outputs(1163) <= not (a or b);
    layer4_outputs(1164) <= b;
    layer4_outputs(1165) <= not b;
    layer4_outputs(1166) <= a xor b;
    layer4_outputs(1167) <= not b;
    layer4_outputs(1168) <= not (a and b);
    layer4_outputs(1169) <= a;
    layer4_outputs(1170) <= not b;
    layer4_outputs(1171) <= not (a or b);
    layer4_outputs(1172) <= a and not b;
    layer4_outputs(1173) <= not a;
    layer4_outputs(1174) <= a xor b;
    layer4_outputs(1175) <= not b or a;
    layer4_outputs(1176) <= b;
    layer4_outputs(1177) <= not b;
    layer4_outputs(1178) <= not a or b;
    layer4_outputs(1179) <= not a;
    layer4_outputs(1180) <= not (a xor b);
    layer4_outputs(1181) <= b;
    layer4_outputs(1182) <= not b;
    layer4_outputs(1183) <= b;
    layer4_outputs(1184) <= a and not b;
    layer4_outputs(1185) <= a xor b;
    layer4_outputs(1186) <= a and b;
    layer4_outputs(1187) <= a;
    layer4_outputs(1188) <= not (a or b);
    layer4_outputs(1189) <= a;
    layer4_outputs(1190) <= b;
    layer4_outputs(1191) <= b;
    layer4_outputs(1192) <= not a;
    layer4_outputs(1193) <= not (a xor b);
    layer4_outputs(1194) <= not b;
    layer4_outputs(1195) <= a;
    layer4_outputs(1196) <= not (a and b);
    layer4_outputs(1197) <= b;
    layer4_outputs(1198) <= a;
    layer4_outputs(1199) <= not a;
    layer4_outputs(1200) <= not (a xor b);
    layer4_outputs(1201) <= a;
    layer4_outputs(1202) <= not a;
    layer4_outputs(1203) <= a xor b;
    layer4_outputs(1204) <= a;
    layer4_outputs(1205) <= not b or a;
    layer4_outputs(1206) <= b;
    layer4_outputs(1207) <= not (a xor b);
    layer4_outputs(1208) <= not (a xor b);
    layer4_outputs(1209) <= a and not b;
    layer4_outputs(1210) <= not b or a;
    layer4_outputs(1211) <= not b;
    layer4_outputs(1212) <= not a;
    layer4_outputs(1213) <= a xor b;
    layer4_outputs(1214) <= a and b;
    layer4_outputs(1215) <= not (a xor b);
    layer4_outputs(1216) <= a;
    layer4_outputs(1217) <= a or b;
    layer4_outputs(1218) <= a;
    layer4_outputs(1219) <= b;
    layer4_outputs(1220) <= a;
    layer4_outputs(1221) <= not (a or b);
    layer4_outputs(1222) <= not (a and b);
    layer4_outputs(1223) <= not a;
    layer4_outputs(1224) <= b;
    layer4_outputs(1225) <= b;
    layer4_outputs(1226) <= b and not a;
    layer4_outputs(1227) <= not (a xor b);
    layer4_outputs(1228) <= b and not a;
    layer4_outputs(1229) <= a or b;
    layer4_outputs(1230) <= not b;
    layer4_outputs(1231) <= a and b;
    layer4_outputs(1232) <= not b;
    layer4_outputs(1233) <= not (a or b);
    layer4_outputs(1234) <= a or b;
    layer4_outputs(1235) <= not b;
    layer4_outputs(1236) <= a xor b;
    layer4_outputs(1237) <= not a;
    layer4_outputs(1238) <= not (a and b);
    layer4_outputs(1239) <= not (a xor b);
    layer4_outputs(1240) <= not a;
    layer4_outputs(1241) <= b;
    layer4_outputs(1242) <= not (a xor b);
    layer4_outputs(1243) <= not a;
    layer4_outputs(1244) <= not b;
    layer4_outputs(1245) <= a and b;
    layer4_outputs(1246) <= not a;
    layer4_outputs(1247) <= not (a and b);
    layer4_outputs(1248) <= a or b;
    layer4_outputs(1249) <= a;
    layer4_outputs(1250) <= not a;
    layer4_outputs(1251) <= b and not a;
    layer4_outputs(1252) <= not b;
    layer4_outputs(1253) <= b;
    layer4_outputs(1254) <= not (a xor b);
    layer4_outputs(1255) <= not (a xor b);
    layer4_outputs(1256) <= a and b;
    layer4_outputs(1257) <= a;
    layer4_outputs(1258) <= not b;
    layer4_outputs(1259) <= a;
    layer4_outputs(1260) <= a;
    layer4_outputs(1261) <= not (a and b);
    layer4_outputs(1262) <= b;
    layer4_outputs(1263) <= not b or a;
    layer4_outputs(1264) <= not b or a;
    layer4_outputs(1265) <= a and not b;
    layer4_outputs(1266) <= not (a or b);
    layer4_outputs(1267) <= a;
    layer4_outputs(1268) <= not (a xor b);
    layer4_outputs(1269) <= not (a xor b);
    layer4_outputs(1270) <= not b;
    layer4_outputs(1271) <= a or b;
    layer4_outputs(1272) <= not b;
    layer4_outputs(1273) <= 1'b1;
    layer4_outputs(1274) <= b;
    layer4_outputs(1275) <= not (a xor b);
    layer4_outputs(1276) <= not b;
    layer4_outputs(1277) <= a or b;
    layer4_outputs(1278) <= b;
    layer4_outputs(1279) <= not a or b;
    layer4_outputs(1280) <= a or b;
    layer4_outputs(1281) <= b;
    layer4_outputs(1282) <= not (a and b);
    layer4_outputs(1283) <= a and b;
    layer4_outputs(1284) <= a;
    layer4_outputs(1285) <= not a or b;
    layer4_outputs(1286) <= b;
    layer4_outputs(1287) <= a;
    layer4_outputs(1288) <= not a;
    layer4_outputs(1289) <= b;
    layer4_outputs(1290) <= a xor b;
    layer4_outputs(1291) <= a;
    layer4_outputs(1292) <= not (a xor b);
    layer4_outputs(1293) <= not (a or b);
    layer4_outputs(1294) <= not b or a;
    layer4_outputs(1295) <= a xor b;
    layer4_outputs(1296) <= not a or b;
    layer4_outputs(1297) <= not b;
    layer4_outputs(1298) <= not a or b;
    layer4_outputs(1299) <= not b or a;
    layer4_outputs(1300) <= a and b;
    layer4_outputs(1301) <= not b;
    layer4_outputs(1302) <= not (a or b);
    layer4_outputs(1303) <= 1'b0;
    layer4_outputs(1304) <= a xor b;
    layer4_outputs(1305) <= a and b;
    layer4_outputs(1306) <= not (a or b);
    layer4_outputs(1307) <= not (a and b);
    layer4_outputs(1308) <= a or b;
    layer4_outputs(1309) <= not b or a;
    layer4_outputs(1310) <= not a;
    layer4_outputs(1311) <= b and not a;
    layer4_outputs(1312) <= a and not b;
    layer4_outputs(1313) <= not a;
    layer4_outputs(1314) <= not a or b;
    layer4_outputs(1315) <= not (a xor b);
    layer4_outputs(1316) <= b and not a;
    layer4_outputs(1317) <= a or b;
    layer4_outputs(1318) <= not (a xor b);
    layer4_outputs(1319) <= b;
    layer4_outputs(1320) <= a;
    layer4_outputs(1321) <= not b;
    layer4_outputs(1322) <= not b;
    layer4_outputs(1323) <= not (a and b);
    layer4_outputs(1324) <= a xor b;
    layer4_outputs(1325) <= b and not a;
    layer4_outputs(1326) <= b;
    layer4_outputs(1327) <= 1'b0;
    layer4_outputs(1328) <= a or b;
    layer4_outputs(1329) <= b;
    layer4_outputs(1330) <= a xor b;
    layer4_outputs(1331) <= not (a or b);
    layer4_outputs(1332) <= a and not b;
    layer4_outputs(1333) <= a xor b;
    layer4_outputs(1334) <= not (a and b);
    layer4_outputs(1335) <= not (a and b);
    layer4_outputs(1336) <= not b or a;
    layer4_outputs(1337) <= b;
    layer4_outputs(1338) <= not b;
    layer4_outputs(1339) <= a;
    layer4_outputs(1340) <= not b;
    layer4_outputs(1341) <= not (a or b);
    layer4_outputs(1342) <= not (a and b);
    layer4_outputs(1343) <= b;
    layer4_outputs(1344) <= not a or b;
    layer4_outputs(1345) <= a and not b;
    layer4_outputs(1346) <= a and not b;
    layer4_outputs(1347) <= not (a xor b);
    layer4_outputs(1348) <= not b or a;
    layer4_outputs(1349) <= not (a xor b);
    layer4_outputs(1350) <= a;
    layer4_outputs(1351) <= a;
    layer4_outputs(1352) <= not a or b;
    layer4_outputs(1353) <= not (a xor b);
    layer4_outputs(1354) <= a xor b;
    layer4_outputs(1355) <= a or b;
    layer4_outputs(1356) <= b;
    layer4_outputs(1357) <= b;
    layer4_outputs(1358) <= 1'b0;
    layer4_outputs(1359) <= not b;
    layer4_outputs(1360) <= b;
    layer4_outputs(1361) <= not a;
    layer4_outputs(1362) <= b and not a;
    layer4_outputs(1363) <= b;
    layer4_outputs(1364) <= b and not a;
    layer4_outputs(1365) <= not (a and b);
    layer4_outputs(1366) <= not (a and b);
    layer4_outputs(1367) <= b;
    layer4_outputs(1368) <= not a;
    layer4_outputs(1369) <= a;
    layer4_outputs(1370) <= b;
    layer4_outputs(1371) <= a and not b;
    layer4_outputs(1372) <= not a;
    layer4_outputs(1373) <= not b;
    layer4_outputs(1374) <= not (a xor b);
    layer4_outputs(1375) <= not b;
    layer4_outputs(1376) <= not (a and b);
    layer4_outputs(1377) <= a or b;
    layer4_outputs(1378) <= a and b;
    layer4_outputs(1379) <= not a;
    layer4_outputs(1380) <= not b;
    layer4_outputs(1381) <= a xor b;
    layer4_outputs(1382) <= b;
    layer4_outputs(1383) <= a and b;
    layer4_outputs(1384) <= a;
    layer4_outputs(1385) <= a;
    layer4_outputs(1386) <= a;
    layer4_outputs(1387) <= b;
    layer4_outputs(1388) <= a xor b;
    layer4_outputs(1389) <= not a or b;
    layer4_outputs(1390) <= not (a and b);
    layer4_outputs(1391) <= not b;
    layer4_outputs(1392) <= a or b;
    layer4_outputs(1393) <= not a;
    layer4_outputs(1394) <= not a;
    layer4_outputs(1395) <= not b;
    layer4_outputs(1396) <= not (a xor b);
    layer4_outputs(1397) <= b and not a;
    layer4_outputs(1398) <= not b;
    layer4_outputs(1399) <= not (a xor b);
    layer4_outputs(1400) <= not (a and b);
    layer4_outputs(1401) <= not b or a;
    layer4_outputs(1402) <= b and not a;
    layer4_outputs(1403) <= a;
    layer4_outputs(1404) <= a;
    layer4_outputs(1405) <= a xor b;
    layer4_outputs(1406) <= a;
    layer4_outputs(1407) <= not (a and b);
    layer4_outputs(1408) <= b and not a;
    layer4_outputs(1409) <= not (a xor b);
    layer4_outputs(1410) <= b and not a;
    layer4_outputs(1411) <= not a;
    layer4_outputs(1412) <= not (a and b);
    layer4_outputs(1413) <= not b;
    layer4_outputs(1414) <= b;
    layer4_outputs(1415) <= b;
    layer4_outputs(1416) <= b;
    layer4_outputs(1417) <= not b or a;
    layer4_outputs(1418) <= not b;
    layer4_outputs(1419) <= not a;
    layer4_outputs(1420) <= a xor b;
    layer4_outputs(1421) <= not b;
    layer4_outputs(1422) <= a;
    layer4_outputs(1423) <= a;
    layer4_outputs(1424) <= b;
    layer4_outputs(1425) <= not a;
    layer4_outputs(1426) <= not b;
    layer4_outputs(1427) <= not b;
    layer4_outputs(1428) <= a;
    layer4_outputs(1429) <= a;
    layer4_outputs(1430) <= a or b;
    layer4_outputs(1431) <= b;
    layer4_outputs(1432) <= not (a xor b);
    layer4_outputs(1433) <= a or b;
    layer4_outputs(1434) <= not a;
    layer4_outputs(1435) <= not (a and b);
    layer4_outputs(1436) <= not (a and b);
    layer4_outputs(1437) <= not a;
    layer4_outputs(1438) <= not b;
    layer4_outputs(1439) <= a;
    layer4_outputs(1440) <= not (a and b);
    layer4_outputs(1441) <= a and b;
    layer4_outputs(1442) <= a and not b;
    layer4_outputs(1443) <= a;
    layer4_outputs(1444) <= not a or b;
    layer4_outputs(1445) <= b and not a;
    layer4_outputs(1446) <= a xor b;
    layer4_outputs(1447) <= not a or b;
    layer4_outputs(1448) <= b;
    layer4_outputs(1449) <= b and not a;
    layer4_outputs(1450) <= a and not b;
    layer4_outputs(1451) <= a and b;
    layer4_outputs(1452) <= not b;
    layer4_outputs(1453) <= a xor b;
    layer4_outputs(1454) <= not (a xor b);
    layer4_outputs(1455) <= b;
    layer4_outputs(1456) <= a;
    layer4_outputs(1457) <= not a;
    layer4_outputs(1458) <= a;
    layer4_outputs(1459) <= b;
    layer4_outputs(1460) <= a xor b;
    layer4_outputs(1461) <= not a or b;
    layer4_outputs(1462) <= a and not b;
    layer4_outputs(1463) <= not a;
    layer4_outputs(1464) <= not a;
    layer4_outputs(1465) <= not a;
    layer4_outputs(1466) <= b;
    layer4_outputs(1467) <= a xor b;
    layer4_outputs(1468) <= a;
    layer4_outputs(1469) <= a and not b;
    layer4_outputs(1470) <= a and b;
    layer4_outputs(1471) <= not a;
    layer4_outputs(1472) <= a or b;
    layer4_outputs(1473) <= not (a or b);
    layer4_outputs(1474) <= a xor b;
    layer4_outputs(1475) <= a or b;
    layer4_outputs(1476) <= b;
    layer4_outputs(1477) <= not a;
    layer4_outputs(1478) <= not (a or b);
    layer4_outputs(1479) <= 1'b0;
    layer4_outputs(1480) <= a and not b;
    layer4_outputs(1481) <= not a or b;
    layer4_outputs(1482) <= not a or b;
    layer4_outputs(1483) <= b;
    layer4_outputs(1484) <= a or b;
    layer4_outputs(1485) <= b and not a;
    layer4_outputs(1486) <= not a or b;
    layer4_outputs(1487) <= not (a xor b);
    layer4_outputs(1488) <= a;
    layer4_outputs(1489) <= not a;
    layer4_outputs(1490) <= not (a or b);
    layer4_outputs(1491) <= a or b;
    layer4_outputs(1492) <= not b;
    layer4_outputs(1493) <= not a or b;
    layer4_outputs(1494) <= not a or b;
    layer4_outputs(1495) <= not b;
    layer4_outputs(1496) <= not (a or b);
    layer4_outputs(1497) <= b;
    layer4_outputs(1498) <= not (a xor b);
    layer4_outputs(1499) <= b;
    layer4_outputs(1500) <= a and not b;
    layer4_outputs(1501) <= a;
    layer4_outputs(1502) <= not b;
    layer4_outputs(1503) <= not b;
    layer4_outputs(1504) <= not (a and b);
    layer4_outputs(1505) <= a and not b;
    layer4_outputs(1506) <= not b;
    layer4_outputs(1507) <= not b or a;
    layer4_outputs(1508) <= not a;
    layer4_outputs(1509) <= not (a and b);
    layer4_outputs(1510) <= not (a xor b);
    layer4_outputs(1511) <= a and not b;
    layer4_outputs(1512) <= a or b;
    layer4_outputs(1513) <= not (a xor b);
    layer4_outputs(1514) <= b;
    layer4_outputs(1515) <= not (a xor b);
    layer4_outputs(1516) <= a;
    layer4_outputs(1517) <= a xor b;
    layer4_outputs(1518) <= not a;
    layer4_outputs(1519) <= not b or a;
    layer4_outputs(1520) <= b;
    layer4_outputs(1521) <= b;
    layer4_outputs(1522) <= b;
    layer4_outputs(1523) <= not b;
    layer4_outputs(1524) <= not (a or b);
    layer4_outputs(1525) <= not b;
    layer4_outputs(1526) <= a;
    layer4_outputs(1527) <= a xor b;
    layer4_outputs(1528) <= a and b;
    layer4_outputs(1529) <= b;
    layer4_outputs(1530) <= not b;
    layer4_outputs(1531) <= not b;
    layer4_outputs(1532) <= a and not b;
    layer4_outputs(1533) <= a xor b;
    layer4_outputs(1534) <= b and not a;
    layer4_outputs(1535) <= a and b;
    layer4_outputs(1536) <= not b;
    layer4_outputs(1537) <= not (a xor b);
    layer4_outputs(1538) <= a xor b;
    layer4_outputs(1539) <= not (a or b);
    layer4_outputs(1540) <= not b or a;
    layer4_outputs(1541) <= a xor b;
    layer4_outputs(1542) <= not a or b;
    layer4_outputs(1543) <= a or b;
    layer4_outputs(1544) <= not a or b;
    layer4_outputs(1545) <= a and b;
    layer4_outputs(1546) <= a xor b;
    layer4_outputs(1547) <= a and not b;
    layer4_outputs(1548) <= not (a xor b);
    layer4_outputs(1549) <= a xor b;
    layer4_outputs(1550) <= not (a and b);
    layer4_outputs(1551) <= not (a or b);
    layer4_outputs(1552) <= not (a xor b);
    layer4_outputs(1553) <= b;
    layer4_outputs(1554) <= not (a xor b);
    layer4_outputs(1555) <= b;
    layer4_outputs(1556) <= a and not b;
    layer4_outputs(1557) <= a;
    layer4_outputs(1558) <= a xor b;
    layer4_outputs(1559) <= a and b;
    layer4_outputs(1560) <= a or b;
    layer4_outputs(1561) <= not (a xor b);
    layer4_outputs(1562) <= not b or a;
    layer4_outputs(1563) <= not a or b;
    layer4_outputs(1564) <= not a;
    layer4_outputs(1565) <= not a;
    layer4_outputs(1566) <= not b;
    layer4_outputs(1567) <= a xor b;
    layer4_outputs(1568) <= a;
    layer4_outputs(1569) <= a and b;
    layer4_outputs(1570) <= a;
    layer4_outputs(1571) <= not (a and b);
    layer4_outputs(1572) <= not (a or b);
    layer4_outputs(1573) <= a and b;
    layer4_outputs(1574) <= b and not a;
    layer4_outputs(1575) <= b;
    layer4_outputs(1576) <= not a;
    layer4_outputs(1577) <= not (a xor b);
    layer4_outputs(1578) <= not b;
    layer4_outputs(1579) <= not a or b;
    layer4_outputs(1580) <= a xor b;
    layer4_outputs(1581) <= not (a and b);
    layer4_outputs(1582) <= b;
    layer4_outputs(1583) <= a xor b;
    layer4_outputs(1584) <= b and not a;
    layer4_outputs(1585) <= not a or b;
    layer4_outputs(1586) <= a and not b;
    layer4_outputs(1587) <= not (a xor b);
    layer4_outputs(1588) <= b;
    layer4_outputs(1589) <= a and b;
    layer4_outputs(1590) <= a and b;
    layer4_outputs(1591) <= b and not a;
    layer4_outputs(1592) <= b;
    layer4_outputs(1593) <= not b;
    layer4_outputs(1594) <= not (a or b);
    layer4_outputs(1595) <= not b;
    layer4_outputs(1596) <= a;
    layer4_outputs(1597) <= not b;
    layer4_outputs(1598) <= not (a and b);
    layer4_outputs(1599) <= a or b;
    layer4_outputs(1600) <= a and b;
    layer4_outputs(1601) <= a xor b;
    layer4_outputs(1602) <= a;
    layer4_outputs(1603) <= not a;
    layer4_outputs(1604) <= a;
    layer4_outputs(1605) <= b;
    layer4_outputs(1606) <= not a;
    layer4_outputs(1607) <= 1'b0;
    layer4_outputs(1608) <= a xor b;
    layer4_outputs(1609) <= a xor b;
    layer4_outputs(1610) <= not b;
    layer4_outputs(1611) <= not (a xor b);
    layer4_outputs(1612) <= not (a xor b);
    layer4_outputs(1613) <= not b;
    layer4_outputs(1614) <= not b;
    layer4_outputs(1615) <= b;
    layer4_outputs(1616) <= not a or b;
    layer4_outputs(1617) <= a;
    layer4_outputs(1618) <= not a;
    layer4_outputs(1619) <= not b;
    layer4_outputs(1620) <= not b;
    layer4_outputs(1621) <= b and not a;
    layer4_outputs(1622) <= not b or a;
    layer4_outputs(1623) <= not a;
    layer4_outputs(1624) <= a xor b;
    layer4_outputs(1625) <= not (a xor b);
    layer4_outputs(1626) <= b;
    layer4_outputs(1627) <= b and not a;
    layer4_outputs(1628) <= a or b;
    layer4_outputs(1629) <= b;
    layer4_outputs(1630) <= not b;
    layer4_outputs(1631) <= not b;
    layer4_outputs(1632) <= b;
    layer4_outputs(1633) <= a xor b;
    layer4_outputs(1634) <= a and not b;
    layer4_outputs(1635) <= b and not a;
    layer4_outputs(1636) <= b;
    layer4_outputs(1637) <= 1'b0;
    layer4_outputs(1638) <= 1'b1;
    layer4_outputs(1639) <= a or b;
    layer4_outputs(1640) <= b and not a;
    layer4_outputs(1641) <= b and not a;
    layer4_outputs(1642) <= not b;
    layer4_outputs(1643) <= a or b;
    layer4_outputs(1644) <= a or b;
    layer4_outputs(1645) <= a;
    layer4_outputs(1646) <= a and not b;
    layer4_outputs(1647) <= a or b;
    layer4_outputs(1648) <= a or b;
    layer4_outputs(1649) <= b and not a;
    layer4_outputs(1650) <= a or b;
    layer4_outputs(1651) <= b;
    layer4_outputs(1652) <= not a;
    layer4_outputs(1653) <= b;
    layer4_outputs(1654) <= a and b;
    layer4_outputs(1655) <= a or b;
    layer4_outputs(1656) <= not a;
    layer4_outputs(1657) <= a xor b;
    layer4_outputs(1658) <= not (a or b);
    layer4_outputs(1659) <= b;
    layer4_outputs(1660) <= not a;
    layer4_outputs(1661) <= not a or b;
    layer4_outputs(1662) <= a;
    layer4_outputs(1663) <= a and not b;
    layer4_outputs(1664) <= not b or a;
    layer4_outputs(1665) <= not b or a;
    layer4_outputs(1666) <= a xor b;
    layer4_outputs(1667) <= a xor b;
    layer4_outputs(1668) <= b;
    layer4_outputs(1669) <= not (a and b);
    layer4_outputs(1670) <= not a;
    layer4_outputs(1671) <= not b;
    layer4_outputs(1672) <= not b;
    layer4_outputs(1673) <= not b or a;
    layer4_outputs(1674) <= b;
    layer4_outputs(1675) <= not (a xor b);
    layer4_outputs(1676) <= b and not a;
    layer4_outputs(1677) <= a xor b;
    layer4_outputs(1678) <= b and not a;
    layer4_outputs(1679) <= not (a and b);
    layer4_outputs(1680) <= not a;
    layer4_outputs(1681) <= not (a xor b);
    layer4_outputs(1682) <= not b;
    layer4_outputs(1683) <= b;
    layer4_outputs(1684) <= not b;
    layer4_outputs(1685) <= b;
    layer4_outputs(1686) <= not a;
    layer4_outputs(1687) <= a or b;
    layer4_outputs(1688) <= not a;
    layer4_outputs(1689) <= not (a xor b);
    layer4_outputs(1690) <= not b;
    layer4_outputs(1691) <= not b or a;
    layer4_outputs(1692) <= a;
    layer4_outputs(1693) <= not (a or b);
    layer4_outputs(1694) <= b and not a;
    layer4_outputs(1695) <= not (a xor b);
    layer4_outputs(1696) <= a or b;
    layer4_outputs(1697) <= not b or a;
    layer4_outputs(1698) <= not b;
    layer4_outputs(1699) <= a xor b;
    layer4_outputs(1700) <= a or b;
    layer4_outputs(1701) <= b;
    layer4_outputs(1702) <= not (a and b);
    layer4_outputs(1703) <= b;
    layer4_outputs(1704) <= not a;
    layer4_outputs(1705) <= not a;
    layer4_outputs(1706) <= not (a xor b);
    layer4_outputs(1707) <= b;
    layer4_outputs(1708) <= a xor b;
    layer4_outputs(1709) <= not b;
    layer4_outputs(1710) <= not b;
    layer4_outputs(1711) <= b;
    layer4_outputs(1712) <= b;
    layer4_outputs(1713) <= not a;
    layer4_outputs(1714) <= b;
    layer4_outputs(1715) <= a or b;
    layer4_outputs(1716) <= not b or a;
    layer4_outputs(1717) <= b;
    layer4_outputs(1718) <= not b or a;
    layer4_outputs(1719) <= not (a or b);
    layer4_outputs(1720) <= b;
    layer4_outputs(1721) <= not b;
    layer4_outputs(1722) <= a or b;
    layer4_outputs(1723) <= not b;
    layer4_outputs(1724) <= a and not b;
    layer4_outputs(1725) <= b;
    layer4_outputs(1726) <= a;
    layer4_outputs(1727) <= not b or a;
    layer4_outputs(1728) <= not b;
    layer4_outputs(1729) <= not a or b;
    layer4_outputs(1730) <= not a;
    layer4_outputs(1731) <= a;
    layer4_outputs(1732) <= not (a or b);
    layer4_outputs(1733) <= not b;
    layer4_outputs(1734) <= not (a xor b);
    layer4_outputs(1735) <= not (a xor b);
    layer4_outputs(1736) <= not a or b;
    layer4_outputs(1737) <= not b;
    layer4_outputs(1738) <= a or b;
    layer4_outputs(1739) <= not (a or b);
    layer4_outputs(1740) <= not b;
    layer4_outputs(1741) <= a;
    layer4_outputs(1742) <= b;
    layer4_outputs(1743) <= not (a xor b);
    layer4_outputs(1744) <= b;
    layer4_outputs(1745) <= not b;
    layer4_outputs(1746) <= a and b;
    layer4_outputs(1747) <= b;
    layer4_outputs(1748) <= not (a or b);
    layer4_outputs(1749) <= a;
    layer4_outputs(1750) <= a xor b;
    layer4_outputs(1751) <= not b or a;
    layer4_outputs(1752) <= a xor b;
    layer4_outputs(1753) <= not a or b;
    layer4_outputs(1754) <= not b;
    layer4_outputs(1755) <= not (a xor b);
    layer4_outputs(1756) <= a xor b;
    layer4_outputs(1757) <= a and b;
    layer4_outputs(1758) <= a xor b;
    layer4_outputs(1759) <= a or b;
    layer4_outputs(1760) <= not (a xor b);
    layer4_outputs(1761) <= a and b;
    layer4_outputs(1762) <= a and b;
    layer4_outputs(1763) <= not (a or b);
    layer4_outputs(1764) <= not b;
    layer4_outputs(1765) <= not a;
    layer4_outputs(1766) <= not (a xor b);
    layer4_outputs(1767) <= not (a or b);
    layer4_outputs(1768) <= a and not b;
    layer4_outputs(1769) <= not a;
    layer4_outputs(1770) <= a and not b;
    layer4_outputs(1771) <= a;
    layer4_outputs(1772) <= not a;
    layer4_outputs(1773) <= not (a and b);
    layer4_outputs(1774) <= not b;
    layer4_outputs(1775) <= not b or a;
    layer4_outputs(1776) <= not b;
    layer4_outputs(1777) <= a xor b;
    layer4_outputs(1778) <= not a or b;
    layer4_outputs(1779) <= not (a and b);
    layer4_outputs(1780) <= not (a xor b);
    layer4_outputs(1781) <= a;
    layer4_outputs(1782) <= a or b;
    layer4_outputs(1783) <= a;
    layer4_outputs(1784) <= b;
    layer4_outputs(1785) <= not (a or b);
    layer4_outputs(1786) <= b;
    layer4_outputs(1787) <= not b;
    layer4_outputs(1788) <= not (a or b);
    layer4_outputs(1789) <= b;
    layer4_outputs(1790) <= not (a xor b);
    layer4_outputs(1791) <= not (a and b);
    layer4_outputs(1792) <= not (a or b);
    layer4_outputs(1793) <= not a;
    layer4_outputs(1794) <= b;
    layer4_outputs(1795) <= not a;
    layer4_outputs(1796) <= not (a and b);
    layer4_outputs(1797) <= not (a xor b);
    layer4_outputs(1798) <= not a;
    layer4_outputs(1799) <= a or b;
    layer4_outputs(1800) <= not (a xor b);
    layer4_outputs(1801) <= a;
    layer4_outputs(1802) <= a;
    layer4_outputs(1803) <= not (a or b);
    layer4_outputs(1804) <= a and not b;
    layer4_outputs(1805) <= a xor b;
    layer4_outputs(1806) <= a;
    layer4_outputs(1807) <= a xor b;
    layer4_outputs(1808) <= a xor b;
    layer4_outputs(1809) <= not (a or b);
    layer4_outputs(1810) <= not (a or b);
    layer4_outputs(1811) <= b;
    layer4_outputs(1812) <= not a;
    layer4_outputs(1813) <= a or b;
    layer4_outputs(1814) <= a or b;
    layer4_outputs(1815) <= not a;
    layer4_outputs(1816) <= a;
    layer4_outputs(1817) <= a;
    layer4_outputs(1818) <= not a;
    layer4_outputs(1819) <= a and not b;
    layer4_outputs(1820) <= not (a xor b);
    layer4_outputs(1821) <= not b;
    layer4_outputs(1822) <= a;
    layer4_outputs(1823) <= not (a xor b);
    layer4_outputs(1824) <= a;
    layer4_outputs(1825) <= b;
    layer4_outputs(1826) <= not (a and b);
    layer4_outputs(1827) <= not b;
    layer4_outputs(1828) <= not (a xor b);
    layer4_outputs(1829) <= not (a or b);
    layer4_outputs(1830) <= a and b;
    layer4_outputs(1831) <= not a;
    layer4_outputs(1832) <= not a;
    layer4_outputs(1833) <= not b;
    layer4_outputs(1834) <= a and not b;
    layer4_outputs(1835) <= a;
    layer4_outputs(1836) <= not b;
    layer4_outputs(1837) <= a and not b;
    layer4_outputs(1838) <= not (a or b);
    layer4_outputs(1839) <= a;
    layer4_outputs(1840) <= not a;
    layer4_outputs(1841) <= not (a xor b);
    layer4_outputs(1842) <= not b;
    layer4_outputs(1843) <= not b;
    layer4_outputs(1844) <= b;
    layer4_outputs(1845) <= a xor b;
    layer4_outputs(1846) <= not a;
    layer4_outputs(1847) <= not b or a;
    layer4_outputs(1848) <= not b or a;
    layer4_outputs(1849) <= a xor b;
    layer4_outputs(1850) <= not (a and b);
    layer4_outputs(1851) <= not b;
    layer4_outputs(1852) <= not b;
    layer4_outputs(1853) <= not (a or b);
    layer4_outputs(1854) <= not b or a;
    layer4_outputs(1855) <= not b or a;
    layer4_outputs(1856) <= b;
    layer4_outputs(1857) <= not b;
    layer4_outputs(1858) <= a and not b;
    layer4_outputs(1859) <= not (a xor b);
    layer4_outputs(1860) <= b and not a;
    layer4_outputs(1861) <= not b;
    layer4_outputs(1862) <= a or b;
    layer4_outputs(1863) <= a;
    layer4_outputs(1864) <= not a;
    layer4_outputs(1865) <= not (a xor b);
    layer4_outputs(1866) <= not (a and b);
    layer4_outputs(1867) <= b;
    layer4_outputs(1868) <= not (a or b);
    layer4_outputs(1869) <= b;
    layer4_outputs(1870) <= not (a or b);
    layer4_outputs(1871) <= a and not b;
    layer4_outputs(1872) <= a;
    layer4_outputs(1873) <= a or b;
    layer4_outputs(1874) <= not (a or b);
    layer4_outputs(1875) <= a and b;
    layer4_outputs(1876) <= a;
    layer4_outputs(1877) <= 1'b0;
    layer4_outputs(1878) <= not a;
    layer4_outputs(1879) <= not (a xor b);
    layer4_outputs(1880) <= b;
    layer4_outputs(1881) <= not b;
    layer4_outputs(1882) <= not b;
    layer4_outputs(1883) <= not a or b;
    layer4_outputs(1884) <= not a or b;
    layer4_outputs(1885) <= not b;
    layer4_outputs(1886) <= b and not a;
    layer4_outputs(1887) <= a xor b;
    layer4_outputs(1888) <= a and b;
    layer4_outputs(1889) <= not (a xor b);
    layer4_outputs(1890) <= not a;
    layer4_outputs(1891) <= not b or a;
    layer4_outputs(1892) <= not b or a;
    layer4_outputs(1893) <= not (a and b);
    layer4_outputs(1894) <= a and b;
    layer4_outputs(1895) <= a or b;
    layer4_outputs(1896) <= a or b;
    layer4_outputs(1897) <= a and b;
    layer4_outputs(1898) <= not b or a;
    layer4_outputs(1899) <= not a;
    layer4_outputs(1900) <= a or b;
    layer4_outputs(1901) <= not a;
    layer4_outputs(1902) <= a xor b;
    layer4_outputs(1903) <= 1'b0;
    layer4_outputs(1904) <= not a;
    layer4_outputs(1905) <= not a;
    layer4_outputs(1906) <= a xor b;
    layer4_outputs(1907) <= not b;
    layer4_outputs(1908) <= a or b;
    layer4_outputs(1909) <= a xor b;
    layer4_outputs(1910) <= a and not b;
    layer4_outputs(1911) <= not b;
    layer4_outputs(1912) <= not b;
    layer4_outputs(1913) <= b;
    layer4_outputs(1914) <= a xor b;
    layer4_outputs(1915) <= not a;
    layer4_outputs(1916) <= not a or b;
    layer4_outputs(1917) <= not (a and b);
    layer4_outputs(1918) <= b and not a;
    layer4_outputs(1919) <= not (a and b);
    layer4_outputs(1920) <= a;
    layer4_outputs(1921) <= a and b;
    layer4_outputs(1922) <= a xor b;
    layer4_outputs(1923) <= not (a xor b);
    layer4_outputs(1924) <= not b or a;
    layer4_outputs(1925) <= a and b;
    layer4_outputs(1926) <= b and not a;
    layer4_outputs(1927) <= not b;
    layer4_outputs(1928) <= b and not a;
    layer4_outputs(1929) <= not (a xor b);
    layer4_outputs(1930) <= a xor b;
    layer4_outputs(1931) <= b;
    layer4_outputs(1932) <= b;
    layer4_outputs(1933) <= a and not b;
    layer4_outputs(1934) <= a;
    layer4_outputs(1935) <= a;
    layer4_outputs(1936) <= not b;
    layer4_outputs(1937) <= not b;
    layer4_outputs(1938) <= not b or a;
    layer4_outputs(1939) <= a;
    layer4_outputs(1940) <= not a;
    layer4_outputs(1941) <= b and not a;
    layer4_outputs(1942) <= not (a or b);
    layer4_outputs(1943) <= a;
    layer4_outputs(1944) <= not b;
    layer4_outputs(1945) <= a and b;
    layer4_outputs(1946) <= not (a xor b);
    layer4_outputs(1947) <= not (a xor b);
    layer4_outputs(1948) <= b and not a;
    layer4_outputs(1949) <= a;
    layer4_outputs(1950) <= a and not b;
    layer4_outputs(1951) <= not a;
    layer4_outputs(1952) <= a;
    layer4_outputs(1953) <= a xor b;
    layer4_outputs(1954) <= a;
    layer4_outputs(1955) <= a;
    layer4_outputs(1956) <= a xor b;
    layer4_outputs(1957) <= not (a xor b);
    layer4_outputs(1958) <= not (a xor b);
    layer4_outputs(1959) <= a xor b;
    layer4_outputs(1960) <= not (a and b);
    layer4_outputs(1961) <= a and b;
    layer4_outputs(1962) <= not (a xor b);
    layer4_outputs(1963) <= a xor b;
    layer4_outputs(1964) <= not a;
    layer4_outputs(1965) <= b;
    layer4_outputs(1966) <= a and not b;
    layer4_outputs(1967) <= not b;
    layer4_outputs(1968) <= not (a and b);
    layer4_outputs(1969) <= not a or b;
    layer4_outputs(1970) <= not (a or b);
    layer4_outputs(1971) <= not b or a;
    layer4_outputs(1972) <= not b;
    layer4_outputs(1973) <= not b;
    layer4_outputs(1974) <= a and not b;
    layer4_outputs(1975) <= a xor b;
    layer4_outputs(1976) <= not (a xor b);
    layer4_outputs(1977) <= not (a xor b);
    layer4_outputs(1978) <= not b;
    layer4_outputs(1979) <= not a or b;
    layer4_outputs(1980) <= a and b;
    layer4_outputs(1981) <= a xor b;
    layer4_outputs(1982) <= not a;
    layer4_outputs(1983) <= not a;
    layer4_outputs(1984) <= b and not a;
    layer4_outputs(1985) <= 1'b1;
    layer4_outputs(1986) <= b and not a;
    layer4_outputs(1987) <= not (a or b);
    layer4_outputs(1988) <= not b;
    layer4_outputs(1989) <= a and b;
    layer4_outputs(1990) <= b;
    layer4_outputs(1991) <= a and not b;
    layer4_outputs(1992) <= a and b;
    layer4_outputs(1993) <= not (a or b);
    layer4_outputs(1994) <= not b;
    layer4_outputs(1995) <= not a;
    layer4_outputs(1996) <= not (a and b);
    layer4_outputs(1997) <= a;
    layer4_outputs(1998) <= a and not b;
    layer4_outputs(1999) <= a and b;
    layer4_outputs(2000) <= not (a or b);
    layer4_outputs(2001) <= not b;
    layer4_outputs(2002) <= b;
    layer4_outputs(2003) <= b and not a;
    layer4_outputs(2004) <= b and not a;
    layer4_outputs(2005) <= a;
    layer4_outputs(2006) <= not a or b;
    layer4_outputs(2007) <= a xor b;
    layer4_outputs(2008) <= a and not b;
    layer4_outputs(2009) <= a xor b;
    layer4_outputs(2010) <= not (a xor b);
    layer4_outputs(2011) <= not a;
    layer4_outputs(2012) <= not b;
    layer4_outputs(2013) <= b;
    layer4_outputs(2014) <= not b;
    layer4_outputs(2015) <= a xor b;
    layer4_outputs(2016) <= not (a xor b);
    layer4_outputs(2017) <= a or b;
    layer4_outputs(2018) <= not a or b;
    layer4_outputs(2019) <= b;
    layer4_outputs(2020) <= a and b;
    layer4_outputs(2021) <= a and b;
    layer4_outputs(2022) <= a and b;
    layer4_outputs(2023) <= a xor b;
    layer4_outputs(2024) <= not (a or b);
    layer4_outputs(2025) <= b;
    layer4_outputs(2026) <= b;
    layer4_outputs(2027) <= not (a and b);
    layer4_outputs(2028) <= a and not b;
    layer4_outputs(2029) <= 1'b1;
    layer4_outputs(2030) <= not b;
    layer4_outputs(2031) <= not a or b;
    layer4_outputs(2032) <= not a;
    layer4_outputs(2033) <= a;
    layer4_outputs(2034) <= b;
    layer4_outputs(2035) <= a and not b;
    layer4_outputs(2036) <= b and not a;
    layer4_outputs(2037) <= not b;
    layer4_outputs(2038) <= a or b;
    layer4_outputs(2039) <= not (a xor b);
    layer4_outputs(2040) <= not a;
    layer4_outputs(2041) <= b and not a;
    layer4_outputs(2042) <= not (a xor b);
    layer4_outputs(2043) <= not (a or b);
    layer4_outputs(2044) <= not a or b;
    layer4_outputs(2045) <= b;
    layer4_outputs(2046) <= not a or b;
    layer4_outputs(2047) <= not a;
    layer4_outputs(2048) <= not b;
    layer4_outputs(2049) <= not b;
    layer4_outputs(2050) <= not b;
    layer4_outputs(2051) <= a;
    layer4_outputs(2052) <= a or b;
    layer4_outputs(2053) <= not b or a;
    layer4_outputs(2054) <= not (a and b);
    layer4_outputs(2055) <= not b or a;
    layer4_outputs(2056) <= a or b;
    layer4_outputs(2057) <= a and b;
    layer4_outputs(2058) <= a and b;
    layer4_outputs(2059) <= not (a and b);
    layer4_outputs(2060) <= a;
    layer4_outputs(2061) <= a xor b;
    layer4_outputs(2062) <= not b or a;
    layer4_outputs(2063) <= not b;
    layer4_outputs(2064) <= not a;
    layer4_outputs(2065) <= not (a xor b);
    layer4_outputs(2066) <= a and b;
    layer4_outputs(2067) <= a xor b;
    layer4_outputs(2068) <= not b or a;
    layer4_outputs(2069) <= 1'b1;
    layer4_outputs(2070) <= not a;
    layer4_outputs(2071) <= not b or a;
    layer4_outputs(2072) <= a or b;
    layer4_outputs(2073) <= a or b;
    layer4_outputs(2074) <= b;
    layer4_outputs(2075) <= a;
    layer4_outputs(2076) <= not b;
    layer4_outputs(2077) <= b;
    layer4_outputs(2078) <= not (a or b);
    layer4_outputs(2079) <= a xor b;
    layer4_outputs(2080) <= not b;
    layer4_outputs(2081) <= not b;
    layer4_outputs(2082) <= b;
    layer4_outputs(2083) <= a;
    layer4_outputs(2084) <= a;
    layer4_outputs(2085) <= a xor b;
    layer4_outputs(2086) <= a or b;
    layer4_outputs(2087) <= not a or b;
    layer4_outputs(2088) <= not a;
    layer4_outputs(2089) <= not a;
    layer4_outputs(2090) <= not (a and b);
    layer4_outputs(2091) <= a or b;
    layer4_outputs(2092) <= not (a xor b);
    layer4_outputs(2093) <= not b or a;
    layer4_outputs(2094) <= not b;
    layer4_outputs(2095) <= not (a or b);
    layer4_outputs(2096) <= not b;
    layer4_outputs(2097) <= b;
    layer4_outputs(2098) <= 1'b0;
    layer4_outputs(2099) <= not b;
    layer4_outputs(2100) <= b;
    layer4_outputs(2101) <= not a;
    layer4_outputs(2102) <= a;
    layer4_outputs(2103) <= a xor b;
    layer4_outputs(2104) <= not a or b;
    layer4_outputs(2105) <= b and not a;
    layer4_outputs(2106) <= not a;
    layer4_outputs(2107) <= b and not a;
    layer4_outputs(2108) <= a xor b;
    layer4_outputs(2109) <= a;
    layer4_outputs(2110) <= a xor b;
    layer4_outputs(2111) <= not b or a;
    layer4_outputs(2112) <= a or b;
    layer4_outputs(2113) <= not (a xor b);
    layer4_outputs(2114) <= not a;
    layer4_outputs(2115) <= not b or a;
    layer4_outputs(2116) <= not b;
    layer4_outputs(2117) <= b;
    layer4_outputs(2118) <= not (a and b);
    layer4_outputs(2119) <= not a;
    layer4_outputs(2120) <= a or b;
    layer4_outputs(2121) <= b;
    layer4_outputs(2122) <= a;
    layer4_outputs(2123) <= not b or a;
    layer4_outputs(2124) <= not (a xor b);
    layer4_outputs(2125) <= a or b;
    layer4_outputs(2126) <= not a;
    layer4_outputs(2127) <= not (a and b);
    layer4_outputs(2128) <= b and not a;
    layer4_outputs(2129) <= a or b;
    layer4_outputs(2130) <= a xor b;
    layer4_outputs(2131) <= a xor b;
    layer4_outputs(2132) <= b;
    layer4_outputs(2133) <= b and not a;
    layer4_outputs(2134) <= a;
    layer4_outputs(2135) <= b and not a;
    layer4_outputs(2136) <= not (a and b);
    layer4_outputs(2137) <= not b;
    layer4_outputs(2138) <= not a;
    layer4_outputs(2139) <= not b;
    layer4_outputs(2140) <= b;
    layer4_outputs(2141) <= a and not b;
    layer4_outputs(2142) <= b and not a;
    layer4_outputs(2143) <= a and b;
    layer4_outputs(2144) <= not a or b;
    layer4_outputs(2145) <= a and b;
    layer4_outputs(2146) <= a;
    layer4_outputs(2147) <= a xor b;
    layer4_outputs(2148) <= not b;
    layer4_outputs(2149) <= a and b;
    layer4_outputs(2150) <= not a;
    layer4_outputs(2151) <= not a;
    layer4_outputs(2152) <= not (a xor b);
    layer4_outputs(2153) <= b and not a;
    layer4_outputs(2154) <= b and not a;
    layer4_outputs(2155) <= a and b;
    layer4_outputs(2156) <= not b;
    layer4_outputs(2157) <= not (a or b);
    layer4_outputs(2158) <= not b;
    layer4_outputs(2159) <= not b;
    layer4_outputs(2160) <= b and not a;
    layer4_outputs(2161) <= not b;
    layer4_outputs(2162) <= a and b;
    layer4_outputs(2163) <= 1'b0;
    layer4_outputs(2164) <= a xor b;
    layer4_outputs(2165) <= a;
    layer4_outputs(2166) <= a;
    layer4_outputs(2167) <= a and b;
    layer4_outputs(2168) <= not (a or b);
    layer4_outputs(2169) <= a;
    layer4_outputs(2170) <= not (a xor b);
    layer4_outputs(2171) <= a;
    layer4_outputs(2172) <= a;
    layer4_outputs(2173) <= b;
    layer4_outputs(2174) <= not a or b;
    layer4_outputs(2175) <= not a or b;
    layer4_outputs(2176) <= not (a xor b);
    layer4_outputs(2177) <= not b;
    layer4_outputs(2178) <= not a;
    layer4_outputs(2179) <= not (a or b);
    layer4_outputs(2180) <= a xor b;
    layer4_outputs(2181) <= a or b;
    layer4_outputs(2182) <= not (a or b);
    layer4_outputs(2183) <= a xor b;
    layer4_outputs(2184) <= not (a or b);
    layer4_outputs(2185) <= not b;
    layer4_outputs(2186) <= a xor b;
    layer4_outputs(2187) <= not b or a;
    layer4_outputs(2188) <= a and b;
    layer4_outputs(2189) <= not a;
    layer4_outputs(2190) <= not a;
    layer4_outputs(2191) <= not (a xor b);
    layer4_outputs(2192) <= a and not b;
    layer4_outputs(2193) <= a;
    layer4_outputs(2194) <= b;
    layer4_outputs(2195) <= a and not b;
    layer4_outputs(2196) <= not b;
    layer4_outputs(2197) <= b;
    layer4_outputs(2198) <= not b;
    layer4_outputs(2199) <= not b;
    layer4_outputs(2200) <= a;
    layer4_outputs(2201) <= not (a xor b);
    layer4_outputs(2202) <= b;
    layer4_outputs(2203) <= not a;
    layer4_outputs(2204) <= a;
    layer4_outputs(2205) <= not a;
    layer4_outputs(2206) <= a;
    layer4_outputs(2207) <= b;
    layer4_outputs(2208) <= not (a xor b);
    layer4_outputs(2209) <= not (a xor b);
    layer4_outputs(2210) <= a xor b;
    layer4_outputs(2211) <= not (a xor b);
    layer4_outputs(2212) <= b and not a;
    layer4_outputs(2213) <= a and b;
    layer4_outputs(2214) <= not (a xor b);
    layer4_outputs(2215) <= not (a xor b);
    layer4_outputs(2216) <= a xor b;
    layer4_outputs(2217) <= not b;
    layer4_outputs(2218) <= not (a xor b);
    layer4_outputs(2219) <= a xor b;
    layer4_outputs(2220) <= a and not b;
    layer4_outputs(2221) <= not a;
    layer4_outputs(2222) <= a and not b;
    layer4_outputs(2223) <= not b;
    layer4_outputs(2224) <= a;
    layer4_outputs(2225) <= not (a xor b);
    layer4_outputs(2226) <= b;
    layer4_outputs(2227) <= not a;
    layer4_outputs(2228) <= not b;
    layer4_outputs(2229) <= b;
    layer4_outputs(2230) <= not b;
    layer4_outputs(2231) <= not (a and b);
    layer4_outputs(2232) <= not b;
    layer4_outputs(2233) <= not a or b;
    layer4_outputs(2234) <= not b;
    layer4_outputs(2235) <= b;
    layer4_outputs(2236) <= not b;
    layer4_outputs(2237) <= not a;
    layer4_outputs(2238) <= a;
    layer4_outputs(2239) <= not a;
    layer4_outputs(2240) <= a xor b;
    layer4_outputs(2241) <= a xor b;
    layer4_outputs(2242) <= a;
    layer4_outputs(2243) <= a;
    layer4_outputs(2244) <= not (a or b);
    layer4_outputs(2245) <= not b or a;
    layer4_outputs(2246) <= a xor b;
    layer4_outputs(2247) <= a or b;
    layer4_outputs(2248) <= b;
    layer4_outputs(2249) <= not (a and b);
    layer4_outputs(2250) <= a xor b;
    layer4_outputs(2251) <= not a or b;
    layer4_outputs(2252) <= not a or b;
    layer4_outputs(2253) <= a and not b;
    layer4_outputs(2254) <= not a;
    layer4_outputs(2255) <= b and not a;
    layer4_outputs(2256) <= not b;
    layer4_outputs(2257) <= a or b;
    layer4_outputs(2258) <= not (a and b);
    layer4_outputs(2259) <= not (a and b);
    layer4_outputs(2260) <= a xor b;
    layer4_outputs(2261) <= b;
    layer4_outputs(2262) <= not (a or b);
    layer4_outputs(2263) <= a xor b;
    layer4_outputs(2264) <= b;
    layer4_outputs(2265) <= not a or b;
    layer4_outputs(2266) <= a;
    layer4_outputs(2267) <= not a;
    layer4_outputs(2268) <= not a;
    layer4_outputs(2269) <= not b;
    layer4_outputs(2270) <= not b;
    layer4_outputs(2271) <= a and b;
    layer4_outputs(2272) <= a or b;
    layer4_outputs(2273) <= not (a xor b);
    layer4_outputs(2274) <= not b or a;
    layer4_outputs(2275) <= a and not b;
    layer4_outputs(2276) <= not a or b;
    layer4_outputs(2277) <= not b;
    layer4_outputs(2278) <= not (a xor b);
    layer4_outputs(2279) <= not b;
    layer4_outputs(2280) <= a;
    layer4_outputs(2281) <= a xor b;
    layer4_outputs(2282) <= not b;
    layer4_outputs(2283) <= not b or a;
    layer4_outputs(2284) <= a;
    layer4_outputs(2285) <= a xor b;
    layer4_outputs(2286) <= b;
    layer4_outputs(2287) <= b and not a;
    layer4_outputs(2288) <= not a;
    layer4_outputs(2289) <= not (a xor b);
    layer4_outputs(2290) <= a xor b;
    layer4_outputs(2291) <= a or b;
    layer4_outputs(2292) <= not a or b;
    layer4_outputs(2293) <= b;
    layer4_outputs(2294) <= b and not a;
    layer4_outputs(2295) <= a and b;
    layer4_outputs(2296) <= not a or b;
    layer4_outputs(2297) <= b;
    layer4_outputs(2298) <= not b;
    layer4_outputs(2299) <= not a;
    layer4_outputs(2300) <= not a or b;
    layer4_outputs(2301) <= not b;
    layer4_outputs(2302) <= not (a xor b);
    layer4_outputs(2303) <= not a or b;
    layer4_outputs(2304) <= a and not b;
    layer4_outputs(2305) <= not b or a;
    layer4_outputs(2306) <= not b;
    layer4_outputs(2307) <= b;
    layer4_outputs(2308) <= not (a or b);
    layer4_outputs(2309) <= a xor b;
    layer4_outputs(2310) <= not a or b;
    layer4_outputs(2311) <= not (a and b);
    layer4_outputs(2312) <= b;
    layer4_outputs(2313) <= a xor b;
    layer4_outputs(2314) <= a;
    layer4_outputs(2315) <= not a;
    layer4_outputs(2316) <= a;
    layer4_outputs(2317) <= a;
    layer4_outputs(2318) <= not b;
    layer4_outputs(2319) <= not a;
    layer4_outputs(2320) <= a and not b;
    layer4_outputs(2321) <= not (a xor b);
    layer4_outputs(2322) <= a;
    layer4_outputs(2323) <= not (a or b);
    layer4_outputs(2324) <= a and not b;
    layer4_outputs(2325) <= not b;
    layer4_outputs(2326) <= b;
    layer4_outputs(2327) <= not a or b;
    layer4_outputs(2328) <= a xor b;
    layer4_outputs(2329) <= a;
    layer4_outputs(2330) <= not a;
    layer4_outputs(2331) <= not (a xor b);
    layer4_outputs(2332) <= not b;
    layer4_outputs(2333) <= not a;
    layer4_outputs(2334) <= b;
    layer4_outputs(2335) <= not (a xor b);
    layer4_outputs(2336) <= b;
    layer4_outputs(2337) <= not (a and b);
    layer4_outputs(2338) <= a and not b;
    layer4_outputs(2339) <= b;
    layer4_outputs(2340) <= not b or a;
    layer4_outputs(2341) <= b;
    layer4_outputs(2342) <= not b;
    layer4_outputs(2343) <= b and not a;
    layer4_outputs(2344) <= not a;
    layer4_outputs(2345) <= a or b;
    layer4_outputs(2346) <= a and b;
    layer4_outputs(2347) <= not (a xor b);
    layer4_outputs(2348) <= not (a and b);
    layer4_outputs(2349) <= a and b;
    layer4_outputs(2350) <= not (a and b);
    layer4_outputs(2351) <= not b;
    layer4_outputs(2352) <= a;
    layer4_outputs(2353) <= a and b;
    layer4_outputs(2354) <= a and b;
    layer4_outputs(2355) <= a or b;
    layer4_outputs(2356) <= not a;
    layer4_outputs(2357) <= b;
    layer4_outputs(2358) <= not a;
    layer4_outputs(2359) <= a;
    layer4_outputs(2360) <= a or b;
    layer4_outputs(2361) <= not (a or b);
    layer4_outputs(2362) <= not b;
    layer4_outputs(2363) <= not b;
    layer4_outputs(2364) <= not (a or b);
    layer4_outputs(2365) <= a;
    layer4_outputs(2366) <= b;
    layer4_outputs(2367) <= a and b;
    layer4_outputs(2368) <= a;
    layer4_outputs(2369) <= not a or b;
    layer4_outputs(2370) <= a xor b;
    layer4_outputs(2371) <= not (a and b);
    layer4_outputs(2372) <= a;
    layer4_outputs(2373) <= not (a or b);
    layer4_outputs(2374) <= not (a or b);
    layer4_outputs(2375) <= b;
    layer4_outputs(2376) <= b;
    layer4_outputs(2377) <= b;
    layer4_outputs(2378) <= not (a xor b);
    layer4_outputs(2379) <= a and not b;
    layer4_outputs(2380) <= not a or b;
    layer4_outputs(2381) <= not (a and b);
    layer4_outputs(2382) <= a xor b;
    layer4_outputs(2383) <= a xor b;
    layer4_outputs(2384) <= not a or b;
    layer4_outputs(2385) <= not a;
    layer4_outputs(2386) <= a;
    layer4_outputs(2387) <= a or b;
    layer4_outputs(2388) <= not (a and b);
    layer4_outputs(2389) <= not (a xor b);
    layer4_outputs(2390) <= b and not a;
    layer4_outputs(2391) <= a;
    layer4_outputs(2392) <= a and not b;
    layer4_outputs(2393) <= not b;
    layer4_outputs(2394) <= b;
    layer4_outputs(2395) <= b;
    layer4_outputs(2396) <= a;
    layer4_outputs(2397) <= not (a xor b);
    layer4_outputs(2398) <= a and not b;
    layer4_outputs(2399) <= not a or b;
    layer4_outputs(2400) <= not a or b;
    layer4_outputs(2401) <= not a or b;
    layer4_outputs(2402) <= a or b;
    layer4_outputs(2403) <= a and b;
    layer4_outputs(2404) <= not (a and b);
    layer4_outputs(2405) <= a xor b;
    layer4_outputs(2406) <= not (a xor b);
    layer4_outputs(2407) <= not (a or b);
    layer4_outputs(2408) <= b;
    layer4_outputs(2409) <= b;
    layer4_outputs(2410) <= b;
    layer4_outputs(2411) <= not b;
    layer4_outputs(2412) <= not (a xor b);
    layer4_outputs(2413) <= not b;
    layer4_outputs(2414) <= not (a and b);
    layer4_outputs(2415) <= a or b;
    layer4_outputs(2416) <= not (a and b);
    layer4_outputs(2417) <= a;
    layer4_outputs(2418) <= b;
    layer4_outputs(2419) <= a or b;
    layer4_outputs(2420) <= a and b;
    layer4_outputs(2421) <= a and b;
    layer4_outputs(2422) <= a xor b;
    layer4_outputs(2423) <= not b or a;
    layer4_outputs(2424) <= not a;
    layer4_outputs(2425) <= not b;
    layer4_outputs(2426) <= not a;
    layer4_outputs(2427) <= not a;
    layer4_outputs(2428) <= a;
    layer4_outputs(2429) <= b and not a;
    layer4_outputs(2430) <= a or b;
    layer4_outputs(2431) <= b and not a;
    layer4_outputs(2432) <= not b;
    layer4_outputs(2433) <= a;
    layer4_outputs(2434) <= b;
    layer4_outputs(2435) <= b and not a;
    layer4_outputs(2436) <= not (a and b);
    layer4_outputs(2437) <= a or b;
    layer4_outputs(2438) <= not (a and b);
    layer4_outputs(2439) <= a and not b;
    layer4_outputs(2440) <= a;
    layer4_outputs(2441) <= not (a xor b);
    layer4_outputs(2442) <= not b or a;
    layer4_outputs(2443) <= not a or b;
    layer4_outputs(2444) <= a and b;
    layer4_outputs(2445) <= a;
    layer4_outputs(2446) <= b;
    layer4_outputs(2447) <= a;
    layer4_outputs(2448) <= a;
    layer4_outputs(2449) <= not (a xor b);
    layer4_outputs(2450) <= not a;
    layer4_outputs(2451) <= not (a xor b);
    layer4_outputs(2452) <= not a;
    layer4_outputs(2453) <= a xor b;
    layer4_outputs(2454) <= not a or b;
    layer4_outputs(2455) <= a and not b;
    layer4_outputs(2456) <= a and b;
    layer4_outputs(2457) <= a xor b;
    layer4_outputs(2458) <= b and not a;
    layer4_outputs(2459) <= not b or a;
    layer4_outputs(2460) <= a or b;
    layer4_outputs(2461) <= not a or b;
    layer4_outputs(2462) <= not b;
    layer4_outputs(2463) <= not (a and b);
    layer4_outputs(2464) <= not a;
    layer4_outputs(2465) <= a xor b;
    layer4_outputs(2466) <= b and not a;
    layer4_outputs(2467) <= not (a xor b);
    layer4_outputs(2468) <= a and b;
    layer4_outputs(2469) <= a;
    layer4_outputs(2470) <= not (a xor b);
    layer4_outputs(2471) <= b and not a;
    layer4_outputs(2472) <= not (a xor b);
    layer4_outputs(2473) <= not b;
    layer4_outputs(2474) <= a;
    layer4_outputs(2475) <= not b or a;
    layer4_outputs(2476) <= not b;
    layer4_outputs(2477) <= b;
    layer4_outputs(2478) <= a xor b;
    layer4_outputs(2479) <= a and b;
    layer4_outputs(2480) <= a and b;
    layer4_outputs(2481) <= not a;
    layer4_outputs(2482) <= a xor b;
    layer4_outputs(2483) <= a;
    layer4_outputs(2484) <= not b;
    layer4_outputs(2485) <= not b or a;
    layer4_outputs(2486) <= not a;
    layer4_outputs(2487) <= a or b;
    layer4_outputs(2488) <= b and not a;
    layer4_outputs(2489) <= b;
    layer4_outputs(2490) <= a;
    layer4_outputs(2491) <= a xor b;
    layer4_outputs(2492) <= a xor b;
    layer4_outputs(2493) <= not a;
    layer4_outputs(2494) <= a;
    layer4_outputs(2495) <= not a or b;
    layer4_outputs(2496) <= not b;
    layer4_outputs(2497) <= a and not b;
    layer4_outputs(2498) <= not (a or b);
    layer4_outputs(2499) <= not a;
    layer4_outputs(2500) <= 1'b0;
    layer4_outputs(2501) <= not b;
    layer4_outputs(2502) <= not a;
    layer4_outputs(2503) <= b;
    layer4_outputs(2504) <= not (a xor b);
    layer4_outputs(2505) <= not b;
    layer4_outputs(2506) <= not b or a;
    layer4_outputs(2507) <= a;
    layer4_outputs(2508) <= a or b;
    layer4_outputs(2509) <= a and b;
    layer4_outputs(2510) <= not (a xor b);
    layer4_outputs(2511) <= not a;
    layer4_outputs(2512) <= not a;
    layer4_outputs(2513) <= b;
    layer4_outputs(2514) <= not a;
    layer4_outputs(2515) <= a;
    layer4_outputs(2516) <= not (a xor b);
    layer4_outputs(2517) <= not b or a;
    layer4_outputs(2518) <= b and not a;
    layer4_outputs(2519) <= b;
    layer4_outputs(2520) <= b;
    layer4_outputs(2521) <= not (a xor b);
    layer4_outputs(2522) <= a xor b;
    layer4_outputs(2523) <= b;
    layer4_outputs(2524) <= a;
    layer4_outputs(2525) <= a or b;
    layer4_outputs(2526) <= a or b;
    layer4_outputs(2527) <= not (a xor b);
    layer4_outputs(2528) <= not b;
    layer4_outputs(2529) <= not a or b;
    layer4_outputs(2530) <= not a;
    layer4_outputs(2531) <= a;
    layer4_outputs(2532) <= not a or b;
    layer4_outputs(2533) <= b;
    layer4_outputs(2534) <= a and not b;
    layer4_outputs(2535) <= b;
    layer4_outputs(2536) <= a;
    layer4_outputs(2537) <= not (a or b);
    layer4_outputs(2538) <= a xor b;
    layer4_outputs(2539) <= a;
    layer4_outputs(2540) <= not (a and b);
    layer4_outputs(2541) <= b;
    layer4_outputs(2542) <= not (a and b);
    layer4_outputs(2543) <= a;
    layer4_outputs(2544) <= b;
    layer4_outputs(2545) <= a and not b;
    layer4_outputs(2546) <= not b;
    layer4_outputs(2547) <= not (a or b);
    layer4_outputs(2548) <= a;
    layer4_outputs(2549) <= not a;
    layer4_outputs(2550) <= not (a xor b);
    layer4_outputs(2551) <= not b or a;
    layer4_outputs(2552) <= a;
    layer4_outputs(2553) <= not (a and b);
    layer4_outputs(2554) <= b;
    layer4_outputs(2555) <= not a or b;
    layer4_outputs(2556) <= b;
    layer4_outputs(2557) <= b and not a;
    layer4_outputs(2558) <= a;
    layer4_outputs(2559) <= not (a xor b);
    layer4_outputs(2560) <= not (a xor b);
    layer4_outputs(2561) <= a and not b;
    layer4_outputs(2562) <= not b;
    layer4_outputs(2563) <= not a;
    layer4_outputs(2564) <= not b;
    layer4_outputs(2565) <= b;
    layer4_outputs(2566) <= not b;
    layer4_outputs(2567) <= not (a and b);
    layer4_outputs(2568) <= a or b;
    layer4_outputs(2569) <= not b;
    layer4_outputs(2570) <= not b or a;
    layer4_outputs(2571) <= not a;
    layer4_outputs(2572) <= not (a or b);
    layer4_outputs(2573) <= not b;
    layer4_outputs(2574) <= not (a xor b);
    layer4_outputs(2575) <= a and b;
    layer4_outputs(2576) <= not b;
    layer4_outputs(2577) <= not b;
    layer4_outputs(2578) <= b;
    layer4_outputs(2579) <= not a;
    layer4_outputs(2580) <= not b;
    layer4_outputs(2581) <= not a or b;
    layer4_outputs(2582) <= a xor b;
    layer4_outputs(2583) <= not a;
    layer4_outputs(2584) <= not b;
    layer4_outputs(2585) <= not a;
    layer4_outputs(2586) <= a or b;
    layer4_outputs(2587) <= b and not a;
    layer4_outputs(2588) <= b;
    layer4_outputs(2589) <= b;
    layer4_outputs(2590) <= not b;
    layer4_outputs(2591) <= not b or a;
    layer4_outputs(2592) <= not (a and b);
    layer4_outputs(2593) <= not (a or b);
    layer4_outputs(2594) <= a;
    layer4_outputs(2595) <= b and not a;
    layer4_outputs(2596) <= not (a xor b);
    layer4_outputs(2597) <= a or b;
    layer4_outputs(2598) <= a and not b;
    layer4_outputs(2599) <= b and not a;
    layer4_outputs(2600) <= a;
    layer4_outputs(2601) <= a and b;
    layer4_outputs(2602) <= not (a xor b);
    layer4_outputs(2603) <= not (a and b);
    layer4_outputs(2604) <= not b;
    layer4_outputs(2605) <= not b or a;
    layer4_outputs(2606) <= not b;
    layer4_outputs(2607) <= b and not a;
    layer4_outputs(2608) <= not a or b;
    layer4_outputs(2609) <= a and not b;
    layer4_outputs(2610) <= b;
    layer4_outputs(2611) <= a;
    layer4_outputs(2612) <= not (a xor b);
    layer4_outputs(2613) <= 1'b1;
    layer4_outputs(2614) <= not (a or b);
    layer4_outputs(2615) <= b;
    layer4_outputs(2616) <= a;
    layer4_outputs(2617) <= not (a or b);
    layer4_outputs(2618) <= not b;
    layer4_outputs(2619) <= a or b;
    layer4_outputs(2620) <= not a;
    layer4_outputs(2621) <= not b;
    layer4_outputs(2622) <= not (a xor b);
    layer4_outputs(2623) <= b and not a;
    layer4_outputs(2624) <= a and not b;
    layer4_outputs(2625) <= not b;
    layer4_outputs(2626) <= a or b;
    layer4_outputs(2627) <= not a;
    layer4_outputs(2628) <= a;
    layer4_outputs(2629) <= a or b;
    layer4_outputs(2630) <= not (a xor b);
    layer4_outputs(2631) <= a;
    layer4_outputs(2632) <= not b;
    layer4_outputs(2633) <= not (a and b);
    layer4_outputs(2634) <= not a;
    layer4_outputs(2635) <= not (a xor b);
    layer4_outputs(2636) <= not a;
    layer4_outputs(2637) <= a and not b;
    layer4_outputs(2638) <= not b;
    layer4_outputs(2639) <= a xor b;
    layer4_outputs(2640) <= not (a xor b);
    layer4_outputs(2641) <= a or b;
    layer4_outputs(2642) <= not a;
    layer4_outputs(2643) <= not b;
    layer4_outputs(2644) <= a;
    layer4_outputs(2645) <= not b;
    layer4_outputs(2646) <= a and b;
    layer4_outputs(2647) <= not (a or b);
    layer4_outputs(2648) <= a;
    layer4_outputs(2649) <= a;
    layer4_outputs(2650) <= b;
    layer4_outputs(2651) <= a;
    layer4_outputs(2652) <= not b or a;
    layer4_outputs(2653) <= a;
    layer4_outputs(2654) <= b;
    layer4_outputs(2655) <= not a;
    layer4_outputs(2656) <= not b;
    layer4_outputs(2657) <= b;
    layer4_outputs(2658) <= not (a and b);
    layer4_outputs(2659) <= a xor b;
    layer4_outputs(2660) <= a;
    layer4_outputs(2661) <= not (a xor b);
    layer4_outputs(2662) <= not (a and b);
    layer4_outputs(2663) <= a or b;
    layer4_outputs(2664) <= not a;
    layer4_outputs(2665) <= not a;
    layer4_outputs(2666) <= not a or b;
    layer4_outputs(2667) <= not b;
    layer4_outputs(2668) <= b;
    layer4_outputs(2669) <= not b;
    layer4_outputs(2670) <= not b;
    layer4_outputs(2671) <= not b;
    layer4_outputs(2672) <= a and b;
    layer4_outputs(2673) <= a;
    layer4_outputs(2674) <= not (a xor b);
    layer4_outputs(2675) <= not a;
    layer4_outputs(2676) <= not a;
    layer4_outputs(2677) <= not b;
    layer4_outputs(2678) <= a;
    layer4_outputs(2679) <= not (a xor b);
    layer4_outputs(2680) <= b;
    layer4_outputs(2681) <= not b;
    layer4_outputs(2682) <= a;
    layer4_outputs(2683) <= not b;
    layer4_outputs(2684) <= a;
    layer4_outputs(2685) <= b;
    layer4_outputs(2686) <= a;
    layer4_outputs(2687) <= not (a and b);
    layer4_outputs(2688) <= not (a or b);
    layer4_outputs(2689) <= b;
    layer4_outputs(2690) <= not (a and b);
    layer4_outputs(2691) <= not (a and b);
    layer4_outputs(2692) <= not a;
    layer4_outputs(2693) <= b;
    layer4_outputs(2694) <= b;
    layer4_outputs(2695) <= not a;
    layer4_outputs(2696) <= a;
    layer4_outputs(2697) <= not (a and b);
    layer4_outputs(2698) <= not (a xor b);
    layer4_outputs(2699) <= a;
    layer4_outputs(2700) <= a;
    layer4_outputs(2701) <= not a or b;
    layer4_outputs(2702) <= a or b;
    layer4_outputs(2703) <= not (a or b);
    layer4_outputs(2704) <= not a;
    layer4_outputs(2705) <= not (a xor b);
    layer4_outputs(2706) <= not a or b;
    layer4_outputs(2707) <= a or b;
    layer4_outputs(2708) <= a or b;
    layer4_outputs(2709) <= not (a xor b);
    layer4_outputs(2710) <= not (a xor b);
    layer4_outputs(2711) <= not a or b;
    layer4_outputs(2712) <= a and b;
    layer4_outputs(2713) <= not b;
    layer4_outputs(2714) <= not (a or b);
    layer4_outputs(2715) <= a;
    layer4_outputs(2716) <= a;
    layer4_outputs(2717) <= b;
    layer4_outputs(2718) <= b;
    layer4_outputs(2719) <= not a;
    layer4_outputs(2720) <= not (a and b);
    layer4_outputs(2721) <= not b or a;
    layer4_outputs(2722) <= not b;
    layer4_outputs(2723) <= not a or b;
    layer4_outputs(2724) <= not a or b;
    layer4_outputs(2725) <= b;
    layer4_outputs(2726) <= a or b;
    layer4_outputs(2727) <= not a or b;
    layer4_outputs(2728) <= a or b;
    layer4_outputs(2729) <= not (a or b);
    layer4_outputs(2730) <= a and not b;
    layer4_outputs(2731) <= not b;
    layer4_outputs(2732) <= a;
    layer4_outputs(2733) <= a;
    layer4_outputs(2734) <= not (a xor b);
    layer4_outputs(2735) <= not b;
    layer4_outputs(2736) <= not (a xor b);
    layer4_outputs(2737) <= a xor b;
    layer4_outputs(2738) <= not a;
    layer4_outputs(2739) <= not (a xor b);
    layer4_outputs(2740) <= a;
    layer4_outputs(2741) <= a and not b;
    layer4_outputs(2742) <= a xor b;
    layer4_outputs(2743) <= b;
    layer4_outputs(2744) <= not b;
    layer4_outputs(2745) <= b;
    layer4_outputs(2746) <= a and b;
    layer4_outputs(2747) <= not (a and b);
    layer4_outputs(2748) <= a xor b;
    layer4_outputs(2749) <= not b;
    layer4_outputs(2750) <= b;
    layer4_outputs(2751) <= a or b;
    layer4_outputs(2752) <= b;
    layer4_outputs(2753) <= not b;
    layer4_outputs(2754) <= a and b;
    layer4_outputs(2755) <= not (a xor b);
    layer4_outputs(2756) <= b and not a;
    layer4_outputs(2757) <= not a;
    layer4_outputs(2758) <= b;
    layer4_outputs(2759) <= b and not a;
    layer4_outputs(2760) <= not (a and b);
    layer4_outputs(2761) <= not b;
    layer4_outputs(2762) <= a and b;
    layer4_outputs(2763) <= not b;
    layer4_outputs(2764) <= not b;
    layer4_outputs(2765) <= a xor b;
    layer4_outputs(2766) <= not a;
    layer4_outputs(2767) <= not (a xor b);
    layer4_outputs(2768) <= not a;
    layer4_outputs(2769) <= not (a xor b);
    layer4_outputs(2770) <= a;
    layer4_outputs(2771) <= b;
    layer4_outputs(2772) <= not a or b;
    layer4_outputs(2773) <= a;
    layer4_outputs(2774) <= b and not a;
    layer4_outputs(2775) <= not (a xor b);
    layer4_outputs(2776) <= 1'b0;
    layer4_outputs(2777) <= a xor b;
    layer4_outputs(2778) <= a or b;
    layer4_outputs(2779) <= b;
    layer4_outputs(2780) <= not a;
    layer4_outputs(2781) <= b;
    layer4_outputs(2782) <= not (a and b);
    layer4_outputs(2783) <= not a or b;
    layer4_outputs(2784) <= a;
    layer4_outputs(2785) <= not (a and b);
    layer4_outputs(2786) <= not a;
    layer4_outputs(2787) <= a or b;
    layer4_outputs(2788) <= a xor b;
    layer4_outputs(2789) <= not a or b;
    layer4_outputs(2790) <= not a;
    layer4_outputs(2791) <= a and b;
    layer4_outputs(2792) <= b;
    layer4_outputs(2793) <= not (a xor b);
    layer4_outputs(2794) <= b;
    layer4_outputs(2795) <= not b;
    layer4_outputs(2796) <= not a;
    layer4_outputs(2797) <= a xor b;
    layer4_outputs(2798) <= not a;
    layer4_outputs(2799) <= not a;
    layer4_outputs(2800) <= a;
    layer4_outputs(2801) <= not (a or b);
    layer4_outputs(2802) <= not (a and b);
    layer4_outputs(2803) <= not a;
    layer4_outputs(2804) <= not (a xor b);
    layer4_outputs(2805) <= not b;
    layer4_outputs(2806) <= b;
    layer4_outputs(2807) <= not (a and b);
    layer4_outputs(2808) <= not (a xor b);
    layer4_outputs(2809) <= not a;
    layer4_outputs(2810) <= a;
    layer4_outputs(2811) <= not a;
    layer4_outputs(2812) <= not a or b;
    layer4_outputs(2813) <= b;
    layer4_outputs(2814) <= a or b;
    layer4_outputs(2815) <= a xor b;
    layer4_outputs(2816) <= not a;
    layer4_outputs(2817) <= not b or a;
    layer4_outputs(2818) <= not (a and b);
    layer4_outputs(2819) <= not b;
    layer4_outputs(2820) <= not (a and b);
    layer4_outputs(2821) <= not b;
    layer4_outputs(2822) <= not (a or b);
    layer4_outputs(2823) <= a;
    layer4_outputs(2824) <= a;
    layer4_outputs(2825) <= a;
    layer4_outputs(2826) <= a;
    layer4_outputs(2827) <= not (a or b);
    layer4_outputs(2828) <= a;
    layer4_outputs(2829) <= not b or a;
    layer4_outputs(2830) <= b;
    layer4_outputs(2831) <= not a;
    layer4_outputs(2832) <= b;
    layer4_outputs(2833) <= not a;
    layer4_outputs(2834) <= not (a xor b);
    layer4_outputs(2835) <= not a or b;
    layer4_outputs(2836) <= a xor b;
    layer4_outputs(2837) <= a and not b;
    layer4_outputs(2838) <= not (a xor b);
    layer4_outputs(2839) <= b;
    layer4_outputs(2840) <= not (a xor b);
    layer4_outputs(2841) <= b;
    layer4_outputs(2842) <= not a;
    layer4_outputs(2843) <= not a or b;
    layer4_outputs(2844) <= not (a or b);
    layer4_outputs(2845) <= not a;
    layer4_outputs(2846) <= not a;
    layer4_outputs(2847) <= not b or a;
    layer4_outputs(2848) <= b;
    layer4_outputs(2849) <= not a or b;
    layer4_outputs(2850) <= not (a or b);
    layer4_outputs(2851) <= not (a and b);
    layer4_outputs(2852) <= not b;
    layer4_outputs(2853) <= a or b;
    layer4_outputs(2854) <= a or b;
    layer4_outputs(2855) <= not b;
    layer4_outputs(2856) <= a xor b;
    layer4_outputs(2857) <= not b or a;
    layer4_outputs(2858) <= a;
    layer4_outputs(2859) <= not b or a;
    layer4_outputs(2860) <= not b;
    layer4_outputs(2861) <= a and not b;
    layer4_outputs(2862) <= b;
    layer4_outputs(2863) <= b;
    layer4_outputs(2864) <= a and not b;
    layer4_outputs(2865) <= a xor b;
    layer4_outputs(2866) <= not a;
    layer4_outputs(2867) <= not b or a;
    layer4_outputs(2868) <= not b;
    layer4_outputs(2869) <= a xor b;
    layer4_outputs(2870) <= b and not a;
    layer4_outputs(2871) <= not a;
    layer4_outputs(2872) <= a;
    layer4_outputs(2873) <= a xor b;
    layer4_outputs(2874) <= b and not a;
    layer4_outputs(2875) <= not b;
    layer4_outputs(2876) <= not (a or b);
    layer4_outputs(2877) <= b;
    layer4_outputs(2878) <= a;
    layer4_outputs(2879) <= not b or a;
    layer4_outputs(2880) <= a;
    layer4_outputs(2881) <= not b;
    layer4_outputs(2882) <= b;
    layer4_outputs(2883) <= not b;
    layer4_outputs(2884) <= not b or a;
    layer4_outputs(2885) <= 1'b0;
    layer4_outputs(2886) <= not b;
    layer4_outputs(2887) <= not (a xor b);
    layer4_outputs(2888) <= not b;
    layer4_outputs(2889) <= a or b;
    layer4_outputs(2890) <= not a;
    layer4_outputs(2891) <= not b or a;
    layer4_outputs(2892) <= not a;
    layer4_outputs(2893) <= not (a xor b);
    layer4_outputs(2894) <= not (a and b);
    layer4_outputs(2895) <= not (a xor b);
    layer4_outputs(2896) <= a xor b;
    layer4_outputs(2897) <= not (a xor b);
    layer4_outputs(2898) <= not b or a;
    layer4_outputs(2899) <= b;
    layer4_outputs(2900) <= not (a and b);
    layer4_outputs(2901) <= a;
    layer4_outputs(2902) <= not b;
    layer4_outputs(2903) <= a;
    layer4_outputs(2904) <= not (a and b);
    layer4_outputs(2905) <= b;
    layer4_outputs(2906) <= b;
    layer4_outputs(2907) <= b and not a;
    layer4_outputs(2908) <= a;
    layer4_outputs(2909) <= b;
    layer4_outputs(2910) <= a;
    layer4_outputs(2911) <= not a;
    layer4_outputs(2912) <= a xor b;
    layer4_outputs(2913) <= a;
    layer4_outputs(2914) <= a xor b;
    layer4_outputs(2915) <= not (a xor b);
    layer4_outputs(2916) <= not b;
    layer4_outputs(2917) <= a;
    layer4_outputs(2918) <= b;
    layer4_outputs(2919) <= b;
    layer4_outputs(2920) <= b;
    layer4_outputs(2921) <= not a;
    layer4_outputs(2922) <= a xor b;
    layer4_outputs(2923) <= not a or b;
    layer4_outputs(2924) <= not b;
    layer4_outputs(2925) <= not (a xor b);
    layer4_outputs(2926) <= not b;
    layer4_outputs(2927) <= b;
    layer4_outputs(2928) <= a xor b;
    layer4_outputs(2929) <= not (a or b);
    layer4_outputs(2930) <= a and b;
    layer4_outputs(2931) <= b;
    layer4_outputs(2932) <= not a;
    layer4_outputs(2933) <= not (a xor b);
    layer4_outputs(2934) <= not b or a;
    layer4_outputs(2935) <= b;
    layer4_outputs(2936) <= a and not b;
    layer4_outputs(2937) <= not b;
    layer4_outputs(2938) <= not (a or b);
    layer4_outputs(2939) <= b;
    layer4_outputs(2940) <= b and not a;
    layer4_outputs(2941) <= b;
    layer4_outputs(2942) <= not b;
    layer4_outputs(2943) <= b and not a;
    layer4_outputs(2944) <= not b or a;
    layer4_outputs(2945) <= not (a or b);
    layer4_outputs(2946) <= a or b;
    layer4_outputs(2947) <= a and not b;
    layer4_outputs(2948) <= a xor b;
    layer4_outputs(2949) <= b and not a;
    layer4_outputs(2950) <= not a;
    layer4_outputs(2951) <= not a;
    layer4_outputs(2952) <= a xor b;
    layer4_outputs(2953) <= a and not b;
    layer4_outputs(2954) <= a or b;
    layer4_outputs(2955) <= a and not b;
    layer4_outputs(2956) <= not (a xor b);
    layer4_outputs(2957) <= b and not a;
    layer4_outputs(2958) <= a xor b;
    layer4_outputs(2959) <= not (a and b);
    layer4_outputs(2960) <= not b or a;
    layer4_outputs(2961) <= not a or b;
    layer4_outputs(2962) <= a;
    layer4_outputs(2963) <= not a;
    layer4_outputs(2964) <= a;
    layer4_outputs(2965) <= a or b;
    layer4_outputs(2966) <= not b or a;
    layer4_outputs(2967) <= b;
    layer4_outputs(2968) <= a and b;
    layer4_outputs(2969) <= not a or b;
    layer4_outputs(2970) <= a;
    layer4_outputs(2971) <= a and b;
    layer4_outputs(2972) <= not a or b;
    layer4_outputs(2973) <= not b;
    layer4_outputs(2974) <= a;
    layer4_outputs(2975) <= not b or a;
    layer4_outputs(2976) <= not (a or b);
    layer4_outputs(2977) <= not a;
    layer4_outputs(2978) <= not (a or b);
    layer4_outputs(2979) <= b and not a;
    layer4_outputs(2980) <= not a or b;
    layer4_outputs(2981) <= not (a xor b);
    layer4_outputs(2982) <= a;
    layer4_outputs(2983) <= a and b;
    layer4_outputs(2984) <= b;
    layer4_outputs(2985) <= a xor b;
    layer4_outputs(2986) <= b;
    layer4_outputs(2987) <= not (a or b);
    layer4_outputs(2988) <= not (a xor b);
    layer4_outputs(2989) <= not b or a;
    layer4_outputs(2990) <= a and not b;
    layer4_outputs(2991) <= b;
    layer4_outputs(2992) <= b and not a;
    layer4_outputs(2993) <= b;
    layer4_outputs(2994) <= b;
    layer4_outputs(2995) <= not b or a;
    layer4_outputs(2996) <= not (a xor b);
    layer4_outputs(2997) <= b and not a;
    layer4_outputs(2998) <= not a;
    layer4_outputs(2999) <= b and not a;
    layer4_outputs(3000) <= a and b;
    layer4_outputs(3001) <= a;
    layer4_outputs(3002) <= a xor b;
    layer4_outputs(3003) <= b and not a;
    layer4_outputs(3004) <= a;
    layer4_outputs(3005) <= a and b;
    layer4_outputs(3006) <= b;
    layer4_outputs(3007) <= a xor b;
    layer4_outputs(3008) <= not a or b;
    layer4_outputs(3009) <= not b;
    layer4_outputs(3010) <= not (a and b);
    layer4_outputs(3011) <= a xor b;
    layer4_outputs(3012) <= not b or a;
    layer4_outputs(3013) <= not a or b;
    layer4_outputs(3014) <= b and not a;
    layer4_outputs(3015) <= not b;
    layer4_outputs(3016) <= not (a or b);
    layer4_outputs(3017) <= b;
    layer4_outputs(3018) <= a or b;
    layer4_outputs(3019) <= not a;
    layer4_outputs(3020) <= not a;
    layer4_outputs(3021) <= not b;
    layer4_outputs(3022) <= 1'b1;
    layer4_outputs(3023) <= a;
    layer4_outputs(3024) <= not b;
    layer4_outputs(3025) <= a;
    layer4_outputs(3026) <= a and b;
    layer4_outputs(3027) <= a or b;
    layer4_outputs(3028) <= not (a or b);
    layer4_outputs(3029) <= b;
    layer4_outputs(3030) <= b and not a;
    layer4_outputs(3031) <= not b;
    layer4_outputs(3032) <= b;
    layer4_outputs(3033) <= not (a or b);
    layer4_outputs(3034) <= a;
    layer4_outputs(3035) <= a;
    layer4_outputs(3036) <= not b;
    layer4_outputs(3037) <= a xor b;
    layer4_outputs(3038) <= not a or b;
    layer4_outputs(3039) <= not b;
    layer4_outputs(3040) <= a or b;
    layer4_outputs(3041) <= a xor b;
    layer4_outputs(3042) <= a;
    layer4_outputs(3043) <= not (a and b);
    layer4_outputs(3044) <= not (a xor b);
    layer4_outputs(3045) <= a;
    layer4_outputs(3046) <= not b;
    layer4_outputs(3047) <= not a;
    layer4_outputs(3048) <= a and b;
    layer4_outputs(3049) <= a and b;
    layer4_outputs(3050) <= not (a or b);
    layer4_outputs(3051) <= b;
    layer4_outputs(3052) <= a xor b;
    layer4_outputs(3053) <= b;
    layer4_outputs(3054) <= not a;
    layer4_outputs(3055) <= not b or a;
    layer4_outputs(3056) <= b and not a;
    layer4_outputs(3057) <= not (a xor b);
    layer4_outputs(3058) <= a;
    layer4_outputs(3059) <= not (a or b);
    layer4_outputs(3060) <= not b;
    layer4_outputs(3061) <= not a;
    layer4_outputs(3062) <= not b;
    layer4_outputs(3063) <= b;
    layer4_outputs(3064) <= not a or b;
    layer4_outputs(3065) <= 1'b1;
    layer4_outputs(3066) <= a and b;
    layer4_outputs(3067) <= a and not b;
    layer4_outputs(3068) <= a or b;
    layer4_outputs(3069) <= not b;
    layer4_outputs(3070) <= not a;
    layer4_outputs(3071) <= a and not b;
    layer4_outputs(3072) <= a xor b;
    layer4_outputs(3073) <= a xor b;
    layer4_outputs(3074) <= b;
    layer4_outputs(3075) <= not b;
    layer4_outputs(3076) <= a and not b;
    layer4_outputs(3077) <= not a;
    layer4_outputs(3078) <= a xor b;
    layer4_outputs(3079) <= a and not b;
    layer4_outputs(3080) <= a;
    layer4_outputs(3081) <= a;
    layer4_outputs(3082) <= b;
    layer4_outputs(3083) <= not a;
    layer4_outputs(3084) <= a or b;
    layer4_outputs(3085) <= not a;
    layer4_outputs(3086) <= a and b;
    layer4_outputs(3087) <= not a;
    layer4_outputs(3088) <= b;
    layer4_outputs(3089) <= not a;
    layer4_outputs(3090) <= not (a or b);
    layer4_outputs(3091) <= not a;
    layer4_outputs(3092) <= b and not a;
    layer4_outputs(3093) <= not a or b;
    layer4_outputs(3094) <= b;
    layer4_outputs(3095) <= not (a xor b);
    layer4_outputs(3096) <= not a;
    layer4_outputs(3097) <= not (a or b);
    layer4_outputs(3098) <= not b;
    layer4_outputs(3099) <= a xor b;
    layer4_outputs(3100) <= not (a or b);
    layer4_outputs(3101) <= a;
    layer4_outputs(3102) <= a and b;
    layer4_outputs(3103) <= a and not b;
    layer4_outputs(3104) <= not a or b;
    layer4_outputs(3105) <= a;
    layer4_outputs(3106) <= a;
    layer4_outputs(3107) <= not a;
    layer4_outputs(3108) <= not a;
    layer4_outputs(3109) <= a xor b;
    layer4_outputs(3110) <= b;
    layer4_outputs(3111) <= not a;
    layer4_outputs(3112) <= not a;
    layer4_outputs(3113) <= not (a or b);
    layer4_outputs(3114) <= a xor b;
    layer4_outputs(3115) <= not a;
    layer4_outputs(3116) <= not b or a;
    layer4_outputs(3117) <= a or b;
    layer4_outputs(3118) <= not (a xor b);
    layer4_outputs(3119) <= a or b;
    layer4_outputs(3120) <= b;
    layer4_outputs(3121) <= b;
    layer4_outputs(3122) <= not (a or b);
    layer4_outputs(3123) <= a and not b;
    layer4_outputs(3124) <= not a;
    layer4_outputs(3125) <= not (a or b);
    layer4_outputs(3126) <= not a;
    layer4_outputs(3127) <= not a;
    layer4_outputs(3128) <= b and not a;
    layer4_outputs(3129) <= not (a and b);
    layer4_outputs(3130) <= not (a and b);
    layer4_outputs(3131) <= a or b;
    layer4_outputs(3132) <= not a;
    layer4_outputs(3133) <= a;
    layer4_outputs(3134) <= 1'b0;
    layer4_outputs(3135) <= not a;
    layer4_outputs(3136) <= not a or b;
    layer4_outputs(3137) <= not b or a;
    layer4_outputs(3138) <= not (a xor b);
    layer4_outputs(3139) <= a;
    layer4_outputs(3140) <= a;
    layer4_outputs(3141) <= a xor b;
    layer4_outputs(3142) <= not b;
    layer4_outputs(3143) <= not a or b;
    layer4_outputs(3144) <= a or b;
    layer4_outputs(3145) <= not (a xor b);
    layer4_outputs(3146) <= not a;
    layer4_outputs(3147) <= a xor b;
    layer4_outputs(3148) <= a and b;
    layer4_outputs(3149) <= a or b;
    layer4_outputs(3150) <= not (a xor b);
    layer4_outputs(3151) <= not (a xor b);
    layer4_outputs(3152) <= a and not b;
    layer4_outputs(3153) <= not (a xor b);
    layer4_outputs(3154) <= b;
    layer4_outputs(3155) <= a;
    layer4_outputs(3156) <= not a;
    layer4_outputs(3157) <= b;
    layer4_outputs(3158) <= not b or a;
    layer4_outputs(3159) <= not a;
    layer4_outputs(3160) <= b;
    layer4_outputs(3161) <= b;
    layer4_outputs(3162) <= a;
    layer4_outputs(3163) <= b and not a;
    layer4_outputs(3164) <= a xor b;
    layer4_outputs(3165) <= not b;
    layer4_outputs(3166) <= b and not a;
    layer4_outputs(3167) <= not b;
    layer4_outputs(3168) <= a and b;
    layer4_outputs(3169) <= a or b;
    layer4_outputs(3170) <= b and not a;
    layer4_outputs(3171) <= not b;
    layer4_outputs(3172) <= not b;
    layer4_outputs(3173) <= not b or a;
    layer4_outputs(3174) <= a;
    layer4_outputs(3175) <= not b or a;
    layer4_outputs(3176) <= not a;
    layer4_outputs(3177) <= a xor b;
    layer4_outputs(3178) <= b;
    layer4_outputs(3179) <= b;
    layer4_outputs(3180) <= not b;
    layer4_outputs(3181) <= b;
    layer4_outputs(3182) <= a and not b;
    layer4_outputs(3183) <= a;
    layer4_outputs(3184) <= not a;
    layer4_outputs(3185) <= not (a xor b);
    layer4_outputs(3186) <= a or b;
    layer4_outputs(3187) <= not (a or b);
    layer4_outputs(3188) <= a xor b;
    layer4_outputs(3189) <= not b or a;
    layer4_outputs(3190) <= a;
    layer4_outputs(3191) <= not b;
    layer4_outputs(3192) <= a and b;
    layer4_outputs(3193) <= not (a or b);
    layer4_outputs(3194) <= a xor b;
    layer4_outputs(3195) <= not b or a;
    layer4_outputs(3196) <= not (a xor b);
    layer4_outputs(3197) <= not (a and b);
    layer4_outputs(3198) <= not b or a;
    layer4_outputs(3199) <= a and b;
    layer4_outputs(3200) <= not (a xor b);
    layer4_outputs(3201) <= a xor b;
    layer4_outputs(3202) <= a xor b;
    layer4_outputs(3203) <= 1'b0;
    layer4_outputs(3204) <= b and not a;
    layer4_outputs(3205) <= not (a or b);
    layer4_outputs(3206) <= a xor b;
    layer4_outputs(3207) <= not a or b;
    layer4_outputs(3208) <= a;
    layer4_outputs(3209) <= b;
    layer4_outputs(3210) <= not (a xor b);
    layer4_outputs(3211) <= not b;
    layer4_outputs(3212) <= not (a xor b);
    layer4_outputs(3213) <= not b or a;
    layer4_outputs(3214) <= not b or a;
    layer4_outputs(3215) <= a or b;
    layer4_outputs(3216) <= not (a xor b);
    layer4_outputs(3217) <= b;
    layer4_outputs(3218) <= b and not a;
    layer4_outputs(3219) <= not a;
    layer4_outputs(3220) <= not b;
    layer4_outputs(3221) <= a;
    layer4_outputs(3222) <= a;
    layer4_outputs(3223) <= a and b;
    layer4_outputs(3224) <= a;
    layer4_outputs(3225) <= not b;
    layer4_outputs(3226) <= a;
    layer4_outputs(3227) <= a or b;
    layer4_outputs(3228) <= not a;
    layer4_outputs(3229) <= not a;
    layer4_outputs(3230) <= a;
    layer4_outputs(3231) <= not b;
    layer4_outputs(3232) <= a;
    layer4_outputs(3233) <= a or b;
    layer4_outputs(3234) <= a;
    layer4_outputs(3235) <= a xor b;
    layer4_outputs(3236) <= not b;
    layer4_outputs(3237) <= b;
    layer4_outputs(3238) <= not (a xor b);
    layer4_outputs(3239) <= not a;
    layer4_outputs(3240) <= not b;
    layer4_outputs(3241) <= not a;
    layer4_outputs(3242) <= a and b;
    layer4_outputs(3243) <= b;
    layer4_outputs(3244) <= not b;
    layer4_outputs(3245) <= b;
    layer4_outputs(3246) <= not (a or b);
    layer4_outputs(3247) <= b;
    layer4_outputs(3248) <= a;
    layer4_outputs(3249) <= a and b;
    layer4_outputs(3250) <= not (a or b);
    layer4_outputs(3251) <= b and not a;
    layer4_outputs(3252) <= b;
    layer4_outputs(3253) <= a and b;
    layer4_outputs(3254) <= not a or b;
    layer4_outputs(3255) <= b and not a;
    layer4_outputs(3256) <= a or b;
    layer4_outputs(3257) <= a;
    layer4_outputs(3258) <= not (a and b);
    layer4_outputs(3259) <= not b or a;
    layer4_outputs(3260) <= not b;
    layer4_outputs(3261) <= a;
    layer4_outputs(3262) <= a;
    layer4_outputs(3263) <= not b;
    layer4_outputs(3264) <= not a;
    layer4_outputs(3265) <= b;
    layer4_outputs(3266) <= a and not b;
    layer4_outputs(3267) <= a;
    layer4_outputs(3268) <= not (a xor b);
    layer4_outputs(3269) <= a xor b;
    layer4_outputs(3270) <= not (a xor b);
    layer4_outputs(3271) <= a xor b;
    layer4_outputs(3272) <= not b;
    layer4_outputs(3273) <= not b;
    layer4_outputs(3274) <= not (a or b);
    layer4_outputs(3275) <= not (a xor b);
    layer4_outputs(3276) <= not (a xor b);
    layer4_outputs(3277) <= not a;
    layer4_outputs(3278) <= b;
    layer4_outputs(3279) <= not a;
    layer4_outputs(3280) <= not b or a;
    layer4_outputs(3281) <= b;
    layer4_outputs(3282) <= not b;
    layer4_outputs(3283) <= not a;
    layer4_outputs(3284) <= a;
    layer4_outputs(3285) <= b;
    layer4_outputs(3286) <= b;
    layer4_outputs(3287) <= b;
    layer4_outputs(3288) <= 1'b0;
    layer4_outputs(3289) <= not a;
    layer4_outputs(3290) <= a and not b;
    layer4_outputs(3291) <= b;
    layer4_outputs(3292) <= a;
    layer4_outputs(3293) <= a or b;
    layer4_outputs(3294) <= a or b;
    layer4_outputs(3295) <= not a;
    layer4_outputs(3296) <= not (a or b);
    layer4_outputs(3297) <= a and not b;
    layer4_outputs(3298) <= not b or a;
    layer4_outputs(3299) <= not (a xor b);
    layer4_outputs(3300) <= not b;
    layer4_outputs(3301) <= not b or a;
    layer4_outputs(3302) <= not a or b;
    layer4_outputs(3303) <= b;
    layer4_outputs(3304) <= b;
    layer4_outputs(3305) <= not b;
    layer4_outputs(3306) <= not b;
    layer4_outputs(3307) <= a or b;
    layer4_outputs(3308) <= a or b;
    layer4_outputs(3309) <= b and not a;
    layer4_outputs(3310) <= b;
    layer4_outputs(3311) <= not b or a;
    layer4_outputs(3312) <= not (a and b);
    layer4_outputs(3313) <= a;
    layer4_outputs(3314) <= not b;
    layer4_outputs(3315) <= b;
    layer4_outputs(3316) <= not (a and b);
    layer4_outputs(3317) <= a and b;
    layer4_outputs(3318) <= not (a xor b);
    layer4_outputs(3319) <= a or b;
    layer4_outputs(3320) <= b and not a;
    layer4_outputs(3321) <= a and b;
    layer4_outputs(3322) <= not (a xor b);
    layer4_outputs(3323) <= a xor b;
    layer4_outputs(3324) <= b;
    layer4_outputs(3325) <= not a;
    layer4_outputs(3326) <= a or b;
    layer4_outputs(3327) <= a or b;
    layer4_outputs(3328) <= a and b;
    layer4_outputs(3329) <= not a or b;
    layer4_outputs(3330) <= not (a xor b);
    layer4_outputs(3331) <= b and not a;
    layer4_outputs(3332) <= not a or b;
    layer4_outputs(3333) <= b and not a;
    layer4_outputs(3334) <= b;
    layer4_outputs(3335) <= not (a or b);
    layer4_outputs(3336) <= not a;
    layer4_outputs(3337) <= not a;
    layer4_outputs(3338) <= not a;
    layer4_outputs(3339) <= not b;
    layer4_outputs(3340) <= not a;
    layer4_outputs(3341) <= a xor b;
    layer4_outputs(3342) <= a;
    layer4_outputs(3343) <= a xor b;
    layer4_outputs(3344) <= a or b;
    layer4_outputs(3345) <= not a or b;
    layer4_outputs(3346) <= not (a xor b);
    layer4_outputs(3347) <= not (a and b);
    layer4_outputs(3348) <= not a;
    layer4_outputs(3349) <= a;
    layer4_outputs(3350) <= not a;
    layer4_outputs(3351) <= a and not b;
    layer4_outputs(3352) <= a;
    layer4_outputs(3353) <= not a or b;
    layer4_outputs(3354) <= b;
    layer4_outputs(3355) <= a xor b;
    layer4_outputs(3356) <= a xor b;
    layer4_outputs(3357) <= not b;
    layer4_outputs(3358) <= not (a and b);
    layer4_outputs(3359) <= b and not a;
    layer4_outputs(3360) <= b;
    layer4_outputs(3361) <= a xor b;
    layer4_outputs(3362) <= not b or a;
    layer4_outputs(3363) <= not b;
    layer4_outputs(3364) <= not a;
    layer4_outputs(3365) <= not b;
    layer4_outputs(3366) <= not (a xor b);
    layer4_outputs(3367) <= not (a xor b);
    layer4_outputs(3368) <= b;
    layer4_outputs(3369) <= b;
    layer4_outputs(3370) <= not (a or b);
    layer4_outputs(3371) <= a and b;
    layer4_outputs(3372) <= not (a xor b);
    layer4_outputs(3373) <= a xor b;
    layer4_outputs(3374) <= b and not a;
    layer4_outputs(3375) <= not a;
    layer4_outputs(3376) <= a;
    layer4_outputs(3377) <= b and not a;
    layer4_outputs(3378) <= b;
    layer4_outputs(3379) <= b and not a;
    layer4_outputs(3380) <= a;
    layer4_outputs(3381) <= a xor b;
    layer4_outputs(3382) <= not (a xor b);
    layer4_outputs(3383) <= not a or b;
    layer4_outputs(3384) <= a xor b;
    layer4_outputs(3385) <= not (a xor b);
    layer4_outputs(3386) <= b and not a;
    layer4_outputs(3387) <= not (a or b);
    layer4_outputs(3388) <= b;
    layer4_outputs(3389) <= a;
    layer4_outputs(3390) <= a or b;
    layer4_outputs(3391) <= not (a xor b);
    layer4_outputs(3392) <= not b or a;
    layer4_outputs(3393) <= a xor b;
    layer4_outputs(3394) <= not (a or b);
    layer4_outputs(3395) <= a;
    layer4_outputs(3396) <= not (a or b);
    layer4_outputs(3397) <= not (a xor b);
    layer4_outputs(3398) <= not (a xor b);
    layer4_outputs(3399) <= not b;
    layer4_outputs(3400) <= not (a xor b);
    layer4_outputs(3401) <= not (a xor b);
    layer4_outputs(3402) <= b;
    layer4_outputs(3403) <= a;
    layer4_outputs(3404) <= a;
    layer4_outputs(3405) <= not a or b;
    layer4_outputs(3406) <= a xor b;
    layer4_outputs(3407) <= not b;
    layer4_outputs(3408) <= not a;
    layer4_outputs(3409) <= b and not a;
    layer4_outputs(3410) <= a xor b;
    layer4_outputs(3411) <= a;
    layer4_outputs(3412) <= a or b;
    layer4_outputs(3413) <= not b or a;
    layer4_outputs(3414) <= not (a xor b);
    layer4_outputs(3415) <= not b;
    layer4_outputs(3416) <= not (a and b);
    layer4_outputs(3417) <= not b;
    layer4_outputs(3418) <= not (a xor b);
    layer4_outputs(3419) <= not a;
    layer4_outputs(3420) <= not b;
    layer4_outputs(3421) <= a xor b;
    layer4_outputs(3422) <= not (a or b);
    layer4_outputs(3423) <= a;
    layer4_outputs(3424) <= a or b;
    layer4_outputs(3425) <= not (a or b);
    layer4_outputs(3426) <= not b or a;
    layer4_outputs(3427) <= a xor b;
    layer4_outputs(3428) <= not (a or b);
    layer4_outputs(3429) <= a or b;
    layer4_outputs(3430) <= not a or b;
    layer4_outputs(3431) <= a;
    layer4_outputs(3432) <= not (a xor b);
    layer4_outputs(3433) <= a xor b;
    layer4_outputs(3434) <= not b or a;
    layer4_outputs(3435) <= b;
    layer4_outputs(3436) <= not (a xor b);
    layer4_outputs(3437) <= b;
    layer4_outputs(3438) <= a and b;
    layer4_outputs(3439) <= a;
    layer4_outputs(3440) <= b;
    layer4_outputs(3441) <= a and b;
    layer4_outputs(3442) <= b;
    layer4_outputs(3443) <= a or b;
    layer4_outputs(3444) <= a;
    layer4_outputs(3445) <= a xor b;
    layer4_outputs(3446) <= a or b;
    layer4_outputs(3447) <= not (a xor b);
    layer4_outputs(3448) <= not a;
    layer4_outputs(3449) <= not b or a;
    layer4_outputs(3450) <= not (a xor b);
    layer4_outputs(3451) <= not b;
    layer4_outputs(3452) <= b and not a;
    layer4_outputs(3453) <= not b or a;
    layer4_outputs(3454) <= not (a xor b);
    layer4_outputs(3455) <= a or b;
    layer4_outputs(3456) <= a xor b;
    layer4_outputs(3457) <= not b or a;
    layer4_outputs(3458) <= a or b;
    layer4_outputs(3459) <= not (a xor b);
    layer4_outputs(3460) <= a and b;
    layer4_outputs(3461) <= not b;
    layer4_outputs(3462) <= not (a xor b);
    layer4_outputs(3463) <= a xor b;
    layer4_outputs(3464) <= not b or a;
    layer4_outputs(3465) <= not (a xor b);
    layer4_outputs(3466) <= not (a xor b);
    layer4_outputs(3467) <= a xor b;
    layer4_outputs(3468) <= a and not b;
    layer4_outputs(3469) <= not b;
    layer4_outputs(3470) <= not a or b;
    layer4_outputs(3471) <= not a;
    layer4_outputs(3472) <= a xor b;
    layer4_outputs(3473) <= a or b;
    layer4_outputs(3474) <= not b;
    layer4_outputs(3475) <= not a or b;
    layer4_outputs(3476) <= not (a and b);
    layer4_outputs(3477) <= a xor b;
    layer4_outputs(3478) <= a and b;
    layer4_outputs(3479) <= a or b;
    layer4_outputs(3480) <= not (a xor b);
    layer4_outputs(3481) <= not (a xor b);
    layer4_outputs(3482) <= a;
    layer4_outputs(3483) <= a;
    layer4_outputs(3484) <= not (a or b);
    layer4_outputs(3485) <= a xor b;
    layer4_outputs(3486) <= b;
    layer4_outputs(3487) <= not (a xor b);
    layer4_outputs(3488) <= a and not b;
    layer4_outputs(3489) <= not (a or b);
    layer4_outputs(3490) <= a or b;
    layer4_outputs(3491) <= not b;
    layer4_outputs(3492) <= a and not b;
    layer4_outputs(3493) <= a and not b;
    layer4_outputs(3494) <= not b or a;
    layer4_outputs(3495) <= not b;
    layer4_outputs(3496) <= a or b;
    layer4_outputs(3497) <= not a;
    layer4_outputs(3498) <= not a or b;
    layer4_outputs(3499) <= a or b;
    layer4_outputs(3500) <= not (a or b);
    layer4_outputs(3501) <= a and b;
    layer4_outputs(3502) <= a;
    layer4_outputs(3503) <= a xor b;
    layer4_outputs(3504) <= not (a xor b);
    layer4_outputs(3505) <= a xor b;
    layer4_outputs(3506) <= not b;
    layer4_outputs(3507) <= b;
    layer4_outputs(3508) <= a and b;
    layer4_outputs(3509) <= not (a and b);
    layer4_outputs(3510) <= not a or b;
    layer4_outputs(3511) <= b;
    layer4_outputs(3512) <= a;
    layer4_outputs(3513) <= a xor b;
    layer4_outputs(3514) <= not (a or b);
    layer4_outputs(3515) <= not (a xor b);
    layer4_outputs(3516) <= not (a xor b);
    layer4_outputs(3517) <= a;
    layer4_outputs(3518) <= a xor b;
    layer4_outputs(3519) <= b;
    layer4_outputs(3520) <= a xor b;
    layer4_outputs(3521) <= a and not b;
    layer4_outputs(3522) <= not b or a;
    layer4_outputs(3523) <= b and not a;
    layer4_outputs(3524) <= a and b;
    layer4_outputs(3525) <= not a or b;
    layer4_outputs(3526) <= not a;
    layer4_outputs(3527) <= b and not a;
    layer4_outputs(3528) <= 1'b0;
    layer4_outputs(3529) <= not a;
    layer4_outputs(3530) <= not a;
    layer4_outputs(3531) <= b and not a;
    layer4_outputs(3532) <= a and b;
    layer4_outputs(3533) <= a or b;
    layer4_outputs(3534) <= a or b;
    layer4_outputs(3535) <= b and not a;
    layer4_outputs(3536) <= a or b;
    layer4_outputs(3537) <= a;
    layer4_outputs(3538) <= not (a or b);
    layer4_outputs(3539) <= b;
    layer4_outputs(3540) <= not b or a;
    layer4_outputs(3541) <= not (a and b);
    layer4_outputs(3542) <= not b;
    layer4_outputs(3543) <= not b;
    layer4_outputs(3544) <= a xor b;
    layer4_outputs(3545) <= not a or b;
    layer4_outputs(3546) <= not a;
    layer4_outputs(3547) <= not a;
    layer4_outputs(3548) <= a or b;
    layer4_outputs(3549) <= not b;
    layer4_outputs(3550) <= b and not a;
    layer4_outputs(3551) <= not (a or b);
    layer4_outputs(3552) <= not (a or b);
    layer4_outputs(3553) <= not (a and b);
    layer4_outputs(3554) <= not a or b;
    layer4_outputs(3555) <= b;
    layer4_outputs(3556) <= not b;
    layer4_outputs(3557) <= a;
    layer4_outputs(3558) <= not a;
    layer4_outputs(3559) <= a;
    layer4_outputs(3560) <= not (a and b);
    layer4_outputs(3561) <= b and not a;
    layer4_outputs(3562) <= a;
    layer4_outputs(3563) <= not (a xor b);
    layer4_outputs(3564) <= b;
    layer4_outputs(3565) <= not b;
    layer4_outputs(3566) <= not a;
    layer4_outputs(3567) <= a;
    layer4_outputs(3568) <= a;
    layer4_outputs(3569) <= a;
    layer4_outputs(3570) <= not b;
    layer4_outputs(3571) <= not (a xor b);
    layer4_outputs(3572) <= not (a xor b);
    layer4_outputs(3573) <= b;
    layer4_outputs(3574) <= b;
    layer4_outputs(3575) <= not (a xor b);
    layer4_outputs(3576) <= not a or b;
    layer4_outputs(3577) <= not (a xor b);
    layer4_outputs(3578) <= b;
    layer4_outputs(3579) <= not (a and b);
    layer4_outputs(3580) <= not (a and b);
    layer4_outputs(3581) <= not b or a;
    layer4_outputs(3582) <= a xor b;
    layer4_outputs(3583) <= a;
    layer4_outputs(3584) <= not b;
    layer4_outputs(3585) <= not b or a;
    layer4_outputs(3586) <= a and not b;
    layer4_outputs(3587) <= not a;
    layer4_outputs(3588) <= not (a xor b);
    layer4_outputs(3589) <= not b or a;
    layer4_outputs(3590) <= a xor b;
    layer4_outputs(3591) <= b;
    layer4_outputs(3592) <= a or b;
    layer4_outputs(3593) <= not a or b;
    layer4_outputs(3594) <= not (a xor b);
    layer4_outputs(3595) <= not a;
    layer4_outputs(3596) <= not (a xor b);
    layer4_outputs(3597) <= a;
    layer4_outputs(3598) <= a or b;
    layer4_outputs(3599) <= not b;
    layer4_outputs(3600) <= a;
    layer4_outputs(3601) <= a;
    layer4_outputs(3602) <= not (a and b);
    layer4_outputs(3603) <= not (a xor b);
    layer4_outputs(3604) <= b;
    layer4_outputs(3605) <= not b;
    layer4_outputs(3606) <= a xor b;
    layer4_outputs(3607) <= not b;
    layer4_outputs(3608) <= a xor b;
    layer4_outputs(3609) <= not (a xor b);
    layer4_outputs(3610) <= not (a and b);
    layer4_outputs(3611) <= b;
    layer4_outputs(3612) <= not a;
    layer4_outputs(3613) <= b and not a;
    layer4_outputs(3614) <= not a;
    layer4_outputs(3615) <= not b;
    layer4_outputs(3616) <= a xor b;
    layer4_outputs(3617) <= not (a and b);
    layer4_outputs(3618) <= a or b;
    layer4_outputs(3619) <= a or b;
    layer4_outputs(3620) <= a and not b;
    layer4_outputs(3621) <= a;
    layer4_outputs(3622) <= not a;
    layer4_outputs(3623) <= not (a xor b);
    layer4_outputs(3624) <= b and not a;
    layer4_outputs(3625) <= not (a and b);
    layer4_outputs(3626) <= not b;
    layer4_outputs(3627) <= not a;
    layer4_outputs(3628) <= not b;
    layer4_outputs(3629) <= a or b;
    layer4_outputs(3630) <= not a;
    layer4_outputs(3631) <= a or b;
    layer4_outputs(3632) <= not a or b;
    layer4_outputs(3633) <= not b or a;
    layer4_outputs(3634) <= a xor b;
    layer4_outputs(3635) <= not (a and b);
    layer4_outputs(3636) <= not b;
    layer4_outputs(3637) <= b and not a;
    layer4_outputs(3638) <= not b;
    layer4_outputs(3639) <= not (a and b);
    layer4_outputs(3640) <= not a or b;
    layer4_outputs(3641) <= not b or a;
    layer4_outputs(3642) <= a and not b;
    layer4_outputs(3643) <= not a or b;
    layer4_outputs(3644) <= b;
    layer4_outputs(3645) <= not a or b;
    layer4_outputs(3646) <= not b;
    layer4_outputs(3647) <= a;
    layer4_outputs(3648) <= a xor b;
    layer4_outputs(3649) <= not b;
    layer4_outputs(3650) <= b;
    layer4_outputs(3651) <= not a;
    layer4_outputs(3652) <= a and not b;
    layer4_outputs(3653) <= b and not a;
    layer4_outputs(3654) <= a;
    layer4_outputs(3655) <= b and not a;
    layer4_outputs(3656) <= not (a xor b);
    layer4_outputs(3657) <= a and not b;
    layer4_outputs(3658) <= a;
    layer4_outputs(3659) <= not b;
    layer4_outputs(3660) <= not b;
    layer4_outputs(3661) <= not a or b;
    layer4_outputs(3662) <= not a;
    layer4_outputs(3663) <= b and not a;
    layer4_outputs(3664) <= a xor b;
    layer4_outputs(3665) <= not (a and b);
    layer4_outputs(3666) <= b;
    layer4_outputs(3667) <= a;
    layer4_outputs(3668) <= a;
    layer4_outputs(3669) <= not a or b;
    layer4_outputs(3670) <= b;
    layer4_outputs(3671) <= not a;
    layer4_outputs(3672) <= not a or b;
    layer4_outputs(3673) <= a xor b;
    layer4_outputs(3674) <= not b;
    layer4_outputs(3675) <= a;
    layer4_outputs(3676) <= not a;
    layer4_outputs(3677) <= not a;
    layer4_outputs(3678) <= not (a xor b);
    layer4_outputs(3679) <= 1'b0;
    layer4_outputs(3680) <= a xor b;
    layer4_outputs(3681) <= not (a or b);
    layer4_outputs(3682) <= a xor b;
    layer4_outputs(3683) <= a and not b;
    layer4_outputs(3684) <= a;
    layer4_outputs(3685) <= not (a xor b);
    layer4_outputs(3686) <= not a;
    layer4_outputs(3687) <= a;
    layer4_outputs(3688) <= not b;
    layer4_outputs(3689) <= a xor b;
    layer4_outputs(3690) <= b;
    layer4_outputs(3691) <= not (a xor b);
    layer4_outputs(3692) <= b;
    layer4_outputs(3693) <= not (a or b);
    layer4_outputs(3694) <= a;
    layer4_outputs(3695) <= b;
    layer4_outputs(3696) <= a and b;
    layer4_outputs(3697) <= a and not b;
    layer4_outputs(3698) <= b;
    layer4_outputs(3699) <= b;
    layer4_outputs(3700) <= a or b;
    layer4_outputs(3701) <= not (a and b);
    layer4_outputs(3702) <= not b;
    layer4_outputs(3703) <= b;
    layer4_outputs(3704) <= not (a and b);
    layer4_outputs(3705) <= not a;
    layer4_outputs(3706) <= a and not b;
    layer4_outputs(3707) <= b;
    layer4_outputs(3708) <= not (a xor b);
    layer4_outputs(3709) <= a and not b;
    layer4_outputs(3710) <= a;
    layer4_outputs(3711) <= a or b;
    layer4_outputs(3712) <= a or b;
    layer4_outputs(3713) <= a xor b;
    layer4_outputs(3714) <= not (a or b);
    layer4_outputs(3715) <= not a;
    layer4_outputs(3716) <= a;
    layer4_outputs(3717) <= a;
    layer4_outputs(3718) <= not b;
    layer4_outputs(3719) <= not (a and b);
    layer4_outputs(3720) <= a and not b;
    layer4_outputs(3721) <= b;
    layer4_outputs(3722) <= not a or b;
    layer4_outputs(3723) <= a;
    layer4_outputs(3724) <= not (a or b);
    layer4_outputs(3725) <= not b or a;
    layer4_outputs(3726) <= not b or a;
    layer4_outputs(3727) <= not b or a;
    layer4_outputs(3728) <= not b or a;
    layer4_outputs(3729) <= a or b;
    layer4_outputs(3730) <= a and not b;
    layer4_outputs(3731) <= a;
    layer4_outputs(3732) <= a and not b;
    layer4_outputs(3733) <= not (a or b);
    layer4_outputs(3734) <= not b;
    layer4_outputs(3735) <= not b or a;
    layer4_outputs(3736) <= not b;
    layer4_outputs(3737) <= a;
    layer4_outputs(3738) <= a and not b;
    layer4_outputs(3739) <= not (a xor b);
    layer4_outputs(3740) <= not b or a;
    layer4_outputs(3741) <= not a;
    layer4_outputs(3742) <= not b;
    layer4_outputs(3743) <= not (a and b);
    layer4_outputs(3744) <= a and b;
    layer4_outputs(3745) <= not (a and b);
    layer4_outputs(3746) <= a and not b;
    layer4_outputs(3747) <= not b;
    layer4_outputs(3748) <= not b;
    layer4_outputs(3749) <= a xor b;
    layer4_outputs(3750) <= not b or a;
    layer4_outputs(3751) <= not b;
    layer4_outputs(3752) <= not b;
    layer4_outputs(3753) <= a xor b;
    layer4_outputs(3754) <= a;
    layer4_outputs(3755) <= not a;
    layer4_outputs(3756) <= a;
    layer4_outputs(3757) <= a xor b;
    layer4_outputs(3758) <= a xor b;
    layer4_outputs(3759) <= not a;
    layer4_outputs(3760) <= not a;
    layer4_outputs(3761) <= not a;
    layer4_outputs(3762) <= not a;
    layer4_outputs(3763) <= not a or b;
    layer4_outputs(3764) <= not (a or b);
    layer4_outputs(3765) <= not (a and b);
    layer4_outputs(3766) <= not b;
    layer4_outputs(3767) <= not a;
    layer4_outputs(3768) <= a;
    layer4_outputs(3769) <= b and not a;
    layer4_outputs(3770) <= a and not b;
    layer4_outputs(3771) <= not (a or b);
    layer4_outputs(3772) <= a or b;
    layer4_outputs(3773) <= not b;
    layer4_outputs(3774) <= not (a xor b);
    layer4_outputs(3775) <= not a or b;
    layer4_outputs(3776) <= b;
    layer4_outputs(3777) <= a;
    layer4_outputs(3778) <= a or b;
    layer4_outputs(3779) <= not a;
    layer4_outputs(3780) <= not a;
    layer4_outputs(3781) <= not (a or b);
    layer4_outputs(3782) <= not a or b;
    layer4_outputs(3783) <= not b;
    layer4_outputs(3784) <= a xor b;
    layer4_outputs(3785) <= b;
    layer4_outputs(3786) <= not a or b;
    layer4_outputs(3787) <= not a or b;
    layer4_outputs(3788) <= a or b;
    layer4_outputs(3789) <= a and b;
    layer4_outputs(3790) <= a;
    layer4_outputs(3791) <= not (a or b);
    layer4_outputs(3792) <= a;
    layer4_outputs(3793) <= a and b;
    layer4_outputs(3794) <= not (a xor b);
    layer4_outputs(3795) <= not a;
    layer4_outputs(3796) <= not b;
    layer4_outputs(3797) <= a xor b;
    layer4_outputs(3798) <= not (a and b);
    layer4_outputs(3799) <= a;
    layer4_outputs(3800) <= b and not a;
    layer4_outputs(3801) <= a and not b;
    layer4_outputs(3802) <= a or b;
    layer4_outputs(3803) <= b;
    layer4_outputs(3804) <= b;
    layer4_outputs(3805) <= not (a or b);
    layer4_outputs(3806) <= not (a xor b);
    layer4_outputs(3807) <= not b or a;
    layer4_outputs(3808) <= not (a xor b);
    layer4_outputs(3809) <= not (a and b);
    layer4_outputs(3810) <= not b or a;
    layer4_outputs(3811) <= a;
    layer4_outputs(3812) <= not b;
    layer4_outputs(3813) <= not a;
    layer4_outputs(3814) <= b and not a;
    layer4_outputs(3815) <= a;
    layer4_outputs(3816) <= b;
    layer4_outputs(3817) <= not b or a;
    layer4_outputs(3818) <= not (a and b);
    layer4_outputs(3819) <= not (a xor b);
    layer4_outputs(3820) <= a and b;
    layer4_outputs(3821) <= not b or a;
    layer4_outputs(3822) <= not (a xor b);
    layer4_outputs(3823) <= not b or a;
    layer4_outputs(3824) <= not b;
    layer4_outputs(3825) <= a xor b;
    layer4_outputs(3826) <= not b or a;
    layer4_outputs(3827) <= a or b;
    layer4_outputs(3828) <= b;
    layer4_outputs(3829) <= not b;
    layer4_outputs(3830) <= not a or b;
    layer4_outputs(3831) <= a;
    layer4_outputs(3832) <= not a or b;
    layer4_outputs(3833) <= b;
    layer4_outputs(3834) <= not a;
    layer4_outputs(3835) <= not a;
    layer4_outputs(3836) <= not a;
    layer4_outputs(3837) <= not (a and b);
    layer4_outputs(3838) <= a xor b;
    layer4_outputs(3839) <= a;
    layer4_outputs(3840) <= not (a xor b);
    layer4_outputs(3841) <= not b or a;
    layer4_outputs(3842) <= b;
    layer4_outputs(3843) <= b;
    layer4_outputs(3844) <= not b;
    layer4_outputs(3845) <= a or b;
    layer4_outputs(3846) <= not (a xor b);
    layer4_outputs(3847) <= not b;
    layer4_outputs(3848) <= not b or a;
    layer4_outputs(3849) <= not (a and b);
    layer4_outputs(3850) <= not (a xor b);
    layer4_outputs(3851) <= not b or a;
    layer4_outputs(3852) <= not b;
    layer4_outputs(3853) <= a;
    layer4_outputs(3854) <= not a;
    layer4_outputs(3855) <= a or b;
    layer4_outputs(3856) <= b;
    layer4_outputs(3857) <= not b;
    layer4_outputs(3858) <= b;
    layer4_outputs(3859) <= not (a and b);
    layer4_outputs(3860) <= a xor b;
    layer4_outputs(3861) <= a;
    layer4_outputs(3862) <= a;
    layer4_outputs(3863) <= not (a xor b);
    layer4_outputs(3864) <= not (a xor b);
    layer4_outputs(3865) <= not b;
    layer4_outputs(3866) <= a;
    layer4_outputs(3867) <= a and not b;
    layer4_outputs(3868) <= a xor b;
    layer4_outputs(3869) <= b;
    layer4_outputs(3870) <= not b;
    layer4_outputs(3871) <= not b;
    layer4_outputs(3872) <= not a;
    layer4_outputs(3873) <= a and not b;
    layer4_outputs(3874) <= b;
    layer4_outputs(3875) <= a and not b;
    layer4_outputs(3876) <= b;
    layer4_outputs(3877) <= a;
    layer4_outputs(3878) <= a;
    layer4_outputs(3879) <= a;
    layer4_outputs(3880) <= not b or a;
    layer4_outputs(3881) <= not b;
    layer4_outputs(3882) <= not (a xor b);
    layer4_outputs(3883) <= not (a or b);
    layer4_outputs(3884) <= not a or b;
    layer4_outputs(3885) <= not a or b;
    layer4_outputs(3886) <= a xor b;
    layer4_outputs(3887) <= not (a xor b);
    layer4_outputs(3888) <= not (a and b);
    layer4_outputs(3889) <= not (a and b);
    layer4_outputs(3890) <= not (a xor b);
    layer4_outputs(3891) <= a xor b;
    layer4_outputs(3892) <= a and b;
    layer4_outputs(3893) <= not b;
    layer4_outputs(3894) <= not a or b;
    layer4_outputs(3895) <= 1'b0;
    layer4_outputs(3896) <= not b or a;
    layer4_outputs(3897) <= not (a and b);
    layer4_outputs(3898) <= a xor b;
    layer4_outputs(3899) <= a or b;
    layer4_outputs(3900) <= a xor b;
    layer4_outputs(3901) <= not b or a;
    layer4_outputs(3902) <= a and not b;
    layer4_outputs(3903) <= not b;
    layer4_outputs(3904) <= b;
    layer4_outputs(3905) <= not a;
    layer4_outputs(3906) <= not (a xor b);
    layer4_outputs(3907) <= not b;
    layer4_outputs(3908) <= a xor b;
    layer4_outputs(3909) <= a or b;
    layer4_outputs(3910) <= not a or b;
    layer4_outputs(3911) <= a;
    layer4_outputs(3912) <= a or b;
    layer4_outputs(3913) <= not (a and b);
    layer4_outputs(3914) <= not a;
    layer4_outputs(3915) <= not b;
    layer4_outputs(3916) <= not b;
    layer4_outputs(3917) <= a xor b;
    layer4_outputs(3918) <= not a;
    layer4_outputs(3919) <= not (a and b);
    layer4_outputs(3920) <= a;
    layer4_outputs(3921) <= b;
    layer4_outputs(3922) <= not a or b;
    layer4_outputs(3923) <= not (a and b);
    layer4_outputs(3924) <= b;
    layer4_outputs(3925) <= not a;
    layer4_outputs(3926) <= a;
    layer4_outputs(3927) <= not b;
    layer4_outputs(3928) <= not (a or b);
    layer4_outputs(3929) <= not b or a;
    layer4_outputs(3930) <= b and not a;
    layer4_outputs(3931) <= a or b;
    layer4_outputs(3932) <= a;
    layer4_outputs(3933) <= a;
    layer4_outputs(3934) <= a xor b;
    layer4_outputs(3935) <= not (a xor b);
    layer4_outputs(3936) <= not (a or b);
    layer4_outputs(3937) <= a;
    layer4_outputs(3938) <= b;
    layer4_outputs(3939) <= not (a and b);
    layer4_outputs(3940) <= not b or a;
    layer4_outputs(3941) <= a and b;
    layer4_outputs(3942) <= b and not a;
    layer4_outputs(3943) <= a and not b;
    layer4_outputs(3944) <= not b or a;
    layer4_outputs(3945) <= a and not b;
    layer4_outputs(3946) <= not (a and b);
    layer4_outputs(3947) <= a xor b;
    layer4_outputs(3948) <= not b;
    layer4_outputs(3949) <= a xor b;
    layer4_outputs(3950) <= not b or a;
    layer4_outputs(3951) <= not (a xor b);
    layer4_outputs(3952) <= not (a and b);
    layer4_outputs(3953) <= b and not a;
    layer4_outputs(3954) <= a xor b;
    layer4_outputs(3955) <= not (a or b);
    layer4_outputs(3956) <= not b;
    layer4_outputs(3957) <= a and not b;
    layer4_outputs(3958) <= b;
    layer4_outputs(3959) <= not (a xor b);
    layer4_outputs(3960) <= a and b;
    layer4_outputs(3961) <= a;
    layer4_outputs(3962) <= not a or b;
    layer4_outputs(3963) <= not b or a;
    layer4_outputs(3964) <= a and b;
    layer4_outputs(3965) <= not (a or b);
    layer4_outputs(3966) <= not b;
    layer4_outputs(3967) <= a or b;
    layer4_outputs(3968) <= not b;
    layer4_outputs(3969) <= a and not b;
    layer4_outputs(3970) <= b;
    layer4_outputs(3971) <= a and b;
    layer4_outputs(3972) <= a and b;
    layer4_outputs(3973) <= not (a xor b);
    layer4_outputs(3974) <= not b or a;
    layer4_outputs(3975) <= not (a or b);
    layer4_outputs(3976) <= not (a and b);
    layer4_outputs(3977) <= not a;
    layer4_outputs(3978) <= a and not b;
    layer4_outputs(3979) <= not a;
    layer4_outputs(3980) <= b;
    layer4_outputs(3981) <= a;
    layer4_outputs(3982) <= not a;
    layer4_outputs(3983) <= a or b;
    layer4_outputs(3984) <= a xor b;
    layer4_outputs(3985) <= a or b;
    layer4_outputs(3986) <= a;
    layer4_outputs(3987) <= a and not b;
    layer4_outputs(3988) <= a;
    layer4_outputs(3989) <= not (a xor b);
    layer4_outputs(3990) <= not (a xor b);
    layer4_outputs(3991) <= not b;
    layer4_outputs(3992) <= not (a xor b);
    layer4_outputs(3993) <= not b;
    layer4_outputs(3994) <= not a or b;
    layer4_outputs(3995) <= not a;
    layer4_outputs(3996) <= not b;
    layer4_outputs(3997) <= a or b;
    layer4_outputs(3998) <= not b;
    layer4_outputs(3999) <= b;
    layer4_outputs(4000) <= b;
    layer4_outputs(4001) <= not a or b;
    layer4_outputs(4002) <= not a or b;
    layer4_outputs(4003) <= not b or a;
    layer4_outputs(4004) <= not (a and b);
    layer4_outputs(4005) <= a and not b;
    layer4_outputs(4006) <= not (a xor b);
    layer4_outputs(4007) <= not a;
    layer4_outputs(4008) <= a;
    layer4_outputs(4009) <= not a;
    layer4_outputs(4010) <= not a;
    layer4_outputs(4011) <= a and not b;
    layer4_outputs(4012) <= not a;
    layer4_outputs(4013) <= a and b;
    layer4_outputs(4014) <= not b;
    layer4_outputs(4015) <= a;
    layer4_outputs(4016) <= a xor b;
    layer4_outputs(4017) <= a;
    layer4_outputs(4018) <= not a;
    layer4_outputs(4019) <= not b;
    layer4_outputs(4020) <= a and b;
    layer4_outputs(4021) <= a;
    layer4_outputs(4022) <= not (a xor b);
    layer4_outputs(4023) <= a;
    layer4_outputs(4024) <= a or b;
    layer4_outputs(4025) <= not a;
    layer4_outputs(4026) <= not a;
    layer4_outputs(4027) <= b and not a;
    layer4_outputs(4028) <= not (a and b);
    layer4_outputs(4029) <= a or b;
    layer4_outputs(4030) <= not (a xor b);
    layer4_outputs(4031) <= b;
    layer4_outputs(4032) <= a xor b;
    layer4_outputs(4033) <= not a;
    layer4_outputs(4034) <= not (a xor b);
    layer4_outputs(4035) <= not a;
    layer4_outputs(4036) <= a and not b;
    layer4_outputs(4037) <= not (a and b);
    layer4_outputs(4038) <= not (a and b);
    layer4_outputs(4039) <= not (a or b);
    layer4_outputs(4040) <= a;
    layer4_outputs(4041) <= a or b;
    layer4_outputs(4042) <= a xor b;
    layer4_outputs(4043) <= a;
    layer4_outputs(4044) <= not a or b;
    layer4_outputs(4045) <= b;
    layer4_outputs(4046) <= b and not a;
    layer4_outputs(4047) <= a;
    layer4_outputs(4048) <= not a;
    layer4_outputs(4049) <= a;
    layer4_outputs(4050) <= not b or a;
    layer4_outputs(4051) <= a and not b;
    layer4_outputs(4052) <= a and b;
    layer4_outputs(4053) <= a and not b;
    layer4_outputs(4054) <= b and not a;
    layer4_outputs(4055) <= not a;
    layer4_outputs(4056) <= not a;
    layer4_outputs(4057) <= a and b;
    layer4_outputs(4058) <= not (a or b);
    layer4_outputs(4059) <= b;
    layer4_outputs(4060) <= a;
    layer4_outputs(4061) <= not a;
    layer4_outputs(4062) <= a or b;
    layer4_outputs(4063) <= a and b;
    layer4_outputs(4064) <= a xor b;
    layer4_outputs(4065) <= a and b;
    layer4_outputs(4066) <= not a or b;
    layer4_outputs(4067) <= not (a and b);
    layer4_outputs(4068) <= b;
    layer4_outputs(4069) <= b;
    layer4_outputs(4070) <= not b;
    layer4_outputs(4071) <= a xor b;
    layer4_outputs(4072) <= b;
    layer4_outputs(4073) <= a xor b;
    layer4_outputs(4074) <= a or b;
    layer4_outputs(4075) <= a and not b;
    layer4_outputs(4076) <= not (a and b);
    layer4_outputs(4077) <= not a or b;
    layer4_outputs(4078) <= not b;
    layer4_outputs(4079) <= not a or b;
    layer4_outputs(4080) <= not a or b;
    layer4_outputs(4081) <= not b or a;
    layer4_outputs(4082) <= b;
    layer4_outputs(4083) <= a and not b;
    layer4_outputs(4084) <= not (a or b);
    layer4_outputs(4085) <= a and not b;
    layer4_outputs(4086) <= not (a or b);
    layer4_outputs(4087) <= a and not b;
    layer4_outputs(4088) <= b;
    layer4_outputs(4089) <= not (a and b);
    layer4_outputs(4090) <= b;
    layer4_outputs(4091) <= a and b;
    layer4_outputs(4092) <= a or b;
    layer4_outputs(4093) <= not (a or b);
    layer4_outputs(4094) <= a or b;
    layer4_outputs(4095) <= a;
    layer4_outputs(4096) <= not a;
    layer4_outputs(4097) <= not b;
    layer4_outputs(4098) <= a xor b;
    layer4_outputs(4099) <= a;
    layer4_outputs(4100) <= a;
    layer4_outputs(4101) <= a xor b;
    layer4_outputs(4102) <= a;
    layer4_outputs(4103) <= not a;
    layer4_outputs(4104) <= a and b;
    layer4_outputs(4105) <= a;
    layer4_outputs(4106) <= b and not a;
    layer4_outputs(4107) <= not b;
    layer4_outputs(4108) <= a or b;
    layer4_outputs(4109) <= a or b;
    layer4_outputs(4110) <= b;
    layer4_outputs(4111) <= a and b;
    layer4_outputs(4112) <= not (a xor b);
    layer4_outputs(4113) <= a and not b;
    layer4_outputs(4114) <= a;
    layer4_outputs(4115) <= not b or a;
    layer4_outputs(4116) <= a;
    layer4_outputs(4117) <= not b;
    layer4_outputs(4118) <= a xor b;
    layer4_outputs(4119) <= not b;
    layer4_outputs(4120) <= b;
    layer4_outputs(4121) <= not a;
    layer4_outputs(4122) <= a and b;
    layer4_outputs(4123) <= a and not b;
    layer4_outputs(4124) <= not (a or b);
    layer4_outputs(4125) <= a and b;
    layer4_outputs(4126) <= a and b;
    layer4_outputs(4127) <= a or b;
    layer4_outputs(4128) <= a and b;
    layer4_outputs(4129) <= a;
    layer4_outputs(4130) <= a;
    layer4_outputs(4131) <= not b or a;
    layer4_outputs(4132) <= not a or b;
    layer4_outputs(4133) <= b;
    layer4_outputs(4134) <= not (a and b);
    layer4_outputs(4135) <= b;
    layer4_outputs(4136) <= not b;
    layer4_outputs(4137) <= b;
    layer4_outputs(4138) <= b;
    layer4_outputs(4139) <= a;
    layer4_outputs(4140) <= a;
    layer4_outputs(4141) <= not (a and b);
    layer4_outputs(4142) <= not a;
    layer4_outputs(4143) <= a and b;
    layer4_outputs(4144) <= not b;
    layer4_outputs(4145) <= not b;
    layer4_outputs(4146) <= not a;
    layer4_outputs(4147) <= a;
    layer4_outputs(4148) <= not b;
    layer4_outputs(4149) <= a;
    layer4_outputs(4150) <= b;
    layer4_outputs(4151) <= a and not b;
    layer4_outputs(4152) <= not a;
    layer4_outputs(4153) <= b;
    layer4_outputs(4154) <= not b or a;
    layer4_outputs(4155) <= not a;
    layer4_outputs(4156) <= not b or a;
    layer4_outputs(4157) <= not a;
    layer4_outputs(4158) <= not b;
    layer4_outputs(4159) <= not (a and b);
    layer4_outputs(4160) <= not b;
    layer4_outputs(4161) <= not b;
    layer4_outputs(4162) <= a xor b;
    layer4_outputs(4163) <= not a;
    layer4_outputs(4164) <= not (a and b);
    layer4_outputs(4165) <= b;
    layer4_outputs(4166) <= not (a xor b);
    layer4_outputs(4167) <= not (a xor b);
    layer4_outputs(4168) <= a xor b;
    layer4_outputs(4169) <= b;
    layer4_outputs(4170) <= not b;
    layer4_outputs(4171) <= a and b;
    layer4_outputs(4172) <= not b;
    layer4_outputs(4173) <= a;
    layer4_outputs(4174) <= not (a or b);
    layer4_outputs(4175) <= a xor b;
    layer4_outputs(4176) <= not (a and b);
    layer4_outputs(4177) <= a;
    layer4_outputs(4178) <= not b;
    layer4_outputs(4179) <= b;
    layer4_outputs(4180) <= not b;
    layer4_outputs(4181) <= not a;
    layer4_outputs(4182) <= not b;
    layer4_outputs(4183) <= a and b;
    layer4_outputs(4184) <= a xor b;
    layer4_outputs(4185) <= a xor b;
    layer4_outputs(4186) <= not b;
    layer4_outputs(4187) <= not (a or b);
    layer4_outputs(4188) <= b;
    layer4_outputs(4189) <= b;
    layer4_outputs(4190) <= a or b;
    layer4_outputs(4191) <= not a;
    layer4_outputs(4192) <= not (a xor b);
    layer4_outputs(4193) <= b;
    layer4_outputs(4194) <= not a or b;
    layer4_outputs(4195) <= not (a and b);
    layer4_outputs(4196) <= not a or b;
    layer4_outputs(4197) <= a xor b;
    layer4_outputs(4198) <= not b or a;
    layer4_outputs(4199) <= not b;
    layer4_outputs(4200) <= not a;
    layer4_outputs(4201) <= not b;
    layer4_outputs(4202) <= a;
    layer4_outputs(4203) <= b;
    layer4_outputs(4204) <= a;
    layer4_outputs(4205) <= not b or a;
    layer4_outputs(4206) <= a;
    layer4_outputs(4207) <= b;
    layer4_outputs(4208) <= not (a and b);
    layer4_outputs(4209) <= not b;
    layer4_outputs(4210) <= b and not a;
    layer4_outputs(4211) <= not a;
    layer4_outputs(4212) <= not b or a;
    layer4_outputs(4213) <= not b;
    layer4_outputs(4214) <= not a or b;
    layer4_outputs(4215) <= not a or b;
    layer4_outputs(4216) <= a xor b;
    layer4_outputs(4217) <= a;
    layer4_outputs(4218) <= a or b;
    layer4_outputs(4219) <= b and not a;
    layer4_outputs(4220) <= a and not b;
    layer4_outputs(4221) <= b;
    layer4_outputs(4222) <= not (a xor b);
    layer4_outputs(4223) <= b;
    layer4_outputs(4224) <= b and not a;
    layer4_outputs(4225) <= not (a xor b);
    layer4_outputs(4226) <= b;
    layer4_outputs(4227) <= not (a or b);
    layer4_outputs(4228) <= 1'b1;
    layer4_outputs(4229) <= not (a or b);
    layer4_outputs(4230) <= a and b;
    layer4_outputs(4231) <= not b;
    layer4_outputs(4232) <= not b or a;
    layer4_outputs(4233) <= a xor b;
    layer4_outputs(4234) <= a and not b;
    layer4_outputs(4235) <= not a;
    layer4_outputs(4236) <= b;
    layer4_outputs(4237) <= a xor b;
    layer4_outputs(4238) <= a or b;
    layer4_outputs(4239) <= not (a xor b);
    layer4_outputs(4240) <= not a;
    layer4_outputs(4241) <= a;
    layer4_outputs(4242) <= not b;
    layer4_outputs(4243) <= not (a xor b);
    layer4_outputs(4244) <= not a;
    layer4_outputs(4245) <= b;
    layer4_outputs(4246) <= not b or a;
    layer4_outputs(4247) <= a or b;
    layer4_outputs(4248) <= not (a or b);
    layer4_outputs(4249) <= a;
    layer4_outputs(4250) <= not (a and b);
    layer4_outputs(4251) <= not (a xor b);
    layer4_outputs(4252) <= a;
    layer4_outputs(4253) <= not b or a;
    layer4_outputs(4254) <= not a or b;
    layer4_outputs(4255) <= not (a or b);
    layer4_outputs(4256) <= a xor b;
    layer4_outputs(4257) <= b and not a;
    layer4_outputs(4258) <= not b or a;
    layer4_outputs(4259) <= not (a xor b);
    layer4_outputs(4260) <= not a;
    layer4_outputs(4261) <= not b;
    layer4_outputs(4262) <= a and b;
    layer4_outputs(4263) <= a or b;
    layer4_outputs(4264) <= a and b;
    layer4_outputs(4265) <= not b or a;
    layer4_outputs(4266) <= not (a or b);
    layer4_outputs(4267) <= a and not b;
    layer4_outputs(4268) <= b and not a;
    layer4_outputs(4269) <= not b;
    layer4_outputs(4270) <= a and b;
    layer4_outputs(4271) <= not (a xor b);
    layer4_outputs(4272) <= a xor b;
    layer4_outputs(4273) <= not b;
    layer4_outputs(4274) <= b;
    layer4_outputs(4275) <= a;
    layer4_outputs(4276) <= not (a or b);
    layer4_outputs(4277) <= not b;
    layer4_outputs(4278) <= a;
    layer4_outputs(4279) <= not b;
    layer4_outputs(4280) <= not a or b;
    layer4_outputs(4281) <= not (a xor b);
    layer4_outputs(4282) <= not (a or b);
    layer4_outputs(4283) <= not (a and b);
    layer4_outputs(4284) <= not b;
    layer4_outputs(4285) <= a;
    layer4_outputs(4286) <= not a;
    layer4_outputs(4287) <= a or b;
    layer4_outputs(4288) <= a or b;
    layer4_outputs(4289) <= not b;
    layer4_outputs(4290) <= not a or b;
    layer4_outputs(4291) <= not b;
    layer4_outputs(4292) <= not (a and b);
    layer4_outputs(4293) <= a and b;
    layer4_outputs(4294) <= not b;
    layer4_outputs(4295) <= a xor b;
    layer4_outputs(4296) <= a;
    layer4_outputs(4297) <= a or b;
    layer4_outputs(4298) <= not a;
    layer4_outputs(4299) <= not a;
    layer4_outputs(4300) <= not (a xor b);
    layer4_outputs(4301) <= not (a xor b);
    layer4_outputs(4302) <= b;
    layer4_outputs(4303) <= not b;
    layer4_outputs(4304) <= not (a and b);
    layer4_outputs(4305) <= a;
    layer4_outputs(4306) <= a;
    layer4_outputs(4307) <= not (a or b);
    layer4_outputs(4308) <= 1'b0;
    layer4_outputs(4309) <= a xor b;
    layer4_outputs(4310) <= not b or a;
    layer4_outputs(4311) <= a xor b;
    layer4_outputs(4312) <= not a or b;
    layer4_outputs(4313) <= a xor b;
    layer4_outputs(4314) <= a;
    layer4_outputs(4315) <= a;
    layer4_outputs(4316) <= not (a and b);
    layer4_outputs(4317) <= a;
    layer4_outputs(4318) <= not (a and b);
    layer4_outputs(4319) <= a xor b;
    layer4_outputs(4320) <= b and not a;
    layer4_outputs(4321) <= not a;
    layer4_outputs(4322) <= not b;
    layer4_outputs(4323) <= not (a or b);
    layer4_outputs(4324) <= a;
    layer4_outputs(4325) <= a xor b;
    layer4_outputs(4326) <= a and b;
    layer4_outputs(4327) <= a and b;
    layer4_outputs(4328) <= not b;
    layer4_outputs(4329) <= a;
    layer4_outputs(4330) <= not b or a;
    layer4_outputs(4331) <= a and b;
    layer4_outputs(4332) <= a;
    layer4_outputs(4333) <= a and b;
    layer4_outputs(4334) <= not b or a;
    layer4_outputs(4335) <= a;
    layer4_outputs(4336) <= a xor b;
    layer4_outputs(4337) <= a;
    layer4_outputs(4338) <= not b;
    layer4_outputs(4339) <= b;
    layer4_outputs(4340) <= a and not b;
    layer4_outputs(4341) <= not b;
    layer4_outputs(4342) <= not a or b;
    layer4_outputs(4343) <= a or b;
    layer4_outputs(4344) <= a;
    layer4_outputs(4345) <= not b;
    layer4_outputs(4346) <= a;
    layer4_outputs(4347) <= not b;
    layer4_outputs(4348) <= not a or b;
    layer4_outputs(4349) <= a and not b;
    layer4_outputs(4350) <= not b;
    layer4_outputs(4351) <= not a;
    layer4_outputs(4352) <= b;
    layer4_outputs(4353) <= not (a or b);
    layer4_outputs(4354) <= a;
    layer4_outputs(4355) <= a xor b;
    layer4_outputs(4356) <= not a or b;
    layer4_outputs(4357) <= not b;
    layer4_outputs(4358) <= not (a or b);
    layer4_outputs(4359) <= not a;
    layer4_outputs(4360) <= not (a and b);
    layer4_outputs(4361) <= a xor b;
    layer4_outputs(4362) <= a;
    layer4_outputs(4363) <= not a;
    layer4_outputs(4364) <= a;
    layer4_outputs(4365) <= not a;
    layer4_outputs(4366) <= a xor b;
    layer4_outputs(4367) <= not a;
    layer4_outputs(4368) <= not b;
    layer4_outputs(4369) <= not (a xor b);
    layer4_outputs(4370) <= a;
    layer4_outputs(4371) <= not b;
    layer4_outputs(4372) <= a and not b;
    layer4_outputs(4373) <= a or b;
    layer4_outputs(4374) <= not b;
    layer4_outputs(4375) <= not (a and b);
    layer4_outputs(4376) <= a xor b;
    layer4_outputs(4377) <= b;
    layer4_outputs(4378) <= not b;
    layer4_outputs(4379) <= not b;
    layer4_outputs(4380) <= a xor b;
    layer4_outputs(4381) <= a;
    layer4_outputs(4382) <= not a;
    layer4_outputs(4383) <= b;
    layer4_outputs(4384) <= not (a xor b);
    layer4_outputs(4385) <= not a;
    layer4_outputs(4386) <= not (a and b);
    layer4_outputs(4387) <= not a;
    layer4_outputs(4388) <= b and not a;
    layer4_outputs(4389) <= b and not a;
    layer4_outputs(4390) <= not a or b;
    layer4_outputs(4391) <= b;
    layer4_outputs(4392) <= b;
    layer4_outputs(4393) <= not b;
    layer4_outputs(4394) <= a xor b;
    layer4_outputs(4395) <= a xor b;
    layer4_outputs(4396) <= not b;
    layer4_outputs(4397) <= a;
    layer4_outputs(4398) <= a and not b;
    layer4_outputs(4399) <= not (a or b);
    layer4_outputs(4400) <= a xor b;
    layer4_outputs(4401) <= b;
    layer4_outputs(4402) <= b and not a;
    layer4_outputs(4403) <= not a;
    layer4_outputs(4404) <= a xor b;
    layer4_outputs(4405) <= not a;
    layer4_outputs(4406) <= not (a xor b);
    layer4_outputs(4407) <= b;
    layer4_outputs(4408) <= a;
    layer4_outputs(4409) <= b;
    layer4_outputs(4410) <= a and not b;
    layer4_outputs(4411) <= a;
    layer4_outputs(4412) <= not a or b;
    layer4_outputs(4413) <= a or b;
    layer4_outputs(4414) <= a and not b;
    layer4_outputs(4415) <= not a;
    layer4_outputs(4416) <= not b or a;
    layer4_outputs(4417) <= a xor b;
    layer4_outputs(4418) <= b and not a;
    layer4_outputs(4419) <= b;
    layer4_outputs(4420) <= a;
    layer4_outputs(4421) <= b;
    layer4_outputs(4422) <= not (a or b);
    layer4_outputs(4423) <= a;
    layer4_outputs(4424) <= not a or b;
    layer4_outputs(4425) <= not b;
    layer4_outputs(4426) <= a or b;
    layer4_outputs(4427) <= not a;
    layer4_outputs(4428) <= not b;
    layer4_outputs(4429) <= b;
    layer4_outputs(4430) <= not a;
    layer4_outputs(4431) <= a;
    layer4_outputs(4432) <= b and not a;
    layer4_outputs(4433) <= b;
    layer4_outputs(4434) <= a and not b;
    layer4_outputs(4435) <= b and not a;
    layer4_outputs(4436) <= not b or a;
    layer4_outputs(4437) <= a or b;
    layer4_outputs(4438) <= not (a xor b);
    layer4_outputs(4439) <= not a or b;
    layer4_outputs(4440) <= a xor b;
    layer4_outputs(4441) <= a;
    layer4_outputs(4442) <= a;
    layer4_outputs(4443) <= not (a or b);
    layer4_outputs(4444) <= a and b;
    layer4_outputs(4445) <= not b or a;
    layer4_outputs(4446) <= b;
    layer4_outputs(4447) <= a or b;
    layer4_outputs(4448) <= a or b;
    layer4_outputs(4449) <= b;
    layer4_outputs(4450) <= b;
    layer4_outputs(4451) <= a xor b;
    layer4_outputs(4452) <= a;
    layer4_outputs(4453) <= a;
    layer4_outputs(4454) <= not a;
    layer4_outputs(4455) <= not a or b;
    layer4_outputs(4456) <= a or b;
    layer4_outputs(4457) <= b;
    layer4_outputs(4458) <= a xor b;
    layer4_outputs(4459) <= not (a xor b);
    layer4_outputs(4460) <= b and not a;
    layer4_outputs(4461) <= 1'b0;
    layer4_outputs(4462) <= a and b;
    layer4_outputs(4463) <= a and b;
    layer4_outputs(4464) <= a;
    layer4_outputs(4465) <= not a or b;
    layer4_outputs(4466) <= not a or b;
    layer4_outputs(4467) <= not (a xor b);
    layer4_outputs(4468) <= a xor b;
    layer4_outputs(4469) <= not a or b;
    layer4_outputs(4470) <= a or b;
    layer4_outputs(4471) <= not a;
    layer4_outputs(4472) <= not a;
    layer4_outputs(4473) <= not b;
    layer4_outputs(4474) <= a;
    layer4_outputs(4475) <= a and b;
    layer4_outputs(4476) <= a and b;
    layer4_outputs(4477) <= not a;
    layer4_outputs(4478) <= a;
    layer4_outputs(4479) <= not (a and b);
    layer4_outputs(4480) <= not b;
    layer4_outputs(4481) <= not b;
    layer4_outputs(4482) <= not a;
    layer4_outputs(4483) <= not b;
    layer4_outputs(4484) <= not (a and b);
    layer4_outputs(4485) <= not a;
    layer4_outputs(4486) <= not (a or b);
    layer4_outputs(4487) <= a;
    layer4_outputs(4488) <= not b or a;
    layer4_outputs(4489) <= not (a xor b);
    layer4_outputs(4490) <= not (a and b);
    layer4_outputs(4491) <= not a;
    layer4_outputs(4492) <= b;
    layer4_outputs(4493) <= not (a and b);
    layer4_outputs(4494) <= not b;
    layer4_outputs(4495) <= b and not a;
    layer4_outputs(4496) <= not a;
    layer4_outputs(4497) <= a xor b;
    layer4_outputs(4498) <= b;
    layer4_outputs(4499) <= not (a or b);
    layer4_outputs(4500) <= a and not b;
    layer4_outputs(4501) <= a xor b;
    layer4_outputs(4502) <= not b or a;
    layer4_outputs(4503) <= a and not b;
    layer4_outputs(4504) <= not b;
    layer4_outputs(4505) <= a and not b;
    layer4_outputs(4506) <= b and not a;
    layer4_outputs(4507) <= b and not a;
    layer4_outputs(4508) <= not (a and b);
    layer4_outputs(4509) <= a and not b;
    layer4_outputs(4510) <= not (a xor b);
    layer4_outputs(4511) <= a xor b;
    layer4_outputs(4512) <= not (a and b);
    layer4_outputs(4513) <= a;
    layer4_outputs(4514) <= not (a xor b);
    layer4_outputs(4515) <= not (a and b);
    layer4_outputs(4516) <= not (a and b);
    layer4_outputs(4517) <= a xor b;
    layer4_outputs(4518) <= a;
    layer4_outputs(4519) <= not (a and b);
    layer4_outputs(4520) <= not a;
    layer4_outputs(4521) <= b and not a;
    layer4_outputs(4522) <= a xor b;
    layer4_outputs(4523) <= not (a or b);
    layer4_outputs(4524) <= not (a xor b);
    layer4_outputs(4525) <= not (a xor b);
    layer4_outputs(4526) <= not (a xor b);
    layer4_outputs(4527) <= not a;
    layer4_outputs(4528) <= a xor b;
    layer4_outputs(4529) <= not b;
    layer4_outputs(4530) <= not a or b;
    layer4_outputs(4531) <= not (a and b);
    layer4_outputs(4532) <= a xor b;
    layer4_outputs(4533) <= not b or a;
    layer4_outputs(4534) <= a;
    layer4_outputs(4535) <= not a;
    layer4_outputs(4536) <= not a;
    layer4_outputs(4537) <= not (a xor b);
    layer4_outputs(4538) <= not b;
    layer4_outputs(4539) <= not (a or b);
    layer4_outputs(4540) <= not (a xor b);
    layer4_outputs(4541) <= not (a or b);
    layer4_outputs(4542) <= b;
    layer4_outputs(4543) <= not b;
    layer4_outputs(4544) <= not (a xor b);
    layer4_outputs(4545) <= not a or b;
    layer4_outputs(4546) <= a;
    layer4_outputs(4547) <= a xor b;
    layer4_outputs(4548) <= not a;
    layer4_outputs(4549) <= a;
    layer4_outputs(4550) <= not b or a;
    layer4_outputs(4551) <= not a;
    layer4_outputs(4552) <= b;
    layer4_outputs(4553) <= b;
    layer4_outputs(4554) <= not (a xor b);
    layer4_outputs(4555) <= not a;
    layer4_outputs(4556) <= not b;
    layer4_outputs(4557) <= not a;
    layer4_outputs(4558) <= b;
    layer4_outputs(4559) <= not a;
    layer4_outputs(4560) <= not (a or b);
    layer4_outputs(4561) <= b;
    layer4_outputs(4562) <= not (a and b);
    layer4_outputs(4563) <= b;
    layer4_outputs(4564) <= a xor b;
    layer4_outputs(4565) <= not a or b;
    layer4_outputs(4566) <= not a;
    layer4_outputs(4567) <= not (a xor b);
    layer4_outputs(4568) <= a and not b;
    layer4_outputs(4569) <= a or b;
    layer4_outputs(4570) <= b and not a;
    layer4_outputs(4571) <= a;
    layer4_outputs(4572) <= not b;
    layer4_outputs(4573) <= not b;
    layer4_outputs(4574) <= b;
    layer4_outputs(4575) <= a xor b;
    layer4_outputs(4576) <= b;
    layer4_outputs(4577) <= a xor b;
    layer4_outputs(4578) <= a xor b;
    layer4_outputs(4579) <= not b;
    layer4_outputs(4580) <= a and b;
    layer4_outputs(4581) <= a and not b;
    layer4_outputs(4582) <= b;
    layer4_outputs(4583) <= not b;
    layer4_outputs(4584) <= not b or a;
    layer4_outputs(4585) <= a or b;
    layer4_outputs(4586) <= not (a xor b);
    layer4_outputs(4587) <= a xor b;
    layer4_outputs(4588) <= not a;
    layer4_outputs(4589) <= a and not b;
    layer4_outputs(4590) <= a or b;
    layer4_outputs(4591) <= a and not b;
    layer4_outputs(4592) <= not b;
    layer4_outputs(4593) <= a xor b;
    layer4_outputs(4594) <= a and not b;
    layer4_outputs(4595) <= a and b;
    layer4_outputs(4596) <= a and b;
    layer4_outputs(4597) <= a;
    layer4_outputs(4598) <= not a;
    layer4_outputs(4599) <= a xor b;
    layer4_outputs(4600) <= not (a and b);
    layer4_outputs(4601) <= not (a xor b);
    layer4_outputs(4602) <= a and not b;
    layer4_outputs(4603) <= not b;
    layer4_outputs(4604) <= a xor b;
    layer4_outputs(4605) <= a;
    layer4_outputs(4606) <= b and not a;
    layer4_outputs(4607) <= not a;
    layer4_outputs(4608) <= b;
    layer4_outputs(4609) <= a or b;
    layer4_outputs(4610) <= not (a xor b);
    layer4_outputs(4611) <= not (a xor b);
    layer4_outputs(4612) <= not a;
    layer4_outputs(4613) <= not (a xor b);
    layer4_outputs(4614) <= a;
    layer4_outputs(4615) <= a or b;
    layer4_outputs(4616) <= a xor b;
    layer4_outputs(4617) <= b;
    layer4_outputs(4618) <= not (a xor b);
    layer4_outputs(4619) <= a;
    layer4_outputs(4620) <= not b;
    layer4_outputs(4621) <= a;
    layer4_outputs(4622) <= not b;
    layer4_outputs(4623) <= not b or a;
    layer4_outputs(4624) <= a;
    layer4_outputs(4625) <= a;
    layer4_outputs(4626) <= not (a xor b);
    layer4_outputs(4627) <= a and b;
    layer4_outputs(4628) <= not (a or b);
    layer4_outputs(4629) <= not (a xor b);
    layer4_outputs(4630) <= a or b;
    layer4_outputs(4631) <= not (a or b);
    layer4_outputs(4632) <= not a;
    layer4_outputs(4633) <= b;
    layer4_outputs(4634) <= not a;
    layer4_outputs(4635) <= not a;
    layer4_outputs(4636) <= a xor b;
    layer4_outputs(4637) <= not (a xor b);
    layer4_outputs(4638) <= a and b;
    layer4_outputs(4639) <= b;
    layer4_outputs(4640) <= not b or a;
    layer4_outputs(4641) <= a or b;
    layer4_outputs(4642) <= a;
    layer4_outputs(4643) <= b;
    layer4_outputs(4644) <= not a or b;
    layer4_outputs(4645) <= a;
    layer4_outputs(4646) <= b and not a;
    layer4_outputs(4647) <= a and not b;
    layer4_outputs(4648) <= not (a xor b);
    layer4_outputs(4649) <= not b;
    layer4_outputs(4650) <= not (a xor b);
    layer4_outputs(4651) <= not a;
    layer4_outputs(4652) <= not b;
    layer4_outputs(4653) <= not b;
    layer4_outputs(4654) <= not b;
    layer4_outputs(4655) <= 1'b1;
    layer4_outputs(4656) <= a or b;
    layer4_outputs(4657) <= a;
    layer4_outputs(4658) <= not a;
    layer4_outputs(4659) <= b and not a;
    layer4_outputs(4660) <= not a or b;
    layer4_outputs(4661) <= a xor b;
    layer4_outputs(4662) <= a;
    layer4_outputs(4663) <= a xor b;
    layer4_outputs(4664) <= b;
    layer4_outputs(4665) <= a and b;
    layer4_outputs(4666) <= a and not b;
    layer4_outputs(4667) <= a xor b;
    layer4_outputs(4668) <= a;
    layer4_outputs(4669) <= b and not a;
    layer4_outputs(4670) <= a;
    layer4_outputs(4671) <= not (a or b);
    layer4_outputs(4672) <= a;
    layer4_outputs(4673) <= b and not a;
    layer4_outputs(4674) <= not (a or b);
    layer4_outputs(4675) <= b;
    layer4_outputs(4676) <= b and not a;
    layer4_outputs(4677) <= a and not b;
    layer4_outputs(4678) <= not b;
    layer4_outputs(4679) <= b;
    layer4_outputs(4680) <= not b;
    layer4_outputs(4681) <= a and not b;
    layer4_outputs(4682) <= not b;
    layer4_outputs(4683) <= a xor b;
    layer4_outputs(4684) <= not a or b;
    layer4_outputs(4685) <= a and b;
    layer4_outputs(4686) <= not (a and b);
    layer4_outputs(4687) <= not b or a;
    layer4_outputs(4688) <= not (a and b);
    layer4_outputs(4689) <= not (a or b);
    layer4_outputs(4690) <= not a;
    layer4_outputs(4691) <= not a;
    layer4_outputs(4692) <= b;
    layer4_outputs(4693) <= a and not b;
    layer4_outputs(4694) <= not (a or b);
    layer4_outputs(4695) <= not b or a;
    layer4_outputs(4696) <= b and not a;
    layer4_outputs(4697) <= b;
    layer4_outputs(4698) <= not a or b;
    layer4_outputs(4699) <= a or b;
    layer4_outputs(4700) <= a xor b;
    layer4_outputs(4701) <= not b;
    layer4_outputs(4702) <= not (a xor b);
    layer4_outputs(4703) <= a xor b;
    layer4_outputs(4704) <= not (a xor b);
    layer4_outputs(4705) <= a and b;
    layer4_outputs(4706) <= not a;
    layer4_outputs(4707) <= b and not a;
    layer4_outputs(4708) <= 1'b0;
    layer4_outputs(4709) <= a xor b;
    layer4_outputs(4710) <= a;
    layer4_outputs(4711) <= b and not a;
    layer4_outputs(4712) <= not a or b;
    layer4_outputs(4713) <= not a;
    layer4_outputs(4714) <= b;
    layer4_outputs(4715) <= not b;
    layer4_outputs(4716) <= a;
    layer4_outputs(4717) <= not (a and b);
    layer4_outputs(4718) <= not (a and b);
    layer4_outputs(4719) <= not (a xor b);
    layer4_outputs(4720) <= not b;
    layer4_outputs(4721) <= not a;
    layer4_outputs(4722) <= a;
    layer4_outputs(4723) <= a xor b;
    layer4_outputs(4724) <= b;
    layer4_outputs(4725) <= not (a and b);
    layer4_outputs(4726) <= a xor b;
    layer4_outputs(4727) <= a or b;
    layer4_outputs(4728) <= not (a and b);
    layer4_outputs(4729) <= not (a and b);
    layer4_outputs(4730) <= a xor b;
    layer4_outputs(4731) <= not a or b;
    layer4_outputs(4732) <= a and not b;
    layer4_outputs(4733) <= not a or b;
    layer4_outputs(4734) <= not (a xor b);
    layer4_outputs(4735) <= a;
    layer4_outputs(4736) <= a and b;
    layer4_outputs(4737) <= not a or b;
    layer4_outputs(4738) <= a xor b;
    layer4_outputs(4739) <= not b;
    layer4_outputs(4740) <= not (a and b);
    layer4_outputs(4741) <= not (a or b);
    layer4_outputs(4742) <= not b or a;
    layer4_outputs(4743) <= not a;
    layer4_outputs(4744) <= not (a xor b);
    layer4_outputs(4745) <= not (a xor b);
    layer4_outputs(4746) <= a;
    layer4_outputs(4747) <= b and not a;
    layer4_outputs(4748) <= a xor b;
    layer4_outputs(4749) <= not (a xor b);
    layer4_outputs(4750) <= not a;
    layer4_outputs(4751) <= b;
    layer4_outputs(4752) <= b and not a;
    layer4_outputs(4753) <= a;
    layer4_outputs(4754) <= not a;
    layer4_outputs(4755) <= a;
    layer4_outputs(4756) <= b;
    layer4_outputs(4757) <= a;
    layer4_outputs(4758) <= b;
    layer4_outputs(4759) <= not b;
    layer4_outputs(4760) <= b;
    layer4_outputs(4761) <= not (a or b);
    layer4_outputs(4762) <= a xor b;
    layer4_outputs(4763) <= a or b;
    layer4_outputs(4764) <= a xor b;
    layer4_outputs(4765) <= not a;
    layer4_outputs(4766) <= a;
    layer4_outputs(4767) <= a xor b;
    layer4_outputs(4768) <= a xor b;
    layer4_outputs(4769) <= a and not b;
    layer4_outputs(4770) <= not b;
    layer4_outputs(4771) <= not b;
    layer4_outputs(4772) <= not b;
    layer4_outputs(4773) <= not b;
    layer4_outputs(4774) <= b;
    layer4_outputs(4775) <= not (a and b);
    layer4_outputs(4776) <= not b or a;
    layer4_outputs(4777) <= a xor b;
    layer4_outputs(4778) <= not b;
    layer4_outputs(4779) <= a;
    layer4_outputs(4780) <= a and not b;
    layer4_outputs(4781) <= b;
    layer4_outputs(4782) <= not a;
    layer4_outputs(4783) <= a and not b;
    layer4_outputs(4784) <= a or b;
    layer4_outputs(4785) <= a;
    layer4_outputs(4786) <= a;
    layer4_outputs(4787) <= not (a xor b);
    layer4_outputs(4788) <= b and not a;
    layer4_outputs(4789) <= a;
    layer4_outputs(4790) <= not (a or b);
    layer4_outputs(4791) <= not a or b;
    layer4_outputs(4792) <= a;
    layer4_outputs(4793) <= not b or a;
    layer4_outputs(4794) <= not b or a;
    layer4_outputs(4795) <= not (a or b);
    layer4_outputs(4796) <= b;
    layer4_outputs(4797) <= a;
    layer4_outputs(4798) <= not a;
    layer4_outputs(4799) <= not b;
    layer4_outputs(4800) <= b;
    layer4_outputs(4801) <= a and not b;
    layer4_outputs(4802) <= not a;
    layer4_outputs(4803) <= a or b;
    layer4_outputs(4804) <= b;
    layer4_outputs(4805) <= not b or a;
    layer4_outputs(4806) <= not b;
    layer4_outputs(4807) <= not a;
    layer4_outputs(4808) <= not a;
    layer4_outputs(4809) <= 1'b0;
    layer4_outputs(4810) <= a;
    layer4_outputs(4811) <= not b;
    layer4_outputs(4812) <= not (a xor b);
    layer4_outputs(4813) <= a xor b;
    layer4_outputs(4814) <= b and not a;
    layer4_outputs(4815) <= a;
    layer4_outputs(4816) <= not (a and b);
    layer4_outputs(4817) <= a and b;
    layer4_outputs(4818) <= not (a xor b);
    layer4_outputs(4819) <= a xor b;
    layer4_outputs(4820) <= not (a and b);
    layer4_outputs(4821) <= not a;
    layer4_outputs(4822) <= not a;
    layer4_outputs(4823) <= a or b;
    layer4_outputs(4824) <= a or b;
    layer4_outputs(4825) <= a and b;
    layer4_outputs(4826) <= not b;
    layer4_outputs(4827) <= not b;
    layer4_outputs(4828) <= not (a or b);
    layer4_outputs(4829) <= not (a xor b);
    layer4_outputs(4830) <= a xor b;
    layer4_outputs(4831) <= not a or b;
    layer4_outputs(4832) <= not a or b;
    layer4_outputs(4833) <= not b;
    layer4_outputs(4834) <= not (a and b);
    layer4_outputs(4835) <= not b;
    layer4_outputs(4836) <= a;
    layer4_outputs(4837) <= a;
    layer4_outputs(4838) <= not b;
    layer4_outputs(4839) <= a and not b;
    layer4_outputs(4840) <= not a;
    layer4_outputs(4841) <= not (a xor b);
    layer4_outputs(4842) <= not b;
    layer4_outputs(4843) <= not b or a;
    layer4_outputs(4844) <= a xor b;
    layer4_outputs(4845) <= not a;
    layer4_outputs(4846) <= a;
    layer4_outputs(4847) <= a or b;
    layer4_outputs(4848) <= b and not a;
    layer4_outputs(4849) <= not a;
    layer4_outputs(4850) <= not (a and b);
    layer4_outputs(4851) <= not b;
    layer4_outputs(4852) <= not a;
    layer4_outputs(4853) <= a;
    layer4_outputs(4854) <= not b;
    layer4_outputs(4855) <= a;
    layer4_outputs(4856) <= a;
    layer4_outputs(4857) <= not a;
    layer4_outputs(4858) <= a or b;
    layer4_outputs(4859) <= a;
    layer4_outputs(4860) <= b;
    layer4_outputs(4861) <= a;
    layer4_outputs(4862) <= not a;
    layer4_outputs(4863) <= not b;
    layer4_outputs(4864) <= b and not a;
    layer4_outputs(4865) <= b and not a;
    layer4_outputs(4866) <= not b;
    layer4_outputs(4867) <= not b or a;
    layer4_outputs(4868) <= b and not a;
    layer4_outputs(4869) <= not b;
    layer4_outputs(4870) <= b;
    layer4_outputs(4871) <= b;
    layer4_outputs(4872) <= not (a and b);
    layer4_outputs(4873) <= b;
    layer4_outputs(4874) <= not b;
    layer4_outputs(4875) <= 1'b0;
    layer4_outputs(4876) <= a;
    layer4_outputs(4877) <= not (a and b);
    layer4_outputs(4878) <= not (a xor b);
    layer4_outputs(4879) <= not (a or b);
    layer4_outputs(4880) <= a;
    layer4_outputs(4881) <= not b;
    layer4_outputs(4882) <= not a or b;
    layer4_outputs(4883) <= not b;
    layer4_outputs(4884) <= a or b;
    layer4_outputs(4885) <= a xor b;
    layer4_outputs(4886) <= b;
    layer4_outputs(4887) <= not (a xor b);
    layer4_outputs(4888) <= a;
    layer4_outputs(4889) <= not b or a;
    layer4_outputs(4890) <= not b or a;
    layer4_outputs(4891) <= not a;
    layer4_outputs(4892) <= not a or b;
    layer4_outputs(4893) <= not b;
    layer4_outputs(4894) <= b;
    layer4_outputs(4895) <= not a;
    layer4_outputs(4896) <= not b;
    layer4_outputs(4897) <= a or b;
    layer4_outputs(4898) <= a xor b;
    layer4_outputs(4899) <= a xor b;
    layer4_outputs(4900) <= not (a and b);
    layer4_outputs(4901) <= not a or b;
    layer4_outputs(4902) <= b and not a;
    layer4_outputs(4903) <= a xor b;
    layer4_outputs(4904) <= not b or a;
    layer4_outputs(4905) <= a and b;
    layer4_outputs(4906) <= not (a or b);
    layer4_outputs(4907) <= a;
    layer4_outputs(4908) <= not (a xor b);
    layer4_outputs(4909) <= not a or b;
    layer4_outputs(4910) <= not (a or b);
    layer4_outputs(4911) <= not a or b;
    layer4_outputs(4912) <= not (a or b);
    layer4_outputs(4913) <= b;
    layer4_outputs(4914) <= b;
    layer4_outputs(4915) <= a and b;
    layer4_outputs(4916) <= not b;
    layer4_outputs(4917) <= b and not a;
    layer4_outputs(4918) <= b;
    layer4_outputs(4919) <= not (a and b);
    layer4_outputs(4920) <= a xor b;
    layer4_outputs(4921) <= not a;
    layer4_outputs(4922) <= a or b;
    layer4_outputs(4923) <= not a or b;
    layer4_outputs(4924) <= b;
    layer4_outputs(4925) <= not b;
    layer4_outputs(4926) <= not b;
    layer4_outputs(4927) <= not (a or b);
    layer4_outputs(4928) <= not (a or b);
    layer4_outputs(4929) <= not a or b;
    layer4_outputs(4930) <= not a or b;
    layer4_outputs(4931) <= not (a or b);
    layer4_outputs(4932) <= not (a xor b);
    layer4_outputs(4933) <= a xor b;
    layer4_outputs(4934) <= a xor b;
    layer4_outputs(4935) <= b;
    layer4_outputs(4936) <= a and b;
    layer4_outputs(4937) <= a xor b;
    layer4_outputs(4938) <= a;
    layer4_outputs(4939) <= not (a and b);
    layer4_outputs(4940) <= not (a or b);
    layer4_outputs(4941) <= a xor b;
    layer4_outputs(4942) <= not a or b;
    layer4_outputs(4943) <= a;
    layer4_outputs(4944) <= not a;
    layer4_outputs(4945) <= a and b;
    layer4_outputs(4946) <= not (a xor b);
    layer4_outputs(4947) <= a;
    layer4_outputs(4948) <= not (a or b);
    layer4_outputs(4949) <= not b;
    layer4_outputs(4950) <= a xor b;
    layer4_outputs(4951) <= not a;
    layer4_outputs(4952) <= a and b;
    layer4_outputs(4953) <= b;
    layer4_outputs(4954) <= b and not a;
    layer4_outputs(4955) <= b;
    layer4_outputs(4956) <= not (a and b);
    layer4_outputs(4957) <= b;
    layer4_outputs(4958) <= not b;
    layer4_outputs(4959) <= not a;
    layer4_outputs(4960) <= a and b;
    layer4_outputs(4961) <= not (a or b);
    layer4_outputs(4962) <= not a or b;
    layer4_outputs(4963) <= b;
    layer4_outputs(4964) <= a xor b;
    layer4_outputs(4965) <= b and not a;
    layer4_outputs(4966) <= a xor b;
    layer4_outputs(4967) <= a;
    layer4_outputs(4968) <= not (a or b);
    layer4_outputs(4969) <= not b or a;
    layer4_outputs(4970) <= a and b;
    layer4_outputs(4971) <= not b;
    layer4_outputs(4972) <= b;
    layer4_outputs(4973) <= b and not a;
    layer4_outputs(4974) <= a;
    layer4_outputs(4975) <= not a or b;
    layer4_outputs(4976) <= not b or a;
    layer4_outputs(4977) <= not b;
    layer4_outputs(4978) <= not b or a;
    layer4_outputs(4979) <= not (a and b);
    layer4_outputs(4980) <= b;
    layer4_outputs(4981) <= not a;
    layer4_outputs(4982) <= b and not a;
    layer4_outputs(4983) <= a xor b;
    layer4_outputs(4984) <= not (a xor b);
    layer4_outputs(4985) <= not (a xor b);
    layer4_outputs(4986) <= not (a xor b);
    layer4_outputs(4987) <= not (a xor b);
    layer4_outputs(4988) <= a;
    layer4_outputs(4989) <= not a or b;
    layer4_outputs(4990) <= not (a and b);
    layer4_outputs(4991) <= a;
    layer4_outputs(4992) <= not a;
    layer4_outputs(4993) <= not a;
    layer4_outputs(4994) <= a and b;
    layer4_outputs(4995) <= not b;
    layer4_outputs(4996) <= b;
    layer4_outputs(4997) <= a;
    layer4_outputs(4998) <= a and b;
    layer4_outputs(4999) <= not (a or b);
    layer4_outputs(5000) <= a or b;
    layer4_outputs(5001) <= b and not a;
    layer4_outputs(5002) <= b;
    layer4_outputs(5003) <= not (a and b);
    layer4_outputs(5004) <= a and b;
    layer4_outputs(5005) <= not (a xor b);
    layer4_outputs(5006) <= not a;
    layer4_outputs(5007) <= a xor b;
    layer4_outputs(5008) <= not (a xor b);
    layer4_outputs(5009) <= a and b;
    layer4_outputs(5010) <= b;
    layer4_outputs(5011) <= b;
    layer4_outputs(5012) <= a xor b;
    layer4_outputs(5013) <= a and not b;
    layer4_outputs(5014) <= not (a xor b);
    layer4_outputs(5015) <= a xor b;
    layer4_outputs(5016) <= b and not a;
    layer4_outputs(5017) <= not a;
    layer4_outputs(5018) <= not (a xor b);
    layer4_outputs(5019) <= not b or a;
    layer4_outputs(5020) <= a or b;
    layer4_outputs(5021) <= not a;
    layer4_outputs(5022) <= b and not a;
    layer4_outputs(5023) <= not (a and b);
    layer4_outputs(5024) <= not b or a;
    layer4_outputs(5025) <= b;
    layer4_outputs(5026) <= not b;
    layer4_outputs(5027) <= not a;
    layer4_outputs(5028) <= a and not b;
    layer4_outputs(5029) <= not (a and b);
    layer4_outputs(5030) <= not a;
    layer4_outputs(5031) <= a xor b;
    layer4_outputs(5032) <= a xor b;
    layer4_outputs(5033) <= not b;
    layer4_outputs(5034) <= not (a and b);
    layer4_outputs(5035) <= b;
    layer4_outputs(5036) <= a or b;
    layer4_outputs(5037) <= not b or a;
    layer4_outputs(5038) <= not a;
    layer4_outputs(5039) <= a;
    layer4_outputs(5040) <= not b;
    layer4_outputs(5041) <= not b;
    layer4_outputs(5042) <= not b;
    layer4_outputs(5043) <= a and b;
    layer4_outputs(5044) <= b;
    layer4_outputs(5045) <= a;
    layer4_outputs(5046) <= not (a and b);
    layer4_outputs(5047) <= a and b;
    layer4_outputs(5048) <= not (a or b);
    layer4_outputs(5049) <= a and not b;
    layer4_outputs(5050) <= a and b;
    layer4_outputs(5051) <= a;
    layer4_outputs(5052) <= not b;
    layer4_outputs(5053) <= a and not b;
    layer4_outputs(5054) <= not a;
    layer4_outputs(5055) <= a and not b;
    layer4_outputs(5056) <= not a or b;
    layer4_outputs(5057) <= b and not a;
    layer4_outputs(5058) <= not a;
    layer4_outputs(5059) <= b;
    layer4_outputs(5060) <= a;
    layer4_outputs(5061) <= a xor b;
    layer4_outputs(5062) <= b and not a;
    layer4_outputs(5063) <= a and b;
    layer4_outputs(5064) <= not a;
    layer4_outputs(5065) <= not (a or b);
    layer4_outputs(5066) <= a;
    layer4_outputs(5067) <= not b;
    layer4_outputs(5068) <= a xor b;
    layer4_outputs(5069) <= b;
    layer4_outputs(5070) <= a xor b;
    layer4_outputs(5071) <= a xor b;
    layer4_outputs(5072) <= not a or b;
    layer4_outputs(5073) <= not (a xor b);
    layer4_outputs(5074) <= not b;
    layer4_outputs(5075) <= b;
    layer4_outputs(5076) <= not (a xor b);
    layer4_outputs(5077) <= not a or b;
    layer4_outputs(5078) <= b;
    layer4_outputs(5079) <= a and not b;
    layer4_outputs(5080) <= a;
    layer4_outputs(5081) <= a or b;
    layer4_outputs(5082) <= a and not b;
    layer4_outputs(5083) <= not b;
    layer4_outputs(5084) <= b and not a;
    layer4_outputs(5085) <= a;
    layer4_outputs(5086) <= a xor b;
    layer4_outputs(5087) <= a;
    layer4_outputs(5088) <= not (a and b);
    layer4_outputs(5089) <= a and b;
    layer4_outputs(5090) <= not b or a;
    layer4_outputs(5091) <= not (a or b);
    layer4_outputs(5092) <= a xor b;
    layer4_outputs(5093) <= a and not b;
    layer4_outputs(5094) <= 1'b0;
    layer4_outputs(5095) <= not (a and b);
    layer4_outputs(5096) <= not (a or b);
    layer4_outputs(5097) <= a xor b;
    layer4_outputs(5098) <= not b;
    layer4_outputs(5099) <= not (a xor b);
    layer4_outputs(5100) <= not (a or b);
    layer4_outputs(5101) <= a;
    layer4_outputs(5102) <= not a;
    layer4_outputs(5103) <= b;
    layer4_outputs(5104) <= a and b;
    layer4_outputs(5105) <= not (a and b);
    layer4_outputs(5106) <= b;
    layer4_outputs(5107) <= not b;
    layer4_outputs(5108) <= a and not b;
    layer4_outputs(5109) <= not a or b;
    layer4_outputs(5110) <= not b;
    layer4_outputs(5111) <= not b;
    layer4_outputs(5112) <= a or b;
    layer4_outputs(5113) <= not (a xor b);
    layer4_outputs(5114) <= not a or b;
    layer4_outputs(5115) <= b;
    layer4_outputs(5116) <= not b;
    layer4_outputs(5117) <= not b or a;
    layer4_outputs(5118) <= not b or a;
    layer4_outputs(5119) <= b;
    layer4_outputs(5120) <= not b or a;
    layer4_outputs(5121) <= not b or a;
    layer4_outputs(5122) <= a and b;
    layer4_outputs(5123) <= b;
    layer4_outputs(5124) <= a and b;
    layer4_outputs(5125) <= a;
    layer4_outputs(5126) <= a and not b;
    layer4_outputs(5127) <= not a;
    layer4_outputs(5128) <= b;
    layer4_outputs(5129) <= a xor b;
    layer4_outputs(5130) <= not a;
    layer4_outputs(5131) <= b and not a;
    layer4_outputs(5132) <= a and not b;
    layer4_outputs(5133) <= a or b;
    layer4_outputs(5134) <= not a or b;
    layer4_outputs(5135) <= b;
    layer4_outputs(5136) <= not a;
    layer4_outputs(5137) <= b;
    layer4_outputs(5138) <= a and not b;
    layer4_outputs(5139) <= not (a xor b);
    layer4_outputs(5140) <= a and not b;
    layer4_outputs(5141) <= a and not b;
    layer4_outputs(5142) <= not b;
    layer4_outputs(5143) <= a xor b;
    layer4_outputs(5144) <= not b;
    layer4_outputs(5145) <= b;
    layer4_outputs(5146) <= not a or b;
    layer4_outputs(5147) <= a or b;
    layer4_outputs(5148) <= not (a xor b);
    layer4_outputs(5149) <= not a;
    layer4_outputs(5150) <= a xor b;
    layer4_outputs(5151) <= a;
    layer4_outputs(5152) <= a and not b;
    layer4_outputs(5153) <= b and not a;
    layer4_outputs(5154) <= not (a xor b);
    layer4_outputs(5155) <= not (a xor b);
    layer4_outputs(5156) <= not (a xor b);
    layer4_outputs(5157) <= a;
    layer4_outputs(5158) <= a xor b;
    layer4_outputs(5159) <= a or b;
    layer4_outputs(5160) <= a xor b;
    layer4_outputs(5161) <= not a;
    layer4_outputs(5162) <= a;
    layer4_outputs(5163) <= not a or b;
    layer4_outputs(5164) <= not (a xor b);
    layer4_outputs(5165) <= not b;
    layer4_outputs(5166) <= a and b;
    layer4_outputs(5167) <= not a;
    layer4_outputs(5168) <= a;
    layer4_outputs(5169) <= not b;
    layer4_outputs(5170) <= not a;
    layer4_outputs(5171) <= not (a and b);
    layer4_outputs(5172) <= not a;
    layer4_outputs(5173) <= not a;
    layer4_outputs(5174) <= not b;
    layer4_outputs(5175) <= b and not a;
    layer4_outputs(5176) <= b;
    layer4_outputs(5177) <= not b;
    layer4_outputs(5178) <= not (a and b);
    layer4_outputs(5179) <= a;
    layer4_outputs(5180) <= a;
    layer4_outputs(5181) <= not (a xor b);
    layer4_outputs(5182) <= a xor b;
    layer4_outputs(5183) <= not a;
    layer4_outputs(5184) <= not (a xor b);
    layer4_outputs(5185) <= not a or b;
    layer4_outputs(5186) <= not a;
    layer4_outputs(5187) <= not (a xor b);
    layer4_outputs(5188) <= not a;
    layer4_outputs(5189) <= b and not a;
    layer4_outputs(5190) <= a;
    layer4_outputs(5191) <= b;
    layer4_outputs(5192) <= not a;
    layer4_outputs(5193) <= a xor b;
    layer4_outputs(5194) <= not a;
    layer4_outputs(5195) <= a and b;
    layer4_outputs(5196) <= not b;
    layer4_outputs(5197) <= not a;
    layer4_outputs(5198) <= a or b;
    layer4_outputs(5199) <= b;
    layer4_outputs(5200) <= b;
    layer4_outputs(5201) <= a and not b;
    layer4_outputs(5202) <= not a;
    layer4_outputs(5203) <= a xor b;
    layer4_outputs(5204) <= not a;
    layer4_outputs(5205) <= not b;
    layer4_outputs(5206) <= a xor b;
    layer4_outputs(5207) <= a xor b;
    layer4_outputs(5208) <= a xor b;
    layer4_outputs(5209) <= b;
    layer4_outputs(5210) <= b;
    layer4_outputs(5211) <= a and b;
    layer4_outputs(5212) <= a xor b;
    layer4_outputs(5213) <= a;
    layer4_outputs(5214) <= a and b;
    layer4_outputs(5215) <= a or b;
    layer4_outputs(5216) <= not b;
    layer4_outputs(5217) <= not b;
    layer4_outputs(5218) <= b;
    layer4_outputs(5219) <= a or b;
    layer4_outputs(5220) <= not (a xor b);
    layer4_outputs(5221) <= not (a xor b);
    layer4_outputs(5222) <= not b;
    layer4_outputs(5223) <= not b or a;
    layer4_outputs(5224) <= b;
    layer4_outputs(5225) <= a xor b;
    layer4_outputs(5226) <= a and not b;
    layer4_outputs(5227) <= b;
    layer4_outputs(5228) <= not (a xor b);
    layer4_outputs(5229) <= a;
    layer4_outputs(5230) <= not a or b;
    layer4_outputs(5231) <= not b;
    layer4_outputs(5232) <= not b;
    layer4_outputs(5233) <= b;
    layer4_outputs(5234) <= b;
    layer4_outputs(5235) <= a;
    layer4_outputs(5236) <= not a;
    layer4_outputs(5237) <= b;
    layer4_outputs(5238) <= not (a or b);
    layer4_outputs(5239) <= not b;
    layer4_outputs(5240) <= a and b;
    layer4_outputs(5241) <= not (a and b);
    layer4_outputs(5242) <= a and b;
    layer4_outputs(5243) <= a;
    layer4_outputs(5244) <= not b or a;
    layer4_outputs(5245) <= a and not b;
    layer4_outputs(5246) <= a and not b;
    layer4_outputs(5247) <= not a;
    layer4_outputs(5248) <= b and not a;
    layer4_outputs(5249) <= a xor b;
    layer4_outputs(5250) <= b;
    layer4_outputs(5251) <= a and b;
    layer4_outputs(5252) <= not b;
    layer4_outputs(5253) <= a or b;
    layer4_outputs(5254) <= b;
    layer4_outputs(5255) <= not a;
    layer4_outputs(5256) <= b and not a;
    layer4_outputs(5257) <= not b;
    layer4_outputs(5258) <= a and b;
    layer4_outputs(5259) <= not b or a;
    layer4_outputs(5260) <= not a or b;
    layer4_outputs(5261) <= not a;
    layer4_outputs(5262) <= a;
    layer4_outputs(5263) <= a;
    layer4_outputs(5264) <= not (a or b);
    layer4_outputs(5265) <= b;
    layer4_outputs(5266) <= a;
    layer4_outputs(5267) <= not b or a;
    layer4_outputs(5268) <= not (a xor b);
    layer4_outputs(5269) <= a xor b;
    layer4_outputs(5270) <= not (a xor b);
    layer4_outputs(5271) <= a and not b;
    layer4_outputs(5272) <= a and not b;
    layer4_outputs(5273) <= a and b;
    layer4_outputs(5274) <= b;
    layer4_outputs(5275) <= not a;
    layer4_outputs(5276) <= not a or b;
    layer4_outputs(5277) <= not a;
    layer4_outputs(5278) <= not b;
    layer4_outputs(5279) <= not b;
    layer4_outputs(5280) <= a;
    layer4_outputs(5281) <= not (a or b);
    layer4_outputs(5282) <= not a;
    layer4_outputs(5283) <= b;
    layer4_outputs(5284) <= a and b;
    layer4_outputs(5285) <= not (a and b);
    layer4_outputs(5286) <= not (a and b);
    layer4_outputs(5287) <= not b;
    layer4_outputs(5288) <= b and not a;
    layer4_outputs(5289) <= not b;
    layer4_outputs(5290) <= a;
    layer4_outputs(5291) <= not (a xor b);
    layer4_outputs(5292) <= not a;
    layer4_outputs(5293) <= a or b;
    layer4_outputs(5294) <= not b or a;
    layer4_outputs(5295) <= not (a xor b);
    layer4_outputs(5296) <= not (a xor b);
    layer4_outputs(5297) <= a or b;
    layer4_outputs(5298) <= a and not b;
    layer4_outputs(5299) <= a;
    layer4_outputs(5300) <= not b or a;
    layer4_outputs(5301) <= a;
    layer4_outputs(5302) <= a xor b;
    layer4_outputs(5303) <= a or b;
    layer4_outputs(5304) <= a;
    layer4_outputs(5305) <= not b or a;
    layer4_outputs(5306) <= a;
    layer4_outputs(5307) <= not b;
    layer4_outputs(5308) <= not b or a;
    layer4_outputs(5309) <= a and not b;
    layer4_outputs(5310) <= not (a or b);
    layer4_outputs(5311) <= a xor b;
    layer4_outputs(5312) <= not (a xor b);
    layer4_outputs(5313) <= a and not b;
    layer4_outputs(5314) <= not b;
    layer4_outputs(5315) <= b and not a;
    layer4_outputs(5316) <= b and not a;
    layer4_outputs(5317) <= b;
    layer4_outputs(5318) <= a;
    layer4_outputs(5319) <= not a;
    layer4_outputs(5320) <= not a;
    layer4_outputs(5321) <= a or b;
    layer4_outputs(5322) <= not b or a;
    layer4_outputs(5323) <= a and not b;
    layer4_outputs(5324) <= a and not b;
    layer4_outputs(5325) <= a and not b;
    layer4_outputs(5326) <= a xor b;
    layer4_outputs(5327) <= not b or a;
    layer4_outputs(5328) <= not a;
    layer4_outputs(5329) <= a xor b;
    layer4_outputs(5330) <= not b;
    layer4_outputs(5331) <= b;
    layer4_outputs(5332) <= not a;
    layer4_outputs(5333) <= not (a or b);
    layer4_outputs(5334) <= not a or b;
    layer4_outputs(5335) <= b;
    layer4_outputs(5336) <= b and not a;
    layer4_outputs(5337) <= not a or b;
    layer4_outputs(5338) <= 1'b0;
    layer4_outputs(5339) <= not b or a;
    layer4_outputs(5340) <= a xor b;
    layer4_outputs(5341) <= not b;
    layer4_outputs(5342) <= not (a or b);
    layer4_outputs(5343) <= b;
    layer4_outputs(5344) <= b and not a;
    layer4_outputs(5345) <= not (a or b);
    layer4_outputs(5346) <= not b;
    layer4_outputs(5347) <= not a or b;
    layer4_outputs(5348) <= a;
    layer4_outputs(5349) <= a and b;
    layer4_outputs(5350) <= not a;
    layer4_outputs(5351) <= b;
    layer4_outputs(5352) <= a or b;
    layer4_outputs(5353) <= b;
    layer4_outputs(5354) <= a xor b;
    layer4_outputs(5355) <= b;
    layer4_outputs(5356) <= not (a xor b);
    layer4_outputs(5357) <= b and not a;
    layer4_outputs(5358) <= b;
    layer4_outputs(5359) <= a;
    layer4_outputs(5360) <= not (a or b);
    layer4_outputs(5361) <= a;
    layer4_outputs(5362) <= not a;
    layer4_outputs(5363) <= not (a and b);
    layer4_outputs(5364) <= b;
    layer4_outputs(5365) <= a xor b;
    layer4_outputs(5366) <= b and not a;
    layer4_outputs(5367) <= a xor b;
    layer4_outputs(5368) <= not (a and b);
    layer4_outputs(5369) <= not a;
    layer4_outputs(5370) <= not b;
    layer4_outputs(5371) <= not a;
    layer4_outputs(5372) <= not (a and b);
    layer4_outputs(5373) <= a;
    layer4_outputs(5374) <= a;
    layer4_outputs(5375) <= a;
    layer4_outputs(5376) <= not (a xor b);
    layer4_outputs(5377) <= not b or a;
    layer4_outputs(5378) <= a and not b;
    layer4_outputs(5379) <= not a;
    layer4_outputs(5380) <= not (a or b);
    layer4_outputs(5381) <= not (a xor b);
    layer4_outputs(5382) <= not b;
    layer4_outputs(5383) <= not (a xor b);
    layer4_outputs(5384) <= a or b;
    layer4_outputs(5385) <= not (a and b);
    layer4_outputs(5386) <= a;
    layer4_outputs(5387) <= a;
    layer4_outputs(5388) <= not b or a;
    layer4_outputs(5389) <= not b;
    layer4_outputs(5390) <= not (a xor b);
    layer4_outputs(5391) <= not a or b;
    layer4_outputs(5392) <= a;
    layer4_outputs(5393) <= b;
    layer4_outputs(5394) <= not b or a;
    layer4_outputs(5395) <= b;
    layer4_outputs(5396) <= not a;
    layer4_outputs(5397) <= not (a xor b);
    layer4_outputs(5398) <= a;
    layer4_outputs(5399) <= b;
    layer4_outputs(5400) <= not a;
    layer4_outputs(5401) <= a;
    layer4_outputs(5402) <= not b;
    layer4_outputs(5403) <= b;
    layer4_outputs(5404) <= not (a and b);
    layer4_outputs(5405) <= not (a or b);
    layer4_outputs(5406) <= b;
    layer4_outputs(5407) <= not b;
    layer4_outputs(5408) <= not a or b;
    layer4_outputs(5409) <= b;
    layer4_outputs(5410) <= a and not b;
    layer4_outputs(5411) <= b;
    layer4_outputs(5412) <= not a;
    layer4_outputs(5413) <= a xor b;
    layer4_outputs(5414) <= a;
    layer4_outputs(5415) <= a or b;
    layer4_outputs(5416) <= a;
    layer4_outputs(5417) <= not b;
    layer4_outputs(5418) <= not (a or b);
    layer4_outputs(5419) <= not b or a;
    layer4_outputs(5420) <= b and not a;
    layer4_outputs(5421) <= not a;
    layer4_outputs(5422) <= not b;
    layer4_outputs(5423) <= not a;
    layer4_outputs(5424) <= a xor b;
    layer4_outputs(5425) <= not b;
    layer4_outputs(5426) <= not (a xor b);
    layer4_outputs(5427) <= a and b;
    layer4_outputs(5428) <= not a;
    layer4_outputs(5429) <= not a;
    layer4_outputs(5430) <= a and not b;
    layer4_outputs(5431) <= b;
    layer4_outputs(5432) <= not b;
    layer4_outputs(5433) <= a;
    layer4_outputs(5434) <= not (a and b);
    layer4_outputs(5435) <= a;
    layer4_outputs(5436) <= b;
    layer4_outputs(5437) <= not a;
    layer4_outputs(5438) <= not a;
    layer4_outputs(5439) <= a or b;
    layer4_outputs(5440) <= not a;
    layer4_outputs(5441) <= a xor b;
    layer4_outputs(5442) <= not (a and b);
    layer4_outputs(5443) <= not a;
    layer4_outputs(5444) <= a and b;
    layer4_outputs(5445) <= not b or a;
    layer4_outputs(5446) <= not (a and b);
    layer4_outputs(5447) <= a;
    layer4_outputs(5448) <= not (a or b);
    layer4_outputs(5449) <= a;
    layer4_outputs(5450) <= b;
    layer4_outputs(5451) <= not a or b;
    layer4_outputs(5452) <= a;
    layer4_outputs(5453) <= not (a xor b);
    layer4_outputs(5454) <= b;
    layer4_outputs(5455) <= a;
    layer4_outputs(5456) <= not b;
    layer4_outputs(5457) <= a and not b;
    layer4_outputs(5458) <= not b;
    layer4_outputs(5459) <= b and not a;
    layer4_outputs(5460) <= not b;
    layer4_outputs(5461) <= a and b;
    layer4_outputs(5462) <= not (a xor b);
    layer4_outputs(5463) <= a or b;
    layer4_outputs(5464) <= a;
    layer4_outputs(5465) <= b;
    layer4_outputs(5466) <= b;
    layer4_outputs(5467) <= not (a xor b);
    layer4_outputs(5468) <= not b;
    layer4_outputs(5469) <= not a or b;
    layer4_outputs(5470) <= b;
    layer4_outputs(5471) <= not b;
    layer4_outputs(5472) <= b;
    layer4_outputs(5473) <= a;
    layer4_outputs(5474) <= not b;
    layer4_outputs(5475) <= not a;
    layer4_outputs(5476) <= not a;
    layer4_outputs(5477) <= not a or b;
    layer4_outputs(5478) <= not (a or b);
    layer4_outputs(5479) <= a xor b;
    layer4_outputs(5480) <= not (a xor b);
    layer4_outputs(5481) <= b;
    layer4_outputs(5482) <= not (a or b);
    layer4_outputs(5483) <= not b or a;
    layer4_outputs(5484) <= not b;
    layer4_outputs(5485) <= not a or b;
    layer4_outputs(5486) <= b;
    layer4_outputs(5487) <= a and not b;
    layer4_outputs(5488) <= b;
    layer4_outputs(5489) <= a or b;
    layer4_outputs(5490) <= a;
    layer4_outputs(5491) <= b;
    layer4_outputs(5492) <= not (a and b);
    layer4_outputs(5493) <= not a;
    layer4_outputs(5494) <= not b;
    layer4_outputs(5495) <= a and not b;
    layer4_outputs(5496) <= not b or a;
    layer4_outputs(5497) <= b and not a;
    layer4_outputs(5498) <= a;
    layer4_outputs(5499) <= not (a and b);
    layer4_outputs(5500) <= a;
    layer4_outputs(5501) <= b;
    layer4_outputs(5502) <= b;
    layer4_outputs(5503) <= b;
    layer4_outputs(5504) <= a xor b;
    layer4_outputs(5505) <= a and b;
    layer4_outputs(5506) <= a;
    layer4_outputs(5507) <= b;
    layer4_outputs(5508) <= a;
    layer4_outputs(5509) <= not b or a;
    layer4_outputs(5510) <= not a or b;
    layer4_outputs(5511) <= a or b;
    layer4_outputs(5512) <= a or b;
    layer4_outputs(5513) <= not (a xor b);
    layer4_outputs(5514) <= not a;
    layer4_outputs(5515) <= a xor b;
    layer4_outputs(5516) <= not b;
    layer4_outputs(5517) <= not a;
    layer4_outputs(5518) <= a and not b;
    layer4_outputs(5519) <= b and not a;
    layer4_outputs(5520) <= not (a xor b);
    layer4_outputs(5521) <= not (a or b);
    layer4_outputs(5522) <= a;
    layer4_outputs(5523) <= not b;
    layer4_outputs(5524) <= b and not a;
    layer4_outputs(5525) <= not (a xor b);
    layer4_outputs(5526) <= a and b;
    layer4_outputs(5527) <= not a;
    layer4_outputs(5528) <= not b;
    layer4_outputs(5529) <= a and b;
    layer4_outputs(5530) <= b;
    layer4_outputs(5531) <= a;
    layer4_outputs(5532) <= b and not a;
    layer4_outputs(5533) <= a or b;
    layer4_outputs(5534) <= not a;
    layer4_outputs(5535) <= not b;
    layer4_outputs(5536) <= a xor b;
    layer4_outputs(5537) <= not (a xor b);
    layer4_outputs(5538) <= b and not a;
    layer4_outputs(5539) <= not a;
    layer4_outputs(5540) <= not (a or b);
    layer4_outputs(5541) <= b;
    layer4_outputs(5542) <= b;
    layer4_outputs(5543) <= a xor b;
    layer4_outputs(5544) <= not b;
    layer4_outputs(5545) <= not b;
    layer4_outputs(5546) <= b;
    layer4_outputs(5547) <= not (a or b);
    layer4_outputs(5548) <= not a;
    layer4_outputs(5549) <= not b or a;
    layer4_outputs(5550) <= not (a or b);
    layer4_outputs(5551) <= a;
    layer4_outputs(5552) <= b;
    layer4_outputs(5553) <= a xor b;
    layer4_outputs(5554) <= not (a and b);
    layer4_outputs(5555) <= not b or a;
    layer4_outputs(5556) <= not (a or b);
    layer4_outputs(5557) <= a xor b;
    layer4_outputs(5558) <= not b or a;
    layer4_outputs(5559) <= not a or b;
    layer4_outputs(5560) <= a xor b;
    layer4_outputs(5561) <= a xor b;
    layer4_outputs(5562) <= not (a xor b);
    layer4_outputs(5563) <= a;
    layer4_outputs(5564) <= a;
    layer4_outputs(5565) <= a and b;
    layer4_outputs(5566) <= not (a xor b);
    layer4_outputs(5567) <= not b or a;
    layer4_outputs(5568) <= b;
    layer4_outputs(5569) <= not a;
    layer4_outputs(5570) <= a xor b;
    layer4_outputs(5571) <= a xor b;
    layer4_outputs(5572) <= a;
    layer4_outputs(5573) <= b;
    layer4_outputs(5574) <= b;
    layer4_outputs(5575) <= a xor b;
    layer4_outputs(5576) <= not (a xor b);
    layer4_outputs(5577) <= a and b;
    layer4_outputs(5578) <= b;
    layer4_outputs(5579) <= a;
    layer4_outputs(5580) <= not a or b;
    layer4_outputs(5581) <= not b;
    layer4_outputs(5582) <= a or b;
    layer4_outputs(5583) <= not a or b;
    layer4_outputs(5584) <= not (a xor b);
    layer4_outputs(5585) <= not b;
    layer4_outputs(5586) <= a;
    layer4_outputs(5587) <= not b;
    layer4_outputs(5588) <= a;
    layer4_outputs(5589) <= not (a xor b);
    layer4_outputs(5590) <= not a or b;
    layer4_outputs(5591) <= a xor b;
    layer4_outputs(5592) <= a;
    layer4_outputs(5593) <= a and b;
    layer4_outputs(5594) <= b;
    layer4_outputs(5595) <= a;
    layer4_outputs(5596) <= not (a and b);
    layer4_outputs(5597) <= b and not a;
    layer4_outputs(5598) <= a or b;
    layer4_outputs(5599) <= a or b;
    layer4_outputs(5600) <= b;
    layer4_outputs(5601) <= a or b;
    layer4_outputs(5602) <= not (a and b);
    layer4_outputs(5603) <= 1'b0;
    layer4_outputs(5604) <= a or b;
    layer4_outputs(5605) <= not b;
    layer4_outputs(5606) <= a and b;
    layer4_outputs(5607) <= not b or a;
    layer4_outputs(5608) <= a and b;
    layer4_outputs(5609) <= a or b;
    layer4_outputs(5610) <= a xor b;
    layer4_outputs(5611) <= not b;
    layer4_outputs(5612) <= not a;
    layer4_outputs(5613) <= not (a xor b);
    layer4_outputs(5614) <= not a or b;
    layer4_outputs(5615) <= b and not a;
    layer4_outputs(5616) <= a;
    layer4_outputs(5617) <= not (a and b);
    layer4_outputs(5618) <= not (a and b);
    layer4_outputs(5619) <= b and not a;
    layer4_outputs(5620) <= not b or a;
    layer4_outputs(5621) <= b and not a;
    layer4_outputs(5622) <= b and not a;
    layer4_outputs(5623) <= a xor b;
    layer4_outputs(5624) <= b;
    layer4_outputs(5625) <= not b;
    layer4_outputs(5626) <= a xor b;
    layer4_outputs(5627) <= not b;
    layer4_outputs(5628) <= not (a and b);
    layer4_outputs(5629) <= b;
    layer4_outputs(5630) <= b;
    layer4_outputs(5631) <= not b;
    layer4_outputs(5632) <= not b;
    layer4_outputs(5633) <= not (a xor b);
    layer4_outputs(5634) <= not (a or b);
    layer4_outputs(5635) <= b;
    layer4_outputs(5636) <= b;
    layer4_outputs(5637) <= a or b;
    layer4_outputs(5638) <= a or b;
    layer4_outputs(5639) <= not (a xor b);
    layer4_outputs(5640) <= not a;
    layer4_outputs(5641) <= not a;
    layer4_outputs(5642) <= not a or b;
    layer4_outputs(5643) <= not b;
    layer4_outputs(5644) <= a xor b;
    layer4_outputs(5645) <= a and not b;
    layer4_outputs(5646) <= not b;
    layer4_outputs(5647) <= b;
    layer4_outputs(5648) <= a and not b;
    layer4_outputs(5649) <= a xor b;
    layer4_outputs(5650) <= b;
    layer4_outputs(5651) <= not (a or b);
    layer4_outputs(5652) <= a;
    layer4_outputs(5653) <= a or b;
    layer4_outputs(5654) <= a or b;
    layer4_outputs(5655) <= a xor b;
    layer4_outputs(5656) <= a;
    layer4_outputs(5657) <= a or b;
    layer4_outputs(5658) <= a and not b;
    layer4_outputs(5659) <= a and not b;
    layer4_outputs(5660) <= not (a xor b);
    layer4_outputs(5661) <= not a;
    layer4_outputs(5662) <= a and not b;
    layer4_outputs(5663) <= b and not a;
    layer4_outputs(5664) <= a xor b;
    layer4_outputs(5665) <= not a;
    layer4_outputs(5666) <= b and not a;
    layer4_outputs(5667) <= not a or b;
    layer4_outputs(5668) <= not a or b;
    layer4_outputs(5669) <= not (a xor b);
    layer4_outputs(5670) <= not b;
    layer4_outputs(5671) <= not a;
    layer4_outputs(5672) <= not a;
    layer4_outputs(5673) <= a and not b;
    layer4_outputs(5674) <= a xor b;
    layer4_outputs(5675) <= not b;
    layer4_outputs(5676) <= b;
    layer4_outputs(5677) <= not b;
    layer4_outputs(5678) <= not b;
    layer4_outputs(5679) <= b and not a;
    layer4_outputs(5680) <= not (a xor b);
    layer4_outputs(5681) <= a;
    layer4_outputs(5682) <= not (a xor b);
    layer4_outputs(5683) <= not b;
    layer4_outputs(5684) <= b and not a;
    layer4_outputs(5685) <= not b;
    layer4_outputs(5686) <= a;
    layer4_outputs(5687) <= not b;
    layer4_outputs(5688) <= b;
    layer4_outputs(5689) <= not b;
    layer4_outputs(5690) <= a and b;
    layer4_outputs(5691) <= not (a and b);
    layer4_outputs(5692) <= b;
    layer4_outputs(5693) <= a and b;
    layer4_outputs(5694) <= not a;
    layer4_outputs(5695) <= not b;
    layer4_outputs(5696) <= a;
    layer4_outputs(5697) <= not a;
    layer4_outputs(5698) <= not a;
    layer4_outputs(5699) <= not b;
    layer4_outputs(5700) <= b;
    layer4_outputs(5701) <= b and not a;
    layer4_outputs(5702) <= a;
    layer4_outputs(5703) <= not a;
    layer4_outputs(5704) <= a xor b;
    layer4_outputs(5705) <= b and not a;
    layer4_outputs(5706) <= a;
    layer4_outputs(5707) <= b;
    layer4_outputs(5708) <= not (a xor b);
    layer4_outputs(5709) <= a;
    layer4_outputs(5710) <= not a;
    layer4_outputs(5711) <= not (a xor b);
    layer4_outputs(5712) <= not a;
    layer4_outputs(5713) <= b;
    layer4_outputs(5714) <= a or b;
    layer4_outputs(5715) <= a xor b;
    layer4_outputs(5716) <= b;
    layer4_outputs(5717) <= a xor b;
    layer4_outputs(5718) <= b;
    layer4_outputs(5719) <= b;
    layer4_outputs(5720) <= b;
    layer4_outputs(5721) <= a or b;
    layer4_outputs(5722) <= a and b;
    layer4_outputs(5723) <= not (a or b);
    layer4_outputs(5724) <= a xor b;
    layer4_outputs(5725) <= a xor b;
    layer4_outputs(5726) <= a;
    layer4_outputs(5727) <= not a;
    layer4_outputs(5728) <= not a;
    layer4_outputs(5729) <= b and not a;
    layer4_outputs(5730) <= not b or a;
    layer4_outputs(5731) <= not b or a;
    layer4_outputs(5732) <= b;
    layer4_outputs(5733) <= not b;
    layer4_outputs(5734) <= a and not b;
    layer4_outputs(5735) <= b;
    layer4_outputs(5736) <= b;
    layer4_outputs(5737) <= not (a or b);
    layer4_outputs(5738) <= b and not a;
    layer4_outputs(5739) <= b and not a;
    layer4_outputs(5740) <= a xor b;
    layer4_outputs(5741) <= a or b;
    layer4_outputs(5742) <= b;
    layer4_outputs(5743) <= not b;
    layer4_outputs(5744) <= b;
    layer4_outputs(5745) <= b and not a;
    layer4_outputs(5746) <= not (a xor b);
    layer4_outputs(5747) <= not (a xor b);
    layer4_outputs(5748) <= not (a xor b);
    layer4_outputs(5749) <= not b or a;
    layer4_outputs(5750) <= a xor b;
    layer4_outputs(5751) <= a;
    layer4_outputs(5752) <= not a;
    layer4_outputs(5753) <= a;
    layer4_outputs(5754) <= a and not b;
    layer4_outputs(5755) <= a xor b;
    layer4_outputs(5756) <= a or b;
    layer4_outputs(5757) <= a;
    layer4_outputs(5758) <= not a;
    layer4_outputs(5759) <= b;
    layer4_outputs(5760) <= not b;
    layer4_outputs(5761) <= a and not b;
    layer4_outputs(5762) <= a or b;
    layer4_outputs(5763) <= b;
    layer4_outputs(5764) <= not a or b;
    layer4_outputs(5765) <= not b;
    layer4_outputs(5766) <= not b;
    layer4_outputs(5767) <= not a;
    layer4_outputs(5768) <= a xor b;
    layer4_outputs(5769) <= not (a or b);
    layer4_outputs(5770) <= not b;
    layer4_outputs(5771) <= a and b;
    layer4_outputs(5772) <= a;
    layer4_outputs(5773) <= not b;
    layer4_outputs(5774) <= not a;
    layer4_outputs(5775) <= not (a xor b);
    layer4_outputs(5776) <= a and not b;
    layer4_outputs(5777) <= not b;
    layer4_outputs(5778) <= a and b;
    layer4_outputs(5779) <= b;
    layer4_outputs(5780) <= not (a and b);
    layer4_outputs(5781) <= b;
    layer4_outputs(5782) <= not b;
    layer4_outputs(5783) <= not a;
    layer4_outputs(5784) <= a and b;
    layer4_outputs(5785) <= a;
    layer4_outputs(5786) <= b and not a;
    layer4_outputs(5787) <= a;
    layer4_outputs(5788) <= a and not b;
    layer4_outputs(5789) <= a xor b;
    layer4_outputs(5790) <= not b or a;
    layer4_outputs(5791) <= not a or b;
    layer4_outputs(5792) <= a;
    layer4_outputs(5793) <= not a or b;
    layer4_outputs(5794) <= a;
    layer4_outputs(5795) <= a or b;
    layer4_outputs(5796) <= a xor b;
    layer4_outputs(5797) <= b;
    layer4_outputs(5798) <= a xor b;
    layer4_outputs(5799) <= not a;
    layer4_outputs(5800) <= a;
    layer4_outputs(5801) <= a;
    layer4_outputs(5802) <= a xor b;
    layer4_outputs(5803) <= a;
    layer4_outputs(5804) <= b;
    layer4_outputs(5805) <= b;
    layer4_outputs(5806) <= a and not b;
    layer4_outputs(5807) <= not (a xor b);
    layer4_outputs(5808) <= not a;
    layer4_outputs(5809) <= b and not a;
    layer4_outputs(5810) <= a and not b;
    layer4_outputs(5811) <= not (a xor b);
    layer4_outputs(5812) <= not (a and b);
    layer4_outputs(5813) <= not (a and b);
    layer4_outputs(5814) <= not a;
    layer4_outputs(5815) <= a xor b;
    layer4_outputs(5816) <= b;
    layer4_outputs(5817) <= not a or b;
    layer4_outputs(5818) <= not a;
    layer4_outputs(5819) <= not (a and b);
    layer4_outputs(5820) <= not a;
    layer4_outputs(5821) <= a and not b;
    layer4_outputs(5822) <= b and not a;
    layer4_outputs(5823) <= a;
    layer4_outputs(5824) <= b;
    layer4_outputs(5825) <= not (a xor b);
    layer4_outputs(5826) <= not (a xor b);
    layer4_outputs(5827) <= not (a xor b);
    layer4_outputs(5828) <= a;
    layer4_outputs(5829) <= b;
    layer4_outputs(5830) <= a and not b;
    layer4_outputs(5831) <= b and not a;
    layer4_outputs(5832) <= a;
    layer4_outputs(5833) <= b;
    layer4_outputs(5834) <= not (a or b);
    layer4_outputs(5835) <= not (a or b);
    layer4_outputs(5836) <= not b;
    layer4_outputs(5837) <= a and b;
    layer4_outputs(5838) <= not (a and b);
    layer4_outputs(5839) <= not a or b;
    layer4_outputs(5840) <= not b;
    layer4_outputs(5841) <= not b;
    layer4_outputs(5842) <= not b or a;
    layer4_outputs(5843) <= b;
    layer4_outputs(5844) <= a;
    layer4_outputs(5845) <= a and b;
    layer4_outputs(5846) <= a;
    layer4_outputs(5847) <= not a;
    layer4_outputs(5848) <= a and not b;
    layer4_outputs(5849) <= a xor b;
    layer4_outputs(5850) <= b;
    layer4_outputs(5851) <= a and not b;
    layer4_outputs(5852) <= a xor b;
    layer4_outputs(5853) <= a xor b;
    layer4_outputs(5854) <= b;
    layer4_outputs(5855) <= not b;
    layer4_outputs(5856) <= not a or b;
    layer4_outputs(5857) <= not b;
    layer4_outputs(5858) <= a xor b;
    layer4_outputs(5859) <= a;
    layer4_outputs(5860) <= not b;
    layer4_outputs(5861) <= not a;
    layer4_outputs(5862) <= b;
    layer4_outputs(5863) <= a and not b;
    layer4_outputs(5864) <= not a;
    layer4_outputs(5865) <= not a or b;
    layer4_outputs(5866) <= a xor b;
    layer4_outputs(5867) <= not a;
    layer4_outputs(5868) <= not (a or b);
    layer4_outputs(5869) <= b;
    layer4_outputs(5870) <= a;
    layer4_outputs(5871) <= a;
    layer4_outputs(5872) <= not (a xor b);
    layer4_outputs(5873) <= not a or b;
    layer4_outputs(5874) <= not b;
    layer4_outputs(5875) <= b;
    layer4_outputs(5876) <= a xor b;
    layer4_outputs(5877) <= b;
    layer4_outputs(5878) <= not a or b;
    layer4_outputs(5879) <= not a or b;
    layer4_outputs(5880) <= not a;
    layer4_outputs(5881) <= a xor b;
    layer4_outputs(5882) <= a;
    layer4_outputs(5883) <= not a or b;
    layer4_outputs(5884) <= not a;
    layer4_outputs(5885) <= a xor b;
    layer4_outputs(5886) <= b;
    layer4_outputs(5887) <= b;
    layer4_outputs(5888) <= not a;
    layer4_outputs(5889) <= not b or a;
    layer4_outputs(5890) <= a xor b;
    layer4_outputs(5891) <= b and not a;
    layer4_outputs(5892) <= b;
    layer4_outputs(5893) <= a xor b;
    layer4_outputs(5894) <= not b or a;
    layer4_outputs(5895) <= not a or b;
    layer4_outputs(5896) <= not a or b;
    layer4_outputs(5897) <= not (a xor b);
    layer4_outputs(5898) <= not b;
    layer4_outputs(5899) <= a xor b;
    layer4_outputs(5900) <= a;
    layer4_outputs(5901) <= not b;
    layer4_outputs(5902) <= b;
    layer4_outputs(5903) <= not (a and b);
    layer4_outputs(5904) <= not a;
    layer4_outputs(5905) <= a xor b;
    layer4_outputs(5906) <= not a;
    layer4_outputs(5907) <= not b;
    layer4_outputs(5908) <= not b or a;
    layer4_outputs(5909) <= b;
    layer4_outputs(5910) <= b;
    layer4_outputs(5911) <= not b or a;
    layer4_outputs(5912) <= a xor b;
    layer4_outputs(5913) <= not (a and b);
    layer4_outputs(5914) <= b;
    layer4_outputs(5915) <= b;
    layer4_outputs(5916) <= not b;
    layer4_outputs(5917) <= a and not b;
    layer4_outputs(5918) <= a;
    layer4_outputs(5919) <= not a;
    layer4_outputs(5920) <= not b;
    layer4_outputs(5921) <= b;
    layer4_outputs(5922) <= b;
    layer4_outputs(5923) <= a;
    layer4_outputs(5924) <= not b or a;
    layer4_outputs(5925) <= a;
    layer4_outputs(5926) <= not a;
    layer4_outputs(5927) <= not a or b;
    layer4_outputs(5928) <= not (a xor b);
    layer4_outputs(5929) <= not (a and b);
    layer4_outputs(5930) <= a and b;
    layer4_outputs(5931) <= b and not a;
    layer4_outputs(5932) <= not (a xor b);
    layer4_outputs(5933) <= not (a and b);
    layer4_outputs(5934) <= not (a xor b);
    layer4_outputs(5935) <= not (a or b);
    layer4_outputs(5936) <= a and not b;
    layer4_outputs(5937) <= a and b;
    layer4_outputs(5938) <= b;
    layer4_outputs(5939) <= a and b;
    layer4_outputs(5940) <= not b;
    layer4_outputs(5941) <= b;
    layer4_outputs(5942) <= a;
    layer4_outputs(5943) <= not (a and b);
    layer4_outputs(5944) <= not b;
    layer4_outputs(5945) <= a;
    layer4_outputs(5946) <= not (a xor b);
    layer4_outputs(5947) <= not a;
    layer4_outputs(5948) <= a;
    layer4_outputs(5949) <= not a;
    layer4_outputs(5950) <= not a or b;
    layer4_outputs(5951) <= not (a xor b);
    layer4_outputs(5952) <= not a;
    layer4_outputs(5953) <= b;
    layer4_outputs(5954) <= not a or b;
    layer4_outputs(5955) <= not (a and b);
    layer4_outputs(5956) <= a and not b;
    layer4_outputs(5957) <= a and not b;
    layer4_outputs(5958) <= a xor b;
    layer4_outputs(5959) <= a xor b;
    layer4_outputs(5960) <= not (a xor b);
    layer4_outputs(5961) <= not (a or b);
    layer4_outputs(5962) <= not a;
    layer4_outputs(5963) <= a and not b;
    layer4_outputs(5964) <= not (a xor b);
    layer4_outputs(5965) <= not (a xor b);
    layer4_outputs(5966) <= not a;
    layer4_outputs(5967) <= not a or b;
    layer4_outputs(5968) <= not b;
    layer4_outputs(5969) <= not a;
    layer4_outputs(5970) <= not b or a;
    layer4_outputs(5971) <= not b or a;
    layer4_outputs(5972) <= b and not a;
    layer4_outputs(5973) <= a xor b;
    layer4_outputs(5974) <= not b;
    layer4_outputs(5975) <= b;
    layer4_outputs(5976) <= not b;
    layer4_outputs(5977) <= not b;
    layer4_outputs(5978) <= not a or b;
    layer4_outputs(5979) <= not b;
    layer4_outputs(5980) <= not b or a;
    layer4_outputs(5981) <= b and not a;
    layer4_outputs(5982) <= a;
    layer4_outputs(5983) <= not b;
    layer4_outputs(5984) <= b;
    layer4_outputs(5985) <= not (a and b);
    layer4_outputs(5986) <= b;
    layer4_outputs(5987) <= b;
    layer4_outputs(5988) <= not (a and b);
    layer4_outputs(5989) <= not (a xor b);
    layer4_outputs(5990) <= a;
    layer4_outputs(5991) <= not a;
    layer4_outputs(5992) <= b;
    layer4_outputs(5993) <= a;
    layer4_outputs(5994) <= not (a and b);
    layer4_outputs(5995) <= not b;
    layer4_outputs(5996) <= a xor b;
    layer4_outputs(5997) <= not b;
    layer4_outputs(5998) <= not (a and b);
    layer4_outputs(5999) <= not a;
    layer4_outputs(6000) <= a and not b;
    layer4_outputs(6001) <= not (a and b);
    layer4_outputs(6002) <= not (a xor b);
    layer4_outputs(6003) <= not (a or b);
    layer4_outputs(6004) <= b;
    layer4_outputs(6005) <= not b;
    layer4_outputs(6006) <= not b or a;
    layer4_outputs(6007) <= a xor b;
    layer4_outputs(6008) <= b;
    layer4_outputs(6009) <= not a;
    layer4_outputs(6010) <= a or b;
    layer4_outputs(6011) <= not (a xor b);
    layer4_outputs(6012) <= a xor b;
    layer4_outputs(6013) <= not a;
    layer4_outputs(6014) <= not a;
    layer4_outputs(6015) <= a;
    layer4_outputs(6016) <= not (a or b);
    layer4_outputs(6017) <= not (a xor b);
    layer4_outputs(6018) <= a;
    layer4_outputs(6019) <= not b;
    layer4_outputs(6020) <= not b;
    layer4_outputs(6021) <= b and not a;
    layer4_outputs(6022) <= a xor b;
    layer4_outputs(6023) <= a;
    layer4_outputs(6024) <= a or b;
    layer4_outputs(6025) <= not a;
    layer4_outputs(6026) <= a and not b;
    layer4_outputs(6027) <= b and not a;
    layer4_outputs(6028) <= b;
    layer4_outputs(6029) <= not b or a;
    layer4_outputs(6030) <= not a;
    layer4_outputs(6031) <= not b;
    layer4_outputs(6032) <= a or b;
    layer4_outputs(6033) <= a;
    layer4_outputs(6034) <= not (a xor b);
    layer4_outputs(6035) <= not (a and b);
    layer4_outputs(6036) <= not a;
    layer4_outputs(6037) <= a;
    layer4_outputs(6038) <= not (a or b);
    layer4_outputs(6039) <= a or b;
    layer4_outputs(6040) <= a and b;
    layer4_outputs(6041) <= b;
    layer4_outputs(6042) <= b;
    layer4_outputs(6043) <= a;
    layer4_outputs(6044) <= b;
    layer4_outputs(6045) <= a xor b;
    layer4_outputs(6046) <= a;
    layer4_outputs(6047) <= a;
    layer4_outputs(6048) <= a;
    layer4_outputs(6049) <= not b or a;
    layer4_outputs(6050) <= not a or b;
    layer4_outputs(6051) <= not a;
    layer4_outputs(6052) <= not b;
    layer4_outputs(6053) <= b;
    layer4_outputs(6054) <= not (a or b);
    layer4_outputs(6055) <= not a;
    layer4_outputs(6056) <= a and b;
    layer4_outputs(6057) <= b and not a;
    layer4_outputs(6058) <= not (a and b);
    layer4_outputs(6059) <= not (a xor b);
    layer4_outputs(6060) <= not (a or b);
    layer4_outputs(6061) <= not a;
    layer4_outputs(6062) <= b and not a;
    layer4_outputs(6063) <= not a or b;
    layer4_outputs(6064) <= not a;
    layer4_outputs(6065) <= a;
    layer4_outputs(6066) <= not a;
    layer4_outputs(6067) <= b and not a;
    layer4_outputs(6068) <= not (a xor b);
    layer4_outputs(6069) <= a;
    layer4_outputs(6070) <= a and not b;
    layer4_outputs(6071) <= not b or a;
    layer4_outputs(6072) <= not (a xor b);
    layer4_outputs(6073) <= not a;
    layer4_outputs(6074) <= not (a xor b);
    layer4_outputs(6075) <= not a or b;
    layer4_outputs(6076) <= b and not a;
    layer4_outputs(6077) <= a;
    layer4_outputs(6078) <= a and b;
    layer4_outputs(6079) <= a;
    layer4_outputs(6080) <= a or b;
    layer4_outputs(6081) <= b;
    layer4_outputs(6082) <= a;
    layer4_outputs(6083) <= a;
    layer4_outputs(6084) <= b;
    layer4_outputs(6085) <= a xor b;
    layer4_outputs(6086) <= not a;
    layer4_outputs(6087) <= not (a or b);
    layer4_outputs(6088) <= not b;
    layer4_outputs(6089) <= not (a xor b);
    layer4_outputs(6090) <= not a;
    layer4_outputs(6091) <= b and not a;
    layer4_outputs(6092) <= b;
    layer4_outputs(6093) <= not (a or b);
    layer4_outputs(6094) <= not b;
    layer4_outputs(6095) <= b;
    layer4_outputs(6096) <= a and not b;
    layer4_outputs(6097) <= a;
    layer4_outputs(6098) <= b;
    layer4_outputs(6099) <= a xor b;
    layer4_outputs(6100) <= a and not b;
    layer4_outputs(6101) <= a and b;
    layer4_outputs(6102) <= a and not b;
    layer4_outputs(6103) <= not a;
    layer4_outputs(6104) <= b and not a;
    layer4_outputs(6105) <= not (a xor b);
    layer4_outputs(6106) <= not a;
    layer4_outputs(6107) <= not b;
    layer4_outputs(6108) <= not b or a;
    layer4_outputs(6109) <= not (a xor b);
    layer4_outputs(6110) <= a;
    layer4_outputs(6111) <= b;
    layer4_outputs(6112) <= b;
    layer4_outputs(6113) <= a;
    layer4_outputs(6114) <= not (a xor b);
    layer4_outputs(6115) <= b;
    layer4_outputs(6116) <= not a or b;
    layer4_outputs(6117) <= not a;
    layer4_outputs(6118) <= not (a or b);
    layer4_outputs(6119) <= not b;
    layer4_outputs(6120) <= not (a xor b);
    layer4_outputs(6121) <= b;
    layer4_outputs(6122) <= not b;
    layer4_outputs(6123) <= not b;
    layer4_outputs(6124) <= not a or b;
    layer4_outputs(6125) <= a and b;
    layer4_outputs(6126) <= b;
    layer4_outputs(6127) <= a;
    layer4_outputs(6128) <= b and not a;
    layer4_outputs(6129) <= not (a and b);
    layer4_outputs(6130) <= not a;
    layer4_outputs(6131) <= not b;
    layer4_outputs(6132) <= a and not b;
    layer4_outputs(6133) <= not (a and b);
    layer4_outputs(6134) <= not a;
    layer4_outputs(6135) <= not (a and b);
    layer4_outputs(6136) <= a;
    layer4_outputs(6137) <= not (a xor b);
    layer4_outputs(6138) <= not b;
    layer4_outputs(6139) <= a;
    layer4_outputs(6140) <= a and not b;
    layer4_outputs(6141) <= 1'b0;
    layer4_outputs(6142) <= b;
    layer4_outputs(6143) <= a and not b;
    layer4_outputs(6144) <= a and b;
    layer4_outputs(6145) <= a;
    layer4_outputs(6146) <= not b;
    layer4_outputs(6147) <= a xor b;
    layer4_outputs(6148) <= b and not a;
    layer4_outputs(6149) <= a;
    layer4_outputs(6150) <= a and b;
    layer4_outputs(6151) <= not (a and b);
    layer4_outputs(6152) <= a xor b;
    layer4_outputs(6153) <= not (a xor b);
    layer4_outputs(6154) <= not a;
    layer4_outputs(6155) <= not (a or b);
    layer4_outputs(6156) <= b;
    layer4_outputs(6157) <= a and b;
    layer4_outputs(6158) <= not (a xor b);
    layer4_outputs(6159) <= not (a xor b);
    layer4_outputs(6160) <= b;
    layer4_outputs(6161) <= a and not b;
    layer4_outputs(6162) <= a;
    layer4_outputs(6163) <= not b;
    layer4_outputs(6164) <= b;
    layer4_outputs(6165) <= b and not a;
    layer4_outputs(6166) <= not b;
    layer4_outputs(6167) <= a xor b;
    layer4_outputs(6168) <= a and not b;
    layer4_outputs(6169) <= a;
    layer4_outputs(6170) <= not (a and b);
    layer4_outputs(6171) <= not b;
    layer4_outputs(6172) <= 1'b0;
    layer4_outputs(6173) <= not a;
    layer4_outputs(6174) <= a or b;
    layer4_outputs(6175) <= a xor b;
    layer4_outputs(6176) <= a xor b;
    layer4_outputs(6177) <= not (a or b);
    layer4_outputs(6178) <= 1'b1;
    layer4_outputs(6179) <= b and not a;
    layer4_outputs(6180) <= a or b;
    layer4_outputs(6181) <= not b;
    layer4_outputs(6182) <= b;
    layer4_outputs(6183) <= a and not b;
    layer4_outputs(6184) <= not a;
    layer4_outputs(6185) <= a;
    layer4_outputs(6186) <= not b;
    layer4_outputs(6187) <= not b;
    layer4_outputs(6188) <= not (a xor b);
    layer4_outputs(6189) <= a and not b;
    layer4_outputs(6190) <= not a;
    layer4_outputs(6191) <= a xor b;
    layer4_outputs(6192) <= a;
    layer4_outputs(6193) <= not a;
    layer4_outputs(6194) <= not a;
    layer4_outputs(6195) <= not a or b;
    layer4_outputs(6196) <= a and not b;
    layer4_outputs(6197) <= b and not a;
    layer4_outputs(6198) <= b;
    layer4_outputs(6199) <= b and not a;
    layer4_outputs(6200) <= not a;
    layer4_outputs(6201) <= not (a xor b);
    layer4_outputs(6202) <= a and not b;
    layer4_outputs(6203) <= not (a xor b);
    layer4_outputs(6204) <= b;
    layer4_outputs(6205) <= not a or b;
    layer4_outputs(6206) <= not (a and b);
    layer4_outputs(6207) <= b;
    layer4_outputs(6208) <= not (a xor b);
    layer4_outputs(6209) <= not (a or b);
    layer4_outputs(6210) <= not b or a;
    layer4_outputs(6211) <= not b;
    layer4_outputs(6212) <= not b;
    layer4_outputs(6213) <= a;
    layer4_outputs(6214) <= not (a xor b);
    layer4_outputs(6215) <= not a or b;
    layer4_outputs(6216) <= b;
    layer4_outputs(6217) <= not a or b;
    layer4_outputs(6218) <= not (a or b);
    layer4_outputs(6219) <= a xor b;
    layer4_outputs(6220) <= a;
    layer4_outputs(6221) <= not b or a;
    layer4_outputs(6222) <= a xor b;
    layer4_outputs(6223) <= b;
    layer4_outputs(6224) <= not b;
    layer4_outputs(6225) <= not (a or b);
    layer4_outputs(6226) <= b;
    layer4_outputs(6227) <= a or b;
    layer4_outputs(6228) <= not (a xor b);
    layer4_outputs(6229) <= a;
    layer4_outputs(6230) <= not (a and b);
    layer4_outputs(6231) <= not b;
    layer4_outputs(6232) <= a or b;
    layer4_outputs(6233) <= not (a and b);
    layer4_outputs(6234) <= not (a or b);
    layer4_outputs(6235) <= not (a and b);
    layer4_outputs(6236) <= b;
    layer4_outputs(6237) <= b;
    layer4_outputs(6238) <= a and b;
    layer4_outputs(6239) <= a xor b;
    layer4_outputs(6240) <= a and not b;
    layer4_outputs(6241) <= not a;
    layer4_outputs(6242) <= not a;
    layer4_outputs(6243) <= b;
    layer4_outputs(6244) <= not b;
    layer4_outputs(6245) <= not a;
    layer4_outputs(6246) <= not a;
    layer4_outputs(6247) <= a xor b;
    layer4_outputs(6248) <= not (a xor b);
    layer4_outputs(6249) <= a or b;
    layer4_outputs(6250) <= b;
    layer4_outputs(6251) <= not a or b;
    layer4_outputs(6252) <= not (a xor b);
    layer4_outputs(6253) <= not (a xor b);
    layer4_outputs(6254) <= a;
    layer4_outputs(6255) <= a and b;
    layer4_outputs(6256) <= not (a or b);
    layer4_outputs(6257) <= not (a and b);
    layer4_outputs(6258) <= a and not b;
    layer4_outputs(6259) <= a;
    layer4_outputs(6260) <= not (a xor b);
    layer4_outputs(6261) <= not (a xor b);
    layer4_outputs(6262) <= not b;
    layer4_outputs(6263) <= not a;
    layer4_outputs(6264) <= a;
    layer4_outputs(6265) <= not (a xor b);
    layer4_outputs(6266) <= not b or a;
    layer4_outputs(6267) <= a;
    layer4_outputs(6268) <= not (a or b);
    layer4_outputs(6269) <= b and not a;
    layer4_outputs(6270) <= not b;
    layer4_outputs(6271) <= b;
    layer4_outputs(6272) <= a or b;
    layer4_outputs(6273) <= not a;
    layer4_outputs(6274) <= not a or b;
    layer4_outputs(6275) <= not a;
    layer4_outputs(6276) <= not (a or b);
    layer4_outputs(6277) <= a xor b;
    layer4_outputs(6278) <= a xor b;
    layer4_outputs(6279) <= not (a or b);
    layer4_outputs(6280) <= a or b;
    layer4_outputs(6281) <= a;
    layer4_outputs(6282) <= not (a and b);
    layer4_outputs(6283) <= not a;
    layer4_outputs(6284) <= a and b;
    layer4_outputs(6285) <= a or b;
    layer4_outputs(6286) <= not a;
    layer4_outputs(6287) <= not (a or b);
    layer4_outputs(6288) <= not a;
    layer4_outputs(6289) <= not b;
    layer4_outputs(6290) <= a xor b;
    layer4_outputs(6291) <= not a;
    layer4_outputs(6292) <= b;
    layer4_outputs(6293) <= b;
    layer4_outputs(6294) <= b and not a;
    layer4_outputs(6295) <= not (a xor b);
    layer4_outputs(6296) <= not (a or b);
    layer4_outputs(6297) <= not b;
    layer4_outputs(6298) <= 1'b0;
    layer4_outputs(6299) <= a xor b;
    layer4_outputs(6300) <= b;
    layer4_outputs(6301) <= a xor b;
    layer4_outputs(6302) <= not a;
    layer4_outputs(6303) <= not b or a;
    layer4_outputs(6304) <= not b;
    layer4_outputs(6305) <= not a or b;
    layer4_outputs(6306) <= not a;
    layer4_outputs(6307) <= a xor b;
    layer4_outputs(6308) <= not b;
    layer4_outputs(6309) <= b;
    layer4_outputs(6310) <= b;
    layer4_outputs(6311) <= not b;
    layer4_outputs(6312) <= a or b;
    layer4_outputs(6313) <= a xor b;
    layer4_outputs(6314) <= b;
    layer4_outputs(6315) <= a;
    layer4_outputs(6316) <= not a;
    layer4_outputs(6317) <= a;
    layer4_outputs(6318) <= a and not b;
    layer4_outputs(6319) <= not b or a;
    layer4_outputs(6320) <= a or b;
    layer4_outputs(6321) <= not (a or b);
    layer4_outputs(6322) <= b;
    layer4_outputs(6323) <= a and b;
    layer4_outputs(6324) <= a and b;
    layer4_outputs(6325) <= not a;
    layer4_outputs(6326) <= not b;
    layer4_outputs(6327) <= not b;
    layer4_outputs(6328) <= a and b;
    layer4_outputs(6329) <= not b;
    layer4_outputs(6330) <= not a;
    layer4_outputs(6331) <= not (a xor b);
    layer4_outputs(6332) <= not (a xor b);
    layer4_outputs(6333) <= not (a or b);
    layer4_outputs(6334) <= not b;
    layer4_outputs(6335) <= b;
    layer4_outputs(6336) <= a;
    layer4_outputs(6337) <= a or b;
    layer4_outputs(6338) <= not a;
    layer4_outputs(6339) <= not b;
    layer4_outputs(6340) <= not b;
    layer4_outputs(6341) <= not (a xor b);
    layer4_outputs(6342) <= not b;
    layer4_outputs(6343) <= not (a xor b);
    layer4_outputs(6344) <= not (a or b);
    layer4_outputs(6345) <= not b;
    layer4_outputs(6346) <= a and b;
    layer4_outputs(6347) <= not a;
    layer4_outputs(6348) <= b;
    layer4_outputs(6349) <= not (a and b);
    layer4_outputs(6350) <= a and b;
    layer4_outputs(6351) <= not a;
    layer4_outputs(6352) <= not b or a;
    layer4_outputs(6353) <= a xor b;
    layer4_outputs(6354) <= a;
    layer4_outputs(6355) <= b;
    layer4_outputs(6356) <= not a;
    layer4_outputs(6357) <= a xor b;
    layer4_outputs(6358) <= a and not b;
    layer4_outputs(6359) <= a and b;
    layer4_outputs(6360) <= a and b;
    layer4_outputs(6361) <= a xor b;
    layer4_outputs(6362) <= a and not b;
    layer4_outputs(6363) <= not b;
    layer4_outputs(6364) <= not (a or b);
    layer4_outputs(6365) <= not a or b;
    layer4_outputs(6366) <= b;
    layer4_outputs(6367) <= a or b;
    layer4_outputs(6368) <= a or b;
    layer4_outputs(6369) <= a and b;
    layer4_outputs(6370) <= a or b;
    layer4_outputs(6371) <= not (a xor b);
    layer4_outputs(6372) <= not (a and b);
    layer4_outputs(6373) <= b and not a;
    layer4_outputs(6374) <= a;
    layer4_outputs(6375) <= not b;
    layer4_outputs(6376) <= b;
    layer4_outputs(6377) <= not (a or b);
    layer4_outputs(6378) <= not b;
    layer4_outputs(6379) <= a;
    layer4_outputs(6380) <= a or b;
    layer4_outputs(6381) <= b and not a;
    layer4_outputs(6382) <= not (a or b);
    layer4_outputs(6383) <= not (a and b);
    layer4_outputs(6384) <= not a;
    layer4_outputs(6385) <= a or b;
    layer4_outputs(6386) <= a xor b;
    layer4_outputs(6387) <= a xor b;
    layer4_outputs(6388) <= not b or a;
    layer4_outputs(6389) <= not (a or b);
    layer4_outputs(6390) <= b;
    layer4_outputs(6391) <= a xor b;
    layer4_outputs(6392) <= not b or a;
    layer4_outputs(6393) <= a and b;
    layer4_outputs(6394) <= not a;
    layer4_outputs(6395) <= a xor b;
    layer4_outputs(6396) <= b;
    layer4_outputs(6397) <= not (a xor b);
    layer4_outputs(6398) <= not a or b;
    layer4_outputs(6399) <= a and not b;
    layer4_outputs(6400) <= not (a or b);
    layer4_outputs(6401) <= a and not b;
    layer4_outputs(6402) <= not (a xor b);
    layer4_outputs(6403) <= a and not b;
    layer4_outputs(6404) <= not a;
    layer4_outputs(6405) <= not a;
    layer4_outputs(6406) <= not b or a;
    layer4_outputs(6407) <= a and not b;
    layer4_outputs(6408) <= not a or b;
    layer4_outputs(6409) <= not b;
    layer4_outputs(6410) <= not a;
    layer4_outputs(6411) <= not a;
    layer4_outputs(6412) <= not (a or b);
    layer4_outputs(6413) <= not a;
    layer4_outputs(6414) <= a xor b;
    layer4_outputs(6415) <= not a;
    layer4_outputs(6416) <= a xor b;
    layer4_outputs(6417) <= b;
    layer4_outputs(6418) <= not b or a;
    layer4_outputs(6419) <= not a;
    layer4_outputs(6420) <= not a or b;
    layer4_outputs(6421) <= not a;
    layer4_outputs(6422) <= not (a or b);
    layer4_outputs(6423) <= a or b;
    layer4_outputs(6424) <= not a or b;
    layer4_outputs(6425) <= not (a xor b);
    layer4_outputs(6426) <= not (a or b);
    layer4_outputs(6427) <= a xor b;
    layer4_outputs(6428) <= a xor b;
    layer4_outputs(6429) <= b;
    layer4_outputs(6430) <= b;
    layer4_outputs(6431) <= not (a xor b);
    layer4_outputs(6432) <= b;
    layer4_outputs(6433) <= a xor b;
    layer4_outputs(6434) <= not (a or b);
    layer4_outputs(6435) <= a or b;
    layer4_outputs(6436) <= b and not a;
    layer4_outputs(6437) <= not (a or b);
    layer4_outputs(6438) <= a or b;
    layer4_outputs(6439) <= not b;
    layer4_outputs(6440) <= a and not b;
    layer4_outputs(6441) <= a xor b;
    layer4_outputs(6442) <= not (a xor b);
    layer4_outputs(6443) <= a xor b;
    layer4_outputs(6444) <= b;
    layer4_outputs(6445) <= a;
    layer4_outputs(6446) <= not a or b;
    layer4_outputs(6447) <= not (a and b);
    layer4_outputs(6448) <= not a;
    layer4_outputs(6449) <= b;
    layer4_outputs(6450) <= a;
    layer4_outputs(6451) <= not (a xor b);
    layer4_outputs(6452) <= a xor b;
    layer4_outputs(6453) <= a;
    layer4_outputs(6454) <= a and b;
    layer4_outputs(6455) <= not b;
    layer4_outputs(6456) <= a;
    layer4_outputs(6457) <= not b;
    layer4_outputs(6458) <= a;
    layer4_outputs(6459) <= not b;
    layer4_outputs(6460) <= not b;
    layer4_outputs(6461) <= not a or b;
    layer4_outputs(6462) <= a;
    layer4_outputs(6463) <= not a;
    layer4_outputs(6464) <= b;
    layer4_outputs(6465) <= not b;
    layer4_outputs(6466) <= not a;
    layer4_outputs(6467) <= not a or b;
    layer4_outputs(6468) <= a and b;
    layer4_outputs(6469) <= a or b;
    layer4_outputs(6470) <= a;
    layer4_outputs(6471) <= a and not b;
    layer4_outputs(6472) <= a;
    layer4_outputs(6473) <= a;
    layer4_outputs(6474) <= b;
    layer4_outputs(6475) <= not b;
    layer4_outputs(6476) <= not a or b;
    layer4_outputs(6477) <= a;
    layer4_outputs(6478) <= b;
    layer4_outputs(6479) <= not b;
    layer4_outputs(6480) <= not b;
    layer4_outputs(6481) <= not (a xor b);
    layer4_outputs(6482) <= not a;
    layer4_outputs(6483) <= a;
    layer4_outputs(6484) <= not a;
    layer4_outputs(6485) <= not a;
    layer4_outputs(6486) <= not (a xor b);
    layer4_outputs(6487) <= not (a xor b);
    layer4_outputs(6488) <= a or b;
    layer4_outputs(6489) <= a or b;
    layer4_outputs(6490) <= not a;
    layer4_outputs(6491) <= not (a xor b);
    layer4_outputs(6492) <= not a or b;
    layer4_outputs(6493) <= a or b;
    layer4_outputs(6494) <= not a or b;
    layer4_outputs(6495) <= not a or b;
    layer4_outputs(6496) <= b and not a;
    layer4_outputs(6497) <= not (a or b);
    layer4_outputs(6498) <= a;
    layer4_outputs(6499) <= not b;
    layer4_outputs(6500) <= b;
    layer4_outputs(6501) <= b;
    layer4_outputs(6502) <= not (a xor b);
    layer4_outputs(6503) <= a xor b;
    layer4_outputs(6504) <= a and not b;
    layer4_outputs(6505) <= not b;
    layer4_outputs(6506) <= not b or a;
    layer4_outputs(6507) <= a or b;
    layer4_outputs(6508) <= a or b;
    layer4_outputs(6509) <= b;
    layer4_outputs(6510) <= a or b;
    layer4_outputs(6511) <= a;
    layer4_outputs(6512) <= a xor b;
    layer4_outputs(6513) <= a or b;
    layer4_outputs(6514) <= not (a xor b);
    layer4_outputs(6515) <= not b;
    layer4_outputs(6516) <= not b or a;
    layer4_outputs(6517) <= not b;
    layer4_outputs(6518) <= not a;
    layer4_outputs(6519) <= a or b;
    layer4_outputs(6520) <= not (a xor b);
    layer4_outputs(6521) <= a xor b;
    layer4_outputs(6522) <= not a or b;
    layer4_outputs(6523) <= not b;
    layer4_outputs(6524) <= b;
    layer4_outputs(6525) <= not a;
    layer4_outputs(6526) <= not b;
    layer4_outputs(6527) <= a;
    layer4_outputs(6528) <= a;
    layer4_outputs(6529) <= not (a or b);
    layer4_outputs(6530) <= b;
    layer4_outputs(6531) <= a and not b;
    layer4_outputs(6532) <= a and b;
    layer4_outputs(6533) <= not a;
    layer4_outputs(6534) <= a;
    layer4_outputs(6535) <= b;
    layer4_outputs(6536) <= not (a xor b);
    layer4_outputs(6537) <= not (a or b);
    layer4_outputs(6538) <= a and b;
    layer4_outputs(6539) <= a xor b;
    layer4_outputs(6540) <= b;
    layer4_outputs(6541) <= a and b;
    layer4_outputs(6542) <= a or b;
    layer4_outputs(6543) <= not (a or b);
    layer4_outputs(6544) <= a and not b;
    layer4_outputs(6545) <= b;
    layer4_outputs(6546) <= a and b;
    layer4_outputs(6547) <= not (a or b);
    layer4_outputs(6548) <= not a or b;
    layer4_outputs(6549) <= b;
    layer4_outputs(6550) <= not (a and b);
    layer4_outputs(6551) <= not (a xor b);
    layer4_outputs(6552) <= b;
    layer4_outputs(6553) <= not (a xor b);
    layer4_outputs(6554) <= a;
    layer4_outputs(6555) <= not b;
    layer4_outputs(6556) <= a or b;
    layer4_outputs(6557) <= a;
    layer4_outputs(6558) <= not a;
    layer4_outputs(6559) <= not (a and b);
    layer4_outputs(6560) <= not (a or b);
    layer4_outputs(6561) <= a and b;
    layer4_outputs(6562) <= b;
    layer4_outputs(6563) <= not a;
    layer4_outputs(6564) <= b;
    layer4_outputs(6565) <= b;
    layer4_outputs(6566) <= not b;
    layer4_outputs(6567) <= a or b;
    layer4_outputs(6568) <= not b;
    layer4_outputs(6569) <= not a;
    layer4_outputs(6570) <= a and b;
    layer4_outputs(6571) <= a and b;
    layer4_outputs(6572) <= a and b;
    layer4_outputs(6573) <= not (a xor b);
    layer4_outputs(6574) <= a and not b;
    layer4_outputs(6575) <= a or b;
    layer4_outputs(6576) <= a;
    layer4_outputs(6577) <= b;
    layer4_outputs(6578) <= b and not a;
    layer4_outputs(6579) <= not (a and b);
    layer4_outputs(6580) <= not b;
    layer4_outputs(6581) <= a;
    layer4_outputs(6582) <= a;
    layer4_outputs(6583) <= b;
    layer4_outputs(6584) <= a or b;
    layer4_outputs(6585) <= not a or b;
    layer4_outputs(6586) <= a xor b;
    layer4_outputs(6587) <= not b or a;
    layer4_outputs(6588) <= not b;
    layer4_outputs(6589) <= not b;
    layer4_outputs(6590) <= not (a xor b);
    layer4_outputs(6591) <= not (a and b);
    layer4_outputs(6592) <= not b or a;
    layer4_outputs(6593) <= a;
    layer4_outputs(6594) <= a;
    layer4_outputs(6595) <= not (a and b);
    layer4_outputs(6596) <= not (a or b);
    layer4_outputs(6597) <= a and b;
    layer4_outputs(6598) <= a and b;
    layer4_outputs(6599) <= a;
    layer4_outputs(6600) <= b;
    layer4_outputs(6601) <= not a or b;
    layer4_outputs(6602) <= a and b;
    layer4_outputs(6603) <= not (a or b);
    layer4_outputs(6604) <= not (a or b);
    layer4_outputs(6605) <= not b;
    layer4_outputs(6606) <= a or b;
    layer4_outputs(6607) <= a or b;
    layer4_outputs(6608) <= not (a or b);
    layer4_outputs(6609) <= not b;
    layer4_outputs(6610) <= not a;
    layer4_outputs(6611) <= not a;
    layer4_outputs(6612) <= not b;
    layer4_outputs(6613) <= a and b;
    layer4_outputs(6614) <= a;
    layer4_outputs(6615) <= not a;
    layer4_outputs(6616) <= not a;
    layer4_outputs(6617) <= not b;
    layer4_outputs(6618) <= not b or a;
    layer4_outputs(6619) <= a or b;
    layer4_outputs(6620) <= not a;
    layer4_outputs(6621) <= not b;
    layer4_outputs(6622) <= b and not a;
    layer4_outputs(6623) <= not (a or b);
    layer4_outputs(6624) <= 1'b1;
    layer4_outputs(6625) <= a xor b;
    layer4_outputs(6626) <= a xor b;
    layer4_outputs(6627) <= not b;
    layer4_outputs(6628) <= a xor b;
    layer4_outputs(6629) <= a and not b;
    layer4_outputs(6630) <= b and not a;
    layer4_outputs(6631) <= b and not a;
    layer4_outputs(6632) <= not (a xor b);
    layer4_outputs(6633) <= not (a xor b);
    layer4_outputs(6634) <= a and b;
    layer4_outputs(6635) <= not a;
    layer4_outputs(6636) <= not (a xor b);
    layer4_outputs(6637) <= a and b;
    layer4_outputs(6638) <= a;
    layer4_outputs(6639) <= a;
    layer4_outputs(6640) <= a or b;
    layer4_outputs(6641) <= not b;
    layer4_outputs(6642) <= not (a xor b);
    layer4_outputs(6643) <= a and not b;
    layer4_outputs(6644) <= not a;
    layer4_outputs(6645) <= a xor b;
    layer4_outputs(6646) <= b and not a;
    layer4_outputs(6647) <= a and b;
    layer4_outputs(6648) <= not (a xor b);
    layer4_outputs(6649) <= not (a xor b);
    layer4_outputs(6650) <= a;
    layer4_outputs(6651) <= a and b;
    layer4_outputs(6652) <= not (a or b);
    layer4_outputs(6653) <= not b or a;
    layer4_outputs(6654) <= not (a and b);
    layer4_outputs(6655) <= b and not a;
    layer4_outputs(6656) <= not b or a;
    layer4_outputs(6657) <= not (a xor b);
    layer4_outputs(6658) <= b and not a;
    layer4_outputs(6659) <= a or b;
    layer4_outputs(6660) <= not a;
    layer4_outputs(6661) <= not b;
    layer4_outputs(6662) <= not b;
    layer4_outputs(6663) <= not (a and b);
    layer4_outputs(6664) <= b and not a;
    layer4_outputs(6665) <= not b;
    layer4_outputs(6666) <= a;
    layer4_outputs(6667) <= b;
    layer4_outputs(6668) <= not a;
    layer4_outputs(6669) <= a;
    layer4_outputs(6670) <= not a;
    layer4_outputs(6671) <= a xor b;
    layer4_outputs(6672) <= not (a and b);
    layer4_outputs(6673) <= not b;
    layer4_outputs(6674) <= b and not a;
    layer4_outputs(6675) <= a and b;
    layer4_outputs(6676) <= a and b;
    layer4_outputs(6677) <= not b;
    layer4_outputs(6678) <= a and not b;
    layer4_outputs(6679) <= not (a xor b);
    layer4_outputs(6680) <= a;
    layer4_outputs(6681) <= a and not b;
    layer4_outputs(6682) <= a;
    layer4_outputs(6683) <= not a;
    layer4_outputs(6684) <= not b;
    layer4_outputs(6685) <= not b;
    layer4_outputs(6686) <= not a or b;
    layer4_outputs(6687) <= not a or b;
    layer4_outputs(6688) <= b;
    layer4_outputs(6689) <= not b;
    layer4_outputs(6690) <= not (a xor b);
    layer4_outputs(6691) <= not b or a;
    layer4_outputs(6692) <= not (a xor b);
    layer4_outputs(6693) <= a or b;
    layer4_outputs(6694) <= not a;
    layer4_outputs(6695) <= a and b;
    layer4_outputs(6696) <= a;
    layer4_outputs(6697) <= a xor b;
    layer4_outputs(6698) <= a and not b;
    layer4_outputs(6699) <= not (a or b);
    layer4_outputs(6700) <= a or b;
    layer4_outputs(6701) <= a and not b;
    layer4_outputs(6702) <= a;
    layer4_outputs(6703) <= not a;
    layer4_outputs(6704) <= a;
    layer4_outputs(6705) <= a and not b;
    layer4_outputs(6706) <= not (a xor b);
    layer4_outputs(6707) <= not a;
    layer4_outputs(6708) <= a;
    layer4_outputs(6709) <= not b or a;
    layer4_outputs(6710) <= a;
    layer4_outputs(6711) <= not b;
    layer4_outputs(6712) <= not b;
    layer4_outputs(6713) <= b;
    layer4_outputs(6714) <= not a;
    layer4_outputs(6715) <= a;
    layer4_outputs(6716) <= b;
    layer4_outputs(6717) <= not (a xor b);
    layer4_outputs(6718) <= not (a or b);
    layer4_outputs(6719) <= not b;
    layer4_outputs(6720) <= a xor b;
    layer4_outputs(6721) <= a xor b;
    layer4_outputs(6722) <= not b;
    layer4_outputs(6723) <= not (a or b);
    layer4_outputs(6724) <= not a;
    layer4_outputs(6725) <= not (a xor b);
    layer4_outputs(6726) <= not (a xor b);
    layer4_outputs(6727) <= 1'b1;
    layer4_outputs(6728) <= not a;
    layer4_outputs(6729) <= a xor b;
    layer4_outputs(6730) <= not b;
    layer4_outputs(6731) <= not b;
    layer4_outputs(6732) <= a xor b;
    layer4_outputs(6733) <= not (a xor b);
    layer4_outputs(6734) <= not (a and b);
    layer4_outputs(6735) <= not (a xor b);
    layer4_outputs(6736) <= not a;
    layer4_outputs(6737) <= not (a or b);
    layer4_outputs(6738) <= not (a or b);
    layer4_outputs(6739) <= not (a xor b);
    layer4_outputs(6740) <= not a;
    layer4_outputs(6741) <= a and not b;
    layer4_outputs(6742) <= not (a and b);
    layer4_outputs(6743) <= not (a or b);
    layer4_outputs(6744) <= not (a and b);
    layer4_outputs(6745) <= b and not a;
    layer4_outputs(6746) <= a or b;
    layer4_outputs(6747) <= not a;
    layer4_outputs(6748) <= a and not b;
    layer4_outputs(6749) <= not (a or b);
    layer4_outputs(6750) <= not (a and b);
    layer4_outputs(6751) <= not b or a;
    layer4_outputs(6752) <= not a;
    layer4_outputs(6753) <= not a;
    layer4_outputs(6754) <= b and not a;
    layer4_outputs(6755) <= b;
    layer4_outputs(6756) <= a;
    layer4_outputs(6757) <= not b;
    layer4_outputs(6758) <= a;
    layer4_outputs(6759) <= a and b;
    layer4_outputs(6760) <= b;
    layer4_outputs(6761) <= not (a and b);
    layer4_outputs(6762) <= not b or a;
    layer4_outputs(6763) <= not b or a;
    layer4_outputs(6764) <= b and not a;
    layer4_outputs(6765) <= b and not a;
    layer4_outputs(6766) <= a xor b;
    layer4_outputs(6767) <= not b or a;
    layer4_outputs(6768) <= a;
    layer4_outputs(6769) <= not b;
    layer4_outputs(6770) <= not b;
    layer4_outputs(6771) <= not b;
    layer4_outputs(6772) <= not b or a;
    layer4_outputs(6773) <= b;
    layer4_outputs(6774) <= a;
    layer4_outputs(6775) <= b;
    layer4_outputs(6776) <= 1'b0;
    layer4_outputs(6777) <= not b;
    layer4_outputs(6778) <= not a or b;
    layer4_outputs(6779) <= not a or b;
    layer4_outputs(6780) <= not (a and b);
    layer4_outputs(6781) <= b and not a;
    layer4_outputs(6782) <= a;
    layer4_outputs(6783) <= a;
    layer4_outputs(6784) <= b and not a;
    layer4_outputs(6785) <= not b;
    layer4_outputs(6786) <= not b;
    layer4_outputs(6787) <= not a;
    layer4_outputs(6788) <= b;
    layer4_outputs(6789) <= a;
    layer4_outputs(6790) <= a or b;
    layer4_outputs(6791) <= not (a or b);
    layer4_outputs(6792) <= b;
    layer4_outputs(6793) <= not b;
    layer4_outputs(6794) <= a and b;
    layer4_outputs(6795) <= not b or a;
    layer4_outputs(6796) <= not a;
    layer4_outputs(6797) <= a and not b;
    layer4_outputs(6798) <= not a or b;
    layer4_outputs(6799) <= a;
    layer4_outputs(6800) <= not (a xor b);
    layer4_outputs(6801) <= a and not b;
    layer4_outputs(6802) <= not (a xor b);
    layer4_outputs(6803) <= a xor b;
    layer4_outputs(6804) <= b and not a;
    layer4_outputs(6805) <= a;
    layer4_outputs(6806) <= a and b;
    layer4_outputs(6807) <= b;
    layer4_outputs(6808) <= a and b;
    layer4_outputs(6809) <= not (a xor b);
    layer4_outputs(6810) <= not b;
    layer4_outputs(6811) <= a or b;
    layer4_outputs(6812) <= not (a and b);
    layer4_outputs(6813) <= not a;
    layer4_outputs(6814) <= b;
    layer4_outputs(6815) <= not a or b;
    layer4_outputs(6816) <= a xor b;
    layer4_outputs(6817) <= b and not a;
    layer4_outputs(6818) <= a and b;
    layer4_outputs(6819) <= not (a and b);
    layer4_outputs(6820) <= not (a or b);
    layer4_outputs(6821) <= a xor b;
    layer4_outputs(6822) <= not b or a;
    layer4_outputs(6823) <= a;
    layer4_outputs(6824) <= 1'b1;
    layer4_outputs(6825) <= b and not a;
    layer4_outputs(6826) <= a or b;
    layer4_outputs(6827) <= not b or a;
    layer4_outputs(6828) <= not b;
    layer4_outputs(6829) <= not b;
    layer4_outputs(6830) <= a or b;
    layer4_outputs(6831) <= a and b;
    layer4_outputs(6832) <= a and not b;
    layer4_outputs(6833) <= b and not a;
    layer4_outputs(6834) <= not a;
    layer4_outputs(6835) <= not a;
    layer4_outputs(6836) <= not b;
    layer4_outputs(6837) <= not b;
    layer4_outputs(6838) <= not b;
    layer4_outputs(6839) <= not a;
    layer4_outputs(6840) <= b;
    layer4_outputs(6841) <= a and not b;
    layer4_outputs(6842) <= a;
    layer4_outputs(6843) <= a and not b;
    layer4_outputs(6844) <= not (a xor b);
    layer4_outputs(6845) <= a xor b;
    layer4_outputs(6846) <= not a;
    layer4_outputs(6847) <= not a;
    layer4_outputs(6848) <= a;
    layer4_outputs(6849) <= not b;
    layer4_outputs(6850) <= not (a and b);
    layer4_outputs(6851) <= a xor b;
    layer4_outputs(6852) <= a xor b;
    layer4_outputs(6853) <= not b or a;
    layer4_outputs(6854) <= 1'b1;
    layer4_outputs(6855) <= not b;
    layer4_outputs(6856) <= a;
    layer4_outputs(6857) <= not b or a;
    layer4_outputs(6858) <= not a or b;
    layer4_outputs(6859) <= not b;
    layer4_outputs(6860) <= not (a and b);
    layer4_outputs(6861) <= a and not b;
    layer4_outputs(6862) <= not b or a;
    layer4_outputs(6863) <= a and not b;
    layer4_outputs(6864) <= not a;
    layer4_outputs(6865) <= not (a or b);
    layer4_outputs(6866) <= a;
    layer4_outputs(6867) <= not (a xor b);
    layer4_outputs(6868) <= not (a xor b);
    layer4_outputs(6869) <= b and not a;
    layer4_outputs(6870) <= not b;
    layer4_outputs(6871) <= not a;
    layer4_outputs(6872) <= not (a or b);
    layer4_outputs(6873) <= a xor b;
    layer4_outputs(6874) <= a and not b;
    layer4_outputs(6875) <= a and b;
    layer4_outputs(6876) <= not b or a;
    layer4_outputs(6877) <= a;
    layer4_outputs(6878) <= not b;
    layer4_outputs(6879) <= b;
    layer4_outputs(6880) <= a xor b;
    layer4_outputs(6881) <= not b;
    layer4_outputs(6882) <= a and b;
    layer4_outputs(6883) <= not b;
    layer4_outputs(6884) <= a xor b;
    layer4_outputs(6885) <= not b;
    layer4_outputs(6886) <= a;
    layer4_outputs(6887) <= not (a and b);
    layer4_outputs(6888) <= not b;
    layer4_outputs(6889) <= not (a or b);
    layer4_outputs(6890) <= not (a or b);
    layer4_outputs(6891) <= a and b;
    layer4_outputs(6892) <= not (a or b);
    layer4_outputs(6893) <= not a;
    layer4_outputs(6894) <= a xor b;
    layer4_outputs(6895) <= not a;
    layer4_outputs(6896) <= not b;
    layer4_outputs(6897) <= not b or a;
    layer4_outputs(6898) <= a and b;
    layer4_outputs(6899) <= a xor b;
    layer4_outputs(6900) <= a and not b;
    layer4_outputs(6901) <= not a;
    layer4_outputs(6902) <= not b or a;
    layer4_outputs(6903) <= a;
    layer4_outputs(6904) <= a xor b;
    layer4_outputs(6905) <= not a;
    layer4_outputs(6906) <= not a;
    layer4_outputs(6907) <= not (a xor b);
    layer4_outputs(6908) <= a xor b;
    layer4_outputs(6909) <= not (a or b);
    layer4_outputs(6910) <= a;
    layer4_outputs(6911) <= b;
    layer4_outputs(6912) <= b;
    layer4_outputs(6913) <= not a;
    layer4_outputs(6914) <= b;
    layer4_outputs(6915) <= a;
    layer4_outputs(6916) <= not a;
    layer4_outputs(6917) <= a and b;
    layer4_outputs(6918) <= a;
    layer4_outputs(6919) <= not (a or b);
    layer4_outputs(6920) <= not (a or b);
    layer4_outputs(6921) <= a;
    layer4_outputs(6922) <= a;
    layer4_outputs(6923) <= b;
    layer4_outputs(6924) <= not (a and b);
    layer4_outputs(6925) <= not b or a;
    layer4_outputs(6926) <= a xor b;
    layer4_outputs(6927) <= not (a or b);
    layer4_outputs(6928) <= not (a xor b);
    layer4_outputs(6929) <= b;
    layer4_outputs(6930) <= a;
    layer4_outputs(6931) <= not a or b;
    layer4_outputs(6932) <= not b;
    layer4_outputs(6933) <= a and b;
    layer4_outputs(6934) <= a xor b;
    layer4_outputs(6935) <= a and not b;
    layer4_outputs(6936) <= not b;
    layer4_outputs(6937) <= a and b;
    layer4_outputs(6938) <= a and not b;
    layer4_outputs(6939) <= b;
    layer4_outputs(6940) <= a or b;
    layer4_outputs(6941) <= a;
    layer4_outputs(6942) <= not b;
    layer4_outputs(6943) <= not b;
    layer4_outputs(6944) <= not (a xor b);
    layer4_outputs(6945) <= not b or a;
    layer4_outputs(6946) <= a;
    layer4_outputs(6947) <= a;
    layer4_outputs(6948) <= b;
    layer4_outputs(6949) <= not b or a;
    layer4_outputs(6950) <= not a;
    layer4_outputs(6951) <= a xor b;
    layer4_outputs(6952) <= b;
    layer4_outputs(6953) <= not (a or b);
    layer4_outputs(6954) <= b and not a;
    layer4_outputs(6955) <= b;
    layer4_outputs(6956) <= not a;
    layer4_outputs(6957) <= a xor b;
    layer4_outputs(6958) <= not (a and b);
    layer4_outputs(6959) <= a;
    layer4_outputs(6960) <= a or b;
    layer4_outputs(6961) <= a xor b;
    layer4_outputs(6962) <= a or b;
    layer4_outputs(6963) <= a;
    layer4_outputs(6964) <= not (a or b);
    layer4_outputs(6965) <= b;
    layer4_outputs(6966) <= not (a xor b);
    layer4_outputs(6967) <= a xor b;
    layer4_outputs(6968) <= not a;
    layer4_outputs(6969) <= a;
    layer4_outputs(6970) <= not (a xor b);
    layer4_outputs(6971) <= not (a xor b);
    layer4_outputs(6972) <= not (a xor b);
    layer4_outputs(6973) <= not (a or b);
    layer4_outputs(6974) <= a;
    layer4_outputs(6975) <= b;
    layer4_outputs(6976) <= not (a or b);
    layer4_outputs(6977) <= not b;
    layer4_outputs(6978) <= not (a or b);
    layer4_outputs(6979) <= not b;
    layer4_outputs(6980) <= not a;
    layer4_outputs(6981) <= a and not b;
    layer4_outputs(6982) <= a xor b;
    layer4_outputs(6983) <= not b;
    layer4_outputs(6984) <= not (a xor b);
    layer4_outputs(6985) <= not (a or b);
    layer4_outputs(6986) <= not (a and b);
    layer4_outputs(6987) <= a;
    layer4_outputs(6988) <= a and not b;
    layer4_outputs(6989) <= not a;
    layer4_outputs(6990) <= not a or b;
    layer4_outputs(6991) <= a and not b;
    layer4_outputs(6992) <= not a;
    layer4_outputs(6993) <= not (a or b);
    layer4_outputs(6994) <= a xor b;
    layer4_outputs(6995) <= a and not b;
    layer4_outputs(6996) <= a xor b;
    layer4_outputs(6997) <= a;
    layer4_outputs(6998) <= b and not a;
    layer4_outputs(6999) <= a and b;
    layer4_outputs(7000) <= a xor b;
    layer4_outputs(7001) <= not b;
    layer4_outputs(7002) <= not (a and b);
    layer4_outputs(7003) <= a;
    layer4_outputs(7004) <= not (a xor b);
    layer4_outputs(7005) <= a xor b;
    layer4_outputs(7006) <= not a or b;
    layer4_outputs(7007) <= a and b;
    layer4_outputs(7008) <= a;
    layer4_outputs(7009) <= a;
    layer4_outputs(7010) <= not b;
    layer4_outputs(7011) <= not (a and b);
    layer4_outputs(7012) <= a;
    layer4_outputs(7013) <= not a;
    layer4_outputs(7014) <= a;
    layer4_outputs(7015) <= a and not b;
    layer4_outputs(7016) <= not b;
    layer4_outputs(7017) <= a and b;
    layer4_outputs(7018) <= not b;
    layer4_outputs(7019) <= not a;
    layer4_outputs(7020) <= a;
    layer4_outputs(7021) <= not a or b;
    layer4_outputs(7022) <= not a;
    layer4_outputs(7023) <= b;
    layer4_outputs(7024) <= a xor b;
    layer4_outputs(7025) <= a or b;
    layer4_outputs(7026) <= not (a xor b);
    layer4_outputs(7027) <= a;
    layer4_outputs(7028) <= not (a or b);
    layer4_outputs(7029) <= not a;
    layer4_outputs(7030) <= a or b;
    layer4_outputs(7031) <= not (a or b);
    layer4_outputs(7032) <= b and not a;
    layer4_outputs(7033) <= a xor b;
    layer4_outputs(7034) <= b;
    layer4_outputs(7035) <= b and not a;
    layer4_outputs(7036) <= b;
    layer4_outputs(7037) <= a xor b;
    layer4_outputs(7038) <= b;
    layer4_outputs(7039) <= not (a xor b);
    layer4_outputs(7040) <= b;
    layer4_outputs(7041) <= a xor b;
    layer4_outputs(7042) <= not b or a;
    layer4_outputs(7043) <= not (a or b);
    layer4_outputs(7044) <= not (a and b);
    layer4_outputs(7045) <= not b;
    layer4_outputs(7046) <= a xor b;
    layer4_outputs(7047) <= a xor b;
    layer4_outputs(7048) <= not (a and b);
    layer4_outputs(7049) <= not (a xor b);
    layer4_outputs(7050) <= b;
    layer4_outputs(7051) <= not a;
    layer4_outputs(7052) <= b and not a;
    layer4_outputs(7053) <= not b;
    layer4_outputs(7054) <= b and not a;
    layer4_outputs(7055) <= not a or b;
    layer4_outputs(7056) <= a xor b;
    layer4_outputs(7057) <= not (a and b);
    layer4_outputs(7058) <= not b;
    layer4_outputs(7059) <= a;
    layer4_outputs(7060) <= a or b;
    layer4_outputs(7061) <= not (a xor b);
    layer4_outputs(7062) <= not a;
    layer4_outputs(7063) <= a and b;
    layer4_outputs(7064) <= not (a and b);
    layer4_outputs(7065) <= not a;
    layer4_outputs(7066) <= not (a and b);
    layer4_outputs(7067) <= a and not b;
    layer4_outputs(7068) <= not (a xor b);
    layer4_outputs(7069) <= not b;
    layer4_outputs(7070) <= b and not a;
    layer4_outputs(7071) <= a and b;
    layer4_outputs(7072) <= not (a and b);
    layer4_outputs(7073) <= not (a and b);
    layer4_outputs(7074) <= not b;
    layer4_outputs(7075) <= b;
    layer4_outputs(7076) <= b;
    layer4_outputs(7077) <= a and b;
    layer4_outputs(7078) <= not (a or b);
    layer4_outputs(7079) <= not b or a;
    layer4_outputs(7080) <= not a or b;
    layer4_outputs(7081) <= a xor b;
    layer4_outputs(7082) <= not a;
    layer4_outputs(7083) <= b;
    layer4_outputs(7084) <= a xor b;
    layer4_outputs(7085) <= not a or b;
    layer4_outputs(7086) <= not a;
    layer4_outputs(7087) <= b;
    layer4_outputs(7088) <= not (a or b);
    layer4_outputs(7089) <= b;
    layer4_outputs(7090) <= b;
    layer4_outputs(7091) <= b;
    layer4_outputs(7092) <= a;
    layer4_outputs(7093) <= not b or a;
    layer4_outputs(7094) <= not b;
    layer4_outputs(7095) <= a;
    layer4_outputs(7096) <= not a or b;
    layer4_outputs(7097) <= b and not a;
    layer4_outputs(7098) <= a;
    layer4_outputs(7099) <= a;
    layer4_outputs(7100) <= not (a or b);
    layer4_outputs(7101) <= a xor b;
    layer4_outputs(7102) <= a and not b;
    layer4_outputs(7103) <= not (a or b);
    layer4_outputs(7104) <= b;
    layer4_outputs(7105) <= not (a and b);
    layer4_outputs(7106) <= a and b;
    layer4_outputs(7107) <= b and not a;
    layer4_outputs(7108) <= b;
    layer4_outputs(7109) <= b and not a;
    layer4_outputs(7110) <= not (a xor b);
    layer4_outputs(7111) <= b;
    layer4_outputs(7112) <= a;
    layer4_outputs(7113) <= not b or a;
    layer4_outputs(7114) <= a xor b;
    layer4_outputs(7115) <= a and not b;
    layer4_outputs(7116) <= not a or b;
    layer4_outputs(7117) <= not a;
    layer4_outputs(7118) <= b;
    layer4_outputs(7119) <= b;
    layer4_outputs(7120) <= not (a or b);
    layer4_outputs(7121) <= not a;
    layer4_outputs(7122) <= not (a and b);
    layer4_outputs(7123) <= not b;
    layer4_outputs(7124) <= a or b;
    layer4_outputs(7125) <= not a;
    layer4_outputs(7126) <= not b;
    layer4_outputs(7127) <= a xor b;
    layer4_outputs(7128) <= not a;
    layer4_outputs(7129) <= b;
    layer4_outputs(7130) <= not (a and b);
    layer4_outputs(7131) <= a or b;
    layer4_outputs(7132) <= a;
    layer4_outputs(7133) <= a;
    layer4_outputs(7134) <= a or b;
    layer4_outputs(7135) <= a;
    layer4_outputs(7136) <= not a;
    layer4_outputs(7137) <= not b;
    layer4_outputs(7138) <= a xor b;
    layer4_outputs(7139) <= a xor b;
    layer4_outputs(7140) <= a;
    layer4_outputs(7141) <= a or b;
    layer4_outputs(7142) <= a;
    layer4_outputs(7143) <= a xor b;
    layer4_outputs(7144) <= not b;
    layer4_outputs(7145) <= not b;
    layer4_outputs(7146) <= a or b;
    layer4_outputs(7147) <= not a or b;
    layer4_outputs(7148) <= not (a or b);
    layer4_outputs(7149) <= a xor b;
    layer4_outputs(7150) <= not (a xor b);
    layer4_outputs(7151) <= a;
    layer4_outputs(7152) <= a or b;
    layer4_outputs(7153) <= not b or a;
    layer4_outputs(7154) <= not a or b;
    layer4_outputs(7155) <= b and not a;
    layer4_outputs(7156) <= not b;
    layer4_outputs(7157) <= a xor b;
    layer4_outputs(7158) <= not (a xor b);
    layer4_outputs(7159) <= b;
    layer4_outputs(7160) <= a or b;
    layer4_outputs(7161) <= not (a and b);
    layer4_outputs(7162) <= b and not a;
    layer4_outputs(7163) <= a;
    layer4_outputs(7164) <= a xor b;
    layer4_outputs(7165) <= a;
    layer4_outputs(7166) <= a and not b;
    layer4_outputs(7167) <= a and not b;
    layer4_outputs(7168) <= a;
    layer4_outputs(7169) <= a;
    layer4_outputs(7170) <= not a or b;
    layer4_outputs(7171) <= a and not b;
    layer4_outputs(7172) <= a and b;
    layer4_outputs(7173) <= b and not a;
    layer4_outputs(7174) <= not a;
    layer4_outputs(7175) <= not (a and b);
    layer4_outputs(7176) <= not (a and b);
    layer4_outputs(7177) <= b and not a;
    layer4_outputs(7178) <= 1'b0;
    layer4_outputs(7179) <= not a;
    layer4_outputs(7180) <= not (a or b);
    layer4_outputs(7181) <= not (a or b);
    layer4_outputs(7182) <= b;
    layer4_outputs(7183) <= not b;
    layer4_outputs(7184) <= not a;
    layer4_outputs(7185) <= not (a or b);
    layer4_outputs(7186) <= not b;
    layer4_outputs(7187) <= not a;
    layer4_outputs(7188) <= b;
    layer4_outputs(7189) <= not b;
    layer4_outputs(7190) <= b and not a;
    layer4_outputs(7191) <= not (a xor b);
    layer4_outputs(7192) <= a and b;
    layer4_outputs(7193) <= a;
    layer4_outputs(7194) <= b and not a;
    layer4_outputs(7195) <= a xor b;
    layer4_outputs(7196) <= a or b;
    layer4_outputs(7197) <= not b;
    layer4_outputs(7198) <= not b or a;
    layer4_outputs(7199) <= a xor b;
    layer4_outputs(7200) <= not (a and b);
    layer4_outputs(7201) <= a;
    layer4_outputs(7202) <= not a;
    layer4_outputs(7203) <= a;
    layer4_outputs(7204) <= b;
    layer4_outputs(7205) <= not a;
    layer4_outputs(7206) <= not (a or b);
    layer4_outputs(7207) <= not b;
    layer4_outputs(7208) <= a;
    layer4_outputs(7209) <= a;
    layer4_outputs(7210) <= not a;
    layer4_outputs(7211) <= not a;
    layer4_outputs(7212) <= not b or a;
    layer4_outputs(7213) <= not a or b;
    layer4_outputs(7214) <= b;
    layer4_outputs(7215) <= a and not b;
    layer4_outputs(7216) <= a;
    layer4_outputs(7217) <= a and not b;
    layer4_outputs(7218) <= a xor b;
    layer4_outputs(7219) <= a xor b;
    layer4_outputs(7220) <= b;
    layer4_outputs(7221) <= a and not b;
    layer4_outputs(7222) <= not a or b;
    layer4_outputs(7223) <= a xor b;
    layer4_outputs(7224) <= not b;
    layer4_outputs(7225) <= not b;
    layer4_outputs(7226) <= a and not b;
    layer4_outputs(7227) <= not a;
    layer4_outputs(7228) <= a and b;
    layer4_outputs(7229) <= not (a xor b);
    layer4_outputs(7230) <= not b;
    layer4_outputs(7231) <= a and b;
    layer4_outputs(7232) <= not a;
    layer4_outputs(7233) <= a xor b;
    layer4_outputs(7234) <= a or b;
    layer4_outputs(7235) <= a and not b;
    layer4_outputs(7236) <= b;
    layer4_outputs(7237) <= a or b;
    layer4_outputs(7238) <= b and not a;
    layer4_outputs(7239) <= not b;
    layer4_outputs(7240) <= a and not b;
    layer4_outputs(7241) <= not a;
    layer4_outputs(7242) <= a xor b;
    layer4_outputs(7243) <= not (a xor b);
    layer4_outputs(7244) <= a and b;
    layer4_outputs(7245) <= b;
    layer4_outputs(7246) <= not a or b;
    layer4_outputs(7247) <= b and not a;
    layer4_outputs(7248) <= a or b;
    layer4_outputs(7249) <= b and not a;
    layer4_outputs(7250) <= not a;
    layer4_outputs(7251) <= b and not a;
    layer4_outputs(7252) <= not (a xor b);
    layer4_outputs(7253) <= a;
    layer4_outputs(7254) <= a xor b;
    layer4_outputs(7255) <= a;
    layer4_outputs(7256) <= a and not b;
    layer4_outputs(7257) <= a xor b;
    layer4_outputs(7258) <= not (a or b);
    layer4_outputs(7259) <= not b;
    layer4_outputs(7260) <= 1'b1;
    layer4_outputs(7261) <= not (a and b);
    layer4_outputs(7262) <= not (a and b);
    layer4_outputs(7263) <= a;
    layer4_outputs(7264) <= not a;
    layer4_outputs(7265) <= not (a or b);
    layer4_outputs(7266) <= not a or b;
    layer4_outputs(7267) <= a;
    layer4_outputs(7268) <= not a;
    layer4_outputs(7269) <= a and not b;
    layer4_outputs(7270) <= a and not b;
    layer4_outputs(7271) <= b;
    layer4_outputs(7272) <= not b;
    layer4_outputs(7273) <= a and b;
    layer4_outputs(7274) <= a;
    layer4_outputs(7275) <= a xor b;
    layer4_outputs(7276) <= a xor b;
    layer4_outputs(7277) <= b and not a;
    layer4_outputs(7278) <= a xor b;
    layer4_outputs(7279) <= not (a xor b);
    layer4_outputs(7280) <= not a;
    layer4_outputs(7281) <= b;
    layer4_outputs(7282) <= not (a xor b);
    layer4_outputs(7283) <= not (a xor b);
    layer4_outputs(7284) <= b;
    layer4_outputs(7285) <= not a;
    layer4_outputs(7286) <= not (a or b);
    layer4_outputs(7287) <= not b or a;
    layer4_outputs(7288) <= b and not a;
    layer4_outputs(7289) <= not (a and b);
    layer4_outputs(7290) <= b;
    layer4_outputs(7291) <= b and not a;
    layer4_outputs(7292) <= a xor b;
    layer4_outputs(7293) <= b;
    layer4_outputs(7294) <= a xor b;
    layer4_outputs(7295) <= not a;
    layer4_outputs(7296) <= not b;
    layer4_outputs(7297) <= not (a or b);
    layer4_outputs(7298) <= b;
    layer4_outputs(7299) <= not a;
    layer4_outputs(7300) <= a xor b;
    layer4_outputs(7301) <= a and not b;
    layer4_outputs(7302) <= not b;
    layer4_outputs(7303) <= not (a xor b);
    layer4_outputs(7304) <= not b;
    layer4_outputs(7305) <= not (a or b);
    layer4_outputs(7306) <= not b;
    layer4_outputs(7307) <= a and b;
    layer4_outputs(7308) <= not a;
    layer4_outputs(7309) <= a;
    layer4_outputs(7310) <= not a;
    layer4_outputs(7311) <= not a;
    layer4_outputs(7312) <= a xor b;
    layer4_outputs(7313) <= a;
    layer4_outputs(7314) <= b;
    layer4_outputs(7315) <= not (a and b);
    layer4_outputs(7316) <= b;
    layer4_outputs(7317) <= not (a or b);
    layer4_outputs(7318) <= not (a xor b);
    layer4_outputs(7319) <= a xor b;
    layer4_outputs(7320) <= not (a or b);
    layer4_outputs(7321) <= a xor b;
    layer4_outputs(7322) <= a and not b;
    layer4_outputs(7323) <= not a or b;
    layer4_outputs(7324) <= not a or b;
    layer4_outputs(7325) <= not a;
    layer4_outputs(7326) <= b;
    layer4_outputs(7327) <= not a or b;
    layer4_outputs(7328) <= a and not b;
    layer4_outputs(7329) <= not a or b;
    layer4_outputs(7330) <= not b or a;
    layer4_outputs(7331) <= b and not a;
    layer4_outputs(7332) <= not (a xor b);
    layer4_outputs(7333) <= a xor b;
    layer4_outputs(7334) <= b;
    layer4_outputs(7335) <= a and b;
    layer4_outputs(7336) <= b;
    layer4_outputs(7337) <= not (a xor b);
    layer4_outputs(7338) <= not b or a;
    layer4_outputs(7339) <= not a;
    layer4_outputs(7340) <= not b;
    layer4_outputs(7341) <= not a;
    layer4_outputs(7342) <= a and b;
    layer4_outputs(7343) <= not b or a;
    layer4_outputs(7344) <= b and not a;
    layer4_outputs(7345) <= a and b;
    layer4_outputs(7346) <= b and not a;
    layer4_outputs(7347) <= not b or a;
    layer4_outputs(7348) <= a and not b;
    layer4_outputs(7349) <= a xor b;
    layer4_outputs(7350) <= not a;
    layer4_outputs(7351) <= not (a and b);
    layer4_outputs(7352) <= not a or b;
    layer4_outputs(7353) <= a;
    layer4_outputs(7354) <= not b;
    layer4_outputs(7355) <= a xor b;
    layer4_outputs(7356) <= a and not b;
    layer4_outputs(7357) <= a xor b;
    layer4_outputs(7358) <= not (a xor b);
    layer4_outputs(7359) <= b and not a;
    layer4_outputs(7360) <= not b;
    layer4_outputs(7361) <= a and b;
    layer4_outputs(7362) <= a and b;
    layer4_outputs(7363) <= a and b;
    layer4_outputs(7364) <= not b;
    layer4_outputs(7365) <= not b;
    layer4_outputs(7366) <= 1'b0;
    layer4_outputs(7367) <= a or b;
    layer4_outputs(7368) <= not b or a;
    layer4_outputs(7369) <= a;
    layer4_outputs(7370) <= a xor b;
    layer4_outputs(7371) <= a and b;
    layer4_outputs(7372) <= a and b;
    layer4_outputs(7373) <= not (a xor b);
    layer4_outputs(7374) <= not (a xor b);
    layer4_outputs(7375) <= a and b;
    layer4_outputs(7376) <= a;
    layer4_outputs(7377) <= a xor b;
    layer4_outputs(7378) <= 1'b0;
    layer4_outputs(7379) <= not a;
    layer4_outputs(7380) <= b and not a;
    layer4_outputs(7381) <= a xor b;
    layer4_outputs(7382) <= not b;
    layer4_outputs(7383) <= not (a or b);
    layer4_outputs(7384) <= not b;
    layer4_outputs(7385) <= not (a xor b);
    layer4_outputs(7386) <= a or b;
    layer4_outputs(7387) <= b;
    layer4_outputs(7388) <= a;
    layer4_outputs(7389) <= not (a or b);
    layer4_outputs(7390) <= a and b;
    layer4_outputs(7391) <= not a;
    layer4_outputs(7392) <= not b;
    layer4_outputs(7393) <= b;
    layer4_outputs(7394) <= b;
    layer4_outputs(7395) <= a;
    layer4_outputs(7396) <= not a;
    layer4_outputs(7397) <= a;
    layer4_outputs(7398) <= not b or a;
    layer4_outputs(7399) <= b;
    layer4_outputs(7400) <= not (a xor b);
    layer4_outputs(7401) <= a;
    layer4_outputs(7402) <= not b;
    layer4_outputs(7403) <= not (a xor b);
    layer4_outputs(7404) <= a xor b;
    layer4_outputs(7405) <= a;
    layer4_outputs(7406) <= a and b;
    layer4_outputs(7407) <= b;
    layer4_outputs(7408) <= not (a and b);
    layer4_outputs(7409) <= not b;
    layer4_outputs(7410) <= not a;
    layer4_outputs(7411) <= a and b;
    layer4_outputs(7412) <= a and b;
    layer4_outputs(7413) <= a or b;
    layer4_outputs(7414) <= a xor b;
    layer4_outputs(7415) <= not b;
    layer4_outputs(7416) <= not a;
    layer4_outputs(7417) <= not a;
    layer4_outputs(7418) <= b;
    layer4_outputs(7419) <= not (a or b);
    layer4_outputs(7420) <= a and not b;
    layer4_outputs(7421) <= not (a or b);
    layer4_outputs(7422) <= a and b;
    layer4_outputs(7423) <= a xor b;
    layer4_outputs(7424) <= a xor b;
    layer4_outputs(7425) <= not a;
    layer4_outputs(7426) <= not (a xor b);
    layer4_outputs(7427) <= a and not b;
    layer4_outputs(7428) <= a;
    layer4_outputs(7429) <= not (a xor b);
    layer4_outputs(7430) <= a xor b;
    layer4_outputs(7431) <= 1'b1;
    layer4_outputs(7432) <= not (a xor b);
    layer4_outputs(7433) <= a and not b;
    layer4_outputs(7434) <= not b or a;
    layer4_outputs(7435) <= b;
    layer4_outputs(7436) <= not (a xor b);
    layer4_outputs(7437) <= not b;
    layer4_outputs(7438) <= not b;
    layer4_outputs(7439) <= a xor b;
    layer4_outputs(7440) <= 1'b1;
    layer4_outputs(7441) <= not a or b;
    layer4_outputs(7442) <= b;
    layer4_outputs(7443) <= 1'b0;
    layer4_outputs(7444) <= a;
    layer4_outputs(7445) <= b;
    layer4_outputs(7446) <= not b or a;
    layer4_outputs(7447) <= not (a xor b);
    layer4_outputs(7448) <= b;
    layer4_outputs(7449) <= b;
    layer4_outputs(7450) <= a;
    layer4_outputs(7451) <= a;
    layer4_outputs(7452) <= a and not b;
    layer4_outputs(7453) <= b;
    layer4_outputs(7454) <= not b or a;
    layer4_outputs(7455) <= not (a and b);
    layer4_outputs(7456) <= a;
    layer4_outputs(7457) <= a and b;
    layer4_outputs(7458) <= not a or b;
    layer4_outputs(7459) <= not (a xor b);
    layer4_outputs(7460) <= a or b;
    layer4_outputs(7461) <= not (a xor b);
    layer4_outputs(7462) <= not a or b;
    layer4_outputs(7463) <= not (a and b);
    layer4_outputs(7464) <= not (a and b);
    layer4_outputs(7465) <= a;
    layer4_outputs(7466) <= a;
    layer4_outputs(7467) <= a xor b;
    layer4_outputs(7468) <= b;
    layer4_outputs(7469) <= a;
    layer4_outputs(7470) <= not a;
    layer4_outputs(7471) <= a;
    layer4_outputs(7472) <= not (a and b);
    layer4_outputs(7473) <= a;
    layer4_outputs(7474) <= not (a and b);
    layer4_outputs(7475) <= a and b;
    layer4_outputs(7476) <= b;
    layer4_outputs(7477) <= not a;
    layer4_outputs(7478) <= not (a or b);
    layer4_outputs(7479) <= not (a xor b);
    layer4_outputs(7480) <= not b or a;
    layer4_outputs(7481) <= b;
    layer4_outputs(7482) <= a and not b;
    layer4_outputs(7483) <= not a;
    layer4_outputs(7484) <= a;
    layer4_outputs(7485) <= a or b;
    layer4_outputs(7486) <= a;
    layer4_outputs(7487) <= not b or a;
    layer4_outputs(7488) <= a xor b;
    layer4_outputs(7489) <= not (a and b);
    layer4_outputs(7490) <= not (a or b);
    layer4_outputs(7491) <= not (a or b);
    layer4_outputs(7492) <= a and b;
    layer4_outputs(7493) <= a;
    layer4_outputs(7494) <= not (a or b);
    layer4_outputs(7495) <= not a;
    layer4_outputs(7496) <= not b or a;
    layer4_outputs(7497) <= a;
    layer4_outputs(7498) <= not (a xor b);
    layer4_outputs(7499) <= a and b;
    layer4_outputs(7500) <= a and b;
    layer4_outputs(7501) <= not a;
    layer4_outputs(7502) <= not b or a;
    layer4_outputs(7503) <= not a;
    layer4_outputs(7504) <= a and b;
    layer4_outputs(7505) <= not a;
    layer4_outputs(7506) <= a xor b;
    layer4_outputs(7507) <= b;
    layer4_outputs(7508) <= b;
    layer4_outputs(7509) <= not b;
    layer4_outputs(7510) <= not b or a;
    layer4_outputs(7511) <= not a;
    layer4_outputs(7512) <= a;
    layer4_outputs(7513) <= a;
    layer4_outputs(7514) <= not a or b;
    layer4_outputs(7515) <= not (a xor b);
    layer4_outputs(7516) <= not a;
    layer4_outputs(7517) <= a or b;
    layer4_outputs(7518) <= not a;
    layer4_outputs(7519) <= not a;
    layer4_outputs(7520) <= a;
    layer4_outputs(7521) <= a and b;
    layer4_outputs(7522) <= a;
    layer4_outputs(7523) <= not a;
    layer4_outputs(7524) <= not a;
    layer4_outputs(7525) <= not a;
    layer4_outputs(7526) <= a and b;
    layer4_outputs(7527) <= not b;
    layer4_outputs(7528) <= a;
    layer4_outputs(7529) <= a;
    layer4_outputs(7530) <= a and not b;
    layer4_outputs(7531) <= a xor b;
    layer4_outputs(7532) <= a;
    layer4_outputs(7533) <= not (a or b);
    layer4_outputs(7534) <= not (a xor b);
    layer4_outputs(7535) <= b;
    layer4_outputs(7536) <= 1'b1;
    layer4_outputs(7537) <= a;
    layer4_outputs(7538) <= b;
    layer4_outputs(7539) <= not b;
    layer4_outputs(7540) <= a xor b;
    layer4_outputs(7541) <= not a;
    layer4_outputs(7542) <= b and not a;
    layer4_outputs(7543) <= a;
    layer4_outputs(7544) <= a and not b;
    layer4_outputs(7545) <= a and b;
    layer4_outputs(7546) <= b;
    layer4_outputs(7547) <= b;
    layer4_outputs(7548) <= 1'b1;
    layer4_outputs(7549) <= a and not b;
    layer4_outputs(7550) <= b;
    layer4_outputs(7551) <= not a;
    layer4_outputs(7552) <= a and not b;
    layer4_outputs(7553) <= a and b;
    layer4_outputs(7554) <= a xor b;
    layer4_outputs(7555) <= not (a and b);
    layer4_outputs(7556) <= not (a and b);
    layer4_outputs(7557) <= b;
    layer4_outputs(7558) <= not b;
    layer4_outputs(7559) <= a;
    layer4_outputs(7560) <= not a;
    layer4_outputs(7561) <= a;
    layer4_outputs(7562) <= not b;
    layer4_outputs(7563) <= a xor b;
    layer4_outputs(7564) <= not b;
    layer4_outputs(7565) <= not a;
    layer4_outputs(7566) <= b;
    layer4_outputs(7567) <= not (a xor b);
    layer4_outputs(7568) <= b and not a;
    layer4_outputs(7569) <= a;
    layer4_outputs(7570) <= b and not a;
    layer4_outputs(7571) <= not b;
    layer4_outputs(7572) <= not a or b;
    layer4_outputs(7573) <= not a;
    layer4_outputs(7574) <= a or b;
    layer4_outputs(7575) <= not (a and b);
    layer4_outputs(7576) <= not (a xor b);
    layer4_outputs(7577) <= not b;
    layer4_outputs(7578) <= not a;
    layer4_outputs(7579) <= a or b;
    layer4_outputs(7580) <= not b;
    layer4_outputs(7581) <= not (a xor b);
    layer4_outputs(7582) <= b;
    layer4_outputs(7583) <= a or b;
    layer4_outputs(7584) <= b and not a;
    layer4_outputs(7585) <= not b;
    layer4_outputs(7586) <= not b;
    layer4_outputs(7587) <= a and b;
    layer4_outputs(7588) <= not b;
    layer4_outputs(7589) <= not (a or b);
    layer4_outputs(7590) <= a;
    layer4_outputs(7591) <= not a or b;
    layer4_outputs(7592) <= not b;
    layer4_outputs(7593) <= not b;
    layer4_outputs(7594) <= b and not a;
    layer4_outputs(7595) <= b and not a;
    layer4_outputs(7596) <= a;
    layer4_outputs(7597) <= a and b;
    layer4_outputs(7598) <= a;
    layer4_outputs(7599) <= b;
    layer4_outputs(7600) <= not (a xor b);
    layer4_outputs(7601) <= a or b;
    layer4_outputs(7602) <= not (a and b);
    layer4_outputs(7603) <= a and b;
    layer4_outputs(7604) <= not (a or b);
    layer4_outputs(7605) <= not b;
    layer4_outputs(7606) <= a and not b;
    layer4_outputs(7607) <= not (a xor b);
    layer4_outputs(7608) <= not a or b;
    layer4_outputs(7609) <= a;
    layer4_outputs(7610) <= a xor b;
    layer4_outputs(7611) <= not a;
    layer4_outputs(7612) <= not a or b;
    layer4_outputs(7613) <= not a;
    layer4_outputs(7614) <= not (a xor b);
    layer4_outputs(7615) <= b;
    layer4_outputs(7616) <= not b;
    layer4_outputs(7617) <= not (a xor b);
    layer4_outputs(7618) <= not (a xor b);
    layer4_outputs(7619) <= a and not b;
    layer4_outputs(7620) <= 1'b0;
    layer4_outputs(7621) <= a;
    layer4_outputs(7622) <= b;
    layer4_outputs(7623) <= a and not b;
    layer4_outputs(7624) <= not a;
    layer4_outputs(7625) <= a and b;
    layer4_outputs(7626) <= a and not b;
    layer4_outputs(7627) <= b;
    layer4_outputs(7628) <= not b;
    layer4_outputs(7629) <= not b;
    layer4_outputs(7630) <= not a;
    layer4_outputs(7631) <= not a;
    layer4_outputs(7632) <= a and b;
    layer4_outputs(7633) <= a xor b;
    layer4_outputs(7634) <= b and not a;
    layer4_outputs(7635) <= not (a and b);
    layer4_outputs(7636) <= not (a or b);
    layer4_outputs(7637) <= a;
    layer4_outputs(7638) <= not a;
    layer4_outputs(7639) <= a;
    layer4_outputs(7640) <= not (a xor b);
    layer4_outputs(7641) <= 1'b1;
    layer4_outputs(7642) <= a and b;
    layer4_outputs(7643) <= not b;
    layer4_outputs(7644) <= a;
    layer4_outputs(7645) <= b;
    layer4_outputs(7646) <= not (a xor b);
    layer4_outputs(7647) <= a;
    layer4_outputs(7648) <= a or b;
    layer4_outputs(7649) <= not (a or b);
    layer4_outputs(7650) <= not b;
    layer4_outputs(7651) <= not a or b;
    layer4_outputs(7652) <= a and b;
    layer4_outputs(7653) <= b and not a;
    layer4_outputs(7654) <= a;
    layer4_outputs(7655) <= not b;
    layer4_outputs(7656) <= a xor b;
    layer4_outputs(7657) <= a xor b;
    layer4_outputs(7658) <= a and not b;
    layer4_outputs(7659) <= not (a xor b);
    layer4_outputs(7660) <= b;
    layer4_outputs(7661) <= a or b;
    layer4_outputs(7662) <= a;
    layer4_outputs(7663) <= a xor b;
    layer4_outputs(7664) <= not b;
    layer4_outputs(7665) <= a;
    layer4_outputs(7666) <= a;
    layer4_outputs(7667) <= a xor b;
    layer4_outputs(7668) <= b;
    layer4_outputs(7669) <= not b or a;
    layer4_outputs(7670) <= not a or b;
    layer4_outputs(7671) <= not (a xor b);
    layer4_outputs(7672) <= b;
    layer4_outputs(7673) <= not a;
    layer4_outputs(7674) <= not a or b;
    layer4_outputs(7675) <= not b or a;
    layer4_outputs(7676) <= not a;
    layer4_outputs(7677) <= not b;
    layer4_outputs(7678) <= a xor b;
    layer4_outputs(7679) <= not (a and b);
    layer4_outputs(7680) <= not a;
    layer4_outputs(7681) <= a xor b;
    layer4_outputs(7682) <= not a or b;
    layer4_outputs(7683) <= not b;
    layer4_outputs(7684) <= not b;
    layer4_outputs(7685) <= not (a and b);
    layer4_outputs(7686) <= not b;
    layer4_outputs(7687) <= b;
    layer4_outputs(7688) <= not a;
    layer4_outputs(7689) <= not a;
    layer4_outputs(7690) <= b;
    layer4_outputs(7691) <= a;
    layer4_outputs(7692) <= a and b;
    layer4_outputs(7693) <= not b or a;
    layer4_outputs(7694) <= a and b;
    layer4_outputs(7695) <= not a;
    layer4_outputs(7696) <= not (a xor b);
    layer4_outputs(7697) <= not a;
    layer4_outputs(7698) <= a;
    layer4_outputs(7699) <= a xor b;
    layer4_outputs(7700) <= not a;
    layer4_outputs(7701) <= a xor b;
    layer4_outputs(7702) <= not b;
    layer4_outputs(7703) <= a or b;
    layer4_outputs(7704) <= a;
    layer4_outputs(7705) <= a xor b;
    layer4_outputs(7706) <= a and not b;
    layer4_outputs(7707) <= a;
    layer4_outputs(7708) <= a;
    layer4_outputs(7709) <= not (a xor b);
    layer4_outputs(7710) <= a and b;
    layer4_outputs(7711) <= a;
    layer4_outputs(7712) <= a or b;
    layer4_outputs(7713) <= a and b;
    layer4_outputs(7714) <= a and b;
    layer4_outputs(7715) <= not b;
    layer4_outputs(7716) <= not b;
    layer4_outputs(7717) <= not a;
    layer4_outputs(7718) <= b and not a;
    layer4_outputs(7719) <= a or b;
    layer4_outputs(7720) <= not (a xor b);
    layer4_outputs(7721) <= a or b;
    layer4_outputs(7722) <= not a or b;
    layer4_outputs(7723) <= not (a or b);
    layer4_outputs(7724) <= a xor b;
    layer4_outputs(7725) <= not b;
    layer4_outputs(7726) <= b;
    layer4_outputs(7727) <= a or b;
    layer4_outputs(7728) <= a;
    layer4_outputs(7729) <= not (a xor b);
    layer4_outputs(7730) <= a;
    layer4_outputs(7731) <= not b;
    layer4_outputs(7732) <= not b;
    layer4_outputs(7733) <= a xor b;
    layer4_outputs(7734) <= a;
    layer4_outputs(7735) <= a and not b;
    layer4_outputs(7736) <= a and not b;
    layer4_outputs(7737) <= a xor b;
    layer4_outputs(7738) <= not (a or b);
    layer4_outputs(7739) <= not b;
    layer4_outputs(7740) <= a xor b;
    layer4_outputs(7741) <= not (a and b);
    layer4_outputs(7742) <= not b;
    layer4_outputs(7743) <= not (a and b);
    layer4_outputs(7744) <= not a;
    layer4_outputs(7745) <= not b;
    layer4_outputs(7746) <= 1'b0;
    layer4_outputs(7747) <= a xor b;
    layer4_outputs(7748) <= a;
    layer4_outputs(7749) <= a xor b;
    layer4_outputs(7750) <= a;
    layer4_outputs(7751) <= a xor b;
    layer4_outputs(7752) <= b;
    layer4_outputs(7753) <= not a;
    layer4_outputs(7754) <= not b or a;
    layer4_outputs(7755) <= a xor b;
    layer4_outputs(7756) <= a xor b;
    layer4_outputs(7757) <= a;
    layer4_outputs(7758) <= a or b;
    layer4_outputs(7759) <= not (a or b);
    layer4_outputs(7760) <= not b;
    layer4_outputs(7761) <= not (a xor b);
    layer4_outputs(7762) <= not b or a;
    layer4_outputs(7763) <= b;
    layer4_outputs(7764) <= a xor b;
    layer4_outputs(7765) <= a or b;
    layer4_outputs(7766) <= b;
    layer4_outputs(7767) <= not (a xor b);
    layer4_outputs(7768) <= b;
    layer4_outputs(7769) <= not a;
    layer4_outputs(7770) <= not (a xor b);
    layer4_outputs(7771) <= a;
    layer4_outputs(7772) <= not (a and b);
    layer4_outputs(7773) <= b;
    layer4_outputs(7774) <= not (a or b);
    layer4_outputs(7775) <= a xor b;
    layer4_outputs(7776) <= b;
    layer4_outputs(7777) <= b;
    layer4_outputs(7778) <= b;
    layer4_outputs(7779) <= not (a and b);
    layer4_outputs(7780) <= not a or b;
    layer4_outputs(7781) <= a and b;
    layer4_outputs(7782) <= b;
    layer4_outputs(7783) <= b;
    layer4_outputs(7784) <= a or b;
    layer4_outputs(7785) <= not (a xor b);
    layer4_outputs(7786) <= not b;
    layer4_outputs(7787) <= a xor b;
    layer4_outputs(7788) <= not (a xor b);
    layer4_outputs(7789) <= not a;
    layer4_outputs(7790) <= b;
    layer4_outputs(7791) <= b and not a;
    layer4_outputs(7792) <= a and b;
    layer4_outputs(7793) <= a;
    layer4_outputs(7794) <= not (a xor b);
    layer4_outputs(7795) <= b;
    layer4_outputs(7796) <= not (a or b);
    layer4_outputs(7797) <= a;
    layer4_outputs(7798) <= not b or a;
    layer4_outputs(7799) <= a;
    layer4_outputs(7800) <= not (a xor b);
    layer4_outputs(7801) <= not b or a;
    layer4_outputs(7802) <= not b;
    layer4_outputs(7803) <= a and not b;
    layer4_outputs(7804) <= not a or b;
    layer4_outputs(7805) <= not b or a;
    layer4_outputs(7806) <= not (a xor b);
    layer4_outputs(7807) <= b;
    layer4_outputs(7808) <= not b;
    layer4_outputs(7809) <= b;
    layer4_outputs(7810) <= 1'b1;
    layer4_outputs(7811) <= not b;
    layer4_outputs(7812) <= a;
    layer4_outputs(7813) <= a;
    layer4_outputs(7814) <= b;
    layer4_outputs(7815) <= not b or a;
    layer4_outputs(7816) <= not a;
    layer4_outputs(7817) <= not (a xor b);
    layer4_outputs(7818) <= not a;
    layer4_outputs(7819) <= not a or b;
    layer4_outputs(7820) <= b;
    layer4_outputs(7821) <= a or b;
    layer4_outputs(7822) <= not (a xor b);
    layer4_outputs(7823) <= a;
    layer4_outputs(7824) <= a;
    layer4_outputs(7825) <= not a or b;
    layer4_outputs(7826) <= a and b;
    layer4_outputs(7827) <= a xor b;
    layer4_outputs(7828) <= a and b;
    layer4_outputs(7829) <= not (a or b);
    layer4_outputs(7830) <= a or b;
    layer4_outputs(7831) <= b;
    layer4_outputs(7832) <= a and not b;
    layer4_outputs(7833) <= a and not b;
    layer4_outputs(7834) <= not b or a;
    layer4_outputs(7835) <= a and b;
    layer4_outputs(7836) <= a xor b;
    layer4_outputs(7837) <= b;
    layer4_outputs(7838) <= a or b;
    layer4_outputs(7839) <= not (a xor b);
    layer4_outputs(7840) <= b;
    layer4_outputs(7841) <= not b;
    layer4_outputs(7842) <= not (a or b);
    layer4_outputs(7843) <= not a;
    layer4_outputs(7844) <= not b or a;
    layer4_outputs(7845) <= not b or a;
    layer4_outputs(7846) <= a;
    layer4_outputs(7847) <= not a;
    layer4_outputs(7848) <= a xor b;
    layer4_outputs(7849) <= a;
    layer4_outputs(7850) <= not (a and b);
    layer4_outputs(7851) <= not a or b;
    layer4_outputs(7852) <= not b or a;
    layer4_outputs(7853) <= a xor b;
    layer4_outputs(7854) <= b;
    layer4_outputs(7855) <= not a;
    layer4_outputs(7856) <= a xor b;
    layer4_outputs(7857) <= not (a xor b);
    layer4_outputs(7858) <= not b or a;
    layer4_outputs(7859) <= a xor b;
    layer4_outputs(7860) <= not a;
    layer4_outputs(7861) <= a and not b;
    layer4_outputs(7862) <= a;
    layer4_outputs(7863) <= not b;
    layer4_outputs(7864) <= 1'b0;
    layer4_outputs(7865) <= a xor b;
    layer4_outputs(7866) <= not (a and b);
    layer4_outputs(7867) <= not (a xor b);
    layer4_outputs(7868) <= not b or a;
    layer4_outputs(7869) <= not (a xor b);
    layer4_outputs(7870) <= not (a and b);
    layer4_outputs(7871) <= b;
    layer4_outputs(7872) <= not b;
    layer4_outputs(7873) <= a;
    layer4_outputs(7874) <= not (a xor b);
    layer4_outputs(7875) <= a or b;
    layer4_outputs(7876) <= b;
    layer4_outputs(7877) <= b;
    layer4_outputs(7878) <= a and not b;
    layer4_outputs(7879) <= a and not b;
    layer4_outputs(7880) <= not b;
    layer4_outputs(7881) <= b;
    layer4_outputs(7882) <= not b;
    layer4_outputs(7883) <= not (a or b);
    layer4_outputs(7884) <= not a;
    layer4_outputs(7885) <= not (a or b);
    layer4_outputs(7886) <= a or b;
    layer4_outputs(7887) <= not a or b;
    layer4_outputs(7888) <= not (a xor b);
    layer4_outputs(7889) <= a xor b;
    layer4_outputs(7890) <= not a;
    layer4_outputs(7891) <= b;
    layer4_outputs(7892) <= a and not b;
    layer4_outputs(7893) <= a;
    layer4_outputs(7894) <= b and not a;
    layer4_outputs(7895) <= b;
    layer4_outputs(7896) <= not a;
    layer4_outputs(7897) <= not a;
    layer4_outputs(7898) <= a;
    layer4_outputs(7899) <= not a;
    layer4_outputs(7900) <= not b;
    layer4_outputs(7901) <= not (a and b);
    layer4_outputs(7902) <= not b;
    layer4_outputs(7903) <= not b;
    layer4_outputs(7904) <= not (a or b);
    layer4_outputs(7905) <= b and not a;
    layer4_outputs(7906) <= a and not b;
    layer4_outputs(7907) <= not (a xor b);
    layer4_outputs(7908) <= b and not a;
    layer4_outputs(7909) <= not a or b;
    layer4_outputs(7910) <= b and not a;
    layer4_outputs(7911) <= a;
    layer4_outputs(7912) <= not (a xor b);
    layer4_outputs(7913) <= b;
    layer4_outputs(7914) <= not b;
    layer4_outputs(7915) <= a xor b;
    layer4_outputs(7916) <= not b;
    layer4_outputs(7917) <= b;
    layer4_outputs(7918) <= not a;
    layer4_outputs(7919) <= not b or a;
    layer4_outputs(7920) <= not a;
    layer4_outputs(7921) <= not (a and b);
    layer4_outputs(7922) <= not b or a;
    layer4_outputs(7923) <= not (a xor b);
    layer4_outputs(7924) <= b;
    layer4_outputs(7925) <= not (a xor b);
    layer4_outputs(7926) <= not (a or b);
    layer4_outputs(7927) <= not a;
    layer4_outputs(7928) <= a;
    layer4_outputs(7929) <= not a;
    layer4_outputs(7930) <= b;
    layer4_outputs(7931) <= not b;
    layer4_outputs(7932) <= not b or a;
    layer4_outputs(7933) <= b;
    layer4_outputs(7934) <= not b or a;
    layer4_outputs(7935) <= not b or a;
    layer4_outputs(7936) <= a or b;
    layer4_outputs(7937) <= not (a xor b);
    layer4_outputs(7938) <= not a or b;
    layer4_outputs(7939) <= b and not a;
    layer4_outputs(7940) <= a;
    layer4_outputs(7941) <= a xor b;
    layer4_outputs(7942) <= b;
    layer4_outputs(7943) <= not (a xor b);
    layer4_outputs(7944) <= a xor b;
    layer4_outputs(7945) <= not b;
    layer4_outputs(7946) <= b and not a;
    layer4_outputs(7947) <= b;
    layer4_outputs(7948) <= b;
    layer4_outputs(7949) <= not b or a;
    layer4_outputs(7950) <= a xor b;
    layer4_outputs(7951) <= b;
    layer4_outputs(7952) <= not (a and b);
    layer4_outputs(7953) <= a or b;
    layer4_outputs(7954) <= not (a xor b);
    layer4_outputs(7955) <= a;
    layer4_outputs(7956) <= not b or a;
    layer4_outputs(7957) <= a;
    layer4_outputs(7958) <= a xor b;
    layer4_outputs(7959) <= a;
    layer4_outputs(7960) <= not b or a;
    layer4_outputs(7961) <= not (a or b);
    layer4_outputs(7962) <= not a or b;
    layer4_outputs(7963) <= b;
    layer4_outputs(7964) <= not b;
    layer4_outputs(7965) <= a or b;
    layer4_outputs(7966) <= a and b;
    layer4_outputs(7967) <= not b;
    layer4_outputs(7968) <= a xor b;
    layer4_outputs(7969) <= b;
    layer4_outputs(7970) <= a and b;
    layer4_outputs(7971) <= not (a and b);
    layer4_outputs(7972) <= a;
    layer4_outputs(7973) <= not a or b;
    layer4_outputs(7974) <= not a;
    layer4_outputs(7975) <= not b;
    layer4_outputs(7976) <= b;
    layer4_outputs(7977) <= not b;
    layer4_outputs(7978) <= not a;
    layer4_outputs(7979) <= not b;
    layer4_outputs(7980) <= not b or a;
    layer4_outputs(7981) <= not a or b;
    layer4_outputs(7982) <= not a;
    layer4_outputs(7983) <= not a;
    layer4_outputs(7984) <= not b;
    layer4_outputs(7985) <= a xor b;
    layer4_outputs(7986) <= not a;
    layer4_outputs(7987) <= not (a or b);
    layer4_outputs(7988) <= not (a xor b);
    layer4_outputs(7989) <= not (a and b);
    layer4_outputs(7990) <= not b or a;
    layer4_outputs(7991) <= b;
    layer4_outputs(7992) <= not a;
    layer4_outputs(7993) <= a;
    layer4_outputs(7994) <= not (a xor b);
    layer4_outputs(7995) <= b;
    layer4_outputs(7996) <= b and not a;
    layer4_outputs(7997) <= not b;
    layer4_outputs(7998) <= not b;
    layer4_outputs(7999) <= a and not b;
    layer4_outputs(8000) <= not b or a;
    layer4_outputs(8001) <= b and not a;
    layer4_outputs(8002) <= a xor b;
    layer4_outputs(8003) <= not (a xor b);
    layer4_outputs(8004) <= a xor b;
    layer4_outputs(8005) <= not b;
    layer4_outputs(8006) <= not b;
    layer4_outputs(8007) <= not b;
    layer4_outputs(8008) <= not (a and b);
    layer4_outputs(8009) <= not a or b;
    layer4_outputs(8010) <= not a;
    layer4_outputs(8011) <= not (a xor b);
    layer4_outputs(8012) <= not a;
    layer4_outputs(8013) <= not b or a;
    layer4_outputs(8014) <= a xor b;
    layer4_outputs(8015) <= a;
    layer4_outputs(8016) <= not (a or b);
    layer4_outputs(8017) <= not b or a;
    layer4_outputs(8018) <= not b;
    layer4_outputs(8019) <= not (a and b);
    layer4_outputs(8020) <= a and not b;
    layer4_outputs(8021) <= a or b;
    layer4_outputs(8022) <= a or b;
    layer4_outputs(8023) <= not (a and b);
    layer4_outputs(8024) <= a xor b;
    layer4_outputs(8025) <= not (a xor b);
    layer4_outputs(8026) <= a or b;
    layer4_outputs(8027) <= not b;
    layer4_outputs(8028) <= b;
    layer4_outputs(8029) <= not b;
    layer4_outputs(8030) <= not a;
    layer4_outputs(8031) <= not a;
    layer4_outputs(8032) <= not b or a;
    layer4_outputs(8033) <= not a;
    layer4_outputs(8034) <= not (a xor b);
    layer4_outputs(8035) <= a;
    layer4_outputs(8036) <= not a or b;
    layer4_outputs(8037) <= not (a or b);
    layer4_outputs(8038) <= not b;
    layer4_outputs(8039) <= b;
    layer4_outputs(8040) <= not b or a;
    layer4_outputs(8041) <= b;
    layer4_outputs(8042) <= not (a xor b);
    layer4_outputs(8043) <= a xor b;
    layer4_outputs(8044) <= not (a and b);
    layer4_outputs(8045) <= a;
    layer4_outputs(8046) <= a;
    layer4_outputs(8047) <= not (a xor b);
    layer4_outputs(8048) <= not a or b;
    layer4_outputs(8049) <= a and not b;
    layer4_outputs(8050) <= a xor b;
    layer4_outputs(8051) <= not a or b;
    layer4_outputs(8052) <= a xor b;
    layer4_outputs(8053) <= not b;
    layer4_outputs(8054) <= not b;
    layer4_outputs(8055) <= not a;
    layer4_outputs(8056) <= b and not a;
    layer4_outputs(8057) <= a and b;
    layer4_outputs(8058) <= a;
    layer4_outputs(8059) <= a xor b;
    layer4_outputs(8060) <= not a;
    layer4_outputs(8061) <= not b or a;
    layer4_outputs(8062) <= not a or b;
    layer4_outputs(8063) <= not (a xor b);
    layer4_outputs(8064) <= a;
    layer4_outputs(8065) <= b;
    layer4_outputs(8066) <= a or b;
    layer4_outputs(8067) <= not b or a;
    layer4_outputs(8068) <= a xor b;
    layer4_outputs(8069) <= a xor b;
    layer4_outputs(8070) <= not (a xor b);
    layer4_outputs(8071) <= not a;
    layer4_outputs(8072) <= b and not a;
    layer4_outputs(8073) <= a;
    layer4_outputs(8074) <= not (a xor b);
    layer4_outputs(8075) <= b;
    layer4_outputs(8076) <= b;
    layer4_outputs(8077) <= a and b;
    layer4_outputs(8078) <= a xor b;
    layer4_outputs(8079) <= b;
    layer4_outputs(8080) <= a xor b;
    layer4_outputs(8081) <= not a or b;
    layer4_outputs(8082) <= not a;
    layer4_outputs(8083) <= not b;
    layer4_outputs(8084) <= not b or a;
    layer4_outputs(8085) <= b and not a;
    layer4_outputs(8086) <= b;
    layer4_outputs(8087) <= not (a and b);
    layer4_outputs(8088) <= not a;
    layer4_outputs(8089) <= b;
    layer4_outputs(8090) <= not b;
    layer4_outputs(8091) <= not (a xor b);
    layer4_outputs(8092) <= not b;
    layer4_outputs(8093) <= b and not a;
    layer4_outputs(8094) <= not (a and b);
    layer4_outputs(8095) <= not a;
    layer4_outputs(8096) <= a;
    layer4_outputs(8097) <= not (a xor b);
    layer4_outputs(8098) <= not a;
    layer4_outputs(8099) <= a and b;
    layer4_outputs(8100) <= a or b;
    layer4_outputs(8101) <= not (a and b);
    layer4_outputs(8102) <= b;
    layer4_outputs(8103) <= not b;
    layer4_outputs(8104) <= not a or b;
    layer4_outputs(8105) <= a;
    layer4_outputs(8106) <= not b;
    layer4_outputs(8107) <= a and b;
    layer4_outputs(8108) <= not b or a;
    layer4_outputs(8109) <= a;
    layer4_outputs(8110) <= a and b;
    layer4_outputs(8111) <= not a;
    layer4_outputs(8112) <= a or b;
    layer4_outputs(8113) <= not b;
    layer4_outputs(8114) <= a;
    layer4_outputs(8115) <= not (a xor b);
    layer4_outputs(8116) <= a;
    layer4_outputs(8117) <= not a;
    layer4_outputs(8118) <= not (a or b);
    layer4_outputs(8119) <= a;
    layer4_outputs(8120) <= a or b;
    layer4_outputs(8121) <= not b;
    layer4_outputs(8122) <= not a;
    layer4_outputs(8123) <= a or b;
    layer4_outputs(8124) <= a xor b;
    layer4_outputs(8125) <= a xor b;
    layer4_outputs(8126) <= b;
    layer4_outputs(8127) <= b;
    layer4_outputs(8128) <= b;
    layer4_outputs(8129) <= b;
    layer4_outputs(8130) <= a and b;
    layer4_outputs(8131) <= not b or a;
    layer4_outputs(8132) <= not b;
    layer4_outputs(8133) <= not (a xor b);
    layer4_outputs(8134) <= a;
    layer4_outputs(8135) <= b and not a;
    layer4_outputs(8136) <= not (a xor b);
    layer4_outputs(8137) <= b;
    layer4_outputs(8138) <= not (a xor b);
    layer4_outputs(8139) <= not b;
    layer4_outputs(8140) <= a xor b;
    layer4_outputs(8141) <= b;
    layer4_outputs(8142) <= not (a xor b);
    layer4_outputs(8143) <= not b;
    layer4_outputs(8144) <= not a;
    layer4_outputs(8145) <= not (a xor b);
    layer4_outputs(8146) <= not b;
    layer4_outputs(8147) <= not a;
    layer4_outputs(8148) <= not b or a;
    layer4_outputs(8149) <= not a or b;
    layer4_outputs(8150) <= a or b;
    layer4_outputs(8151) <= a and b;
    layer4_outputs(8152) <= a or b;
    layer4_outputs(8153) <= b;
    layer4_outputs(8154) <= a;
    layer4_outputs(8155) <= a xor b;
    layer4_outputs(8156) <= not b;
    layer4_outputs(8157) <= not a;
    layer4_outputs(8158) <= a xor b;
    layer4_outputs(8159) <= a and not b;
    layer4_outputs(8160) <= a;
    layer4_outputs(8161) <= not a;
    layer4_outputs(8162) <= b;
    layer4_outputs(8163) <= not b;
    layer4_outputs(8164) <= a xor b;
    layer4_outputs(8165) <= a and b;
    layer4_outputs(8166) <= not b;
    layer4_outputs(8167) <= not (a and b);
    layer4_outputs(8168) <= a;
    layer4_outputs(8169) <= not a or b;
    layer4_outputs(8170) <= not (a xor b);
    layer4_outputs(8171) <= not (a or b);
    layer4_outputs(8172) <= not b;
    layer4_outputs(8173) <= not a or b;
    layer4_outputs(8174) <= b;
    layer4_outputs(8175) <= not a;
    layer4_outputs(8176) <= not (a or b);
    layer4_outputs(8177) <= a;
    layer4_outputs(8178) <= not a;
    layer4_outputs(8179) <= b;
    layer4_outputs(8180) <= b;
    layer4_outputs(8181) <= a and b;
    layer4_outputs(8182) <= a;
    layer4_outputs(8183) <= b and not a;
    layer4_outputs(8184) <= a;
    layer4_outputs(8185) <= not a or b;
    layer4_outputs(8186) <= not b;
    layer4_outputs(8187) <= a and not b;
    layer4_outputs(8188) <= a xor b;
    layer4_outputs(8189) <= not (a or b);
    layer4_outputs(8190) <= a;
    layer4_outputs(8191) <= b;
    layer4_outputs(8192) <= not a;
    layer4_outputs(8193) <= a xor b;
    layer4_outputs(8194) <= not b;
    layer4_outputs(8195) <= a and b;
    layer4_outputs(8196) <= b and not a;
    layer4_outputs(8197) <= a xor b;
    layer4_outputs(8198) <= a or b;
    layer4_outputs(8199) <= a or b;
    layer4_outputs(8200) <= b;
    layer4_outputs(8201) <= not (a xor b);
    layer4_outputs(8202) <= not (a xor b);
    layer4_outputs(8203) <= a;
    layer4_outputs(8204) <= b;
    layer4_outputs(8205) <= not a;
    layer4_outputs(8206) <= not (a and b);
    layer4_outputs(8207) <= not (a or b);
    layer4_outputs(8208) <= not a;
    layer4_outputs(8209) <= b;
    layer4_outputs(8210) <= not a or b;
    layer4_outputs(8211) <= not a;
    layer4_outputs(8212) <= a xor b;
    layer4_outputs(8213) <= not a or b;
    layer4_outputs(8214) <= not (a xor b);
    layer4_outputs(8215) <= b and not a;
    layer4_outputs(8216) <= not a or b;
    layer4_outputs(8217) <= not a or b;
    layer4_outputs(8218) <= a xor b;
    layer4_outputs(8219) <= not a;
    layer4_outputs(8220) <= not (a xor b);
    layer4_outputs(8221) <= a;
    layer4_outputs(8222) <= not b;
    layer4_outputs(8223) <= b and not a;
    layer4_outputs(8224) <= a and b;
    layer4_outputs(8225) <= not a or b;
    layer4_outputs(8226) <= not b or a;
    layer4_outputs(8227) <= not (a xor b);
    layer4_outputs(8228) <= b;
    layer4_outputs(8229) <= not b;
    layer4_outputs(8230) <= not (a and b);
    layer4_outputs(8231) <= not b;
    layer4_outputs(8232) <= not b or a;
    layer4_outputs(8233) <= not (a or b);
    layer4_outputs(8234) <= not (a xor b);
    layer4_outputs(8235) <= b;
    layer4_outputs(8236) <= not a or b;
    layer4_outputs(8237) <= not (a xor b);
    layer4_outputs(8238) <= a xor b;
    layer4_outputs(8239) <= a;
    layer4_outputs(8240) <= a;
    layer4_outputs(8241) <= not a or b;
    layer4_outputs(8242) <= not a;
    layer4_outputs(8243) <= a and b;
    layer4_outputs(8244) <= a xor b;
    layer4_outputs(8245) <= a xor b;
    layer4_outputs(8246) <= b and not a;
    layer4_outputs(8247) <= not a;
    layer4_outputs(8248) <= a;
    layer4_outputs(8249) <= not (a and b);
    layer4_outputs(8250) <= not b or a;
    layer4_outputs(8251) <= a xor b;
    layer4_outputs(8252) <= a xor b;
    layer4_outputs(8253) <= a or b;
    layer4_outputs(8254) <= a;
    layer4_outputs(8255) <= not (a and b);
    layer4_outputs(8256) <= b and not a;
    layer4_outputs(8257) <= b and not a;
    layer4_outputs(8258) <= not b;
    layer4_outputs(8259) <= a and b;
    layer4_outputs(8260) <= not (a xor b);
    layer4_outputs(8261) <= a;
    layer4_outputs(8262) <= a and not b;
    layer4_outputs(8263) <= a xor b;
    layer4_outputs(8264) <= not (a and b);
    layer4_outputs(8265) <= b;
    layer4_outputs(8266) <= a and not b;
    layer4_outputs(8267) <= not a or b;
    layer4_outputs(8268) <= a xor b;
    layer4_outputs(8269) <= not (a or b);
    layer4_outputs(8270) <= not a;
    layer4_outputs(8271) <= b;
    layer4_outputs(8272) <= not b;
    layer4_outputs(8273) <= not a;
    layer4_outputs(8274) <= a and b;
    layer4_outputs(8275) <= not a or b;
    layer4_outputs(8276) <= not b;
    layer4_outputs(8277) <= not (a xor b);
    layer4_outputs(8278) <= b;
    layer4_outputs(8279) <= a;
    layer4_outputs(8280) <= b;
    layer4_outputs(8281) <= not (a and b);
    layer4_outputs(8282) <= b;
    layer4_outputs(8283) <= not (a and b);
    layer4_outputs(8284) <= a and not b;
    layer4_outputs(8285) <= not b;
    layer4_outputs(8286) <= not (a xor b);
    layer4_outputs(8287) <= a;
    layer4_outputs(8288) <= not b or a;
    layer4_outputs(8289) <= a or b;
    layer4_outputs(8290) <= not b;
    layer4_outputs(8291) <= b and not a;
    layer4_outputs(8292) <= not b;
    layer4_outputs(8293) <= not (a xor b);
    layer4_outputs(8294) <= not a;
    layer4_outputs(8295) <= not b or a;
    layer4_outputs(8296) <= not b;
    layer4_outputs(8297) <= not (a xor b);
    layer4_outputs(8298) <= not (a or b);
    layer4_outputs(8299) <= not (a and b);
    layer4_outputs(8300) <= b;
    layer4_outputs(8301) <= not (a and b);
    layer4_outputs(8302) <= not b;
    layer4_outputs(8303) <= a or b;
    layer4_outputs(8304) <= a and not b;
    layer4_outputs(8305) <= a xor b;
    layer4_outputs(8306) <= not b;
    layer4_outputs(8307) <= not b;
    layer4_outputs(8308) <= a and not b;
    layer4_outputs(8309) <= not a;
    layer4_outputs(8310) <= not a;
    layer4_outputs(8311) <= not a;
    layer4_outputs(8312) <= a;
    layer4_outputs(8313) <= not (a xor b);
    layer4_outputs(8314) <= b and not a;
    layer4_outputs(8315) <= b;
    layer4_outputs(8316) <= a and b;
    layer4_outputs(8317) <= a or b;
    layer4_outputs(8318) <= b and not a;
    layer4_outputs(8319) <= a xor b;
    layer4_outputs(8320) <= not b;
    layer4_outputs(8321) <= b and not a;
    layer4_outputs(8322) <= not a or b;
    layer4_outputs(8323) <= not (a or b);
    layer4_outputs(8324) <= not (a and b);
    layer4_outputs(8325) <= not (a and b);
    layer4_outputs(8326) <= a;
    layer4_outputs(8327) <= not (a xor b);
    layer4_outputs(8328) <= not (a and b);
    layer4_outputs(8329) <= a;
    layer4_outputs(8330) <= a or b;
    layer4_outputs(8331) <= not (a xor b);
    layer4_outputs(8332) <= not a;
    layer4_outputs(8333) <= not b;
    layer4_outputs(8334) <= not b or a;
    layer4_outputs(8335) <= not (a or b);
    layer4_outputs(8336) <= not (a xor b);
    layer4_outputs(8337) <= not a or b;
    layer4_outputs(8338) <= not b;
    layer4_outputs(8339) <= b;
    layer4_outputs(8340) <= a xor b;
    layer4_outputs(8341) <= not a;
    layer4_outputs(8342) <= not (a xor b);
    layer4_outputs(8343) <= a or b;
    layer4_outputs(8344) <= a and b;
    layer4_outputs(8345) <= not a;
    layer4_outputs(8346) <= a;
    layer4_outputs(8347) <= a;
    layer4_outputs(8348) <= a or b;
    layer4_outputs(8349) <= a and b;
    layer4_outputs(8350) <= b;
    layer4_outputs(8351) <= not a;
    layer4_outputs(8352) <= not b or a;
    layer4_outputs(8353) <= not (a xor b);
    layer4_outputs(8354) <= a;
    layer4_outputs(8355) <= b;
    layer4_outputs(8356) <= a;
    layer4_outputs(8357) <= b;
    layer4_outputs(8358) <= not (a or b);
    layer4_outputs(8359) <= a;
    layer4_outputs(8360) <= not a;
    layer4_outputs(8361) <= not b;
    layer4_outputs(8362) <= a and not b;
    layer4_outputs(8363) <= a;
    layer4_outputs(8364) <= a or b;
    layer4_outputs(8365) <= not b;
    layer4_outputs(8366) <= a;
    layer4_outputs(8367) <= a and b;
    layer4_outputs(8368) <= b;
    layer4_outputs(8369) <= not a;
    layer4_outputs(8370) <= not b;
    layer4_outputs(8371) <= not (a xor b);
    layer4_outputs(8372) <= not b;
    layer4_outputs(8373) <= not b;
    layer4_outputs(8374) <= b;
    layer4_outputs(8375) <= a;
    layer4_outputs(8376) <= not b;
    layer4_outputs(8377) <= a;
    layer4_outputs(8378) <= a or b;
    layer4_outputs(8379) <= not a;
    layer4_outputs(8380) <= not (a or b);
    layer4_outputs(8381) <= not a or b;
    layer4_outputs(8382) <= not a;
    layer4_outputs(8383) <= not a;
    layer4_outputs(8384) <= a xor b;
    layer4_outputs(8385) <= not b;
    layer4_outputs(8386) <= a and not b;
    layer4_outputs(8387) <= not a;
    layer4_outputs(8388) <= not (a or b);
    layer4_outputs(8389) <= not b;
    layer4_outputs(8390) <= a and b;
    layer4_outputs(8391) <= a and b;
    layer4_outputs(8392) <= a or b;
    layer4_outputs(8393) <= a;
    layer4_outputs(8394) <= not a;
    layer4_outputs(8395) <= not a;
    layer4_outputs(8396) <= a;
    layer4_outputs(8397) <= a xor b;
    layer4_outputs(8398) <= not a;
    layer4_outputs(8399) <= a or b;
    layer4_outputs(8400) <= not (a xor b);
    layer4_outputs(8401) <= not (a or b);
    layer4_outputs(8402) <= b and not a;
    layer4_outputs(8403) <= a xor b;
    layer4_outputs(8404) <= a and b;
    layer4_outputs(8405) <= not b;
    layer4_outputs(8406) <= b;
    layer4_outputs(8407) <= not b;
    layer4_outputs(8408) <= b;
    layer4_outputs(8409) <= not b or a;
    layer4_outputs(8410) <= not b;
    layer4_outputs(8411) <= b;
    layer4_outputs(8412) <= a and not b;
    layer4_outputs(8413) <= not b;
    layer4_outputs(8414) <= a;
    layer4_outputs(8415) <= not a;
    layer4_outputs(8416) <= not a or b;
    layer4_outputs(8417) <= not b or a;
    layer4_outputs(8418) <= not a;
    layer4_outputs(8419) <= a;
    layer4_outputs(8420) <= not (a xor b);
    layer4_outputs(8421) <= not b;
    layer4_outputs(8422) <= not b;
    layer4_outputs(8423) <= b;
    layer4_outputs(8424) <= b;
    layer4_outputs(8425) <= not (a and b);
    layer4_outputs(8426) <= not (a or b);
    layer4_outputs(8427) <= b;
    layer4_outputs(8428) <= not (a or b);
    layer4_outputs(8429) <= a or b;
    layer4_outputs(8430) <= b;
    layer4_outputs(8431) <= not a or b;
    layer4_outputs(8432) <= not b;
    layer4_outputs(8433) <= a and b;
    layer4_outputs(8434) <= a and b;
    layer4_outputs(8435) <= not b or a;
    layer4_outputs(8436) <= not (a or b);
    layer4_outputs(8437) <= a xor b;
    layer4_outputs(8438) <= not a;
    layer4_outputs(8439) <= not a;
    layer4_outputs(8440) <= a and b;
    layer4_outputs(8441) <= a xor b;
    layer4_outputs(8442) <= not a;
    layer4_outputs(8443) <= not (a or b);
    layer4_outputs(8444) <= b;
    layer4_outputs(8445) <= a xor b;
    layer4_outputs(8446) <= a or b;
    layer4_outputs(8447) <= not (a or b);
    layer4_outputs(8448) <= not b;
    layer4_outputs(8449) <= a and b;
    layer4_outputs(8450) <= b;
    layer4_outputs(8451) <= not (a or b);
    layer4_outputs(8452) <= not (a xor b);
    layer4_outputs(8453) <= not (a or b);
    layer4_outputs(8454) <= not a or b;
    layer4_outputs(8455) <= not a;
    layer4_outputs(8456) <= 1'b0;
    layer4_outputs(8457) <= not (a xor b);
    layer4_outputs(8458) <= not (a or b);
    layer4_outputs(8459) <= not (a xor b);
    layer4_outputs(8460) <= b;
    layer4_outputs(8461) <= not (a xor b);
    layer4_outputs(8462) <= not a;
    layer4_outputs(8463) <= a and b;
    layer4_outputs(8464) <= a and b;
    layer4_outputs(8465) <= b and not a;
    layer4_outputs(8466) <= not b or a;
    layer4_outputs(8467) <= not b;
    layer4_outputs(8468) <= not (a xor b);
    layer4_outputs(8469) <= b;
    layer4_outputs(8470) <= a xor b;
    layer4_outputs(8471) <= a xor b;
    layer4_outputs(8472) <= not b or a;
    layer4_outputs(8473) <= a and b;
    layer4_outputs(8474) <= b;
    layer4_outputs(8475) <= b;
    layer4_outputs(8476) <= not a;
    layer4_outputs(8477) <= a;
    layer4_outputs(8478) <= not a;
    layer4_outputs(8479) <= b;
    layer4_outputs(8480) <= b;
    layer4_outputs(8481) <= a xor b;
    layer4_outputs(8482) <= not a or b;
    layer4_outputs(8483) <= a or b;
    layer4_outputs(8484) <= not (a xor b);
    layer4_outputs(8485) <= a;
    layer4_outputs(8486) <= not a;
    layer4_outputs(8487) <= b;
    layer4_outputs(8488) <= b;
    layer4_outputs(8489) <= a xor b;
    layer4_outputs(8490) <= not (a xor b);
    layer4_outputs(8491) <= not b;
    layer4_outputs(8492) <= not b;
    layer4_outputs(8493) <= b and not a;
    layer4_outputs(8494) <= not (a xor b);
    layer4_outputs(8495) <= a xor b;
    layer4_outputs(8496) <= a xor b;
    layer4_outputs(8497) <= not a;
    layer4_outputs(8498) <= a xor b;
    layer4_outputs(8499) <= not b;
    layer4_outputs(8500) <= not (a and b);
    layer4_outputs(8501) <= a;
    layer4_outputs(8502) <= a xor b;
    layer4_outputs(8503) <= not a;
    layer4_outputs(8504) <= a xor b;
    layer4_outputs(8505) <= not (a and b);
    layer4_outputs(8506) <= b;
    layer4_outputs(8507) <= 1'b1;
    layer4_outputs(8508) <= a;
    layer4_outputs(8509) <= not a;
    layer4_outputs(8510) <= a xor b;
    layer4_outputs(8511) <= not a or b;
    layer4_outputs(8512) <= not (a and b);
    layer4_outputs(8513) <= not (a xor b);
    layer4_outputs(8514) <= a xor b;
    layer4_outputs(8515) <= not b;
    layer4_outputs(8516) <= not b;
    layer4_outputs(8517) <= not b;
    layer4_outputs(8518) <= a xor b;
    layer4_outputs(8519) <= not b;
    layer4_outputs(8520) <= not b;
    layer4_outputs(8521) <= a;
    layer4_outputs(8522) <= 1'b1;
    layer4_outputs(8523) <= not (a xor b);
    layer4_outputs(8524) <= not b or a;
    layer4_outputs(8525) <= not b;
    layer4_outputs(8526) <= not (a and b);
    layer4_outputs(8527) <= not a;
    layer4_outputs(8528) <= not b;
    layer4_outputs(8529) <= a;
    layer4_outputs(8530) <= not b or a;
    layer4_outputs(8531) <= a xor b;
    layer4_outputs(8532) <= not b;
    layer4_outputs(8533) <= a or b;
    layer4_outputs(8534) <= a and b;
    layer4_outputs(8535) <= a;
    layer4_outputs(8536) <= b;
    layer4_outputs(8537) <= not a or b;
    layer4_outputs(8538) <= not b;
    layer4_outputs(8539) <= not (a xor b);
    layer4_outputs(8540) <= a;
    layer4_outputs(8541) <= not a;
    layer4_outputs(8542) <= not (a xor b);
    layer4_outputs(8543) <= a xor b;
    layer4_outputs(8544) <= not b or a;
    layer4_outputs(8545) <= b and not a;
    layer4_outputs(8546) <= not (a or b);
    layer4_outputs(8547) <= not b or a;
    layer4_outputs(8548) <= a;
    layer4_outputs(8549) <= not b or a;
    layer4_outputs(8550) <= not b;
    layer4_outputs(8551) <= a;
    layer4_outputs(8552) <= a and b;
    layer4_outputs(8553) <= a;
    layer4_outputs(8554) <= not b;
    layer4_outputs(8555) <= a or b;
    layer4_outputs(8556) <= b and not a;
    layer4_outputs(8557) <= b;
    layer4_outputs(8558) <= not b;
    layer4_outputs(8559) <= a or b;
    layer4_outputs(8560) <= not (a xor b);
    layer4_outputs(8561) <= b and not a;
    layer4_outputs(8562) <= not (a xor b);
    layer4_outputs(8563) <= not (a xor b);
    layer4_outputs(8564) <= a xor b;
    layer4_outputs(8565) <= a and not b;
    layer4_outputs(8566) <= not a or b;
    layer4_outputs(8567) <= not b;
    layer4_outputs(8568) <= a;
    layer4_outputs(8569) <= not b;
    layer4_outputs(8570) <= not b;
    layer4_outputs(8571) <= not a or b;
    layer4_outputs(8572) <= not b;
    layer4_outputs(8573) <= a xor b;
    layer4_outputs(8574) <= a or b;
    layer4_outputs(8575) <= not a;
    layer4_outputs(8576) <= b;
    layer4_outputs(8577) <= not b;
    layer4_outputs(8578) <= a xor b;
    layer4_outputs(8579) <= not (a or b);
    layer4_outputs(8580) <= not a;
    layer4_outputs(8581) <= not (a xor b);
    layer4_outputs(8582) <= not b or a;
    layer4_outputs(8583) <= a or b;
    layer4_outputs(8584) <= not (a xor b);
    layer4_outputs(8585) <= not (a xor b);
    layer4_outputs(8586) <= 1'b1;
    layer4_outputs(8587) <= not (a xor b);
    layer4_outputs(8588) <= not b;
    layer4_outputs(8589) <= a and b;
    layer4_outputs(8590) <= not (a xor b);
    layer4_outputs(8591) <= not (a xor b);
    layer4_outputs(8592) <= not a;
    layer4_outputs(8593) <= not a;
    layer4_outputs(8594) <= not b;
    layer4_outputs(8595) <= a;
    layer4_outputs(8596) <= b;
    layer4_outputs(8597) <= not (a xor b);
    layer4_outputs(8598) <= a and b;
    layer4_outputs(8599) <= a and not b;
    layer4_outputs(8600) <= b and not a;
    layer4_outputs(8601) <= a and b;
    layer4_outputs(8602) <= not (a and b);
    layer4_outputs(8603) <= a xor b;
    layer4_outputs(8604) <= a;
    layer4_outputs(8605) <= not a or b;
    layer4_outputs(8606) <= not b or a;
    layer4_outputs(8607) <= a;
    layer4_outputs(8608) <= b;
    layer4_outputs(8609) <= not a;
    layer4_outputs(8610) <= not b;
    layer4_outputs(8611) <= not b;
    layer4_outputs(8612) <= a or b;
    layer4_outputs(8613) <= not (a xor b);
    layer4_outputs(8614) <= not a;
    layer4_outputs(8615) <= a or b;
    layer4_outputs(8616) <= not a;
    layer4_outputs(8617) <= a and b;
    layer4_outputs(8618) <= a and b;
    layer4_outputs(8619) <= not b or a;
    layer4_outputs(8620) <= not a;
    layer4_outputs(8621) <= not a;
    layer4_outputs(8622) <= a;
    layer4_outputs(8623) <= not (a and b);
    layer4_outputs(8624) <= a;
    layer4_outputs(8625) <= b;
    layer4_outputs(8626) <= not (a xor b);
    layer4_outputs(8627) <= not b or a;
    layer4_outputs(8628) <= not a;
    layer4_outputs(8629) <= not b;
    layer4_outputs(8630) <= a;
    layer4_outputs(8631) <= a;
    layer4_outputs(8632) <= a;
    layer4_outputs(8633) <= not b;
    layer4_outputs(8634) <= not a;
    layer4_outputs(8635) <= b and not a;
    layer4_outputs(8636) <= a;
    layer4_outputs(8637) <= a;
    layer4_outputs(8638) <= b and not a;
    layer4_outputs(8639) <= a and b;
    layer4_outputs(8640) <= a or b;
    layer4_outputs(8641) <= not b or a;
    layer4_outputs(8642) <= b;
    layer4_outputs(8643) <= a xor b;
    layer4_outputs(8644) <= not a;
    layer4_outputs(8645) <= a;
    layer4_outputs(8646) <= not b;
    layer4_outputs(8647) <= a;
    layer4_outputs(8648) <= not b;
    layer4_outputs(8649) <= b;
    layer4_outputs(8650) <= not a;
    layer4_outputs(8651) <= not a or b;
    layer4_outputs(8652) <= a and b;
    layer4_outputs(8653) <= not (a xor b);
    layer4_outputs(8654) <= not (a xor b);
    layer4_outputs(8655) <= a;
    layer4_outputs(8656) <= a xor b;
    layer4_outputs(8657) <= a;
    layer4_outputs(8658) <= not (a xor b);
    layer4_outputs(8659) <= a or b;
    layer4_outputs(8660) <= b;
    layer4_outputs(8661) <= not a;
    layer4_outputs(8662) <= a and not b;
    layer4_outputs(8663) <= not b or a;
    layer4_outputs(8664) <= b;
    layer4_outputs(8665) <= not a;
    layer4_outputs(8666) <= not a;
    layer4_outputs(8667) <= not b;
    layer4_outputs(8668) <= a and not b;
    layer4_outputs(8669) <= a and b;
    layer4_outputs(8670) <= not (a and b);
    layer4_outputs(8671) <= a xor b;
    layer4_outputs(8672) <= not (a and b);
    layer4_outputs(8673) <= a;
    layer4_outputs(8674) <= a;
    layer4_outputs(8675) <= not b;
    layer4_outputs(8676) <= a or b;
    layer4_outputs(8677) <= a;
    layer4_outputs(8678) <= not a;
    layer4_outputs(8679) <= not a;
    layer4_outputs(8680) <= not (a xor b);
    layer4_outputs(8681) <= not a or b;
    layer4_outputs(8682) <= b;
    layer4_outputs(8683) <= not a;
    layer4_outputs(8684) <= not (a xor b);
    layer4_outputs(8685) <= not (a and b);
    layer4_outputs(8686) <= not b;
    layer4_outputs(8687) <= b;
    layer4_outputs(8688) <= a and not b;
    layer4_outputs(8689) <= not a or b;
    layer4_outputs(8690) <= a;
    layer4_outputs(8691) <= b;
    layer4_outputs(8692) <= not a;
    layer4_outputs(8693) <= a and not b;
    layer4_outputs(8694) <= not b;
    layer4_outputs(8695) <= b;
    layer4_outputs(8696) <= not a;
    layer4_outputs(8697) <= not (a and b);
    layer4_outputs(8698) <= not (a and b);
    layer4_outputs(8699) <= a and not b;
    layer4_outputs(8700) <= not b;
    layer4_outputs(8701) <= not b;
    layer4_outputs(8702) <= a and b;
    layer4_outputs(8703) <= b;
    layer4_outputs(8704) <= a;
    layer4_outputs(8705) <= not a;
    layer4_outputs(8706) <= b;
    layer4_outputs(8707) <= a xor b;
    layer4_outputs(8708) <= not (a and b);
    layer4_outputs(8709) <= b;
    layer4_outputs(8710) <= b;
    layer4_outputs(8711) <= not (a and b);
    layer4_outputs(8712) <= a and not b;
    layer4_outputs(8713) <= b;
    layer4_outputs(8714) <= not b;
    layer4_outputs(8715) <= a and b;
    layer4_outputs(8716) <= b;
    layer4_outputs(8717) <= a xor b;
    layer4_outputs(8718) <= not (a xor b);
    layer4_outputs(8719) <= a xor b;
    layer4_outputs(8720) <= a xor b;
    layer4_outputs(8721) <= not (a or b);
    layer4_outputs(8722) <= not a or b;
    layer4_outputs(8723) <= not a;
    layer4_outputs(8724) <= a;
    layer4_outputs(8725) <= not a;
    layer4_outputs(8726) <= not b;
    layer4_outputs(8727) <= not a or b;
    layer4_outputs(8728) <= not a;
    layer4_outputs(8729) <= b;
    layer4_outputs(8730) <= b and not a;
    layer4_outputs(8731) <= a or b;
    layer4_outputs(8732) <= b;
    layer4_outputs(8733) <= not (a and b);
    layer4_outputs(8734) <= not b or a;
    layer4_outputs(8735) <= a xor b;
    layer4_outputs(8736) <= not (a xor b);
    layer4_outputs(8737) <= a and not b;
    layer4_outputs(8738) <= a and not b;
    layer4_outputs(8739) <= a;
    layer4_outputs(8740) <= a and b;
    layer4_outputs(8741) <= a or b;
    layer4_outputs(8742) <= a and b;
    layer4_outputs(8743) <= not (a and b);
    layer4_outputs(8744) <= not (a xor b);
    layer4_outputs(8745) <= not (a xor b);
    layer4_outputs(8746) <= not b or a;
    layer4_outputs(8747) <= not b;
    layer4_outputs(8748) <= not (a or b);
    layer4_outputs(8749) <= b;
    layer4_outputs(8750) <= not (a xor b);
    layer4_outputs(8751) <= a and b;
    layer4_outputs(8752) <= b;
    layer4_outputs(8753) <= not b;
    layer4_outputs(8754) <= not (a or b);
    layer4_outputs(8755) <= b and not a;
    layer4_outputs(8756) <= b;
    layer4_outputs(8757) <= b;
    layer4_outputs(8758) <= not (a and b);
    layer4_outputs(8759) <= not a or b;
    layer4_outputs(8760) <= not (a xor b);
    layer4_outputs(8761) <= a or b;
    layer4_outputs(8762) <= a;
    layer4_outputs(8763) <= not (a xor b);
    layer4_outputs(8764) <= a and not b;
    layer4_outputs(8765) <= not (a or b);
    layer4_outputs(8766) <= a;
    layer4_outputs(8767) <= a or b;
    layer4_outputs(8768) <= not (a and b);
    layer4_outputs(8769) <= a xor b;
    layer4_outputs(8770) <= b;
    layer4_outputs(8771) <= not a;
    layer4_outputs(8772) <= not (a or b);
    layer4_outputs(8773) <= a and b;
    layer4_outputs(8774) <= not b;
    layer4_outputs(8775) <= a and b;
    layer4_outputs(8776) <= not b;
    layer4_outputs(8777) <= a and not b;
    layer4_outputs(8778) <= a and b;
    layer4_outputs(8779) <= not (a or b);
    layer4_outputs(8780) <= a and b;
    layer4_outputs(8781) <= a;
    layer4_outputs(8782) <= not b;
    layer4_outputs(8783) <= a;
    layer4_outputs(8784) <= not (a xor b);
    layer4_outputs(8785) <= not b or a;
    layer4_outputs(8786) <= b;
    layer4_outputs(8787) <= a xor b;
    layer4_outputs(8788) <= a;
    layer4_outputs(8789) <= not a or b;
    layer4_outputs(8790) <= a;
    layer4_outputs(8791) <= a and b;
    layer4_outputs(8792) <= not (a xor b);
    layer4_outputs(8793) <= not a;
    layer4_outputs(8794) <= not b;
    layer4_outputs(8795) <= not (a or b);
    layer4_outputs(8796) <= a xor b;
    layer4_outputs(8797) <= not (a and b);
    layer4_outputs(8798) <= not b or a;
    layer4_outputs(8799) <= a;
    layer4_outputs(8800) <= a;
    layer4_outputs(8801) <= b;
    layer4_outputs(8802) <= not b or a;
    layer4_outputs(8803) <= a and not b;
    layer4_outputs(8804) <= a xor b;
    layer4_outputs(8805) <= b;
    layer4_outputs(8806) <= b;
    layer4_outputs(8807) <= not (a xor b);
    layer4_outputs(8808) <= a xor b;
    layer4_outputs(8809) <= a;
    layer4_outputs(8810) <= a;
    layer4_outputs(8811) <= a and b;
    layer4_outputs(8812) <= b;
    layer4_outputs(8813) <= not (a xor b);
    layer4_outputs(8814) <= not b;
    layer4_outputs(8815) <= not a or b;
    layer4_outputs(8816) <= not (a xor b);
    layer4_outputs(8817) <= not a;
    layer4_outputs(8818) <= a or b;
    layer4_outputs(8819) <= a xor b;
    layer4_outputs(8820) <= a and not b;
    layer4_outputs(8821) <= not (a xor b);
    layer4_outputs(8822) <= not b;
    layer4_outputs(8823) <= not b;
    layer4_outputs(8824) <= a;
    layer4_outputs(8825) <= not (a xor b);
    layer4_outputs(8826) <= a xor b;
    layer4_outputs(8827) <= not b;
    layer4_outputs(8828) <= a;
    layer4_outputs(8829) <= a;
    layer4_outputs(8830) <= a or b;
    layer4_outputs(8831) <= not (a and b);
    layer4_outputs(8832) <= a;
    layer4_outputs(8833) <= a;
    layer4_outputs(8834) <= a;
    layer4_outputs(8835) <= not (a and b);
    layer4_outputs(8836) <= a and b;
    layer4_outputs(8837) <= a;
    layer4_outputs(8838) <= b;
    layer4_outputs(8839) <= not (a xor b);
    layer4_outputs(8840) <= a and b;
    layer4_outputs(8841) <= not (a and b);
    layer4_outputs(8842) <= b;
    layer4_outputs(8843) <= not b;
    layer4_outputs(8844) <= a;
    layer4_outputs(8845) <= not (a and b);
    layer4_outputs(8846) <= not (a xor b);
    layer4_outputs(8847) <= a;
    layer4_outputs(8848) <= not a or b;
    layer4_outputs(8849) <= not b or a;
    layer4_outputs(8850) <= not b;
    layer4_outputs(8851) <= not (a xor b);
    layer4_outputs(8852) <= not b;
    layer4_outputs(8853) <= a xor b;
    layer4_outputs(8854) <= not (a or b);
    layer4_outputs(8855) <= not b;
    layer4_outputs(8856) <= a xor b;
    layer4_outputs(8857) <= b and not a;
    layer4_outputs(8858) <= not b;
    layer4_outputs(8859) <= b;
    layer4_outputs(8860) <= not (a xor b);
    layer4_outputs(8861) <= not a;
    layer4_outputs(8862) <= not (a xor b);
    layer4_outputs(8863) <= b;
    layer4_outputs(8864) <= not (a xor b);
    layer4_outputs(8865) <= not (a or b);
    layer4_outputs(8866) <= a;
    layer4_outputs(8867) <= not b;
    layer4_outputs(8868) <= not a;
    layer4_outputs(8869) <= not a;
    layer4_outputs(8870) <= not a;
    layer4_outputs(8871) <= not a;
    layer4_outputs(8872) <= a;
    layer4_outputs(8873) <= not (a xor b);
    layer4_outputs(8874) <= not b;
    layer4_outputs(8875) <= not b or a;
    layer4_outputs(8876) <= a;
    layer4_outputs(8877) <= b;
    layer4_outputs(8878) <= b;
    layer4_outputs(8879) <= b and not a;
    layer4_outputs(8880) <= a;
    layer4_outputs(8881) <= not b or a;
    layer4_outputs(8882) <= a;
    layer4_outputs(8883) <= a;
    layer4_outputs(8884) <= b and not a;
    layer4_outputs(8885) <= a or b;
    layer4_outputs(8886) <= a xor b;
    layer4_outputs(8887) <= not a;
    layer4_outputs(8888) <= a and b;
    layer4_outputs(8889) <= a;
    layer4_outputs(8890) <= not a or b;
    layer4_outputs(8891) <= not a or b;
    layer4_outputs(8892) <= not a;
    layer4_outputs(8893) <= not b;
    layer4_outputs(8894) <= b;
    layer4_outputs(8895) <= not a;
    layer4_outputs(8896) <= a xor b;
    layer4_outputs(8897) <= a and not b;
    layer4_outputs(8898) <= b;
    layer4_outputs(8899) <= a xor b;
    layer4_outputs(8900) <= not b;
    layer4_outputs(8901) <= not b;
    layer4_outputs(8902) <= not (a xor b);
    layer4_outputs(8903) <= a;
    layer4_outputs(8904) <= not (a xor b);
    layer4_outputs(8905) <= a xor b;
    layer4_outputs(8906) <= not a;
    layer4_outputs(8907) <= b;
    layer4_outputs(8908) <= not (a or b);
    layer4_outputs(8909) <= a;
    layer4_outputs(8910) <= not a;
    layer4_outputs(8911) <= b and not a;
    layer4_outputs(8912) <= not b or a;
    layer4_outputs(8913) <= not (a xor b);
    layer4_outputs(8914) <= not a;
    layer4_outputs(8915) <= a and not b;
    layer4_outputs(8916) <= a or b;
    layer4_outputs(8917) <= not b or a;
    layer4_outputs(8918) <= not a;
    layer4_outputs(8919) <= a and not b;
    layer4_outputs(8920) <= a;
    layer4_outputs(8921) <= not a;
    layer4_outputs(8922) <= b;
    layer4_outputs(8923) <= b;
    layer4_outputs(8924) <= a;
    layer4_outputs(8925) <= a;
    layer4_outputs(8926) <= b and not a;
    layer4_outputs(8927) <= not a;
    layer4_outputs(8928) <= b;
    layer4_outputs(8929) <= a xor b;
    layer4_outputs(8930) <= b;
    layer4_outputs(8931) <= a;
    layer4_outputs(8932) <= b;
    layer4_outputs(8933) <= not a;
    layer4_outputs(8934) <= not a;
    layer4_outputs(8935) <= not (a and b);
    layer4_outputs(8936) <= not a or b;
    layer4_outputs(8937) <= b;
    layer4_outputs(8938) <= b;
    layer4_outputs(8939) <= not (a or b);
    layer4_outputs(8940) <= not a;
    layer4_outputs(8941) <= not (a and b);
    layer4_outputs(8942) <= not a;
    layer4_outputs(8943) <= not a;
    layer4_outputs(8944) <= a or b;
    layer4_outputs(8945) <= b and not a;
    layer4_outputs(8946) <= not b;
    layer4_outputs(8947) <= a xor b;
    layer4_outputs(8948) <= not b;
    layer4_outputs(8949) <= not a;
    layer4_outputs(8950) <= a and b;
    layer4_outputs(8951) <= not (a or b);
    layer4_outputs(8952) <= not a;
    layer4_outputs(8953) <= a;
    layer4_outputs(8954) <= b;
    layer4_outputs(8955) <= a xor b;
    layer4_outputs(8956) <= b;
    layer4_outputs(8957) <= b;
    layer4_outputs(8958) <= not (a and b);
    layer4_outputs(8959) <= 1'b0;
    layer4_outputs(8960) <= not a;
    layer4_outputs(8961) <= not a;
    layer4_outputs(8962) <= b;
    layer4_outputs(8963) <= not b;
    layer4_outputs(8964) <= b and not a;
    layer4_outputs(8965) <= b;
    layer4_outputs(8966) <= a xor b;
    layer4_outputs(8967) <= not a or b;
    layer4_outputs(8968) <= not (a xor b);
    layer4_outputs(8969) <= a;
    layer4_outputs(8970) <= not a or b;
    layer4_outputs(8971) <= a;
    layer4_outputs(8972) <= not b;
    layer4_outputs(8973) <= a xor b;
    layer4_outputs(8974) <= a or b;
    layer4_outputs(8975) <= a or b;
    layer4_outputs(8976) <= not a;
    layer4_outputs(8977) <= a and b;
    layer4_outputs(8978) <= a and not b;
    layer4_outputs(8979) <= a;
    layer4_outputs(8980) <= a xor b;
    layer4_outputs(8981) <= not (a or b);
    layer4_outputs(8982) <= a;
    layer4_outputs(8983) <= not a;
    layer4_outputs(8984) <= a or b;
    layer4_outputs(8985) <= b and not a;
    layer4_outputs(8986) <= not (a or b);
    layer4_outputs(8987) <= not (a xor b);
    layer4_outputs(8988) <= not (a xor b);
    layer4_outputs(8989) <= b;
    layer4_outputs(8990) <= a;
    layer4_outputs(8991) <= a xor b;
    layer4_outputs(8992) <= not b;
    layer4_outputs(8993) <= b and not a;
    layer4_outputs(8994) <= b and not a;
    layer4_outputs(8995) <= b and not a;
    layer4_outputs(8996) <= b;
    layer4_outputs(8997) <= not b or a;
    layer4_outputs(8998) <= not b;
    layer4_outputs(8999) <= not a;
    layer4_outputs(9000) <= a and not b;
    layer4_outputs(9001) <= a or b;
    layer4_outputs(9002) <= not a;
    layer4_outputs(9003) <= not a;
    layer4_outputs(9004) <= not b or a;
    layer4_outputs(9005) <= a;
    layer4_outputs(9006) <= not a;
    layer4_outputs(9007) <= a and not b;
    layer4_outputs(9008) <= not b;
    layer4_outputs(9009) <= not a;
    layer4_outputs(9010) <= not (a or b);
    layer4_outputs(9011) <= not (a and b);
    layer4_outputs(9012) <= not (a xor b);
    layer4_outputs(9013) <= a or b;
    layer4_outputs(9014) <= b and not a;
    layer4_outputs(9015) <= not a;
    layer4_outputs(9016) <= not a;
    layer4_outputs(9017) <= b;
    layer4_outputs(9018) <= a;
    layer4_outputs(9019) <= a and b;
    layer4_outputs(9020) <= not (a xor b);
    layer4_outputs(9021) <= a xor b;
    layer4_outputs(9022) <= b;
    layer4_outputs(9023) <= b and not a;
    layer4_outputs(9024) <= a;
    layer4_outputs(9025) <= a xor b;
    layer4_outputs(9026) <= not b;
    layer4_outputs(9027) <= a and b;
    layer4_outputs(9028) <= a and not b;
    layer4_outputs(9029) <= b;
    layer4_outputs(9030) <= not a or b;
    layer4_outputs(9031) <= a or b;
    layer4_outputs(9032) <= not (a xor b);
    layer4_outputs(9033) <= b;
    layer4_outputs(9034) <= not a or b;
    layer4_outputs(9035) <= not a;
    layer4_outputs(9036) <= not b or a;
    layer4_outputs(9037) <= a;
    layer4_outputs(9038) <= b;
    layer4_outputs(9039) <= not a or b;
    layer4_outputs(9040) <= b;
    layer4_outputs(9041) <= a;
    layer4_outputs(9042) <= b and not a;
    layer4_outputs(9043) <= a and b;
    layer4_outputs(9044) <= not b or a;
    layer4_outputs(9045) <= b and not a;
    layer4_outputs(9046) <= not a;
    layer4_outputs(9047) <= not a;
    layer4_outputs(9048) <= a xor b;
    layer4_outputs(9049) <= not b;
    layer4_outputs(9050) <= b and not a;
    layer4_outputs(9051) <= b and not a;
    layer4_outputs(9052) <= not (a or b);
    layer4_outputs(9053) <= not b;
    layer4_outputs(9054) <= not a;
    layer4_outputs(9055) <= not (a and b);
    layer4_outputs(9056) <= not (a and b);
    layer4_outputs(9057) <= not a;
    layer4_outputs(9058) <= b and not a;
    layer4_outputs(9059) <= not b or a;
    layer4_outputs(9060) <= b and not a;
    layer4_outputs(9061) <= not a;
    layer4_outputs(9062) <= not b;
    layer4_outputs(9063) <= not a or b;
    layer4_outputs(9064) <= not a;
    layer4_outputs(9065) <= b;
    layer4_outputs(9066) <= a;
    layer4_outputs(9067) <= not (a or b);
    layer4_outputs(9068) <= a and not b;
    layer4_outputs(9069) <= 1'b0;
    layer4_outputs(9070) <= a;
    layer4_outputs(9071) <= not b;
    layer4_outputs(9072) <= not a;
    layer4_outputs(9073) <= b;
    layer4_outputs(9074) <= a xor b;
    layer4_outputs(9075) <= a and b;
    layer4_outputs(9076) <= not b;
    layer4_outputs(9077) <= b;
    layer4_outputs(9078) <= a xor b;
    layer4_outputs(9079) <= not b or a;
    layer4_outputs(9080) <= a;
    layer4_outputs(9081) <= a and b;
    layer4_outputs(9082) <= a;
    layer4_outputs(9083) <= a or b;
    layer4_outputs(9084) <= a;
    layer4_outputs(9085) <= a xor b;
    layer4_outputs(9086) <= not b or a;
    layer4_outputs(9087) <= a xor b;
    layer4_outputs(9088) <= not b;
    layer4_outputs(9089) <= b;
    layer4_outputs(9090) <= not a or b;
    layer4_outputs(9091) <= not (a or b);
    layer4_outputs(9092) <= not b or a;
    layer4_outputs(9093) <= not (a xor b);
    layer4_outputs(9094) <= not (a or b);
    layer4_outputs(9095) <= b;
    layer4_outputs(9096) <= not (a and b);
    layer4_outputs(9097) <= not a or b;
    layer4_outputs(9098) <= not a;
    layer4_outputs(9099) <= not b;
    layer4_outputs(9100) <= b;
    layer4_outputs(9101) <= a;
    layer4_outputs(9102) <= not b;
    layer4_outputs(9103) <= not (a xor b);
    layer4_outputs(9104) <= a;
    layer4_outputs(9105) <= not b;
    layer4_outputs(9106) <= a;
    layer4_outputs(9107) <= a and not b;
    layer4_outputs(9108) <= not a;
    layer4_outputs(9109) <= not (a or b);
    layer4_outputs(9110) <= b and not a;
    layer4_outputs(9111) <= b;
    layer4_outputs(9112) <= not b;
    layer4_outputs(9113) <= not (a xor b);
    layer4_outputs(9114) <= b;
    layer4_outputs(9115) <= not (a or b);
    layer4_outputs(9116) <= a xor b;
    layer4_outputs(9117) <= a and not b;
    layer4_outputs(9118) <= not (a xor b);
    layer4_outputs(9119) <= a and not b;
    layer4_outputs(9120) <= not (a and b);
    layer4_outputs(9121) <= not (a xor b);
    layer4_outputs(9122) <= not (a xor b);
    layer4_outputs(9123) <= b;
    layer4_outputs(9124) <= not a or b;
    layer4_outputs(9125) <= a xor b;
    layer4_outputs(9126) <= not a or b;
    layer4_outputs(9127) <= not a;
    layer4_outputs(9128) <= a;
    layer4_outputs(9129) <= not b;
    layer4_outputs(9130) <= not b;
    layer4_outputs(9131) <= a or b;
    layer4_outputs(9132) <= b;
    layer4_outputs(9133) <= not a;
    layer4_outputs(9134) <= not (a xor b);
    layer4_outputs(9135) <= b and not a;
    layer4_outputs(9136) <= a;
    layer4_outputs(9137) <= not (a xor b);
    layer4_outputs(9138) <= a xor b;
    layer4_outputs(9139) <= b;
    layer4_outputs(9140) <= a xor b;
    layer4_outputs(9141) <= a xor b;
    layer4_outputs(9142) <= not a;
    layer4_outputs(9143) <= a xor b;
    layer4_outputs(9144) <= not b;
    layer4_outputs(9145) <= not a;
    layer4_outputs(9146) <= a;
    layer4_outputs(9147) <= not (a and b);
    layer4_outputs(9148) <= b and not a;
    layer4_outputs(9149) <= a and b;
    layer4_outputs(9150) <= b;
    layer4_outputs(9151) <= a and not b;
    layer4_outputs(9152) <= a or b;
    layer4_outputs(9153) <= b;
    layer4_outputs(9154) <= a;
    layer4_outputs(9155) <= not (a or b);
    layer4_outputs(9156) <= b;
    layer4_outputs(9157) <= not b;
    layer4_outputs(9158) <= not a;
    layer4_outputs(9159) <= a and not b;
    layer4_outputs(9160) <= not (a and b);
    layer4_outputs(9161) <= a and not b;
    layer4_outputs(9162) <= a xor b;
    layer4_outputs(9163) <= 1'b0;
    layer4_outputs(9164) <= not b or a;
    layer4_outputs(9165) <= b and not a;
    layer4_outputs(9166) <= not a;
    layer4_outputs(9167) <= a and not b;
    layer4_outputs(9168) <= not b;
    layer4_outputs(9169) <= b;
    layer4_outputs(9170) <= not (a xor b);
    layer4_outputs(9171) <= not a;
    layer4_outputs(9172) <= not (a xor b);
    layer4_outputs(9173) <= a or b;
    layer4_outputs(9174) <= not a or b;
    layer4_outputs(9175) <= not a;
    layer4_outputs(9176) <= a;
    layer4_outputs(9177) <= not b;
    layer4_outputs(9178) <= not a;
    layer4_outputs(9179) <= not b;
    layer4_outputs(9180) <= not a or b;
    layer4_outputs(9181) <= not (a xor b);
    layer4_outputs(9182) <= not (a xor b);
    layer4_outputs(9183) <= a xor b;
    layer4_outputs(9184) <= b and not a;
    layer4_outputs(9185) <= b;
    layer4_outputs(9186) <= a or b;
    layer4_outputs(9187) <= not (a and b);
    layer4_outputs(9188) <= not a or b;
    layer4_outputs(9189) <= a;
    layer4_outputs(9190) <= not (a xor b);
    layer4_outputs(9191) <= not b or a;
    layer4_outputs(9192) <= not a;
    layer4_outputs(9193) <= not a;
    layer4_outputs(9194) <= not b;
    layer4_outputs(9195) <= a or b;
    layer4_outputs(9196) <= a and b;
    layer4_outputs(9197) <= b and not a;
    layer4_outputs(9198) <= a;
    layer4_outputs(9199) <= a and not b;
    layer4_outputs(9200) <= a;
    layer4_outputs(9201) <= a xor b;
    layer4_outputs(9202) <= b and not a;
    layer4_outputs(9203) <= not a;
    layer4_outputs(9204) <= a or b;
    layer4_outputs(9205) <= a xor b;
    layer4_outputs(9206) <= a or b;
    layer4_outputs(9207) <= a and b;
    layer4_outputs(9208) <= not (a and b);
    layer4_outputs(9209) <= not (a xor b);
    layer4_outputs(9210) <= not a;
    layer4_outputs(9211) <= not b or a;
    layer4_outputs(9212) <= b;
    layer4_outputs(9213) <= a and b;
    layer4_outputs(9214) <= not b;
    layer4_outputs(9215) <= not (a and b);
    layer4_outputs(9216) <= not a;
    layer4_outputs(9217) <= not b;
    layer4_outputs(9218) <= not a or b;
    layer4_outputs(9219) <= not a;
    layer4_outputs(9220) <= not a or b;
    layer4_outputs(9221) <= a and b;
    layer4_outputs(9222) <= not (a xor b);
    layer4_outputs(9223) <= not (a xor b);
    layer4_outputs(9224) <= not (a and b);
    layer4_outputs(9225) <= not (a or b);
    layer4_outputs(9226) <= a or b;
    layer4_outputs(9227) <= not a;
    layer4_outputs(9228) <= a and not b;
    layer4_outputs(9229) <= not (a and b);
    layer4_outputs(9230) <= a or b;
    layer4_outputs(9231) <= b;
    layer4_outputs(9232) <= a and b;
    layer4_outputs(9233) <= a xor b;
    layer4_outputs(9234) <= b;
    layer4_outputs(9235) <= not (a and b);
    layer4_outputs(9236) <= a;
    layer4_outputs(9237) <= not b;
    layer4_outputs(9238) <= not (a xor b);
    layer4_outputs(9239) <= not (a or b);
    layer4_outputs(9240) <= b;
    layer4_outputs(9241) <= not b or a;
    layer4_outputs(9242) <= not (a or b);
    layer4_outputs(9243) <= a xor b;
    layer4_outputs(9244) <= b;
    layer4_outputs(9245) <= not b or a;
    layer4_outputs(9246) <= b;
    layer4_outputs(9247) <= a;
    layer4_outputs(9248) <= a and b;
    layer4_outputs(9249) <= a and not b;
    layer4_outputs(9250) <= a and not b;
    layer4_outputs(9251) <= not a;
    layer4_outputs(9252) <= not (a and b);
    layer4_outputs(9253) <= not b;
    layer4_outputs(9254) <= not a;
    layer4_outputs(9255) <= b and not a;
    layer4_outputs(9256) <= not (a xor b);
    layer4_outputs(9257) <= not (a or b);
    layer4_outputs(9258) <= b and not a;
    layer4_outputs(9259) <= b and not a;
    layer4_outputs(9260) <= not b;
    layer4_outputs(9261) <= not b;
    layer4_outputs(9262) <= a;
    layer4_outputs(9263) <= not (a xor b);
    layer4_outputs(9264) <= not (a or b);
    layer4_outputs(9265) <= a xor b;
    layer4_outputs(9266) <= not (a xor b);
    layer4_outputs(9267) <= not b or a;
    layer4_outputs(9268) <= b and not a;
    layer4_outputs(9269) <= a and not b;
    layer4_outputs(9270) <= a xor b;
    layer4_outputs(9271) <= not a;
    layer4_outputs(9272) <= not b;
    layer4_outputs(9273) <= b;
    layer4_outputs(9274) <= a and b;
    layer4_outputs(9275) <= a;
    layer4_outputs(9276) <= not (a or b);
    layer4_outputs(9277) <= not (a xor b);
    layer4_outputs(9278) <= a;
    layer4_outputs(9279) <= a xor b;
    layer4_outputs(9280) <= not (a xor b);
    layer4_outputs(9281) <= not a;
    layer4_outputs(9282) <= a xor b;
    layer4_outputs(9283) <= not b;
    layer4_outputs(9284) <= not b or a;
    layer4_outputs(9285) <= not b;
    layer4_outputs(9286) <= a or b;
    layer4_outputs(9287) <= not a;
    layer4_outputs(9288) <= not (a xor b);
    layer4_outputs(9289) <= not b;
    layer4_outputs(9290) <= not a;
    layer4_outputs(9291) <= a and b;
    layer4_outputs(9292) <= not b or a;
    layer4_outputs(9293) <= not a;
    layer4_outputs(9294) <= a and b;
    layer4_outputs(9295) <= not (a or b);
    layer4_outputs(9296) <= a xor b;
    layer4_outputs(9297) <= not (a xor b);
    layer4_outputs(9298) <= not (a and b);
    layer4_outputs(9299) <= not b or a;
    layer4_outputs(9300) <= not a;
    layer4_outputs(9301) <= a xor b;
    layer4_outputs(9302) <= b;
    layer4_outputs(9303) <= not (a xor b);
    layer4_outputs(9304) <= not a;
    layer4_outputs(9305) <= a;
    layer4_outputs(9306) <= b and not a;
    layer4_outputs(9307) <= b;
    layer4_outputs(9308) <= a xor b;
    layer4_outputs(9309) <= not b;
    layer4_outputs(9310) <= a xor b;
    layer4_outputs(9311) <= not a or b;
    layer4_outputs(9312) <= not (a or b);
    layer4_outputs(9313) <= b;
    layer4_outputs(9314) <= a;
    layer4_outputs(9315) <= not b;
    layer4_outputs(9316) <= not b;
    layer4_outputs(9317) <= b;
    layer4_outputs(9318) <= a;
    layer4_outputs(9319) <= b;
    layer4_outputs(9320) <= not a;
    layer4_outputs(9321) <= not b;
    layer4_outputs(9322) <= not a or b;
    layer4_outputs(9323) <= not (a xor b);
    layer4_outputs(9324) <= not (a and b);
    layer4_outputs(9325) <= not a;
    layer4_outputs(9326) <= a xor b;
    layer4_outputs(9327) <= not (a or b);
    layer4_outputs(9328) <= not (a xor b);
    layer4_outputs(9329) <= b;
    layer4_outputs(9330) <= a and b;
    layer4_outputs(9331) <= a and b;
    layer4_outputs(9332) <= not b;
    layer4_outputs(9333) <= not b;
    layer4_outputs(9334) <= a;
    layer4_outputs(9335) <= a;
    layer4_outputs(9336) <= 1'b0;
    layer4_outputs(9337) <= a;
    layer4_outputs(9338) <= not a or b;
    layer4_outputs(9339) <= not b or a;
    layer4_outputs(9340) <= a xor b;
    layer4_outputs(9341) <= a or b;
    layer4_outputs(9342) <= b;
    layer4_outputs(9343) <= a and b;
    layer4_outputs(9344) <= not b;
    layer4_outputs(9345) <= not (a xor b);
    layer4_outputs(9346) <= a xor b;
    layer4_outputs(9347) <= a and b;
    layer4_outputs(9348) <= a or b;
    layer4_outputs(9349) <= a xor b;
    layer4_outputs(9350) <= a and not b;
    layer4_outputs(9351) <= a or b;
    layer4_outputs(9352) <= not b;
    layer4_outputs(9353) <= not b or a;
    layer4_outputs(9354) <= b and not a;
    layer4_outputs(9355) <= a xor b;
    layer4_outputs(9356) <= b;
    layer4_outputs(9357) <= not b or a;
    layer4_outputs(9358) <= not a;
    layer4_outputs(9359) <= a or b;
    layer4_outputs(9360) <= b;
    layer4_outputs(9361) <= not (a and b);
    layer4_outputs(9362) <= not b;
    layer4_outputs(9363) <= not b or a;
    layer4_outputs(9364) <= not b or a;
    layer4_outputs(9365) <= a xor b;
    layer4_outputs(9366) <= not (a xor b);
    layer4_outputs(9367) <= a and not b;
    layer4_outputs(9368) <= b and not a;
    layer4_outputs(9369) <= not b or a;
    layer4_outputs(9370) <= not (a xor b);
    layer4_outputs(9371) <= not a;
    layer4_outputs(9372) <= a xor b;
    layer4_outputs(9373) <= b;
    layer4_outputs(9374) <= not a;
    layer4_outputs(9375) <= a;
    layer4_outputs(9376) <= not (a and b);
    layer4_outputs(9377) <= not b;
    layer4_outputs(9378) <= not a;
    layer4_outputs(9379) <= b and not a;
    layer4_outputs(9380) <= not a or b;
    layer4_outputs(9381) <= not b;
    layer4_outputs(9382) <= b;
    layer4_outputs(9383) <= not b;
    layer4_outputs(9384) <= not b;
    layer4_outputs(9385) <= not b;
    layer4_outputs(9386) <= not b;
    layer4_outputs(9387) <= a;
    layer4_outputs(9388) <= not (a or b);
    layer4_outputs(9389) <= not (a and b);
    layer4_outputs(9390) <= not b;
    layer4_outputs(9391) <= not a;
    layer4_outputs(9392) <= a xor b;
    layer4_outputs(9393) <= not (a xor b);
    layer4_outputs(9394) <= not a or b;
    layer4_outputs(9395) <= not (a xor b);
    layer4_outputs(9396) <= b and not a;
    layer4_outputs(9397) <= b;
    layer4_outputs(9398) <= b;
    layer4_outputs(9399) <= b;
    layer4_outputs(9400) <= not (a and b);
    layer4_outputs(9401) <= a;
    layer4_outputs(9402) <= not a or b;
    layer4_outputs(9403) <= not a or b;
    layer4_outputs(9404) <= not a;
    layer4_outputs(9405) <= a or b;
    layer4_outputs(9406) <= not (a xor b);
    layer4_outputs(9407) <= not a;
    layer4_outputs(9408) <= not b;
    layer4_outputs(9409) <= a or b;
    layer4_outputs(9410) <= b;
    layer4_outputs(9411) <= not b;
    layer4_outputs(9412) <= b;
    layer4_outputs(9413) <= a xor b;
    layer4_outputs(9414) <= b;
    layer4_outputs(9415) <= a and not b;
    layer4_outputs(9416) <= not b;
    layer4_outputs(9417) <= b and not a;
    layer4_outputs(9418) <= a or b;
    layer4_outputs(9419) <= b;
    layer4_outputs(9420) <= a xor b;
    layer4_outputs(9421) <= not b;
    layer4_outputs(9422) <= a;
    layer4_outputs(9423) <= not b;
    layer4_outputs(9424) <= not a;
    layer4_outputs(9425) <= b;
    layer4_outputs(9426) <= not a;
    layer4_outputs(9427) <= not b;
    layer4_outputs(9428) <= not a;
    layer4_outputs(9429) <= not (a and b);
    layer4_outputs(9430) <= a and b;
    layer4_outputs(9431) <= not b;
    layer4_outputs(9432) <= not (a xor b);
    layer4_outputs(9433) <= a;
    layer4_outputs(9434) <= not a or b;
    layer4_outputs(9435) <= not b or a;
    layer4_outputs(9436) <= a or b;
    layer4_outputs(9437) <= b;
    layer4_outputs(9438) <= not (a xor b);
    layer4_outputs(9439) <= not b;
    layer4_outputs(9440) <= b;
    layer4_outputs(9441) <= not b or a;
    layer4_outputs(9442) <= a;
    layer4_outputs(9443) <= b;
    layer4_outputs(9444) <= not a;
    layer4_outputs(9445) <= not a or b;
    layer4_outputs(9446) <= not (a xor b);
    layer4_outputs(9447) <= a xor b;
    layer4_outputs(9448) <= not b;
    layer4_outputs(9449) <= b;
    layer4_outputs(9450) <= a or b;
    layer4_outputs(9451) <= a xor b;
    layer4_outputs(9452) <= a xor b;
    layer4_outputs(9453) <= b;
    layer4_outputs(9454) <= a;
    layer4_outputs(9455) <= not b or a;
    layer4_outputs(9456) <= a;
    layer4_outputs(9457) <= not (a and b);
    layer4_outputs(9458) <= not (a xor b);
    layer4_outputs(9459) <= b;
    layer4_outputs(9460) <= a;
    layer4_outputs(9461) <= not (a or b);
    layer4_outputs(9462) <= a xor b;
    layer4_outputs(9463) <= not a or b;
    layer4_outputs(9464) <= not a;
    layer4_outputs(9465) <= not b;
    layer4_outputs(9466) <= a and not b;
    layer4_outputs(9467) <= a xor b;
    layer4_outputs(9468) <= not b;
    layer4_outputs(9469) <= not a;
    layer4_outputs(9470) <= not b or a;
    layer4_outputs(9471) <= a and b;
    layer4_outputs(9472) <= not b;
    layer4_outputs(9473) <= not (a and b);
    layer4_outputs(9474) <= not (a or b);
    layer4_outputs(9475) <= a and b;
    layer4_outputs(9476) <= not (a and b);
    layer4_outputs(9477) <= b;
    layer4_outputs(9478) <= not a;
    layer4_outputs(9479) <= not a or b;
    layer4_outputs(9480) <= a;
    layer4_outputs(9481) <= not (a xor b);
    layer4_outputs(9482) <= a and not b;
    layer4_outputs(9483) <= a;
    layer4_outputs(9484) <= a;
    layer4_outputs(9485) <= b and not a;
    layer4_outputs(9486) <= not a or b;
    layer4_outputs(9487) <= not b;
    layer4_outputs(9488) <= not (a xor b);
    layer4_outputs(9489) <= b and not a;
    layer4_outputs(9490) <= not b or a;
    layer4_outputs(9491) <= a and b;
    layer4_outputs(9492) <= not b;
    layer4_outputs(9493) <= a;
    layer4_outputs(9494) <= a xor b;
    layer4_outputs(9495) <= not (a xor b);
    layer4_outputs(9496) <= not a;
    layer4_outputs(9497) <= b;
    layer4_outputs(9498) <= not a or b;
    layer4_outputs(9499) <= not a or b;
    layer4_outputs(9500) <= not a or b;
    layer4_outputs(9501) <= a;
    layer4_outputs(9502) <= a and b;
    layer4_outputs(9503) <= 1'b1;
    layer4_outputs(9504) <= not b;
    layer4_outputs(9505) <= b;
    layer4_outputs(9506) <= not a;
    layer4_outputs(9507) <= a;
    layer4_outputs(9508) <= not (a xor b);
    layer4_outputs(9509) <= not b;
    layer4_outputs(9510) <= not b;
    layer4_outputs(9511) <= a xor b;
    layer4_outputs(9512) <= not b or a;
    layer4_outputs(9513) <= b;
    layer4_outputs(9514) <= not a or b;
    layer4_outputs(9515) <= not (a or b);
    layer4_outputs(9516) <= b;
    layer4_outputs(9517) <= a xor b;
    layer4_outputs(9518) <= a and b;
    layer4_outputs(9519) <= a and b;
    layer4_outputs(9520) <= a or b;
    layer4_outputs(9521) <= b and not a;
    layer4_outputs(9522) <= b;
    layer4_outputs(9523) <= a or b;
    layer4_outputs(9524) <= not (a and b);
    layer4_outputs(9525) <= a and not b;
    layer4_outputs(9526) <= not a;
    layer4_outputs(9527) <= a xor b;
    layer4_outputs(9528) <= not b;
    layer4_outputs(9529) <= a xor b;
    layer4_outputs(9530) <= a;
    layer4_outputs(9531) <= a and not b;
    layer4_outputs(9532) <= not a;
    layer4_outputs(9533) <= not b;
    layer4_outputs(9534) <= a xor b;
    layer4_outputs(9535) <= not a;
    layer4_outputs(9536) <= not a;
    layer4_outputs(9537) <= a and b;
    layer4_outputs(9538) <= not b;
    layer4_outputs(9539) <= not (a or b);
    layer4_outputs(9540) <= a or b;
    layer4_outputs(9541) <= not a;
    layer4_outputs(9542) <= a xor b;
    layer4_outputs(9543) <= a and b;
    layer4_outputs(9544) <= 1'b1;
    layer4_outputs(9545) <= a xor b;
    layer4_outputs(9546) <= a;
    layer4_outputs(9547) <= not b;
    layer4_outputs(9548) <= not a;
    layer4_outputs(9549) <= a or b;
    layer4_outputs(9550) <= a;
    layer4_outputs(9551) <= a or b;
    layer4_outputs(9552) <= a and b;
    layer4_outputs(9553) <= a xor b;
    layer4_outputs(9554) <= not b;
    layer4_outputs(9555) <= not a;
    layer4_outputs(9556) <= a xor b;
    layer4_outputs(9557) <= not a or b;
    layer4_outputs(9558) <= b;
    layer4_outputs(9559) <= a and not b;
    layer4_outputs(9560) <= a and b;
    layer4_outputs(9561) <= not b;
    layer4_outputs(9562) <= not a;
    layer4_outputs(9563) <= not a;
    layer4_outputs(9564) <= not (a and b);
    layer4_outputs(9565) <= not a or b;
    layer4_outputs(9566) <= not a or b;
    layer4_outputs(9567) <= a xor b;
    layer4_outputs(9568) <= b;
    layer4_outputs(9569) <= a xor b;
    layer4_outputs(9570) <= b;
    layer4_outputs(9571) <= not a;
    layer4_outputs(9572) <= not b;
    layer4_outputs(9573) <= not a or b;
    layer4_outputs(9574) <= a and b;
    layer4_outputs(9575) <= not a;
    layer4_outputs(9576) <= not a or b;
    layer4_outputs(9577) <= a xor b;
    layer4_outputs(9578) <= not b or a;
    layer4_outputs(9579) <= not a;
    layer4_outputs(9580) <= not (a xor b);
    layer4_outputs(9581) <= not (a or b);
    layer4_outputs(9582) <= not a;
    layer4_outputs(9583) <= not (a or b);
    layer4_outputs(9584) <= a;
    layer4_outputs(9585) <= not (a xor b);
    layer4_outputs(9586) <= a;
    layer4_outputs(9587) <= a and not b;
    layer4_outputs(9588) <= not (a or b);
    layer4_outputs(9589) <= not a;
    layer4_outputs(9590) <= not a;
    layer4_outputs(9591) <= a xor b;
    layer4_outputs(9592) <= a or b;
    layer4_outputs(9593) <= not (a xor b);
    layer4_outputs(9594) <= not a;
    layer4_outputs(9595) <= not a or b;
    layer4_outputs(9596) <= not (a and b);
    layer4_outputs(9597) <= a xor b;
    layer4_outputs(9598) <= a xor b;
    layer4_outputs(9599) <= not b;
    layer4_outputs(9600) <= b;
    layer4_outputs(9601) <= not b;
    layer4_outputs(9602) <= not a;
    layer4_outputs(9603) <= a and not b;
    layer4_outputs(9604) <= a;
    layer4_outputs(9605) <= not (a and b);
    layer4_outputs(9606) <= not (a and b);
    layer4_outputs(9607) <= a;
    layer4_outputs(9608) <= b;
    layer4_outputs(9609) <= b;
    layer4_outputs(9610) <= not (a xor b);
    layer4_outputs(9611) <= a and not b;
    layer4_outputs(9612) <= not (a or b);
    layer4_outputs(9613) <= not b;
    layer4_outputs(9614) <= not b;
    layer4_outputs(9615) <= not a;
    layer4_outputs(9616) <= not (a or b);
    layer4_outputs(9617) <= not b;
    layer4_outputs(9618) <= not b or a;
    layer4_outputs(9619) <= a;
    layer4_outputs(9620) <= not b;
    layer4_outputs(9621) <= b;
    layer4_outputs(9622) <= a and b;
    layer4_outputs(9623) <= a and not b;
    layer4_outputs(9624) <= not (a xor b);
    layer4_outputs(9625) <= not a;
    layer4_outputs(9626) <= not b or a;
    layer4_outputs(9627) <= not a;
    layer4_outputs(9628) <= not a;
    layer4_outputs(9629) <= not b;
    layer4_outputs(9630) <= not (a and b);
    layer4_outputs(9631) <= not b or a;
    layer4_outputs(9632) <= not b or a;
    layer4_outputs(9633) <= not (a or b);
    layer4_outputs(9634) <= not (a or b);
    layer4_outputs(9635) <= a and not b;
    layer4_outputs(9636) <= a;
    layer4_outputs(9637) <= not (a xor b);
    layer4_outputs(9638) <= not (a xor b);
    layer4_outputs(9639) <= a or b;
    layer4_outputs(9640) <= b and not a;
    layer4_outputs(9641) <= a and not b;
    layer4_outputs(9642) <= not b or a;
    layer4_outputs(9643) <= a xor b;
    layer4_outputs(9644) <= a;
    layer4_outputs(9645) <= a;
    layer4_outputs(9646) <= a and b;
    layer4_outputs(9647) <= not b;
    layer4_outputs(9648) <= not (a xor b);
    layer4_outputs(9649) <= b;
    layer4_outputs(9650) <= a xor b;
    layer4_outputs(9651) <= a;
    layer4_outputs(9652) <= a xor b;
    layer4_outputs(9653) <= not (a and b);
    layer4_outputs(9654) <= not (a or b);
    layer4_outputs(9655) <= a and not b;
    layer4_outputs(9656) <= b and not a;
    layer4_outputs(9657) <= not (a or b);
    layer4_outputs(9658) <= a;
    layer4_outputs(9659) <= b;
    layer4_outputs(9660) <= a and not b;
    layer4_outputs(9661) <= a or b;
    layer4_outputs(9662) <= a and b;
    layer4_outputs(9663) <= not b or a;
    layer4_outputs(9664) <= b and not a;
    layer4_outputs(9665) <= a and b;
    layer4_outputs(9666) <= not a;
    layer4_outputs(9667) <= b;
    layer4_outputs(9668) <= b;
    layer4_outputs(9669) <= a;
    layer4_outputs(9670) <= not b;
    layer4_outputs(9671) <= b and not a;
    layer4_outputs(9672) <= b and not a;
    layer4_outputs(9673) <= a xor b;
    layer4_outputs(9674) <= not b;
    layer4_outputs(9675) <= a and not b;
    layer4_outputs(9676) <= b;
    layer4_outputs(9677) <= b and not a;
    layer4_outputs(9678) <= not (a xor b);
    layer4_outputs(9679) <= not a;
    layer4_outputs(9680) <= a or b;
    layer4_outputs(9681) <= not a;
    layer4_outputs(9682) <= b;
    layer4_outputs(9683) <= not a or b;
    layer4_outputs(9684) <= not b or a;
    layer4_outputs(9685) <= not b;
    layer4_outputs(9686) <= a;
    layer4_outputs(9687) <= a and b;
    layer4_outputs(9688) <= not a or b;
    layer4_outputs(9689) <= not b;
    layer4_outputs(9690) <= not (a and b);
    layer4_outputs(9691) <= a;
    layer4_outputs(9692) <= a and b;
    layer4_outputs(9693) <= a and b;
    layer4_outputs(9694) <= b;
    layer4_outputs(9695) <= a xor b;
    layer4_outputs(9696) <= a and b;
    layer4_outputs(9697) <= not b;
    layer4_outputs(9698) <= a or b;
    layer4_outputs(9699) <= a;
    layer4_outputs(9700) <= a;
    layer4_outputs(9701) <= not b;
    layer4_outputs(9702) <= a and not b;
    layer4_outputs(9703) <= a and b;
    layer4_outputs(9704) <= a xor b;
    layer4_outputs(9705) <= a and b;
    layer4_outputs(9706) <= a;
    layer4_outputs(9707) <= not a;
    layer4_outputs(9708) <= a or b;
    layer4_outputs(9709) <= not b;
    layer4_outputs(9710) <= b and not a;
    layer4_outputs(9711) <= a;
    layer4_outputs(9712) <= a and b;
    layer4_outputs(9713) <= a and b;
    layer4_outputs(9714) <= not a or b;
    layer4_outputs(9715) <= a xor b;
    layer4_outputs(9716) <= not (a and b);
    layer4_outputs(9717) <= a;
    layer4_outputs(9718) <= b;
    layer4_outputs(9719) <= a or b;
    layer4_outputs(9720) <= a xor b;
    layer4_outputs(9721) <= a xor b;
    layer4_outputs(9722) <= a or b;
    layer4_outputs(9723) <= not a or b;
    layer4_outputs(9724) <= a xor b;
    layer4_outputs(9725) <= a and b;
    layer4_outputs(9726) <= b;
    layer4_outputs(9727) <= a;
    layer4_outputs(9728) <= 1'b1;
    layer4_outputs(9729) <= a xor b;
    layer4_outputs(9730) <= b and not a;
    layer4_outputs(9731) <= b;
    layer4_outputs(9732) <= b;
    layer4_outputs(9733) <= not a or b;
    layer4_outputs(9734) <= not (a or b);
    layer4_outputs(9735) <= b and not a;
    layer4_outputs(9736) <= a;
    layer4_outputs(9737) <= not b;
    layer4_outputs(9738) <= not (a xor b);
    layer4_outputs(9739) <= not a or b;
    layer4_outputs(9740) <= a or b;
    layer4_outputs(9741) <= not (a xor b);
    layer4_outputs(9742) <= b and not a;
    layer4_outputs(9743) <= not a;
    layer4_outputs(9744) <= b;
    layer4_outputs(9745) <= a or b;
    layer4_outputs(9746) <= a;
    layer4_outputs(9747) <= a;
    layer4_outputs(9748) <= not b or a;
    layer4_outputs(9749) <= a xor b;
    layer4_outputs(9750) <= not b;
    layer4_outputs(9751) <= not (a and b);
    layer4_outputs(9752) <= not b or a;
    layer4_outputs(9753) <= not a;
    layer4_outputs(9754) <= not b or a;
    layer4_outputs(9755) <= not (a xor b);
    layer4_outputs(9756) <= not b;
    layer4_outputs(9757) <= not a or b;
    layer4_outputs(9758) <= not a;
    layer4_outputs(9759) <= not (a or b);
    layer4_outputs(9760) <= a and b;
    layer4_outputs(9761) <= not b;
    layer4_outputs(9762) <= not (a or b);
    layer4_outputs(9763) <= a;
    layer4_outputs(9764) <= not b;
    layer4_outputs(9765) <= a;
    layer4_outputs(9766) <= b;
    layer4_outputs(9767) <= not (a xor b);
    layer4_outputs(9768) <= b;
    layer4_outputs(9769) <= a or b;
    layer4_outputs(9770) <= not (a or b);
    layer4_outputs(9771) <= b;
    layer4_outputs(9772) <= not (a or b);
    layer4_outputs(9773) <= a;
    layer4_outputs(9774) <= not a;
    layer4_outputs(9775) <= not (a xor b);
    layer4_outputs(9776) <= not a or b;
    layer4_outputs(9777) <= not b;
    layer4_outputs(9778) <= b;
    layer4_outputs(9779) <= a xor b;
    layer4_outputs(9780) <= not b;
    layer4_outputs(9781) <= not (a xor b);
    layer4_outputs(9782) <= a;
    layer4_outputs(9783) <= b;
    layer4_outputs(9784) <= a and not b;
    layer4_outputs(9785) <= not b or a;
    layer4_outputs(9786) <= b;
    layer4_outputs(9787) <= b;
    layer4_outputs(9788) <= b;
    layer4_outputs(9789) <= not a;
    layer4_outputs(9790) <= a and b;
    layer4_outputs(9791) <= not (a xor b);
    layer4_outputs(9792) <= b;
    layer4_outputs(9793) <= b;
    layer4_outputs(9794) <= a;
    layer4_outputs(9795) <= not b;
    layer4_outputs(9796) <= not b;
    layer4_outputs(9797) <= not a;
    layer4_outputs(9798) <= a or b;
    layer4_outputs(9799) <= not a or b;
    layer4_outputs(9800) <= a;
    layer4_outputs(9801) <= b;
    layer4_outputs(9802) <= b;
    layer4_outputs(9803) <= not a or b;
    layer4_outputs(9804) <= not (a or b);
    layer4_outputs(9805) <= not a;
    layer4_outputs(9806) <= not b;
    layer4_outputs(9807) <= a;
    layer4_outputs(9808) <= a;
    layer4_outputs(9809) <= not a;
    layer4_outputs(9810) <= a;
    layer4_outputs(9811) <= a;
    layer4_outputs(9812) <= a xor b;
    layer4_outputs(9813) <= not b or a;
    layer4_outputs(9814) <= not (a xor b);
    layer4_outputs(9815) <= not (a or b);
    layer4_outputs(9816) <= a xor b;
    layer4_outputs(9817) <= b;
    layer4_outputs(9818) <= not b;
    layer4_outputs(9819) <= not b or a;
    layer4_outputs(9820) <= not a;
    layer4_outputs(9821) <= a;
    layer4_outputs(9822) <= not (a or b);
    layer4_outputs(9823) <= a xor b;
    layer4_outputs(9824) <= a and b;
    layer4_outputs(9825) <= not a;
    layer4_outputs(9826) <= a;
    layer4_outputs(9827) <= b;
    layer4_outputs(9828) <= 1'b0;
    layer4_outputs(9829) <= not b;
    layer4_outputs(9830) <= a and not b;
    layer4_outputs(9831) <= not b;
    layer4_outputs(9832) <= a;
    layer4_outputs(9833) <= a;
    layer4_outputs(9834) <= not a or b;
    layer4_outputs(9835) <= b and not a;
    layer4_outputs(9836) <= not a;
    layer4_outputs(9837) <= not b;
    layer4_outputs(9838) <= not b;
    layer4_outputs(9839) <= b;
    layer4_outputs(9840) <= not b or a;
    layer4_outputs(9841) <= not b or a;
    layer4_outputs(9842) <= 1'b0;
    layer4_outputs(9843) <= not (a xor b);
    layer4_outputs(9844) <= not (a and b);
    layer4_outputs(9845) <= not (a xor b);
    layer4_outputs(9846) <= b;
    layer4_outputs(9847) <= b;
    layer4_outputs(9848) <= not a;
    layer4_outputs(9849) <= not (a xor b);
    layer4_outputs(9850) <= not b or a;
    layer4_outputs(9851) <= not a;
    layer4_outputs(9852) <= a;
    layer4_outputs(9853) <= not b or a;
    layer4_outputs(9854) <= not a or b;
    layer4_outputs(9855) <= b;
    layer4_outputs(9856) <= not (a and b);
    layer4_outputs(9857) <= not a;
    layer4_outputs(9858) <= not (a xor b);
    layer4_outputs(9859) <= not b;
    layer4_outputs(9860) <= a or b;
    layer4_outputs(9861) <= a;
    layer4_outputs(9862) <= a xor b;
    layer4_outputs(9863) <= a;
    layer4_outputs(9864) <= a and not b;
    layer4_outputs(9865) <= a;
    layer4_outputs(9866) <= a or b;
    layer4_outputs(9867) <= not a;
    layer4_outputs(9868) <= a and not b;
    layer4_outputs(9869) <= a;
    layer4_outputs(9870) <= not a or b;
    layer4_outputs(9871) <= not (a xor b);
    layer4_outputs(9872) <= b and not a;
    layer4_outputs(9873) <= not a or b;
    layer4_outputs(9874) <= not a;
    layer4_outputs(9875) <= b;
    layer4_outputs(9876) <= b;
    layer4_outputs(9877) <= not (a xor b);
    layer4_outputs(9878) <= b;
    layer4_outputs(9879) <= not b or a;
    layer4_outputs(9880) <= a;
    layer4_outputs(9881) <= not (a xor b);
    layer4_outputs(9882) <= not a;
    layer4_outputs(9883) <= a and b;
    layer4_outputs(9884) <= not b;
    layer4_outputs(9885) <= not a;
    layer4_outputs(9886) <= b;
    layer4_outputs(9887) <= a xor b;
    layer4_outputs(9888) <= not b or a;
    layer4_outputs(9889) <= a;
    layer4_outputs(9890) <= a xor b;
    layer4_outputs(9891) <= not (a and b);
    layer4_outputs(9892) <= a and b;
    layer4_outputs(9893) <= not b;
    layer4_outputs(9894) <= not (a xor b);
    layer4_outputs(9895) <= a or b;
    layer4_outputs(9896) <= not (a or b);
    layer4_outputs(9897) <= b;
    layer4_outputs(9898) <= not a;
    layer4_outputs(9899) <= not (a xor b);
    layer4_outputs(9900) <= not b;
    layer4_outputs(9901) <= not (a and b);
    layer4_outputs(9902) <= not a or b;
    layer4_outputs(9903) <= not b;
    layer4_outputs(9904) <= a xor b;
    layer4_outputs(9905) <= a or b;
    layer4_outputs(9906) <= a;
    layer4_outputs(9907) <= not (a and b);
    layer4_outputs(9908) <= b;
    layer4_outputs(9909) <= a xor b;
    layer4_outputs(9910) <= not (a xor b);
    layer4_outputs(9911) <= not b or a;
    layer4_outputs(9912) <= b;
    layer4_outputs(9913) <= b;
    layer4_outputs(9914) <= not (a or b);
    layer4_outputs(9915) <= a and not b;
    layer4_outputs(9916) <= a and b;
    layer4_outputs(9917) <= not b;
    layer4_outputs(9918) <= a and not b;
    layer4_outputs(9919) <= not b;
    layer4_outputs(9920) <= not (a or b);
    layer4_outputs(9921) <= a;
    layer4_outputs(9922) <= a;
    layer4_outputs(9923) <= not (a or b);
    layer4_outputs(9924) <= not a;
    layer4_outputs(9925) <= a;
    layer4_outputs(9926) <= a and not b;
    layer4_outputs(9927) <= a and b;
    layer4_outputs(9928) <= not b;
    layer4_outputs(9929) <= a and b;
    layer4_outputs(9930) <= a or b;
    layer4_outputs(9931) <= not a;
    layer4_outputs(9932) <= not (a and b);
    layer4_outputs(9933) <= b;
    layer4_outputs(9934) <= not a;
    layer4_outputs(9935) <= a or b;
    layer4_outputs(9936) <= a;
    layer4_outputs(9937) <= a;
    layer4_outputs(9938) <= a;
    layer4_outputs(9939) <= b;
    layer4_outputs(9940) <= a or b;
    layer4_outputs(9941) <= b and not a;
    layer4_outputs(9942) <= b and not a;
    layer4_outputs(9943) <= a xor b;
    layer4_outputs(9944) <= b and not a;
    layer4_outputs(9945) <= a or b;
    layer4_outputs(9946) <= a and not b;
    layer4_outputs(9947) <= a;
    layer4_outputs(9948) <= a xor b;
    layer4_outputs(9949) <= not (a and b);
    layer4_outputs(9950) <= not (a or b);
    layer4_outputs(9951) <= not (a xor b);
    layer4_outputs(9952) <= a xor b;
    layer4_outputs(9953) <= a and b;
    layer4_outputs(9954) <= not a;
    layer4_outputs(9955) <= not a;
    layer4_outputs(9956) <= a;
    layer4_outputs(9957) <= a and not b;
    layer4_outputs(9958) <= a;
    layer4_outputs(9959) <= not (a xor b);
    layer4_outputs(9960) <= a or b;
    layer4_outputs(9961) <= not b;
    layer4_outputs(9962) <= not a;
    layer4_outputs(9963) <= not (a or b);
    layer4_outputs(9964) <= not (a xor b);
    layer4_outputs(9965) <= b;
    layer4_outputs(9966) <= not (a or b);
    layer4_outputs(9967) <= not b;
    layer4_outputs(9968) <= b and not a;
    layer4_outputs(9969) <= a xor b;
    layer4_outputs(9970) <= b;
    layer4_outputs(9971) <= not b;
    layer4_outputs(9972) <= 1'b1;
    layer4_outputs(9973) <= not (a xor b);
    layer4_outputs(9974) <= not a;
    layer4_outputs(9975) <= a and b;
    layer4_outputs(9976) <= b;
    layer4_outputs(9977) <= a and b;
    layer4_outputs(9978) <= not b or a;
    layer4_outputs(9979) <= a xor b;
    layer4_outputs(9980) <= a xor b;
    layer4_outputs(9981) <= 1'b0;
    layer4_outputs(9982) <= a and b;
    layer4_outputs(9983) <= a and not b;
    layer4_outputs(9984) <= not a or b;
    layer4_outputs(9985) <= a;
    layer4_outputs(9986) <= not b or a;
    layer4_outputs(9987) <= b;
    layer4_outputs(9988) <= a and not b;
    layer4_outputs(9989) <= b and not a;
    layer4_outputs(9990) <= a or b;
    layer4_outputs(9991) <= b and not a;
    layer4_outputs(9992) <= a and not b;
    layer4_outputs(9993) <= b;
    layer4_outputs(9994) <= not a;
    layer4_outputs(9995) <= b and not a;
    layer4_outputs(9996) <= b and not a;
    layer4_outputs(9997) <= not (a or b);
    layer4_outputs(9998) <= not a or b;
    layer4_outputs(9999) <= a and not b;
    layer4_outputs(10000) <= a and b;
    layer4_outputs(10001) <= a and not b;
    layer4_outputs(10002) <= not (a or b);
    layer4_outputs(10003) <= a xor b;
    layer4_outputs(10004) <= a and not b;
    layer4_outputs(10005) <= not (a and b);
    layer4_outputs(10006) <= not b;
    layer4_outputs(10007) <= not (a xor b);
    layer4_outputs(10008) <= not b;
    layer4_outputs(10009) <= b and not a;
    layer4_outputs(10010) <= not (a xor b);
    layer4_outputs(10011) <= not a;
    layer4_outputs(10012) <= b;
    layer4_outputs(10013) <= not (a or b);
    layer4_outputs(10014) <= not b;
    layer4_outputs(10015) <= a xor b;
    layer4_outputs(10016) <= a xor b;
    layer4_outputs(10017) <= not b or a;
    layer4_outputs(10018) <= a and b;
    layer4_outputs(10019) <= a xor b;
    layer4_outputs(10020) <= a or b;
    layer4_outputs(10021) <= b;
    layer4_outputs(10022) <= b;
    layer4_outputs(10023) <= a xor b;
    layer4_outputs(10024) <= b and not a;
    layer4_outputs(10025) <= a or b;
    layer4_outputs(10026) <= not b or a;
    layer4_outputs(10027) <= b and not a;
    layer4_outputs(10028) <= a;
    layer4_outputs(10029) <= a and b;
    layer4_outputs(10030) <= not (a or b);
    layer4_outputs(10031) <= not a;
    layer4_outputs(10032) <= a and not b;
    layer4_outputs(10033) <= b;
    layer4_outputs(10034) <= b;
    layer4_outputs(10035) <= not (a xor b);
    layer4_outputs(10036) <= not a or b;
    layer4_outputs(10037) <= not b;
    layer4_outputs(10038) <= a and b;
    layer4_outputs(10039) <= not b;
    layer4_outputs(10040) <= b;
    layer4_outputs(10041) <= not (a and b);
    layer4_outputs(10042) <= not a or b;
    layer4_outputs(10043) <= b;
    layer4_outputs(10044) <= not (a xor b);
    layer4_outputs(10045) <= b;
    layer4_outputs(10046) <= b and not a;
    layer4_outputs(10047) <= not a or b;
    layer4_outputs(10048) <= not a or b;
    layer4_outputs(10049) <= not a;
    layer4_outputs(10050) <= a;
    layer4_outputs(10051) <= a or b;
    layer4_outputs(10052) <= not (a or b);
    layer4_outputs(10053) <= b and not a;
    layer4_outputs(10054) <= not a;
    layer4_outputs(10055) <= b;
    layer4_outputs(10056) <= a and not b;
    layer4_outputs(10057) <= not a;
    layer4_outputs(10058) <= not (a and b);
    layer4_outputs(10059) <= not a;
    layer4_outputs(10060) <= not (a xor b);
    layer4_outputs(10061) <= not a or b;
    layer4_outputs(10062) <= b;
    layer4_outputs(10063) <= not (a and b);
    layer4_outputs(10064) <= not b;
    layer4_outputs(10065) <= not (a or b);
    layer4_outputs(10066) <= not (a xor b);
    layer4_outputs(10067) <= a and not b;
    layer4_outputs(10068) <= not (a xor b);
    layer4_outputs(10069) <= a xor b;
    layer4_outputs(10070) <= b;
    layer4_outputs(10071) <= a;
    layer4_outputs(10072) <= not b;
    layer4_outputs(10073) <= a or b;
    layer4_outputs(10074) <= a;
    layer4_outputs(10075) <= a xor b;
    layer4_outputs(10076) <= not b;
    layer4_outputs(10077) <= not b or a;
    layer4_outputs(10078) <= not a;
    layer4_outputs(10079) <= a;
    layer4_outputs(10080) <= a;
    layer4_outputs(10081) <= not b or a;
    layer4_outputs(10082) <= a or b;
    layer4_outputs(10083) <= a and not b;
    layer4_outputs(10084) <= not a;
    layer4_outputs(10085) <= not b or a;
    layer4_outputs(10086) <= a or b;
    layer4_outputs(10087) <= a and not b;
    layer4_outputs(10088) <= not b;
    layer4_outputs(10089) <= a xor b;
    layer4_outputs(10090) <= not b;
    layer4_outputs(10091) <= not a or b;
    layer4_outputs(10092) <= a;
    layer4_outputs(10093) <= not a;
    layer4_outputs(10094) <= a xor b;
    layer4_outputs(10095) <= not b;
    layer4_outputs(10096) <= not (a and b);
    layer4_outputs(10097) <= not a or b;
    layer4_outputs(10098) <= b;
    layer4_outputs(10099) <= b;
    layer4_outputs(10100) <= not b or a;
    layer4_outputs(10101) <= not (a xor b);
    layer4_outputs(10102) <= not b or a;
    layer4_outputs(10103) <= a xor b;
    layer4_outputs(10104) <= a or b;
    layer4_outputs(10105) <= not b;
    layer4_outputs(10106) <= a xor b;
    layer4_outputs(10107) <= b;
    layer4_outputs(10108) <= b and not a;
    layer4_outputs(10109) <= a and not b;
    layer4_outputs(10110) <= b and not a;
    layer4_outputs(10111) <= b;
    layer4_outputs(10112) <= a xor b;
    layer4_outputs(10113) <= not b or a;
    layer4_outputs(10114) <= not (a or b);
    layer4_outputs(10115) <= a;
    layer4_outputs(10116) <= not a or b;
    layer4_outputs(10117) <= not (a xor b);
    layer4_outputs(10118) <= b;
    layer4_outputs(10119) <= not a or b;
    layer4_outputs(10120) <= a;
    layer4_outputs(10121) <= not a or b;
    layer4_outputs(10122) <= b and not a;
    layer4_outputs(10123) <= b and not a;
    layer4_outputs(10124) <= not a or b;
    layer4_outputs(10125) <= not b or a;
    layer4_outputs(10126) <= not b;
    layer4_outputs(10127) <= not a;
    layer4_outputs(10128) <= 1'b0;
    layer4_outputs(10129) <= a xor b;
    layer4_outputs(10130) <= not b;
    layer4_outputs(10131) <= a and not b;
    layer4_outputs(10132) <= not a;
    layer4_outputs(10133) <= not a;
    layer4_outputs(10134) <= b;
    layer4_outputs(10135) <= not a;
    layer4_outputs(10136) <= not a;
    layer4_outputs(10137) <= not b;
    layer4_outputs(10138) <= a xor b;
    layer4_outputs(10139) <= not (a xor b);
    layer4_outputs(10140) <= a;
    layer4_outputs(10141) <= b and not a;
    layer4_outputs(10142) <= not a or b;
    layer4_outputs(10143) <= a and not b;
    layer4_outputs(10144) <= a xor b;
    layer4_outputs(10145) <= not a;
    layer4_outputs(10146) <= not b;
    layer4_outputs(10147) <= not a or b;
    layer4_outputs(10148) <= not (a or b);
    layer4_outputs(10149) <= not b;
    layer4_outputs(10150) <= not a;
    layer4_outputs(10151) <= not (a xor b);
    layer4_outputs(10152) <= a;
    layer4_outputs(10153) <= a and not b;
    layer4_outputs(10154) <= a xor b;
    layer4_outputs(10155) <= b and not a;
    layer4_outputs(10156) <= a xor b;
    layer4_outputs(10157) <= b;
    layer4_outputs(10158) <= a and not b;
    layer4_outputs(10159) <= a;
    layer4_outputs(10160) <= a;
    layer4_outputs(10161) <= not (a or b);
    layer4_outputs(10162) <= a xor b;
    layer4_outputs(10163) <= not b or a;
    layer4_outputs(10164) <= not (a xor b);
    layer4_outputs(10165) <= not (a xor b);
    layer4_outputs(10166) <= not b;
    layer4_outputs(10167) <= b;
    layer4_outputs(10168) <= not a;
    layer4_outputs(10169) <= b;
    layer4_outputs(10170) <= not a;
    layer4_outputs(10171) <= not b;
    layer4_outputs(10172) <= a and b;
    layer4_outputs(10173) <= not b;
    layer4_outputs(10174) <= a or b;
    layer4_outputs(10175) <= a and b;
    layer4_outputs(10176) <= a;
    layer4_outputs(10177) <= b;
    layer4_outputs(10178) <= not (a or b);
    layer4_outputs(10179) <= a and not b;
    layer4_outputs(10180) <= b;
    layer4_outputs(10181) <= not a;
    layer4_outputs(10182) <= not (a or b);
    layer4_outputs(10183) <= not b;
    layer4_outputs(10184) <= a;
    layer4_outputs(10185) <= not a;
    layer4_outputs(10186) <= a or b;
    layer4_outputs(10187) <= not a or b;
    layer4_outputs(10188) <= not a;
    layer4_outputs(10189) <= a or b;
    layer4_outputs(10190) <= b and not a;
    layer4_outputs(10191) <= not (a xor b);
    layer4_outputs(10192) <= a and b;
    layer4_outputs(10193) <= a or b;
    layer4_outputs(10194) <= not a;
    layer4_outputs(10195) <= not (a or b);
    layer4_outputs(10196) <= not a or b;
    layer4_outputs(10197) <= not a or b;
    layer4_outputs(10198) <= not a;
    layer4_outputs(10199) <= a;
    layer4_outputs(10200) <= a and b;
    layer4_outputs(10201) <= b;
    layer4_outputs(10202) <= not a;
    layer4_outputs(10203) <= a xor b;
    layer4_outputs(10204) <= not a or b;
    layer4_outputs(10205) <= not a or b;
    layer4_outputs(10206) <= a;
    layer4_outputs(10207) <= a;
    layer4_outputs(10208) <= a and b;
    layer4_outputs(10209) <= b;
    layer4_outputs(10210) <= not (a and b);
    layer4_outputs(10211) <= a;
    layer4_outputs(10212) <= not a or b;
    layer4_outputs(10213) <= a or b;
    layer4_outputs(10214) <= not b or a;
    layer4_outputs(10215) <= not (a xor b);
    layer4_outputs(10216) <= a or b;
    layer4_outputs(10217) <= not a;
    layer4_outputs(10218) <= not b;
    layer4_outputs(10219) <= a and b;
    layer4_outputs(10220) <= not b;
    layer4_outputs(10221) <= not (a and b);
    layer4_outputs(10222) <= b;
    layer4_outputs(10223) <= not (a and b);
    layer4_outputs(10224) <= not a or b;
    layer4_outputs(10225) <= not (a xor b);
    layer4_outputs(10226) <= b and not a;
    layer4_outputs(10227) <= b;
    layer4_outputs(10228) <= b;
    layer4_outputs(10229) <= a;
    layer4_outputs(10230) <= a and not b;
    layer4_outputs(10231) <= b;
    layer4_outputs(10232) <= not (a and b);
    layer4_outputs(10233) <= not (a and b);
    layer4_outputs(10234) <= not (a xor b);
    layer4_outputs(10235) <= a;
    layer4_outputs(10236) <= not (a xor b);
    layer4_outputs(10237) <= a;
    layer4_outputs(10238) <= not b;
    layer4_outputs(10239) <= b;
    outputs(0) <= not a or b;
    outputs(1) <= b;
    outputs(2) <= b and not a;
    outputs(3) <= a and not b;
    outputs(4) <= not a or b;
    outputs(5) <= not b;
    outputs(6) <= a xor b;
    outputs(7) <= not (a or b);
    outputs(8) <= not (a and b);
    outputs(9) <= not a;
    outputs(10) <= not a or b;
    outputs(11) <= not a;
    outputs(12) <= b;
    outputs(13) <= not (a and b);
    outputs(14) <= a xor b;
    outputs(15) <= not (a and b);
    outputs(16) <= not a;
    outputs(17) <= not b;
    outputs(18) <= not (a and b);
    outputs(19) <= a xor b;
    outputs(20) <= a xor b;
    outputs(21) <= not (a xor b);
    outputs(22) <= not b;
    outputs(23) <= not b or a;
    outputs(24) <= not (a xor b);
    outputs(25) <= not (a or b);
    outputs(26) <= a and b;
    outputs(27) <= not b;
    outputs(28) <= a xor b;
    outputs(29) <= a and b;
    outputs(30) <= b;
    outputs(31) <= a xor b;
    outputs(32) <= b;
    outputs(33) <= not b;
    outputs(34) <= not a;
    outputs(35) <= not (a and b);
    outputs(36) <= b;
    outputs(37) <= b;
    outputs(38) <= not (a xor b);
    outputs(39) <= b;
    outputs(40) <= b;
    outputs(41) <= not b;
    outputs(42) <= b;
    outputs(43) <= b;
    outputs(44) <= b and not a;
    outputs(45) <= a;
    outputs(46) <= b;
    outputs(47) <= not (a and b);
    outputs(48) <= a or b;
    outputs(49) <= b;
    outputs(50) <= a and not b;
    outputs(51) <= a;
    outputs(52) <= b;
    outputs(53) <= a;
    outputs(54) <= not (a xor b);
    outputs(55) <= b and not a;
    outputs(56) <= b;
    outputs(57) <= not (a or b);
    outputs(58) <= a;
    outputs(59) <= a;
    outputs(60) <= not (a xor b);
    outputs(61) <= not a;
    outputs(62) <= a and b;
    outputs(63) <= not (a xor b);
    outputs(64) <= not (a or b);
    outputs(65) <= a and b;
    outputs(66) <= a xor b;
    outputs(67) <= a and b;
    outputs(68) <= b;
    outputs(69) <= a;
    outputs(70) <= b and not a;
    outputs(71) <= a;
    outputs(72) <= not a;
    outputs(73) <= not (a xor b);
    outputs(74) <= b;
    outputs(75) <= not (a xor b);
    outputs(76) <= a and b;
    outputs(77) <= a xor b;
    outputs(78) <= not (a or b);
    outputs(79) <= b;
    outputs(80) <= not (a or b);
    outputs(81) <= b;
    outputs(82) <= a;
    outputs(83) <= not b;
    outputs(84) <= a and not b;
    outputs(85) <= not b;
    outputs(86) <= b and not a;
    outputs(87) <= not (a xor b);
    outputs(88) <= not b;
    outputs(89) <= not (a xor b);
    outputs(90) <= a xor b;
    outputs(91) <= b;
    outputs(92) <= a;
    outputs(93) <= b;
    outputs(94) <= not b;
    outputs(95) <= not (a xor b);
    outputs(96) <= not b;
    outputs(97) <= not a;
    outputs(98) <= not (a xor b);
    outputs(99) <= a xor b;
    outputs(100) <= not b;
    outputs(101) <= a xor b;
    outputs(102) <= a xor b;
    outputs(103) <= not b;
    outputs(104) <= b and not a;
    outputs(105) <= not (a xor b);
    outputs(106) <= a and not b;
    outputs(107) <= not (a xor b);
    outputs(108) <= not a or b;
    outputs(109) <= not (a or b);
    outputs(110) <= a and b;
    outputs(111) <= a xor b;
    outputs(112) <= not (a xor b);
    outputs(113) <= a xor b;
    outputs(114) <= a;
    outputs(115) <= a xor b;
    outputs(116) <= not (a and b);
    outputs(117) <= a;
    outputs(118) <= a or b;
    outputs(119) <= not b;
    outputs(120) <= not (a or b);
    outputs(121) <= not a or b;
    outputs(122) <= a xor b;
    outputs(123) <= b;
    outputs(124) <= not b;
    outputs(125) <= a;
    outputs(126) <= a xor b;
    outputs(127) <= b;
    outputs(128) <= not a;
    outputs(129) <= not a;
    outputs(130) <= a;
    outputs(131) <= a and not b;
    outputs(132) <= not a;
    outputs(133) <= a xor b;
    outputs(134) <= not (a xor b);
    outputs(135) <= not (a xor b);
    outputs(136) <= not b;
    outputs(137) <= b;
    outputs(138) <= not b;
    outputs(139) <= not b;
    outputs(140) <= not b;
    outputs(141) <= not b;
    outputs(142) <= b and not a;
    outputs(143) <= b and not a;
    outputs(144) <= not (a and b);
    outputs(145) <= not (a xor b);
    outputs(146) <= not b;
    outputs(147) <= b and not a;
    outputs(148) <= not a;
    outputs(149) <= not (a xor b);
    outputs(150) <= a xor b;
    outputs(151) <= not (a xor b);
    outputs(152) <= b;
    outputs(153) <= a and b;
    outputs(154) <= a and b;
    outputs(155) <= not b;
    outputs(156) <= not (a and b);
    outputs(157) <= not b or a;
    outputs(158) <= not (a xor b);
    outputs(159) <= a;
    outputs(160) <= b;
    outputs(161) <= not a;
    outputs(162) <= a and not b;
    outputs(163) <= a and b;
    outputs(164) <= not a or b;
    outputs(165) <= not (a xor b);
    outputs(166) <= a;
    outputs(167) <= not (a xor b);
    outputs(168) <= b;
    outputs(169) <= b and not a;
    outputs(170) <= not b;
    outputs(171) <= not (a xor b);
    outputs(172) <= not (a xor b);
    outputs(173) <= not a;
    outputs(174) <= a;
    outputs(175) <= a and not b;
    outputs(176) <= b and not a;
    outputs(177) <= a and not b;
    outputs(178) <= b;
    outputs(179) <= not (a xor b);
    outputs(180) <= a and not b;
    outputs(181) <= not (a xor b);
    outputs(182) <= not a;
    outputs(183) <= not a;
    outputs(184) <= not (a xor b);
    outputs(185) <= a;
    outputs(186) <= a xor b;
    outputs(187) <= not (a xor b);
    outputs(188) <= not a;
    outputs(189) <= b;
    outputs(190) <= not a;
    outputs(191) <= a;
    outputs(192) <= b;
    outputs(193) <= not b or a;
    outputs(194) <= a;
    outputs(195) <= b;
    outputs(196) <= a;
    outputs(197) <= a and b;
    outputs(198) <= not (a xor b);
    outputs(199) <= not (a xor b);
    outputs(200) <= b and not a;
    outputs(201) <= b and not a;
    outputs(202) <= b and not a;
    outputs(203) <= a xor b;
    outputs(204) <= a;
    outputs(205) <= a and not b;
    outputs(206) <= not (a xor b);
    outputs(207) <= b;
    outputs(208) <= not (a or b);
    outputs(209) <= a;
    outputs(210) <= not (a xor b);
    outputs(211) <= not a or b;
    outputs(212) <= not (a xor b);
    outputs(213) <= a and not b;
    outputs(214) <= not b;
    outputs(215) <= a;
    outputs(216) <= a xor b;
    outputs(217) <= not (a xor b);
    outputs(218) <= b;
    outputs(219) <= a or b;
    outputs(220) <= a;
    outputs(221) <= not (a xor b);
    outputs(222) <= a;
    outputs(223) <= a and b;
    outputs(224) <= b;
    outputs(225) <= not b;
    outputs(226) <= not a or b;
    outputs(227) <= not (a xor b);
    outputs(228) <= b and not a;
    outputs(229) <= not a or b;
    outputs(230) <= not b;
    outputs(231) <= not (a or b);
    outputs(232) <= b;
    outputs(233) <= a and b;
    outputs(234) <= not (a and b);
    outputs(235) <= a and b;
    outputs(236) <= not (a xor b);
    outputs(237) <= not a or b;
    outputs(238) <= a and not b;
    outputs(239) <= b;
    outputs(240) <= not b;
    outputs(241) <= not (a or b);
    outputs(242) <= b;
    outputs(243) <= not (a xor b);
    outputs(244) <= not b;
    outputs(245) <= a and b;
    outputs(246) <= not a;
    outputs(247) <= a xor b;
    outputs(248) <= b;
    outputs(249) <= not b;
    outputs(250) <= b and not a;
    outputs(251) <= not b;
    outputs(252) <= a;
    outputs(253) <= b;
    outputs(254) <= not a;
    outputs(255) <= a;
    outputs(256) <= not b;
    outputs(257) <= a or b;
    outputs(258) <= a;
    outputs(259) <= b;
    outputs(260) <= not a;
    outputs(261) <= a;
    outputs(262) <= b;
    outputs(263) <= not (a xor b);
    outputs(264) <= not b or a;
    outputs(265) <= b;
    outputs(266) <= not (a or b);
    outputs(267) <= not (a xor b);
    outputs(268) <= b;
    outputs(269) <= a and not b;
    outputs(270) <= not a;
    outputs(271) <= not (a xor b);
    outputs(272) <= b;
    outputs(273) <= b and not a;
    outputs(274) <= not b;
    outputs(275) <= not b;
    outputs(276) <= a;
    outputs(277) <= a or b;
    outputs(278) <= a xor b;
    outputs(279) <= not b;
    outputs(280) <= not a;
    outputs(281) <= not b;
    outputs(282) <= not (a or b);
    outputs(283) <= not (a xor b);
    outputs(284) <= a xor b;
    outputs(285) <= a xor b;
    outputs(286) <= a;
    outputs(287) <= not a;
    outputs(288) <= not b;
    outputs(289) <= a xor b;
    outputs(290) <= b;
    outputs(291) <= b;
    outputs(292) <= not (a xor b);
    outputs(293) <= b and not a;
    outputs(294) <= b;
    outputs(295) <= a;
    outputs(296) <= not (a and b);
    outputs(297) <= a;
    outputs(298) <= not b;
    outputs(299) <= not (a and b);
    outputs(300) <= not a or b;
    outputs(301) <= a xor b;
    outputs(302) <= not b;
    outputs(303) <= not a;
    outputs(304) <= not a or b;
    outputs(305) <= not (a xor b);
    outputs(306) <= not (a and b);
    outputs(307) <= not a;
    outputs(308) <= a;
    outputs(309) <= not a;
    outputs(310) <= not b;
    outputs(311) <= not (a xor b);
    outputs(312) <= not a;
    outputs(313) <= not a;
    outputs(314) <= not a;
    outputs(315) <= not b;
    outputs(316) <= not b;
    outputs(317) <= a xor b;
    outputs(318) <= not a;
    outputs(319) <= not (a or b);
    outputs(320) <= a xor b;
    outputs(321) <= not b;
    outputs(322) <= a and b;
    outputs(323) <= not b;
    outputs(324) <= a;
    outputs(325) <= not a;
    outputs(326) <= b and not a;
    outputs(327) <= not b;
    outputs(328) <= not (a or b);
    outputs(329) <= not b;
    outputs(330) <= not b;
    outputs(331) <= a;
    outputs(332) <= not b;
    outputs(333) <= a and not b;
    outputs(334) <= a xor b;
    outputs(335) <= not a or b;
    outputs(336) <= b and not a;
    outputs(337) <= a xor b;
    outputs(338) <= b;
    outputs(339) <= not (a or b);
    outputs(340) <= not a;
    outputs(341) <= not b;
    outputs(342) <= not a;
    outputs(343) <= a and b;
    outputs(344) <= not (a or b);
    outputs(345) <= a;
    outputs(346) <= b;
    outputs(347) <= not b;
    outputs(348) <= a xor b;
    outputs(349) <= not b or a;
    outputs(350) <= not b;
    outputs(351) <= b and not a;
    outputs(352) <= not a or b;
    outputs(353) <= a xor b;
    outputs(354) <= a xor b;
    outputs(355) <= not b;
    outputs(356) <= a;
    outputs(357) <= a xor b;
    outputs(358) <= a xor b;
    outputs(359) <= not a;
    outputs(360) <= not (a or b);
    outputs(361) <= not (a or b);
    outputs(362) <= a and not b;
    outputs(363) <= a and not b;
    outputs(364) <= not b;
    outputs(365) <= not b;
    outputs(366) <= not b;
    outputs(367) <= not b;
    outputs(368) <= not b;
    outputs(369) <= b;
    outputs(370) <= a and not b;
    outputs(371) <= b;
    outputs(372) <= a and b;
    outputs(373) <= not b;
    outputs(374) <= not b;
    outputs(375) <= a xor b;
    outputs(376) <= not b;
    outputs(377) <= a xor b;
    outputs(378) <= not (a or b);
    outputs(379) <= not (a xor b);
    outputs(380) <= not (a xor b);
    outputs(381) <= b and not a;
    outputs(382) <= b;
    outputs(383) <= a xor b;
    outputs(384) <= not (a or b);
    outputs(385) <= not a or b;
    outputs(386) <= b;
    outputs(387) <= a xor b;
    outputs(388) <= a xor b;
    outputs(389) <= a;
    outputs(390) <= a or b;
    outputs(391) <= a;
    outputs(392) <= not a;
    outputs(393) <= a;
    outputs(394) <= a;
    outputs(395) <= a;
    outputs(396) <= not b;
    outputs(397) <= a xor b;
    outputs(398) <= not (a xor b);
    outputs(399) <= not b;
    outputs(400) <= a and not b;
    outputs(401) <= b and not a;
    outputs(402) <= b;
    outputs(403) <= not (a xor b);
    outputs(404) <= not a;
    outputs(405) <= a or b;
    outputs(406) <= not b;
    outputs(407) <= not a or b;
    outputs(408) <= a;
    outputs(409) <= not b;
    outputs(410) <= b;
    outputs(411) <= not b;
    outputs(412) <= a;
    outputs(413) <= a;
    outputs(414) <= not (a xor b);
    outputs(415) <= b;
    outputs(416) <= not a;
    outputs(417) <= a xor b;
    outputs(418) <= a xor b;
    outputs(419) <= not (a or b);
    outputs(420) <= b;
    outputs(421) <= a xor b;
    outputs(422) <= b;
    outputs(423) <= b;
    outputs(424) <= not b;
    outputs(425) <= not a;
    outputs(426) <= b;
    outputs(427) <= not a;
    outputs(428) <= a;
    outputs(429) <= a;
    outputs(430) <= a;
    outputs(431) <= not a;
    outputs(432) <= a;
    outputs(433) <= not b;
    outputs(434) <= not (a or b);
    outputs(435) <= not b;
    outputs(436) <= a xor b;
    outputs(437) <= b;
    outputs(438) <= b;
    outputs(439) <= a;
    outputs(440) <= b;
    outputs(441) <= not (a and b);
    outputs(442) <= not a;
    outputs(443) <= not (a xor b);
    outputs(444) <= not a;
    outputs(445) <= not (a xor b);
    outputs(446) <= a and b;
    outputs(447) <= b;
    outputs(448) <= a;
    outputs(449) <= not (a xor b);
    outputs(450) <= not b;
    outputs(451) <= a and b;
    outputs(452) <= a;
    outputs(453) <= b;
    outputs(454) <= not a;
    outputs(455) <= not a;
    outputs(456) <= b;
    outputs(457) <= not a or b;
    outputs(458) <= not b;
    outputs(459) <= not b;
    outputs(460) <= a and not b;
    outputs(461) <= a;
    outputs(462) <= not a or b;
    outputs(463) <= not (a or b);
    outputs(464) <= not (a or b);
    outputs(465) <= not (a xor b);
    outputs(466) <= not b or a;
    outputs(467) <= not (a xor b);
    outputs(468) <= b;
    outputs(469) <= a;
    outputs(470) <= not a;
    outputs(471) <= a and b;
    outputs(472) <= a;
    outputs(473) <= a xor b;
    outputs(474) <= not a;
    outputs(475) <= not (a or b);
    outputs(476) <= not b or a;
    outputs(477) <= b and not a;
    outputs(478) <= a;
    outputs(479) <= a and b;
    outputs(480) <= not b;
    outputs(481) <= a;
    outputs(482) <= not a or b;
    outputs(483) <= not (a xor b);
    outputs(484) <= b;
    outputs(485) <= b;
    outputs(486) <= a and b;
    outputs(487) <= a xor b;
    outputs(488) <= not a;
    outputs(489) <= not (a and b);
    outputs(490) <= b;
    outputs(491) <= not (a and b);
    outputs(492) <= a;
    outputs(493) <= a;
    outputs(494) <= a and not b;
    outputs(495) <= a xor b;
    outputs(496) <= not (a xor b);
    outputs(497) <= b;
    outputs(498) <= a and b;
    outputs(499) <= not b;
    outputs(500) <= not b;
    outputs(501) <= a and b;
    outputs(502) <= not b;
    outputs(503) <= a;
    outputs(504) <= a and not b;
    outputs(505) <= b;
    outputs(506) <= a;
    outputs(507) <= b and not a;
    outputs(508) <= not (a or b);
    outputs(509) <= b;
    outputs(510) <= a;
    outputs(511) <= b;
    outputs(512) <= a and not b;
    outputs(513) <= a or b;
    outputs(514) <= a;
    outputs(515) <= a xor b;
    outputs(516) <= not (a xor b);
    outputs(517) <= a;
    outputs(518) <= not (a xor b);
    outputs(519) <= not b;
    outputs(520) <= b;
    outputs(521) <= b;
    outputs(522) <= b;
    outputs(523) <= not a or b;
    outputs(524) <= not (a xor b);
    outputs(525) <= not (a or b);
    outputs(526) <= a xor b;
    outputs(527) <= not a;
    outputs(528) <= a;
    outputs(529) <= not a;
    outputs(530) <= b;
    outputs(531) <= not b;
    outputs(532) <= not (a xor b);
    outputs(533) <= a or b;
    outputs(534) <= b;
    outputs(535) <= b;
    outputs(536) <= a;
    outputs(537) <= not b;
    outputs(538) <= a xor b;
    outputs(539) <= not b;
    outputs(540) <= not (a xor b);
    outputs(541) <= not (a and b);
    outputs(542) <= a;
    outputs(543) <= a;
    outputs(544) <= not (a xor b);
    outputs(545) <= a;
    outputs(546) <= not (a and b);
    outputs(547) <= not b or a;
    outputs(548) <= a and not b;
    outputs(549) <= not a;
    outputs(550) <= b;
    outputs(551) <= a and b;
    outputs(552) <= b;
    outputs(553) <= b;
    outputs(554) <= not (a xor b);
    outputs(555) <= b;
    outputs(556) <= not b;
    outputs(557) <= a;
    outputs(558) <= not b;
    outputs(559) <= not b;
    outputs(560) <= a and b;
    outputs(561) <= a and b;
    outputs(562) <= not (a xor b);
    outputs(563) <= a;
    outputs(564) <= a or b;
    outputs(565) <= a;
    outputs(566) <= a and not b;
    outputs(567) <= a and not b;
    outputs(568) <= a xor b;
    outputs(569) <= not (a and b);
    outputs(570) <= b;
    outputs(571) <= a xor b;
    outputs(572) <= not b;
    outputs(573) <= b;
    outputs(574) <= not b;
    outputs(575) <= a;
    outputs(576) <= not b;
    outputs(577) <= a xor b;
    outputs(578) <= not a;
    outputs(579) <= not (a xor b);
    outputs(580) <= not b or a;
    outputs(581) <= not b;
    outputs(582) <= not (a xor b);
    outputs(583) <= not a;
    outputs(584) <= not (a xor b);
    outputs(585) <= not a or b;
    outputs(586) <= not b;
    outputs(587) <= a or b;
    outputs(588) <= not (a xor b);
    outputs(589) <= b;
    outputs(590) <= not (a xor b);
    outputs(591) <= not (a or b);
    outputs(592) <= a and not b;
    outputs(593) <= b and not a;
    outputs(594) <= a and b;
    outputs(595) <= not b;
    outputs(596) <= a;
    outputs(597) <= a;
    outputs(598) <= not (a xor b);
    outputs(599) <= a;
    outputs(600) <= not (a and b);
    outputs(601) <= not (a xor b);
    outputs(602) <= not (a xor b);
    outputs(603) <= a;
    outputs(604) <= not b;
    outputs(605) <= a xor b;
    outputs(606) <= a and not b;
    outputs(607) <= a and not b;
    outputs(608) <= a xor b;
    outputs(609) <= not a;
    outputs(610) <= a and not b;
    outputs(611) <= not a;
    outputs(612) <= not (a xor b);
    outputs(613) <= not (a and b);
    outputs(614) <= not (a xor b);
    outputs(615) <= not b or a;
    outputs(616) <= not a;
    outputs(617) <= not (a or b);
    outputs(618) <= a;
    outputs(619) <= a xor b;
    outputs(620) <= a;
    outputs(621) <= not (a xor b);
    outputs(622) <= a and b;
    outputs(623) <= a and b;
    outputs(624) <= not a;
    outputs(625) <= b;
    outputs(626) <= not (a xor b);
    outputs(627) <= a;
    outputs(628) <= a and b;
    outputs(629) <= b;
    outputs(630) <= not (a xor b);
    outputs(631) <= not b;
    outputs(632) <= not (a xor b);
    outputs(633) <= not (a and b);
    outputs(634) <= not b;
    outputs(635) <= a xor b;
    outputs(636) <= a or b;
    outputs(637) <= b;
    outputs(638) <= not (a xor b);
    outputs(639) <= not b;
    outputs(640) <= a;
    outputs(641) <= not (a xor b);
    outputs(642) <= not b;
    outputs(643) <= not (a or b);
    outputs(644) <= not a;
    outputs(645) <= b;
    outputs(646) <= a and not b;
    outputs(647) <= b;
    outputs(648) <= a;
    outputs(649) <= a;
    outputs(650) <= a xor b;
    outputs(651) <= not (a xor b);
    outputs(652) <= not (a xor b);
    outputs(653) <= not (a or b);
    outputs(654) <= not b or a;
    outputs(655) <= a and not b;
    outputs(656) <= not b;
    outputs(657) <= a;
    outputs(658) <= a;
    outputs(659) <= not (a or b);
    outputs(660) <= a xor b;
    outputs(661) <= a xor b;
    outputs(662) <= not a;
    outputs(663) <= not a;
    outputs(664) <= not (a and b);
    outputs(665) <= b and not a;
    outputs(666) <= b;
    outputs(667) <= not a;
    outputs(668) <= not b;
    outputs(669) <= a xor b;
    outputs(670) <= a and not b;
    outputs(671) <= not b;
    outputs(672) <= a xor b;
    outputs(673) <= not (a xor b);
    outputs(674) <= a;
    outputs(675) <= a and not b;
    outputs(676) <= a xor b;
    outputs(677) <= a;
    outputs(678) <= a and not b;
    outputs(679) <= a xor b;
    outputs(680) <= b;
    outputs(681) <= not a;
    outputs(682) <= a xor b;
    outputs(683) <= a xor b;
    outputs(684) <= not a;
    outputs(685) <= a and not b;
    outputs(686) <= not (a or b);
    outputs(687) <= b;
    outputs(688) <= not (a xor b);
    outputs(689) <= not b;
    outputs(690) <= not (a or b);
    outputs(691) <= not (a or b);
    outputs(692) <= a or b;
    outputs(693) <= not (a or b);
    outputs(694) <= 1'b0;
    outputs(695) <= b;
    outputs(696) <= a and not b;
    outputs(697) <= not a;
    outputs(698) <= a xor b;
    outputs(699) <= not (a xor b);
    outputs(700) <= not (a or b);
    outputs(701) <= a;
    outputs(702) <= not b;
    outputs(703) <= b;
    outputs(704) <= not (a or b);
    outputs(705) <= a;
    outputs(706) <= not a;
    outputs(707) <= not b;
    outputs(708) <= b;
    outputs(709) <= not (a or b);
    outputs(710) <= a xor b;
    outputs(711) <= a and b;
    outputs(712) <= a;
    outputs(713) <= a xor b;
    outputs(714) <= not (a or b);
    outputs(715) <= b and not a;
    outputs(716) <= not (a and b);
    outputs(717) <= a;
    outputs(718) <= not a;
    outputs(719) <= not a;
    outputs(720) <= a and b;
    outputs(721) <= not b;
    outputs(722) <= b;
    outputs(723) <= not a;
    outputs(724) <= not a;
    outputs(725) <= a;
    outputs(726) <= b and not a;
    outputs(727) <= a and not b;
    outputs(728) <= not (a xor b);
    outputs(729) <= not (a or b);
    outputs(730) <= not a;
    outputs(731) <= a and b;
    outputs(732) <= a xor b;
    outputs(733) <= not a;
    outputs(734) <= not a or b;
    outputs(735) <= a xor b;
    outputs(736) <= a;
    outputs(737) <= a xor b;
    outputs(738) <= not a;
    outputs(739) <= a xor b;
    outputs(740) <= not (a xor b);
    outputs(741) <= not (a xor b);
    outputs(742) <= not b;
    outputs(743) <= not a;
    outputs(744) <= b and not a;
    outputs(745) <= not (a or b);
    outputs(746) <= a;
    outputs(747) <= a;
    outputs(748) <= not b;
    outputs(749) <= not a;
    outputs(750) <= not (a or b);
    outputs(751) <= a xor b;
    outputs(752) <= not a;
    outputs(753) <= not b;
    outputs(754) <= not (a xor b);
    outputs(755) <= not a;
    outputs(756) <= not b or a;
    outputs(757) <= not b;
    outputs(758) <= not (a or b);
    outputs(759) <= b;
    outputs(760) <= a xor b;
    outputs(761) <= b and not a;
    outputs(762) <= not b or a;
    outputs(763) <= a xor b;
    outputs(764) <= b;
    outputs(765) <= b;
    outputs(766) <= a and b;
    outputs(767) <= not (a xor b);
    outputs(768) <= a and b;
    outputs(769) <= a xor b;
    outputs(770) <= not (a or b);
    outputs(771) <= not a;
    outputs(772) <= not a;
    outputs(773) <= not b;
    outputs(774) <= b and not a;
    outputs(775) <= b;
    outputs(776) <= not b;
    outputs(777) <= not (a and b);
    outputs(778) <= not b or a;
    outputs(779) <= not (a and b);
    outputs(780) <= a and not b;
    outputs(781) <= not a;
    outputs(782) <= not b;
    outputs(783) <= not (a xor b);
    outputs(784) <= not b;
    outputs(785) <= not a;
    outputs(786) <= b and not a;
    outputs(787) <= not (a xor b);
    outputs(788) <= not a;
    outputs(789) <= a and not b;
    outputs(790) <= not (a xor b);
    outputs(791) <= b;
    outputs(792) <= b;
    outputs(793) <= a;
    outputs(794) <= not (a xor b);
    outputs(795) <= not (a xor b);
    outputs(796) <= not a;
    outputs(797) <= a and b;
    outputs(798) <= not a;
    outputs(799) <= not a;
    outputs(800) <= a or b;
    outputs(801) <= a xor b;
    outputs(802) <= a xor b;
    outputs(803) <= a or b;
    outputs(804) <= not a;
    outputs(805) <= a and not b;
    outputs(806) <= not b;
    outputs(807) <= not a;
    outputs(808) <= b;
    outputs(809) <= not (a xor b);
    outputs(810) <= not (a xor b);
    outputs(811) <= not b;
    outputs(812) <= a;
    outputs(813) <= not b;
    outputs(814) <= a;
    outputs(815) <= a or b;
    outputs(816) <= not (a or b);
    outputs(817) <= not a;
    outputs(818) <= not (a or b);
    outputs(819) <= not (a xor b);
    outputs(820) <= not b or a;
    outputs(821) <= a;
    outputs(822) <= not (a or b);
    outputs(823) <= a;
    outputs(824) <= not b;
    outputs(825) <= not (a and b);
    outputs(826) <= not b or a;
    outputs(827) <= not (a xor b);
    outputs(828) <= a;
    outputs(829) <= b;
    outputs(830) <= b and not a;
    outputs(831) <= b;
    outputs(832) <= a;
    outputs(833) <= not (a xor b);
    outputs(834) <= b and not a;
    outputs(835) <= b and not a;
    outputs(836) <= a xor b;
    outputs(837) <= b;
    outputs(838) <= a;
    outputs(839) <= not b;
    outputs(840) <= a;
    outputs(841) <= not (a and b);
    outputs(842) <= b;
    outputs(843) <= a xor b;
    outputs(844) <= not (a xor b);
    outputs(845) <= b;
    outputs(846) <= a and not b;
    outputs(847) <= b;
    outputs(848) <= a and not b;
    outputs(849) <= a;
    outputs(850) <= not a;
    outputs(851) <= not b;
    outputs(852) <= not b;
    outputs(853) <= not (a or b);
    outputs(854) <= a;
    outputs(855) <= a;
    outputs(856) <= b;
    outputs(857) <= a;
    outputs(858) <= a xor b;
    outputs(859) <= a and not b;
    outputs(860) <= not b;
    outputs(861) <= a and b;
    outputs(862) <= not (a xor b);
    outputs(863) <= not b;
    outputs(864) <= not a;
    outputs(865) <= not b;
    outputs(866) <= not (a xor b);
    outputs(867) <= not a;
    outputs(868) <= not b;
    outputs(869) <= not a or b;
    outputs(870) <= not b;
    outputs(871) <= not b;
    outputs(872) <= not (a and b);
    outputs(873) <= not (a xor b);
    outputs(874) <= a xor b;
    outputs(875) <= a;
    outputs(876) <= not (a xor b);
    outputs(877) <= not b;
    outputs(878) <= not a;
    outputs(879) <= a xor b;
    outputs(880) <= a;
    outputs(881) <= not (a and b);
    outputs(882) <= b;
    outputs(883) <= not a;
    outputs(884) <= b;
    outputs(885) <= not (a xor b);
    outputs(886) <= b and not a;
    outputs(887) <= not a;
    outputs(888) <= not (a or b);
    outputs(889) <= b and not a;
    outputs(890) <= a and b;
    outputs(891) <= a xor b;
    outputs(892) <= a or b;
    outputs(893) <= not a or b;
    outputs(894) <= a;
    outputs(895) <= not (a xor b);
    outputs(896) <= not a;
    outputs(897) <= a and b;
    outputs(898) <= not (a xor b);
    outputs(899) <= b and not a;
    outputs(900) <= a and not b;
    outputs(901) <= a and not b;
    outputs(902) <= a and b;
    outputs(903) <= not a;
    outputs(904) <= not a or b;
    outputs(905) <= a;
    outputs(906) <= a;
    outputs(907) <= not b;
    outputs(908) <= a xor b;
    outputs(909) <= b;
    outputs(910) <= not b;
    outputs(911) <= not (a xor b);
    outputs(912) <= a xor b;
    outputs(913) <= b and not a;
    outputs(914) <= not a;
    outputs(915) <= a xor b;
    outputs(916) <= a;
    outputs(917) <= a;
    outputs(918) <= b and not a;
    outputs(919) <= not a or b;
    outputs(920) <= a xor b;
    outputs(921) <= b;
    outputs(922) <= not (a and b);
    outputs(923) <= not a;
    outputs(924) <= not a;
    outputs(925) <= not b;
    outputs(926) <= b;
    outputs(927) <= not (a or b);
    outputs(928) <= not (a or b);
    outputs(929) <= b;
    outputs(930) <= not (a xor b);
    outputs(931) <= a;
    outputs(932) <= b;
    outputs(933) <= a xor b;
    outputs(934) <= a and b;
    outputs(935) <= b and not a;
    outputs(936) <= not a;
    outputs(937) <= b;
    outputs(938) <= a xor b;
    outputs(939) <= not (a and b);
    outputs(940) <= b;
    outputs(941) <= not b;
    outputs(942) <= a xor b;
    outputs(943) <= a xor b;
    outputs(944) <= b and not a;
    outputs(945) <= a;
    outputs(946) <= b and not a;
    outputs(947) <= not a;
    outputs(948) <= a;
    outputs(949) <= not b or a;
    outputs(950) <= a xor b;
    outputs(951) <= not a;
    outputs(952) <= not a;
    outputs(953) <= not b or a;
    outputs(954) <= not (a xor b);
    outputs(955) <= a;
    outputs(956) <= a and b;
    outputs(957) <= not (a and b);
    outputs(958) <= not a;
    outputs(959) <= not b or a;
    outputs(960) <= a and not b;
    outputs(961) <= not a;
    outputs(962) <= not a or b;
    outputs(963) <= not a;
    outputs(964) <= b and not a;
    outputs(965) <= b;
    outputs(966) <= a or b;
    outputs(967) <= b;
    outputs(968) <= not b;
    outputs(969) <= a or b;
    outputs(970) <= a;
    outputs(971) <= not a;
    outputs(972) <= a and not b;
    outputs(973) <= not a or b;
    outputs(974) <= b and not a;
    outputs(975) <= a;
    outputs(976) <= b;
    outputs(977) <= a;
    outputs(978) <= not b or a;
    outputs(979) <= a;
    outputs(980) <= a and b;
    outputs(981) <= not (a xor b);
    outputs(982) <= b;
    outputs(983) <= b;
    outputs(984) <= b and not a;
    outputs(985) <= not a;
    outputs(986) <= a;
    outputs(987) <= not b or a;
    outputs(988) <= b and not a;
    outputs(989) <= not (a xor b);
    outputs(990) <= not (a xor b);
    outputs(991) <= not a;
    outputs(992) <= a or b;
    outputs(993) <= not (a and b);
    outputs(994) <= b and not a;
    outputs(995) <= not a;
    outputs(996) <= not a;
    outputs(997) <= a and b;
    outputs(998) <= b;
    outputs(999) <= a and not b;
    outputs(1000) <= not a;
    outputs(1001) <= not (a and b);
    outputs(1002) <= a and not b;
    outputs(1003) <= a;
    outputs(1004) <= not a;
    outputs(1005) <= b;
    outputs(1006) <= b;
    outputs(1007) <= not b;
    outputs(1008) <= a;
    outputs(1009) <= a and b;
    outputs(1010) <= not a;
    outputs(1011) <= not a or b;
    outputs(1012) <= not (a and b);
    outputs(1013) <= a or b;
    outputs(1014) <= not a;
    outputs(1015) <= not (a and b);
    outputs(1016) <= not (a or b);
    outputs(1017) <= not a;
    outputs(1018) <= not a;
    outputs(1019) <= a and not b;
    outputs(1020) <= not a;
    outputs(1021) <= b;
    outputs(1022) <= not b;
    outputs(1023) <= b;
    outputs(1024) <= not (a or b);
    outputs(1025) <= a xor b;
    outputs(1026) <= not (a xor b);
    outputs(1027) <= a xor b;
    outputs(1028) <= not b;
    outputs(1029) <= not b;
    outputs(1030) <= not a;
    outputs(1031) <= not (a xor b);
    outputs(1032) <= b and not a;
    outputs(1033) <= a and not b;
    outputs(1034) <= b;
    outputs(1035) <= not (a or b);
    outputs(1036) <= not (a xor b);
    outputs(1037) <= b;
    outputs(1038) <= not (a and b);
    outputs(1039) <= a xor b;
    outputs(1040) <= a;
    outputs(1041) <= not (a xor b);
    outputs(1042) <= b and not a;
    outputs(1043) <= a;
    outputs(1044) <= a xor b;
    outputs(1045) <= a;
    outputs(1046) <= a xor b;
    outputs(1047) <= not (a xor b);
    outputs(1048) <= b;
    outputs(1049) <= not (a xor b);
    outputs(1050) <= a and not b;
    outputs(1051) <= a;
    outputs(1052) <= b and not a;
    outputs(1053) <= b and not a;
    outputs(1054) <= a and b;
    outputs(1055) <= not a;
    outputs(1056) <= a xor b;
    outputs(1057) <= a;
    outputs(1058) <= a;
    outputs(1059) <= a;
    outputs(1060) <= a and b;
    outputs(1061) <= a xor b;
    outputs(1062) <= not (a xor b);
    outputs(1063) <= not a;
    outputs(1064) <= not (a or b);
    outputs(1065) <= a and b;
    outputs(1066) <= b;
    outputs(1067) <= not b;
    outputs(1068) <= b;
    outputs(1069) <= not a;
    outputs(1070) <= not b;
    outputs(1071) <= not (a xor b);
    outputs(1072) <= not (a xor b);
    outputs(1073) <= a and not b;
    outputs(1074) <= a xor b;
    outputs(1075) <= a xor b;
    outputs(1076) <= not a;
    outputs(1077) <= 1'b0;
    outputs(1078) <= not b;
    outputs(1079) <= not b;
    outputs(1080) <= not (a or b);
    outputs(1081) <= a;
    outputs(1082) <= not (a xor b);
    outputs(1083) <= a and not b;
    outputs(1084) <= a;
    outputs(1085) <= not (a xor b);
    outputs(1086) <= not b;
    outputs(1087) <= a xor b;
    outputs(1088) <= a xor b;
    outputs(1089) <= not (a xor b);
    outputs(1090) <= a and not b;
    outputs(1091) <= not b;
    outputs(1092) <= not b;
    outputs(1093) <= not (a xor b);
    outputs(1094) <= a xor b;
    outputs(1095) <= b;
    outputs(1096) <= a and b;
    outputs(1097) <= a and b;
    outputs(1098) <= not b;
    outputs(1099) <= a xor b;
    outputs(1100) <= a xor b;
    outputs(1101) <= not (a xor b);
    outputs(1102) <= a xor b;
    outputs(1103) <= a and not b;
    outputs(1104) <= not b;
    outputs(1105) <= b;
    outputs(1106) <= not (a xor b);
    outputs(1107) <= not (a xor b);
    outputs(1108) <= b;
    outputs(1109) <= a and not b;
    outputs(1110) <= not (a xor b);
    outputs(1111) <= a;
    outputs(1112) <= a and b;
    outputs(1113) <= b;
    outputs(1114) <= not a;
    outputs(1115) <= a xor b;
    outputs(1116) <= not a;
    outputs(1117) <= a and b;
    outputs(1118) <= a and not b;
    outputs(1119) <= not a;
    outputs(1120) <= b and not a;
    outputs(1121) <= a xor b;
    outputs(1122) <= not b;
    outputs(1123) <= not a;
    outputs(1124) <= not a;
    outputs(1125) <= not a;
    outputs(1126) <= a;
    outputs(1127) <= a;
    outputs(1128) <= not (a xor b);
    outputs(1129) <= a xor b;
    outputs(1130) <= not (a or b);
    outputs(1131) <= a and b;
    outputs(1132) <= not b;
    outputs(1133) <= not a;
    outputs(1134) <= a xor b;
    outputs(1135) <= b;
    outputs(1136) <= b and not a;
    outputs(1137) <= a and b;
    outputs(1138) <= not (a and b);
    outputs(1139) <= a and not b;
    outputs(1140) <= a xor b;
    outputs(1141) <= a and not b;
    outputs(1142) <= a;
    outputs(1143) <= a and not b;
    outputs(1144) <= b;
    outputs(1145) <= not (a xor b);
    outputs(1146) <= not (a xor b);
    outputs(1147) <= a and b;
    outputs(1148) <= a xor b;
    outputs(1149) <= a and b;
    outputs(1150) <= not (a or b);
    outputs(1151) <= a xor b;
    outputs(1152) <= b;
    outputs(1153) <= b and not a;
    outputs(1154) <= not a;
    outputs(1155) <= b and not a;
    outputs(1156) <= a or b;
    outputs(1157) <= not (a xor b);
    outputs(1158) <= a xor b;
    outputs(1159) <= not (a xor b);
    outputs(1160) <= b and not a;
    outputs(1161) <= not (a xor b);
    outputs(1162) <= a xor b;
    outputs(1163) <= not (a xor b);
    outputs(1164) <= not a;
    outputs(1165) <= b;
    outputs(1166) <= a and not b;
    outputs(1167) <= a xor b;
    outputs(1168) <= a xor b;
    outputs(1169) <= a xor b;
    outputs(1170) <= a xor b;
    outputs(1171) <= not (a xor b);
    outputs(1172) <= a and b;
    outputs(1173) <= not b;
    outputs(1174) <= a xor b;
    outputs(1175) <= not (a and b);
    outputs(1176) <= a xor b;
    outputs(1177) <= b;
    outputs(1178) <= not (a or b);
    outputs(1179) <= a;
    outputs(1180) <= a xor b;
    outputs(1181) <= not (a or b);
    outputs(1182) <= not (a xor b);
    outputs(1183) <= a and b;
    outputs(1184) <= a and b;
    outputs(1185) <= b;
    outputs(1186) <= a;
    outputs(1187) <= not b;
    outputs(1188) <= a and not b;
    outputs(1189) <= not (a or b);
    outputs(1190) <= a or b;
    outputs(1191) <= b;
    outputs(1192) <= not a;
    outputs(1193) <= not a;
    outputs(1194) <= a or b;
    outputs(1195) <= a and b;
    outputs(1196) <= not b;
    outputs(1197) <= not b;
    outputs(1198) <= b;
    outputs(1199) <= not b;
    outputs(1200) <= a xor b;
    outputs(1201) <= a xor b;
    outputs(1202) <= a and b;
    outputs(1203) <= not (a xor b);
    outputs(1204) <= not (a xor b);
    outputs(1205) <= not (a xor b);
    outputs(1206) <= a;
    outputs(1207) <= a xor b;
    outputs(1208) <= not (a or b);
    outputs(1209) <= not (a xor b);
    outputs(1210) <= not a;
    outputs(1211) <= a;
    outputs(1212) <= a and not b;
    outputs(1213) <= b and not a;
    outputs(1214) <= b;
    outputs(1215) <= not (a xor b);
    outputs(1216) <= not b;
    outputs(1217) <= b and not a;
    outputs(1218) <= a and not b;
    outputs(1219) <= a;
    outputs(1220) <= not a;
    outputs(1221) <= not b;
    outputs(1222) <= not (a or b);
    outputs(1223) <= not (a or b);
    outputs(1224) <= a xor b;
    outputs(1225) <= a xor b;
    outputs(1226) <= b;
    outputs(1227) <= b and not a;
    outputs(1228) <= a xor b;
    outputs(1229) <= not (a xor b);
    outputs(1230) <= a and b;
    outputs(1231) <= b;
    outputs(1232) <= b;
    outputs(1233) <= a or b;
    outputs(1234) <= not (a xor b);
    outputs(1235) <= not (a xor b);
    outputs(1236) <= not (a or b);
    outputs(1237) <= not (a or b);
    outputs(1238) <= b;
    outputs(1239) <= not a or b;
    outputs(1240) <= not (a xor b);
    outputs(1241) <= not b;
    outputs(1242) <= a xor b;
    outputs(1243) <= not (a xor b);
    outputs(1244) <= a and not b;
    outputs(1245) <= not b;
    outputs(1246) <= not (a xor b);
    outputs(1247) <= b and not a;
    outputs(1248) <= a xor b;
    outputs(1249) <= b;
    outputs(1250) <= b and not a;
    outputs(1251) <= a and not b;
    outputs(1252) <= not a;
    outputs(1253) <= a and not b;
    outputs(1254) <= b and not a;
    outputs(1255) <= a xor b;
    outputs(1256) <= a and b;
    outputs(1257) <= not a;
    outputs(1258) <= b and not a;
    outputs(1259) <= a;
    outputs(1260) <= a and b;
    outputs(1261) <= a xor b;
    outputs(1262) <= not b;
    outputs(1263) <= a and b;
    outputs(1264) <= a xor b;
    outputs(1265) <= not b;
    outputs(1266) <= not a;
    outputs(1267) <= not (a xor b);
    outputs(1268) <= a;
    outputs(1269) <= not b;
    outputs(1270) <= not (a or b);
    outputs(1271) <= a and not b;
    outputs(1272) <= b;
    outputs(1273) <= not (a xor b);
    outputs(1274) <= b;
    outputs(1275) <= not (a xor b);
    outputs(1276) <= not (a or b);
    outputs(1277) <= b;
    outputs(1278) <= b;
    outputs(1279) <= not a or b;
    outputs(1280) <= not a;
    outputs(1281) <= not b;
    outputs(1282) <= a;
    outputs(1283) <= not (a xor b);
    outputs(1284) <= not (a or b);
    outputs(1285) <= a xor b;
    outputs(1286) <= not (a or b);
    outputs(1287) <= not (a xor b);
    outputs(1288) <= not (a or b);
    outputs(1289) <= a xor b;
    outputs(1290) <= b;
    outputs(1291) <= not a;
    outputs(1292) <= a or b;
    outputs(1293) <= not (a or b);
    outputs(1294) <= a xor b;
    outputs(1295) <= a and not b;
    outputs(1296) <= not (a or b);
    outputs(1297) <= a and b;
    outputs(1298) <= not (a xor b);
    outputs(1299) <= not (a or b);
    outputs(1300) <= a xor b;
    outputs(1301) <= not (a and b);
    outputs(1302) <= not (a or b);
    outputs(1303) <= not (a xor b);
    outputs(1304) <= not a;
    outputs(1305) <= a and b;
    outputs(1306) <= a;
    outputs(1307) <= a and b;
    outputs(1308) <= not a;
    outputs(1309) <= a;
    outputs(1310) <= not (a or b);
    outputs(1311) <= a and b;
    outputs(1312) <= a or b;
    outputs(1313) <= a or b;
    outputs(1314) <= a and b;
    outputs(1315) <= not (a or b);
    outputs(1316) <= not (a xor b);
    outputs(1317) <= not b;
    outputs(1318) <= a and b;
    outputs(1319) <= not a;
    outputs(1320) <= a and b;
    outputs(1321) <= not (a or b);
    outputs(1322) <= not (a or b);
    outputs(1323) <= not (a or b);
    outputs(1324) <= not (a or b);
    outputs(1325) <= a and not b;
    outputs(1326) <= a and b;
    outputs(1327) <= not b;
    outputs(1328) <= not (a or b);
    outputs(1329) <= a and not b;
    outputs(1330) <= not b;
    outputs(1331) <= a xor b;
    outputs(1332) <= b and not a;
    outputs(1333) <= not b;
    outputs(1334) <= not b;
    outputs(1335) <= not (a xor b);
    outputs(1336) <= a xor b;
    outputs(1337) <= b and not a;
    outputs(1338) <= not a;
    outputs(1339) <= a and not b;
    outputs(1340) <= b;
    outputs(1341) <= b and not a;
    outputs(1342) <= a and not b;
    outputs(1343) <= b;
    outputs(1344) <= not b;
    outputs(1345) <= a xor b;
    outputs(1346) <= a xor b;
    outputs(1347) <= not (a xor b);
    outputs(1348) <= b;
    outputs(1349) <= not (a xor b);
    outputs(1350) <= not a;
    outputs(1351) <= not a;
    outputs(1352) <= not (a xor b);
    outputs(1353) <= a xor b;
    outputs(1354) <= not (a or b);
    outputs(1355) <= a;
    outputs(1356) <= a and not b;
    outputs(1357) <= a and b;
    outputs(1358) <= not (a or b);
    outputs(1359) <= not a;
    outputs(1360) <= not b;
    outputs(1361) <= not b;
    outputs(1362) <= not (a xor b);
    outputs(1363) <= not b or a;
    outputs(1364) <= not (a xor b);
    outputs(1365) <= a xor b;
    outputs(1366) <= a xor b;
    outputs(1367) <= b and not a;
    outputs(1368) <= not (a xor b);
    outputs(1369) <= not (a xor b);
    outputs(1370) <= not a;
    outputs(1371) <= a and not b;
    outputs(1372) <= not (a xor b);
    outputs(1373) <= a xor b;
    outputs(1374) <= a xor b;
    outputs(1375) <= not (a xor b);
    outputs(1376) <= not b;
    outputs(1377) <= not a;
    outputs(1378) <= a and not b;
    outputs(1379) <= not (a xor b);
    outputs(1380) <= b;
    outputs(1381) <= a xor b;
    outputs(1382) <= a and not b;
    outputs(1383) <= not (a xor b);
    outputs(1384) <= a;
    outputs(1385) <= a;
    outputs(1386) <= a;
    outputs(1387) <= a xor b;
    outputs(1388) <= not b;
    outputs(1389) <= a;
    outputs(1390) <= not (a or b);
    outputs(1391) <= not (a xor b);
    outputs(1392) <= not (a or b);
    outputs(1393) <= a;
    outputs(1394) <= a and not b;
    outputs(1395) <= a and not b;
    outputs(1396) <= b and not a;
    outputs(1397) <= b and not a;
    outputs(1398) <= a and b;
    outputs(1399) <= not (a xor b);
    outputs(1400) <= a xor b;
    outputs(1401) <= a and not b;
    outputs(1402) <= not a;
    outputs(1403) <= not b;
    outputs(1404) <= not a;
    outputs(1405) <= not (a xor b);
    outputs(1406) <= a and not b;
    outputs(1407) <= not (a xor b);
    outputs(1408) <= b and not a;
    outputs(1409) <= b;
    outputs(1410) <= a xor b;
    outputs(1411) <= b and not a;
    outputs(1412) <= not (a or b);
    outputs(1413) <= not (a xor b);
    outputs(1414) <= not b;
    outputs(1415) <= not (a xor b);
    outputs(1416) <= a;
    outputs(1417) <= a and not b;
    outputs(1418) <= a xor b;
    outputs(1419) <= a xor b;
    outputs(1420) <= not a;
    outputs(1421) <= not a;
    outputs(1422) <= not (a or b);
    outputs(1423) <= not (a xor b);
    outputs(1424) <= not (a and b);
    outputs(1425) <= not b;
    outputs(1426) <= 1'b0;
    outputs(1427) <= a;
    outputs(1428) <= not (a xor b);
    outputs(1429) <= not (a or b);
    outputs(1430) <= b;
    outputs(1431) <= b;
    outputs(1432) <= a;
    outputs(1433) <= b and not a;
    outputs(1434) <= a xor b;
    outputs(1435) <= not b;
    outputs(1436) <= a xor b;
    outputs(1437) <= a and b;
    outputs(1438) <= a and b;
    outputs(1439) <= not a;
    outputs(1440) <= a and not b;
    outputs(1441) <= a xor b;
    outputs(1442) <= not a;
    outputs(1443) <= not (a xor b);
    outputs(1444) <= a;
    outputs(1445) <= b;
    outputs(1446) <= a xor b;
    outputs(1447) <= not (a xor b);
    outputs(1448) <= b;
    outputs(1449) <= b;
    outputs(1450) <= a xor b;
    outputs(1451) <= not (a xor b);
    outputs(1452) <= not b;
    outputs(1453) <= b and not a;
    outputs(1454) <= a xor b;
    outputs(1455) <= not (a xor b);
    outputs(1456) <= not b;
    outputs(1457) <= 1'b0;
    outputs(1458) <= not (a or b);
    outputs(1459) <= a;
    outputs(1460) <= not (a or b);
    outputs(1461) <= not b;
    outputs(1462) <= a xor b;
    outputs(1463) <= b and not a;
    outputs(1464) <= not a;
    outputs(1465) <= not (a or b);
    outputs(1466) <= not (a xor b);
    outputs(1467) <= a xor b;
    outputs(1468) <= a and b;
    outputs(1469) <= b and not a;
    outputs(1470) <= not (a xor b);
    outputs(1471) <= a and not b;
    outputs(1472) <= a;
    outputs(1473) <= not (a xor b);
    outputs(1474) <= a xor b;
    outputs(1475) <= not b;
    outputs(1476) <= a;
    outputs(1477) <= not (a xor b);
    outputs(1478) <= not (a or b);
    outputs(1479) <= not (a xor b);
    outputs(1480) <= not a;
    outputs(1481) <= a and not b;
    outputs(1482) <= a and not b;
    outputs(1483) <= not (a or b);
    outputs(1484) <= not (a xor b);
    outputs(1485) <= a and b;
    outputs(1486) <= not b or a;
    outputs(1487) <= a xor b;
    outputs(1488) <= not a;
    outputs(1489) <= a xor b;
    outputs(1490) <= a and not b;
    outputs(1491) <= b;
    outputs(1492) <= not b or a;
    outputs(1493) <= not b;
    outputs(1494) <= not a;
    outputs(1495) <= a xor b;
    outputs(1496) <= a and not b;
    outputs(1497) <= b;
    outputs(1498) <= not b;
    outputs(1499) <= a and b;
    outputs(1500) <= b;
    outputs(1501) <= not a or b;
    outputs(1502) <= a xor b;
    outputs(1503) <= b;
    outputs(1504) <= b and not a;
    outputs(1505) <= b;
    outputs(1506) <= a;
    outputs(1507) <= not b;
    outputs(1508) <= a and not b;
    outputs(1509) <= a and b;
    outputs(1510) <= b and not a;
    outputs(1511) <= not b;
    outputs(1512) <= not (a or b);
    outputs(1513) <= not (a or b);
    outputs(1514) <= not (a xor b);
    outputs(1515) <= not (a xor b);
    outputs(1516) <= b and not a;
    outputs(1517) <= not (a xor b);
    outputs(1518) <= a and not b;
    outputs(1519) <= not b or a;
    outputs(1520) <= a xor b;
    outputs(1521) <= not (a xor b);
    outputs(1522) <= b and not a;
    outputs(1523) <= b;
    outputs(1524) <= not a;
    outputs(1525) <= not (a xor b);
    outputs(1526) <= a and not b;
    outputs(1527) <= b and not a;
    outputs(1528) <= not (a xor b);
    outputs(1529) <= a xor b;
    outputs(1530) <= a;
    outputs(1531) <= a and b;
    outputs(1532) <= not b;
    outputs(1533) <= a and b;
    outputs(1534) <= b and not a;
    outputs(1535) <= not b;
    outputs(1536) <= a and not b;
    outputs(1537) <= not (a or b);
    outputs(1538) <= not a;
    outputs(1539) <= not (a xor b);
    outputs(1540) <= a and b;
    outputs(1541) <= not (a xor b);
    outputs(1542) <= not (a or b);
    outputs(1543) <= a and not b;
    outputs(1544) <= a xor b;
    outputs(1545) <= a xor b;
    outputs(1546) <= not b;
    outputs(1547) <= not (a xor b);
    outputs(1548) <= a;
    outputs(1549) <= b;
    outputs(1550) <= not a;
    outputs(1551) <= a and not b;
    outputs(1552) <= not (a xor b);
    outputs(1553) <= not (a or b);
    outputs(1554) <= a and b;
    outputs(1555) <= not b;
    outputs(1556) <= a xor b;
    outputs(1557) <= a or b;
    outputs(1558) <= a xor b;
    outputs(1559) <= a and b;
    outputs(1560) <= not (a xor b);
    outputs(1561) <= a and b;
    outputs(1562) <= b and not a;
    outputs(1563) <= a xor b;
    outputs(1564) <= not b;
    outputs(1565) <= b and not a;
    outputs(1566) <= a and not b;
    outputs(1567) <= a xor b;
    outputs(1568) <= not a;
    outputs(1569) <= a xor b;
    outputs(1570) <= a and not b;
    outputs(1571) <= not b;
    outputs(1572) <= not (a or b);
    outputs(1573) <= b and not a;
    outputs(1574) <= not (a xor b);
    outputs(1575) <= a and not b;
    outputs(1576) <= not (a or b);
    outputs(1577) <= not b;
    outputs(1578) <= b and not a;
    outputs(1579) <= a xor b;
    outputs(1580) <= not a or b;
    outputs(1581) <= b;
    outputs(1582) <= not b;
    outputs(1583) <= not b;
    outputs(1584) <= b;
    outputs(1585) <= a and not b;
    outputs(1586) <= b and not a;
    outputs(1587) <= a and not b;
    outputs(1588) <= not (a or b);
    outputs(1589) <= a;
    outputs(1590) <= a xor b;
    outputs(1591) <= not (a xor b);
    outputs(1592) <= a and not b;
    outputs(1593) <= not (a or b);
    outputs(1594) <= a;
    outputs(1595) <= not (a xor b);
    outputs(1596) <= not b;
    outputs(1597) <= b;
    outputs(1598) <= a;
    outputs(1599) <= not (a xor b);
    outputs(1600) <= a;
    outputs(1601) <= b;
    outputs(1602) <= a xor b;
    outputs(1603) <= a and b;
    outputs(1604) <= a;
    outputs(1605) <= a and not b;
    outputs(1606) <= not (a xor b);
    outputs(1607) <= a and b;
    outputs(1608) <= b;
    outputs(1609) <= not a;
    outputs(1610) <= a and not b;
    outputs(1611) <= b;
    outputs(1612) <= a;
    outputs(1613) <= a and b;
    outputs(1614) <= b and not a;
    outputs(1615) <= not (a or b);
    outputs(1616) <= not (a or b);
    outputs(1617) <= b;
    outputs(1618) <= not (a xor b);
    outputs(1619) <= a xor b;
    outputs(1620) <= a xor b;
    outputs(1621) <= not a;
    outputs(1622) <= not (a xor b);
    outputs(1623) <= a and not b;
    outputs(1624) <= a;
    outputs(1625) <= a and not b;
    outputs(1626) <= b;
    outputs(1627) <= a;
    outputs(1628) <= not (a xor b);
    outputs(1629) <= a;
    outputs(1630) <= not (a xor b);
    outputs(1631) <= not (a xor b);
    outputs(1632) <= a xor b;
    outputs(1633) <= not (a xor b);
    outputs(1634) <= not b;
    outputs(1635) <= not b;
    outputs(1636) <= not (a xor b);
    outputs(1637) <= a xor b;
    outputs(1638) <= a and b;
    outputs(1639) <= not (a xor b);
    outputs(1640) <= a xor b;
    outputs(1641) <= not b;
    outputs(1642) <= not (a xor b);
    outputs(1643) <= b;
    outputs(1644) <= not b;
    outputs(1645) <= a and not b;
    outputs(1646) <= a and not b;
    outputs(1647) <= a xor b;
    outputs(1648) <= b and not a;
    outputs(1649) <= a and not b;
    outputs(1650) <= not a or b;
    outputs(1651) <= a;
    outputs(1652) <= a xor b;
    outputs(1653) <= not (a xor b);
    outputs(1654) <= a and not b;
    outputs(1655) <= a;
    outputs(1656) <= a;
    outputs(1657) <= b and not a;
    outputs(1658) <= not b;
    outputs(1659) <= not (a xor b);
    outputs(1660) <= not b;
    outputs(1661) <= not (a or b);
    outputs(1662) <= a and not b;
    outputs(1663) <= a xor b;
    outputs(1664) <= a xor b;
    outputs(1665) <= a and not b;
    outputs(1666) <= not (a or b);
    outputs(1667) <= b and not a;
    outputs(1668) <= not (a xor b);
    outputs(1669) <= not a;
    outputs(1670) <= not (a or b);
    outputs(1671) <= a and not b;
    outputs(1672) <= a xor b;
    outputs(1673) <= not a;
    outputs(1674) <= not (a xor b);
    outputs(1675) <= not (a or b);
    outputs(1676) <= a xor b;
    outputs(1677) <= a xor b;
    outputs(1678) <= not (a xor b);
    outputs(1679) <= a xor b;
    outputs(1680) <= not (a xor b);
    outputs(1681) <= not (a xor b);
    outputs(1682) <= not a;
    outputs(1683) <= not b;
    outputs(1684) <= b;
    outputs(1685) <= a;
    outputs(1686) <= not (a xor b);
    outputs(1687) <= not (a xor b);
    outputs(1688) <= a and not b;
    outputs(1689) <= not (a xor b);
    outputs(1690) <= a;
    outputs(1691) <= not a;
    outputs(1692) <= a and b;
    outputs(1693) <= a and not b;
    outputs(1694) <= a and not b;
    outputs(1695) <= not a;
    outputs(1696) <= a and b;
    outputs(1697) <= a and not b;
    outputs(1698) <= a and b;
    outputs(1699) <= not b;
    outputs(1700) <= a;
    outputs(1701) <= a and not b;
    outputs(1702) <= not a;
    outputs(1703) <= not (a or b);
    outputs(1704) <= not (a or b);
    outputs(1705) <= not a;
    outputs(1706) <= not a;
    outputs(1707) <= a and not b;
    outputs(1708) <= not a or b;
    outputs(1709) <= a;
    outputs(1710) <= not b;
    outputs(1711) <= not (a xor b);
    outputs(1712) <= not (a xor b);
    outputs(1713) <= not (a xor b);
    outputs(1714) <= a and b;
    outputs(1715) <= a and not b;
    outputs(1716) <= not a;
    outputs(1717) <= b;
    outputs(1718) <= not a;
    outputs(1719) <= b;
    outputs(1720) <= a xor b;
    outputs(1721) <= not (a xor b);
    outputs(1722) <= not b;
    outputs(1723) <= not (a or b);
    outputs(1724) <= b and not a;
    outputs(1725) <= a xor b;
    outputs(1726) <= not a;
    outputs(1727) <= not b or a;
    outputs(1728) <= a and b;
    outputs(1729) <= b;
    outputs(1730) <= a and b;
    outputs(1731) <= b;
    outputs(1732) <= a xor b;
    outputs(1733) <= not (a or b);
    outputs(1734) <= not (a xor b);
    outputs(1735) <= a and b;
    outputs(1736) <= b;
    outputs(1737) <= not (a and b);
    outputs(1738) <= a xor b;
    outputs(1739) <= a or b;
    outputs(1740) <= b;
    outputs(1741) <= a xor b;
    outputs(1742) <= a and not b;
    outputs(1743) <= a xor b;
    outputs(1744) <= a and b;
    outputs(1745) <= not (a xor b);
    outputs(1746) <= a and b;
    outputs(1747) <= not b;
    outputs(1748) <= a xor b;
    outputs(1749) <= a;
    outputs(1750) <= a and b;
    outputs(1751) <= a xor b;
    outputs(1752) <= a and b;
    outputs(1753) <= a xor b;
    outputs(1754) <= a xor b;
    outputs(1755) <= not b;
    outputs(1756) <= a xor b;
    outputs(1757) <= a and b;
    outputs(1758) <= not b;
    outputs(1759) <= a xor b;
    outputs(1760) <= a xor b;
    outputs(1761) <= not (a xor b);
    outputs(1762) <= a;
    outputs(1763) <= a xor b;
    outputs(1764) <= a and not b;
    outputs(1765) <= a xor b;
    outputs(1766) <= a xor b;
    outputs(1767) <= a;
    outputs(1768) <= not (a or b);
    outputs(1769) <= not b;
    outputs(1770) <= not a;
    outputs(1771) <= a;
    outputs(1772) <= b;
    outputs(1773) <= a and b;
    outputs(1774) <= not (a and b);
    outputs(1775) <= a xor b;
    outputs(1776) <= a and b;
    outputs(1777) <= not (a or b);
    outputs(1778) <= b;
    outputs(1779) <= a and not b;
    outputs(1780) <= a and b;
    outputs(1781) <= not a;
    outputs(1782) <= b;
    outputs(1783) <= a and b;
    outputs(1784) <= not a;
    outputs(1785) <= not (a or b);
    outputs(1786) <= a or b;
    outputs(1787) <= b and not a;
    outputs(1788) <= a and not b;
    outputs(1789) <= not (a xor b);
    outputs(1790) <= not a or b;
    outputs(1791) <= not b;
    outputs(1792) <= a xor b;
    outputs(1793) <= a;
    outputs(1794) <= not (a xor b);
    outputs(1795) <= a;
    outputs(1796) <= b;
    outputs(1797) <= a;
    outputs(1798) <= not (a xor b);
    outputs(1799) <= b;
    outputs(1800) <= not b;
    outputs(1801) <= not (a or b);
    outputs(1802) <= not (a xor b);
    outputs(1803) <= not (a and b);
    outputs(1804) <= not b;
    outputs(1805) <= b;
    outputs(1806) <= a xor b;
    outputs(1807) <= b;
    outputs(1808) <= not b;
    outputs(1809) <= a;
    outputs(1810) <= a or b;
    outputs(1811) <= b;
    outputs(1812) <= not (a or b);
    outputs(1813) <= not (a or b);
    outputs(1814) <= b and not a;
    outputs(1815) <= a;
    outputs(1816) <= a and not b;
    outputs(1817) <= not a;
    outputs(1818) <= a;
    outputs(1819) <= b and not a;
    outputs(1820) <= not (a xor b);
    outputs(1821) <= not b;
    outputs(1822) <= not a;
    outputs(1823) <= b and not a;
    outputs(1824) <= not (a xor b);
    outputs(1825) <= not b;
    outputs(1826) <= a and b;
    outputs(1827) <= a;
    outputs(1828) <= not (a or b);
    outputs(1829) <= not b;
    outputs(1830) <= not (a xor b);
    outputs(1831) <= b and not a;
    outputs(1832) <= not (a xor b);
    outputs(1833) <= a xor b;
    outputs(1834) <= a;
    outputs(1835) <= a xor b;
    outputs(1836) <= not b;
    outputs(1837) <= b and not a;
    outputs(1838) <= a and not b;
    outputs(1839) <= a and b;
    outputs(1840) <= not a;
    outputs(1841) <= a xor b;
    outputs(1842) <= a xor b;
    outputs(1843) <= a xor b;
    outputs(1844) <= b and not a;
    outputs(1845) <= not b;
    outputs(1846) <= not a;
    outputs(1847) <= b;
    outputs(1848) <= a;
    outputs(1849) <= not (a or b);
    outputs(1850) <= a;
    outputs(1851) <= a xor b;
    outputs(1852) <= not (a or b);
    outputs(1853) <= a and not b;
    outputs(1854) <= not (a xor b);
    outputs(1855) <= not b;
    outputs(1856) <= a and not b;
    outputs(1857) <= a and not b;
    outputs(1858) <= not (a xor b);
    outputs(1859) <= not (a xor b);
    outputs(1860) <= not (a xor b);
    outputs(1861) <= not (a or b);
    outputs(1862) <= b;
    outputs(1863) <= not (a xor b);
    outputs(1864) <= a;
    outputs(1865) <= not a;
    outputs(1866) <= not a;
    outputs(1867) <= not a or b;
    outputs(1868) <= not a;
    outputs(1869) <= not (a xor b);
    outputs(1870) <= b;
    outputs(1871) <= a xor b;
    outputs(1872) <= b and not a;
    outputs(1873) <= a and b;
    outputs(1874) <= not (a or b);
    outputs(1875) <= b;
    outputs(1876) <= a and not b;
    outputs(1877) <= a and not b;
    outputs(1878) <= a and b;
    outputs(1879) <= not a;
    outputs(1880) <= a xor b;
    outputs(1881) <= a and b;
    outputs(1882) <= a xor b;
    outputs(1883) <= b and not a;
    outputs(1884) <= b and not a;
    outputs(1885) <= b and not a;
    outputs(1886) <= a and not b;
    outputs(1887) <= a xor b;
    outputs(1888) <= not (a and b);
    outputs(1889) <= a and b;
    outputs(1890) <= a xor b;
    outputs(1891) <= not (a xor b);
    outputs(1892) <= a;
    outputs(1893) <= b and not a;
    outputs(1894) <= a xor b;
    outputs(1895) <= a xor b;
    outputs(1896) <= not a;
    outputs(1897) <= a xor b;
    outputs(1898) <= a xor b;
    outputs(1899) <= a xor b;
    outputs(1900) <= b;
    outputs(1901) <= not (a xor b);
    outputs(1902) <= a and not b;
    outputs(1903) <= not b or a;
    outputs(1904) <= not b;
    outputs(1905) <= not b or a;
    outputs(1906) <= not a;
    outputs(1907) <= not (a xor b);
    outputs(1908) <= not (a xor b);
    outputs(1909) <= not b;
    outputs(1910) <= not a;
    outputs(1911) <= not a;
    outputs(1912) <= a;
    outputs(1913) <= a or b;
    outputs(1914) <= b;
    outputs(1915) <= not (a xor b);
    outputs(1916) <= a xor b;
    outputs(1917) <= a xor b;
    outputs(1918) <= a xor b;
    outputs(1919) <= a;
    outputs(1920) <= not a;
    outputs(1921) <= not a;
    outputs(1922) <= b;
    outputs(1923) <= not a;
    outputs(1924) <= not (a xor b);
    outputs(1925) <= a and not b;
    outputs(1926) <= not (a xor b);
    outputs(1927) <= a or b;
    outputs(1928) <= not (a xor b);
    outputs(1929) <= a xor b;
    outputs(1930) <= a and not b;
    outputs(1931) <= a xor b;
    outputs(1932) <= not b;
    outputs(1933) <= b;
    outputs(1934) <= not a or b;
    outputs(1935) <= not (a xor b);
    outputs(1936) <= not (a xor b);
    outputs(1937) <= not a;
    outputs(1938) <= b;
    outputs(1939) <= not (a or b);
    outputs(1940) <= a or b;
    outputs(1941) <= not (a xor b);
    outputs(1942) <= b and not a;
    outputs(1943) <= a;
    outputs(1944) <= not b;
    outputs(1945) <= not a;
    outputs(1946) <= a xor b;
    outputs(1947) <= a and b;
    outputs(1948) <= not (a xor b);
    outputs(1949) <= not (a xor b);
    outputs(1950) <= b and not a;
    outputs(1951) <= not (a or b);
    outputs(1952) <= b and not a;
    outputs(1953) <= not (a xor b);
    outputs(1954) <= b;
    outputs(1955) <= not a;
    outputs(1956) <= a xor b;
    outputs(1957) <= not (a xor b);
    outputs(1958) <= not (a or b);
    outputs(1959) <= not b;
    outputs(1960) <= not b;
    outputs(1961) <= a and b;
    outputs(1962) <= not (a xor b);
    outputs(1963) <= not b;
    outputs(1964) <= a and not b;
    outputs(1965) <= a and b;
    outputs(1966) <= b and not a;
    outputs(1967) <= not b;
    outputs(1968) <= a and b;
    outputs(1969) <= b;
    outputs(1970) <= b;
    outputs(1971) <= not b;
    outputs(1972) <= not (a or b);
    outputs(1973) <= not (a xor b);
    outputs(1974) <= a xor b;
    outputs(1975) <= not a;
    outputs(1976) <= a and b;
    outputs(1977) <= not (a xor b);
    outputs(1978) <= not (a or b);
    outputs(1979) <= a xor b;
    outputs(1980) <= a and not b;
    outputs(1981) <= not a;
    outputs(1982) <= a and b;
    outputs(1983) <= a and b;
    outputs(1984) <= a and not b;
    outputs(1985) <= not (a or b);
    outputs(1986) <= a and b;
    outputs(1987) <= a and b;
    outputs(1988) <= b and not a;
    outputs(1989) <= a;
    outputs(1990) <= a and b;
    outputs(1991) <= not (a xor b);
    outputs(1992) <= a and not b;
    outputs(1993) <= a xor b;
    outputs(1994) <= a and b;
    outputs(1995) <= not (a and b);
    outputs(1996) <= not (a or b);
    outputs(1997) <= b and not a;
    outputs(1998) <= a xor b;
    outputs(1999) <= not (a xor b);
    outputs(2000) <= 1'b0;
    outputs(2001) <= not b or a;
    outputs(2002) <= not (a or b);
    outputs(2003) <= not a;
    outputs(2004) <= a xor b;
    outputs(2005) <= not a;
    outputs(2006) <= a xor b;
    outputs(2007) <= not a;
    outputs(2008) <= not (a xor b);
    outputs(2009) <= a xor b;
    outputs(2010) <= b and not a;
    outputs(2011) <= not (a or b);
    outputs(2012) <= not (a or b);
    outputs(2013) <= a;
    outputs(2014) <= not b;
    outputs(2015) <= not (a or b);
    outputs(2016) <= a xor b;
    outputs(2017) <= a and b;
    outputs(2018) <= b and not a;
    outputs(2019) <= a and b;
    outputs(2020) <= not b;
    outputs(2021) <= not b;
    outputs(2022) <= a and not b;
    outputs(2023) <= a and b;
    outputs(2024) <= a;
    outputs(2025) <= a xor b;
    outputs(2026) <= a;
    outputs(2027) <= b;
    outputs(2028) <= not (a or b);
    outputs(2029) <= a;
    outputs(2030) <= a xor b;
    outputs(2031) <= a and b;
    outputs(2032) <= a;
    outputs(2033) <= not a;
    outputs(2034) <= not b;
    outputs(2035) <= not b;
    outputs(2036) <= b and not a;
    outputs(2037) <= not (a xor b);
    outputs(2038) <= a;
    outputs(2039) <= a;
    outputs(2040) <= a and not b;
    outputs(2041) <= a and b;
    outputs(2042) <= not (a or b);
    outputs(2043) <= a xor b;
    outputs(2044) <= a;
    outputs(2045) <= b;
    outputs(2046) <= a xor b;
    outputs(2047) <= not (a or b);
    outputs(2048) <= not b;
    outputs(2049) <= a xor b;
    outputs(2050) <= not a;
    outputs(2051) <= b;
    outputs(2052) <= not b or a;
    outputs(2053) <= not b;
    outputs(2054) <= not (a or b);
    outputs(2055) <= not (a xor b);
    outputs(2056) <= b and not a;
    outputs(2057) <= not a;
    outputs(2058) <= not a or b;
    outputs(2059) <= b;
    outputs(2060) <= b;
    outputs(2061) <= not (a xor b);
    outputs(2062) <= not (a or b);
    outputs(2063) <= a and not b;
    outputs(2064) <= not a;
    outputs(2065) <= not (a xor b);
    outputs(2066) <= not a;
    outputs(2067) <= b;
    outputs(2068) <= a and not b;
    outputs(2069) <= not (a and b);
    outputs(2070) <= not (a or b);
    outputs(2071) <= a and b;
    outputs(2072) <= not (a xor b);
    outputs(2073) <= not (a xor b);
    outputs(2074) <= not b;
    outputs(2075) <= a or b;
    outputs(2076) <= not (a and b);
    outputs(2077) <= a and not b;
    outputs(2078) <= a xor b;
    outputs(2079) <= a xor b;
    outputs(2080) <= b;
    outputs(2081) <= a and b;
    outputs(2082) <= not (a xor b);
    outputs(2083) <= b and not a;
    outputs(2084) <= a and b;
    outputs(2085) <= not b;
    outputs(2086) <= b and not a;
    outputs(2087) <= not (a xor b);
    outputs(2088) <= a xor b;
    outputs(2089) <= not (a xor b);
    outputs(2090) <= not a or b;
    outputs(2091) <= not b;
    outputs(2092) <= a xor b;
    outputs(2093) <= not (a xor b);
    outputs(2094) <= a xor b;
    outputs(2095) <= not b or a;
    outputs(2096) <= a xor b;
    outputs(2097) <= a and b;
    outputs(2098) <= a xor b;
    outputs(2099) <= not (a xor b);
    outputs(2100) <= b;
    outputs(2101) <= a or b;
    outputs(2102) <= a and b;
    outputs(2103) <= not b;
    outputs(2104) <= not b;
    outputs(2105) <= not (a xor b);
    outputs(2106) <= not b;
    outputs(2107) <= not a;
    outputs(2108) <= not (a and b);
    outputs(2109) <= not a;
    outputs(2110) <= a and b;
    outputs(2111) <= a;
    outputs(2112) <= not (a xor b);
    outputs(2113) <= a xor b;
    outputs(2114) <= a;
    outputs(2115) <= not a;
    outputs(2116) <= a;
    outputs(2117) <= b;
    outputs(2118) <= not (a or b);
    outputs(2119) <= not b;
    outputs(2120) <= not a;
    outputs(2121) <= not (a xor b);
    outputs(2122) <= not a or b;
    outputs(2123) <= not a;
    outputs(2124) <= not a;
    outputs(2125) <= not b or a;
    outputs(2126) <= b and not a;
    outputs(2127) <= a xor b;
    outputs(2128) <= not a;
    outputs(2129) <= not (a xor b);
    outputs(2130) <= not b;
    outputs(2131) <= a and b;
    outputs(2132) <= not a;
    outputs(2133) <= not b;
    outputs(2134) <= b;
    outputs(2135) <= not (a xor b);
    outputs(2136) <= a xor b;
    outputs(2137) <= a or b;
    outputs(2138) <= not b;
    outputs(2139) <= not a;
    outputs(2140) <= a and b;
    outputs(2141) <= a;
    outputs(2142) <= b;
    outputs(2143) <= not b;
    outputs(2144) <= not (a and b);
    outputs(2145) <= b;
    outputs(2146) <= not (a xor b);
    outputs(2147) <= a;
    outputs(2148) <= a;
    outputs(2149) <= b;
    outputs(2150) <= not (a xor b);
    outputs(2151) <= not b;
    outputs(2152) <= not b or a;
    outputs(2153) <= b and not a;
    outputs(2154) <= not a;
    outputs(2155) <= b;
    outputs(2156) <= not a or b;
    outputs(2157) <= not b or a;
    outputs(2158) <= not a;
    outputs(2159) <= a xor b;
    outputs(2160) <= not b;
    outputs(2161) <= not (a xor b);
    outputs(2162) <= a;
    outputs(2163) <= b and not a;
    outputs(2164) <= b and not a;
    outputs(2165) <= not a;
    outputs(2166) <= a xor b;
    outputs(2167) <= a and b;
    outputs(2168) <= a xor b;
    outputs(2169) <= not (a xor b);
    outputs(2170) <= not (a xor b);
    outputs(2171) <= not b;
    outputs(2172) <= a;
    outputs(2173) <= not b;
    outputs(2174) <= b and not a;
    outputs(2175) <= not (a xor b);
    outputs(2176) <= a xor b;
    outputs(2177) <= b;
    outputs(2178) <= not a or b;
    outputs(2179) <= a;
    outputs(2180) <= a or b;
    outputs(2181) <= not b;
    outputs(2182) <= a;
    outputs(2183) <= not (a xor b);
    outputs(2184) <= b and not a;
    outputs(2185) <= not a;
    outputs(2186) <= not a;
    outputs(2187) <= a xor b;
    outputs(2188) <= b and not a;
    outputs(2189) <= not a or b;
    outputs(2190) <= b;
    outputs(2191) <= not b;
    outputs(2192) <= a xor b;
    outputs(2193) <= a;
    outputs(2194) <= a and not b;
    outputs(2195) <= a and not b;
    outputs(2196) <= not a;
    outputs(2197) <= a;
    outputs(2198) <= not (a xor b);
    outputs(2199) <= a;
    outputs(2200) <= a xor b;
    outputs(2201) <= not b or a;
    outputs(2202) <= not (a xor b);
    outputs(2203) <= not (a xor b);
    outputs(2204) <= b;
    outputs(2205) <= a;
    outputs(2206) <= a xor b;
    outputs(2207) <= not b;
    outputs(2208) <= b;
    outputs(2209) <= b and not a;
    outputs(2210) <= a and b;
    outputs(2211) <= not (a xor b);
    outputs(2212) <= a xor b;
    outputs(2213) <= a and b;
    outputs(2214) <= a xor b;
    outputs(2215) <= not (a xor b);
    outputs(2216) <= a xor b;
    outputs(2217) <= not b;
    outputs(2218) <= not b or a;
    outputs(2219) <= not b;
    outputs(2220) <= not b or a;
    outputs(2221) <= b;
    outputs(2222) <= not a or b;
    outputs(2223) <= b and not a;
    outputs(2224) <= not b or a;
    outputs(2225) <= not a;
    outputs(2226) <= not (a or b);
    outputs(2227) <= b;
    outputs(2228) <= a xor b;
    outputs(2229) <= not b;
    outputs(2230) <= not (a and b);
    outputs(2231) <= not a;
    outputs(2232) <= not b or a;
    outputs(2233) <= b;
    outputs(2234) <= a;
    outputs(2235) <= a xor b;
    outputs(2236) <= b and not a;
    outputs(2237) <= not (a xor b);
    outputs(2238) <= not a;
    outputs(2239) <= b;
    outputs(2240) <= a and b;
    outputs(2241) <= not b or a;
    outputs(2242) <= a xor b;
    outputs(2243) <= not (a or b);
    outputs(2244) <= a;
    outputs(2245) <= not b;
    outputs(2246) <= b;
    outputs(2247) <= not (a xor b);
    outputs(2248) <= b;
    outputs(2249) <= a;
    outputs(2250) <= not (a xor b);
    outputs(2251) <= a xor b;
    outputs(2252) <= a;
    outputs(2253) <= not a or b;
    outputs(2254) <= b;
    outputs(2255) <= not (a or b);
    outputs(2256) <= a xor b;
    outputs(2257) <= not b;
    outputs(2258) <= b;
    outputs(2259) <= a and b;
    outputs(2260) <= not a;
    outputs(2261) <= not (a xor b);
    outputs(2262) <= a and not b;
    outputs(2263) <= not a or b;
    outputs(2264) <= a or b;
    outputs(2265) <= b and not a;
    outputs(2266) <= not (a and b);
    outputs(2267) <= not a or b;
    outputs(2268) <= b;
    outputs(2269) <= a;
    outputs(2270) <= b;
    outputs(2271) <= a or b;
    outputs(2272) <= a;
    outputs(2273) <= not (a and b);
    outputs(2274) <= not a;
    outputs(2275) <= b;
    outputs(2276) <= not (a or b);
    outputs(2277) <= a;
    outputs(2278) <= a;
    outputs(2279) <= a or b;
    outputs(2280) <= a;
    outputs(2281) <= a and not b;
    outputs(2282) <= b;
    outputs(2283) <= not a;
    outputs(2284) <= not a;
    outputs(2285) <= not a or b;
    outputs(2286) <= a xor b;
    outputs(2287) <= not b;
    outputs(2288) <= a xor b;
    outputs(2289) <= not b;
    outputs(2290) <= a xor b;
    outputs(2291) <= a;
    outputs(2292) <= b and not a;
    outputs(2293) <= not b;
    outputs(2294) <= not b;
    outputs(2295) <= a and b;
    outputs(2296) <= a xor b;
    outputs(2297) <= a;
    outputs(2298) <= a;
    outputs(2299) <= not b or a;
    outputs(2300) <= a;
    outputs(2301) <= a and b;
    outputs(2302) <= not a;
    outputs(2303) <= a or b;
    outputs(2304) <= not (a or b);
    outputs(2305) <= not b or a;
    outputs(2306) <= not a;
    outputs(2307) <= a xor b;
    outputs(2308) <= b;
    outputs(2309) <= b;
    outputs(2310) <= a;
    outputs(2311) <= b;
    outputs(2312) <= a;
    outputs(2313) <= a or b;
    outputs(2314) <= not (a and b);
    outputs(2315) <= a and b;
    outputs(2316) <= a xor b;
    outputs(2317) <= not (a and b);
    outputs(2318) <= not (a xor b);
    outputs(2319) <= not a;
    outputs(2320) <= b;
    outputs(2321) <= a xor b;
    outputs(2322) <= not a;
    outputs(2323) <= not a or b;
    outputs(2324) <= not a;
    outputs(2325) <= not (a xor b);
    outputs(2326) <= b and not a;
    outputs(2327) <= b;
    outputs(2328) <= b;
    outputs(2329) <= a or b;
    outputs(2330) <= not a;
    outputs(2331) <= a;
    outputs(2332) <= a xor b;
    outputs(2333) <= not b;
    outputs(2334) <= not (a and b);
    outputs(2335) <= a;
    outputs(2336) <= not (a xor b);
    outputs(2337) <= not a or b;
    outputs(2338) <= not a;
    outputs(2339) <= b;
    outputs(2340) <= b;
    outputs(2341) <= not (a xor b);
    outputs(2342) <= not (a xor b);
    outputs(2343) <= a;
    outputs(2344) <= not b;
    outputs(2345) <= not (a xor b);
    outputs(2346) <= not (a or b);
    outputs(2347) <= not b;
    outputs(2348) <= not (a xor b);
    outputs(2349) <= a xor b;
    outputs(2350) <= not (a xor b);
    outputs(2351) <= not a;
    outputs(2352) <= a;
    outputs(2353) <= not (a or b);
    outputs(2354) <= a and not b;
    outputs(2355) <= a xor b;
    outputs(2356) <= not b;
    outputs(2357) <= a xor b;
    outputs(2358) <= a;
    outputs(2359) <= b;
    outputs(2360) <= not (a xor b);
    outputs(2361) <= a xor b;
    outputs(2362) <= b and not a;
    outputs(2363) <= a or b;
    outputs(2364) <= not b;
    outputs(2365) <= a;
    outputs(2366) <= not a or b;
    outputs(2367) <= a and not b;
    outputs(2368) <= a and b;
    outputs(2369) <= not a;
    outputs(2370) <= not (a or b);
    outputs(2371) <= a;
    outputs(2372) <= a or b;
    outputs(2373) <= a;
    outputs(2374) <= b and not a;
    outputs(2375) <= not b;
    outputs(2376) <= not a or b;
    outputs(2377) <= a;
    outputs(2378) <= a xor b;
    outputs(2379) <= not (a and b);
    outputs(2380) <= a and b;
    outputs(2381) <= not b;
    outputs(2382) <= a xor b;
    outputs(2383) <= not b;
    outputs(2384) <= a;
    outputs(2385) <= not (a xor b);
    outputs(2386) <= not (a and b);
    outputs(2387) <= a;
    outputs(2388) <= a or b;
    outputs(2389) <= not (a xor b);
    outputs(2390) <= not (a and b);
    outputs(2391) <= a and not b;
    outputs(2392) <= a and b;
    outputs(2393) <= b and not a;
    outputs(2394) <= not a;
    outputs(2395) <= not a or b;
    outputs(2396) <= a;
    outputs(2397) <= a;
    outputs(2398) <= a xor b;
    outputs(2399) <= a and b;
    outputs(2400) <= not b;
    outputs(2401) <= a;
    outputs(2402) <= b and not a;
    outputs(2403) <= not a;
    outputs(2404) <= not a or b;
    outputs(2405) <= b;
    outputs(2406) <= a and b;
    outputs(2407) <= b;
    outputs(2408) <= a or b;
    outputs(2409) <= not (a xor b);
    outputs(2410) <= not b;
    outputs(2411) <= b and not a;
    outputs(2412) <= b;
    outputs(2413) <= a xor b;
    outputs(2414) <= not b or a;
    outputs(2415) <= not a;
    outputs(2416) <= not b;
    outputs(2417) <= not b or a;
    outputs(2418) <= not a;
    outputs(2419) <= not (a xor b);
    outputs(2420) <= a xor b;
    outputs(2421) <= not a;
    outputs(2422) <= not a;
    outputs(2423) <= a and not b;
    outputs(2424) <= a xor b;
    outputs(2425) <= not (a and b);
    outputs(2426) <= not a;
    outputs(2427) <= a xor b;
    outputs(2428) <= not b or a;
    outputs(2429) <= not a;
    outputs(2430) <= not b;
    outputs(2431) <= a xor b;
    outputs(2432) <= a xor b;
    outputs(2433) <= not (a and b);
    outputs(2434) <= not a;
    outputs(2435) <= a xor b;
    outputs(2436) <= not (a and b);
    outputs(2437) <= not b;
    outputs(2438) <= a xor b;
    outputs(2439) <= not a or b;
    outputs(2440) <= not b or a;
    outputs(2441) <= not a or b;
    outputs(2442) <= a xor b;
    outputs(2443) <= not b;
    outputs(2444) <= not a;
    outputs(2445) <= not a or b;
    outputs(2446) <= not b;
    outputs(2447) <= b;
    outputs(2448) <= not (a xor b);
    outputs(2449) <= a xor b;
    outputs(2450) <= not (a and b);
    outputs(2451) <= a;
    outputs(2452) <= b;
    outputs(2453) <= not b;
    outputs(2454) <= a xor b;
    outputs(2455) <= a or b;
    outputs(2456) <= not a;
    outputs(2457) <= a or b;
    outputs(2458) <= not b;
    outputs(2459) <= not (a or b);
    outputs(2460) <= not b;
    outputs(2461) <= b;
    outputs(2462) <= not b;
    outputs(2463) <= not b or a;
    outputs(2464) <= not b or a;
    outputs(2465) <= b and not a;
    outputs(2466) <= b and not a;
    outputs(2467) <= a xor b;
    outputs(2468) <= a xor b;
    outputs(2469) <= a;
    outputs(2470) <= not b;
    outputs(2471) <= not (a and b);
    outputs(2472) <= a xor b;
    outputs(2473) <= a xor b;
    outputs(2474) <= not b or a;
    outputs(2475) <= not (a xor b);
    outputs(2476) <= not a or b;
    outputs(2477) <= not b;
    outputs(2478) <= not b;
    outputs(2479) <= not b;
    outputs(2480) <= not (a and b);
    outputs(2481) <= not (a xor b);
    outputs(2482) <= b;
    outputs(2483) <= not b;
    outputs(2484) <= a;
    outputs(2485) <= a and b;
    outputs(2486) <= not b;
    outputs(2487) <= not (a xor b);
    outputs(2488) <= not a or b;
    outputs(2489) <= not a;
    outputs(2490) <= a or b;
    outputs(2491) <= b and not a;
    outputs(2492) <= a xor b;
    outputs(2493) <= a;
    outputs(2494) <= b;
    outputs(2495) <= not (a or b);
    outputs(2496) <= not (a and b);
    outputs(2497) <= not (a and b);
    outputs(2498) <= a xor b;
    outputs(2499) <= not b;
    outputs(2500) <= a and not b;
    outputs(2501) <= not b;
    outputs(2502) <= not a;
    outputs(2503) <= b;
    outputs(2504) <= a xor b;
    outputs(2505) <= a;
    outputs(2506) <= a xor b;
    outputs(2507) <= b;
    outputs(2508) <= not (a xor b);
    outputs(2509) <= not b;
    outputs(2510) <= not (a xor b);
    outputs(2511) <= not a;
    outputs(2512) <= b;
    outputs(2513) <= b and not a;
    outputs(2514) <= not b or a;
    outputs(2515) <= not (a xor b);
    outputs(2516) <= not a;
    outputs(2517) <= a;
    outputs(2518) <= not (a or b);
    outputs(2519) <= not b;
    outputs(2520) <= a and not b;
    outputs(2521) <= a;
    outputs(2522) <= a;
    outputs(2523) <= not (a and b);
    outputs(2524) <= a or b;
    outputs(2525) <= not (a xor b);
    outputs(2526) <= not b;
    outputs(2527) <= a or b;
    outputs(2528) <= not (a and b);
    outputs(2529) <= a;
    outputs(2530) <= a xor b;
    outputs(2531) <= not (a xor b);
    outputs(2532) <= not a;
    outputs(2533) <= not b;
    outputs(2534) <= a xor b;
    outputs(2535) <= not a or b;
    outputs(2536) <= not a;
    outputs(2537) <= not a or b;
    outputs(2538) <= not a or b;
    outputs(2539) <= a and b;
    outputs(2540) <= a;
    outputs(2541) <= a or b;
    outputs(2542) <= a and not b;
    outputs(2543) <= a and not b;
    outputs(2544) <= a;
    outputs(2545) <= not a;
    outputs(2546) <= a and b;
    outputs(2547) <= not (a xor b);
    outputs(2548) <= a xor b;
    outputs(2549) <= not b;
    outputs(2550) <= not a;
    outputs(2551) <= not (a or b);
    outputs(2552) <= not b;
    outputs(2553) <= not b;
    outputs(2554) <= a;
    outputs(2555) <= a and not b;
    outputs(2556) <= not (a and b);
    outputs(2557) <= not b;
    outputs(2558) <= a;
    outputs(2559) <= b;
    outputs(2560) <= not (a xor b);
    outputs(2561) <= a;
    outputs(2562) <= b;
    outputs(2563) <= not (a xor b);
    outputs(2564) <= not (a xor b);
    outputs(2565) <= not (a xor b);
    outputs(2566) <= not (a xor b);
    outputs(2567) <= not a;
    outputs(2568) <= a xor b;
    outputs(2569) <= b;
    outputs(2570) <= not a;
    outputs(2571) <= b and not a;
    outputs(2572) <= a;
    outputs(2573) <= not (a xor b);
    outputs(2574) <= b;
    outputs(2575) <= a or b;
    outputs(2576) <= not b or a;
    outputs(2577) <= not a;
    outputs(2578) <= a xor b;
    outputs(2579) <= b;
    outputs(2580) <= not a;
    outputs(2581) <= not a;
    outputs(2582) <= a;
    outputs(2583) <= not b;
    outputs(2584) <= a or b;
    outputs(2585) <= not b;
    outputs(2586) <= not a or b;
    outputs(2587) <= a xor b;
    outputs(2588) <= not a;
    outputs(2589) <= a;
    outputs(2590) <= a;
    outputs(2591) <= b and not a;
    outputs(2592) <= not (a and b);
    outputs(2593) <= not a;
    outputs(2594) <= not (a xor b);
    outputs(2595) <= not b or a;
    outputs(2596) <= b;
    outputs(2597) <= b and not a;
    outputs(2598) <= not a or b;
    outputs(2599) <= not b or a;
    outputs(2600) <= b;
    outputs(2601) <= not (a xor b);
    outputs(2602) <= b;
    outputs(2603) <= a;
    outputs(2604) <= a xor b;
    outputs(2605) <= not b;
    outputs(2606) <= a xor b;
    outputs(2607) <= a xor b;
    outputs(2608) <= b and not a;
    outputs(2609) <= a;
    outputs(2610) <= not (a xor b);
    outputs(2611) <= b and not a;
    outputs(2612) <= not a;
    outputs(2613) <= a;
    outputs(2614) <= a xor b;
    outputs(2615) <= a xor b;
    outputs(2616) <= not (a and b);
    outputs(2617) <= a and not b;
    outputs(2618) <= not a;
    outputs(2619) <= a;
    outputs(2620) <= not (a xor b);
    outputs(2621) <= a;
    outputs(2622) <= a;
    outputs(2623) <= b;
    outputs(2624) <= not b;
    outputs(2625) <= not b;
    outputs(2626) <= a;
    outputs(2627) <= not a or b;
    outputs(2628) <= not (a and b);
    outputs(2629) <= not a;
    outputs(2630) <= a;
    outputs(2631) <= b;
    outputs(2632) <= a xor b;
    outputs(2633) <= a or b;
    outputs(2634) <= a or b;
    outputs(2635) <= not (a xor b);
    outputs(2636) <= a xor b;
    outputs(2637) <= not b;
    outputs(2638) <= a xor b;
    outputs(2639) <= not (a xor b);
    outputs(2640) <= b;
    outputs(2641) <= not (a xor b);
    outputs(2642) <= b;
    outputs(2643) <= a or b;
    outputs(2644) <= not b or a;
    outputs(2645) <= b;
    outputs(2646) <= not (a xor b);
    outputs(2647) <= not (a and b);
    outputs(2648) <= a xor b;
    outputs(2649) <= a;
    outputs(2650) <= a or b;
    outputs(2651) <= a xor b;
    outputs(2652) <= a and b;
    outputs(2653) <= a;
    outputs(2654) <= not (a xor b);
    outputs(2655) <= not a or b;
    outputs(2656) <= not (a xor b);
    outputs(2657) <= not a or b;
    outputs(2658) <= a and b;
    outputs(2659) <= not (a and b);
    outputs(2660) <= a;
    outputs(2661) <= b and not a;
    outputs(2662) <= a xor b;
    outputs(2663) <= b and not a;
    outputs(2664) <= a;
    outputs(2665) <= not b;
    outputs(2666) <= b;
    outputs(2667) <= not (a or b);
    outputs(2668) <= a and b;
    outputs(2669) <= a and not b;
    outputs(2670) <= not a or b;
    outputs(2671) <= b;
    outputs(2672) <= not (a xor b);
    outputs(2673) <= not b;
    outputs(2674) <= a xor b;
    outputs(2675) <= not (a xor b);
    outputs(2676) <= not (a and b);
    outputs(2677) <= not a or b;
    outputs(2678) <= not b;
    outputs(2679) <= a and not b;
    outputs(2680) <= b;
    outputs(2681) <= b;
    outputs(2682) <= not b or a;
    outputs(2683) <= a xor b;
    outputs(2684) <= a;
    outputs(2685) <= b;
    outputs(2686) <= not b or a;
    outputs(2687) <= not (a xor b);
    outputs(2688) <= a xor b;
    outputs(2689) <= not (a and b);
    outputs(2690) <= not a;
    outputs(2691) <= not b or a;
    outputs(2692) <= not (a and b);
    outputs(2693) <= a xor b;
    outputs(2694) <= not (a xor b);
    outputs(2695) <= not a;
    outputs(2696) <= not a;
    outputs(2697) <= not a;
    outputs(2698) <= not a;
    outputs(2699) <= not b;
    outputs(2700) <= not (a xor b);
    outputs(2701) <= b and not a;
    outputs(2702) <= not b;
    outputs(2703) <= not a;
    outputs(2704) <= not b;
    outputs(2705) <= a and not b;
    outputs(2706) <= b and not a;
    outputs(2707) <= not a;
    outputs(2708) <= b;
    outputs(2709) <= not (a xor b);
    outputs(2710) <= a and not b;
    outputs(2711) <= not a or b;
    outputs(2712) <= b and not a;
    outputs(2713) <= a or b;
    outputs(2714) <= b and not a;
    outputs(2715) <= b and not a;
    outputs(2716) <= not a;
    outputs(2717) <= not a;
    outputs(2718) <= not b or a;
    outputs(2719) <= not b;
    outputs(2720) <= b;
    outputs(2721) <= not (a and b);
    outputs(2722) <= a xor b;
    outputs(2723) <= not (a xor b);
    outputs(2724) <= not (a xor b);
    outputs(2725) <= a xor b;
    outputs(2726) <= not (a xor b);
    outputs(2727) <= a;
    outputs(2728) <= not b;
    outputs(2729) <= not (a xor b);
    outputs(2730) <= not (a xor b);
    outputs(2731) <= a and b;
    outputs(2732) <= a xor b;
    outputs(2733) <= not a;
    outputs(2734) <= a or b;
    outputs(2735) <= not a;
    outputs(2736) <= a;
    outputs(2737) <= not a or b;
    outputs(2738) <= a xor b;
    outputs(2739) <= a;
    outputs(2740) <= a xor b;
    outputs(2741) <= not a or b;
    outputs(2742) <= not b or a;
    outputs(2743) <= not (a xor b);
    outputs(2744) <= not a;
    outputs(2745) <= a xor b;
    outputs(2746) <= not (a and b);
    outputs(2747) <= not (a xor b);
    outputs(2748) <= a or b;
    outputs(2749) <= not (a xor b);
    outputs(2750) <= b;
    outputs(2751) <= b;
    outputs(2752) <= not (a xor b);
    outputs(2753) <= a;
    outputs(2754) <= not b;
    outputs(2755) <= not (a or b);
    outputs(2756) <= a;
    outputs(2757) <= b and not a;
    outputs(2758) <= not (a xor b);
    outputs(2759) <= a or b;
    outputs(2760) <= not (a xor b);
    outputs(2761) <= a;
    outputs(2762) <= not (a and b);
    outputs(2763) <= a;
    outputs(2764) <= a and not b;
    outputs(2765) <= a;
    outputs(2766) <= not (a xor b);
    outputs(2767) <= not (a xor b);
    outputs(2768) <= a and not b;
    outputs(2769) <= a xor b;
    outputs(2770) <= not a;
    outputs(2771) <= not (a xor b);
    outputs(2772) <= not (a xor b);
    outputs(2773) <= a;
    outputs(2774) <= not (a xor b);
    outputs(2775) <= a and b;
    outputs(2776) <= b and not a;
    outputs(2777) <= a xor b;
    outputs(2778) <= b;
    outputs(2779) <= a and not b;
    outputs(2780) <= b and not a;
    outputs(2781) <= a;
    outputs(2782) <= not (a xor b);
    outputs(2783) <= not (a xor b);
    outputs(2784) <= a and b;
    outputs(2785) <= a xor b;
    outputs(2786) <= a and not b;
    outputs(2787) <= not (a and b);
    outputs(2788) <= not (a xor b);
    outputs(2789) <= not a;
    outputs(2790) <= not (a and b);
    outputs(2791) <= not b;
    outputs(2792) <= not b;
    outputs(2793) <= a or b;
    outputs(2794) <= not (a xor b);
    outputs(2795) <= not (a xor b);
    outputs(2796) <= not a;
    outputs(2797) <= not (a xor b);
    outputs(2798) <= not (a xor b);
    outputs(2799) <= a;
    outputs(2800) <= not a;
    outputs(2801) <= a xor b;
    outputs(2802) <= a;
    outputs(2803) <= a and b;
    outputs(2804) <= a and not b;
    outputs(2805) <= not a;
    outputs(2806) <= not b;
    outputs(2807) <= not (a and b);
    outputs(2808) <= b;
    outputs(2809) <= not (a and b);
    outputs(2810) <= a;
    outputs(2811) <= not a;
    outputs(2812) <= a or b;
    outputs(2813) <= a and not b;
    outputs(2814) <= not a;
    outputs(2815) <= b;
    outputs(2816) <= not b;
    outputs(2817) <= not (a xor b);
    outputs(2818) <= b and not a;
    outputs(2819) <= b;
    outputs(2820) <= not a;
    outputs(2821) <= not (a or b);
    outputs(2822) <= b;
    outputs(2823) <= not a;
    outputs(2824) <= not a;
    outputs(2825) <= not b;
    outputs(2826) <= not (a or b);
    outputs(2827) <= b;
    outputs(2828) <= not b;
    outputs(2829) <= a and not b;
    outputs(2830) <= a xor b;
    outputs(2831) <= not a;
    outputs(2832) <= not (a or b);
    outputs(2833) <= b;
    outputs(2834) <= a;
    outputs(2835) <= b;
    outputs(2836) <= a and b;
    outputs(2837) <= a xor b;
    outputs(2838) <= not (a xor b);
    outputs(2839) <= a and not b;
    outputs(2840) <= a or b;
    outputs(2841) <= a xor b;
    outputs(2842) <= not (a xor b);
    outputs(2843) <= a and not b;
    outputs(2844) <= a xor b;
    outputs(2845) <= not (a or b);
    outputs(2846) <= b;
    outputs(2847) <= not b;
    outputs(2848) <= not a or b;
    outputs(2849) <= not (a xor b);
    outputs(2850) <= not (a xor b);
    outputs(2851) <= b;
    outputs(2852) <= not (a or b);
    outputs(2853) <= not a or b;
    outputs(2854) <= b;
    outputs(2855) <= not b;
    outputs(2856) <= b;
    outputs(2857) <= a xor b;
    outputs(2858) <= not a;
    outputs(2859) <= not (a or b);
    outputs(2860) <= not b;
    outputs(2861) <= not (a xor b);
    outputs(2862) <= a and b;
    outputs(2863) <= a xor b;
    outputs(2864) <= not a or b;
    outputs(2865) <= a;
    outputs(2866) <= not a;
    outputs(2867) <= not (a and b);
    outputs(2868) <= not (a and b);
    outputs(2869) <= not a;
    outputs(2870) <= a xor b;
    outputs(2871) <= b and not a;
    outputs(2872) <= not (a xor b);
    outputs(2873) <= b;
    outputs(2874) <= a;
    outputs(2875) <= not (a xor b);
    outputs(2876) <= b;
    outputs(2877) <= a and not b;
    outputs(2878) <= a;
    outputs(2879) <= not a;
    outputs(2880) <= a xor b;
    outputs(2881) <= a;
    outputs(2882) <= a;
    outputs(2883) <= a;
    outputs(2884) <= a;
    outputs(2885) <= a xor b;
    outputs(2886) <= b;
    outputs(2887) <= a and not b;
    outputs(2888) <= not b;
    outputs(2889) <= b;
    outputs(2890) <= a;
    outputs(2891) <= not b;
    outputs(2892) <= not a or b;
    outputs(2893) <= a xor b;
    outputs(2894) <= not (a xor b);
    outputs(2895) <= not (a and b);
    outputs(2896) <= not b or a;
    outputs(2897) <= not a;
    outputs(2898) <= not a or b;
    outputs(2899) <= a;
    outputs(2900) <= b;
    outputs(2901) <= a;
    outputs(2902) <= not (a and b);
    outputs(2903) <= b;
    outputs(2904) <= a xor b;
    outputs(2905) <= not a;
    outputs(2906) <= not b or a;
    outputs(2907) <= not b or a;
    outputs(2908) <= a;
    outputs(2909) <= not (a xor b);
    outputs(2910) <= a or b;
    outputs(2911) <= not (a or b);
    outputs(2912) <= not b;
    outputs(2913) <= not (a and b);
    outputs(2914) <= b and not a;
    outputs(2915) <= not b;
    outputs(2916) <= a xor b;
    outputs(2917) <= not b or a;
    outputs(2918) <= not b or a;
    outputs(2919) <= a;
    outputs(2920) <= not a or b;
    outputs(2921) <= a xor b;
    outputs(2922) <= b and not a;
    outputs(2923) <= a;
    outputs(2924) <= not (a xor b);
    outputs(2925) <= not (a and b);
    outputs(2926) <= not a;
    outputs(2927) <= a xor b;
    outputs(2928) <= b and not a;
    outputs(2929) <= a xor b;
    outputs(2930) <= not a or b;
    outputs(2931) <= not b;
    outputs(2932) <= not a;
    outputs(2933) <= not b;
    outputs(2934) <= not (a and b);
    outputs(2935) <= not (a xor b);
    outputs(2936) <= not a;
    outputs(2937) <= a or b;
    outputs(2938) <= b and not a;
    outputs(2939) <= not a;
    outputs(2940) <= not b;
    outputs(2941) <= not b;
    outputs(2942) <= not b;
    outputs(2943) <= a;
    outputs(2944) <= not (a and b);
    outputs(2945) <= a;
    outputs(2946) <= b;
    outputs(2947) <= not a;
    outputs(2948) <= a;
    outputs(2949) <= not a;
    outputs(2950) <= not a or b;
    outputs(2951) <= not b or a;
    outputs(2952) <= a and b;
    outputs(2953) <= a and not b;
    outputs(2954) <= not (a xor b);
    outputs(2955) <= a xor b;
    outputs(2956) <= a;
    outputs(2957) <= a and b;
    outputs(2958) <= b and not a;
    outputs(2959) <= not (a xor b);
    outputs(2960) <= a and not b;
    outputs(2961) <= b;
    outputs(2962) <= not a;
    outputs(2963) <= a;
    outputs(2964) <= a or b;
    outputs(2965) <= not (a and b);
    outputs(2966) <= not (a xor b);
    outputs(2967) <= a xor b;
    outputs(2968) <= not b or a;
    outputs(2969) <= a;
    outputs(2970) <= a xor b;
    outputs(2971) <= not (a xor b);
    outputs(2972) <= b;
    outputs(2973) <= b;
    outputs(2974) <= not a or b;
    outputs(2975) <= not (a xor b);
    outputs(2976) <= a xor b;
    outputs(2977) <= not a or b;
    outputs(2978) <= not (a and b);
    outputs(2979) <= not (a xor b);
    outputs(2980) <= not (a xor b);
    outputs(2981) <= a and not b;
    outputs(2982) <= not a or b;
    outputs(2983) <= b;
    outputs(2984) <= not (a xor b);
    outputs(2985) <= a or b;
    outputs(2986) <= a xor b;
    outputs(2987) <= a;
    outputs(2988) <= a;
    outputs(2989) <= not b;
    outputs(2990) <= not b;
    outputs(2991) <= a or b;
    outputs(2992) <= b and not a;
    outputs(2993) <= a;
    outputs(2994) <= b;
    outputs(2995) <= not (a xor b);
    outputs(2996) <= not b;
    outputs(2997) <= b;
    outputs(2998) <= not b;
    outputs(2999) <= not b or a;
    outputs(3000) <= not (a xor b);
    outputs(3001) <= a;
    outputs(3002) <= a xor b;
    outputs(3003) <= a xor b;
    outputs(3004) <= not a or b;
    outputs(3005) <= not b or a;
    outputs(3006) <= b;
    outputs(3007) <= not a;
    outputs(3008) <= a and b;
    outputs(3009) <= not (a and b);
    outputs(3010) <= not b or a;
    outputs(3011) <= a and not b;
    outputs(3012) <= not (a or b);
    outputs(3013) <= b and not a;
    outputs(3014) <= not (a xor b);
    outputs(3015) <= not b;
    outputs(3016) <= not a or b;
    outputs(3017) <= not (a or b);
    outputs(3018) <= a xor b;
    outputs(3019) <= a xor b;
    outputs(3020) <= not (a and b);
    outputs(3021) <= not b;
    outputs(3022) <= not (a xor b);
    outputs(3023) <= not (a xor b);
    outputs(3024) <= not a or b;
    outputs(3025) <= b;
    outputs(3026) <= a;
    outputs(3027) <= not (a or b);
    outputs(3028) <= not (a or b);
    outputs(3029) <= a and not b;
    outputs(3030) <= not b;
    outputs(3031) <= not a or b;
    outputs(3032) <= not b or a;
    outputs(3033) <= b;
    outputs(3034) <= not a;
    outputs(3035) <= not a;
    outputs(3036) <= not (a xor b);
    outputs(3037) <= not a;
    outputs(3038) <= a;
    outputs(3039) <= not b;
    outputs(3040) <= b;
    outputs(3041) <= not b or a;
    outputs(3042) <= a and b;
    outputs(3043) <= a;
    outputs(3044) <= not a;
    outputs(3045) <= a and b;
    outputs(3046) <= b;
    outputs(3047) <= a xor b;
    outputs(3048) <= not (a xor b);
    outputs(3049) <= not b;
    outputs(3050) <= not (a xor b);
    outputs(3051) <= a;
    outputs(3052) <= not (a or b);
    outputs(3053) <= not (a xor b);
    outputs(3054) <= not b;
    outputs(3055) <= not a;
    outputs(3056) <= not (a and b);
    outputs(3057) <= not (a xor b);
    outputs(3058) <= not (a xor b);
    outputs(3059) <= b and not a;
    outputs(3060) <= not a;
    outputs(3061) <= not b;
    outputs(3062) <= b and not a;
    outputs(3063) <= not a or b;
    outputs(3064) <= a;
    outputs(3065) <= a xor b;
    outputs(3066) <= b;
    outputs(3067) <= b;
    outputs(3068) <= not b;
    outputs(3069) <= a and b;
    outputs(3070) <= not (a xor b);
    outputs(3071) <= a;
    outputs(3072) <= not (a xor b);
    outputs(3073) <= b;
    outputs(3074) <= not (a xor b);
    outputs(3075) <= not (a xor b);
    outputs(3076) <= not (a xor b);
    outputs(3077) <= not a;
    outputs(3078) <= a;
    outputs(3079) <= not a;
    outputs(3080) <= a and not b;
    outputs(3081) <= not b or a;
    outputs(3082) <= not (a xor b);
    outputs(3083) <= not (a and b);
    outputs(3084) <= a;
    outputs(3085) <= not (a xor b);
    outputs(3086) <= not a;
    outputs(3087) <= not a or b;
    outputs(3088) <= not (a xor b);
    outputs(3089) <= a or b;
    outputs(3090) <= b;
    outputs(3091) <= not (a or b);
    outputs(3092) <= b;
    outputs(3093) <= not (a and b);
    outputs(3094) <= not b;
    outputs(3095) <= not a;
    outputs(3096) <= a and not b;
    outputs(3097) <= not b;
    outputs(3098) <= a xor b;
    outputs(3099) <= not a or b;
    outputs(3100) <= a and b;
    outputs(3101) <= not a;
    outputs(3102) <= a xor b;
    outputs(3103) <= a and b;
    outputs(3104) <= not (a and b);
    outputs(3105) <= not b;
    outputs(3106) <= a and b;
    outputs(3107) <= not (a xor b);
    outputs(3108) <= a;
    outputs(3109) <= a xor b;
    outputs(3110) <= not a;
    outputs(3111) <= not b;
    outputs(3112) <= a or b;
    outputs(3113) <= a;
    outputs(3114) <= not a;
    outputs(3115) <= not a;
    outputs(3116) <= not a;
    outputs(3117) <= b and not a;
    outputs(3118) <= b;
    outputs(3119) <= a xor b;
    outputs(3120) <= not a or b;
    outputs(3121) <= not a;
    outputs(3122) <= not (a xor b);
    outputs(3123) <= a xor b;
    outputs(3124) <= not (a or b);
    outputs(3125) <= a xor b;
    outputs(3126) <= not (a and b);
    outputs(3127) <= not b;
    outputs(3128) <= not (a xor b);
    outputs(3129) <= not (a xor b);
    outputs(3130) <= not b;
    outputs(3131) <= not (a xor b);
    outputs(3132) <= a xor b;
    outputs(3133) <= a xor b;
    outputs(3134) <= a or b;
    outputs(3135) <= not (a and b);
    outputs(3136) <= b;
    outputs(3137) <= a xor b;
    outputs(3138) <= not a;
    outputs(3139) <= b and not a;
    outputs(3140) <= not b or a;
    outputs(3141) <= b;
    outputs(3142) <= b and not a;
    outputs(3143) <= a;
    outputs(3144) <= not (a or b);
    outputs(3145) <= not (a xor b);
    outputs(3146) <= a xor b;
    outputs(3147) <= b;
    outputs(3148) <= b and not a;
    outputs(3149) <= a;
    outputs(3150) <= not (a xor b);
    outputs(3151) <= not a;
    outputs(3152) <= not (a or b);
    outputs(3153) <= not a or b;
    outputs(3154) <= a xor b;
    outputs(3155) <= a or b;
    outputs(3156) <= not (a and b);
    outputs(3157) <= not (a xor b);
    outputs(3158) <= not a or b;
    outputs(3159) <= a and not b;
    outputs(3160) <= not b;
    outputs(3161) <= not b;
    outputs(3162) <= not b;
    outputs(3163) <= a;
    outputs(3164) <= not a or b;
    outputs(3165) <= b;
    outputs(3166) <= a and not b;
    outputs(3167) <= a xor b;
    outputs(3168) <= a xor b;
    outputs(3169) <= a xor b;
    outputs(3170) <= a;
    outputs(3171) <= b;
    outputs(3172) <= not b;
    outputs(3173) <= not b;
    outputs(3174) <= b;
    outputs(3175) <= b;
    outputs(3176) <= not a;
    outputs(3177) <= a and not b;
    outputs(3178) <= a;
    outputs(3179) <= a xor b;
    outputs(3180) <= not a;
    outputs(3181) <= a;
    outputs(3182) <= a xor b;
    outputs(3183) <= a;
    outputs(3184) <= a;
    outputs(3185) <= not a or b;
    outputs(3186) <= not a;
    outputs(3187) <= not (a or b);
    outputs(3188) <= a;
    outputs(3189) <= not a or b;
    outputs(3190) <= a or b;
    outputs(3191) <= not a;
    outputs(3192) <= a;
    outputs(3193) <= not b or a;
    outputs(3194) <= a or b;
    outputs(3195) <= not (a xor b);
    outputs(3196) <= not b or a;
    outputs(3197) <= not (a or b);
    outputs(3198) <= not (a xor b);
    outputs(3199) <= a xor b;
    outputs(3200) <= not a;
    outputs(3201) <= not (a or b);
    outputs(3202) <= not (a xor b);
    outputs(3203) <= not (a xor b);
    outputs(3204) <= not (a and b);
    outputs(3205) <= not b;
    outputs(3206) <= not (a xor b);
    outputs(3207) <= a xor b;
    outputs(3208) <= b;
    outputs(3209) <= a and b;
    outputs(3210) <= not b;
    outputs(3211) <= a or b;
    outputs(3212) <= not b;
    outputs(3213) <= not (a or b);
    outputs(3214) <= not (a or b);
    outputs(3215) <= a xor b;
    outputs(3216) <= not (a or b);
    outputs(3217) <= a;
    outputs(3218) <= not a;
    outputs(3219) <= b;
    outputs(3220) <= a xor b;
    outputs(3221) <= a;
    outputs(3222) <= a xor b;
    outputs(3223) <= not (a or b);
    outputs(3224) <= not a;
    outputs(3225) <= a and b;
    outputs(3226) <= not (a xor b);
    outputs(3227) <= not (a xor b);
    outputs(3228) <= a and b;
    outputs(3229) <= b;
    outputs(3230) <= b;
    outputs(3231) <= a and not b;
    outputs(3232) <= b and not a;
    outputs(3233) <= b;
    outputs(3234) <= not (a or b);
    outputs(3235) <= not a;
    outputs(3236) <= a;
    outputs(3237) <= not b or a;
    outputs(3238) <= not (a and b);
    outputs(3239) <= not (a xor b);
    outputs(3240) <= a or b;
    outputs(3241) <= b;
    outputs(3242) <= a xor b;
    outputs(3243) <= not a or b;
    outputs(3244) <= a and b;
    outputs(3245) <= not b or a;
    outputs(3246) <= not a;
    outputs(3247) <= not a;
    outputs(3248) <= not (a or b);
    outputs(3249) <= a or b;
    outputs(3250) <= a xor b;
    outputs(3251) <= not (a xor b);
    outputs(3252) <= a xor b;
    outputs(3253) <= not a;
    outputs(3254) <= not (a xor b);
    outputs(3255) <= not (a and b);
    outputs(3256) <= not a;
    outputs(3257) <= b;
    outputs(3258) <= not b;
    outputs(3259) <= a;
    outputs(3260) <= not b;
    outputs(3261) <= a xor b;
    outputs(3262) <= not (a and b);
    outputs(3263) <= not b;
    outputs(3264) <= b;
    outputs(3265) <= a and not b;
    outputs(3266) <= a;
    outputs(3267) <= b;
    outputs(3268) <= not (a or b);
    outputs(3269) <= b and not a;
    outputs(3270) <= not (a xor b);
    outputs(3271) <= not a;
    outputs(3272) <= not b;
    outputs(3273) <= not b;
    outputs(3274) <= b;
    outputs(3275) <= not (a xor b);
    outputs(3276) <= a and b;
    outputs(3277) <= b;
    outputs(3278) <= not b;
    outputs(3279) <= not a or b;
    outputs(3280) <= not (a xor b);
    outputs(3281) <= not a;
    outputs(3282) <= b and not a;
    outputs(3283) <= not (a xor b);
    outputs(3284) <= b;
    outputs(3285) <= b and not a;
    outputs(3286) <= a;
    outputs(3287) <= not a or b;
    outputs(3288) <= not b;
    outputs(3289) <= not a;
    outputs(3290) <= a xor b;
    outputs(3291) <= b and not a;
    outputs(3292) <= b;
    outputs(3293) <= not a;
    outputs(3294) <= a;
    outputs(3295) <= a xor b;
    outputs(3296) <= b;
    outputs(3297) <= a;
    outputs(3298) <= not (a xor b);
    outputs(3299) <= not b;
    outputs(3300) <= a;
    outputs(3301) <= not a or b;
    outputs(3302) <= not a;
    outputs(3303) <= a and b;
    outputs(3304) <= a xor b;
    outputs(3305) <= a xor b;
    outputs(3306) <= b;
    outputs(3307) <= a xor b;
    outputs(3308) <= a;
    outputs(3309) <= not (a xor b);
    outputs(3310) <= b and not a;
    outputs(3311) <= not (a xor b);
    outputs(3312) <= not a or b;
    outputs(3313) <= not (a xor b);
    outputs(3314) <= b;
    outputs(3315) <= a xor b;
    outputs(3316) <= not (a xor b);
    outputs(3317) <= a;
    outputs(3318) <= b;
    outputs(3319) <= a and b;
    outputs(3320) <= a;
    outputs(3321) <= a;
    outputs(3322) <= a xor b;
    outputs(3323) <= not b;
    outputs(3324) <= not (a or b);
    outputs(3325) <= b;
    outputs(3326) <= not (a or b);
    outputs(3327) <= b;
    outputs(3328) <= not (a xor b);
    outputs(3329) <= not (a xor b);
    outputs(3330) <= not a;
    outputs(3331) <= a xor b;
    outputs(3332) <= not a or b;
    outputs(3333) <= a xor b;
    outputs(3334) <= not (a xor b);
    outputs(3335) <= a xor b;
    outputs(3336) <= not (a or b);
    outputs(3337) <= a xor b;
    outputs(3338) <= not a;
    outputs(3339) <= a or b;
    outputs(3340) <= a xor b;
    outputs(3341) <= not b;
    outputs(3342) <= a;
    outputs(3343) <= not a;
    outputs(3344) <= not b or a;
    outputs(3345) <= a;
    outputs(3346) <= b;
    outputs(3347) <= not a;
    outputs(3348) <= a or b;
    outputs(3349) <= a xor b;
    outputs(3350) <= a xor b;
    outputs(3351) <= a and not b;
    outputs(3352) <= not a;
    outputs(3353) <= a xor b;
    outputs(3354) <= not a;
    outputs(3355) <= not b;
    outputs(3356) <= a and b;
    outputs(3357) <= not a;
    outputs(3358) <= b;
    outputs(3359) <= not a;
    outputs(3360) <= not a;
    outputs(3361) <= a or b;
    outputs(3362) <= not (a xor b);
    outputs(3363) <= not a;
    outputs(3364) <= not b;
    outputs(3365) <= a xor b;
    outputs(3366) <= a xor b;
    outputs(3367) <= b;
    outputs(3368) <= not (a or b);
    outputs(3369) <= not (a or b);
    outputs(3370) <= not a;
    outputs(3371) <= not (a xor b);
    outputs(3372) <= not b or a;
    outputs(3373) <= a xor b;
    outputs(3374) <= a xor b;
    outputs(3375) <= not a;
    outputs(3376) <= not a;
    outputs(3377) <= b and not a;
    outputs(3378) <= b;
    outputs(3379) <= b and not a;
    outputs(3380) <= not a;
    outputs(3381) <= b;
    outputs(3382) <= not (a xor b);
    outputs(3383) <= not a;
    outputs(3384) <= not a or b;
    outputs(3385) <= a and b;
    outputs(3386) <= a or b;
    outputs(3387) <= a xor b;
    outputs(3388) <= b;
    outputs(3389) <= a xor b;
    outputs(3390) <= b;
    outputs(3391) <= not b or a;
    outputs(3392) <= b;
    outputs(3393) <= a or b;
    outputs(3394) <= a and not b;
    outputs(3395) <= a and b;
    outputs(3396) <= a and not b;
    outputs(3397) <= a;
    outputs(3398) <= not b;
    outputs(3399) <= b;
    outputs(3400) <= not (a xor b);
    outputs(3401) <= b;
    outputs(3402) <= b;
    outputs(3403) <= a and b;
    outputs(3404) <= not b;
    outputs(3405) <= not (a or b);
    outputs(3406) <= not b;
    outputs(3407) <= a;
    outputs(3408) <= b;
    outputs(3409) <= not (a xor b);
    outputs(3410) <= a xor b;
    outputs(3411) <= a xor b;
    outputs(3412) <= not a;
    outputs(3413) <= not b;
    outputs(3414) <= a and b;
    outputs(3415) <= a and not b;
    outputs(3416) <= a;
    outputs(3417) <= not (a xor b);
    outputs(3418) <= not (a or b);
    outputs(3419) <= not a;
    outputs(3420) <= b;
    outputs(3421) <= not a;
    outputs(3422) <= not b;
    outputs(3423) <= b and not a;
    outputs(3424) <= a xor b;
    outputs(3425) <= a xor b;
    outputs(3426) <= not b;
    outputs(3427) <= not (a xor b);
    outputs(3428) <= not a;
    outputs(3429) <= not (a xor b);
    outputs(3430) <= not b or a;
    outputs(3431) <= b;
    outputs(3432) <= b and not a;
    outputs(3433) <= a;
    outputs(3434) <= a and not b;
    outputs(3435) <= not a;
    outputs(3436) <= not (a xor b);
    outputs(3437) <= not b;
    outputs(3438) <= not (a xor b);
    outputs(3439) <= a;
    outputs(3440) <= a xor b;
    outputs(3441) <= b;
    outputs(3442) <= not (a and b);
    outputs(3443) <= a or b;
    outputs(3444) <= a or b;
    outputs(3445) <= a;
    outputs(3446) <= a xor b;
    outputs(3447) <= b;
    outputs(3448) <= not (a and b);
    outputs(3449) <= not (a xor b);
    outputs(3450) <= not b;
    outputs(3451) <= a and not b;
    outputs(3452) <= a xor b;
    outputs(3453) <= not (a xor b);
    outputs(3454) <= a and not b;
    outputs(3455) <= b;
    outputs(3456) <= b;
    outputs(3457) <= not a;
    outputs(3458) <= not (a xor b);
    outputs(3459) <= a xor b;
    outputs(3460) <= not b;
    outputs(3461) <= a and b;
    outputs(3462) <= not a;
    outputs(3463) <= not (a xor b);
    outputs(3464) <= not (a or b);
    outputs(3465) <= not a;
    outputs(3466) <= a xor b;
    outputs(3467) <= not (a xor b);
    outputs(3468) <= not b;
    outputs(3469) <= not b;
    outputs(3470) <= not b or a;
    outputs(3471) <= a xor b;
    outputs(3472) <= not a;
    outputs(3473) <= not (a xor b);
    outputs(3474) <= a and b;
    outputs(3475) <= b;
    outputs(3476) <= b;
    outputs(3477) <= b;
    outputs(3478) <= b;
    outputs(3479) <= not (a xor b);
    outputs(3480) <= not (a or b);
    outputs(3481) <= not a or b;
    outputs(3482) <= b;
    outputs(3483) <= not a or b;
    outputs(3484) <= not b;
    outputs(3485) <= a;
    outputs(3486) <= not b;
    outputs(3487) <= a and not b;
    outputs(3488) <= a;
    outputs(3489) <= b;
    outputs(3490) <= not b;
    outputs(3491) <= b;
    outputs(3492) <= not (a xor b);
    outputs(3493) <= b and not a;
    outputs(3494) <= a and b;
    outputs(3495) <= not a;
    outputs(3496) <= a xor b;
    outputs(3497) <= a or b;
    outputs(3498) <= b and not a;
    outputs(3499) <= a;
    outputs(3500) <= a xor b;
    outputs(3501) <= not a or b;
    outputs(3502) <= b and not a;
    outputs(3503) <= b and not a;
    outputs(3504) <= b;
    outputs(3505) <= not (a xor b);
    outputs(3506) <= a xor b;
    outputs(3507) <= not b;
    outputs(3508) <= not (a xor b);
    outputs(3509) <= not (a xor b);
    outputs(3510) <= not (a and b);
    outputs(3511) <= not a;
    outputs(3512) <= b;
    outputs(3513) <= not (a and b);
    outputs(3514) <= a;
    outputs(3515) <= not b or a;
    outputs(3516) <= not a;
    outputs(3517) <= not (a and b);
    outputs(3518) <= not a;
    outputs(3519) <= not a;
    outputs(3520) <= not a;
    outputs(3521) <= a xor b;
    outputs(3522) <= a and not b;
    outputs(3523) <= not a;
    outputs(3524) <= not a;
    outputs(3525) <= a;
    outputs(3526) <= a;
    outputs(3527) <= a xor b;
    outputs(3528) <= a xor b;
    outputs(3529) <= not (a or b);
    outputs(3530) <= not (a and b);
    outputs(3531) <= not (a xor b);
    outputs(3532) <= not b;
    outputs(3533) <= not (a xor b);
    outputs(3534) <= not (a xor b);
    outputs(3535) <= not b;
    outputs(3536) <= a and b;
    outputs(3537) <= not a;
    outputs(3538) <= a;
    outputs(3539) <= not (a or b);
    outputs(3540) <= a;
    outputs(3541) <= not a;
    outputs(3542) <= b;
    outputs(3543) <= a and not b;
    outputs(3544) <= b and not a;
    outputs(3545) <= not b or a;
    outputs(3546) <= not b;
    outputs(3547) <= a;
    outputs(3548) <= not (a or b);
    outputs(3549) <= not (a and b);
    outputs(3550) <= a xor b;
    outputs(3551) <= not (a xor b);
    outputs(3552) <= not (a xor b);
    outputs(3553) <= not a;
    outputs(3554) <= a xor b;
    outputs(3555) <= not (a xor b);
    outputs(3556) <= not (a xor b);
    outputs(3557) <= not (a xor b);
    outputs(3558) <= not (a and b);
    outputs(3559) <= b and not a;
    outputs(3560) <= not a or b;
    outputs(3561) <= not b;
    outputs(3562) <= not a or b;
    outputs(3563) <= not b or a;
    outputs(3564) <= a and b;
    outputs(3565) <= a xor b;
    outputs(3566) <= b;
    outputs(3567) <= a;
    outputs(3568) <= a;
    outputs(3569) <= a xor b;
    outputs(3570) <= not a;
    outputs(3571) <= b;
    outputs(3572) <= not (a xor b);
    outputs(3573) <= a and b;
    outputs(3574) <= not a;
    outputs(3575) <= b;
    outputs(3576) <= b;
    outputs(3577) <= b;
    outputs(3578) <= b;
    outputs(3579) <= a xor b;
    outputs(3580) <= not (a xor b);
    outputs(3581) <= a and not b;
    outputs(3582) <= not b;
    outputs(3583) <= not (a or b);
    outputs(3584) <= not a;
    outputs(3585) <= a xor b;
    outputs(3586) <= a xor b;
    outputs(3587) <= not (a xor b);
    outputs(3588) <= b and not a;
    outputs(3589) <= not a or b;
    outputs(3590) <= not (a xor b);
    outputs(3591) <= not a;
    outputs(3592) <= a and b;
    outputs(3593) <= not a;
    outputs(3594) <= a xor b;
    outputs(3595) <= not (a xor b);
    outputs(3596) <= b;
    outputs(3597) <= not (a xor b);
    outputs(3598) <= a;
    outputs(3599) <= b;
    outputs(3600) <= a xor b;
    outputs(3601) <= not a;
    outputs(3602) <= a;
    outputs(3603) <= not (a or b);
    outputs(3604) <= not a;
    outputs(3605) <= not a;
    outputs(3606) <= a or b;
    outputs(3607) <= b;
    outputs(3608) <= a and not b;
    outputs(3609) <= not b;
    outputs(3610) <= a xor b;
    outputs(3611) <= not b;
    outputs(3612) <= b;
    outputs(3613) <= not a;
    outputs(3614) <= a xor b;
    outputs(3615) <= a xor b;
    outputs(3616) <= not b;
    outputs(3617) <= a;
    outputs(3618) <= b;
    outputs(3619) <= a;
    outputs(3620) <= not (a xor b);
    outputs(3621) <= not a;
    outputs(3622) <= b;
    outputs(3623) <= not b;
    outputs(3624) <= not (a xor b);
    outputs(3625) <= a or b;
    outputs(3626) <= a and not b;
    outputs(3627) <= not (a xor b);
    outputs(3628) <= not b or a;
    outputs(3629) <= not a;
    outputs(3630) <= b and not a;
    outputs(3631) <= a and b;
    outputs(3632) <= a;
    outputs(3633) <= b and not a;
    outputs(3634) <= not b or a;
    outputs(3635) <= not (a xor b);
    outputs(3636) <= not (a xor b);
    outputs(3637) <= a xor b;
    outputs(3638) <= not (a xor b);
    outputs(3639) <= not (a xor b);
    outputs(3640) <= b and not a;
    outputs(3641) <= b;
    outputs(3642) <= b;
    outputs(3643) <= a;
    outputs(3644) <= not b;
    outputs(3645) <= a;
    outputs(3646) <= not a;
    outputs(3647) <= a xor b;
    outputs(3648) <= not (a or b);
    outputs(3649) <= a and not b;
    outputs(3650) <= not a;
    outputs(3651) <= not b or a;
    outputs(3652) <= not a or b;
    outputs(3653) <= b;
    outputs(3654) <= not b;
    outputs(3655) <= a and not b;
    outputs(3656) <= a;
    outputs(3657) <= a xor b;
    outputs(3658) <= not a;
    outputs(3659) <= a;
    outputs(3660) <= not a;
    outputs(3661) <= not a or b;
    outputs(3662) <= a xor b;
    outputs(3663) <= a;
    outputs(3664) <= a or b;
    outputs(3665) <= not b;
    outputs(3666) <= b;
    outputs(3667) <= a xor b;
    outputs(3668) <= a xor b;
    outputs(3669) <= a xor b;
    outputs(3670) <= not (a xor b);
    outputs(3671) <= not b;
    outputs(3672) <= a xor b;
    outputs(3673) <= not a or b;
    outputs(3674) <= not b or a;
    outputs(3675) <= a and not b;
    outputs(3676) <= a xor b;
    outputs(3677) <= not (a xor b);
    outputs(3678) <= a;
    outputs(3679) <= a;
    outputs(3680) <= not a;
    outputs(3681) <= not (a xor b);
    outputs(3682) <= a and b;
    outputs(3683) <= a;
    outputs(3684) <= b and not a;
    outputs(3685) <= not a or b;
    outputs(3686) <= a or b;
    outputs(3687) <= not (a or b);
    outputs(3688) <= a xor b;
    outputs(3689) <= b;
    outputs(3690) <= not (a or b);
    outputs(3691) <= not a;
    outputs(3692) <= b;
    outputs(3693) <= not (a or b);
    outputs(3694) <= a and b;
    outputs(3695) <= not (a xor b);
    outputs(3696) <= not (a xor b);
    outputs(3697) <= not b or a;
    outputs(3698) <= not (a or b);
    outputs(3699) <= not (a xor b);
    outputs(3700) <= not b;
    outputs(3701) <= not b;
    outputs(3702) <= a;
    outputs(3703) <= not b;
    outputs(3704) <= not b;
    outputs(3705) <= b;
    outputs(3706) <= not (a xor b);
    outputs(3707) <= b;
    outputs(3708) <= b and not a;
    outputs(3709) <= b;
    outputs(3710) <= not b or a;
    outputs(3711) <= b and not a;
    outputs(3712) <= a or b;
    outputs(3713) <= not (a xor b);
    outputs(3714) <= a;
    outputs(3715) <= not a;
    outputs(3716) <= a;
    outputs(3717) <= not a;
    outputs(3718) <= a xor b;
    outputs(3719) <= not a;
    outputs(3720) <= a xor b;
    outputs(3721) <= not (a or b);
    outputs(3722) <= not a;
    outputs(3723) <= a;
    outputs(3724) <= a xor b;
    outputs(3725) <= b and not a;
    outputs(3726) <= a and not b;
    outputs(3727) <= not (a or b);
    outputs(3728) <= not (a xor b);
    outputs(3729) <= a;
    outputs(3730) <= a or b;
    outputs(3731) <= not (a xor b);
    outputs(3732) <= b and not a;
    outputs(3733) <= a xor b;
    outputs(3734) <= not b;
    outputs(3735) <= not b or a;
    outputs(3736) <= not a;
    outputs(3737) <= b and not a;
    outputs(3738) <= a and not b;
    outputs(3739) <= not b;
    outputs(3740) <= not (a or b);
    outputs(3741) <= not a;
    outputs(3742) <= not (a or b);
    outputs(3743) <= a;
    outputs(3744) <= b;
    outputs(3745) <= a or b;
    outputs(3746) <= not b;
    outputs(3747) <= a xor b;
    outputs(3748) <= a;
    outputs(3749) <= not b;
    outputs(3750) <= a and not b;
    outputs(3751) <= a xor b;
    outputs(3752) <= not (a and b);
    outputs(3753) <= b;
    outputs(3754) <= not b;
    outputs(3755) <= a and not b;
    outputs(3756) <= a xor b;
    outputs(3757) <= a xor b;
    outputs(3758) <= not b;
    outputs(3759) <= a and not b;
    outputs(3760) <= a;
    outputs(3761) <= not a;
    outputs(3762) <= b;
    outputs(3763) <= b;
    outputs(3764) <= not (a or b);
    outputs(3765) <= not b;
    outputs(3766) <= not (a or b);
    outputs(3767) <= not b or a;
    outputs(3768) <= not a or b;
    outputs(3769) <= not b;
    outputs(3770) <= a;
    outputs(3771) <= a and not b;
    outputs(3772) <= a xor b;
    outputs(3773) <= a or b;
    outputs(3774) <= b;
    outputs(3775) <= not a;
    outputs(3776) <= b;
    outputs(3777) <= not a;
    outputs(3778) <= a and b;
    outputs(3779) <= not (a and b);
    outputs(3780) <= a xor b;
    outputs(3781) <= not b;
    outputs(3782) <= b;
    outputs(3783) <= a;
    outputs(3784) <= not (a xor b);
    outputs(3785) <= b;
    outputs(3786) <= a xor b;
    outputs(3787) <= a xor b;
    outputs(3788) <= not a;
    outputs(3789) <= not (a or b);
    outputs(3790) <= b;
    outputs(3791) <= a and b;
    outputs(3792) <= a;
    outputs(3793) <= not (a and b);
    outputs(3794) <= not (a and b);
    outputs(3795) <= a;
    outputs(3796) <= not b or a;
    outputs(3797) <= not (a xor b);
    outputs(3798) <= not b or a;
    outputs(3799) <= a xor b;
    outputs(3800) <= not a or b;
    outputs(3801) <= a or b;
    outputs(3802) <= a;
    outputs(3803) <= b;
    outputs(3804) <= a xor b;
    outputs(3805) <= a xor b;
    outputs(3806) <= not b;
    outputs(3807) <= a xor b;
    outputs(3808) <= not b or a;
    outputs(3809) <= a xor b;
    outputs(3810) <= a;
    outputs(3811) <= a and not b;
    outputs(3812) <= not a;
    outputs(3813) <= b;
    outputs(3814) <= not b;
    outputs(3815) <= a or b;
    outputs(3816) <= a xor b;
    outputs(3817) <= not a;
    outputs(3818) <= a xor b;
    outputs(3819) <= not a or b;
    outputs(3820) <= a;
    outputs(3821) <= not (a xor b);
    outputs(3822) <= not a;
    outputs(3823) <= not a;
    outputs(3824) <= not (a xor b);
    outputs(3825) <= a;
    outputs(3826) <= not (a and b);
    outputs(3827) <= a and b;
    outputs(3828) <= b;
    outputs(3829) <= a;
    outputs(3830) <= not b;
    outputs(3831) <= a;
    outputs(3832) <= not a;
    outputs(3833) <= not (a xor b);
    outputs(3834) <= b;
    outputs(3835) <= a and not b;
    outputs(3836) <= not a;
    outputs(3837) <= not b;
    outputs(3838) <= a or b;
    outputs(3839) <= not a;
    outputs(3840) <= not a;
    outputs(3841) <= not a;
    outputs(3842) <= not a;
    outputs(3843) <= b;
    outputs(3844) <= b;
    outputs(3845) <= a or b;
    outputs(3846) <= not a;
    outputs(3847) <= a;
    outputs(3848) <= a xor b;
    outputs(3849) <= b;
    outputs(3850) <= b;
    outputs(3851) <= not a;
    outputs(3852) <= not a;
    outputs(3853) <= not a;
    outputs(3854) <= b and not a;
    outputs(3855) <= not b or a;
    outputs(3856) <= b;
    outputs(3857) <= a xor b;
    outputs(3858) <= b;
    outputs(3859) <= a and not b;
    outputs(3860) <= not a;
    outputs(3861) <= not b;
    outputs(3862) <= a;
    outputs(3863) <= not (a and b);
    outputs(3864) <= a xor b;
    outputs(3865) <= not a;
    outputs(3866) <= b;
    outputs(3867) <= b and not a;
    outputs(3868) <= a;
    outputs(3869) <= b and not a;
    outputs(3870) <= a and not b;
    outputs(3871) <= b;
    outputs(3872) <= not a;
    outputs(3873) <= not b;
    outputs(3874) <= not (a xor b);
    outputs(3875) <= not a;
    outputs(3876) <= a xor b;
    outputs(3877) <= a and b;
    outputs(3878) <= not a;
    outputs(3879) <= b;
    outputs(3880) <= b;
    outputs(3881) <= not (a xor b);
    outputs(3882) <= b;
    outputs(3883) <= not (a xor b);
    outputs(3884) <= a and not b;
    outputs(3885) <= a;
    outputs(3886) <= not b;
    outputs(3887) <= not b;
    outputs(3888) <= not b;
    outputs(3889) <= b;
    outputs(3890) <= not b;
    outputs(3891) <= b and not a;
    outputs(3892) <= not (a xor b);
    outputs(3893) <= not b;
    outputs(3894) <= not (a xor b);
    outputs(3895) <= not b;
    outputs(3896) <= a xor b;
    outputs(3897) <= not (a xor b);
    outputs(3898) <= b;
    outputs(3899) <= not b;
    outputs(3900) <= not (a xor b);
    outputs(3901) <= not a;
    outputs(3902) <= not (a xor b);
    outputs(3903) <= not (a and b);
    outputs(3904) <= not (a or b);
    outputs(3905) <= not (a xor b);
    outputs(3906) <= not b;
    outputs(3907) <= not (a xor b);
    outputs(3908) <= a;
    outputs(3909) <= a or b;
    outputs(3910) <= a xor b;
    outputs(3911) <= b;
    outputs(3912) <= not b or a;
    outputs(3913) <= not (a or b);
    outputs(3914) <= b;
    outputs(3915) <= not a;
    outputs(3916) <= b;
    outputs(3917) <= not b or a;
    outputs(3918) <= b and not a;
    outputs(3919) <= not (a xor b);
    outputs(3920) <= a;
    outputs(3921) <= not b;
    outputs(3922) <= not a;
    outputs(3923) <= b;
    outputs(3924) <= not (a or b);
    outputs(3925) <= a;
    outputs(3926) <= not b;
    outputs(3927) <= not b or a;
    outputs(3928) <= not a;
    outputs(3929) <= not b;
    outputs(3930) <= not (a and b);
    outputs(3931) <= not b;
    outputs(3932) <= not (a or b);
    outputs(3933) <= not b;
    outputs(3934) <= a;
    outputs(3935) <= not (a xor b);
    outputs(3936) <= not (a xor b);
    outputs(3937) <= b and not a;
    outputs(3938) <= b;
    outputs(3939) <= a;
    outputs(3940) <= not b;
    outputs(3941) <= not (a or b);
    outputs(3942) <= not a or b;
    outputs(3943) <= a and b;
    outputs(3944) <= a;
    outputs(3945) <= not a;
    outputs(3946) <= b;
    outputs(3947) <= b;
    outputs(3948) <= not (a or b);
    outputs(3949) <= not b or a;
    outputs(3950) <= not a;
    outputs(3951) <= a xor b;
    outputs(3952) <= b and not a;
    outputs(3953) <= a xor b;
    outputs(3954) <= not a;
    outputs(3955) <= not (a xor b);
    outputs(3956) <= b and not a;
    outputs(3957) <= a;
    outputs(3958) <= not (a xor b);
    outputs(3959) <= not a;
    outputs(3960) <= a and b;
    outputs(3961) <= a;
    outputs(3962) <= a or b;
    outputs(3963) <= not a;
    outputs(3964) <= a xor b;
    outputs(3965) <= not (a or b);
    outputs(3966) <= a or b;
    outputs(3967) <= a and not b;
    outputs(3968) <= not (a and b);
    outputs(3969) <= a and b;
    outputs(3970) <= a xor b;
    outputs(3971) <= b;
    outputs(3972) <= not a;
    outputs(3973) <= a and b;
    outputs(3974) <= not (a xor b);
    outputs(3975) <= not (a or b);
    outputs(3976) <= a and not b;
    outputs(3977) <= not a;
    outputs(3978) <= not (a xor b);
    outputs(3979) <= a and b;
    outputs(3980) <= not a or b;
    outputs(3981) <= not (a xor b);
    outputs(3982) <= a;
    outputs(3983) <= not a;
    outputs(3984) <= b;
    outputs(3985) <= a and not b;
    outputs(3986) <= not b;
    outputs(3987) <= a xor b;
    outputs(3988) <= a xor b;
    outputs(3989) <= a xor b;
    outputs(3990) <= b;
    outputs(3991) <= not a or b;
    outputs(3992) <= b and not a;
    outputs(3993) <= a and not b;
    outputs(3994) <= not (a xor b);
    outputs(3995) <= not b;
    outputs(3996) <= b;
    outputs(3997) <= not b;
    outputs(3998) <= not b;
    outputs(3999) <= a;
    outputs(4000) <= a or b;
    outputs(4001) <= not a;
    outputs(4002) <= not (a xor b);
    outputs(4003) <= a xor b;
    outputs(4004) <= not (a and b);
    outputs(4005) <= b;
    outputs(4006) <= not b;
    outputs(4007) <= b and not a;
    outputs(4008) <= b;
    outputs(4009) <= a and b;
    outputs(4010) <= a;
    outputs(4011) <= a and b;
    outputs(4012) <= b;
    outputs(4013) <= not (a xor b);
    outputs(4014) <= a xor b;
    outputs(4015) <= not (a or b);
    outputs(4016) <= not b;
    outputs(4017) <= not b;
    outputs(4018) <= not b or a;
    outputs(4019) <= b;
    outputs(4020) <= a xor b;
    outputs(4021) <= a or b;
    outputs(4022) <= not a or b;
    outputs(4023) <= a xor b;
    outputs(4024) <= not (a xor b);
    outputs(4025) <= a xor b;
    outputs(4026) <= not b;
    outputs(4027) <= a and not b;
    outputs(4028) <= a;
    outputs(4029) <= a;
    outputs(4030) <= a and not b;
    outputs(4031) <= not (a xor b);
    outputs(4032) <= not (a and b);
    outputs(4033) <= b;
    outputs(4034) <= a and b;
    outputs(4035) <= a;
    outputs(4036) <= not a;
    outputs(4037) <= b;
    outputs(4038) <= not a;
    outputs(4039) <= b;
    outputs(4040) <= not b or a;
    outputs(4041) <= a and b;
    outputs(4042) <= b;
    outputs(4043) <= not (a xor b);
    outputs(4044) <= not (a xor b);
    outputs(4045) <= not b;
    outputs(4046) <= not a or b;
    outputs(4047) <= a;
    outputs(4048) <= not (a xor b);
    outputs(4049) <= not a;
    outputs(4050) <= not a;
    outputs(4051) <= not b or a;
    outputs(4052) <= a and not b;
    outputs(4053) <= a;
    outputs(4054) <= not b or a;
    outputs(4055) <= not a;
    outputs(4056) <= a;
    outputs(4057) <= not (a xor b);
    outputs(4058) <= a xor b;
    outputs(4059) <= a or b;
    outputs(4060) <= not (a and b);
    outputs(4061) <= a or b;
    outputs(4062) <= not (a xor b);
    outputs(4063) <= not (a xor b);
    outputs(4064) <= a or b;
    outputs(4065) <= a or b;
    outputs(4066) <= a;
    outputs(4067) <= not a;
    outputs(4068) <= a or b;
    outputs(4069) <= not b;
    outputs(4070) <= a xor b;
    outputs(4071) <= not b;
    outputs(4072) <= not (a or b);
    outputs(4073) <= not a;
    outputs(4074) <= a xor b;
    outputs(4075) <= not (a and b);
    outputs(4076) <= a or b;
    outputs(4077) <= not (a or b);
    outputs(4078) <= a and b;
    outputs(4079) <= not a or b;
    outputs(4080) <= not a;
    outputs(4081) <= not a;
    outputs(4082) <= b;
    outputs(4083) <= not a or b;
    outputs(4084) <= not a;
    outputs(4085) <= b and not a;
    outputs(4086) <= b;
    outputs(4087) <= a;
    outputs(4088) <= not a;
    outputs(4089) <= not (a or b);
    outputs(4090) <= not a;
    outputs(4091) <= b;
    outputs(4092) <= a;
    outputs(4093) <= not (a xor b);
    outputs(4094) <= a and b;
    outputs(4095) <= not b;
    outputs(4096) <= not a;
    outputs(4097) <= not a;
    outputs(4098) <= not (a xor b);
    outputs(4099) <= a xor b;
    outputs(4100) <= not (a xor b);
    outputs(4101) <= not a;
    outputs(4102) <= b;
    outputs(4103) <= a and not b;
    outputs(4104) <= a and b;
    outputs(4105) <= not (a xor b);
    outputs(4106) <= not (a xor b);
    outputs(4107) <= not (a xor b);
    outputs(4108) <= not a or b;
    outputs(4109) <= not b or a;
    outputs(4110) <= not b;
    outputs(4111) <= b;
    outputs(4112) <= a and b;
    outputs(4113) <= not (a xor b);
    outputs(4114) <= not b;
    outputs(4115) <= not a or b;
    outputs(4116) <= not a;
    outputs(4117) <= not b;
    outputs(4118) <= not b;
    outputs(4119) <= b;
    outputs(4120) <= not (a xor b);
    outputs(4121) <= a;
    outputs(4122) <= not a;
    outputs(4123) <= not a or b;
    outputs(4124) <= not b;
    outputs(4125) <= not a;
    outputs(4126) <= a xor b;
    outputs(4127) <= not a;
    outputs(4128) <= not (a and b);
    outputs(4129) <= b;
    outputs(4130) <= not b;
    outputs(4131) <= a xor b;
    outputs(4132) <= not (a xor b);
    outputs(4133) <= not a;
    outputs(4134) <= b;
    outputs(4135) <= a or b;
    outputs(4136) <= a xor b;
    outputs(4137) <= not b;
    outputs(4138) <= a;
    outputs(4139) <= not (a xor b);
    outputs(4140) <= not (a xor b);
    outputs(4141) <= b;
    outputs(4142) <= a and b;
    outputs(4143) <= b and not a;
    outputs(4144) <= a xor b;
    outputs(4145) <= b and not a;
    outputs(4146) <= a;
    outputs(4147) <= a;
    outputs(4148) <= b and not a;
    outputs(4149) <= not (a xor b);
    outputs(4150) <= not (a xor b);
    outputs(4151) <= not a;
    outputs(4152) <= not (a xor b);
    outputs(4153) <= a xor b;
    outputs(4154) <= b;
    outputs(4155) <= not b or a;
    outputs(4156) <= b and not a;
    outputs(4157) <= b and not a;
    outputs(4158) <= not a;
    outputs(4159) <= not (a xor b);
    outputs(4160) <= not a;
    outputs(4161) <= not a;
    outputs(4162) <= a xor b;
    outputs(4163) <= not b or a;
    outputs(4164) <= a;
    outputs(4165) <= not (a xor b);
    outputs(4166) <= not a;
    outputs(4167) <= not (a and b);
    outputs(4168) <= not a;
    outputs(4169) <= not b or a;
    outputs(4170) <= not a;
    outputs(4171) <= a;
    outputs(4172) <= a xor b;
    outputs(4173) <= not (a or b);
    outputs(4174) <= not (a xor b);
    outputs(4175) <= a and not b;
    outputs(4176) <= not a;
    outputs(4177) <= not a;
    outputs(4178) <= not b;
    outputs(4179) <= b;
    outputs(4180) <= not (a xor b);
    outputs(4181) <= not b;
    outputs(4182) <= b;
    outputs(4183) <= b and not a;
    outputs(4184) <= not b;
    outputs(4185) <= a and not b;
    outputs(4186) <= not b;
    outputs(4187) <= a and not b;
    outputs(4188) <= b;
    outputs(4189) <= not b;
    outputs(4190) <= a xor b;
    outputs(4191) <= not (a xor b);
    outputs(4192) <= not b;
    outputs(4193) <= b and not a;
    outputs(4194) <= not (a xor b);
    outputs(4195) <= a and b;
    outputs(4196) <= not (a and b);
    outputs(4197) <= not a;
    outputs(4198) <= not (a or b);
    outputs(4199) <= a xor b;
    outputs(4200) <= not (a xor b);
    outputs(4201) <= a;
    outputs(4202) <= a;
    outputs(4203) <= b;
    outputs(4204) <= not b;
    outputs(4205) <= b and not a;
    outputs(4206) <= not b;
    outputs(4207) <= a xor b;
    outputs(4208) <= b and not a;
    outputs(4209) <= not a;
    outputs(4210) <= not (a xor b);
    outputs(4211) <= a;
    outputs(4212) <= not (a xor b);
    outputs(4213) <= b;
    outputs(4214) <= a xor b;
    outputs(4215) <= b;
    outputs(4216) <= not b;
    outputs(4217) <= a;
    outputs(4218) <= a and not b;
    outputs(4219) <= b;
    outputs(4220) <= b;
    outputs(4221) <= not (a xor b);
    outputs(4222) <= b;
    outputs(4223) <= not (a and b);
    outputs(4224) <= not a;
    outputs(4225) <= a and b;
    outputs(4226) <= a;
    outputs(4227) <= not a;
    outputs(4228) <= b;
    outputs(4229) <= not a;
    outputs(4230) <= not a;
    outputs(4231) <= not (a and b);
    outputs(4232) <= b;
    outputs(4233) <= a xor b;
    outputs(4234) <= b;
    outputs(4235) <= not a or b;
    outputs(4236) <= not (a or b);
    outputs(4237) <= not a;
    outputs(4238) <= b and not a;
    outputs(4239) <= not (a xor b);
    outputs(4240) <= a xor b;
    outputs(4241) <= not (a or b);
    outputs(4242) <= not b;
    outputs(4243) <= b;
    outputs(4244) <= not (a xor b);
    outputs(4245) <= not (a xor b);
    outputs(4246) <= a;
    outputs(4247) <= not (a xor b);
    outputs(4248) <= not (a and b);
    outputs(4249) <= a;
    outputs(4250) <= not (a or b);
    outputs(4251) <= not b;
    outputs(4252) <= not (a or b);
    outputs(4253) <= a and not b;
    outputs(4254) <= b;
    outputs(4255) <= a xor b;
    outputs(4256) <= not b;
    outputs(4257) <= b;
    outputs(4258) <= not (a or b);
    outputs(4259) <= b;
    outputs(4260) <= not (a xor b);
    outputs(4261) <= b and not a;
    outputs(4262) <= not (a or b);
    outputs(4263) <= not a or b;
    outputs(4264) <= not (a xor b);
    outputs(4265) <= not (a or b);
    outputs(4266) <= not (a xor b);
    outputs(4267) <= b and not a;
    outputs(4268) <= a xor b;
    outputs(4269) <= not (a or b);
    outputs(4270) <= not b;
    outputs(4271) <= not a;
    outputs(4272) <= not a;
    outputs(4273) <= a;
    outputs(4274) <= not (a xor b);
    outputs(4275) <= not a;
    outputs(4276) <= not b;
    outputs(4277) <= b;
    outputs(4278) <= not b;
    outputs(4279) <= not a;
    outputs(4280) <= b and not a;
    outputs(4281) <= not b;
    outputs(4282) <= not a;
    outputs(4283) <= not (a xor b);
    outputs(4284) <= not (a xor b);
    outputs(4285) <= not a;
    outputs(4286) <= a and not b;
    outputs(4287) <= not (a or b);
    outputs(4288) <= not (a or b);
    outputs(4289) <= not b or a;
    outputs(4290) <= a;
    outputs(4291) <= not a;
    outputs(4292) <= a xor b;
    outputs(4293) <= not b;
    outputs(4294) <= b and not a;
    outputs(4295) <= a and b;
    outputs(4296) <= a;
    outputs(4297) <= not (a xor b);
    outputs(4298) <= not (a or b);
    outputs(4299) <= not a;
    outputs(4300) <= a;
    outputs(4301) <= b;
    outputs(4302) <= b;
    outputs(4303) <= a or b;
    outputs(4304) <= not a;
    outputs(4305) <= a;
    outputs(4306) <= a and not b;
    outputs(4307) <= a and not b;
    outputs(4308) <= a and b;
    outputs(4309) <= not a;
    outputs(4310) <= not b;
    outputs(4311) <= b;
    outputs(4312) <= not (a xor b);
    outputs(4313) <= a and not b;
    outputs(4314) <= not (a or b);
    outputs(4315) <= b;
    outputs(4316) <= a;
    outputs(4317) <= not a;
    outputs(4318) <= a and not b;
    outputs(4319) <= not (a or b);
    outputs(4320) <= b;
    outputs(4321) <= b;
    outputs(4322) <= a xor b;
    outputs(4323) <= a;
    outputs(4324) <= a xor b;
    outputs(4325) <= not b;
    outputs(4326) <= b;
    outputs(4327) <= not (a xor b);
    outputs(4328) <= a;
    outputs(4329) <= not a;
    outputs(4330) <= a xor b;
    outputs(4331) <= a and b;
    outputs(4332) <= not (a xor b);
    outputs(4333) <= a or b;
    outputs(4334) <= a and b;
    outputs(4335) <= a xor b;
    outputs(4336) <= not (a xor b);
    outputs(4337) <= b;
    outputs(4338) <= not b;
    outputs(4339) <= not a;
    outputs(4340) <= a;
    outputs(4341) <= not b;
    outputs(4342) <= not (a or b);
    outputs(4343) <= not b;
    outputs(4344) <= b;
    outputs(4345) <= not (a or b);
    outputs(4346) <= a or b;
    outputs(4347) <= b and not a;
    outputs(4348) <= not (a xor b);
    outputs(4349) <= not a or b;
    outputs(4350) <= a xor b;
    outputs(4351) <= a and not b;
    outputs(4352) <= not a;
    outputs(4353) <= b;
    outputs(4354) <= not a;
    outputs(4355) <= a and not b;
    outputs(4356) <= a xor b;
    outputs(4357) <= b;
    outputs(4358) <= not b;
    outputs(4359) <= not b;
    outputs(4360) <= b;
    outputs(4361) <= a;
    outputs(4362) <= not b;
    outputs(4363) <= a xor b;
    outputs(4364) <= not a;
    outputs(4365) <= a xor b;
    outputs(4366) <= not b;
    outputs(4367) <= not b or a;
    outputs(4368) <= a and b;
    outputs(4369) <= a;
    outputs(4370) <= not b;
    outputs(4371) <= not (a xor b);
    outputs(4372) <= not b or a;
    outputs(4373) <= not (a xor b);
    outputs(4374) <= a;
    outputs(4375) <= not (a xor b);
    outputs(4376) <= b;
    outputs(4377) <= not a;
    outputs(4378) <= a;
    outputs(4379) <= not a or b;
    outputs(4380) <= b;
    outputs(4381) <= not b;
    outputs(4382) <= a xor b;
    outputs(4383) <= a;
    outputs(4384) <= a;
    outputs(4385) <= b;
    outputs(4386) <= not b;
    outputs(4387) <= a xor b;
    outputs(4388) <= b;
    outputs(4389) <= not a;
    outputs(4390) <= not (a xor b);
    outputs(4391) <= b;
    outputs(4392) <= a;
    outputs(4393) <= not a or b;
    outputs(4394) <= not b;
    outputs(4395) <= a;
    outputs(4396) <= not b;
    outputs(4397) <= b;
    outputs(4398) <= not (a xor b);
    outputs(4399) <= a;
    outputs(4400) <= a and b;
    outputs(4401) <= a;
    outputs(4402) <= a and b;
    outputs(4403) <= not b;
    outputs(4404) <= not (a xor b);
    outputs(4405) <= b;
    outputs(4406) <= b and not a;
    outputs(4407) <= not b;
    outputs(4408) <= not (a or b);
    outputs(4409) <= a;
    outputs(4410) <= a;
    outputs(4411) <= not a;
    outputs(4412) <= not a;
    outputs(4413) <= a;
    outputs(4414) <= b;
    outputs(4415) <= not (a xor b);
    outputs(4416) <= b and not a;
    outputs(4417) <= not (a or b);
    outputs(4418) <= a xor b;
    outputs(4419) <= a xor b;
    outputs(4420) <= not b;
    outputs(4421) <= not b;
    outputs(4422) <= not a or b;
    outputs(4423) <= a and not b;
    outputs(4424) <= not (a xor b);
    outputs(4425) <= a xor b;
    outputs(4426) <= not a;
    outputs(4427) <= not a;
    outputs(4428) <= a and not b;
    outputs(4429) <= a;
    outputs(4430) <= not (a xor b);
    outputs(4431) <= b;
    outputs(4432) <= not a;
    outputs(4433) <= not a or b;
    outputs(4434) <= a and b;
    outputs(4435) <= b;
    outputs(4436) <= b;
    outputs(4437) <= not a;
    outputs(4438) <= not (a or b);
    outputs(4439) <= not b;
    outputs(4440) <= not b;
    outputs(4441) <= b and not a;
    outputs(4442) <= not a or b;
    outputs(4443) <= not b;
    outputs(4444) <= a;
    outputs(4445) <= not (a xor b);
    outputs(4446) <= a and not b;
    outputs(4447) <= not (a or b);
    outputs(4448) <= not b;
    outputs(4449) <= a;
    outputs(4450) <= b;
    outputs(4451) <= b;
    outputs(4452) <= b;
    outputs(4453) <= not a;
    outputs(4454) <= a xor b;
    outputs(4455) <= a;
    outputs(4456) <= b and not a;
    outputs(4457) <= not (a or b);
    outputs(4458) <= not (a or b);
    outputs(4459) <= not b or a;
    outputs(4460) <= b;
    outputs(4461) <= a xor b;
    outputs(4462) <= b;
    outputs(4463) <= a;
    outputs(4464) <= not a;
    outputs(4465) <= a;
    outputs(4466) <= not b;
    outputs(4467) <= a or b;
    outputs(4468) <= a and not b;
    outputs(4469) <= not a or b;
    outputs(4470) <= a xor b;
    outputs(4471) <= b;
    outputs(4472) <= not (a xor b);
    outputs(4473) <= b;
    outputs(4474) <= not b;
    outputs(4475) <= not b;
    outputs(4476) <= not (a xor b);
    outputs(4477) <= not a;
    outputs(4478) <= b;
    outputs(4479) <= not b;
    outputs(4480) <= not (a and b);
    outputs(4481) <= not a or b;
    outputs(4482) <= a and not b;
    outputs(4483) <= b;
    outputs(4484) <= not a or b;
    outputs(4485) <= not (a xor b);
    outputs(4486) <= a and b;
    outputs(4487) <= not (a xor b);
    outputs(4488) <= a;
    outputs(4489) <= not (a or b);
    outputs(4490) <= not b;
    outputs(4491) <= b;
    outputs(4492) <= b;
    outputs(4493) <= a;
    outputs(4494) <= a and not b;
    outputs(4495) <= a;
    outputs(4496) <= not a;
    outputs(4497) <= b;
    outputs(4498) <= not b;
    outputs(4499) <= a xor b;
    outputs(4500) <= a or b;
    outputs(4501) <= not b;
    outputs(4502) <= not a;
    outputs(4503) <= a xor b;
    outputs(4504) <= b and not a;
    outputs(4505) <= not b;
    outputs(4506) <= not a;
    outputs(4507) <= not a;
    outputs(4508) <= not b;
    outputs(4509) <= not (a xor b);
    outputs(4510) <= a xor b;
    outputs(4511) <= not (a xor b);
    outputs(4512) <= a xor b;
    outputs(4513) <= not (a xor b);
    outputs(4514) <= b;
    outputs(4515) <= b;
    outputs(4516) <= a;
    outputs(4517) <= a and b;
    outputs(4518) <= not (a or b);
    outputs(4519) <= b;
    outputs(4520) <= a and not b;
    outputs(4521) <= b;
    outputs(4522) <= a and not b;
    outputs(4523) <= b;
    outputs(4524) <= b;
    outputs(4525) <= not b;
    outputs(4526) <= a;
    outputs(4527) <= b and not a;
    outputs(4528) <= a xor b;
    outputs(4529) <= not (a xor b);
    outputs(4530) <= b and not a;
    outputs(4531) <= not a;
    outputs(4532) <= not b;
    outputs(4533) <= not a;
    outputs(4534) <= not a;
    outputs(4535) <= a xor b;
    outputs(4536) <= a xor b;
    outputs(4537) <= not a or b;
    outputs(4538) <= a or b;
    outputs(4539) <= a;
    outputs(4540) <= b;
    outputs(4541) <= a xor b;
    outputs(4542) <= a or b;
    outputs(4543) <= a and b;
    outputs(4544) <= b;
    outputs(4545) <= a xor b;
    outputs(4546) <= not (a or b);
    outputs(4547) <= a;
    outputs(4548) <= a;
    outputs(4549) <= a and not b;
    outputs(4550) <= not b;
    outputs(4551) <= b and not a;
    outputs(4552) <= b;
    outputs(4553) <= not a;
    outputs(4554) <= not (a xor b);
    outputs(4555) <= not a or b;
    outputs(4556) <= a;
    outputs(4557) <= a;
    outputs(4558) <= b;
    outputs(4559) <= a xor b;
    outputs(4560) <= a xor b;
    outputs(4561) <= not (a xor b);
    outputs(4562) <= a;
    outputs(4563) <= not b;
    outputs(4564) <= a;
    outputs(4565) <= not (a or b);
    outputs(4566) <= not (a xor b);
    outputs(4567) <= a and not b;
    outputs(4568) <= a xor b;
    outputs(4569) <= a xor b;
    outputs(4570) <= b;
    outputs(4571) <= a xor b;
    outputs(4572) <= a;
    outputs(4573) <= not a;
    outputs(4574) <= a;
    outputs(4575) <= not (a xor b);
    outputs(4576) <= b;
    outputs(4577) <= not b;
    outputs(4578) <= not b;
    outputs(4579) <= not a;
    outputs(4580) <= not (a xor b);
    outputs(4581) <= b;
    outputs(4582) <= not b;
    outputs(4583) <= a;
    outputs(4584) <= not (a xor b);
    outputs(4585) <= b and not a;
    outputs(4586) <= a and b;
    outputs(4587) <= b;
    outputs(4588) <= not b;
    outputs(4589) <= b;
    outputs(4590) <= not b;
    outputs(4591) <= not (a and b);
    outputs(4592) <= not (a and b);
    outputs(4593) <= not (a xor b);
    outputs(4594) <= not a;
    outputs(4595) <= not (a xor b);
    outputs(4596) <= b;
    outputs(4597) <= a and b;
    outputs(4598) <= not (a xor b);
    outputs(4599) <= not (a or b);
    outputs(4600) <= b;
    outputs(4601) <= a xor b;
    outputs(4602) <= not (a and b);
    outputs(4603) <= not a;
    outputs(4604) <= b;
    outputs(4605) <= a and b;
    outputs(4606) <= b;
    outputs(4607) <= a and b;
    outputs(4608) <= not (a and b);
    outputs(4609) <= not b or a;
    outputs(4610) <= a;
    outputs(4611) <= b and not a;
    outputs(4612) <= not (a and b);
    outputs(4613) <= not (a xor b);
    outputs(4614) <= not (a or b);
    outputs(4615) <= not (a xor b);
    outputs(4616) <= not b;
    outputs(4617) <= not (a or b);
    outputs(4618) <= b and not a;
    outputs(4619) <= a xor b;
    outputs(4620) <= b;
    outputs(4621) <= not a;
    outputs(4622) <= a;
    outputs(4623) <= not b;
    outputs(4624) <= not (a xor b);
    outputs(4625) <= not a;
    outputs(4626) <= a;
    outputs(4627) <= a or b;
    outputs(4628) <= a and not b;
    outputs(4629) <= not (a or b);
    outputs(4630) <= a and b;
    outputs(4631) <= not a;
    outputs(4632) <= a xor b;
    outputs(4633) <= a and not b;
    outputs(4634) <= not a;
    outputs(4635) <= a;
    outputs(4636) <= a and not b;
    outputs(4637) <= not b or a;
    outputs(4638) <= not b;
    outputs(4639) <= a and b;
    outputs(4640) <= b and not a;
    outputs(4641) <= not a;
    outputs(4642) <= not b;
    outputs(4643) <= not (a xor b);
    outputs(4644) <= b and not a;
    outputs(4645) <= b and not a;
    outputs(4646) <= not a;
    outputs(4647) <= not a;
    outputs(4648) <= b and not a;
    outputs(4649) <= b and not a;
    outputs(4650) <= a and b;
    outputs(4651) <= not (a xor b);
    outputs(4652) <= a and b;
    outputs(4653) <= a xor b;
    outputs(4654) <= not b;
    outputs(4655) <= not (a xor b);
    outputs(4656) <= b;
    outputs(4657) <= a;
    outputs(4658) <= a or b;
    outputs(4659) <= not a;
    outputs(4660) <= not a;
    outputs(4661) <= not a or b;
    outputs(4662) <= a;
    outputs(4663) <= not b;
    outputs(4664) <= a;
    outputs(4665) <= not b;
    outputs(4666) <= not b;
    outputs(4667) <= not b;
    outputs(4668) <= not (a xor b);
    outputs(4669) <= a xor b;
    outputs(4670) <= not a;
    outputs(4671) <= b;
    outputs(4672) <= a xor b;
    outputs(4673) <= a;
    outputs(4674) <= not (a or b);
    outputs(4675) <= not a;
    outputs(4676) <= a;
    outputs(4677) <= not a;
    outputs(4678) <= not (a xor b);
    outputs(4679) <= not a;
    outputs(4680) <= not (a xor b);
    outputs(4681) <= not b;
    outputs(4682) <= b;
    outputs(4683) <= not (a xor b);
    outputs(4684) <= a;
    outputs(4685) <= not (a xor b);
    outputs(4686) <= b;
    outputs(4687) <= a and b;
    outputs(4688) <= not (a and b);
    outputs(4689) <= not (a or b);
    outputs(4690) <= a xor b;
    outputs(4691) <= a;
    outputs(4692) <= a or b;
    outputs(4693) <= b;
    outputs(4694) <= a;
    outputs(4695) <= a and not b;
    outputs(4696) <= a xor b;
    outputs(4697) <= b and not a;
    outputs(4698) <= not a;
    outputs(4699) <= not (a xor b);
    outputs(4700) <= a xor b;
    outputs(4701) <= not (a or b);
    outputs(4702) <= a and not b;
    outputs(4703) <= a;
    outputs(4704) <= not b;
    outputs(4705) <= b and not a;
    outputs(4706) <= a;
    outputs(4707) <= b;
    outputs(4708) <= not a;
    outputs(4709) <= not a;
    outputs(4710) <= a;
    outputs(4711) <= not a;
    outputs(4712) <= not a;
    outputs(4713) <= a xor b;
    outputs(4714) <= not a;
    outputs(4715) <= a and b;
    outputs(4716) <= a and not b;
    outputs(4717) <= not (a xor b);
    outputs(4718) <= a xor b;
    outputs(4719) <= not b;
    outputs(4720) <= not (a xor b);
    outputs(4721) <= a and b;
    outputs(4722) <= b;
    outputs(4723) <= a;
    outputs(4724) <= not a;
    outputs(4725) <= not b;
    outputs(4726) <= not a;
    outputs(4727) <= not (a xor b);
    outputs(4728) <= not a;
    outputs(4729) <= a;
    outputs(4730) <= not a;
    outputs(4731) <= a and not b;
    outputs(4732) <= not (a xor b);
    outputs(4733) <= a xor b;
    outputs(4734) <= a;
    outputs(4735) <= not a;
    outputs(4736) <= a xor b;
    outputs(4737) <= not b;
    outputs(4738) <= b;
    outputs(4739) <= a and b;
    outputs(4740) <= a;
    outputs(4741) <= not (a and b);
    outputs(4742) <= not b;
    outputs(4743) <= a;
    outputs(4744) <= b and not a;
    outputs(4745) <= not b;
    outputs(4746) <= not (a xor b);
    outputs(4747) <= a;
    outputs(4748) <= b;
    outputs(4749) <= a and not b;
    outputs(4750) <= not (a or b);
    outputs(4751) <= a and b;
    outputs(4752) <= not (a or b);
    outputs(4753) <= b and not a;
    outputs(4754) <= a;
    outputs(4755) <= not a;
    outputs(4756) <= not b or a;
    outputs(4757) <= not b;
    outputs(4758) <= not a;
    outputs(4759) <= a xor b;
    outputs(4760) <= b;
    outputs(4761) <= not (a xor b);
    outputs(4762) <= a and b;
    outputs(4763) <= b;
    outputs(4764) <= not b or a;
    outputs(4765) <= a;
    outputs(4766) <= not a or b;
    outputs(4767) <= a xor b;
    outputs(4768) <= b;
    outputs(4769) <= a;
    outputs(4770) <= a;
    outputs(4771) <= not b or a;
    outputs(4772) <= a xor b;
    outputs(4773) <= not (a and b);
    outputs(4774) <= a and b;
    outputs(4775) <= not (a and b);
    outputs(4776) <= b and not a;
    outputs(4777) <= not (a xor b);
    outputs(4778) <= b and not a;
    outputs(4779) <= a;
    outputs(4780) <= not b;
    outputs(4781) <= not (a xor b);
    outputs(4782) <= a and not b;
    outputs(4783) <= a xor b;
    outputs(4784) <= not a;
    outputs(4785) <= a;
    outputs(4786) <= a;
    outputs(4787) <= not a or b;
    outputs(4788) <= not a or b;
    outputs(4789) <= not a;
    outputs(4790) <= a;
    outputs(4791) <= b and not a;
    outputs(4792) <= not a;
    outputs(4793) <= not b;
    outputs(4794) <= not (a xor b);
    outputs(4795) <= b and not a;
    outputs(4796) <= a and not b;
    outputs(4797) <= b;
    outputs(4798) <= a;
    outputs(4799) <= not b or a;
    outputs(4800) <= not (a xor b);
    outputs(4801) <= not b;
    outputs(4802) <= b;
    outputs(4803) <= not a;
    outputs(4804) <= b and not a;
    outputs(4805) <= not a;
    outputs(4806) <= a;
    outputs(4807) <= not (a xor b);
    outputs(4808) <= not a;
    outputs(4809) <= not a;
    outputs(4810) <= not a;
    outputs(4811) <= a xor b;
    outputs(4812) <= not b;
    outputs(4813) <= a;
    outputs(4814) <= b;
    outputs(4815) <= a xor b;
    outputs(4816) <= not (a xor b);
    outputs(4817) <= not a or b;
    outputs(4818) <= not (a xor b);
    outputs(4819) <= a or b;
    outputs(4820) <= b and not a;
    outputs(4821) <= a xor b;
    outputs(4822) <= a;
    outputs(4823) <= not b;
    outputs(4824) <= a xor b;
    outputs(4825) <= a or b;
    outputs(4826) <= a xor b;
    outputs(4827) <= a xor b;
    outputs(4828) <= a xor b;
    outputs(4829) <= a and not b;
    outputs(4830) <= not a;
    outputs(4831) <= b;
    outputs(4832) <= not (a xor b);
    outputs(4833) <= a and not b;
    outputs(4834) <= a;
    outputs(4835) <= a and not b;
    outputs(4836) <= not a;
    outputs(4837) <= a;
    outputs(4838) <= a xor b;
    outputs(4839) <= a and not b;
    outputs(4840) <= a;
    outputs(4841) <= not (a or b);
    outputs(4842) <= b and not a;
    outputs(4843) <= a xor b;
    outputs(4844) <= a;
    outputs(4845) <= b;
    outputs(4846) <= not (a xor b);
    outputs(4847) <= not (a or b);
    outputs(4848) <= b and not a;
    outputs(4849) <= not b;
    outputs(4850) <= a xor b;
    outputs(4851) <= b;
    outputs(4852) <= b;
    outputs(4853) <= a xor b;
    outputs(4854) <= not a or b;
    outputs(4855) <= a;
    outputs(4856) <= not b;
    outputs(4857) <= not (a and b);
    outputs(4858) <= not (a xor b);
    outputs(4859) <= a;
    outputs(4860) <= a;
    outputs(4861) <= b and not a;
    outputs(4862) <= not (a or b);
    outputs(4863) <= a xor b;
    outputs(4864) <= not (a or b);
    outputs(4865) <= not a;
    outputs(4866) <= a;
    outputs(4867) <= not (a xor b);
    outputs(4868) <= a;
    outputs(4869) <= a;
    outputs(4870) <= a xor b;
    outputs(4871) <= a xor b;
    outputs(4872) <= not (a xor b);
    outputs(4873) <= not (a or b);
    outputs(4874) <= not a;
    outputs(4875) <= a xor b;
    outputs(4876) <= not a;
    outputs(4877) <= not a;
    outputs(4878) <= not (a xor b);
    outputs(4879) <= not b;
    outputs(4880) <= not b;
    outputs(4881) <= not (a xor b);
    outputs(4882) <= not a;
    outputs(4883) <= b;
    outputs(4884) <= not a;
    outputs(4885) <= b;
    outputs(4886) <= not a;
    outputs(4887) <= a xor b;
    outputs(4888) <= not (a xor b);
    outputs(4889) <= a and b;
    outputs(4890) <= b;
    outputs(4891) <= a and not b;
    outputs(4892) <= a and not b;
    outputs(4893) <= not b;
    outputs(4894) <= not b;
    outputs(4895) <= a xor b;
    outputs(4896) <= a;
    outputs(4897) <= b;
    outputs(4898) <= b;
    outputs(4899) <= not b;
    outputs(4900) <= not (a xor b);
    outputs(4901) <= not a;
    outputs(4902) <= b;
    outputs(4903) <= a and b;
    outputs(4904) <= a and not b;
    outputs(4905) <= a xor b;
    outputs(4906) <= b;
    outputs(4907) <= b and not a;
    outputs(4908) <= not a;
    outputs(4909) <= a and not b;
    outputs(4910) <= b;
    outputs(4911) <= not (a or b);
    outputs(4912) <= a and not b;
    outputs(4913) <= a and b;
    outputs(4914) <= b;
    outputs(4915) <= not (a xor b);
    outputs(4916) <= not a;
    outputs(4917) <= not a;
    outputs(4918) <= not (a xor b);
    outputs(4919) <= a;
    outputs(4920) <= not (a and b);
    outputs(4921) <= not b;
    outputs(4922) <= a;
    outputs(4923) <= not (a xor b);
    outputs(4924) <= a and b;
    outputs(4925) <= not b;
    outputs(4926) <= a;
    outputs(4927) <= a and b;
    outputs(4928) <= a;
    outputs(4929) <= not a;
    outputs(4930) <= not (a or b);
    outputs(4931) <= a xor b;
    outputs(4932) <= not (a or b);
    outputs(4933) <= b;
    outputs(4934) <= a xor b;
    outputs(4935) <= not a;
    outputs(4936) <= not (a and b);
    outputs(4937) <= a;
    outputs(4938) <= b and not a;
    outputs(4939) <= not (a xor b);
    outputs(4940) <= a;
    outputs(4941) <= b;
    outputs(4942) <= not (a xor b);
    outputs(4943) <= not (a or b);
    outputs(4944) <= not a;
    outputs(4945) <= b and not a;
    outputs(4946) <= not a;
    outputs(4947) <= not (a or b);
    outputs(4948) <= a;
    outputs(4949) <= not b or a;
    outputs(4950) <= a xor b;
    outputs(4951) <= not a;
    outputs(4952) <= not (a or b);
    outputs(4953) <= not b;
    outputs(4954) <= a xor b;
    outputs(4955) <= a and b;
    outputs(4956) <= a xor b;
    outputs(4957) <= not a;
    outputs(4958) <= not b;
    outputs(4959) <= b;
    outputs(4960) <= a xor b;
    outputs(4961) <= not a;
    outputs(4962) <= b and not a;
    outputs(4963) <= not a;
    outputs(4964) <= a and b;
    outputs(4965) <= a and b;
    outputs(4966) <= a xor b;
    outputs(4967) <= not (a or b);
    outputs(4968) <= a and b;
    outputs(4969) <= not b;
    outputs(4970) <= not a;
    outputs(4971) <= a or b;
    outputs(4972) <= not a;
    outputs(4973) <= a xor b;
    outputs(4974) <= not a;
    outputs(4975) <= a xor b;
    outputs(4976) <= not b;
    outputs(4977) <= a and b;
    outputs(4978) <= not (a or b);
    outputs(4979) <= not (a xor b);
    outputs(4980) <= a xor b;
    outputs(4981) <= a and b;
    outputs(4982) <= not b;
    outputs(4983) <= a;
    outputs(4984) <= not a;
    outputs(4985) <= b;
    outputs(4986) <= not (a or b);
    outputs(4987) <= not a;
    outputs(4988) <= not a;
    outputs(4989) <= not (a xor b);
    outputs(4990) <= not (a xor b);
    outputs(4991) <= not b;
    outputs(4992) <= a xor b;
    outputs(4993) <= a;
    outputs(4994) <= not a or b;
    outputs(4995) <= not b;
    outputs(4996) <= a or b;
    outputs(4997) <= not (a or b);
    outputs(4998) <= a xor b;
    outputs(4999) <= b;
    outputs(5000) <= not (a xor b);
    outputs(5001) <= b;
    outputs(5002) <= b and not a;
    outputs(5003) <= not (a xor b);
    outputs(5004) <= a and b;
    outputs(5005) <= not a;
    outputs(5006) <= b and not a;
    outputs(5007) <= not b;
    outputs(5008) <= not b;
    outputs(5009) <= not (a or b);
    outputs(5010) <= not b or a;
    outputs(5011) <= not a;
    outputs(5012) <= not (a xor b);
    outputs(5013) <= a and b;
    outputs(5014) <= a;
    outputs(5015) <= a;
    outputs(5016) <= b;
    outputs(5017) <= a and not b;
    outputs(5018) <= not (a xor b);
    outputs(5019) <= a and b;
    outputs(5020) <= not (a or b);
    outputs(5021) <= not a;
    outputs(5022) <= a or b;
    outputs(5023) <= not b;
    outputs(5024) <= a and b;
    outputs(5025) <= a xor b;
    outputs(5026) <= not a or b;
    outputs(5027) <= a or b;
    outputs(5028) <= not (a xor b);
    outputs(5029) <= not (a or b);
    outputs(5030) <= b;
    outputs(5031) <= not (a xor b);
    outputs(5032) <= a and b;
    outputs(5033) <= a;
    outputs(5034) <= b;
    outputs(5035) <= not (a xor b);
    outputs(5036) <= not (a xor b);
    outputs(5037) <= not (a xor b);
    outputs(5038) <= a and not b;
    outputs(5039) <= a xor b;
    outputs(5040) <= a xor b;
    outputs(5041) <= not a;
    outputs(5042) <= not b;
    outputs(5043) <= not (a xor b);
    outputs(5044) <= a xor b;
    outputs(5045) <= not a;
    outputs(5046) <= a;
    outputs(5047) <= not a;
    outputs(5048) <= not (a and b);
    outputs(5049) <= a or b;
    outputs(5050) <= not (a xor b);
    outputs(5051) <= not (a xor b);
    outputs(5052) <= a;
    outputs(5053) <= not (a xor b);
    outputs(5054) <= not (a xor b);
    outputs(5055) <= not a;
    outputs(5056) <= not a;
    outputs(5057) <= b and not a;
    outputs(5058) <= not b;
    outputs(5059) <= b;
    outputs(5060) <= b;
    outputs(5061) <= a and b;
    outputs(5062) <= not a;
    outputs(5063) <= a xor b;
    outputs(5064) <= a xor b;
    outputs(5065) <= not (a xor b);
    outputs(5066) <= a xor b;
    outputs(5067) <= not a;
    outputs(5068) <= not b;
    outputs(5069) <= not a;
    outputs(5070) <= not a;
    outputs(5071) <= not (a and b);
    outputs(5072) <= not a;
    outputs(5073) <= a;
    outputs(5074) <= not a;
    outputs(5075) <= b and not a;
    outputs(5076) <= a;
    outputs(5077) <= not (a or b);
    outputs(5078) <= a;
    outputs(5079) <= a or b;
    outputs(5080) <= a and not b;
    outputs(5081) <= a;
    outputs(5082) <= not a;
    outputs(5083) <= not (a xor b);
    outputs(5084) <= a;
    outputs(5085) <= not a;
    outputs(5086) <= a;
    outputs(5087) <= not (a xor b);
    outputs(5088) <= not (a xor b);
    outputs(5089) <= a;
    outputs(5090) <= b and not a;
    outputs(5091) <= not (a or b);
    outputs(5092) <= b;
    outputs(5093) <= a and b;
    outputs(5094) <= not b;
    outputs(5095) <= a and b;
    outputs(5096) <= b;
    outputs(5097) <= not a;
    outputs(5098) <= not (a xor b);
    outputs(5099) <= a and not b;
    outputs(5100) <= a;
    outputs(5101) <= a;
    outputs(5102) <= b and not a;
    outputs(5103) <= not (a xor b);
    outputs(5104) <= not a;
    outputs(5105) <= b;
    outputs(5106) <= a;
    outputs(5107) <= not b;
    outputs(5108) <= a;
    outputs(5109) <= not a;
    outputs(5110) <= a;
    outputs(5111) <= not (a and b);
    outputs(5112) <= a xor b;
    outputs(5113) <= not (a xor b);
    outputs(5114) <= b;
    outputs(5115) <= a xor b;
    outputs(5116) <= a and not b;
    outputs(5117) <= not b;
    outputs(5118) <= a xor b;
    outputs(5119) <= not b;
    outputs(5120) <= a;
    outputs(5121) <= not (a or b);
    outputs(5122) <= b;
    outputs(5123) <= not (a xor b);
    outputs(5124) <= a;
    outputs(5125) <= b;
    outputs(5126) <= a xor b;
    outputs(5127) <= not a;
    outputs(5128) <= b;
    outputs(5129) <= a xor b;
    outputs(5130) <= a xor b;
    outputs(5131) <= b;
    outputs(5132) <= a;
    outputs(5133) <= a xor b;
    outputs(5134) <= not (a xor b);
    outputs(5135) <= a xor b;
    outputs(5136) <= not a;
    outputs(5137) <= a xor b;
    outputs(5138) <= a;
    outputs(5139) <= a;
    outputs(5140) <= a xor b;
    outputs(5141) <= not (a xor b);
    outputs(5142) <= not (a xor b);
    outputs(5143) <= not a or b;
    outputs(5144) <= not b;
    outputs(5145) <= not (a xor b);
    outputs(5146) <= not (a or b);
    outputs(5147) <= not a or b;
    outputs(5148) <= a xor b;
    outputs(5149) <= not a or b;
    outputs(5150) <= not (a xor b);
    outputs(5151) <= not (a and b);
    outputs(5152) <= not a;
    outputs(5153) <= b and not a;
    outputs(5154) <= a xor b;
    outputs(5155) <= not (a xor b);
    outputs(5156) <= not b;
    outputs(5157) <= a xor b;
    outputs(5158) <= not (a or b);
    outputs(5159) <= b;
    outputs(5160) <= not b or a;
    outputs(5161) <= a;
    outputs(5162) <= a;
    outputs(5163) <= a;
    outputs(5164) <= a xor b;
    outputs(5165) <= a;
    outputs(5166) <= not (a xor b);
    outputs(5167) <= not (a xor b);
    outputs(5168) <= not (a xor b);
    outputs(5169) <= b and not a;
    outputs(5170) <= a xor b;
    outputs(5171) <= b;
    outputs(5172) <= b;
    outputs(5173) <= b and not a;
    outputs(5174) <= not (a or b);
    outputs(5175) <= a and b;
    outputs(5176) <= not (a xor b);
    outputs(5177) <= not b or a;
    outputs(5178) <= b and not a;
    outputs(5179) <= not a;
    outputs(5180) <= b;
    outputs(5181) <= b;
    outputs(5182) <= a xor b;
    outputs(5183) <= not (a xor b);
    outputs(5184) <= a and not b;
    outputs(5185) <= not b or a;
    outputs(5186) <= a xor b;
    outputs(5187) <= b;
    outputs(5188) <= not (a or b);
    outputs(5189) <= a;
    outputs(5190) <= not (a xor b);
    outputs(5191) <= not a;
    outputs(5192) <= not (a xor b);
    outputs(5193) <= not b or a;
    outputs(5194) <= a;
    outputs(5195) <= a and b;
    outputs(5196) <= not (a or b);
    outputs(5197) <= a or b;
    outputs(5198) <= not (a xor b);
    outputs(5199) <= a xor b;
    outputs(5200) <= not b;
    outputs(5201) <= not b;
    outputs(5202) <= b;
    outputs(5203) <= a xor b;
    outputs(5204) <= not a;
    outputs(5205) <= not (a and b);
    outputs(5206) <= a;
    outputs(5207) <= not b;
    outputs(5208) <= not a;
    outputs(5209) <= b;
    outputs(5210) <= b;
    outputs(5211) <= not a;
    outputs(5212) <= b;
    outputs(5213) <= a;
    outputs(5214) <= not a;
    outputs(5215) <= a xor b;
    outputs(5216) <= b;
    outputs(5217) <= not (a and b);
    outputs(5218) <= not b;
    outputs(5219) <= a;
    outputs(5220) <= a;
    outputs(5221) <= not (a xor b);
    outputs(5222) <= not a;
    outputs(5223) <= not (a xor b);
    outputs(5224) <= a;
    outputs(5225) <= not b or a;
    outputs(5226) <= not (a xor b);
    outputs(5227) <= a xor b;
    outputs(5228) <= b and not a;
    outputs(5229) <= not (a and b);
    outputs(5230) <= a xor b;
    outputs(5231) <= a xor b;
    outputs(5232) <= not a or b;
    outputs(5233) <= not (a xor b);
    outputs(5234) <= not (a xor b);
    outputs(5235) <= not (a xor b);
    outputs(5236) <= a and not b;
    outputs(5237) <= not (a xor b);
    outputs(5238) <= not b;
    outputs(5239) <= not (a xor b);
    outputs(5240) <= not (a xor b);
    outputs(5241) <= b;
    outputs(5242) <= not b;
    outputs(5243) <= a and not b;
    outputs(5244) <= not (a and b);
    outputs(5245) <= a xor b;
    outputs(5246) <= not (a xor b);
    outputs(5247) <= not (a xor b);
    outputs(5248) <= not (a and b);
    outputs(5249) <= not (a and b);
    outputs(5250) <= a xor b;
    outputs(5251) <= a;
    outputs(5252) <= b;
    outputs(5253) <= not b or a;
    outputs(5254) <= a;
    outputs(5255) <= a xor b;
    outputs(5256) <= b;
    outputs(5257) <= b;
    outputs(5258) <= a;
    outputs(5259) <= not b or a;
    outputs(5260) <= a xor b;
    outputs(5261) <= not (a xor b);
    outputs(5262) <= b;
    outputs(5263) <= a and b;
    outputs(5264) <= a xor b;
    outputs(5265) <= a and b;
    outputs(5266) <= b;
    outputs(5267) <= not (a xor b);
    outputs(5268) <= not (a xor b);
    outputs(5269) <= a xor b;
    outputs(5270) <= b;
    outputs(5271) <= not a;
    outputs(5272) <= not (a xor b);
    outputs(5273) <= not (a and b);
    outputs(5274) <= a xor b;
    outputs(5275) <= not b;
    outputs(5276) <= not (a xor b);
    outputs(5277) <= not (a xor b);
    outputs(5278) <= not b;
    outputs(5279) <= a and b;
    outputs(5280) <= a xor b;
    outputs(5281) <= a or b;
    outputs(5282) <= b;
    outputs(5283) <= b;
    outputs(5284) <= b;
    outputs(5285) <= a xor b;
    outputs(5286) <= a xor b;
    outputs(5287) <= a xor b;
    outputs(5288) <= not a;
    outputs(5289) <= not b or a;
    outputs(5290) <= not (a xor b);
    outputs(5291) <= not b;
    outputs(5292) <= a xor b;
    outputs(5293) <= not b;
    outputs(5294) <= a;
    outputs(5295) <= not a;
    outputs(5296) <= a xor b;
    outputs(5297) <= not a;
    outputs(5298) <= not b;
    outputs(5299) <= a xor b;
    outputs(5300) <= not (a xor b);
    outputs(5301) <= b;
    outputs(5302) <= b and not a;
    outputs(5303) <= not a or b;
    outputs(5304) <= b and not a;
    outputs(5305) <= not b;
    outputs(5306) <= not b;
    outputs(5307) <= not (a xor b);
    outputs(5308) <= a and b;
    outputs(5309) <= not (a and b);
    outputs(5310) <= not a or b;
    outputs(5311) <= a;
    outputs(5312) <= not b;
    outputs(5313) <= not (a xor b);
    outputs(5314) <= a and b;
    outputs(5315) <= a xor b;
    outputs(5316) <= not a or b;
    outputs(5317) <= a xor b;
    outputs(5318) <= b;
    outputs(5319) <= a xor b;
    outputs(5320) <= not b;
    outputs(5321) <= not a;
    outputs(5322) <= b;
    outputs(5323) <= not a;
    outputs(5324) <= a;
    outputs(5325) <= a and not b;
    outputs(5326) <= not (a xor b);
    outputs(5327) <= b;
    outputs(5328) <= a;
    outputs(5329) <= b and not a;
    outputs(5330) <= a and b;
    outputs(5331) <= a;
    outputs(5332) <= not a;
    outputs(5333) <= b;
    outputs(5334) <= a and not b;
    outputs(5335) <= a xor b;
    outputs(5336) <= not a;
    outputs(5337) <= not (a xor b);
    outputs(5338) <= a;
    outputs(5339) <= not a;
    outputs(5340) <= a and not b;
    outputs(5341) <= b and not a;
    outputs(5342) <= not b;
    outputs(5343) <= a xor b;
    outputs(5344) <= not (a xor b);
    outputs(5345) <= not (a xor b);
    outputs(5346) <= a xor b;
    outputs(5347) <= a xor b;
    outputs(5348) <= not (a xor b);
    outputs(5349) <= not a;
    outputs(5350) <= a;
    outputs(5351) <= a and not b;
    outputs(5352) <= a;
    outputs(5353) <= not (a xor b);
    outputs(5354) <= a xor b;
    outputs(5355) <= b;
    outputs(5356) <= a or b;
    outputs(5357) <= a;
    outputs(5358) <= a and b;
    outputs(5359) <= not (a xor b);
    outputs(5360) <= a or b;
    outputs(5361) <= a or b;
    outputs(5362) <= not b;
    outputs(5363) <= a xor b;
    outputs(5364) <= a or b;
    outputs(5365) <= not (a xor b);
    outputs(5366) <= a;
    outputs(5367) <= a xor b;
    outputs(5368) <= a;
    outputs(5369) <= a and b;
    outputs(5370) <= not b;
    outputs(5371) <= not (a xor b);
    outputs(5372) <= not (a xor b);
    outputs(5373) <= not b;
    outputs(5374) <= a;
    outputs(5375) <= a xor b;
    outputs(5376) <= a xor b;
    outputs(5377) <= b;
    outputs(5378) <= b and not a;
    outputs(5379) <= a xor b;
    outputs(5380) <= a;
    outputs(5381) <= not a;
    outputs(5382) <= not a;
    outputs(5383) <= not b;
    outputs(5384) <= a;
    outputs(5385) <= a;
    outputs(5386) <= not b;
    outputs(5387) <= not a;
    outputs(5388) <= not (a or b);
    outputs(5389) <= a xor b;
    outputs(5390) <= b;
    outputs(5391) <= a;
    outputs(5392) <= b;
    outputs(5393) <= b and not a;
    outputs(5394) <= a or b;
    outputs(5395) <= a xor b;
    outputs(5396) <= a xor b;
    outputs(5397) <= a;
    outputs(5398) <= a xor b;
    outputs(5399) <= a xor b;
    outputs(5400) <= b;
    outputs(5401) <= not (a xor b);
    outputs(5402) <= not (a xor b);
    outputs(5403) <= a xor b;
    outputs(5404) <= a xor b;
    outputs(5405) <= not b;
    outputs(5406) <= not (a xor b);
    outputs(5407) <= a;
    outputs(5408) <= not (a xor b);
    outputs(5409) <= not (a xor b);
    outputs(5410) <= a xor b;
    outputs(5411) <= a xor b;
    outputs(5412) <= not (a xor b);
    outputs(5413) <= b;
    outputs(5414) <= not b;
    outputs(5415) <= not (a xor b);
    outputs(5416) <= not (a xor b);
    outputs(5417) <= not (a and b);
    outputs(5418) <= not (a xor b);
    outputs(5419) <= b;
    outputs(5420) <= not a;
    outputs(5421) <= not (a xor b);
    outputs(5422) <= not (a and b);
    outputs(5423) <= a xor b;
    outputs(5424) <= a and b;
    outputs(5425) <= not (a xor b);
    outputs(5426) <= a;
    outputs(5427) <= b;
    outputs(5428) <= not b;
    outputs(5429) <= a xor b;
    outputs(5430) <= not (a or b);
    outputs(5431) <= not (a and b);
    outputs(5432) <= not b;
    outputs(5433) <= not (a xor b);
    outputs(5434) <= not a;
    outputs(5435) <= not b;
    outputs(5436) <= a;
    outputs(5437) <= not b;
    outputs(5438) <= not (a xor b);
    outputs(5439) <= a;
    outputs(5440) <= not b;
    outputs(5441) <= a xor b;
    outputs(5442) <= b;
    outputs(5443) <= a and not b;
    outputs(5444) <= not b;
    outputs(5445) <= not b or a;
    outputs(5446) <= not a;
    outputs(5447) <= b;
    outputs(5448) <= b;
    outputs(5449) <= b;
    outputs(5450) <= a or b;
    outputs(5451) <= a;
    outputs(5452) <= not (a or b);
    outputs(5453) <= b;
    outputs(5454) <= not a;
    outputs(5455) <= not a;
    outputs(5456) <= not a;
    outputs(5457) <= not a or b;
    outputs(5458) <= b;
    outputs(5459) <= a or b;
    outputs(5460) <= not a or b;
    outputs(5461) <= not a;
    outputs(5462) <= not (a xor b);
    outputs(5463) <= b and not a;
    outputs(5464) <= a;
    outputs(5465) <= not a;
    outputs(5466) <= not a;
    outputs(5467) <= a;
    outputs(5468) <= not b;
    outputs(5469) <= not (a and b);
    outputs(5470) <= not a;
    outputs(5471) <= not b;
    outputs(5472) <= not (a xor b);
    outputs(5473) <= b;
    outputs(5474) <= not (a xor b);
    outputs(5475) <= not (a and b);
    outputs(5476) <= a;
    outputs(5477) <= not b;
    outputs(5478) <= b and not a;
    outputs(5479) <= b;
    outputs(5480) <= not (a xor b);
    outputs(5481) <= a xor b;
    outputs(5482) <= not a;
    outputs(5483) <= not (a xor b);
    outputs(5484) <= not (a xor b);
    outputs(5485) <= not (a xor b);
    outputs(5486) <= not a;
    outputs(5487) <= a;
    outputs(5488) <= a xor b;
    outputs(5489) <= a xor b;
    outputs(5490) <= not a;
    outputs(5491) <= a xor b;
    outputs(5492) <= not (a or b);
    outputs(5493) <= a xor b;
    outputs(5494) <= b;
    outputs(5495) <= a xor b;
    outputs(5496) <= not (a and b);
    outputs(5497) <= not b;
    outputs(5498) <= not (a xor b);
    outputs(5499) <= a xor b;
    outputs(5500) <= a and b;
    outputs(5501) <= a xor b;
    outputs(5502) <= b;
    outputs(5503) <= a xor b;
    outputs(5504) <= not b;
    outputs(5505) <= a and not b;
    outputs(5506) <= b;
    outputs(5507) <= a xor b;
    outputs(5508) <= not a or b;
    outputs(5509) <= not (a xor b);
    outputs(5510) <= a;
    outputs(5511) <= not (a or b);
    outputs(5512) <= not a or b;
    outputs(5513) <= not a;
    outputs(5514) <= b;
    outputs(5515) <= not b;
    outputs(5516) <= not a;
    outputs(5517) <= not b;
    outputs(5518) <= a;
    outputs(5519) <= b;
    outputs(5520) <= a xor b;
    outputs(5521) <= b;
    outputs(5522) <= b;
    outputs(5523) <= a xor b;
    outputs(5524) <= b;
    outputs(5525) <= a;
    outputs(5526) <= not b;
    outputs(5527) <= not a;
    outputs(5528) <= a;
    outputs(5529) <= not b;
    outputs(5530) <= a xor b;
    outputs(5531) <= b and not a;
    outputs(5532) <= a or b;
    outputs(5533) <= a xor b;
    outputs(5534) <= not a;
    outputs(5535) <= a;
    outputs(5536) <= a;
    outputs(5537) <= a xor b;
    outputs(5538) <= a xor b;
    outputs(5539) <= a;
    outputs(5540) <= a and not b;
    outputs(5541) <= a xor b;
    outputs(5542) <= a xor b;
    outputs(5543) <= a xor b;
    outputs(5544) <= a xor b;
    outputs(5545) <= not (a or b);
    outputs(5546) <= not b;
    outputs(5547) <= b;
    outputs(5548) <= not (a xor b);
    outputs(5549) <= b;
    outputs(5550) <= not (a xor b);
    outputs(5551) <= a xor b;
    outputs(5552) <= not (a or b);
    outputs(5553) <= not (a xor b);
    outputs(5554) <= a xor b;
    outputs(5555) <= not (a or b);
    outputs(5556) <= not b;
    outputs(5557) <= a xor b;
    outputs(5558) <= b;
    outputs(5559) <= a or b;
    outputs(5560) <= b;
    outputs(5561) <= not (a xor b);
    outputs(5562) <= not (a xor b);
    outputs(5563) <= not (a and b);
    outputs(5564) <= a xor b;
    outputs(5565) <= a;
    outputs(5566) <= not (a xor b);
    outputs(5567) <= a;
    outputs(5568) <= a xor b;
    outputs(5569) <= a xor b;
    outputs(5570) <= not b or a;
    outputs(5571) <= a;
    outputs(5572) <= not a;
    outputs(5573) <= b;
    outputs(5574) <= not (a and b);
    outputs(5575) <= b;
    outputs(5576) <= b;
    outputs(5577) <= not (a xor b);
    outputs(5578) <= a;
    outputs(5579) <= not b;
    outputs(5580) <= b;
    outputs(5581) <= not b;
    outputs(5582) <= a xor b;
    outputs(5583) <= not a or b;
    outputs(5584) <= not (a xor b);
    outputs(5585) <= b;
    outputs(5586) <= not b;
    outputs(5587) <= not (a or b);
    outputs(5588) <= not b;
    outputs(5589) <= a xor b;
    outputs(5590) <= a xor b;
    outputs(5591) <= not (a xor b);
    outputs(5592) <= not (a xor b);
    outputs(5593) <= not (a xor b);
    outputs(5594) <= not (a xor b);
    outputs(5595) <= a xor b;
    outputs(5596) <= a and not b;
    outputs(5597) <= a;
    outputs(5598) <= not b or a;
    outputs(5599) <= not (a xor b);
    outputs(5600) <= a xor b;
    outputs(5601) <= a xor b;
    outputs(5602) <= a xor b;
    outputs(5603) <= a and b;
    outputs(5604) <= a xor b;
    outputs(5605) <= not a;
    outputs(5606) <= not (a xor b);
    outputs(5607) <= not (a or b);
    outputs(5608) <= b;
    outputs(5609) <= not (a xor b);
    outputs(5610) <= not a;
    outputs(5611) <= b;
    outputs(5612) <= b and not a;
    outputs(5613) <= not a;
    outputs(5614) <= not (a or b);
    outputs(5615) <= a;
    outputs(5616) <= a;
    outputs(5617) <= b and not a;
    outputs(5618) <= not (a and b);
    outputs(5619) <= b and not a;
    outputs(5620) <= a and not b;
    outputs(5621) <= b;
    outputs(5622) <= not (a xor b);
    outputs(5623) <= a and not b;
    outputs(5624) <= b;
    outputs(5625) <= a xor b;
    outputs(5626) <= not b;
    outputs(5627) <= not b;
    outputs(5628) <= b;
    outputs(5629) <= a;
    outputs(5630) <= a or b;
    outputs(5631) <= not a;
    outputs(5632) <= b and not a;
    outputs(5633) <= not b;
    outputs(5634) <= not (a xor b);
    outputs(5635) <= a and b;
    outputs(5636) <= not b;
    outputs(5637) <= a xor b;
    outputs(5638) <= a and b;
    outputs(5639) <= not a;
    outputs(5640) <= not a;
    outputs(5641) <= not a;
    outputs(5642) <= not b;
    outputs(5643) <= not b;
    outputs(5644) <= a xor b;
    outputs(5645) <= not (a xor b);
    outputs(5646) <= not b or a;
    outputs(5647) <= b;
    outputs(5648) <= a xor b;
    outputs(5649) <= a xor b;
    outputs(5650) <= a xor b;
    outputs(5651) <= not b;
    outputs(5652) <= a;
    outputs(5653) <= not b;
    outputs(5654) <= not (a or b);
    outputs(5655) <= not b;
    outputs(5656) <= not b;
    outputs(5657) <= a and b;
    outputs(5658) <= a xor b;
    outputs(5659) <= a xor b;
    outputs(5660) <= not (a or b);
    outputs(5661) <= not (a xor b);
    outputs(5662) <= a xor b;
    outputs(5663) <= a or b;
    outputs(5664) <= b and not a;
    outputs(5665) <= b;
    outputs(5666) <= not (a and b);
    outputs(5667) <= not a;
    outputs(5668) <= a xor b;
    outputs(5669) <= not b;
    outputs(5670) <= not (a or b);
    outputs(5671) <= a;
    outputs(5672) <= a xor b;
    outputs(5673) <= a;
    outputs(5674) <= not (a xor b);
    outputs(5675) <= a xor b;
    outputs(5676) <= not a;
    outputs(5677) <= a and b;
    outputs(5678) <= a and b;
    outputs(5679) <= a xor b;
    outputs(5680) <= not b;
    outputs(5681) <= a xor b;
    outputs(5682) <= a;
    outputs(5683) <= not (a xor b);
    outputs(5684) <= a xor b;
    outputs(5685) <= b;
    outputs(5686) <= a and not b;
    outputs(5687) <= b;
    outputs(5688) <= a or b;
    outputs(5689) <= not b;
    outputs(5690) <= not b or a;
    outputs(5691) <= b;
    outputs(5692) <= a;
    outputs(5693) <= a and b;
    outputs(5694) <= not a or b;
    outputs(5695) <= b;
    outputs(5696) <= a;
    outputs(5697) <= a;
    outputs(5698) <= not b or a;
    outputs(5699) <= a xor b;
    outputs(5700) <= not b or a;
    outputs(5701) <= not a or b;
    outputs(5702) <= b and not a;
    outputs(5703) <= a xor b;
    outputs(5704) <= not a;
    outputs(5705) <= not (a or b);
    outputs(5706) <= not b;
    outputs(5707) <= b;
    outputs(5708) <= not (a and b);
    outputs(5709) <= not b;
    outputs(5710) <= not b;
    outputs(5711) <= not a;
    outputs(5712) <= not a;
    outputs(5713) <= a and b;
    outputs(5714) <= not b;
    outputs(5715) <= not (a or b);
    outputs(5716) <= a xor b;
    outputs(5717) <= not b;
    outputs(5718) <= not a;
    outputs(5719) <= not (a xor b);
    outputs(5720) <= not b;
    outputs(5721) <= a xor b;
    outputs(5722) <= not b;
    outputs(5723) <= a xor b;
    outputs(5724) <= not (a xor b);
    outputs(5725) <= b;
    outputs(5726) <= a;
    outputs(5727) <= a xor b;
    outputs(5728) <= a xor b;
    outputs(5729) <= a and b;
    outputs(5730) <= b and not a;
    outputs(5731) <= not b;
    outputs(5732) <= a or b;
    outputs(5733) <= not (a and b);
    outputs(5734) <= not (a xor b);
    outputs(5735) <= not (a xor b);
    outputs(5736) <= a;
    outputs(5737) <= a xor b;
    outputs(5738) <= not b;
    outputs(5739) <= b and not a;
    outputs(5740) <= b and not a;
    outputs(5741) <= a xor b;
    outputs(5742) <= a xor b;
    outputs(5743) <= not (a xor b);
    outputs(5744) <= a xor b;
    outputs(5745) <= not a;
    outputs(5746) <= not b;
    outputs(5747) <= b;
    outputs(5748) <= not (a or b);
    outputs(5749) <= not (a xor b);
    outputs(5750) <= not b;
    outputs(5751) <= not a;
    outputs(5752) <= not (a xor b);
    outputs(5753) <= a;
    outputs(5754) <= b;
    outputs(5755) <= a or b;
    outputs(5756) <= a xor b;
    outputs(5757) <= b and not a;
    outputs(5758) <= not (a or b);
    outputs(5759) <= a xor b;
    outputs(5760) <= a xor b;
    outputs(5761) <= not a;
    outputs(5762) <= not a or b;
    outputs(5763) <= not a or b;
    outputs(5764) <= a xor b;
    outputs(5765) <= b and not a;
    outputs(5766) <= a xor b;
    outputs(5767) <= not (a xor b);
    outputs(5768) <= b;
    outputs(5769) <= b;
    outputs(5770) <= not a;
    outputs(5771) <= not a;
    outputs(5772) <= a and not b;
    outputs(5773) <= b;
    outputs(5774) <= a;
    outputs(5775) <= not a or b;
    outputs(5776) <= not (a and b);
    outputs(5777) <= not a;
    outputs(5778) <= not a or b;
    outputs(5779) <= not a;
    outputs(5780) <= not (a xor b);
    outputs(5781) <= not (a xor b);
    outputs(5782) <= a xor b;
    outputs(5783) <= not (a xor b);
    outputs(5784) <= not a;
    outputs(5785) <= b;
    outputs(5786) <= a xor b;
    outputs(5787) <= a and b;
    outputs(5788) <= not a;
    outputs(5789) <= a xor b;
    outputs(5790) <= not (a xor b);
    outputs(5791) <= not (a xor b);
    outputs(5792) <= not a;
    outputs(5793) <= not b;
    outputs(5794) <= a;
    outputs(5795) <= not a;
    outputs(5796) <= not (a xor b);
    outputs(5797) <= not b;
    outputs(5798) <= not (a xor b);
    outputs(5799) <= not (a xor b);
    outputs(5800) <= a xor b;
    outputs(5801) <= not b;
    outputs(5802) <= b;
    outputs(5803) <= a;
    outputs(5804) <= not (a or b);
    outputs(5805) <= b;
    outputs(5806) <= not (a xor b);
    outputs(5807) <= a and b;
    outputs(5808) <= not (a xor b);
    outputs(5809) <= not b;
    outputs(5810) <= not (a xor b);
    outputs(5811) <= a;
    outputs(5812) <= not (a xor b);
    outputs(5813) <= a and b;
    outputs(5814) <= not (a or b);
    outputs(5815) <= not (a xor b);
    outputs(5816) <= b;
    outputs(5817) <= b and not a;
    outputs(5818) <= not a;
    outputs(5819) <= not (a xor b);
    outputs(5820) <= not a;
    outputs(5821) <= a xor b;
    outputs(5822) <= not b;
    outputs(5823) <= a xor b;
    outputs(5824) <= not (a xor b);
    outputs(5825) <= not (a or b);
    outputs(5826) <= not a or b;
    outputs(5827) <= a;
    outputs(5828) <= a;
    outputs(5829) <= not b;
    outputs(5830) <= not (a xor b);
    outputs(5831) <= a;
    outputs(5832) <= not (a xor b);
    outputs(5833) <= b;
    outputs(5834) <= not (a xor b);
    outputs(5835) <= b;
    outputs(5836) <= b;
    outputs(5837) <= not a;
    outputs(5838) <= b and not a;
    outputs(5839) <= b;
    outputs(5840) <= a and not b;
    outputs(5841) <= not (a or b);
    outputs(5842) <= not b;
    outputs(5843) <= a;
    outputs(5844) <= not (a or b);
    outputs(5845) <= a;
    outputs(5846) <= b;
    outputs(5847) <= a;
    outputs(5848) <= a;
    outputs(5849) <= a and not b;
    outputs(5850) <= a xor b;
    outputs(5851) <= not (a xor b);
    outputs(5852) <= not (a and b);
    outputs(5853) <= a and not b;
    outputs(5854) <= not b;
    outputs(5855) <= not (a xor b);
    outputs(5856) <= not (a xor b);
    outputs(5857) <= not b;
    outputs(5858) <= not b;
    outputs(5859) <= not a;
    outputs(5860) <= a and b;
    outputs(5861) <= not b;
    outputs(5862) <= a xor b;
    outputs(5863) <= a;
    outputs(5864) <= b;
    outputs(5865) <= a xor b;
    outputs(5866) <= a xor b;
    outputs(5867) <= not (a xor b);
    outputs(5868) <= not a or b;
    outputs(5869) <= a xor b;
    outputs(5870) <= not (a or b);
    outputs(5871) <= not a;
    outputs(5872) <= not (a xor b);
    outputs(5873) <= not (a xor b);
    outputs(5874) <= not (a xor b);
    outputs(5875) <= not a;
    outputs(5876) <= not b;
    outputs(5877) <= a xor b;
    outputs(5878) <= not (a and b);
    outputs(5879) <= b and not a;
    outputs(5880) <= a xor b;
    outputs(5881) <= not a;
    outputs(5882) <= a;
    outputs(5883) <= a xor b;
    outputs(5884) <= not a or b;
    outputs(5885) <= a xor b;
    outputs(5886) <= b and not a;
    outputs(5887) <= not a;
    outputs(5888) <= not a or b;
    outputs(5889) <= b;
    outputs(5890) <= b;
    outputs(5891) <= not (a xor b);
    outputs(5892) <= not a;
    outputs(5893) <= a;
    outputs(5894) <= not a or b;
    outputs(5895) <= a;
    outputs(5896) <= not (a xor b);
    outputs(5897) <= a;
    outputs(5898) <= not a or b;
    outputs(5899) <= not a;
    outputs(5900) <= b;
    outputs(5901) <= not (a xor b);
    outputs(5902) <= a xor b;
    outputs(5903) <= not b;
    outputs(5904) <= not b;
    outputs(5905) <= not (a or b);
    outputs(5906) <= a;
    outputs(5907) <= a xor b;
    outputs(5908) <= a xor b;
    outputs(5909) <= b;
    outputs(5910) <= a;
    outputs(5911) <= a;
    outputs(5912) <= not (a xor b);
    outputs(5913) <= not a;
    outputs(5914) <= a and not b;
    outputs(5915) <= not (a and b);
    outputs(5916) <= not (a xor b);
    outputs(5917) <= a;
    outputs(5918) <= a;
    outputs(5919) <= not (a xor b);
    outputs(5920) <= not a;
    outputs(5921) <= a;
    outputs(5922) <= a;
    outputs(5923) <= not a;
    outputs(5924) <= a and b;
    outputs(5925) <= a;
    outputs(5926) <= a xor b;
    outputs(5927) <= b;
    outputs(5928) <= not a;
    outputs(5929) <= a xor b;
    outputs(5930) <= not (a xor b);
    outputs(5931) <= b;
    outputs(5932) <= b;
    outputs(5933) <= not b;
    outputs(5934) <= b;
    outputs(5935) <= a xor b;
    outputs(5936) <= a xor b;
    outputs(5937) <= a xor b;
    outputs(5938) <= not b;
    outputs(5939) <= not b;
    outputs(5940) <= b and not a;
    outputs(5941) <= a xor b;
    outputs(5942) <= not (a and b);
    outputs(5943) <= not a or b;
    outputs(5944) <= not (a or b);
    outputs(5945) <= not (a xor b);
    outputs(5946) <= not b;
    outputs(5947) <= not a or b;
    outputs(5948) <= b;
    outputs(5949) <= not (a xor b);
    outputs(5950) <= not a;
    outputs(5951) <= b;
    outputs(5952) <= not a;
    outputs(5953) <= not a;
    outputs(5954) <= a;
    outputs(5955) <= not (a xor b);
    outputs(5956) <= a xor b;
    outputs(5957) <= b;
    outputs(5958) <= a;
    outputs(5959) <= not (a xor b);
    outputs(5960) <= not a;
    outputs(5961) <= not b or a;
    outputs(5962) <= a xor b;
    outputs(5963) <= not b;
    outputs(5964) <= a;
    outputs(5965) <= not b;
    outputs(5966) <= not b or a;
    outputs(5967) <= b and not a;
    outputs(5968) <= not b;
    outputs(5969) <= not b;
    outputs(5970) <= a xor b;
    outputs(5971) <= a xor b;
    outputs(5972) <= not b or a;
    outputs(5973) <= b;
    outputs(5974) <= not (a xor b);
    outputs(5975) <= b;
    outputs(5976) <= not (a and b);
    outputs(5977) <= a and b;
    outputs(5978) <= a xor b;
    outputs(5979) <= not a or b;
    outputs(5980) <= a;
    outputs(5981) <= not (a xor b);
    outputs(5982) <= not (a xor b);
    outputs(5983) <= a or b;
    outputs(5984) <= a or b;
    outputs(5985) <= not a or b;
    outputs(5986) <= not a;
    outputs(5987) <= a xor b;
    outputs(5988) <= b;
    outputs(5989) <= a;
    outputs(5990) <= a and b;
    outputs(5991) <= not (a xor b);
    outputs(5992) <= not b;
    outputs(5993) <= b;
    outputs(5994) <= not b or a;
    outputs(5995) <= a xor b;
    outputs(5996) <= a;
    outputs(5997) <= not (a xor b);
    outputs(5998) <= b and not a;
    outputs(5999) <= b;
    outputs(6000) <= not a;
    outputs(6001) <= a and not b;
    outputs(6002) <= a;
    outputs(6003) <= a;
    outputs(6004) <= not (a xor b);
    outputs(6005) <= a xor b;
    outputs(6006) <= not (a xor b);
    outputs(6007) <= not (a and b);
    outputs(6008) <= not (a xor b);
    outputs(6009) <= a;
    outputs(6010) <= not (a and b);
    outputs(6011) <= a and b;
    outputs(6012) <= a;
    outputs(6013) <= not a or b;
    outputs(6014) <= not a;
    outputs(6015) <= a;
    outputs(6016) <= a;
    outputs(6017) <= a and not b;
    outputs(6018) <= not (a xor b);
    outputs(6019) <= b and not a;
    outputs(6020) <= not a or b;
    outputs(6021) <= not (a xor b);
    outputs(6022) <= not b;
    outputs(6023) <= a xor b;
    outputs(6024) <= a xor b;
    outputs(6025) <= not a;
    outputs(6026) <= not a;
    outputs(6027) <= a xor b;
    outputs(6028) <= not (a xor b);
    outputs(6029) <= not (a xor b);
    outputs(6030) <= a;
    outputs(6031) <= b;
    outputs(6032) <= not (a xor b);
    outputs(6033) <= b;
    outputs(6034) <= b;
    outputs(6035) <= a and not b;
    outputs(6036) <= not (a or b);
    outputs(6037) <= b;
    outputs(6038) <= not (a or b);
    outputs(6039) <= a xor b;
    outputs(6040) <= not (a xor b);
    outputs(6041) <= not a;
    outputs(6042) <= a;
    outputs(6043) <= not b;
    outputs(6044) <= b and not a;
    outputs(6045) <= a xor b;
    outputs(6046) <= not (a xor b);
    outputs(6047) <= not (a xor b);
    outputs(6048) <= a xor b;
    outputs(6049) <= not a or b;
    outputs(6050) <= a xor b;
    outputs(6051) <= not a;
    outputs(6052) <= not (a xor b);
    outputs(6053) <= b;
    outputs(6054) <= a or b;
    outputs(6055) <= b and not a;
    outputs(6056) <= a or b;
    outputs(6057) <= b;
    outputs(6058) <= a and not b;
    outputs(6059) <= a or b;
    outputs(6060) <= a xor b;
    outputs(6061) <= a and not b;
    outputs(6062) <= not (a xor b);
    outputs(6063) <= not a;
    outputs(6064) <= a and b;
    outputs(6065) <= b;
    outputs(6066) <= not (a or b);
    outputs(6067) <= not b;
    outputs(6068) <= a xor b;
    outputs(6069) <= b;
    outputs(6070) <= a xor b;
    outputs(6071) <= not (a xor b);
    outputs(6072) <= not (a xor b);
    outputs(6073) <= a;
    outputs(6074) <= not a;
    outputs(6075) <= not b;
    outputs(6076) <= a;
    outputs(6077) <= not b;
    outputs(6078) <= not (a xor b);
    outputs(6079) <= a xor b;
    outputs(6080) <= not b;
    outputs(6081) <= b;
    outputs(6082) <= not (a xor b);
    outputs(6083) <= b;
    outputs(6084) <= a xor b;
    outputs(6085) <= not (a xor b);
    outputs(6086) <= not a;
    outputs(6087) <= a xor b;
    outputs(6088) <= a;
    outputs(6089) <= not a;
    outputs(6090) <= not (a or b);
    outputs(6091) <= a;
    outputs(6092) <= not (a or b);
    outputs(6093) <= not (a xor b);
    outputs(6094) <= a xor b;
    outputs(6095) <= not b;
    outputs(6096) <= not (a xor b);
    outputs(6097) <= a or b;
    outputs(6098) <= not b;
    outputs(6099) <= a;
    outputs(6100) <= a and b;
    outputs(6101) <= not a;
    outputs(6102) <= b;
    outputs(6103) <= a xor b;
    outputs(6104) <= a xor b;
    outputs(6105) <= a xor b;
    outputs(6106) <= not b;
    outputs(6107) <= not a or b;
    outputs(6108) <= not b;
    outputs(6109) <= b;
    outputs(6110) <= b;
    outputs(6111) <= not (a or b);
    outputs(6112) <= a;
    outputs(6113) <= not (a xor b);
    outputs(6114) <= a xor b;
    outputs(6115) <= a xor b;
    outputs(6116) <= a xor b;
    outputs(6117) <= a xor b;
    outputs(6118) <= not b;
    outputs(6119) <= not (a or b);
    outputs(6120) <= a xor b;
    outputs(6121) <= not b;
    outputs(6122) <= a xor b;
    outputs(6123) <= a;
    outputs(6124) <= a;
    outputs(6125) <= not b;
    outputs(6126) <= a and b;
    outputs(6127) <= a and not b;
    outputs(6128) <= a and b;
    outputs(6129) <= b;
    outputs(6130) <= a and not b;
    outputs(6131) <= a xor b;
    outputs(6132) <= b;
    outputs(6133) <= b;
    outputs(6134) <= a;
    outputs(6135) <= b;
    outputs(6136) <= a;
    outputs(6137) <= not (a xor b);
    outputs(6138) <= b and not a;
    outputs(6139) <= a xor b;
    outputs(6140) <= a or b;
    outputs(6141) <= a xor b;
    outputs(6142) <= not (a xor b);
    outputs(6143) <= a and b;
    outputs(6144) <= not b or a;
    outputs(6145) <= a xor b;
    outputs(6146) <= a;
    outputs(6147) <= a and not b;
    outputs(6148) <= not (a or b);
    outputs(6149) <= not (a xor b);
    outputs(6150) <= not a;
    outputs(6151) <= not b;
    outputs(6152) <= not (a xor b);
    outputs(6153) <= b and not a;
    outputs(6154) <= not (a xor b);
    outputs(6155) <= not a or b;
    outputs(6156) <= b;
    outputs(6157) <= not a;
    outputs(6158) <= a and b;
    outputs(6159) <= not (a xor b);
    outputs(6160) <= not a;
    outputs(6161) <= a xor b;
    outputs(6162) <= not (a or b);
    outputs(6163) <= a xor b;
    outputs(6164) <= a;
    outputs(6165) <= b;
    outputs(6166) <= a;
    outputs(6167) <= a and b;
    outputs(6168) <= not a;
    outputs(6169) <= not b;
    outputs(6170) <= b;
    outputs(6171) <= not a;
    outputs(6172) <= b;
    outputs(6173) <= not (a xor b);
    outputs(6174) <= not b;
    outputs(6175) <= not (a xor b);
    outputs(6176) <= not (a xor b);
    outputs(6177) <= b;
    outputs(6178) <= b and not a;
    outputs(6179) <= not (a xor b);
    outputs(6180) <= not (a and b);
    outputs(6181) <= a and not b;
    outputs(6182) <= not a;
    outputs(6183) <= a and b;
    outputs(6184) <= b;
    outputs(6185) <= not (a or b);
    outputs(6186) <= b;
    outputs(6187) <= a xor b;
    outputs(6188) <= not (a and b);
    outputs(6189) <= a;
    outputs(6190) <= not a or b;
    outputs(6191) <= not (a xor b);
    outputs(6192) <= not b;
    outputs(6193) <= not (a xor b);
    outputs(6194) <= a;
    outputs(6195) <= not a;
    outputs(6196) <= b;
    outputs(6197) <= not (a or b);
    outputs(6198) <= a xor b;
    outputs(6199) <= a and b;
    outputs(6200) <= not a;
    outputs(6201) <= b;
    outputs(6202) <= not (a or b);
    outputs(6203) <= a;
    outputs(6204) <= not b;
    outputs(6205) <= a xor b;
    outputs(6206) <= not a or b;
    outputs(6207) <= b;
    outputs(6208) <= b and not a;
    outputs(6209) <= a;
    outputs(6210) <= b;
    outputs(6211) <= not (a xor b);
    outputs(6212) <= not (a and b);
    outputs(6213) <= a;
    outputs(6214) <= a and b;
    outputs(6215) <= b and not a;
    outputs(6216) <= a;
    outputs(6217) <= not a;
    outputs(6218) <= b and not a;
    outputs(6219) <= not (a or b);
    outputs(6220) <= b;
    outputs(6221) <= not a;
    outputs(6222) <= not b;
    outputs(6223) <= b;
    outputs(6224) <= not a;
    outputs(6225) <= a;
    outputs(6226) <= b;
    outputs(6227) <= b;
    outputs(6228) <= not (a xor b);
    outputs(6229) <= not a or b;
    outputs(6230) <= b;
    outputs(6231) <= a;
    outputs(6232) <= not (a or b);
    outputs(6233) <= a and b;
    outputs(6234) <= a xor b;
    outputs(6235) <= not b;
    outputs(6236) <= not (a or b);
    outputs(6237) <= not a;
    outputs(6238) <= not a or b;
    outputs(6239) <= a xor b;
    outputs(6240) <= not (a or b);
    outputs(6241) <= not a;
    outputs(6242) <= not (a xor b);
    outputs(6243) <= a and not b;
    outputs(6244) <= not (a or b);
    outputs(6245) <= not b;
    outputs(6246) <= not b;
    outputs(6247) <= not (a xor b);
    outputs(6248) <= b;
    outputs(6249) <= not a;
    outputs(6250) <= not (a and b);
    outputs(6251) <= not a;
    outputs(6252) <= a;
    outputs(6253) <= a;
    outputs(6254) <= not a;
    outputs(6255) <= a xor b;
    outputs(6256) <= not a;
    outputs(6257) <= b;
    outputs(6258) <= a and b;
    outputs(6259) <= a and not b;
    outputs(6260) <= a xor b;
    outputs(6261) <= a xor b;
    outputs(6262) <= not b;
    outputs(6263) <= a and not b;
    outputs(6264) <= a and not b;
    outputs(6265) <= a;
    outputs(6266) <= b and not a;
    outputs(6267) <= not b or a;
    outputs(6268) <= not a;
    outputs(6269) <= a and b;
    outputs(6270) <= not (a or b);
    outputs(6271) <= not a or b;
    outputs(6272) <= not (a xor b);
    outputs(6273) <= a and b;
    outputs(6274) <= b;
    outputs(6275) <= b and not a;
    outputs(6276) <= not a;
    outputs(6277) <= b;
    outputs(6278) <= a xor b;
    outputs(6279) <= a xor b;
    outputs(6280) <= not b;
    outputs(6281) <= a and not b;
    outputs(6282) <= a and b;
    outputs(6283) <= a and b;
    outputs(6284) <= a and b;
    outputs(6285) <= not (a xor b);
    outputs(6286) <= a xor b;
    outputs(6287) <= a;
    outputs(6288) <= a xor b;
    outputs(6289) <= not b or a;
    outputs(6290) <= a xor b;
    outputs(6291) <= not a;
    outputs(6292) <= not (a or b);
    outputs(6293) <= a xor b;
    outputs(6294) <= a and not b;
    outputs(6295) <= a xor b;
    outputs(6296) <= not (a xor b);
    outputs(6297) <= not a or b;
    outputs(6298) <= not a;
    outputs(6299) <= not (a xor b);
    outputs(6300) <= not b;
    outputs(6301) <= a;
    outputs(6302) <= a;
    outputs(6303) <= not b;
    outputs(6304) <= b and not a;
    outputs(6305) <= not (a xor b);
    outputs(6306) <= not a;
    outputs(6307) <= b;
    outputs(6308) <= not a;
    outputs(6309) <= not b;
    outputs(6310) <= not a;
    outputs(6311) <= not b;
    outputs(6312) <= not (a xor b);
    outputs(6313) <= a and not b;
    outputs(6314) <= a and b;
    outputs(6315) <= a;
    outputs(6316) <= not (a or b);
    outputs(6317) <= not b;
    outputs(6318) <= a;
    outputs(6319) <= a xor b;
    outputs(6320) <= a and b;
    outputs(6321) <= a;
    outputs(6322) <= b and not a;
    outputs(6323) <= b and not a;
    outputs(6324) <= not b;
    outputs(6325) <= a;
    outputs(6326) <= not (a and b);
    outputs(6327) <= a and not b;
    outputs(6328) <= a and b;
    outputs(6329) <= not (a xor b);
    outputs(6330) <= not b;
    outputs(6331) <= not a;
    outputs(6332) <= not a;
    outputs(6333) <= b;
    outputs(6334) <= not b;
    outputs(6335) <= not b;
    outputs(6336) <= a and b;
    outputs(6337) <= a xor b;
    outputs(6338) <= not (a xor b);
    outputs(6339) <= not b or a;
    outputs(6340) <= not b or a;
    outputs(6341) <= b;
    outputs(6342) <= not (a xor b);
    outputs(6343) <= b;
    outputs(6344) <= not (a or b);
    outputs(6345) <= not (a and b);
    outputs(6346) <= b;
    outputs(6347) <= not (a xor b);
    outputs(6348) <= b;
    outputs(6349) <= a xor b;
    outputs(6350) <= not a or b;
    outputs(6351) <= not (a xor b);
    outputs(6352) <= a;
    outputs(6353) <= not a;
    outputs(6354) <= a;
    outputs(6355) <= a xor b;
    outputs(6356) <= not b;
    outputs(6357) <= not b;
    outputs(6358) <= a and not b;
    outputs(6359) <= not b;
    outputs(6360) <= b;
    outputs(6361) <= not (a or b);
    outputs(6362) <= a;
    outputs(6363) <= not a or b;
    outputs(6364) <= not (a xor b);
    outputs(6365) <= a;
    outputs(6366) <= not (a xor b);
    outputs(6367) <= a and b;
    outputs(6368) <= a;
    outputs(6369) <= b and not a;
    outputs(6370) <= b and not a;
    outputs(6371) <= a;
    outputs(6372) <= a and not b;
    outputs(6373) <= not (a and b);
    outputs(6374) <= not (a xor b);
    outputs(6375) <= not (a xor b);
    outputs(6376) <= not b or a;
    outputs(6377) <= b;
    outputs(6378) <= not a;
    outputs(6379) <= b;
    outputs(6380) <= not b;
    outputs(6381) <= not b;
    outputs(6382) <= b and not a;
    outputs(6383) <= not (a or b);
    outputs(6384) <= not b or a;
    outputs(6385) <= b and not a;
    outputs(6386) <= a;
    outputs(6387) <= not b;
    outputs(6388) <= b;
    outputs(6389) <= not b;
    outputs(6390) <= not b or a;
    outputs(6391) <= b;
    outputs(6392) <= not (a xor b);
    outputs(6393) <= not b;
    outputs(6394) <= b;
    outputs(6395) <= a and not b;
    outputs(6396) <= a;
    outputs(6397) <= a xor b;
    outputs(6398) <= a and b;
    outputs(6399) <= a and b;
    outputs(6400) <= not b;
    outputs(6401) <= not (a and b);
    outputs(6402) <= a xor b;
    outputs(6403) <= not a;
    outputs(6404) <= b;
    outputs(6405) <= a;
    outputs(6406) <= a xor b;
    outputs(6407) <= b;
    outputs(6408) <= not b;
    outputs(6409) <= not a or b;
    outputs(6410) <= not (a and b);
    outputs(6411) <= a;
    outputs(6412) <= not a;
    outputs(6413) <= not (a xor b);
    outputs(6414) <= b and not a;
    outputs(6415) <= not a or b;
    outputs(6416) <= b and not a;
    outputs(6417) <= a xor b;
    outputs(6418) <= not (a xor b);
    outputs(6419) <= not b;
    outputs(6420) <= a;
    outputs(6421) <= not b;
    outputs(6422) <= not a;
    outputs(6423) <= a;
    outputs(6424) <= not (a and b);
    outputs(6425) <= a;
    outputs(6426) <= a xor b;
    outputs(6427) <= b;
    outputs(6428) <= a and not b;
    outputs(6429) <= not (a xor b);
    outputs(6430) <= not b;
    outputs(6431) <= not (a or b);
    outputs(6432) <= not b;
    outputs(6433) <= a xor b;
    outputs(6434) <= a xor b;
    outputs(6435) <= a and not b;
    outputs(6436) <= a or b;
    outputs(6437) <= b;
    outputs(6438) <= not b;
    outputs(6439) <= a;
    outputs(6440) <= a;
    outputs(6441) <= not a;
    outputs(6442) <= a and not b;
    outputs(6443) <= not b;
    outputs(6444) <= a and not b;
    outputs(6445) <= a xor b;
    outputs(6446) <= b and not a;
    outputs(6447) <= a;
    outputs(6448) <= not (a xor b);
    outputs(6449) <= not b or a;
    outputs(6450) <= not (a and b);
    outputs(6451) <= b;
    outputs(6452) <= a xor b;
    outputs(6453) <= not a;
    outputs(6454) <= not (a xor b);
    outputs(6455) <= b and not a;
    outputs(6456) <= not (a and b);
    outputs(6457) <= not b;
    outputs(6458) <= not a;
    outputs(6459) <= a;
    outputs(6460) <= not b;
    outputs(6461) <= a xor b;
    outputs(6462) <= not b;
    outputs(6463) <= b and not a;
    outputs(6464) <= a and b;
    outputs(6465) <= not (a xor b);
    outputs(6466) <= a;
    outputs(6467) <= b;
    outputs(6468) <= b;
    outputs(6469) <= not (a xor b);
    outputs(6470) <= a;
    outputs(6471) <= a and not b;
    outputs(6472) <= not b or a;
    outputs(6473) <= not b;
    outputs(6474) <= a;
    outputs(6475) <= a xor b;
    outputs(6476) <= a and not b;
    outputs(6477) <= not b;
    outputs(6478) <= not a;
    outputs(6479) <= a and not b;
    outputs(6480) <= not b;
    outputs(6481) <= a xor b;
    outputs(6482) <= not (a or b);
    outputs(6483) <= a and b;
    outputs(6484) <= b;
    outputs(6485) <= a;
    outputs(6486) <= a;
    outputs(6487) <= not b or a;
    outputs(6488) <= a xor b;
    outputs(6489) <= not a;
    outputs(6490) <= a xor b;
    outputs(6491) <= not b;
    outputs(6492) <= a;
    outputs(6493) <= a xor b;
    outputs(6494) <= a;
    outputs(6495) <= b and not a;
    outputs(6496) <= not (a xor b);
    outputs(6497) <= not b;
    outputs(6498) <= not b;
    outputs(6499) <= not a;
    outputs(6500) <= not (a or b);
    outputs(6501) <= not (a xor b);
    outputs(6502) <= a xor b;
    outputs(6503) <= not b;
    outputs(6504) <= a xor b;
    outputs(6505) <= a and b;
    outputs(6506) <= a xor b;
    outputs(6507) <= not b;
    outputs(6508) <= b;
    outputs(6509) <= not (a xor b);
    outputs(6510) <= a;
    outputs(6511) <= not (a or b);
    outputs(6512) <= a;
    outputs(6513) <= b;
    outputs(6514) <= not (a xor b);
    outputs(6515) <= not b;
    outputs(6516) <= not a;
    outputs(6517) <= a and not b;
    outputs(6518) <= not (a xor b);
    outputs(6519) <= b;
    outputs(6520) <= not (a or b);
    outputs(6521) <= a and not b;
    outputs(6522) <= not a;
    outputs(6523) <= a and b;
    outputs(6524) <= not (a xor b);
    outputs(6525) <= b;
    outputs(6526) <= a;
    outputs(6527) <= not (a xor b);
    outputs(6528) <= a and not b;
    outputs(6529) <= a;
    outputs(6530) <= a or b;
    outputs(6531) <= not a;
    outputs(6532) <= a xor b;
    outputs(6533) <= not (a or b);
    outputs(6534) <= b;
    outputs(6535) <= a;
    outputs(6536) <= not (a or b);
    outputs(6537) <= not (a xor b);
    outputs(6538) <= not a;
    outputs(6539) <= b and not a;
    outputs(6540) <= a;
    outputs(6541) <= a;
    outputs(6542) <= b;
    outputs(6543) <= a;
    outputs(6544) <= a or b;
    outputs(6545) <= not (a xor b);
    outputs(6546) <= not (a or b);
    outputs(6547) <= b and not a;
    outputs(6548) <= a and b;
    outputs(6549) <= not (a or b);
    outputs(6550) <= b and not a;
    outputs(6551) <= not (a or b);
    outputs(6552) <= not (a xor b);
    outputs(6553) <= a xor b;
    outputs(6554) <= a xor b;
    outputs(6555) <= not b;
    outputs(6556) <= a xor b;
    outputs(6557) <= a and not b;
    outputs(6558) <= not b;
    outputs(6559) <= not a or b;
    outputs(6560) <= b;
    outputs(6561) <= a;
    outputs(6562) <= not b;
    outputs(6563) <= a;
    outputs(6564) <= not b;
    outputs(6565) <= not (a xor b);
    outputs(6566) <= a and not b;
    outputs(6567) <= not a;
    outputs(6568) <= a;
    outputs(6569) <= a and not b;
    outputs(6570) <= not a;
    outputs(6571) <= not b;
    outputs(6572) <= not b;
    outputs(6573) <= not (a xor b);
    outputs(6574) <= not b;
    outputs(6575) <= a;
    outputs(6576) <= not b;
    outputs(6577) <= not (a xor b);
    outputs(6578) <= a or b;
    outputs(6579) <= not a;
    outputs(6580) <= not a;
    outputs(6581) <= not b;
    outputs(6582) <= not (a xor b);
    outputs(6583) <= not b;
    outputs(6584) <= not (a xor b);
    outputs(6585) <= a xor b;
    outputs(6586) <= not (a xor b);
    outputs(6587) <= a;
    outputs(6588) <= a and b;
    outputs(6589) <= not (a xor b);
    outputs(6590) <= not (a xor b);
    outputs(6591) <= not a;
    outputs(6592) <= a;
    outputs(6593) <= not a or b;
    outputs(6594) <= a xor b;
    outputs(6595) <= a xor b;
    outputs(6596) <= not (a or b);
    outputs(6597) <= a;
    outputs(6598) <= b;
    outputs(6599) <= a;
    outputs(6600) <= not b;
    outputs(6601) <= not b;
    outputs(6602) <= a and b;
    outputs(6603) <= not a;
    outputs(6604) <= a;
    outputs(6605) <= not b;
    outputs(6606) <= a xor b;
    outputs(6607) <= not (a xor b);
    outputs(6608) <= not (a and b);
    outputs(6609) <= b;
    outputs(6610) <= not a;
    outputs(6611) <= a or b;
    outputs(6612) <= not (a xor b);
    outputs(6613) <= not b;
    outputs(6614) <= not b;
    outputs(6615) <= not a;
    outputs(6616) <= not a;
    outputs(6617) <= not b;
    outputs(6618) <= a and b;
    outputs(6619) <= not a;
    outputs(6620) <= b and not a;
    outputs(6621) <= not (a xor b);
    outputs(6622) <= not a;
    outputs(6623) <= a;
    outputs(6624) <= not a;
    outputs(6625) <= not a;
    outputs(6626) <= not a;
    outputs(6627) <= b;
    outputs(6628) <= b;
    outputs(6629) <= not a or b;
    outputs(6630) <= b;
    outputs(6631) <= not a;
    outputs(6632) <= not b;
    outputs(6633) <= not b;
    outputs(6634) <= not a or b;
    outputs(6635) <= not b;
    outputs(6636) <= a and not b;
    outputs(6637) <= a xor b;
    outputs(6638) <= not b;
    outputs(6639) <= b and not a;
    outputs(6640) <= not (a xor b);
    outputs(6641) <= not (a xor b);
    outputs(6642) <= not a;
    outputs(6643) <= a xor b;
    outputs(6644) <= not (a xor b);
    outputs(6645) <= a or b;
    outputs(6646) <= a;
    outputs(6647) <= a and not b;
    outputs(6648) <= not a;
    outputs(6649) <= a xor b;
    outputs(6650) <= b and not a;
    outputs(6651) <= a xor b;
    outputs(6652) <= a;
    outputs(6653) <= not a;
    outputs(6654) <= not a or b;
    outputs(6655) <= not b;
    outputs(6656) <= a;
    outputs(6657) <= not b;
    outputs(6658) <= a;
    outputs(6659) <= a xor b;
    outputs(6660) <= a xor b;
    outputs(6661) <= not a;
    outputs(6662) <= not (a xor b);
    outputs(6663) <= a;
    outputs(6664) <= not (a xor b);
    outputs(6665) <= a and not b;
    outputs(6666) <= b;
    outputs(6667) <= not (a or b);
    outputs(6668) <= not b;
    outputs(6669) <= a xor b;
    outputs(6670) <= not (a xor b);
    outputs(6671) <= a;
    outputs(6672) <= not a;
    outputs(6673) <= a;
    outputs(6674) <= b;
    outputs(6675) <= a xor b;
    outputs(6676) <= not a;
    outputs(6677) <= b;
    outputs(6678) <= not (a or b);
    outputs(6679) <= not (a or b);
    outputs(6680) <= a xor b;
    outputs(6681) <= not a;
    outputs(6682) <= a;
    outputs(6683) <= not (a or b);
    outputs(6684) <= not (a or b);
    outputs(6685) <= b;
    outputs(6686) <= b;
    outputs(6687) <= not (a or b);
    outputs(6688) <= a xor b;
    outputs(6689) <= a;
    outputs(6690) <= not a;
    outputs(6691) <= b;
    outputs(6692) <= b;
    outputs(6693) <= a;
    outputs(6694) <= b;
    outputs(6695) <= not (a xor b);
    outputs(6696) <= a xor b;
    outputs(6697) <= not (a or b);
    outputs(6698) <= not (a xor b);
    outputs(6699) <= b;
    outputs(6700) <= not (a or b);
    outputs(6701) <= a and b;
    outputs(6702) <= not (a and b);
    outputs(6703) <= b and not a;
    outputs(6704) <= a;
    outputs(6705) <= not b;
    outputs(6706) <= b;
    outputs(6707) <= not (a or b);
    outputs(6708) <= not b or a;
    outputs(6709) <= not (a xor b);
    outputs(6710) <= a;
    outputs(6711) <= not (a xor b);
    outputs(6712) <= b;
    outputs(6713) <= a and not b;
    outputs(6714) <= not b or a;
    outputs(6715) <= not b;
    outputs(6716) <= not (a xor b);
    outputs(6717) <= not b;
    outputs(6718) <= not a;
    outputs(6719) <= not a;
    outputs(6720) <= b;
    outputs(6721) <= a or b;
    outputs(6722) <= b and not a;
    outputs(6723) <= not (a or b);
    outputs(6724) <= a;
    outputs(6725) <= not a;
    outputs(6726) <= not a;
    outputs(6727) <= b;
    outputs(6728) <= not a;
    outputs(6729) <= not (a xor b);
    outputs(6730) <= b;
    outputs(6731) <= a;
    outputs(6732) <= b and not a;
    outputs(6733) <= a xor b;
    outputs(6734) <= not (a or b);
    outputs(6735) <= b;
    outputs(6736) <= not a;
    outputs(6737) <= a xor b;
    outputs(6738) <= not a;
    outputs(6739) <= a and not b;
    outputs(6740) <= not b;
    outputs(6741) <= not b;
    outputs(6742) <= a xor b;
    outputs(6743) <= a and not b;
    outputs(6744) <= a;
    outputs(6745) <= b;
    outputs(6746) <= not (a or b);
    outputs(6747) <= a and b;
    outputs(6748) <= not (a xor b);
    outputs(6749) <= not a;
    outputs(6750) <= not a or b;
    outputs(6751) <= not (a xor b);
    outputs(6752) <= not b;
    outputs(6753) <= a and not b;
    outputs(6754) <= not b;
    outputs(6755) <= not (a xor b);
    outputs(6756) <= b and not a;
    outputs(6757) <= not b;
    outputs(6758) <= not b;
    outputs(6759) <= a;
    outputs(6760) <= not (a xor b);
    outputs(6761) <= a xor b;
    outputs(6762) <= b and not a;
    outputs(6763) <= b;
    outputs(6764) <= b;
    outputs(6765) <= not a;
    outputs(6766) <= not (a or b);
    outputs(6767) <= not b or a;
    outputs(6768) <= not b;
    outputs(6769) <= a and b;
    outputs(6770) <= a;
    outputs(6771) <= a and not b;
    outputs(6772) <= a and b;
    outputs(6773) <= not (a xor b);
    outputs(6774) <= a;
    outputs(6775) <= a;
    outputs(6776) <= b;
    outputs(6777) <= not (a xor b);
    outputs(6778) <= not a;
    outputs(6779) <= not b;
    outputs(6780) <= not b;
    outputs(6781) <= not (a xor b);
    outputs(6782) <= not a;
    outputs(6783) <= a and b;
    outputs(6784) <= not a;
    outputs(6785) <= a and b;
    outputs(6786) <= a and b;
    outputs(6787) <= b;
    outputs(6788) <= not a or b;
    outputs(6789) <= b;
    outputs(6790) <= a xor b;
    outputs(6791) <= a xor b;
    outputs(6792) <= a xor b;
    outputs(6793) <= a;
    outputs(6794) <= not (a xor b);
    outputs(6795) <= a or b;
    outputs(6796) <= not a;
    outputs(6797) <= a;
    outputs(6798) <= not (a or b);
    outputs(6799) <= not b;
    outputs(6800) <= a xor b;
    outputs(6801) <= not (a and b);
    outputs(6802) <= not (a xor b);
    outputs(6803) <= not a;
    outputs(6804) <= not b;
    outputs(6805) <= b;
    outputs(6806) <= not a;
    outputs(6807) <= not a or b;
    outputs(6808) <= b;
    outputs(6809) <= b and not a;
    outputs(6810) <= not b;
    outputs(6811) <= not b;
    outputs(6812) <= not b;
    outputs(6813) <= b and not a;
    outputs(6814) <= not a;
    outputs(6815) <= not a or b;
    outputs(6816) <= not b;
    outputs(6817) <= not b;
    outputs(6818) <= b;
    outputs(6819) <= not b;
    outputs(6820) <= not (a and b);
    outputs(6821) <= not (a xor b);
    outputs(6822) <= not (a or b);
    outputs(6823) <= a;
    outputs(6824) <= a;
    outputs(6825) <= not b or a;
    outputs(6826) <= a and not b;
    outputs(6827) <= not (a or b);
    outputs(6828) <= a and b;
    outputs(6829) <= not a;
    outputs(6830) <= a xor b;
    outputs(6831) <= a;
    outputs(6832) <= not (a or b);
    outputs(6833) <= a xor b;
    outputs(6834) <= a xor b;
    outputs(6835) <= a and not b;
    outputs(6836) <= not a;
    outputs(6837) <= b and not a;
    outputs(6838) <= not b;
    outputs(6839) <= not (a xor b);
    outputs(6840) <= not (a xor b);
    outputs(6841) <= a xor b;
    outputs(6842) <= not a;
    outputs(6843) <= not b or a;
    outputs(6844) <= a xor b;
    outputs(6845) <= a;
    outputs(6846) <= not b;
    outputs(6847) <= b;
    outputs(6848) <= a xor b;
    outputs(6849) <= a;
    outputs(6850) <= not a;
    outputs(6851) <= not a;
    outputs(6852) <= not (a xor b);
    outputs(6853) <= not a or b;
    outputs(6854) <= a;
    outputs(6855) <= not b or a;
    outputs(6856) <= a and b;
    outputs(6857) <= not b;
    outputs(6858) <= not b;
    outputs(6859) <= b;
    outputs(6860) <= b;
    outputs(6861) <= a or b;
    outputs(6862) <= a or b;
    outputs(6863) <= a;
    outputs(6864) <= b;
    outputs(6865) <= not (a xor b);
    outputs(6866) <= not (a or b);
    outputs(6867) <= not (a xor b);
    outputs(6868) <= not (a xor b);
    outputs(6869) <= a or b;
    outputs(6870) <= b and not a;
    outputs(6871) <= a or b;
    outputs(6872) <= a xor b;
    outputs(6873) <= not b;
    outputs(6874) <= not (a xor b);
    outputs(6875) <= b;
    outputs(6876) <= a;
    outputs(6877) <= b;
    outputs(6878) <= not a;
    outputs(6879) <= not a;
    outputs(6880) <= not (a xor b);
    outputs(6881) <= not a;
    outputs(6882) <= not b or a;
    outputs(6883) <= not b;
    outputs(6884) <= not (a or b);
    outputs(6885) <= b and not a;
    outputs(6886) <= b;
    outputs(6887) <= a;
    outputs(6888) <= b and not a;
    outputs(6889) <= a or b;
    outputs(6890) <= a xor b;
    outputs(6891) <= b;
    outputs(6892) <= b;
    outputs(6893) <= a or b;
    outputs(6894) <= not a;
    outputs(6895) <= a xor b;
    outputs(6896) <= a xor b;
    outputs(6897) <= a;
    outputs(6898) <= b;
    outputs(6899) <= a;
    outputs(6900) <= not (a xor b);
    outputs(6901) <= not a;
    outputs(6902) <= not (a xor b);
    outputs(6903) <= not b;
    outputs(6904) <= a and b;
    outputs(6905) <= not a;
    outputs(6906) <= not b;
    outputs(6907) <= not b;
    outputs(6908) <= b;
    outputs(6909) <= b and not a;
    outputs(6910) <= not b;
    outputs(6911) <= a and not b;
    outputs(6912) <= not (a xor b);
    outputs(6913) <= not a;
    outputs(6914) <= not a;
    outputs(6915) <= a;
    outputs(6916) <= not b;
    outputs(6917) <= not a;
    outputs(6918) <= not (a xor b);
    outputs(6919) <= b;
    outputs(6920) <= not a or b;
    outputs(6921) <= a;
    outputs(6922) <= not a;
    outputs(6923) <= a or b;
    outputs(6924) <= not b;
    outputs(6925) <= a and b;
    outputs(6926) <= not a or b;
    outputs(6927) <= a or b;
    outputs(6928) <= a and b;
    outputs(6929) <= b;
    outputs(6930) <= a xor b;
    outputs(6931) <= not a;
    outputs(6932) <= not a;
    outputs(6933) <= not b;
    outputs(6934) <= not (a or b);
    outputs(6935) <= not a;
    outputs(6936) <= not b;
    outputs(6937) <= b;
    outputs(6938) <= a xor b;
    outputs(6939) <= b;
    outputs(6940) <= a and not b;
    outputs(6941) <= a xor b;
    outputs(6942) <= a;
    outputs(6943) <= not b;
    outputs(6944) <= a and not b;
    outputs(6945) <= not (a xor b);
    outputs(6946) <= not b;
    outputs(6947) <= a;
    outputs(6948) <= not (a xor b);
    outputs(6949) <= a;
    outputs(6950) <= not (a xor b);
    outputs(6951) <= a and not b;
    outputs(6952) <= a xor b;
    outputs(6953) <= a xor b;
    outputs(6954) <= not (a or b);
    outputs(6955) <= a;
    outputs(6956) <= not (a xor b);
    outputs(6957) <= a;
    outputs(6958) <= a;
    outputs(6959) <= a xor b;
    outputs(6960) <= a and not b;
    outputs(6961) <= a xor b;
    outputs(6962) <= not a;
    outputs(6963) <= a or b;
    outputs(6964) <= not b;
    outputs(6965) <= not (a xor b);
    outputs(6966) <= not a;
    outputs(6967) <= a xor b;
    outputs(6968) <= not b;
    outputs(6969) <= not a;
    outputs(6970) <= not b;
    outputs(6971) <= not (a xor b);
    outputs(6972) <= not (a or b);
    outputs(6973) <= a and not b;
    outputs(6974) <= a or b;
    outputs(6975) <= a xor b;
    outputs(6976) <= b;
    outputs(6977) <= not a or b;
    outputs(6978) <= b;
    outputs(6979) <= not (a or b);
    outputs(6980) <= a and b;
    outputs(6981) <= not a;
    outputs(6982) <= a;
    outputs(6983) <= not b;
    outputs(6984) <= not a or b;
    outputs(6985) <= a and b;
    outputs(6986) <= not (a xor b);
    outputs(6987) <= not (a or b);
    outputs(6988) <= not a;
    outputs(6989) <= a and b;
    outputs(6990) <= a;
    outputs(6991) <= b;
    outputs(6992) <= not a;
    outputs(6993) <= a;
    outputs(6994) <= not b;
    outputs(6995) <= not (a or b);
    outputs(6996) <= not (a or b);
    outputs(6997) <= not (a xor b);
    outputs(6998) <= a;
    outputs(6999) <= a and not b;
    outputs(7000) <= not b;
    outputs(7001) <= a;
    outputs(7002) <= a xor b;
    outputs(7003) <= not (a xor b);
    outputs(7004) <= not b;
    outputs(7005) <= not (a xor b);
    outputs(7006) <= not a;
    outputs(7007) <= not a;
    outputs(7008) <= a xor b;
    outputs(7009) <= not (a xor b);
    outputs(7010) <= not b;
    outputs(7011) <= not a;
    outputs(7012) <= not (a and b);
    outputs(7013) <= not a;
    outputs(7014) <= b;
    outputs(7015) <= not b;
    outputs(7016) <= a and b;
    outputs(7017) <= a;
    outputs(7018) <= a;
    outputs(7019) <= not a;
    outputs(7020) <= not a;
    outputs(7021) <= a xor b;
    outputs(7022) <= not a;
    outputs(7023) <= a;
    outputs(7024) <= a;
    outputs(7025) <= not (a xor b);
    outputs(7026) <= a xor b;
    outputs(7027) <= not a;
    outputs(7028) <= a xor b;
    outputs(7029) <= not b;
    outputs(7030) <= not a;
    outputs(7031) <= a;
    outputs(7032) <= not (a xor b);
    outputs(7033) <= a xor b;
    outputs(7034) <= not (a or b);
    outputs(7035) <= not b or a;
    outputs(7036) <= a or b;
    outputs(7037) <= b;
    outputs(7038) <= b and not a;
    outputs(7039) <= not b or a;
    outputs(7040) <= b and not a;
    outputs(7041) <= not (a xor b);
    outputs(7042) <= b;
    outputs(7043) <= not a;
    outputs(7044) <= a and not b;
    outputs(7045) <= not a;
    outputs(7046) <= not (a xor b);
    outputs(7047) <= not a;
    outputs(7048) <= not a;
    outputs(7049) <= not b or a;
    outputs(7050) <= b;
    outputs(7051) <= a and b;
    outputs(7052) <= not (a xor b);
    outputs(7053) <= b and not a;
    outputs(7054) <= a xor b;
    outputs(7055) <= not (a or b);
    outputs(7056) <= not b;
    outputs(7057) <= not b;
    outputs(7058) <= not a;
    outputs(7059) <= not a;
    outputs(7060) <= a;
    outputs(7061) <= not (a and b);
    outputs(7062) <= not b;
    outputs(7063) <= a;
    outputs(7064) <= not (a and b);
    outputs(7065) <= a;
    outputs(7066) <= not b;
    outputs(7067) <= b and not a;
    outputs(7068) <= not a;
    outputs(7069) <= not a;
    outputs(7070) <= a xor b;
    outputs(7071) <= a;
    outputs(7072) <= not (a and b);
    outputs(7073) <= a;
    outputs(7074) <= not b;
    outputs(7075) <= not a;
    outputs(7076) <= b;
    outputs(7077) <= not (a or b);
    outputs(7078) <= not (a or b);
    outputs(7079) <= not (a or b);
    outputs(7080) <= not (a xor b);
    outputs(7081) <= a;
    outputs(7082) <= not (a xor b);
    outputs(7083) <= b;
    outputs(7084) <= not b;
    outputs(7085) <= not (a xor b);
    outputs(7086) <= a and not b;
    outputs(7087) <= a and not b;
    outputs(7088) <= a xor b;
    outputs(7089) <= b;
    outputs(7090) <= a;
    outputs(7091) <= b;
    outputs(7092) <= b;
    outputs(7093) <= not b or a;
    outputs(7094) <= a;
    outputs(7095) <= a;
    outputs(7096) <= not a;
    outputs(7097) <= not b;
    outputs(7098) <= a and not b;
    outputs(7099) <= a;
    outputs(7100) <= not a or b;
    outputs(7101) <= not b;
    outputs(7102) <= not b;
    outputs(7103) <= a and not b;
    outputs(7104) <= a and not b;
    outputs(7105) <= a;
    outputs(7106) <= not (a xor b);
    outputs(7107) <= a;
    outputs(7108) <= not b;
    outputs(7109) <= not b;
    outputs(7110) <= not b;
    outputs(7111) <= not a;
    outputs(7112) <= not a;
    outputs(7113) <= not (a xor b);
    outputs(7114) <= not (a xor b);
    outputs(7115) <= b;
    outputs(7116) <= a;
    outputs(7117) <= not b;
    outputs(7118) <= not b;
    outputs(7119) <= a and b;
    outputs(7120) <= a xor b;
    outputs(7121) <= not b;
    outputs(7122) <= not a;
    outputs(7123) <= a;
    outputs(7124) <= not (a or b);
    outputs(7125) <= not b or a;
    outputs(7126) <= a and b;
    outputs(7127) <= b and not a;
    outputs(7128) <= a xor b;
    outputs(7129) <= not a;
    outputs(7130) <= not b;
    outputs(7131) <= not (a xor b);
    outputs(7132) <= not a;
    outputs(7133) <= b;
    outputs(7134) <= a;
    outputs(7135) <= not (a or b);
    outputs(7136) <= b;
    outputs(7137) <= b;
    outputs(7138) <= not b;
    outputs(7139) <= a;
    outputs(7140) <= b;
    outputs(7141) <= not b;
    outputs(7142) <= a xor b;
    outputs(7143) <= not b;
    outputs(7144) <= b;
    outputs(7145) <= not a or b;
    outputs(7146) <= not b;
    outputs(7147) <= b;
    outputs(7148) <= a xor b;
    outputs(7149) <= not a;
    outputs(7150) <= not b;
    outputs(7151) <= not (a or b);
    outputs(7152) <= a xor b;
    outputs(7153) <= not b;
    outputs(7154) <= not b;
    outputs(7155) <= b;
    outputs(7156) <= not b or a;
    outputs(7157) <= a and b;
    outputs(7158) <= not a;
    outputs(7159) <= not b;
    outputs(7160) <= not a;
    outputs(7161) <= not a;
    outputs(7162) <= a and b;
    outputs(7163) <= a and b;
    outputs(7164) <= not b;
    outputs(7165) <= a xor b;
    outputs(7166) <= not b;
    outputs(7167) <= not a or b;
    outputs(7168) <= b;
    outputs(7169) <= b;
    outputs(7170) <= a xor b;
    outputs(7171) <= a and not b;
    outputs(7172) <= not b;
    outputs(7173) <= a and b;
    outputs(7174) <= not (a or b);
    outputs(7175) <= not a or b;
    outputs(7176) <= not (a or b);
    outputs(7177) <= not a or b;
    outputs(7178) <= a xor b;
    outputs(7179) <= not a;
    outputs(7180) <= not a;
    outputs(7181) <= a and not b;
    outputs(7182) <= b;
    outputs(7183) <= not a;
    outputs(7184) <= not b;
    outputs(7185) <= a and b;
    outputs(7186) <= a;
    outputs(7187) <= b and not a;
    outputs(7188) <= a;
    outputs(7189) <= a xor b;
    outputs(7190) <= not a or b;
    outputs(7191) <= a and b;
    outputs(7192) <= a and not b;
    outputs(7193) <= a and not b;
    outputs(7194) <= a and not b;
    outputs(7195) <= not a;
    outputs(7196) <= a xor b;
    outputs(7197) <= not a;
    outputs(7198) <= b and not a;
    outputs(7199) <= not b;
    outputs(7200) <= a;
    outputs(7201) <= a xor b;
    outputs(7202) <= a and b;
    outputs(7203) <= a and b;
    outputs(7204) <= a;
    outputs(7205) <= a xor b;
    outputs(7206) <= a and not b;
    outputs(7207) <= not (a xor b);
    outputs(7208) <= a and b;
    outputs(7209) <= b and not a;
    outputs(7210) <= not (a and b);
    outputs(7211) <= a and b;
    outputs(7212) <= not a or b;
    outputs(7213) <= not a;
    outputs(7214) <= not b or a;
    outputs(7215) <= not a;
    outputs(7216) <= b;
    outputs(7217) <= a xor b;
    outputs(7218) <= not (a xor b);
    outputs(7219) <= not (a or b);
    outputs(7220) <= a xor b;
    outputs(7221) <= not a;
    outputs(7222) <= not (a xor b);
    outputs(7223) <= a and not b;
    outputs(7224) <= b;
    outputs(7225) <= b and not a;
    outputs(7226) <= a;
    outputs(7227) <= a;
    outputs(7228) <= not a;
    outputs(7229) <= a;
    outputs(7230) <= not a;
    outputs(7231) <= b;
    outputs(7232) <= not (a or b);
    outputs(7233) <= not a;
    outputs(7234) <= not a;
    outputs(7235) <= a and b;
    outputs(7236) <= a;
    outputs(7237) <= not (a xor b);
    outputs(7238) <= not (a and b);
    outputs(7239) <= not b;
    outputs(7240) <= not b;
    outputs(7241) <= b and not a;
    outputs(7242) <= b and not a;
    outputs(7243) <= not b or a;
    outputs(7244) <= a;
    outputs(7245) <= b;
    outputs(7246) <= not a;
    outputs(7247) <= a xor b;
    outputs(7248) <= a xor b;
    outputs(7249) <= a or b;
    outputs(7250) <= not (a or b);
    outputs(7251) <= a xor b;
    outputs(7252) <= a xor b;
    outputs(7253) <= a xor b;
    outputs(7254) <= not (a xor b);
    outputs(7255) <= a;
    outputs(7256) <= not a;
    outputs(7257) <= not a;
    outputs(7258) <= not b;
    outputs(7259) <= a;
    outputs(7260) <= a;
    outputs(7261) <= not (a or b);
    outputs(7262) <= not b or a;
    outputs(7263) <= a;
    outputs(7264) <= not (a or b);
    outputs(7265) <= a xor b;
    outputs(7266) <= not (a or b);
    outputs(7267) <= a xor b;
    outputs(7268) <= not (a xor b);
    outputs(7269) <= a and b;
    outputs(7270) <= a xor b;
    outputs(7271) <= b;
    outputs(7272) <= not (a or b);
    outputs(7273) <= not (a xor b);
    outputs(7274) <= not (a or b);
    outputs(7275) <= a and not b;
    outputs(7276) <= not (a xor b);
    outputs(7277) <= not b;
    outputs(7278) <= a and not b;
    outputs(7279) <= not (a xor b);
    outputs(7280) <= a xor b;
    outputs(7281) <= b;
    outputs(7282) <= a or b;
    outputs(7283) <= a xor b;
    outputs(7284) <= not (a or b);
    outputs(7285) <= a and not b;
    outputs(7286) <= not a;
    outputs(7287) <= not b;
    outputs(7288) <= b;
    outputs(7289) <= not (a and b);
    outputs(7290) <= not a;
    outputs(7291) <= a and not b;
    outputs(7292) <= not (a or b);
    outputs(7293) <= b and not a;
    outputs(7294) <= not b;
    outputs(7295) <= not a;
    outputs(7296) <= not b;
    outputs(7297) <= a xor b;
    outputs(7298) <= b;
    outputs(7299) <= not a or b;
    outputs(7300) <= not b;
    outputs(7301) <= a;
    outputs(7302) <= b;
    outputs(7303) <= a xor b;
    outputs(7304) <= b;
    outputs(7305) <= not a;
    outputs(7306) <= a xor b;
    outputs(7307) <= a and b;
    outputs(7308) <= a xor b;
    outputs(7309) <= not b;
    outputs(7310) <= b;
    outputs(7311) <= a xor b;
    outputs(7312) <= not (a xor b);
    outputs(7313) <= a xor b;
    outputs(7314) <= a or b;
    outputs(7315) <= a;
    outputs(7316) <= b and not a;
    outputs(7317) <= a xor b;
    outputs(7318) <= a xor b;
    outputs(7319) <= a and not b;
    outputs(7320) <= b;
    outputs(7321) <= a and not b;
    outputs(7322) <= a;
    outputs(7323) <= b;
    outputs(7324) <= not a;
    outputs(7325) <= not a;
    outputs(7326) <= not a;
    outputs(7327) <= a and b;
    outputs(7328) <= b;
    outputs(7329) <= a and b;
    outputs(7330) <= b and not a;
    outputs(7331) <= a;
    outputs(7332) <= a and not b;
    outputs(7333) <= a;
    outputs(7334) <= not a;
    outputs(7335) <= a;
    outputs(7336) <= not a;
    outputs(7337) <= not b;
    outputs(7338) <= a and b;
    outputs(7339) <= a and not b;
    outputs(7340) <= b and not a;
    outputs(7341) <= b and not a;
    outputs(7342) <= a;
    outputs(7343) <= not (a xor b);
    outputs(7344) <= not (a or b);
    outputs(7345) <= a and b;
    outputs(7346) <= a and b;
    outputs(7347) <= not (a or b);
    outputs(7348) <= not (a and b);
    outputs(7349) <= a;
    outputs(7350) <= a xor b;
    outputs(7351) <= a and b;
    outputs(7352) <= a and not b;
    outputs(7353) <= not b;
    outputs(7354) <= not a;
    outputs(7355) <= not (a or b);
    outputs(7356) <= b;
    outputs(7357) <= not a;
    outputs(7358) <= a or b;
    outputs(7359) <= a and b;
    outputs(7360) <= a xor b;
    outputs(7361) <= not a;
    outputs(7362) <= b and not a;
    outputs(7363) <= a;
    outputs(7364) <= not a;
    outputs(7365) <= a and b;
    outputs(7366) <= b;
    outputs(7367) <= not a;
    outputs(7368) <= a and not b;
    outputs(7369) <= not (a xor b);
    outputs(7370) <= a;
    outputs(7371) <= a xor b;
    outputs(7372) <= b;
    outputs(7373) <= b;
    outputs(7374) <= not (a or b);
    outputs(7375) <= a xor b;
    outputs(7376) <= not a;
    outputs(7377) <= not (a xor b);
    outputs(7378) <= a;
    outputs(7379) <= not b;
    outputs(7380) <= not b or a;
    outputs(7381) <= not b;
    outputs(7382) <= not a;
    outputs(7383) <= a and not b;
    outputs(7384) <= not a;
    outputs(7385) <= a;
    outputs(7386) <= a and not b;
    outputs(7387) <= not (a xor b);
    outputs(7388) <= not b;
    outputs(7389) <= b;
    outputs(7390) <= not a;
    outputs(7391) <= a;
    outputs(7392) <= b;
    outputs(7393) <= a and not b;
    outputs(7394) <= a xor b;
    outputs(7395) <= a xor b;
    outputs(7396) <= not b;
    outputs(7397) <= not a;
    outputs(7398) <= not (a xor b);
    outputs(7399) <= not b;
    outputs(7400) <= not a or b;
    outputs(7401) <= not (a xor b);
    outputs(7402) <= not (a xor b);
    outputs(7403) <= not (a or b);
    outputs(7404) <= not b;
    outputs(7405) <= a xor b;
    outputs(7406) <= b and not a;
    outputs(7407) <= not (a xor b);
    outputs(7408) <= not (a xor b);
    outputs(7409) <= a;
    outputs(7410) <= not b;
    outputs(7411) <= not b;
    outputs(7412) <= not (a xor b);
    outputs(7413) <= not (a xor b);
    outputs(7414) <= b;
    outputs(7415) <= not a;
    outputs(7416) <= a;
    outputs(7417) <= not b;
    outputs(7418) <= not (a xor b);
    outputs(7419) <= a xor b;
    outputs(7420) <= b;
    outputs(7421) <= not a;
    outputs(7422) <= not b;
    outputs(7423) <= not b;
    outputs(7424) <= not b or a;
    outputs(7425) <= a;
    outputs(7426) <= a;
    outputs(7427) <= a xor b;
    outputs(7428) <= not a;
    outputs(7429) <= not b;
    outputs(7430) <= b and not a;
    outputs(7431) <= not a;
    outputs(7432) <= not b;
    outputs(7433) <= not (a xor b);
    outputs(7434) <= not (a and b);
    outputs(7435) <= b and not a;
    outputs(7436) <= not a;
    outputs(7437) <= b and not a;
    outputs(7438) <= not b or a;
    outputs(7439) <= a and b;
    outputs(7440) <= a;
    outputs(7441) <= a and not b;
    outputs(7442) <= not (a or b);
    outputs(7443) <= not a;
    outputs(7444) <= not (a or b);
    outputs(7445) <= a;
    outputs(7446) <= not b;
    outputs(7447) <= b;
    outputs(7448) <= a xor b;
    outputs(7449) <= not a;
    outputs(7450) <= not a;
    outputs(7451) <= b;
    outputs(7452) <= not (a xor b);
    outputs(7453) <= a xor b;
    outputs(7454) <= not (a xor b);
    outputs(7455) <= not b or a;
    outputs(7456) <= not a;
    outputs(7457) <= not b;
    outputs(7458) <= not a or b;
    outputs(7459) <= a or b;
    outputs(7460) <= not a;
    outputs(7461) <= not b;
    outputs(7462) <= not (a xor b);
    outputs(7463) <= b;
    outputs(7464) <= a xor b;
    outputs(7465) <= a and not b;
    outputs(7466) <= not b;
    outputs(7467) <= not (a xor b);
    outputs(7468) <= not (a xor b);
    outputs(7469) <= b and not a;
    outputs(7470) <= a;
    outputs(7471) <= a xor b;
    outputs(7472) <= not b;
    outputs(7473) <= not a;
    outputs(7474) <= b and not a;
    outputs(7475) <= not (a xor b);
    outputs(7476) <= a xor b;
    outputs(7477) <= b;
    outputs(7478) <= a;
    outputs(7479) <= a xor b;
    outputs(7480) <= not b;
    outputs(7481) <= b and not a;
    outputs(7482) <= not b;
    outputs(7483) <= a;
    outputs(7484) <= not (a or b);
    outputs(7485) <= not b;
    outputs(7486) <= b;
    outputs(7487) <= not (a and b);
    outputs(7488) <= b;
    outputs(7489) <= not a;
    outputs(7490) <= not (a xor b);
    outputs(7491) <= not (a or b);
    outputs(7492) <= not (a or b);
    outputs(7493) <= a and b;
    outputs(7494) <= a xor b;
    outputs(7495) <= a and b;
    outputs(7496) <= a and not b;
    outputs(7497) <= not (a xor b);
    outputs(7498) <= a xor b;
    outputs(7499) <= b and not a;
    outputs(7500) <= not (a xor b);
    outputs(7501) <= not (a xor b);
    outputs(7502) <= b;
    outputs(7503) <= a;
    outputs(7504) <= not a;
    outputs(7505) <= not a;
    outputs(7506) <= a xor b;
    outputs(7507) <= a and not b;
    outputs(7508) <= b;
    outputs(7509) <= a or b;
    outputs(7510) <= a;
    outputs(7511) <= a and b;
    outputs(7512) <= a and b;
    outputs(7513) <= not a;
    outputs(7514) <= a xor b;
    outputs(7515) <= not b;
    outputs(7516) <= not b or a;
    outputs(7517) <= not (a xor b);
    outputs(7518) <= not a;
    outputs(7519) <= not b;
    outputs(7520) <= b;
    outputs(7521) <= not (a and b);
    outputs(7522) <= a xor b;
    outputs(7523) <= not (a xor b);
    outputs(7524) <= a and b;
    outputs(7525) <= not a;
    outputs(7526) <= a and b;
    outputs(7527) <= not (a or b);
    outputs(7528) <= a and b;
    outputs(7529) <= not b or a;
    outputs(7530) <= not b;
    outputs(7531) <= not a;
    outputs(7532) <= b and not a;
    outputs(7533) <= not (a or b);
    outputs(7534) <= a;
    outputs(7535) <= a;
    outputs(7536) <= a or b;
    outputs(7537) <= not (a xor b);
    outputs(7538) <= a and b;
    outputs(7539) <= a and b;
    outputs(7540) <= b and not a;
    outputs(7541) <= not (a or b);
    outputs(7542) <= not (a xor b);
    outputs(7543) <= b;
    outputs(7544) <= not b;
    outputs(7545) <= not (a xor b);
    outputs(7546) <= a or b;
    outputs(7547) <= not a;
    outputs(7548) <= not b or a;
    outputs(7549) <= not a;
    outputs(7550) <= a;
    outputs(7551) <= b;
    outputs(7552) <= a xor b;
    outputs(7553) <= a and b;
    outputs(7554) <= not a;
    outputs(7555) <= not a;
    outputs(7556) <= a xor b;
    outputs(7557) <= a and not b;
    outputs(7558) <= not b;
    outputs(7559) <= not (a xor b);
    outputs(7560) <= a xor b;
    outputs(7561) <= a;
    outputs(7562) <= a and not b;
    outputs(7563) <= a;
    outputs(7564) <= a;
    outputs(7565) <= not (a or b);
    outputs(7566) <= a and b;
    outputs(7567) <= not (a xor b);
    outputs(7568) <= not a or b;
    outputs(7569) <= not a;
    outputs(7570) <= not (a xor b);
    outputs(7571) <= not a;
    outputs(7572) <= a and b;
    outputs(7573) <= not (a or b);
    outputs(7574) <= a;
    outputs(7575) <= b;
    outputs(7576) <= not a or b;
    outputs(7577) <= not a or b;
    outputs(7578) <= a and b;
    outputs(7579) <= b and not a;
    outputs(7580) <= not a;
    outputs(7581) <= a or b;
    outputs(7582) <= a and not b;
    outputs(7583) <= not a or b;
    outputs(7584) <= a and not b;
    outputs(7585) <= a xor b;
    outputs(7586) <= b and not a;
    outputs(7587) <= not (a or b);
    outputs(7588) <= not a;
    outputs(7589) <= not b;
    outputs(7590) <= not (a xor b);
    outputs(7591) <= not a;
    outputs(7592) <= a and b;
    outputs(7593) <= a;
    outputs(7594) <= a or b;
    outputs(7595) <= not (a xor b);
    outputs(7596) <= a;
    outputs(7597) <= a and not b;
    outputs(7598) <= not b;
    outputs(7599) <= not b;
    outputs(7600) <= b;
    outputs(7601) <= not (a or b);
    outputs(7602) <= a;
    outputs(7603) <= a xor b;
    outputs(7604) <= a xor b;
    outputs(7605) <= not b;
    outputs(7606) <= a and b;
    outputs(7607) <= not a;
    outputs(7608) <= b;
    outputs(7609) <= not (a or b);
    outputs(7610) <= b and not a;
    outputs(7611) <= not (a or b);
    outputs(7612) <= a and b;
    outputs(7613) <= a xor b;
    outputs(7614) <= not (a or b);
    outputs(7615) <= not (a xor b);
    outputs(7616) <= a xor b;
    outputs(7617) <= a;
    outputs(7618) <= a and not b;
    outputs(7619) <= b;
    outputs(7620) <= a xor b;
    outputs(7621) <= not (a xor b);
    outputs(7622) <= a xor b;
    outputs(7623) <= not b;
    outputs(7624) <= a and not b;
    outputs(7625) <= not (a or b);
    outputs(7626) <= a xor b;
    outputs(7627) <= b and not a;
    outputs(7628) <= a and not b;
    outputs(7629) <= not (a xor b);
    outputs(7630) <= not a;
    outputs(7631) <= not (a or b);
    outputs(7632) <= a;
    outputs(7633) <= a;
    outputs(7634) <= not (a xor b);
    outputs(7635) <= a;
    outputs(7636) <= not (a xor b);
    outputs(7637) <= a;
    outputs(7638) <= not a;
    outputs(7639) <= not a;
    outputs(7640) <= not b or a;
    outputs(7641) <= not (a xor b);
    outputs(7642) <= a xor b;
    outputs(7643) <= b and not a;
    outputs(7644) <= not (a xor b);
    outputs(7645) <= not a;
    outputs(7646) <= not b;
    outputs(7647) <= not a;
    outputs(7648) <= not (a xor b);
    outputs(7649) <= a;
    outputs(7650) <= b;
    outputs(7651) <= b and not a;
    outputs(7652) <= a;
    outputs(7653) <= not a;
    outputs(7654) <= not b;
    outputs(7655) <= b;
    outputs(7656) <= a and not b;
    outputs(7657) <= not (a or b);
    outputs(7658) <= not b or a;
    outputs(7659) <= not (a xor b);
    outputs(7660) <= a;
    outputs(7661) <= b;
    outputs(7662) <= a;
    outputs(7663) <= not a;
    outputs(7664) <= not (a xor b);
    outputs(7665) <= a xor b;
    outputs(7666) <= not (a xor b);
    outputs(7667) <= b and not a;
    outputs(7668) <= not b;
    outputs(7669) <= not a;
    outputs(7670) <= a or b;
    outputs(7671) <= not (a xor b);
    outputs(7672) <= b;
    outputs(7673) <= a;
    outputs(7674) <= b;
    outputs(7675) <= not b;
    outputs(7676) <= a or b;
    outputs(7677) <= not (a xor b);
    outputs(7678) <= not b or a;
    outputs(7679) <= a and not b;
    outputs(7680) <= not (a and b);
    outputs(7681) <= a and b;
    outputs(7682) <= b and not a;
    outputs(7683) <= a;
    outputs(7684) <= a and b;
    outputs(7685) <= not b;
    outputs(7686) <= a;
    outputs(7687) <= a;
    outputs(7688) <= not (a xor b);
    outputs(7689) <= not b;
    outputs(7690) <= a;
    outputs(7691) <= not a;
    outputs(7692) <= not (a xor b);
    outputs(7693) <= not (a xor b);
    outputs(7694) <= not a;
    outputs(7695) <= a and b;
    outputs(7696) <= not b or a;
    outputs(7697) <= b;
    outputs(7698) <= not (a or b);
    outputs(7699) <= not (a xor b);
    outputs(7700) <= not a;
    outputs(7701) <= a;
    outputs(7702) <= not b or a;
    outputs(7703) <= not (a and b);
    outputs(7704) <= not b;
    outputs(7705) <= not (a xor b);
    outputs(7706) <= b;
    outputs(7707) <= a xor b;
    outputs(7708) <= a xor b;
    outputs(7709) <= not a;
    outputs(7710) <= a and b;
    outputs(7711) <= a xor b;
    outputs(7712) <= b;
    outputs(7713) <= b;
    outputs(7714) <= not (a xor b);
    outputs(7715) <= a and not b;
    outputs(7716) <= a;
    outputs(7717) <= not (a xor b);
    outputs(7718) <= not (a xor b);
    outputs(7719) <= not (a and b);
    outputs(7720) <= not b;
    outputs(7721) <= a xor b;
    outputs(7722) <= a and b;
    outputs(7723) <= a xor b;
    outputs(7724) <= b;
    outputs(7725) <= a and b;
    outputs(7726) <= not a;
    outputs(7727) <= b and not a;
    outputs(7728) <= a xor b;
    outputs(7729) <= not (a xor b);
    outputs(7730) <= not (a xor b);
    outputs(7731) <= a;
    outputs(7732) <= b;
    outputs(7733) <= not a;
    outputs(7734) <= a;
    outputs(7735) <= a xor b;
    outputs(7736) <= a and not b;
    outputs(7737) <= not (a or b);
    outputs(7738) <= a and b;
    outputs(7739) <= not b;
    outputs(7740) <= b and not a;
    outputs(7741) <= a xor b;
    outputs(7742) <= a xor b;
    outputs(7743) <= a;
    outputs(7744) <= b;
    outputs(7745) <= not a or b;
    outputs(7746) <= a xor b;
    outputs(7747) <= a;
    outputs(7748) <= a xor b;
    outputs(7749) <= not (a xor b);
    outputs(7750) <= a;
    outputs(7751) <= a xor b;
    outputs(7752) <= not (a and b);
    outputs(7753) <= b;
    outputs(7754) <= not a;
    outputs(7755) <= not a;
    outputs(7756) <= a;
    outputs(7757) <= a and b;
    outputs(7758) <= not (a xor b);
    outputs(7759) <= not a or b;
    outputs(7760) <= a xor b;
    outputs(7761) <= a xor b;
    outputs(7762) <= not (a xor b);
    outputs(7763) <= a xor b;
    outputs(7764) <= a xor b;
    outputs(7765) <= not b;
    outputs(7766) <= not a;
    outputs(7767) <= not b;
    outputs(7768) <= not (a xor b);
    outputs(7769) <= a xor b;
    outputs(7770) <= a xor b;
    outputs(7771) <= b;
    outputs(7772) <= a xor b;
    outputs(7773) <= not a;
    outputs(7774) <= a xor b;
    outputs(7775) <= not b;
    outputs(7776) <= a and not b;
    outputs(7777) <= not b;
    outputs(7778) <= a and not b;
    outputs(7779) <= a or b;
    outputs(7780) <= not (a xor b);
    outputs(7781) <= not a or b;
    outputs(7782) <= not (a xor b);
    outputs(7783) <= a;
    outputs(7784) <= not a;
    outputs(7785) <= a or b;
    outputs(7786) <= not (a or b);
    outputs(7787) <= not (a xor b);
    outputs(7788) <= a and not b;
    outputs(7789) <= a and b;
    outputs(7790) <= not a or b;
    outputs(7791) <= not b;
    outputs(7792) <= not b;
    outputs(7793) <= not a;
    outputs(7794) <= not b;
    outputs(7795) <= a and not b;
    outputs(7796) <= a xor b;
    outputs(7797) <= not (a xor b);
    outputs(7798) <= b and not a;
    outputs(7799) <= b;
    outputs(7800) <= a xor b;
    outputs(7801) <= not b;
    outputs(7802) <= not a;
    outputs(7803) <= a xor b;
    outputs(7804) <= not (a xor b);
    outputs(7805) <= a or b;
    outputs(7806) <= a;
    outputs(7807) <= not a or b;
    outputs(7808) <= a or b;
    outputs(7809) <= not (a xor b);
    outputs(7810) <= not (a xor b);
    outputs(7811) <= not (a xor b);
    outputs(7812) <= not b;
    outputs(7813) <= a;
    outputs(7814) <= a;
    outputs(7815) <= not b;
    outputs(7816) <= not a;
    outputs(7817) <= b;
    outputs(7818) <= a;
    outputs(7819) <= a and b;
    outputs(7820) <= b and not a;
    outputs(7821) <= not (a xor b);
    outputs(7822) <= not (a xor b);
    outputs(7823) <= not b;
    outputs(7824) <= a or b;
    outputs(7825) <= not (a xor b);
    outputs(7826) <= a xor b;
    outputs(7827) <= a and not b;
    outputs(7828) <= a;
    outputs(7829) <= b;
    outputs(7830) <= not b;
    outputs(7831) <= b;
    outputs(7832) <= not (a or b);
    outputs(7833) <= not b;
    outputs(7834) <= a xor b;
    outputs(7835) <= a and b;
    outputs(7836) <= a or b;
    outputs(7837) <= a;
    outputs(7838) <= a xor b;
    outputs(7839) <= b;
    outputs(7840) <= a xor b;
    outputs(7841) <= not b;
    outputs(7842) <= not (a xor b);
    outputs(7843) <= not b;
    outputs(7844) <= not a or b;
    outputs(7845) <= a and b;
    outputs(7846) <= not a;
    outputs(7847) <= not (a xor b);
    outputs(7848) <= a;
    outputs(7849) <= a xor b;
    outputs(7850) <= b;
    outputs(7851) <= a;
    outputs(7852) <= not (a xor b);
    outputs(7853) <= a xor b;
    outputs(7854) <= not b;
    outputs(7855) <= not b;
    outputs(7856) <= b and not a;
    outputs(7857) <= a;
    outputs(7858) <= a and not b;
    outputs(7859) <= not (a xor b);
    outputs(7860) <= not b;
    outputs(7861) <= not (a and b);
    outputs(7862) <= a;
    outputs(7863) <= not (a xor b);
    outputs(7864) <= not (a or b);
    outputs(7865) <= not a;
    outputs(7866) <= b;
    outputs(7867) <= b;
    outputs(7868) <= a and b;
    outputs(7869) <= b and not a;
    outputs(7870) <= not (a and b);
    outputs(7871) <= not (a xor b);
    outputs(7872) <= not (a or b);
    outputs(7873) <= b;
    outputs(7874) <= a;
    outputs(7875) <= a xor b;
    outputs(7876) <= not a;
    outputs(7877) <= b;
    outputs(7878) <= a xor b;
    outputs(7879) <= not a;
    outputs(7880) <= a and not b;
    outputs(7881) <= a xor b;
    outputs(7882) <= a xor b;
    outputs(7883) <= not (a and b);
    outputs(7884) <= not (a and b);
    outputs(7885) <= not a;
    outputs(7886) <= b;
    outputs(7887) <= not a;
    outputs(7888) <= a;
    outputs(7889) <= b;
    outputs(7890) <= b and not a;
    outputs(7891) <= a;
    outputs(7892) <= not (a xor b);
    outputs(7893) <= a;
    outputs(7894) <= not b;
    outputs(7895) <= not a;
    outputs(7896) <= a;
    outputs(7897) <= not (a or b);
    outputs(7898) <= not b;
    outputs(7899) <= a;
    outputs(7900) <= a xor b;
    outputs(7901) <= a and b;
    outputs(7902) <= a and not b;
    outputs(7903) <= not a;
    outputs(7904) <= not (a xor b);
    outputs(7905) <= a;
    outputs(7906) <= b and not a;
    outputs(7907) <= a and not b;
    outputs(7908) <= a and b;
    outputs(7909) <= a and not b;
    outputs(7910) <= a and b;
    outputs(7911) <= a xor b;
    outputs(7912) <= b and not a;
    outputs(7913) <= a xor b;
    outputs(7914) <= not b;
    outputs(7915) <= a and not b;
    outputs(7916) <= not a;
    outputs(7917) <= not (a or b);
    outputs(7918) <= b and not a;
    outputs(7919) <= a and b;
    outputs(7920) <= a and not b;
    outputs(7921) <= not b;
    outputs(7922) <= not (a xor b);
    outputs(7923) <= a;
    outputs(7924) <= not (a and b);
    outputs(7925) <= not a;
    outputs(7926) <= not b;
    outputs(7927) <= a;
    outputs(7928) <= not (a xor b);
    outputs(7929) <= not a;
    outputs(7930) <= not (a xor b);
    outputs(7931) <= a and b;
    outputs(7932) <= a;
    outputs(7933) <= not (a xor b);
    outputs(7934) <= b;
    outputs(7935) <= not a;
    outputs(7936) <= a and not b;
    outputs(7937) <= not b;
    outputs(7938) <= a;
    outputs(7939) <= a and not b;
    outputs(7940) <= b;
    outputs(7941) <= b;
    outputs(7942) <= a;
    outputs(7943) <= not b;
    outputs(7944) <= b;
    outputs(7945) <= a xor b;
    outputs(7946) <= b and not a;
    outputs(7947) <= not a;
    outputs(7948) <= a and b;
    outputs(7949) <= not b;
    outputs(7950) <= b;
    outputs(7951) <= not (a or b);
    outputs(7952) <= a xor b;
    outputs(7953) <= a;
    outputs(7954) <= a;
    outputs(7955) <= a;
    outputs(7956) <= a and not b;
    outputs(7957) <= a;
    outputs(7958) <= a;
    outputs(7959) <= not b;
    outputs(7960) <= not b;
    outputs(7961) <= a;
    outputs(7962) <= not a;
    outputs(7963) <= not (a xor b);
    outputs(7964) <= not (a and b);
    outputs(7965) <= b and not a;
    outputs(7966) <= a and b;
    outputs(7967) <= a;
    outputs(7968) <= a and b;
    outputs(7969) <= not a;
    outputs(7970) <= a and not b;
    outputs(7971) <= a and not b;
    outputs(7972) <= a and b;
    outputs(7973) <= b;
    outputs(7974) <= b;
    outputs(7975) <= a and not b;
    outputs(7976) <= not (a xor b);
    outputs(7977) <= not (a xor b);
    outputs(7978) <= b;
    outputs(7979) <= not b;
    outputs(7980) <= b;
    outputs(7981) <= not (a xor b);
    outputs(7982) <= b;
    outputs(7983) <= a and b;
    outputs(7984) <= b and not a;
    outputs(7985) <= b and not a;
    outputs(7986) <= not (a xor b);
    outputs(7987) <= b;
    outputs(7988) <= a xor b;
    outputs(7989) <= a xor b;
    outputs(7990) <= not b;
    outputs(7991) <= not (a or b);
    outputs(7992) <= b;
    outputs(7993) <= not a;
    outputs(7994) <= a or b;
    outputs(7995) <= b and not a;
    outputs(7996) <= a xor b;
    outputs(7997) <= not a;
    outputs(7998) <= a;
    outputs(7999) <= not (a xor b);
    outputs(8000) <= not a;
    outputs(8001) <= not a or b;
    outputs(8002) <= not b;
    outputs(8003) <= a and not b;
    outputs(8004) <= a and not b;
    outputs(8005) <= a xor b;
    outputs(8006) <= not b;
    outputs(8007) <= not a;
    outputs(8008) <= a;
    outputs(8009) <= not (a and b);
    outputs(8010) <= a;
    outputs(8011) <= not (a and b);
    outputs(8012) <= a xor b;
    outputs(8013) <= not (a and b);
    outputs(8014) <= a xor b;
    outputs(8015) <= a and not b;
    outputs(8016) <= not b or a;
    outputs(8017) <= b;
    outputs(8018) <= a;
    outputs(8019) <= b;
    outputs(8020) <= a xor b;
    outputs(8021) <= a;
    outputs(8022) <= a and b;
    outputs(8023) <= a or b;
    outputs(8024) <= b;
    outputs(8025) <= b;
    outputs(8026) <= a xor b;
    outputs(8027) <= b;
    outputs(8028) <= not a;
    outputs(8029) <= b;
    outputs(8030) <= not (a or b);
    outputs(8031) <= not a;
    outputs(8032) <= a and b;
    outputs(8033) <= not a;
    outputs(8034) <= a and b;
    outputs(8035) <= a xor b;
    outputs(8036) <= a;
    outputs(8037) <= not (a xor b);
    outputs(8038) <= a and not b;
    outputs(8039) <= not a;
    outputs(8040) <= not (a xor b);
    outputs(8041) <= not b;
    outputs(8042) <= b;
    outputs(8043) <= a;
    outputs(8044) <= a and not b;
    outputs(8045) <= a;
    outputs(8046) <= not b;
    outputs(8047) <= a;
    outputs(8048) <= a xor b;
    outputs(8049) <= not (a or b);
    outputs(8050) <= not b or a;
    outputs(8051) <= b;
    outputs(8052) <= not a;
    outputs(8053) <= not a;
    outputs(8054) <= not a;
    outputs(8055) <= a xor b;
    outputs(8056) <= a xor b;
    outputs(8057) <= a xor b;
    outputs(8058) <= a and not b;
    outputs(8059) <= a;
    outputs(8060) <= not a or b;
    outputs(8061) <= not a;
    outputs(8062) <= b;
    outputs(8063) <= a xor b;
    outputs(8064) <= a xor b;
    outputs(8065) <= not b;
    outputs(8066) <= b and not a;
    outputs(8067) <= b;
    outputs(8068) <= b;
    outputs(8069) <= b;
    outputs(8070) <= not b;
    outputs(8071) <= not b;
    outputs(8072) <= not b;
    outputs(8073) <= a xor b;
    outputs(8074) <= not (a or b);
    outputs(8075) <= a and not b;
    outputs(8076) <= a and not b;
    outputs(8077) <= not a;
    outputs(8078) <= not (a xor b);
    outputs(8079) <= b and not a;
    outputs(8080) <= not b;
    outputs(8081) <= not (a xor b);
    outputs(8082) <= not b;
    outputs(8083) <= a;
    outputs(8084) <= not (a and b);
    outputs(8085) <= b;
    outputs(8086) <= a xor b;
    outputs(8087) <= not a;
    outputs(8088) <= a;
    outputs(8089) <= not b;
    outputs(8090) <= b;
    outputs(8091) <= b and not a;
    outputs(8092) <= a xor b;
    outputs(8093) <= not b;
    outputs(8094) <= not (a or b);
    outputs(8095) <= b and not a;
    outputs(8096) <= not (a xor b);
    outputs(8097) <= b and not a;
    outputs(8098) <= b and not a;
    outputs(8099) <= a xor b;
    outputs(8100) <= not b;
    outputs(8101) <= a xor b;
    outputs(8102) <= b;
    outputs(8103) <= not (a xor b);
    outputs(8104) <= a and b;
    outputs(8105) <= not b;
    outputs(8106) <= b;
    outputs(8107) <= not (a xor b);
    outputs(8108) <= a xor b;
    outputs(8109) <= not b;
    outputs(8110) <= not (a xor b);
    outputs(8111) <= a xor b;
    outputs(8112) <= not a;
    outputs(8113) <= not b;
    outputs(8114) <= b;
    outputs(8115) <= a or b;
    outputs(8116) <= a and not b;
    outputs(8117) <= a xor b;
    outputs(8118) <= a and b;
    outputs(8119) <= not (a xor b);
    outputs(8120) <= a xor b;
    outputs(8121) <= not b;
    outputs(8122) <= not a;
    outputs(8123) <= not (a and b);
    outputs(8124) <= not b or a;
    outputs(8125) <= a and b;
    outputs(8126) <= a and not b;
    outputs(8127) <= a xor b;
    outputs(8128) <= a and not b;
    outputs(8129) <= a;
    outputs(8130) <= not b;
    outputs(8131) <= not b or a;
    outputs(8132) <= not b;
    outputs(8133) <= a;
    outputs(8134) <= not b;
    outputs(8135) <= not b;
    outputs(8136) <= a and b;
    outputs(8137) <= not a;
    outputs(8138) <= b;
    outputs(8139) <= not a;
    outputs(8140) <= a;
    outputs(8141) <= a xor b;
    outputs(8142) <= a;
    outputs(8143) <= not a;
    outputs(8144) <= a and not b;
    outputs(8145) <= b;
    outputs(8146) <= a;
    outputs(8147) <= a xor b;
    outputs(8148) <= a;
    outputs(8149) <= not (a or b);
    outputs(8150) <= not b;
    outputs(8151) <= not b;
    outputs(8152) <= a xor b;
    outputs(8153) <= not b or a;
    outputs(8154) <= not (a xor b);
    outputs(8155) <= b;
    outputs(8156) <= not b;
    outputs(8157) <= not b or a;
    outputs(8158) <= b;
    outputs(8159) <= not (a xor b);
    outputs(8160) <= a;
    outputs(8161) <= a and b;
    outputs(8162) <= a and b;
    outputs(8163) <= not (a xor b);
    outputs(8164) <= not b;
    outputs(8165) <= a and not b;
    outputs(8166) <= not a;
    outputs(8167) <= not (a xor b);
    outputs(8168) <= not b;
    outputs(8169) <= not a;
    outputs(8170) <= not (a or b);
    outputs(8171) <= not b;
    outputs(8172) <= not (a xor b);
    outputs(8173) <= not a;
    outputs(8174) <= b;
    outputs(8175) <= not (a xor b);
    outputs(8176) <= a and b;
    outputs(8177) <= not (a xor b);
    outputs(8178) <= not b;
    outputs(8179) <= not a;
    outputs(8180) <= a and not b;
    outputs(8181) <= a xor b;
    outputs(8182) <= a;
    outputs(8183) <= a xor b;
    outputs(8184) <= not (a or b);
    outputs(8185) <= a xor b;
    outputs(8186) <= not (a or b);
    outputs(8187) <= not a or b;
    outputs(8188) <= a;
    outputs(8189) <= not a;
    outputs(8190) <= a and b;
    outputs(8191) <= a;
    outputs(8192) <= not (a and b);
    outputs(8193) <= a;
    outputs(8194) <= not b;
    outputs(8195) <= not a;
    outputs(8196) <= a xor b;
    outputs(8197) <= not (a xor b);
    outputs(8198) <= a or b;
    outputs(8199) <= not (a xor b);
    outputs(8200) <= not a;
    outputs(8201) <= a xor b;
    outputs(8202) <= not a;
    outputs(8203) <= not b;
    outputs(8204) <= a;
    outputs(8205) <= not (a xor b);
    outputs(8206) <= not b;
    outputs(8207) <= a;
    outputs(8208) <= not a;
    outputs(8209) <= not b;
    outputs(8210) <= a xor b;
    outputs(8211) <= not (a and b);
    outputs(8212) <= a xor b;
    outputs(8213) <= not (a xor b);
    outputs(8214) <= not (a and b);
    outputs(8215) <= a xor b;
    outputs(8216) <= not (a xor b);
    outputs(8217) <= not (a xor b);
    outputs(8218) <= not (a xor b);
    outputs(8219) <= not (a or b);
    outputs(8220) <= not a;
    outputs(8221) <= a and not b;
    outputs(8222) <= a xor b;
    outputs(8223) <= not a;
    outputs(8224) <= a xor b;
    outputs(8225) <= not b;
    outputs(8226) <= not (a or b);
    outputs(8227) <= not (a and b);
    outputs(8228) <= not (a xor b);
    outputs(8229) <= not a;
    outputs(8230) <= not (a and b);
    outputs(8231) <= b;
    outputs(8232) <= a;
    outputs(8233) <= not a;
    outputs(8234) <= a;
    outputs(8235) <= not (a xor b);
    outputs(8236) <= not (a xor b);
    outputs(8237) <= not b;
    outputs(8238) <= not b;
    outputs(8239) <= b;
    outputs(8240) <= b;
    outputs(8241) <= b;
    outputs(8242) <= b;
    outputs(8243) <= a or b;
    outputs(8244) <= not (a xor b);
    outputs(8245) <= a;
    outputs(8246) <= a xor b;
    outputs(8247) <= not (a xor b);
    outputs(8248) <= a;
    outputs(8249) <= not a or b;
    outputs(8250) <= not (a xor b);
    outputs(8251) <= not (a xor b);
    outputs(8252) <= a xor b;
    outputs(8253) <= b;
    outputs(8254) <= b;
    outputs(8255) <= not b;
    outputs(8256) <= not a;
    outputs(8257) <= b;
    outputs(8258) <= not (a or b);
    outputs(8259) <= not (a or b);
    outputs(8260) <= not a;
    outputs(8261) <= a;
    outputs(8262) <= not (a or b);
    outputs(8263) <= not a;
    outputs(8264) <= a xor b;
    outputs(8265) <= not (a xor b);
    outputs(8266) <= a;
    outputs(8267) <= a and b;
    outputs(8268) <= not b or a;
    outputs(8269) <= not (a xor b);
    outputs(8270) <= not (a and b);
    outputs(8271) <= a xor b;
    outputs(8272) <= a and not b;
    outputs(8273) <= a xor b;
    outputs(8274) <= a xor b;
    outputs(8275) <= not a;
    outputs(8276) <= not a;
    outputs(8277) <= not (a xor b);
    outputs(8278) <= b;
    outputs(8279) <= not b;
    outputs(8280) <= not (a xor b);
    outputs(8281) <= not b;
    outputs(8282) <= not (a xor b);
    outputs(8283) <= not a;
    outputs(8284) <= b;
    outputs(8285) <= a xor b;
    outputs(8286) <= not b or a;
    outputs(8287) <= not (a xor b);
    outputs(8288) <= b;
    outputs(8289) <= a xor b;
    outputs(8290) <= not b or a;
    outputs(8291) <= not a;
    outputs(8292) <= not a;
    outputs(8293) <= not b;
    outputs(8294) <= not a or b;
    outputs(8295) <= a xor b;
    outputs(8296) <= not b;
    outputs(8297) <= a;
    outputs(8298) <= not (a xor b);
    outputs(8299) <= not a or b;
    outputs(8300) <= not (a and b);
    outputs(8301) <= not (a xor b);
    outputs(8302) <= not (a and b);
    outputs(8303) <= not (a xor b);
    outputs(8304) <= a;
    outputs(8305) <= a;
    outputs(8306) <= not b;
    outputs(8307) <= a xor b;
    outputs(8308) <= not a or b;
    outputs(8309) <= not (a xor b);
    outputs(8310) <= not a;
    outputs(8311) <= not (a xor b);
    outputs(8312) <= not (a xor b);
    outputs(8313) <= not (a xor b);
    outputs(8314) <= a;
    outputs(8315) <= a xor b;
    outputs(8316) <= a xor b;
    outputs(8317) <= a xor b;
    outputs(8318) <= a xor b;
    outputs(8319) <= a xor b;
    outputs(8320) <= a xor b;
    outputs(8321) <= not (a xor b);
    outputs(8322) <= not b;
    outputs(8323) <= a xor b;
    outputs(8324) <= a xor b;
    outputs(8325) <= a;
    outputs(8326) <= not b;
    outputs(8327) <= not a;
    outputs(8328) <= a;
    outputs(8329) <= not b or a;
    outputs(8330) <= a;
    outputs(8331) <= not a;
    outputs(8332) <= not (a or b);
    outputs(8333) <= not a;
    outputs(8334) <= a or b;
    outputs(8335) <= not a;
    outputs(8336) <= a xor b;
    outputs(8337) <= not a;
    outputs(8338) <= a xor b;
    outputs(8339) <= b;
    outputs(8340) <= a xor b;
    outputs(8341) <= a;
    outputs(8342) <= not a or b;
    outputs(8343) <= a;
    outputs(8344) <= a xor b;
    outputs(8345) <= not (a xor b);
    outputs(8346) <= not (a or b);
    outputs(8347) <= not a;
    outputs(8348) <= not (a xor b);
    outputs(8349) <= a xor b;
    outputs(8350) <= a;
    outputs(8351) <= not a or b;
    outputs(8352) <= not (a or b);
    outputs(8353) <= a xor b;
    outputs(8354) <= a;
    outputs(8355) <= not b;
    outputs(8356) <= not a;
    outputs(8357) <= not (a xor b);
    outputs(8358) <= not a;
    outputs(8359) <= not b or a;
    outputs(8360) <= a xor b;
    outputs(8361) <= not (a xor b);
    outputs(8362) <= not b;
    outputs(8363) <= a or b;
    outputs(8364) <= not a;
    outputs(8365) <= not (a xor b);
    outputs(8366) <= not b;
    outputs(8367) <= not (a xor b);
    outputs(8368) <= not b or a;
    outputs(8369) <= a;
    outputs(8370) <= not a;
    outputs(8371) <= a;
    outputs(8372) <= a xor b;
    outputs(8373) <= not (a xor b);
    outputs(8374) <= not a;
    outputs(8375) <= not b;
    outputs(8376) <= not b;
    outputs(8377) <= not (a xor b);
    outputs(8378) <= a;
    outputs(8379) <= not a;
    outputs(8380) <= a or b;
    outputs(8381) <= not a or b;
    outputs(8382) <= a xor b;
    outputs(8383) <= not (a xor b);
    outputs(8384) <= a xor b;
    outputs(8385) <= a xor b;
    outputs(8386) <= not (a xor b);
    outputs(8387) <= not a;
    outputs(8388) <= not (a and b);
    outputs(8389) <= not (a xor b);
    outputs(8390) <= a or b;
    outputs(8391) <= not b;
    outputs(8392) <= not (a xor b);
    outputs(8393) <= not b;
    outputs(8394) <= not (a xor b);
    outputs(8395) <= not a or b;
    outputs(8396) <= a xor b;
    outputs(8397) <= b and not a;
    outputs(8398) <= a and not b;
    outputs(8399) <= not a;
    outputs(8400) <= not b or a;
    outputs(8401) <= a and b;
    outputs(8402) <= not a or b;
    outputs(8403) <= a or b;
    outputs(8404) <= a xor b;
    outputs(8405) <= b;
    outputs(8406) <= not (a xor b);
    outputs(8407) <= a or b;
    outputs(8408) <= not (a xor b);
    outputs(8409) <= not b;
    outputs(8410) <= not a;
    outputs(8411) <= b and not a;
    outputs(8412) <= not b or a;
    outputs(8413) <= not (a or b);
    outputs(8414) <= not (a and b);
    outputs(8415) <= not b;
    outputs(8416) <= a xor b;
    outputs(8417) <= not b;
    outputs(8418) <= a;
    outputs(8419) <= not (a xor b);
    outputs(8420) <= not (a xor b);
    outputs(8421) <= not (a xor b);
    outputs(8422) <= not (a xor b);
    outputs(8423) <= a and not b;
    outputs(8424) <= a;
    outputs(8425) <= a xor b;
    outputs(8426) <= not a;
    outputs(8427) <= not (a xor b);
    outputs(8428) <= not (a or b);
    outputs(8429) <= a xor b;
    outputs(8430) <= not b;
    outputs(8431) <= b and not a;
    outputs(8432) <= a xor b;
    outputs(8433) <= not (a xor b);
    outputs(8434) <= not b;
    outputs(8435) <= not (a and b);
    outputs(8436) <= not (a and b);
    outputs(8437) <= b;
    outputs(8438) <= a xor b;
    outputs(8439) <= not b;
    outputs(8440) <= not a or b;
    outputs(8441) <= not b;
    outputs(8442) <= a;
    outputs(8443) <= b;
    outputs(8444) <= not a;
    outputs(8445) <= a and not b;
    outputs(8446) <= b;
    outputs(8447) <= b;
    outputs(8448) <= a xor b;
    outputs(8449) <= not (a xor b);
    outputs(8450) <= not a;
    outputs(8451) <= not a;
    outputs(8452) <= not (a and b);
    outputs(8453) <= a;
    outputs(8454) <= a;
    outputs(8455) <= a xor b;
    outputs(8456) <= not (a xor b);
    outputs(8457) <= not (a xor b);
    outputs(8458) <= not (a or b);
    outputs(8459) <= a xor b;
    outputs(8460) <= a xor b;
    outputs(8461) <= a xor b;
    outputs(8462) <= not (a or b);
    outputs(8463) <= not b;
    outputs(8464) <= not (a or b);
    outputs(8465) <= a xor b;
    outputs(8466) <= a xor b;
    outputs(8467) <= not (a xor b);
    outputs(8468) <= b;
    outputs(8469) <= not a;
    outputs(8470) <= not a;
    outputs(8471) <= a and not b;
    outputs(8472) <= not b;
    outputs(8473) <= not (a xor b);
    outputs(8474) <= a;
    outputs(8475) <= b;
    outputs(8476) <= b;
    outputs(8477) <= not (a xor b);
    outputs(8478) <= not a or b;
    outputs(8479) <= b;
    outputs(8480) <= not (a xor b);
    outputs(8481) <= not (a xor b);
    outputs(8482) <= not a or b;
    outputs(8483) <= b;
    outputs(8484) <= a xor b;
    outputs(8485) <= not a;
    outputs(8486) <= a and b;
    outputs(8487) <= not a or b;
    outputs(8488) <= a xor b;
    outputs(8489) <= not (a xor b);
    outputs(8490) <= a;
    outputs(8491) <= not (a xor b);
    outputs(8492) <= not (a xor b);
    outputs(8493) <= not (a xor b);
    outputs(8494) <= a xor b;
    outputs(8495) <= not b or a;
    outputs(8496) <= not b;
    outputs(8497) <= not b;
    outputs(8498) <= not b;
    outputs(8499) <= not (a xor b);
    outputs(8500) <= a xor b;
    outputs(8501) <= a and b;
    outputs(8502) <= not (a xor b);
    outputs(8503) <= not a;
    outputs(8504) <= b;
    outputs(8505) <= not a;
    outputs(8506) <= a xor b;
    outputs(8507) <= b;
    outputs(8508) <= a xor b;
    outputs(8509) <= not a;
    outputs(8510) <= not b;
    outputs(8511) <= not (a xor b);
    outputs(8512) <= not a;
    outputs(8513) <= b;
    outputs(8514) <= a and b;
    outputs(8515) <= not a;
    outputs(8516) <= not a;
    outputs(8517) <= a or b;
    outputs(8518) <= not (a xor b);
    outputs(8519) <= not a or b;
    outputs(8520) <= b;
    outputs(8521) <= b;
    outputs(8522) <= a and not b;
    outputs(8523) <= b;
    outputs(8524) <= a;
    outputs(8525) <= a or b;
    outputs(8526) <= not b;
    outputs(8527) <= a;
    outputs(8528) <= a;
    outputs(8529) <= not (a xor b);
    outputs(8530) <= a;
    outputs(8531) <= b;
    outputs(8532) <= not a or b;
    outputs(8533) <= not (a xor b);
    outputs(8534) <= not (a xor b);
    outputs(8535) <= not (a xor b);
    outputs(8536) <= not b;
    outputs(8537) <= not b;
    outputs(8538) <= a xor b;
    outputs(8539) <= not b;
    outputs(8540) <= not b;
    outputs(8541) <= not a;
    outputs(8542) <= not (a xor b);
    outputs(8543) <= b;
    outputs(8544) <= not b;
    outputs(8545) <= not (a xor b);
    outputs(8546) <= not a or b;
    outputs(8547) <= b and not a;
    outputs(8548) <= not (a xor b);
    outputs(8549) <= b;
    outputs(8550) <= not a;
    outputs(8551) <= not a or b;
    outputs(8552) <= a;
    outputs(8553) <= not a or b;
    outputs(8554) <= not b or a;
    outputs(8555) <= a xor b;
    outputs(8556) <= a;
    outputs(8557) <= not a;
    outputs(8558) <= a and not b;
    outputs(8559) <= not b;
    outputs(8560) <= not (a xor b);
    outputs(8561) <= b;
    outputs(8562) <= not b;
    outputs(8563) <= not a;
    outputs(8564) <= not a;
    outputs(8565) <= a or b;
    outputs(8566) <= not (a xor b);
    outputs(8567) <= not (a xor b);
    outputs(8568) <= not (a and b);
    outputs(8569) <= a or b;
    outputs(8570) <= not b;
    outputs(8571) <= not (a xor b);
    outputs(8572) <= b;
    outputs(8573) <= not (a xor b);
    outputs(8574) <= a xor b;
    outputs(8575) <= not (a xor b);
    outputs(8576) <= not (a xor b);
    outputs(8577) <= not a;
    outputs(8578) <= a or b;
    outputs(8579) <= not b;
    outputs(8580) <= a and not b;
    outputs(8581) <= a xor b;
    outputs(8582) <= not b or a;
    outputs(8583) <= b;
    outputs(8584) <= not (a xor b);
    outputs(8585) <= b and not a;
    outputs(8586) <= not (a xor b);
    outputs(8587) <= a or b;
    outputs(8588) <= a;
    outputs(8589) <= not (a xor b);
    outputs(8590) <= not (a and b);
    outputs(8591) <= a xor b;
    outputs(8592) <= not b;
    outputs(8593) <= not (a xor b);
    outputs(8594) <= a xor b;
    outputs(8595) <= not (a xor b);
    outputs(8596) <= not (a and b);
    outputs(8597) <= not b;
    outputs(8598) <= not b;
    outputs(8599) <= a;
    outputs(8600) <= not (a xor b);
    outputs(8601) <= a xor b;
    outputs(8602) <= not (a and b);
    outputs(8603) <= not (a xor b);
    outputs(8604) <= not (a xor b);
    outputs(8605) <= not b;
    outputs(8606) <= not (a xor b);
    outputs(8607) <= a and not b;
    outputs(8608) <= not b;
    outputs(8609) <= a;
    outputs(8610) <= a xor b;
    outputs(8611) <= not (a and b);
    outputs(8612) <= a xor b;
    outputs(8613) <= not (a xor b);
    outputs(8614) <= a xor b;
    outputs(8615) <= a xor b;
    outputs(8616) <= not b;
    outputs(8617) <= b;
    outputs(8618) <= not (a or b);
    outputs(8619) <= b;
    outputs(8620) <= not a or b;
    outputs(8621) <= not a;
    outputs(8622) <= not a;
    outputs(8623) <= b;
    outputs(8624) <= b and not a;
    outputs(8625) <= not a or b;
    outputs(8626) <= not b;
    outputs(8627) <= a xor b;
    outputs(8628) <= not (a xor b);
    outputs(8629) <= a xor b;
    outputs(8630) <= not (a or b);
    outputs(8631) <= not (a xor b);
    outputs(8632) <= not b or a;
    outputs(8633) <= a;
    outputs(8634) <= b;
    outputs(8635) <= not a;
    outputs(8636) <= not b or a;
    outputs(8637) <= not a;
    outputs(8638) <= not a;
    outputs(8639) <= not a;
    outputs(8640) <= not a or b;
    outputs(8641) <= not a;
    outputs(8642) <= b;
    outputs(8643) <= not b;
    outputs(8644) <= not a;
    outputs(8645) <= a;
    outputs(8646) <= not b;
    outputs(8647) <= not b;
    outputs(8648) <= b;
    outputs(8649) <= a xor b;
    outputs(8650) <= a xor b;
    outputs(8651) <= not b;
    outputs(8652) <= not (a xor b);
    outputs(8653) <= not b;
    outputs(8654) <= not a;
    outputs(8655) <= b;
    outputs(8656) <= not (a xor b);
    outputs(8657) <= a;
    outputs(8658) <= a xor b;
    outputs(8659) <= not b;
    outputs(8660) <= a;
    outputs(8661) <= not a or b;
    outputs(8662) <= not b;
    outputs(8663) <= not (a xor b);
    outputs(8664) <= a xor b;
    outputs(8665) <= not b;
    outputs(8666) <= a xor b;
    outputs(8667) <= not (a xor b);
    outputs(8668) <= not (a xor b);
    outputs(8669) <= not a;
    outputs(8670) <= not (a xor b);
    outputs(8671) <= a;
    outputs(8672) <= not a;
    outputs(8673) <= a;
    outputs(8674) <= a xor b;
    outputs(8675) <= a;
    outputs(8676) <= b;
    outputs(8677) <= not b;
    outputs(8678) <= not (a and b);
    outputs(8679) <= not a or b;
    outputs(8680) <= not a;
    outputs(8681) <= not a;
    outputs(8682) <= a xor b;
    outputs(8683) <= not (a xor b);
    outputs(8684) <= not (a xor b);
    outputs(8685) <= not a;
    outputs(8686) <= a and not b;
    outputs(8687) <= not (a or b);
    outputs(8688) <= a xor b;
    outputs(8689) <= a xor b;
    outputs(8690) <= not a;
    outputs(8691) <= not (a or b);
    outputs(8692) <= not b;
    outputs(8693) <= a;
    outputs(8694) <= not a or b;
    outputs(8695) <= a and not b;
    outputs(8696) <= not (a xor b);
    outputs(8697) <= not a;
    outputs(8698) <= b;
    outputs(8699) <= a xor b;
    outputs(8700) <= not a;
    outputs(8701) <= not (a or b);
    outputs(8702) <= not (a xor b);
    outputs(8703) <= a xor b;
    outputs(8704) <= not b;
    outputs(8705) <= not b;
    outputs(8706) <= b;
    outputs(8707) <= not (a xor b);
    outputs(8708) <= b and not a;
    outputs(8709) <= b and not a;
    outputs(8710) <= a and b;
    outputs(8711) <= not b;
    outputs(8712) <= not (a or b);
    outputs(8713) <= not (a xor b);
    outputs(8714) <= a xor b;
    outputs(8715) <= not (a and b);
    outputs(8716) <= a xor b;
    outputs(8717) <= not b;
    outputs(8718) <= a xor b;
    outputs(8719) <= not (a xor b);
    outputs(8720) <= a xor b;
    outputs(8721) <= not a;
    outputs(8722) <= a xor b;
    outputs(8723) <= not a;
    outputs(8724) <= not (a xor b);
    outputs(8725) <= a and not b;
    outputs(8726) <= a xor b;
    outputs(8727) <= not b;
    outputs(8728) <= not (a or b);
    outputs(8729) <= a;
    outputs(8730) <= a or b;
    outputs(8731) <= a and b;
    outputs(8732) <= not b or a;
    outputs(8733) <= b;
    outputs(8734) <= a;
    outputs(8735) <= b;
    outputs(8736) <= a;
    outputs(8737) <= not a;
    outputs(8738) <= a or b;
    outputs(8739) <= b;
    outputs(8740) <= a;
    outputs(8741) <= a or b;
    outputs(8742) <= b;
    outputs(8743) <= a xor b;
    outputs(8744) <= not (a xor b);
    outputs(8745) <= not (a xor b);
    outputs(8746) <= b;
    outputs(8747) <= not a or b;
    outputs(8748) <= b;
    outputs(8749) <= not b;
    outputs(8750) <= a;
    outputs(8751) <= b;
    outputs(8752) <= a xor b;
    outputs(8753) <= not a;
    outputs(8754) <= not a;
    outputs(8755) <= b;
    outputs(8756) <= a xor b;
    outputs(8757) <= not b or a;
    outputs(8758) <= a or b;
    outputs(8759) <= not b;
    outputs(8760) <= a xor b;
    outputs(8761) <= not (a xor b);
    outputs(8762) <= b;
    outputs(8763) <= not a;
    outputs(8764) <= not b or a;
    outputs(8765) <= a xor b;
    outputs(8766) <= not (a or b);
    outputs(8767) <= a;
    outputs(8768) <= not a;
    outputs(8769) <= not b or a;
    outputs(8770) <= a;
    outputs(8771) <= not (a and b);
    outputs(8772) <= not (a xor b);
    outputs(8773) <= not (a xor b);
    outputs(8774) <= b;
    outputs(8775) <= a and b;
    outputs(8776) <= not a;
    outputs(8777) <= a xor b;
    outputs(8778) <= b;
    outputs(8779) <= a or b;
    outputs(8780) <= a;
    outputs(8781) <= not a;
    outputs(8782) <= a xor b;
    outputs(8783) <= a;
    outputs(8784) <= not (a xor b);
    outputs(8785) <= a xor b;
    outputs(8786) <= not b or a;
    outputs(8787) <= not (a or b);
    outputs(8788) <= a xor b;
    outputs(8789) <= not a;
    outputs(8790) <= a xor b;
    outputs(8791) <= not b;
    outputs(8792) <= a;
    outputs(8793) <= b;
    outputs(8794) <= not a;
    outputs(8795) <= not (a xor b);
    outputs(8796) <= not a;
    outputs(8797) <= a xor b;
    outputs(8798) <= a or b;
    outputs(8799) <= a and not b;
    outputs(8800) <= not a or b;
    outputs(8801) <= not b;
    outputs(8802) <= a xor b;
    outputs(8803) <= not (a xor b);
    outputs(8804) <= a xor b;
    outputs(8805) <= a or b;
    outputs(8806) <= a xor b;
    outputs(8807) <= not a;
    outputs(8808) <= a xor b;
    outputs(8809) <= not (a and b);
    outputs(8810) <= not (a and b);
    outputs(8811) <= a;
    outputs(8812) <= not a;
    outputs(8813) <= a;
    outputs(8814) <= a and not b;
    outputs(8815) <= a xor b;
    outputs(8816) <= not b;
    outputs(8817) <= not b;
    outputs(8818) <= not a or b;
    outputs(8819) <= b;
    outputs(8820) <= not b;
    outputs(8821) <= not a or b;
    outputs(8822) <= not a;
    outputs(8823) <= a and not b;
    outputs(8824) <= not (a xor b);
    outputs(8825) <= not (a xor b);
    outputs(8826) <= a;
    outputs(8827) <= not (a xor b);
    outputs(8828) <= not b or a;
    outputs(8829) <= not (a xor b);
    outputs(8830) <= a xor b;
    outputs(8831) <= a xor b;
    outputs(8832) <= not b;
    outputs(8833) <= a and b;
    outputs(8834) <= b and not a;
    outputs(8835) <= not b;
    outputs(8836) <= b;
    outputs(8837) <= not (a xor b);
    outputs(8838) <= not b or a;
    outputs(8839) <= not (a or b);
    outputs(8840) <= a xor b;
    outputs(8841) <= a xor b;
    outputs(8842) <= a xor b;
    outputs(8843) <= not (a xor b);
    outputs(8844) <= not (a and b);
    outputs(8845) <= a xor b;
    outputs(8846) <= not (a xor b);
    outputs(8847) <= a xor b;
    outputs(8848) <= a or b;
    outputs(8849) <= not (a xor b);
    outputs(8850) <= a or b;
    outputs(8851) <= a xor b;
    outputs(8852) <= not a;
    outputs(8853) <= a or b;
    outputs(8854) <= a xor b;
    outputs(8855) <= a xor b;
    outputs(8856) <= a or b;
    outputs(8857) <= not (a xor b);
    outputs(8858) <= a;
    outputs(8859) <= a;
    outputs(8860) <= a xor b;
    outputs(8861) <= not b;
    outputs(8862) <= not b;
    outputs(8863) <= not a;
    outputs(8864) <= not a;
    outputs(8865) <= b;
    outputs(8866) <= b;
    outputs(8867) <= not (a xor b);
    outputs(8868) <= a xor b;
    outputs(8869) <= not b;
    outputs(8870) <= not a or b;
    outputs(8871) <= b and not a;
    outputs(8872) <= a xor b;
    outputs(8873) <= not (a xor b);
    outputs(8874) <= not (a xor b);
    outputs(8875) <= not a or b;
    outputs(8876) <= not (a xor b);
    outputs(8877) <= not (a xor b);
    outputs(8878) <= a;
    outputs(8879) <= not (a xor b);
    outputs(8880) <= not (a xor b);
    outputs(8881) <= a;
    outputs(8882) <= not b or a;
    outputs(8883) <= not b;
    outputs(8884) <= b;
    outputs(8885) <= not (a xor b);
    outputs(8886) <= a;
    outputs(8887) <= a or b;
    outputs(8888) <= a or b;
    outputs(8889) <= a;
    outputs(8890) <= a and not b;
    outputs(8891) <= a xor b;
    outputs(8892) <= not a;
    outputs(8893) <= not (a xor b);
    outputs(8894) <= not (a and b);
    outputs(8895) <= not a;
    outputs(8896) <= not b;
    outputs(8897) <= not a;
    outputs(8898) <= not (a and b);
    outputs(8899) <= not (a xor b);
    outputs(8900) <= not b;
    outputs(8901) <= b and not a;
    outputs(8902) <= a xor b;
    outputs(8903) <= not (a or b);
    outputs(8904) <= a xor b;
    outputs(8905) <= a;
    outputs(8906) <= a xor b;
    outputs(8907) <= a;
    outputs(8908) <= a xor b;
    outputs(8909) <= not b;
    outputs(8910) <= b;
    outputs(8911) <= not b;
    outputs(8912) <= a and b;
    outputs(8913) <= a xor b;
    outputs(8914) <= a;
    outputs(8915) <= not b;
    outputs(8916) <= a and not b;
    outputs(8917) <= b;
    outputs(8918) <= not b;
    outputs(8919) <= not (a xor b);
    outputs(8920) <= b;
    outputs(8921) <= not (a xor b);
    outputs(8922) <= not b;
    outputs(8923) <= not b;
    outputs(8924) <= a xor b;
    outputs(8925) <= not b or a;
    outputs(8926) <= a xor b;
    outputs(8927) <= a;
    outputs(8928) <= a xor b;
    outputs(8929) <= not (a xor b);
    outputs(8930) <= not b;
    outputs(8931) <= b;
    outputs(8932) <= not a;
    outputs(8933) <= not (a or b);
    outputs(8934) <= a;
    outputs(8935) <= b;
    outputs(8936) <= a;
    outputs(8937) <= a xor b;
    outputs(8938) <= not b;
    outputs(8939) <= a xor b;
    outputs(8940) <= not b;
    outputs(8941) <= not (a xor b);
    outputs(8942) <= not (a xor b);
    outputs(8943) <= not (a xor b);
    outputs(8944) <= b;
    outputs(8945) <= not (a xor b);
    outputs(8946) <= not (a xor b);
    outputs(8947) <= a xor b;
    outputs(8948) <= a;
    outputs(8949) <= not (a xor b);
    outputs(8950) <= not a;
    outputs(8951) <= a and not b;
    outputs(8952) <= not (a or b);
    outputs(8953) <= not (a xor b);
    outputs(8954) <= a xor b;
    outputs(8955) <= b and not a;
    outputs(8956) <= not a;
    outputs(8957) <= a and b;
    outputs(8958) <= not a;
    outputs(8959) <= a;
    outputs(8960) <= a xor b;
    outputs(8961) <= not a or b;
    outputs(8962) <= not b;
    outputs(8963) <= a and b;
    outputs(8964) <= a and not b;
    outputs(8965) <= b;
    outputs(8966) <= not a or b;
    outputs(8967) <= not (a xor b);
    outputs(8968) <= a xor b;
    outputs(8969) <= a;
    outputs(8970) <= b;
    outputs(8971) <= not a;
    outputs(8972) <= not a;
    outputs(8973) <= not b;
    outputs(8974) <= not (a xor b);
    outputs(8975) <= a and not b;
    outputs(8976) <= a;
    outputs(8977) <= not (a and b);
    outputs(8978) <= not a;
    outputs(8979) <= a and not b;
    outputs(8980) <= not (a xor b);
    outputs(8981) <= not b;
    outputs(8982) <= a xor b;
    outputs(8983) <= not (a xor b);
    outputs(8984) <= not b;
    outputs(8985) <= b;
    outputs(8986) <= not (a xor b);
    outputs(8987) <= not a;
    outputs(8988) <= b;
    outputs(8989) <= a xor b;
    outputs(8990) <= not a or b;
    outputs(8991) <= not b;
    outputs(8992) <= b and not a;
    outputs(8993) <= a;
    outputs(8994) <= a or b;
    outputs(8995) <= not b;
    outputs(8996) <= not a;
    outputs(8997) <= not (a xor b);
    outputs(8998) <= not a or b;
    outputs(8999) <= not b;
    outputs(9000) <= not b;
    outputs(9001) <= a;
    outputs(9002) <= a or b;
    outputs(9003) <= not (a xor b);
    outputs(9004) <= b;
    outputs(9005) <= a or b;
    outputs(9006) <= a xor b;
    outputs(9007) <= a;
    outputs(9008) <= a xor b;
    outputs(9009) <= a or b;
    outputs(9010) <= not b;
    outputs(9011) <= not b;
    outputs(9012) <= a;
    outputs(9013) <= not b;
    outputs(9014) <= b;
    outputs(9015) <= not (a xor b);
    outputs(9016) <= not (a xor b);
    outputs(9017) <= a;
    outputs(9018) <= not (a and b);
    outputs(9019) <= a;
    outputs(9020) <= a xor b;
    outputs(9021) <= a xor b;
    outputs(9022) <= a xor b;
    outputs(9023) <= not b or a;
    outputs(9024) <= not (a xor b);
    outputs(9025) <= b;
    outputs(9026) <= b;
    outputs(9027) <= a xor b;
    outputs(9028) <= not (a xor b);
    outputs(9029) <= not a;
    outputs(9030) <= not (a xor b);
    outputs(9031) <= a xor b;
    outputs(9032) <= not (a and b);
    outputs(9033) <= a xor b;
    outputs(9034) <= a and b;
    outputs(9035) <= not (a xor b);
    outputs(9036) <= a and not b;
    outputs(9037) <= not (a xor b);
    outputs(9038) <= not (a xor b);
    outputs(9039) <= b;
    outputs(9040) <= not b;
    outputs(9041) <= not b;
    outputs(9042) <= not (a xor b);
    outputs(9043) <= not b;
    outputs(9044) <= a;
    outputs(9045) <= not (a xor b);
    outputs(9046) <= a and not b;
    outputs(9047) <= a xor b;
    outputs(9048) <= not b;
    outputs(9049) <= not (a xor b);
    outputs(9050) <= a xor b;
    outputs(9051) <= a xor b;
    outputs(9052) <= not (a xor b);
    outputs(9053) <= not b;
    outputs(9054) <= a xor b;
    outputs(9055) <= not b or a;
    outputs(9056) <= not (a xor b);
    outputs(9057) <= a;
    outputs(9058) <= not b;
    outputs(9059) <= b and not a;
    outputs(9060) <= a;
    outputs(9061) <= a and not b;
    outputs(9062) <= a or b;
    outputs(9063) <= b and not a;
    outputs(9064) <= not (a xor b);
    outputs(9065) <= b;
    outputs(9066) <= b;
    outputs(9067) <= not (a xor b);
    outputs(9068) <= not (a xor b);
    outputs(9069) <= a xor b;
    outputs(9070) <= not (a xor b);
    outputs(9071) <= not (a xor b);
    outputs(9072) <= a xor b;
    outputs(9073) <= not a;
    outputs(9074) <= b and not a;
    outputs(9075) <= not b;
    outputs(9076) <= b;
    outputs(9077) <= not b;
    outputs(9078) <= b;
    outputs(9079) <= not (a xor b);
    outputs(9080) <= a;
    outputs(9081) <= b;
    outputs(9082) <= a xor b;
    outputs(9083) <= a xor b;
    outputs(9084) <= not (a and b);
    outputs(9085) <= a xor b;
    outputs(9086) <= not (a xor b);
    outputs(9087) <= a;
    outputs(9088) <= not (a xor b);
    outputs(9089) <= a or b;
    outputs(9090) <= a xor b;
    outputs(9091) <= not a;
    outputs(9092) <= b;
    outputs(9093) <= a xor b;
    outputs(9094) <= not b;
    outputs(9095) <= not (a xor b);
    outputs(9096) <= not b or a;
    outputs(9097) <= b;
    outputs(9098) <= a xor b;
    outputs(9099) <= not (a xor b);
    outputs(9100) <= b;
    outputs(9101) <= a and not b;
    outputs(9102) <= b;
    outputs(9103) <= a xor b;
    outputs(9104) <= not (a xor b);
    outputs(9105) <= a xor b;
    outputs(9106) <= b;
    outputs(9107) <= a or b;
    outputs(9108) <= not b;
    outputs(9109) <= not a or b;
    outputs(9110) <= b;
    outputs(9111) <= a;
    outputs(9112) <= b;
    outputs(9113) <= not (a and b);
    outputs(9114) <= a;
    outputs(9115) <= not a;
    outputs(9116) <= a xor b;
    outputs(9117) <= not (a xor b);
    outputs(9118) <= not b;
    outputs(9119) <= not a or b;
    outputs(9120) <= not b;
    outputs(9121) <= a or b;
    outputs(9122) <= b;
    outputs(9123) <= a;
    outputs(9124) <= a or b;
    outputs(9125) <= not b;
    outputs(9126) <= a xor b;
    outputs(9127) <= b;
    outputs(9128) <= b and not a;
    outputs(9129) <= a xor b;
    outputs(9130) <= not b;
    outputs(9131) <= a;
    outputs(9132) <= a or b;
    outputs(9133) <= b;
    outputs(9134) <= a xor b;
    outputs(9135) <= a xor b;
    outputs(9136) <= a or b;
    outputs(9137) <= not a;
    outputs(9138) <= not b;
    outputs(9139) <= a xor b;
    outputs(9140) <= b;
    outputs(9141) <= not b;
    outputs(9142) <= a xor b;
    outputs(9143) <= a xor b;
    outputs(9144) <= a xor b;
    outputs(9145) <= a xor b;
    outputs(9146) <= not a or b;
    outputs(9147) <= b and not a;
    outputs(9148) <= not b;
    outputs(9149) <= a and b;
    outputs(9150) <= not (a xor b);
    outputs(9151) <= a and not b;
    outputs(9152) <= not (a or b);
    outputs(9153) <= not (a and b);
    outputs(9154) <= a;
    outputs(9155) <= not a or b;
    outputs(9156) <= not b;
    outputs(9157) <= b;
    outputs(9158) <= not b;
    outputs(9159) <= not b;
    outputs(9160) <= not a;
    outputs(9161) <= not (a xor b);
    outputs(9162) <= not (a xor b);
    outputs(9163) <= not b;
    outputs(9164) <= a xor b;
    outputs(9165) <= a xor b;
    outputs(9166) <= not a;
    outputs(9167) <= a;
    outputs(9168) <= not (a xor b);
    outputs(9169) <= not (a xor b);
    outputs(9170) <= not (a xor b);
    outputs(9171) <= not (a xor b);
    outputs(9172) <= a;
    outputs(9173) <= b;
    outputs(9174) <= not (a xor b);
    outputs(9175) <= a xor b;
    outputs(9176) <= not (a and b);
    outputs(9177) <= not (a xor b);
    outputs(9178) <= a xor b;
    outputs(9179) <= not a;
    outputs(9180) <= not a;
    outputs(9181) <= a;
    outputs(9182) <= not a;
    outputs(9183) <= not b;
    outputs(9184) <= not a;
    outputs(9185) <= a xor b;
    outputs(9186) <= not (a xor b);
    outputs(9187) <= not (a xor b);
    outputs(9188) <= a or b;
    outputs(9189) <= not (a or b);
    outputs(9190) <= not (a or b);
    outputs(9191) <= a;
    outputs(9192) <= a or b;
    outputs(9193) <= not a or b;
    outputs(9194) <= a xor b;
    outputs(9195) <= a and not b;
    outputs(9196) <= b;
    outputs(9197) <= not a;
    outputs(9198) <= a;
    outputs(9199) <= not a or b;
    outputs(9200) <= not a;
    outputs(9201) <= not (a xor b);
    outputs(9202) <= a;
    outputs(9203) <= a xor b;
    outputs(9204) <= not (a xor b);
    outputs(9205) <= not (a xor b);
    outputs(9206) <= not b;
    outputs(9207) <= b;
    outputs(9208) <= a and b;
    outputs(9209) <= not (a or b);
    outputs(9210) <= not a or b;
    outputs(9211) <= b;
    outputs(9212) <= a xor b;
    outputs(9213) <= not (a and b);
    outputs(9214) <= not a;
    outputs(9215) <= a xor b;
    outputs(9216) <= not (a or b);
    outputs(9217) <= a or b;
    outputs(9218) <= not (a and b);
    outputs(9219) <= not a;
    outputs(9220) <= a;
    outputs(9221) <= not a;
    outputs(9222) <= b and not a;
    outputs(9223) <= a;
    outputs(9224) <= a and not b;
    outputs(9225) <= b;
    outputs(9226) <= not (a or b);
    outputs(9227) <= not b or a;
    outputs(9228) <= a xor b;
    outputs(9229) <= a xor b;
    outputs(9230) <= a;
    outputs(9231) <= not (a xor b);
    outputs(9232) <= a xor b;
    outputs(9233) <= a;
    outputs(9234) <= a xor b;
    outputs(9235) <= b;
    outputs(9236) <= b;
    outputs(9237) <= not (a xor b);
    outputs(9238) <= not (a or b);
    outputs(9239) <= a or b;
    outputs(9240) <= b;
    outputs(9241) <= not (a or b);
    outputs(9242) <= not (a or b);
    outputs(9243) <= a xor b;
    outputs(9244) <= not (a xor b);
    outputs(9245) <= not (a and b);
    outputs(9246) <= a;
    outputs(9247) <= a xor b;
    outputs(9248) <= not a;
    outputs(9249) <= b;
    outputs(9250) <= b;
    outputs(9251) <= b;
    outputs(9252) <= not (a or b);
    outputs(9253) <= b;
    outputs(9254) <= a xor b;
    outputs(9255) <= b;
    outputs(9256) <= a and not b;
    outputs(9257) <= a;
    outputs(9258) <= not a;
    outputs(9259) <= a and b;
    outputs(9260) <= a xor b;
    outputs(9261) <= a or b;
    outputs(9262) <= not (a xor b);
    outputs(9263) <= not (a xor b);
    outputs(9264) <= a and b;
    outputs(9265) <= not b;
    outputs(9266) <= a xor b;
    outputs(9267) <= a and b;
    outputs(9268) <= not (a xor b);
    outputs(9269) <= not (a or b);
    outputs(9270) <= not (a and b);
    outputs(9271) <= not (a xor b);
    outputs(9272) <= a;
    outputs(9273) <= not (a xor b);
    outputs(9274) <= not b;
    outputs(9275) <= a;
    outputs(9276) <= b;
    outputs(9277) <= not b;
    outputs(9278) <= not a;
    outputs(9279) <= a xor b;
    outputs(9280) <= a xor b;
    outputs(9281) <= a;
    outputs(9282) <= not (a xor b);
    outputs(9283) <= a;
    outputs(9284) <= not (a xor b);
    outputs(9285) <= a;
    outputs(9286) <= a and b;
    outputs(9287) <= a and b;
    outputs(9288) <= a xor b;
    outputs(9289) <= not (a xor b);
    outputs(9290) <= not a;
    outputs(9291) <= a and b;
    outputs(9292) <= a and b;
    outputs(9293) <= a xor b;
    outputs(9294) <= not (a xor b);
    outputs(9295) <= a xor b;
    outputs(9296) <= a;
    outputs(9297) <= not a;
    outputs(9298) <= not (a xor b);
    outputs(9299) <= not b or a;
    outputs(9300) <= not (a and b);
    outputs(9301) <= not b;
    outputs(9302) <= b;
    outputs(9303) <= not (a xor b);
    outputs(9304) <= a;
    outputs(9305) <= not (a xor b);
    outputs(9306) <= not b;
    outputs(9307) <= not a;
    outputs(9308) <= not (a and b);
    outputs(9309) <= b and not a;
    outputs(9310) <= a;
    outputs(9311) <= not b;
    outputs(9312) <= a xor b;
    outputs(9313) <= a xor b;
    outputs(9314) <= a;
    outputs(9315) <= not (a or b);
    outputs(9316) <= b;
    outputs(9317) <= a and not b;
    outputs(9318) <= b;
    outputs(9319) <= not b or a;
    outputs(9320) <= not b;
    outputs(9321) <= b;
    outputs(9322) <= not (a xor b);
    outputs(9323) <= not (a or b);
    outputs(9324) <= not b;
    outputs(9325) <= not b;
    outputs(9326) <= not (a xor b);
    outputs(9327) <= a and not b;
    outputs(9328) <= 1'b1;
    outputs(9329) <= not (a xor b);
    outputs(9330) <= not b;
    outputs(9331) <= b and not a;
    outputs(9332) <= not a;
    outputs(9333) <= not (a or b);
    outputs(9334) <= a xor b;
    outputs(9335) <= a xor b;
    outputs(9336) <= not (a xor b);
    outputs(9337) <= a xor b;
    outputs(9338) <= a and b;
    outputs(9339) <= b and not a;
    outputs(9340) <= b and not a;
    outputs(9341) <= a and b;
    outputs(9342) <= not a;
    outputs(9343) <= not b;
    outputs(9344) <= b;
    outputs(9345) <= a xor b;
    outputs(9346) <= a xor b;
    outputs(9347) <= a xor b;
    outputs(9348) <= not b;
    outputs(9349) <= a xor b;
    outputs(9350) <= a xor b;
    outputs(9351) <= not a;
    outputs(9352) <= not (a or b);
    outputs(9353) <= b;
    outputs(9354) <= a and not b;
    outputs(9355) <= a and not b;
    outputs(9356) <= a or b;
    outputs(9357) <= a;
    outputs(9358) <= b and not a;
    outputs(9359) <= a xor b;
    outputs(9360) <= not a;
    outputs(9361) <= b and not a;
    outputs(9362) <= a and b;
    outputs(9363) <= b;
    outputs(9364) <= a xor b;
    outputs(9365) <= a xor b;
    outputs(9366) <= a and b;
    outputs(9367) <= a or b;
    outputs(9368) <= not a;
    outputs(9369) <= a;
    outputs(9370) <= a xor b;
    outputs(9371) <= a xor b;
    outputs(9372) <= a and not b;
    outputs(9373) <= not (a xor b);
    outputs(9374) <= a;
    outputs(9375) <= a and b;
    outputs(9376) <= not a;
    outputs(9377) <= not b;
    outputs(9378) <= a and not b;
    outputs(9379) <= not (a xor b);
    outputs(9380) <= not (a xor b);
    outputs(9381) <= not a;
    outputs(9382) <= not (a xor b);
    outputs(9383) <= not b;
    outputs(9384) <= a and b;
    outputs(9385) <= not b;
    outputs(9386) <= not (a xor b);
    outputs(9387) <= a and b;
    outputs(9388) <= b and not a;
    outputs(9389) <= a or b;
    outputs(9390) <= not (a xor b);
    outputs(9391) <= not a;
    outputs(9392) <= a and b;
    outputs(9393) <= not (a xor b);
    outputs(9394) <= not a;
    outputs(9395) <= b and not a;
    outputs(9396) <= not b or a;
    outputs(9397) <= a and b;
    outputs(9398) <= not b;
    outputs(9399) <= a;
    outputs(9400) <= b and not a;
    outputs(9401) <= not a;
    outputs(9402) <= a or b;
    outputs(9403) <= not (a xor b);
    outputs(9404) <= a xor b;
    outputs(9405) <= b and not a;
    outputs(9406) <= not (a or b);
    outputs(9407) <= not b or a;
    outputs(9408) <= not (a and b);
    outputs(9409) <= not (a xor b);
    outputs(9410) <= a xor b;
    outputs(9411) <= a;
    outputs(9412) <= b;
    outputs(9413) <= not a;
    outputs(9414) <= a and not b;
    outputs(9415) <= b;
    outputs(9416) <= not (a or b);
    outputs(9417) <= b;
    outputs(9418) <= not (a xor b);
    outputs(9419) <= b;
    outputs(9420) <= a xor b;
    outputs(9421) <= b;
    outputs(9422) <= not b;
    outputs(9423) <= a xor b;
    outputs(9424) <= not (a xor b);
    outputs(9425) <= a xor b;
    outputs(9426) <= not (a xor b);
    outputs(9427) <= a and not b;
    outputs(9428) <= not a;
    outputs(9429) <= not (a xor b);
    outputs(9430) <= not a;
    outputs(9431) <= b;
    outputs(9432) <= a and b;
    outputs(9433) <= a xor b;
    outputs(9434) <= not (a xor b);
    outputs(9435) <= not (a and b);
    outputs(9436) <= a;
    outputs(9437) <= not (a xor b);
    outputs(9438) <= a;
    outputs(9439) <= a;
    outputs(9440) <= a xor b;
    outputs(9441) <= a xor b;
    outputs(9442) <= a xor b;
    outputs(9443) <= a xor b;
    outputs(9444) <= not a;
    outputs(9445) <= not b;
    outputs(9446) <= not (a xor b);
    outputs(9447) <= not b or a;
    outputs(9448) <= not a;
    outputs(9449) <= a;
    outputs(9450) <= not (a and b);
    outputs(9451) <= b;
    outputs(9452) <= not (a and b);
    outputs(9453) <= a;
    outputs(9454) <= not a or b;
    outputs(9455) <= not b;
    outputs(9456) <= b;
    outputs(9457) <= a;
    outputs(9458) <= not b or a;
    outputs(9459) <= b and not a;
    outputs(9460) <= a xor b;
    outputs(9461) <= b and not a;
    outputs(9462) <= not (a or b);
    outputs(9463) <= not a;
    outputs(9464) <= not a;
    outputs(9465) <= a and not b;
    outputs(9466) <= b;
    outputs(9467) <= a and not b;
    outputs(9468) <= not b;
    outputs(9469) <= not (a xor b);
    outputs(9470) <= not b;
    outputs(9471) <= not (a xor b);
    outputs(9472) <= not (a xor b);
    outputs(9473) <= a;
    outputs(9474) <= b;
    outputs(9475) <= a xor b;
    outputs(9476) <= a;
    outputs(9477) <= a xor b;
    outputs(9478) <= not a or b;
    outputs(9479) <= not (a xor b);
    outputs(9480) <= not b;
    outputs(9481) <= not (a xor b);
    outputs(9482) <= b and not a;
    outputs(9483) <= b and not a;
    outputs(9484) <= not (a xor b);
    outputs(9485) <= a and b;
    outputs(9486) <= not (a xor b);
    outputs(9487) <= not b;
    outputs(9488) <= a;
    outputs(9489) <= not a;
    outputs(9490) <= not b;
    outputs(9491) <= a xor b;
    outputs(9492) <= a and not b;
    outputs(9493) <= not a;
    outputs(9494) <= a;
    outputs(9495) <= not a or b;
    outputs(9496) <= b and not a;
    outputs(9497) <= not b;
    outputs(9498) <= b and not a;
    outputs(9499) <= not a;
    outputs(9500) <= a;
    outputs(9501) <= a and not b;
    outputs(9502) <= not (a and b);
    outputs(9503) <= not a or b;
    outputs(9504) <= not (a or b);
    outputs(9505) <= not a;
    outputs(9506) <= not b or a;
    outputs(9507) <= a;
    outputs(9508) <= b;
    outputs(9509) <= not (a xor b);
    outputs(9510) <= not b;
    outputs(9511) <= not b;
    outputs(9512) <= a and not b;
    outputs(9513) <= not b;
    outputs(9514) <= a and not b;
    outputs(9515) <= a;
    outputs(9516) <= not (a xor b);
    outputs(9517) <= not b or a;
    outputs(9518) <= a and not b;
    outputs(9519) <= a xor b;
    outputs(9520) <= not b or a;
    outputs(9521) <= not (a xor b);
    outputs(9522) <= not a;
    outputs(9523) <= a xor b;
    outputs(9524) <= b;
    outputs(9525) <= not b;
    outputs(9526) <= a;
    outputs(9527) <= a xor b;
    outputs(9528) <= not b;
    outputs(9529) <= not a or b;
    outputs(9530) <= a xor b;
    outputs(9531) <= not a;
    outputs(9532) <= b;
    outputs(9533) <= a and not b;
    outputs(9534) <= not a or b;
    outputs(9535) <= not (a xor b);
    outputs(9536) <= not (a xor b);
    outputs(9537) <= not a;
    outputs(9538) <= not b;
    outputs(9539) <= not b or a;
    outputs(9540) <= b;
    outputs(9541) <= not (a xor b);
    outputs(9542) <= a xor b;
    outputs(9543) <= b;
    outputs(9544) <= a and b;
    outputs(9545) <= b;
    outputs(9546) <= not a;
    outputs(9547) <= not a;
    outputs(9548) <= a or b;
    outputs(9549) <= a and b;
    outputs(9550) <= not a;
    outputs(9551) <= not (a xor b);
    outputs(9552) <= not a;
    outputs(9553) <= not a;
    outputs(9554) <= a xor b;
    outputs(9555) <= not (a xor b);
    outputs(9556) <= a xor b;
    outputs(9557) <= not (a and b);
    outputs(9558) <= not b;
    outputs(9559) <= not (a xor b);
    outputs(9560) <= b;
    outputs(9561) <= not b;
    outputs(9562) <= b;
    outputs(9563) <= not b;
    outputs(9564) <= not a;
    outputs(9565) <= a xor b;
    outputs(9566) <= not b;
    outputs(9567) <= b;
    outputs(9568) <= a and b;
    outputs(9569) <= a xor b;
    outputs(9570) <= not (a or b);
    outputs(9571) <= not a;
    outputs(9572) <= not a;
    outputs(9573) <= not (a xor b);
    outputs(9574) <= not (a and b);
    outputs(9575) <= not a;
    outputs(9576) <= a and b;
    outputs(9577) <= a xor b;
    outputs(9578) <= not a;
    outputs(9579) <= not b;
    outputs(9580) <= b;
    outputs(9581) <= a;
    outputs(9582) <= not b;
    outputs(9583) <= not (a xor b);
    outputs(9584) <= not (a xor b);
    outputs(9585) <= not b;
    outputs(9586) <= a xor b;
    outputs(9587) <= b;
    outputs(9588) <= a xor b;
    outputs(9589) <= a;
    outputs(9590) <= a and not b;
    outputs(9591) <= not (a or b);
    outputs(9592) <= b;
    outputs(9593) <= not a;
    outputs(9594) <= a and b;
    outputs(9595) <= a or b;
    outputs(9596) <= a xor b;
    outputs(9597) <= b and not a;
    outputs(9598) <= not (a xor b);
    outputs(9599) <= a xor b;
    outputs(9600) <= b;
    outputs(9601) <= not a;
    outputs(9602) <= not b;
    outputs(9603) <= a;
    outputs(9604) <= b;
    outputs(9605) <= not a;
    outputs(9606) <= a xor b;
    outputs(9607) <= not (a or b);
    outputs(9608) <= not a;
    outputs(9609) <= not a;
    outputs(9610) <= not b;
    outputs(9611) <= not a;
    outputs(9612) <= not (a and b);
    outputs(9613) <= not (a xor b);
    outputs(9614) <= not a;
    outputs(9615) <= not (a or b);
    outputs(9616) <= b;
    outputs(9617) <= a and not b;
    outputs(9618) <= a xor b;
    outputs(9619) <= not (a xor b);
    outputs(9620) <= not (a xor b);
    outputs(9621) <= a xor b;
    outputs(9622) <= not (a or b);
    outputs(9623) <= a and not b;
    outputs(9624) <= b;
    outputs(9625) <= not (a or b);
    outputs(9626) <= not (a and b);
    outputs(9627) <= b;
    outputs(9628) <= not (a or b);
    outputs(9629) <= a xor b;
    outputs(9630) <= a xor b;
    outputs(9631) <= a;
    outputs(9632) <= not (a or b);
    outputs(9633) <= not a;
    outputs(9634) <= a or b;
    outputs(9635) <= a and not b;
    outputs(9636) <= not (a xor b);
    outputs(9637) <= not (a xor b);
    outputs(9638) <= not a or b;
    outputs(9639) <= a;
    outputs(9640) <= not (a and b);
    outputs(9641) <= a and b;
    outputs(9642) <= not a;
    outputs(9643) <= not b or a;
    outputs(9644) <= a and b;
    outputs(9645) <= not (a xor b);
    outputs(9646) <= not (a xor b);
    outputs(9647) <= a xor b;
    outputs(9648) <= a xor b;
    outputs(9649) <= a and b;
    outputs(9650) <= not a;
    outputs(9651) <= a;
    outputs(9652) <= a;
    outputs(9653) <= not a;
    outputs(9654) <= not b;
    outputs(9655) <= a;
    outputs(9656) <= a;
    outputs(9657) <= a xor b;
    outputs(9658) <= a xor b;
    outputs(9659) <= not (a xor b);
    outputs(9660) <= a and b;
    outputs(9661) <= a xor b;
    outputs(9662) <= a xor b;
    outputs(9663) <= not a or b;
    outputs(9664) <= a;
    outputs(9665) <= b and not a;
    outputs(9666) <= not a;
    outputs(9667) <= not (a xor b);
    outputs(9668) <= a;
    outputs(9669) <= b and not a;
    outputs(9670) <= not b;
    outputs(9671) <= not b;
    outputs(9672) <= a xor b;
    outputs(9673) <= a xor b;
    outputs(9674) <= not b;
    outputs(9675) <= not (a xor b);
    outputs(9676) <= b and not a;
    outputs(9677) <= a and b;
    outputs(9678) <= a and not b;
    outputs(9679) <= not (a xor b);
    outputs(9680) <= b;
    outputs(9681) <= b;
    outputs(9682) <= not (a and b);
    outputs(9683) <= b;
    outputs(9684) <= not a;
    outputs(9685) <= not b;
    outputs(9686) <= not (a or b);
    outputs(9687) <= a or b;
    outputs(9688) <= not b or a;
    outputs(9689) <= a;
    outputs(9690) <= not (a xor b);
    outputs(9691) <= not (a xor b);
    outputs(9692) <= a xor b;
    outputs(9693) <= not (a and b);
    outputs(9694) <= a xor b;
    outputs(9695) <= not a;
    outputs(9696) <= not (a or b);
    outputs(9697) <= not b or a;
    outputs(9698) <= not a;
    outputs(9699) <= a or b;
    outputs(9700) <= b and not a;
    outputs(9701) <= b and not a;
    outputs(9702) <= not b;
    outputs(9703) <= not (a xor b);
    outputs(9704) <= not (a xor b);
    outputs(9705) <= a;
    outputs(9706) <= not a;
    outputs(9707) <= a and b;
    outputs(9708) <= not b;
    outputs(9709) <= b;
    outputs(9710) <= a xor b;
    outputs(9711) <= not a or b;
    outputs(9712) <= not b;
    outputs(9713) <= a xor b;
    outputs(9714) <= not a or b;
    outputs(9715) <= b;
    outputs(9716) <= a and b;
    outputs(9717) <= not b;
    outputs(9718) <= not (a xor b);
    outputs(9719) <= b;
    outputs(9720) <= a and b;
    outputs(9721) <= a xor b;
    outputs(9722) <= a xor b;
    outputs(9723) <= not b;
    outputs(9724) <= not a;
    outputs(9725) <= a;
    outputs(9726) <= not (a xor b);
    outputs(9727) <= a or b;
    outputs(9728) <= a and not b;
    outputs(9729) <= a xor b;
    outputs(9730) <= a xor b;
    outputs(9731) <= not (a or b);
    outputs(9732) <= not (a or b);
    outputs(9733) <= a or b;
    outputs(9734) <= a xor b;
    outputs(9735) <= b;
    outputs(9736) <= a and b;
    outputs(9737) <= not a or b;
    outputs(9738) <= a xor b;
    outputs(9739) <= b;
    outputs(9740) <= a xor b;
    outputs(9741) <= not (a and b);
    outputs(9742) <= a or b;
    outputs(9743) <= not (a or b);
    outputs(9744) <= not b;
    outputs(9745) <= b;
    outputs(9746) <= a;
    outputs(9747) <= not (a or b);
    outputs(9748) <= b;
    outputs(9749) <= not (a xor b);
    outputs(9750) <= a xor b;
    outputs(9751) <= not (a and b);
    outputs(9752) <= a and not b;
    outputs(9753) <= a;
    outputs(9754) <= not b;
    outputs(9755) <= not (a and b);
    outputs(9756) <= not b;
    outputs(9757) <= a and not b;
    outputs(9758) <= a;
    outputs(9759) <= a xor b;
    outputs(9760) <= not b;
    outputs(9761) <= b;
    outputs(9762) <= a;
    outputs(9763) <= b;
    outputs(9764) <= not (a or b);
    outputs(9765) <= not b;
    outputs(9766) <= not a;
    outputs(9767) <= a;
    outputs(9768) <= not b;
    outputs(9769) <= b;
    outputs(9770) <= not b;
    outputs(9771) <= not a;
    outputs(9772) <= a xor b;
    outputs(9773) <= a xor b;
    outputs(9774) <= a and b;
    outputs(9775) <= not a;
    outputs(9776) <= a and b;
    outputs(9777) <= a and b;
    outputs(9778) <= not a;
    outputs(9779) <= not b or a;
    outputs(9780) <= not (a or b);
    outputs(9781) <= a xor b;
    outputs(9782) <= not (a or b);
    outputs(9783) <= not (a xor b);
    outputs(9784) <= a and not b;
    outputs(9785) <= not (a xor b);
    outputs(9786) <= not b;
    outputs(9787) <= not (a xor b);
    outputs(9788) <= not (a xor b);
    outputs(9789) <= a xor b;
    outputs(9790) <= not (a xor b);
    outputs(9791) <= a and not b;
    outputs(9792) <= b;
    outputs(9793) <= a and not b;
    outputs(9794) <= a or b;
    outputs(9795) <= a xor b;
    outputs(9796) <= a;
    outputs(9797) <= a xor b;
    outputs(9798) <= not (a or b);
    outputs(9799) <= a xor b;
    outputs(9800) <= a xor b;
    outputs(9801) <= b;
    outputs(9802) <= b;
    outputs(9803) <= b;
    outputs(9804) <= b and not a;
    outputs(9805) <= b;
    outputs(9806) <= not (a xor b);
    outputs(9807) <= not b;
    outputs(9808) <= a xor b;
    outputs(9809) <= a and b;
    outputs(9810) <= not b;
    outputs(9811) <= not (a or b);
    outputs(9812) <= not a;
    outputs(9813) <= not a or b;
    outputs(9814) <= b;
    outputs(9815) <= a and b;
    outputs(9816) <= a xor b;
    outputs(9817) <= not (a xor b);
    outputs(9818) <= b;
    outputs(9819) <= b and not a;
    outputs(9820) <= b and not a;
    outputs(9821) <= not a;
    outputs(9822) <= b;
    outputs(9823) <= not (a xor b);
    outputs(9824) <= not (a and b);
    outputs(9825) <= a xor b;
    outputs(9826) <= not (a xor b);
    outputs(9827) <= a xor b;
    outputs(9828) <= not (a xor b);
    outputs(9829) <= a xor b;
    outputs(9830) <= a xor b;
    outputs(9831) <= a;
    outputs(9832) <= not b or a;
    outputs(9833) <= not b;
    outputs(9834) <= not (a and b);
    outputs(9835) <= b;
    outputs(9836) <= not a;
    outputs(9837) <= not (a xor b);
    outputs(9838) <= not (a or b);
    outputs(9839) <= a xor b;
    outputs(9840) <= not (a xor b);
    outputs(9841) <= a xor b;
    outputs(9842) <= not b;
    outputs(9843) <= not (a or b);
    outputs(9844) <= a xor b;
    outputs(9845) <= not a;
    outputs(9846) <= a and not b;
    outputs(9847) <= b;
    outputs(9848) <= a;
    outputs(9849) <= not a;
    outputs(9850) <= a or b;
    outputs(9851) <= b and not a;
    outputs(9852) <= a and not b;
    outputs(9853) <= a xor b;
    outputs(9854) <= not (a xor b);
    outputs(9855) <= a and b;
    outputs(9856) <= a;
    outputs(9857) <= not b;
    outputs(9858) <= not (a or b);
    outputs(9859) <= a;
    outputs(9860) <= b and not a;
    outputs(9861) <= not a;
    outputs(9862) <= not a;
    outputs(9863) <= not (a xor b);
    outputs(9864) <= not a;
    outputs(9865) <= a xor b;
    outputs(9866) <= a or b;
    outputs(9867) <= not (a and b);
    outputs(9868) <= a xor b;
    outputs(9869) <= a and b;
    outputs(9870) <= b;
    outputs(9871) <= a and not b;
    outputs(9872) <= b;
    outputs(9873) <= b and not a;
    outputs(9874) <= not b;
    outputs(9875) <= not a;
    outputs(9876) <= b;
    outputs(9877) <= a;
    outputs(9878) <= not a;
    outputs(9879) <= not (a xor b);
    outputs(9880) <= a and not b;
    outputs(9881) <= a;
    outputs(9882) <= b and not a;
    outputs(9883) <= a;
    outputs(9884) <= not (a and b);
    outputs(9885) <= a;
    outputs(9886) <= b;
    outputs(9887) <= not (a xor b);
    outputs(9888) <= a xor b;
    outputs(9889) <= a xor b;
    outputs(9890) <= not a;
    outputs(9891) <= a;
    outputs(9892) <= not (a xor b);
    outputs(9893) <= not b;
    outputs(9894) <= a xor b;
    outputs(9895) <= not (a and b);
    outputs(9896) <= not b;
    outputs(9897) <= a and b;
    outputs(9898) <= b;
    outputs(9899) <= not (a or b);
    outputs(9900) <= a xor b;
    outputs(9901) <= not (a xor b);
    outputs(9902) <= b;
    outputs(9903) <= a xor b;
    outputs(9904) <= a;
    outputs(9905) <= not b;
    outputs(9906) <= b;
    outputs(9907) <= not (a xor b);
    outputs(9908) <= a xor b;
    outputs(9909) <= not (a xor b);
    outputs(9910) <= not b;
    outputs(9911) <= a or b;
    outputs(9912) <= b and not a;
    outputs(9913) <= not a;
    outputs(9914) <= a xor b;
    outputs(9915) <= not b;
    outputs(9916) <= not (a xor b);
    outputs(9917) <= a;
    outputs(9918) <= b;
    outputs(9919) <= not b or a;
    outputs(9920) <= not b;
    outputs(9921) <= a xor b;
    outputs(9922) <= a;
    outputs(9923) <= a and b;
    outputs(9924) <= a;
    outputs(9925) <= a or b;
    outputs(9926) <= a xor b;
    outputs(9927) <= b;
    outputs(9928) <= a and not b;
    outputs(9929) <= not (a and b);
    outputs(9930) <= a and b;
    outputs(9931) <= a xor b;
    outputs(9932) <= not (a xor b);
    outputs(9933) <= a xor b;
    outputs(9934) <= a;
    outputs(9935) <= not a;
    outputs(9936) <= a xor b;
    outputs(9937) <= b;
    outputs(9938) <= b;
    outputs(9939) <= a xor b;
    outputs(9940) <= b and not a;
    outputs(9941) <= a;
    outputs(9942) <= not (a xor b);
    outputs(9943) <= not (a xor b);
    outputs(9944) <= a xor b;
    outputs(9945) <= not b;
    outputs(9946) <= not b;
    outputs(9947) <= not b;
    outputs(9948) <= not (a xor b);
    outputs(9949) <= not (a xor b);
    outputs(9950) <= not (a xor b);
    outputs(9951) <= a and not b;
    outputs(9952) <= not a;
    outputs(9953) <= not a;
    outputs(9954) <= b and not a;
    outputs(9955) <= a and b;
    outputs(9956) <= not (a and b);
    outputs(9957) <= b;
    outputs(9958) <= a xor b;
    outputs(9959) <= not a;
    outputs(9960) <= b and not a;
    outputs(9961) <= a;
    outputs(9962) <= not b;
    outputs(9963) <= not a;
    outputs(9964) <= not (a xor b);
    outputs(9965) <= a xor b;
    outputs(9966) <= not (a xor b);
    outputs(9967) <= not (a xor b);
    outputs(9968) <= a xor b;
    outputs(9969) <= a;
    outputs(9970) <= b;
    outputs(9971) <= not b;
    outputs(9972) <= b and not a;
    outputs(9973) <= not (a xor b);
    outputs(9974) <= b and not a;
    outputs(9975) <= b;
    outputs(9976) <= a xor b;
    outputs(9977) <= b;
    outputs(9978) <= not a;
    outputs(9979) <= b;
    outputs(9980) <= b;
    outputs(9981) <= not a;
    outputs(9982) <= b and not a;
    outputs(9983) <= not a;
    outputs(9984) <= b and not a;
    outputs(9985) <= a;
    outputs(9986) <= a;
    outputs(9987) <= b;
    outputs(9988) <= not b or a;
    outputs(9989) <= a;
    outputs(9990) <= a;
    outputs(9991) <= not b or a;
    outputs(9992) <= not a or b;
    outputs(9993) <= a and not b;
    outputs(9994) <= a xor b;
    outputs(9995) <= not (a or b);
    outputs(9996) <= a;
    outputs(9997) <= not b;
    outputs(9998) <= not a;
    outputs(9999) <= a;
    outputs(10000) <= not (a xor b);
    outputs(10001) <= not (a xor b);
    outputs(10002) <= not b;
    outputs(10003) <= not (a xor b);
    outputs(10004) <= not a or b;
    outputs(10005) <= a xor b;
    outputs(10006) <= not (a xor b);
    outputs(10007) <= a;
    outputs(10008) <= a and b;
    outputs(10009) <= not (a and b);
    outputs(10010) <= not (a or b);
    outputs(10011) <= a and b;
    outputs(10012) <= not a;
    outputs(10013) <= not b;
    outputs(10014) <= a xor b;
    outputs(10015) <= a;
    outputs(10016) <= not b;
    outputs(10017) <= a;
    outputs(10018) <= not b;
    outputs(10019) <= a;
    outputs(10020) <= not (a and b);
    outputs(10021) <= b;
    outputs(10022) <= not (a or b);
    outputs(10023) <= a;
    outputs(10024) <= a and not b;
    outputs(10025) <= not a or b;
    outputs(10026) <= not (a xor b);
    outputs(10027) <= a xor b;
    outputs(10028) <= b;
    outputs(10029) <= b;
    outputs(10030) <= not b;
    outputs(10031) <= b;
    outputs(10032) <= not (a and b);
    outputs(10033) <= a xor b;
    outputs(10034) <= not (a or b);
    outputs(10035) <= a;
    outputs(10036) <= b and not a;
    outputs(10037) <= a and not b;
    outputs(10038) <= a;
    outputs(10039) <= not (a or b);
    outputs(10040) <= not a;
    outputs(10041) <= not (a or b);
    outputs(10042) <= a xor b;
    outputs(10043) <= not b or a;
    outputs(10044) <= b;
    outputs(10045) <= not (a and b);
    outputs(10046) <= a and not b;
    outputs(10047) <= b and not a;
    outputs(10048) <= b;
    outputs(10049) <= not b;
    outputs(10050) <= not (a xor b);
    outputs(10051) <= not a;
    outputs(10052) <= not (a and b);
    outputs(10053) <= a xor b;
    outputs(10054) <= not (a or b);
    outputs(10055) <= not (a or b);
    outputs(10056) <= a;
    outputs(10057) <= a xor b;
    outputs(10058) <= not a;
    outputs(10059) <= b;
    outputs(10060) <= not b;
    outputs(10061) <= not (a xor b);
    outputs(10062) <= not (a xor b);
    outputs(10063) <= not (a xor b);
    outputs(10064) <= not b or a;
    outputs(10065) <= not a or b;
    outputs(10066) <= a and b;
    outputs(10067) <= not (a or b);
    outputs(10068) <= a xor b;
    outputs(10069) <= a xor b;
    outputs(10070) <= a xor b;
    outputs(10071) <= a xor b;
    outputs(10072) <= not (a xor b);
    outputs(10073) <= not b;
    outputs(10074) <= b;
    outputs(10075) <= not b;
    outputs(10076) <= not a or b;
    outputs(10077) <= not (a or b);
    outputs(10078) <= a;
    outputs(10079) <= not (a xor b);
    outputs(10080) <= not (a xor b);
    outputs(10081) <= b and not a;
    outputs(10082) <= a xor b;
    outputs(10083) <= b and not a;
    outputs(10084) <= not a;
    outputs(10085) <= a xor b;
    outputs(10086) <= not b;
    outputs(10087) <= a;
    outputs(10088) <= not (a xor b);
    outputs(10089) <= not a or b;
    outputs(10090) <= not a;
    outputs(10091) <= not b;
    outputs(10092) <= not (a xor b);
    outputs(10093) <= a and b;
    outputs(10094) <= not a;
    outputs(10095) <= not a;
    outputs(10096) <= not a;
    outputs(10097) <= not (a xor b);
    outputs(10098) <= not b or a;
    outputs(10099) <= not (a or b);
    outputs(10100) <= not a;
    outputs(10101) <= a xor b;
    outputs(10102) <= b and not a;
    outputs(10103) <= not a;
    outputs(10104) <= not (a xor b);
    outputs(10105) <= b;
    outputs(10106) <= a and not b;
    outputs(10107) <= not (a and b);
    outputs(10108) <= not (a xor b);
    outputs(10109) <= not b or a;
    outputs(10110) <= a and b;
    outputs(10111) <= b and not a;
    outputs(10112) <= a;
    outputs(10113) <= a xor b;
    outputs(10114) <= not b;
    outputs(10115) <= not (a xor b);
    outputs(10116) <= not a or b;
    outputs(10117) <= not a or b;
    outputs(10118) <= not a;
    outputs(10119) <= not b or a;
    outputs(10120) <= not (a or b);
    outputs(10121) <= not a;
    outputs(10122) <= not (a or b);
    outputs(10123) <= b;
    outputs(10124) <= not a or b;
    outputs(10125) <= not a;
    outputs(10126) <= not (a xor b);
    outputs(10127) <= not (a xor b);
    outputs(10128) <= b and not a;
    outputs(10129) <= not (a or b);
    outputs(10130) <= a;
    outputs(10131) <= a xor b;
    outputs(10132) <= not (a xor b);
    outputs(10133) <= not a;
    outputs(10134) <= b;
    outputs(10135) <= not (a xor b);
    outputs(10136) <= not b;
    outputs(10137) <= a xor b;
    outputs(10138) <= not (a or b);
    outputs(10139) <= a and b;
    outputs(10140) <= b;
    outputs(10141) <= a xor b;
    outputs(10142) <= b;
    outputs(10143) <= a and b;
    outputs(10144) <= b and not a;
    outputs(10145) <= b;
    outputs(10146) <= not b or a;
    outputs(10147) <= a;
    outputs(10148) <= not (a xor b);
    outputs(10149) <= not b;
    outputs(10150) <= not b;
    outputs(10151) <= not (a xor b);
    outputs(10152) <= not a;
    outputs(10153) <= not b;
    outputs(10154) <= not a;
    outputs(10155) <= not (a or b);
    outputs(10156) <= b;
    outputs(10157) <= not (a xor b);
    outputs(10158) <= a;
    outputs(10159) <= not (a and b);
    outputs(10160) <= b;
    outputs(10161) <= not a;
    outputs(10162) <= b;
    outputs(10163) <= not b;
    outputs(10164) <= not (a xor b);
    outputs(10165) <= b;
    outputs(10166) <= not b;
    outputs(10167) <= a xor b;
    outputs(10168) <= not (a xor b);
    outputs(10169) <= a and not b;
    outputs(10170) <= not b;
    outputs(10171) <= not a;
    outputs(10172) <= not a;
    outputs(10173) <= b;
    outputs(10174) <= not (a xor b);
    outputs(10175) <= not (a or b);
    outputs(10176) <= a or b;
    outputs(10177) <= a and b;
    outputs(10178) <= not (a xor b);
    outputs(10179) <= not (a or b);
    outputs(10180) <= a;
    outputs(10181) <= b;
    outputs(10182) <= a xor b;
    outputs(10183) <= a;
    outputs(10184) <= b and not a;
    outputs(10185) <= not b or a;
    outputs(10186) <= b and not a;
    outputs(10187) <= not (a or b);
    outputs(10188) <= not a;
    outputs(10189) <= not (a xor b);
    outputs(10190) <= b and not a;
    outputs(10191) <= not b;
    outputs(10192) <= a;
    outputs(10193) <= not (a or b);
    outputs(10194) <= b and not a;
    outputs(10195) <= not (a and b);
    outputs(10196) <= a xor b;
    outputs(10197) <= not (a xor b);
    outputs(10198) <= not (a xor b);
    outputs(10199) <= b;
    outputs(10200) <= b;
    outputs(10201) <= b and not a;
    outputs(10202) <= a xor b;
    outputs(10203) <= not a;
    outputs(10204) <= not (a or b);
    outputs(10205) <= b and not a;
    outputs(10206) <= b;
    outputs(10207) <= not b;
    outputs(10208) <= b;
    outputs(10209) <= a;
    outputs(10210) <= b and not a;
    outputs(10211) <= b and not a;
    outputs(10212) <= not (a or b);
    outputs(10213) <= b;
    outputs(10214) <= b;
    outputs(10215) <= a and b;
    outputs(10216) <= not a;
    outputs(10217) <= b;
    outputs(10218) <= a xor b;
    outputs(10219) <= a;
    outputs(10220) <= not b;
    outputs(10221) <= a xor b;
    outputs(10222) <= b;
    outputs(10223) <= a;
    outputs(10224) <= not a;
    outputs(10225) <= not b;
    outputs(10226) <= not b;
    outputs(10227) <= not b;
    outputs(10228) <= a xor b;
    outputs(10229) <= a;
    outputs(10230) <= not (a or b);
    outputs(10231) <= not a;
    outputs(10232) <= a xor b;
    outputs(10233) <= not b or a;
    outputs(10234) <= b and not a;
    outputs(10235) <= a xor b;
    outputs(10236) <= b;
    outputs(10237) <= a;
    outputs(10238) <= a;
    outputs(10239) <= a;
end Behavioral;
