library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(12799 downto 0);

begin

    layer0_outputs(0) <= not(inputs(74));
    layer0_outputs(1) <= not((inputs(53)) xor (inputs(45)));
    layer0_outputs(2) <= not(inputs(43)) or (inputs(19));
    layer0_outputs(3) <= (inputs(228)) or (inputs(173));
    layer0_outputs(4) <= not(inputs(39)) or (inputs(33));
    layer0_outputs(5) <= (inputs(15)) xor (inputs(4));
    layer0_outputs(6) <= '0';
    layer0_outputs(7) <= '1';
    layer0_outputs(8) <= not(inputs(251)) or (inputs(45));
    layer0_outputs(9) <= not(inputs(153));
    layer0_outputs(10) <= (inputs(137)) or (inputs(167));
    layer0_outputs(11) <= (inputs(0)) or (inputs(153));
    layer0_outputs(12) <= (inputs(237)) or (inputs(24));
    layer0_outputs(13) <= not((inputs(253)) or (inputs(85)));
    layer0_outputs(14) <= not(inputs(50)) or (inputs(225));
    layer0_outputs(15) <= (inputs(213)) or (inputs(192));
    layer0_outputs(16) <= inputs(192);
    layer0_outputs(17) <= not(inputs(219));
    layer0_outputs(18) <= (inputs(8)) and (inputs(53));
    layer0_outputs(19) <= not(inputs(229));
    layer0_outputs(20) <= not((inputs(177)) xor (inputs(209)));
    layer0_outputs(21) <= not((inputs(50)) or (inputs(171)));
    layer0_outputs(22) <= (inputs(37)) xor (inputs(119));
    layer0_outputs(23) <= (inputs(209)) xor (inputs(114));
    layer0_outputs(24) <= (inputs(155)) and not (inputs(33));
    layer0_outputs(25) <= not(inputs(121)) or (inputs(178));
    layer0_outputs(26) <= not((inputs(173)) xor (inputs(240)));
    layer0_outputs(27) <= (inputs(201)) or (inputs(254));
    layer0_outputs(28) <= not(inputs(232));
    layer0_outputs(29) <= not((inputs(52)) and (inputs(107)));
    layer0_outputs(30) <= (inputs(96)) xor (inputs(72));
    layer0_outputs(31) <= (inputs(247)) and not (inputs(176));
    layer0_outputs(32) <= (inputs(206)) or (inputs(150));
    layer0_outputs(33) <= not((inputs(67)) or (inputs(168)));
    layer0_outputs(34) <= (inputs(140)) or (inputs(14));
    layer0_outputs(35) <= not((inputs(188)) or (inputs(141)));
    layer0_outputs(36) <= not(inputs(223)) or (inputs(34));
    layer0_outputs(37) <= not((inputs(83)) or (inputs(255)));
    layer0_outputs(38) <= (inputs(188)) and not (inputs(95));
    layer0_outputs(39) <= inputs(168);
    layer0_outputs(40) <= inputs(162);
    layer0_outputs(41) <= inputs(192);
    layer0_outputs(42) <= not((inputs(199)) xor (inputs(30)));
    layer0_outputs(43) <= (inputs(108)) or (inputs(223));
    layer0_outputs(44) <= (inputs(58)) or (inputs(130));
    layer0_outputs(45) <= not((inputs(147)) xor (inputs(81)));
    layer0_outputs(46) <= (inputs(64)) or (inputs(27));
    layer0_outputs(47) <= (inputs(46)) and not (inputs(223));
    layer0_outputs(48) <= (inputs(195)) or (inputs(189));
    layer0_outputs(49) <= not((inputs(142)) xor (inputs(20)));
    layer0_outputs(50) <= not(inputs(48)) or (inputs(115));
    layer0_outputs(51) <= not((inputs(92)) xor (inputs(13)));
    layer0_outputs(52) <= not((inputs(241)) or (inputs(13)));
    layer0_outputs(53) <= not((inputs(25)) or (inputs(254)));
    layer0_outputs(54) <= (inputs(10)) and not (inputs(205));
    layer0_outputs(55) <= (inputs(89)) and not (inputs(141));
    layer0_outputs(56) <= not((inputs(32)) or (inputs(61)));
    layer0_outputs(57) <= not((inputs(33)) xor (inputs(209)));
    layer0_outputs(58) <= (inputs(34)) or (inputs(60));
    layer0_outputs(59) <= not(inputs(173));
    layer0_outputs(60) <= (inputs(195)) and not (inputs(207));
    layer0_outputs(61) <= not((inputs(58)) or (inputs(67)));
    layer0_outputs(62) <= (inputs(245)) and not (inputs(47));
    layer0_outputs(63) <= not(inputs(246)) or (inputs(145));
    layer0_outputs(64) <= (inputs(179)) and (inputs(59));
    layer0_outputs(65) <= not(inputs(36));
    layer0_outputs(66) <= (inputs(87)) and not (inputs(34));
    layer0_outputs(67) <= not(inputs(182));
    layer0_outputs(68) <= inputs(8);
    layer0_outputs(69) <= (inputs(125)) xor (inputs(3));
    layer0_outputs(70) <= inputs(180);
    layer0_outputs(71) <= '0';
    layer0_outputs(72) <= not((inputs(98)) or (inputs(241)));
    layer0_outputs(73) <= (inputs(194)) or (inputs(220));
    layer0_outputs(74) <= inputs(213);
    layer0_outputs(75) <= not(inputs(4));
    layer0_outputs(76) <= not(inputs(232));
    layer0_outputs(77) <= (inputs(163)) xor (inputs(125));
    layer0_outputs(78) <= (inputs(55)) and not (inputs(204));
    layer0_outputs(79) <= not(inputs(145)) or (inputs(64));
    layer0_outputs(80) <= not((inputs(226)) or (inputs(6)));
    layer0_outputs(81) <= (inputs(77)) or (inputs(92));
    layer0_outputs(82) <= inputs(248);
    layer0_outputs(83) <= (inputs(235)) or (inputs(3));
    layer0_outputs(84) <= not((inputs(255)) xor (inputs(86)));
    layer0_outputs(85) <= not((inputs(82)) xor (inputs(102)));
    layer0_outputs(86) <= not(inputs(121));
    layer0_outputs(87) <= inputs(103);
    layer0_outputs(88) <= not(inputs(195)) or (inputs(110));
    layer0_outputs(89) <= inputs(130);
    layer0_outputs(90) <= not(inputs(131));
    layer0_outputs(91) <= not((inputs(180)) xor (inputs(149)));
    layer0_outputs(92) <= (inputs(112)) and not (inputs(91));
    layer0_outputs(93) <= (inputs(72)) and not (inputs(132));
    layer0_outputs(94) <= not((inputs(254)) or (inputs(195)));
    layer0_outputs(95) <= not((inputs(8)) xor (inputs(120)));
    layer0_outputs(96) <= not(inputs(65)) or (inputs(167));
    layer0_outputs(97) <= not((inputs(236)) or (inputs(223)));
    layer0_outputs(98) <= (inputs(100)) and not (inputs(244));
    layer0_outputs(99) <= not(inputs(106));
    layer0_outputs(100) <= not(inputs(206));
    layer0_outputs(101) <= not(inputs(115));
    layer0_outputs(102) <= (inputs(239)) or (inputs(168));
    layer0_outputs(103) <= (inputs(216)) and not (inputs(70));
    layer0_outputs(104) <= inputs(148);
    layer0_outputs(105) <= (inputs(74)) and not (inputs(36));
    layer0_outputs(106) <= inputs(69);
    layer0_outputs(107) <= (inputs(1)) or (inputs(231));
    layer0_outputs(108) <= not((inputs(158)) or (inputs(187)));
    layer0_outputs(109) <= not(inputs(53)) or (inputs(189));
    layer0_outputs(110) <= not((inputs(52)) xor (inputs(209)));
    layer0_outputs(111) <= not((inputs(43)) xor (inputs(31)));
    layer0_outputs(112) <= not(inputs(5));
    layer0_outputs(113) <= (inputs(23)) and not (inputs(243));
    layer0_outputs(114) <= inputs(29);
    layer0_outputs(115) <= not(inputs(234));
    layer0_outputs(116) <= inputs(74);
    layer0_outputs(117) <= (inputs(129)) xor (inputs(229));
    layer0_outputs(118) <= (inputs(247)) xor (inputs(188));
    layer0_outputs(119) <= not((inputs(112)) or (inputs(108)));
    layer0_outputs(120) <= (inputs(197)) xor (inputs(81));
    layer0_outputs(121) <= not((inputs(4)) or (inputs(184)));
    layer0_outputs(122) <= (inputs(86)) xor (inputs(200));
    layer0_outputs(123) <= not(inputs(182));
    layer0_outputs(124) <= (inputs(238)) or (inputs(130));
    layer0_outputs(125) <= (inputs(3)) xor (inputs(128));
    layer0_outputs(126) <= inputs(91);
    layer0_outputs(127) <= (inputs(163)) or (inputs(65));
    layer0_outputs(128) <= not((inputs(155)) xor (inputs(169)));
    layer0_outputs(129) <= (inputs(132)) or (inputs(46));
    layer0_outputs(130) <= (inputs(254)) or (inputs(151));
    layer0_outputs(131) <= inputs(198);
    layer0_outputs(132) <= not(inputs(192)) or (inputs(73));
    layer0_outputs(133) <= not((inputs(28)) or (inputs(147)));
    layer0_outputs(134) <= inputs(173);
    layer0_outputs(135) <= (inputs(224)) or (inputs(39));
    layer0_outputs(136) <= (inputs(86)) xor (inputs(65));
    layer0_outputs(137) <= not(inputs(102));
    layer0_outputs(138) <= (inputs(96)) xor (inputs(34));
    layer0_outputs(139) <= not((inputs(2)) or (inputs(241)));
    layer0_outputs(140) <= inputs(219);
    layer0_outputs(141) <= inputs(216);
    layer0_outputs(142) <= not(inputs(207));
    layer0_outputs(143) <= (inputs(187)) or (inputs(219));
    layer0_outputs(144) <= (inputs(93)) and (inputs(1));
    layer0_outputs(145) <= inputs(13);
    layer0_outputs(146) <= inputs(230);
    layer0_outputs(147) <= not((inputs(0)) or (inputs(9)));
    layer0_outputs(148) <= not((inputs(35)) or (inputs(129)));
    layer0_outputs(149) <= '1';
    layer0_outputs(150) <= inputs(5);
    layer0_outputs(151) <= not((inputs(194)) or (inputs(162)));
    layer0_outputs(152) <= inputs(83);
    layer0_outputs(153) <= inputs(57);
    layer0_outputs(154) <= not((inputs(168)) and (inputs(89)));
    layer0_outputs(155) <= (inputs(140)) and not (inputs(65));
    layer0_outputs(156) <= (inputs(209)) xor (inputs(32));
    layer0_outputs(157) <= not(inputs(83));
    layer0_outputs(158) <= not(inputs(189));
    layer0_outputs(159) <= inputs(61);
    layer0_outputs(160) <= (inputs(110)) or (inputs(68));
    layer0_outputs(161) <= not(inputs(227)) or (inputs(127));
    layer0_outputs(162) <= (inputs(143)) or (inputs(31));
    layer0_outputs(163) <= not((inputs(132)) or (inputs(47)));
    layer0_outputs(164) <= not((inputs(186)) xor (inputs(234)));
    layer0_outputs(165) <= inputs(3);
    layer0_outputs(166) <= inputs(103);
    layer0_outputs(167) <= not((inputs(150)) xor (inputs(212)));
    layer0_outputs(168) <= '0';
    layer0_outputs(169) <= not(inputs(59)) or (inputs(174));
    layer0_outputs(170) <= not(inputs(84));
    layer0_outputs(171) <= not(inputs(101));
    layer0_outputs(172) <= inputs(66);
    layer0_outputs(173) <= not(inputs(144));
    layer0_outputs(174) <= not(inputs(197));
    layer0_outputs(175) <= not(inputs(29)) or (inputs(195));
    layer0_outputs(176) <= not((inputs(37)) or (inputs(77)));
    layer0_outputs(177) <= not((inputs(48)) xor (inputs(4)));
    layer0_outputs(178) <= not((inputs(75)) or (inputs(77)));
    layer0_outputs(179) <= not((inputs(70)) or (inputs(5)));
    layer0_outputs(180) <= not(inputs(45)) or (inputs(194));
    layer0_outputs(181) <= (inputs(151)) and not (inputs(138));
    layer0_outputs(182) <= not((inputs(77)) or (inputs(36)));
    layer0_outputs(183) <= not((inputs(196)) and (inputs(156)));
    layer0_outputs(184) <= not((inputs(102)) xor (inputs(114)));
    layer0_outputs(185) <= (inputs(64)) and (inputs(70));
    layer0_outputs(186) <= inputs(135);
    layer0_outputs(187) <= not((inputs(176)) xor (inputs(139)));
    layer0_outputs(188) <= not(inputs(83));
    layer0_outputs(189) <= not(inputs(90)) or (inputs(0));
    layer0_outputs(190) <= not((inputs(13)) or (inputs(184)));
    layer0_outputs(191) <= (inputs(157)) and not (inputs(47));
    layer0_outputs(192) <= (inputs(58)) or (inputs(122));
    layer0_outputs(193) <= (inputs(127)) or (inputs(79));
    layer0_outputs(194) <= not(inputs(231));
    layer0_outputs(195) <= not((inputs(227)) xor (inputs(204)));
    layer0_outputs(196) <= not(inputs(23));
    layer0_outputs(197) <= (inputs(193)) or (inputs(238));
    layer0_outputs(198) <= (inputs(250)) xor (inputs(220));
    layer0_outputs(199) <= (inputs(107)) and not (inputs(33));
    layer0_outputs(200) <= inputs(120);
    layer0_outputs(201) <= (inputs(38)) and not (inputs(212));
    layer0_outputs(202) <= (inputs(153)) and (inputs(30));
    layer0_outputs(203) <= not((inputs(145)) xor (inputs(166)));
    layer0_outputs(204) <= '1';
    layer0_outputs(205) <= inputs(76);
    layer0_outputs(206) <= (inputs(62)) xor (inputs(73));
    layer0_outputs(207) <= inputs(34);
    layer0_outputs(208) <= inputs(86);
    layer0_outputs(209) <= (inputs(120)) xor (inputs(236));
    layer0_outputs(210) <= not((inputs(184)) or (inputs(237)));
    layer0_outputs(211) <= (inputs(231)) and not (inputs(163));
    layer0_outputs(212) <= not(inputs(56));
    layer0_outputs(213) <= inputs(177);
    layer0_outputs(214) <= not(inputs(249));
    layer0_outputs(215) <= '1';
    layer0_outputs(216) <= (inputs(165)) or (inputs(250));
    layer0_outputs(217) <= not((inputs(137)) or (inputs(6)));
    layer0_outputs(218) <= not(inputs(52)) or (inputs(198));
    layer0_outputs(219) <= (inputs(190)) and not (inputs(200));
    layer0_outputs(220) <= not(inputs(57));
    layer0_outputs(221) <= (inputs(176)) or (inputs(246));
    layer0_outputs(222) <= (inputs(86)) xor (inputs(24));
    layer0_outputs(223) <= inputs(35);
    layer0_outputs(224) <= inputs(126);
    layer0_outputs(225) <= '1';
    layer0_outputs(226) <= (inputs(80)) and not (inputs(14));
    layer0_outputs(227) <= not(inputs(196)) or (inputs(62));
    layer0_outputs(228) <= not((inputs(119)) xor (inputs(157)));
    layer0_outputs(229) <= inputs(78);
    layer0_outputs(230) <= (inputs(8)) xor (inputs(54));
    layer0_outputs(231) <= not((inputs(104)) xor (inputs(42)));
    layer0_outputs(232) <= (inputs(203)) and not (inputs(114));
    layer0_outputs(233) <= not((inputs(68)) and (inputs(25)));
    layer0_outputs(234) <= not((inputs(72)) and (inputs(207)));
    layer0_outputs(235) <= not(inputs(72));
    layer0_outputs(236) <= not(inputs(222));
    layer0_outputs(237) <= not(inputs(201));
    layer0_outputs(238) <= inputs(104);
    layer0_outputs(239) <= not(inputs(114));
    layer0_outputs(240) <= (inputs(26)) and not (inputs(246));
    layer0_outputs(241) <= (inputs(110)) xor (inputs(84));
    layer0_outputs(242) <= not(inputs(102));
    layer0_outputs(243) <= not((inputs(187)) xor (inputs(1)));
    layer0_outputs(244) <= (inputs(101)) and not (inputs(208));
    layer0_outputs(245) <= not(inputs(82)) or (inputs(95));
    layer0_outputs(246) <= (inputs(4)) or (inputs(194));
    layer0_outputs(247) <= inputs(16);
    layer0_outputs(248) <= inputs(92);
    layer0_outputs(249) <= (inputs(20)) xor (inputs(71));
    layer0_outputs(250) <= (inputs(151)) and not (inputs(31));
    layer0_outputs(251) <= inputs(227);
    layer0_outputs(252) <= inputs(217);
    layer0_outputs(253) <= (inputs(16)) xor (inputs(197));
    layer0_outputs(254) <= inputs(246);
    layer0_outputs(255) <= not(inputs(53)) or (inputs(158));
    layer0_outputs(256) <= (inputs(53)) and not (inputs(251));
    layer0_outputs(257) <= (inputs(23)) or (inputs(61));
    layer0_outputs(258) <= (inputs(64)) xor (inputs(95));
    layer0_outputs(259) <= (inputs(100)) and not (inputs(239));
    layer0_outputs(260) <= inputs(213);
    layer0_outputs(261) <= '1';
    layer0_outputs(262) <= (inputs(195)) or (inputs(131));
    layer0_outputs(263) <= (inputs(246)) or (inputs(99));
    layer0_outputs(264) <= not((inputs(192)) or (inputs(138)));
    layer0_outputs(265) <= not((inputs(244)) and (inputs(246)));
    layer0_outputs(266) <= not(inputs(230)) or (inputs(237));
    layer0_outputs(267) <= (inputs(155)) and not (inputs(205));
    layer0_outputs(268) <= '0';
    layer0_outputs(269) <= (inputs(201)) or (inputs(246));
    layer0_outputs(270) <= inputs(160);
    layer0_outputs(271) <= (inputs(68)) and not (inputs(29));
    layer0_outputs(272) <= not(inputs(39)) or (inputs(220));
    layer0_outputs(273) <= not((inputs(157)) xor (inputs(11)));
    layer0_outputs(274) <= not(inputs(99));
    layer0_outputs(275) <= not(inputs(204));
    layer0_outputs(276) <= not((inputs(122)) or (inputs(225)));
    layer0_outputs(277) <= (inputs(242)) and (inputs(172));
    layer0_outputs(278) <= (inputs(73)) and (inputs(176));
    layer0_outputs(279) <= (inputs(177)) xor (inputs(232));
    layer0_outputs(280) <= not(inputs(115)) or (inputs(62));
    layer0_outputs(281) <= not(inputs(85));
    layer0_outputs(282) <= not(inputs(238)) or (inputs(159));
    layer0_outputs(283) <= inputs(166);
    layer0_outputs(284) <= inputs(194);
    layer0_outputs(285) <= inputs(200);
    layer0_outputs(286) <= not((inputs(254)) or (inputs(221)));
    layer0_outputs(287) <= not((inputs(176)) or (inputs(85)));
    layer0_outputs(288) <= not((inputs(223)) or (inputs(10)));
    layer0_outputs(289) <= (inputs(72)) xor (inputs(40));
    layer0_outputs(290) <= not(inputs(78));
    layer0_outputs(291) <= not(inputs(238));
    layer0_outputs(292) <= not(inputs(39)) or (inputs(175));
    layer0_outputs(293) <= (inputs(177)) or (inputs(192));
    layer0_outputs(294) <= not(inputs(120)) or (inputs(255));
    layer0_outputs(295) <= not(inputs(172));
    layer0_outputs(296) <= (inputs(42)) and (inputs(120));
    layer0_outputs(297) <= not(inputs(90));
    layer0_outputs(298) <= not(inputs(181));
    layer0_outputs(299) <= not(inputs(66)) or (inputs(250));
    layer0_outputs(300) <= not(inputs(69)) or (inputs(147));
    layer0_outputs(301) <= inputs(209);
    layer0_outputs(302) <= not(inputs(217)) or (inputs(235));
    layer0_outputs(303) <= (inputs(54)) and not (inputs(30));
    layer0_outputs(304) <= (inputs(128)) or (inputs(71));
    layer0_outputs(305) <= inputs(220);
    layer0_outputs(306) <= not((inputs(252)) or (inputs(195)));
    layer0_outputs(307) <= not(inputs(188)) or (inputs(99));
    layer0_outputs(308) <= (inputs(213)) and not (inputs(1));
    layer0_outputs(309) <= not((inputs(64)) or (inputs(149)));
    layer0_outputs(310) <= (inputs(61)) and not (inputs(143));
    layer0_outputs(311) <= not(inputs(165));
    layer0_outputs(312) <= '0';
    layer0_outputs(313) <= not(inputs(123));
    layer0_outputs(314) <= not(inputs(165)) or (inputs(109));
    layer0_outputs(315) <= not(inputs(135));
    layer0_outputs(316) <= inputs(211);
    layer0_outputs(317) <= not(inputs(34)) or (inputs(214));
    layer0_outputs(318) <= not(inputs(77)) or (inputs(30));
    layer0_outputs(319) <= (inputs(24)) and (inputs(117));
    layer0_outputs(320) <= (inputs(197)) xor (inputs(243));
    layer0_outputs(321) <= (inputs(66)) or (inputs(80));
    layer0_outputs(322) <= (inputs(106)) xor (inputs(236));
    layer0_outputs(323) <= (inputs(183)) or (inputs(167));
    layer0_outputs(324) <= not(inputs(219));
    layer0_outputs(325) <= (inputs(6)) or (inputs(215));
    layer0_outputs(326) <= (inputs(77)) and not (inputs(208));
    layer0_outputs(327) <= not(inputs(241));
    layer0_outputs(328) <= (inputs(6)) or (inputs(39));
    layer0_outputs(329) <= not((inputs(2)) or (inputs(202)));
    layer0_outputs(330) <= not(inputs(62));
    layer0_outputs(331) <= (inputs(63)) xor (inputs(178));
    layer0_outputs(332) <= not((inputs(145)) or (inputs(158)));
    layer0_outputs(333) <= (inputs(74)) and not (inputs(255));
    layer0_outputs(334) <= inputs(169);
    layer0_outputs(335) <= not((inputs(230)) or (inputs(151)));
    layer0_outputs(336) <= (inputs(14)) and not (inputs(224));
    layer0_outputs(337) <= (inputs(204)) and not (inputs(94));
    layer0_outputs(338) <= (inputs(8)) xor (inputs(245));
    layer0_outputs(339) <= not((inputs(128)) or (inputs(30)));
    layer0_outputs(340) <= not(inputs(181)) or (inputs(79));
    layer0_outputs(341) <= inputs(173);
    layer0_outputs(342) <= not(inputs(124));
    layer0_outputs(343) <= not((inputs(246)) or (inputs(126)));
    layer0_outputs(344) <= not((inputs(188)) xor (inputs(124)));
    layer0_outputs(345) <= not(inputs(60));
    layer0_outputs(346) <= (inputs(224)) or (inputs(42));
    layer0_outputs(347) <= not((inputs(123)) or (inputs(34)));
    layer0_outputs(348) <= (inputs(117)) and not (inputs(81));
    layer0_outputs(349) <= inputs(236);
    layer0_outputs(350) <= not((inputs(111)) xor (inputs(9)));
    layer0_outputs(351) <= inputs(26);
    layer0_outputs(352) <= not((inputs(234)) or (inputs(251)));
    layer0_outputs(353) <= (inputs(102)) and not (inputs(160));
    layer0_outputs(354) <= not((inputs(112)) xor (inputs(101)));
    layer0_outputs(355) <= (inputs(52)) or (inputs(52));
    layer0_outputs(356) <= (inputs(221)) xor (inputs(126));
    layer0_outputs(357) <= inputs(131);
    layer0_outputs(358) <= (inputs(75)) xor (inputs(13));
    layer0_outputs(359) <= inputs(59);
    layer0_outputs(360) <= (inputs(166)) and not (inputs(231));
    layer0_outputs(361) <= not((inputs(28)) xor (inputs(6)));
    layer0_outputs(362) <= not(inputs(50)) or (inputs(92));
    layer0_outputs(363) <= (inputs(93)) or (inputs(243));
    layer0_outputs(364) <= not((inputs(167)) or (inputs(182)));
    layer0_outputs(365) <= not((inputs(178)) xor (inputs(204)));
    layer0_outputs(366) <= inputs(38);
    layer0_outputs(367) <= not((inputs(164)) xor (inputs(84)));
    layer0_outputs(368) <= not(inputs(71)) or (inputs(105));
    layer0_outputs(369) <= inputs(109);
    layer0_outputs(370) <= (inputs(225)) and not (inputs(130));
    layer0_outputs(371) <= not(inputs(178)) or (inputs(34));
    layer0_outputs(372) <= not((inputs(103)) xor (inputs(242)));
    layer0_outputs(373) <= not(inputs(81));
    layer0_outputs(374) <= (inputs(186)) and not (inputs(193));
    layer0_outputs(375) <= inputs(131);
    layer0_outputs(376) <= inputs(233);
    layer0_outputs(377) <= not((inputs(253)) or (inputs(198)));
    layer0_outputs(378) <= inputs(149);
    layer0_outputs(379) <= '1';
    layer0_outputs(380) <= (inputs(169)) and not (inputs(94));
    layer0_outputs(381) <= (inputs(167)) xor (inputs(150));
    layer0_outputs(382) <= (inputs(230)) or (inputs(175));
    layer0_outputs(383) <= inputs(164);
    layer0_outputs(384) <= not(inputs(115)) or (inputs(240));
    layer0_outputs(385) <= (inputs(88)) xor (inputs(97));
    layer0_outputs(386) <= not(inputs(9));
    layer0_outputs(387) <= not(inputs(56)) or (inputs(140));
    layer0_outputs(388) <= (inputs(193)) or (inputs(46));
    layer0_outputs(389) <= (inputs(178)) xor (inputs(144));
    layer0_outputs(390) <= (inputs(7)) or (inputs(132));
    layer0_outputs(391) <= not((inputs(153)) or (inputs(254)));
    layer0_outputs(392) <= (inputs(202)) or (inputs(9));
    layer0_outputs(393) <= not((inputs(145)) xor (inputs(180)));
    layer0_outputs(394) <= not(inputs(194));
    layer0_outputs(395) <= inputs(102);
    layer0_outputs(396) <= not((inputs(109)) or (inputs(43)));
    layer0_outputs(397) <= inputs(4);
    layer0_outputs(398) <= not(inputs(155)) or (inputs(33));
    layer0_outputs(399) <= (inputs(204)) xor (inputs(224));
    layer0_outputs(400) <= not(inputs(235)) or (inputs(142));
    layer0_outputs(401) <= (inputs(61)) and not (inputs(169));
    layer0_outputs(402) <= (inputs(208)) xor (inputs(185));
    layer0_outputs(403) <= '0';
    layer0_outputs(404) <= inputs(215);
    layer0_outputs(405) <= (inputs(131)) and (inputs(57));
    layer0_outputs(406) <= not(inputs(15)) or (inputs(217));
    layer0_outputs(407) <= (inputs(162)) and not (inputs(16));
    layer0_outputs(408) <= not(inputs(53)) or (inputs(72));
    layer0_outputs(409) <= (inputs(4)) or (inputs(129));
    layer0_outputs(410) <= not(inputs(207)) or (inputs(199));
    layer0_outputs(411) <= (inputs(238)) or (inputs(106));
    layer0_outputs(412) <= (inputs(54)) xor (inputs(49));
    layer0_outputs(413) <= inputs(56);
    layer0_outputs(414) <= (inputs(210)) and (inputs(161));
    layer0_outputs(415) <= not(inputs(252));
    layer0_outputs(416) <= not((inputs(95)) or (inputs(85)));
    layer0_outputs(417) <= inputs(88);
    layer0_outputs(418) <= inputs(147);
    layer0_outputs(419) <= inputs(24);
    layer0_outputs(420) <= (inputs(27)) or (inputs(68));
    layer0_outputs(421) <= (inputs(104)) or (inputs(191));
    layer0_outputs(422) <= not(inputs(215)) or (inputs(168));
    layer0_outputs(423) <= (inputs(189)) or (inputs(44));
    layer0_outputs(424) <= inputs(142);
    layer0_outputs(425) <= not(inputs(75)) or (inputs(16));
    layer0_outputs(426) <= '1';
    layer0_outputs(427) <= not((inputs(111)) or (inputs(229)));
    layer0_outputs(428) <= (inputs(52)) or (inputs(10));
    layer0_outputs(429) <= not((inputs(255)) xor (inputs(177)));
    layer0_outputs(430) <= (inputs(247)) xor (inputs(12));
    layer0_outputs(431) <= inputs(61);
    layer0_outputs(432) <= not((inputs(148)) xor (inputs(201)));
    layer0_outputs(433) <= not((inputs(143)) and (inputs(144)));
    layer0_outputs(434) <= (inputs(153)) or (inputs(48));
    layer0_outputs(435) <= '1';
    layer0_outputs(436) <= not(inputs(75)) or (inputs(14));
    layer0_outputs(437) <= not(inputs(7)) or (inputs(247));
    layer0_outputs(438) <= (inputs(183)) xor (inputs(79));
    layer0_outputs(439) <= (inputs(157)) or (inputs(180));
    layer0_outputs(440) <= not(inputs(41)) or (inputs(178));
    layer0_outputs(441) <= (inputs(56)) and (inputs(145));
    layer0_outputs(442) <= not(inputs(231));
    layer0_outputs(443) <= inputs(94);
    layer0_outputs(444) <= not(inputs(222)) or (inputs(11));
    layer0_outputs(445) <= '1';
    layer0_outputs(446) <= inputs(60);
    layer0_outputs(447) <= inputs(23);
    layer0_outputs(448) <= not(inputs(74));
    layer0_outputs(449) <= (inputs(236)) or (inputs(3));
    layer0_outputs(450) <= '0';
    layer0_outputs(451) <= inputs(107);
    layer0_outputs(452) <= (inputs(26)) and not (inputs(178));
    layer0_outputs(453) <= not(inputs(82));
    layer0_outputs(454) <= (inputs(44)) and not (inputs(146));
    layer0_outputs(455) <= not(inputs(53));
    layer0_outputs(456) <= not(inputs(146));
    layer0_outputs(457) <= (inputs(42)) xor (inputs(240));
    layer0_outputs(458) <= not(inputs(39));
    layer0_outputs(459) <= not(inputs(43)) or (inputs(187));
    layer0_outputs(460) <= not((inputs(64)) and (inputs(19)));
    layer0_outputs(461) <= not(inputs(164)) or (inputs(31));
    layer0_outputs(462) <= not(inputs(94));
    layer0_outputs(463) <= not((inputs(26)) and (inputs(215)));
    layer0_outputs(464) <= (inputs(177)) xor (inputs(197));
    layer0_outputs(465) <= not((inputs(178)) xor (inputs(245)));
    layer0_outputs(466) <= inputs(105);
    layer0_outputs(467) <= (inputs(82)) and not (inputs(50));
    layer0_outputs(468) <= (inputs(18)) or (inputs(24));
    layer0_outputs(469) <= not((inputs(77)) or (inputs(189)));
    layer0_outputs(470) <= (inputs(199)) or (inputs(191));
    layer0_outputs(471) <= not((inputs(25)) or (inputs(207)));
    layer0_outputs(472) <= not((inputs(38)) or (inputs(78)));
    layer0_outputs(473) <= not((inputs(85)) xor (inputs(65)));
    layer0_outputs(474) <= (inputs(26)) xor (inputs(107));
    layer0_outputs(475) <= not((inputs(238)) or (inputs(213)));
    layer0_outputs(476) <= (inputs(104)) xor (inputs(166));
    layer0_outputs(477) <= not((inputs(140)) or (inputs(14)));
    layer0_outputs(478) <= (inputs(0)) xor (inputs(7));
    layer0_outputs(479) <= not((inputs(194)) or (inputs(199)));
    layer0_outputs(480) <= not(inputs(192)) or (inputs(142));
    layer0_outputs(481) <= not((inputs(231)) xor (inputs(105)));
    layer0_outputs(482) <= not(inputs(243)) or (inputs(4));
    layer0_outputs(483) <= inputs(96);
    layer0_outputs(484) <= not((inputs(33)) or (inputs(184)));
    layer0_outputs(485) <= (inputs(18)) or (inputs(111));
    layer0_outputs(486) <= (inputs(182)) or (inputs(115));
    layer0_outputs(487) <= not(inputs(35));
    layer0_outputs(488) <= inputs(136);
    layer0_outputs(489) <= not((inputs(36)) xor (inputs(51)));
    layer0_outputs(490) <= not(inputs(7));
    layer0_outputs(491) <= not(inputs(55));
    layer0_outputs(492) <= not(inputs(106));
    layer0_outputs(493) <= (inputs(12)) xor (inputs(20));
    layer0_outputs(494) <= inputs(76);
    layer0_outputs(495) <= (inputs(83)) xor (inputs(219));
    layer0_outputs(496) <= inputs(40);
    layer0_outputs(497) <= not((inputs(3)) or (inputs(94)));
    layer0_outputs(498) <= not(inputs(213)) or (inputs(125));
    layer0_outputs(499) <= (inputs(249)) and not (inputs(196));
    layer0_outputs(500) <= (inputs(36)) and not (inputs(230));
    layer0_outputs(501) <= not(inputs(38));
    layer0_outputs(502) <= not(inputs(106));
    layer0_outputs(503) <= not(inputs(103)) or (inputs(177));
    layer0_outputs(504) <= (inputs(77)) and not (inputs(203));
    layer0_outputs(505) <= (inputs(221)) or (inputs(207));
    layer0_outputs(506) <= not((inputs(24)) or (inputs(223)));
    layer0_outputs(507) <= (inputs(84)) xor (inputs(178));
    layer0_outputs(508) <= (inputs(20)) and not (inputs(144));
    layer0_outputs(509) <= inputs(102);
    layer0_outputs(510) <= not(inputs(29)) or (inputs(79));
    layer0_outputs(511) <= not((inputs(20)) xor (inputs(38)));
    layer0_outputs(512) <= (inputs(190)) or (inputs(66));
    layer0_outputs(513) <= (inputs(86)) or (inputs(247));
    layer0_outputs(514) <= not((inputs(122)) xor (inputs(93)));
    layer0_outputs(515) <= not(inputs(135)) or (inputs(111));
    layer0_outputs(516) <= not((inputs(33)) or (inputs(203)));
    layer0_outputs(517) <= (inputs(189)) or (inputs(254));
    layer0_outputs(518) <= not((inputs(23)) xor (inputs(56)));
    layer0_outputs(519) <= inputs(165);
    layer0_outputs(520) <= not(inputs(230));
    layer0_outputs(521) <= not((inputs(133)) xor (inputs(70)));
    layer0_outputs(522) <= not((inputs(22)) xor (inputs(245)));
    layer0_outputs(523) <= inputs(133);
    layer0_outputs(524) <= (inputs(110)) or (inputs(39));
    layer0_outputs(525) <= not(inputs(12)) or (inputs(91));
    layer0_outputs(526) <= not((inputs(139)) or (inputs(58)));
    layer0_outputs(527) <= not(inputs(89));
    layer0_outputs(528) <= not(inputs(167));
    layer0_outputs(529) <= not((inputs(163)) or (inputs(255)));
    layer0_outputs(530) <= not((inputs(51)) and (inputs(113)));
    layer0_outputs(531) <= (inputs(162)) xor (inputs(99));
    layer0_outputs(532) <= not(inputs(114)) or (inputs(81));
    layer0_outputs(533) <= not(inputs(75));
    layer0_outputs(534) <= not((inputs(178)) xor (inputs(252)));
    layer0_outputs(535) <= inputs(86);
    layer0_outputs(536) <= not((inputs(205)) xor (inputs(201)));
    layer0_outputs(537) <= '0';
    layer0_outputs(538) <= (inputs(193)) and not (inputs(202));
    layer0_outputs(539) <= '0';
    layer0_outputs(540) <= not(inputs(136)) or (inputs(12));
    layer0_outputs(541) <= not(inputs(149)) or (inputs(138));
    layer0_outputs(542) <= not(inputs(9));
    layer0_outputs(543) <= (inputs(92)) and (inputs(186));
    layer0_outputs(544) <= not(inputs(21));
    layer0_outputs(545) <= (inputs(253)) or (inputs(211));
    layer0_outputs(546) <= inputs(7);
    layer0_outputs(547) <= inputs(119);
    layer0_outputs(548) <= not(inputs(77));
    layer0_outputs(549) <= not(inputs(241));
    layer0_outputs(550) <= (inputs(21)) or (inputs(19));
    layer0_outputs(551) <= (inputs(171)) and not (inputs(121));
    layer0_outputs(552) <= inputs(237);
    layer0_outputs(553) <= not(inputs(42)) or (inputs(177));
    layer0_outputs(554) <= not(inputs(94));
    layer0_outputs(555) <= (inputs(105)) and not (inputs(14));
    layer0_outputs(556) <= (inputs(202)) xor (inputs(122));
    layer0_outputs(557) <= inputs(186);
    layer0_outputs(558) <= not((inputs(219)) or (inputs(90)));
    layer0_outputs(559) <= (inputs(209)) or (inputs(181));
    layer0_outputs(560) <= inputs(14);
    layer0_outputs(561) <= inputs(82);
    layer0_outputs(562) <= not(inputs(147));
    layer0_outputs(563) <= '1';
    layer0_outputs(564) <= (inputs(34)) or (inputs(218));
    layer0_outputs(565) <= not((inputs(220)) or (inputs(21)));
    layer0_outputs(566) <= not((inputs(214)) or (inputs(244)));
    layer0_outputs(567) <= inputs(105);
    layer0_outputs(568) <= (inputs(244)) or (inputs(89));
    layer0_outputs(569) <= not(inputs(191));
    layer0_outputs(570) <= not(inputs(182));
    layer0_outputs(571) <= not(inputs(136));
    layer0_outputs(572) <= inputs(96);
    layer0_outputs(573) <= inputs(116);
    layer0_outputs(574) <= inputs(88);
    layer0_outputs(575) <= (inputs(70)) xor (inputs(72));
    layer0_outputs(576) <= (inputs(187)) and not (inputs(253));
    layer0_outputs(577) <= not(inputs(54));
    layer0_outputs(578) <= inputs(65);
    layer0_outputs(579) <= (inputs(133)) xor (inputs(156));
    layer0_outputs(580) <= not((inputs(204)) or (inputs(188)));
    layer0_outputs(581) <= (inputs(32)) or (inputs(73));
    layer0_outputs(582) <= (inputs(80)) and not (inputs(138));
    layer0_outputs(583) <= (inputs(210)) xor (inputs(219));
    layer0_outputs(584) <= (inputs(212)) and not (inputs(239));
    layer0_outputs(585) <= not(inputs(93));
    layer0_outputs(586) <= (inputs(121)) and (inputs(75));
    layer0_outputs(587) <= not(inputs(47));
    layer0_outputs(588) <= not(inputs(212));
    layer0_outputs(589) <= (inputs(49)) and (inputs(175));
    layer0_outputs(590) <= not((inputs(1)) or (inputs(222)));
    layer0_outputs(591) <= '1';
    layer0_outputs(592) <= (inputs(146)) xor (inputs(97));
    layer0_outputs(593) <= inputs(208);
    layer0_outputs(594) <= not((inputs(83)) xor (inputs(158)));
    layer0_outputs(595) <= inputs(118);
    layer0_outputs(596) <= (inputs(185)) or (inputs(112));
    layer0_outputs(597) <= (inputs(228)) and not (inputs(241));
    layer0_outputs(598) <= not(inputs(129));
    layer0_outputs(599) <= not(inputs(73));
    layer0_outputs(600) <= not(inputs(101)) or (inputs(220));
    layer0_outputs(601) <= not(inputs(246));
    layer0_outputs(602) <= not((inputs(78)) or (inputs(59)));
    layer0_outputs(603) <= not((inputs(40)) or (inputs(48)));
    layer0_outputs(604) <= inputs(119);
    layer0_outputs(605) <= not((inputs(17)) xor (inputs(190)));
    layer0_outputs(606) <= not((inputs(132)) or (inputs(115)));
    layer0_outputs(607) <= not((inputs(214)) or (inputs(211)));
    layer0_outputs(608) <= not(inputs(214)) or (inputs(78));
    layer0_outputs(609) <= (inputs(92)) and (inputs(173));
    layer0_outputs(610) <= not(inputs(40)) or (inputs(189));
    layer0_outputs(611) <= not((inputs(170)) xor (inputs(48)));
    layer0_outputs(612) <= (inputs(177)) or (inputs(176));
    layer0_outputs(613) <= not((inputs(28)) and (inputs(212)));
    layer0_outputs(614) <= not(inputs(87));
    layer0_outputs(615) <= inputs(214);
    layer0_outputs(616) <= not(inputs(126));
    layer0_outputs(617) <= not(inputs(199));
    layer0_outputs(618) <= inputs(243);
    layer0_outputs(619) <= not((inputs(227)) or (inputs(94)));
    layer0_outputs(620) <= not(inputs(116)) or (inputs(125));
    layer0_outputs(621) <= inputs(114);
    layer0_outputs(622) <= not(inputs(78));
    layer0_outputs(623) <= not((inputs(206)) or (inputs(100)));
    layer0_outputs(624) <= inputs(216);
    layer0_outputs(625) <= not((inputs(34)) or (inputs(143)));
    layer0_outputs(626) <= not(inputs(75));
    layer0_outputs(627) <= (inputs(239)) or (inputs(34));
    layer0_outputs(628) <= not((inputs(30)) and (inputs(248)));
    layer0_outputs(629) <= (inputs(247)) and (inputs(253));
    layer0_outputs(630) <= not((inputs(5)) xor (inputs(176)));
    layer0_outputs(631) <= '1';
    layer0_outputs(632) <= (inputs(128)) or (inputs(55));
    layer0_outputs(633) <= not(inputs(165));
    layer0_outputs(634) <= (inputs(135)) or (inputs(175));
    layer0_outputs(635) <= (inputs(130)) xor (inputs(180));
    layer0_outputs(636) <= (inputs(77)) or (inputs(72));
    layer0_outputs(637) <= (inputs(84)) or (inputs(203));
    layer0_outputs(638) <= not(inputs(187)) or (inputs(45));
    layer0_outputs(639) <= (inputs(231)) xor (inputs(235));
    layer0_outputs(640) <= inputs(250);
    layer0_outputs(641) <= (inputs(127)) or (inputs(143));
    layer0_outputs(642) <= inputs(26);
    layer0_outputs(643) <= (inputs(106)) xor (inputs(236));
    layer0_outputs(644) <= (inputs(165)) and not (inputs(123));
    layer0_outputs(645) <= not((inputs(61)) or (inputs(201)));
    layer0_outputs(646) <= not((inputs(251)) and (inputs(188)));
    layer0_outputs(647) <= (inputs(107)) xor (inputs(182));
    layer0_outputs(648) <= not((inputs(207)) or (inputs(243)));
    layer0_outputs(649) <= inputs(11);
    layer0_outputs(650) <= (inputs(91)) and (inputs(230));
    layer0_outputs(651) <= (inputs(238)) xor (inputs(26));
    layer0_outputs(652) <= not((inputs(159)) and (inputs(187)));
    layer0_outputs(653) <= inputs(62);
    layer0_outputs(654) <= (inputs(245)) and not (inputs(13));
    layer0_outputs(655) <= not(inputs(118));
    layer0_outputs(656) <= inputs(8);
    layer0_outputs(657) <= not(inputs(248));
    layer0_outputs(658) <= not((inputs(136)) xor (inputs(233)));
    layer0_outputs(659) <= (inputs(168)) and not (inputs(26));
    layer0_outputs(660) <= not(inputs(101));
    layer0_outputs(661) <= not(inputs(30)) or (inputs(47));
    layer0_outputs(662) <= inputs(227);
    layer0_outputs(663) <= inputs(137);
    layer0_outputs(664) <= inputs(236);
    layer0_outputs(665) <= inputs(164);
    layer0_outputs(666) <= not(inputs(30));
    layer0_outputs(667) <= not((inputs(170)) or (inputs(192)));
    layer0_outputs(668) <= (inputs(247)) xor (inputs(62));
    layer0_outputs(669) <= inputs(165);
    layer0_outputs(670) <= '1';
    layer0_outputs(671) <= (inputs(155)) and not (inputs(183));
    layer0_outputs(672) <= not((inputs(66)) or (inputs(123)));
    layer0_outputs(673) <= not((inputs(156)) xor (inputs(65)));
    layer0_outputs(674) <= not(inputs(158)) or (inputs(159));
    layer0_outputs(675) <= not((inputs(192)) or (inputs(56)));
    layer0_outputs(676) <= (inputs(5)) or (inputs(186));
    layer0_outputs(677) <= not((inputs(42)) or (inputs(28)));
    layer0_outputs(678) <= (inputs(191)) and (inputs(214));
    layer0_outputs(679) <= not(inputs(64)) or (inputs(123));
    layer0_outputs(680) <= (inputs(154)) and not (inputs(175));
    layer0_outputs(681) <= not(inputs(210));
    layer0_outputs(682) <= not(inputs(39)) or (inputs(100));
    layer0_outputs(683) <= (inputs(74)) xor (inputs(208));
    layer0_outputs(684) <= (inputs(253)) or (inputs(132));
    layer0_outputs(685) <= not(inputs(13)) or (inputs(235));
    layer0_outputs(686) <= (inputs(160)) or (inputs(243));
    layer0_outputs(687) <= (inputs(41)) xor (inputs(72));
    layer0_outputs(688) <= (inputs(91)) or (inputs(170));
    layer0_outputs(689) <= not(inputs(36)) or (inputs(231));
    layer0_outputs(690) <= (inputs(138)) and not (inputs(39));
    layer0_outputs(691) <= not(inputs(73)) or (inputs(126));
    layer0_outputs(692) <= not((inputs(36)) xor (inputs(22)));
    layer0_outputs(693) <= not(inputs(126));
    layer0_outputs(694) <= not(inputs(155));
    layer0_outputs(695) <= not(inputs(90));
    layer0_outputs(696) <= not(inputs(245));
    layer0_outputs(697) <= not(inputs(232)) or (inputs(226));
    layer0_outputs(698) <= inputs(118);
    layer0_outputs(699) <= (inputs(240)) or (inputs(75));
    layer0_outputs(700) <= not((inputs(14)) xor (inputs(238)));
    layer0_outputs(701) <= not((inputs(206)) or (inputs(158)));
    layer0_outputs(702) <= not(inputs(104));
    layer0_outputs(703) <= (inputs(175)) and not (inputs(191));
    layer0_outputs(704) <= (inputs(127)) or (inputs(182));
    layer0_outputs(705) <= (inputs(138)) and not (inputs(216));
    layer0_outputs(706) <= (inputs(38)) and not (inputs(205));
    layer0_outputs(707) <= inputs(110);
    layer0_outputs(708) <= (inputs(171)) xor (inputs(189));
    layer0_outputs(709) <= not((inputs(150)) xor (inputs(221)));
    layer0_outputs(710) <= inputs(229);
    layer0_outputs(711) <= not(inputs(27));
    layer0_outputs(712) <= not((inputs(236)) xor (inputs(44)));
    layer0_outputs(713) <= (inputs(168)) and not (inputs(225));
    layer0_outputs(714) <= (inputs(46)) or (inputs(95));
    layer0_outputs(715) <= not((inputs(40)) xor (inputs(43)));
    layer0_outputs(716) <= not((inputs(67)) or (inputs(188)));
    layer0_outputs(717) <= not((inputs(75)) xor (inputs(28)));
    layer0_outputs(718) <= inputs(119);
    layer0_outputs(719) <= (inputs(101)) and not (inputs(220));
    layer0_outputs(720) <= (inputs(235)) or (inputs(127));
    layer0_outputs(721) <= not(inputs(166)) or (inputs(1));
    layer0_outputs(722) <= inputs(87);
    layer0_outputs(723) <= not(inputs(163)) or (inputs(18));
    layer0_outputs(724) <= (inputs(196)) or (inputs(173));
    layer0_outputs(725) <= inputs(149);
    layer0_outputs(726) <= not(inputs(208)) or (inputs(162));
    layer0_outputs(727) <= not(inputs(62));
    layer0_outputs(728) <= (inputs(75)) xor (inputs(248));
    layer0_outputs(729) <= not(inputs(143)) or (inputs(123));
    layer0_outputs(730) <= (inputs(28)) or (inputs(108));
    layer0_outputs(731) <= (inputs(53)) xor (inputs(32));
    layer0_outputs(732) <= not((inputs(32)) or (inputs(248)));
    layer0_outputs(733) <= not(inputs(244));
    layer0_outputs(734) <= not((inputs(167)) and (inputs(75)));
    layer0_outputs(735) <= inputs(245);
    layer0_outputs(736) <= not((inputs(20)) or (inputs(18)));
    layer0_outputs(737) <= (inputs(76)) xor (inputs(6));
    layer0_outputs(738) <= not((inputs(44)) or (inputs(148)));
    layer0_outputs(739) <= not((inputs(54)) xor (inputs(0)));
    layer0_outputs(740) <= not((inputs(2)) xor (inputs(108)));
    layer0_outputs(741) <= (inputs(3)) or (inputs(192));
    layer0_outputs(742) <= (inputs(65)) xor (inputs(132));
    layer0_outputs(743) <= inputs(186);
    layer0_outputs(744) <= not(inputs(110));
    layer0_outputs(745) <= inputs(52);
    layer0_outputs(746) <= '0';
    layer0_outputs(747) <= inputs(108);
    layer0_outputs(748) <= (inputs(61)) or (inputs(166));
    layer0_outputs(749) <= inputs(70);
    layer0_outputs(750) <= not((inputs(185)) and (inputs(50)));
    layer0_outputs(751) <= (inputs(19)) or (inputs(178));
    layer0_outputs(752) <= (inputs(60)) and (inputs(100));
    layer0_outputs(753) <= inputs(32);
    layer0_outputs(754) <= (inputs(93)) and not (inputs(118));
    layer0_outputs(755) <= (inputs(181)) xor (inputs(30));
    layer0_outputs(756) <= not(inputs(135)) or (inputs(107));
    layer0_outputs(757) <= not(inputs(204));
    layer0_outputs(758) <= not(inputs(195)) or (inputs(51));
    layer0_outputs(759) <= (inputs(44)) and (inputs(66));
    layer0_outputs(760) <= not((inputs(204)) xor (inputs(21)));
    layer0_outputs(761) <= inputs(246);
    layer0_outputs(762) <= not(inputs(175));
    layer0_outputs(763) <= (inputs(252)) or (inputs(230));
    layer0_outputs(764) <= (inputs(199)) and not (inputs(66));
    layer0_outputs(765) <= inputs(10);
    layer0_outputs(766) <= not(inputs(143));
    layer0_outputs(767) <= inputs(41);
    layer0_outputs(768) <= (inputs(225)) xor (inputs(74));
    layer0_outputs(769) <= not((inputs(157)) or (inputs(128)));
    layer0_outputs(770) <= (inputs(197)) or (inputs(61));
    layer0_outputs(771) <= inputs(71);
    layer0_outputs(772) <= (inputs(227)) or (inputs(202));
    layer0_outputs(773) <= (inputs(25)) and not (inputs(172));
    layer0_outputs(774) <= not(inputs(121)) or (inputs(64));
    layer0_outputs(775) <= not(inputs(134));
    layer0_outputs(776) <= not(inputs(40)) or (inputs(129));
    layer0_outputs(777) <= not(inputs(100));
    layer0_outputs(778) <= inputs(69);
    layer0_outputs(779) <= not((inputs(177)) and (inputs(240)));
    layer0_outputs(780) <= not(inputs(86));
    layer0_outputs(781) <= '0';
    layer0_outputs(782) <= (inputs(50)) xor (inputs(54));
    layer0_outputs(783) <= not(inputs(229)) or (inputs(66));
    layer0_outputs(784) <= (inputs(120)) or (inputs(150));
    layer0_outputs(785) <= inputs(249);
    layer0_outputs(786) <= not(inputs(231)) or (inputs(67));
    layer0_outputs(787) <= not((inputs(140)) xor (inputs(206)));
    layer0_outputs(788) <= not(inputs(105));
    layer0_outputs(789) <= (inputs(76)) and not (inputs(195));
    layer0_outputs(790) <= (inputs(149)) xor (inputs(197));
    layer0_outputs(791) <= (inputs(117)) xor (inputs(71));
    layer0_outputs(792) <= inputs(60);
    layer0_outputs(793) <= not(inputs(36));
    layer0_outputs(794) <= (inputs(186)) and (inputs(134));
    layer0_outputs(795) <= not(inputs(248));
    layer0_outputs(796) <= not(inputs(86));
    layer0_outputs(797) <= not(inputs(252));
    layer0_outputs(798) <= not((inputs(108)) and (inputs(231)));
    layer0_outputs(799) <= not((inputs(98)) or (inputs(22)));
    layer0_outputs(800) <= inputs(76);
    layer0_outputs(801) <= not(inputs(15));
    layer0_outputs(802) <= (inputs(191)) or (inputs(141));
    layer0_outputs(803) <= not((inputs(98)) or (inputs(112)));
    layer0_outputs(804) <= '0';
    layer0_outputs(805) <= not((inputs(167)) xor (inputs(70)));
    layer0_outputs(806) <= '1';
    layer0_outputs(807) <= not(inputs(155)) or (inputs(96));
    layer0_outputs(808) <= not(inputs(230)) or (inputs(88));
    layer0_outputs(809) <= not(inputs(189)) or (inputs(51));
    layer0_outputs(810) <= inputs(114);
    layer0_outputs(811) <= not((inputs(126)) xor (inputs(9)));
    layer0_outputs(812) <= not(inputs(73)) or (inputs(84));
    layer0_outputs(813) <= (inputs(173)) or (inputs(228));
    layer0_outputs(814) <= not((inputs(238)) xor (inputs(156)));
    layer0_outputs(815) <= not(inputs(158));
    layer0_outputs(816) <= not((inputs(17)) or (inputs(238)));
    layer0_outputs(817) <= inputs(85);
    layer0_outputs(818) <= (inputs(132)) and not (inputs(242));
    layer0_outputs(819) <= not(inputs(166));
    layer0_outputs(820) <= not((inputs(12)) xor (inputs(42)));
    layer0_outputs(821) <= not((inputs(11)) and (inputs(149)));
    layer0_outputs(822) <= (inputs(127)) and not (inputs(118));
    layer0_outputs(823) <= not((inputs(173)) xor (inputs(120)));
    layer0_outputs(824) <= not(inputs(68));
    layer0_outputs(825) <= (inputs(41)) or (inputs(27));
    layer0_outputs(826) <= not((inputs(222)) xor (inputs(125)));
    layer0_outputs(827) <= inputs(219);
    layer0_outputs(828) <= (inputs(223)) and not (inputs(141));
    layer0_outputs(829) <= inputs(111);
    layer0_outputs(830) <= not(inputs(22));
    layer0_outputs(831) <= (inputs(195)) and not (inputs(96));
    layer0_outputs(832) <= not((inputs(194)) xor (inputs(240)));
    layer0_outputs(833) <= not((inputs(219)) and (inputs(90)));
    layer0_outputs(834) <= not(inputs(231));
    layer0_outputs(835) <= '0';
    layer0_outputs(836) <= not((inputs(245)) xor (inputs(159)));
    layer0_outputs(837) <= inputs(178);
    layer0_outputs(838) <= inputs(233);
    layer0_outputs(839) <= not(inputs(55));
    layer0_outputs(840) <= not(inputs(146));
    layer0_outputs(841) <= (inputs(222)) xor (inputs(3));
    layer0_outputs(842) <= (inputs(152)) and not (inputs(11));
    layer0_outputs(843) <= not(inputs(110));
    layer0_outputs(844) <= not((inputs(80)) or (inputs(169)));
    layer0_outputs(845) <= (inputs(122)) and (inputs(189));
    layer0_outputs(846) <= not(inputs(124)) or (inputs(17));
    layer0_outputs(847) <= (inputs(91)) xor (inputs(141));
    layer0_outputs(848) <= (inputs(26)) xor (inputs(76));
    layer0_outputs(849) <= not((inputs(246)) xor (inputs(5)));
    layer0_outputs(850) <= not(inputs(94));
    layer0_outputs(851) <= not((inputs(81)) xor (inputs(172)));
    layer0_outputs(852) <= inputs(127);
    layer0_outputs(853) <= not((inputs(0)) or (inputs(221)));
    layer0_outputs(854) <= (inputs(85)) and not (inputs(32));
    layer0_outputs(855) <= not(inputs(33)) or (inputs(198));
    layer0_outputs(856) <= not(inputs(213));
    layer0_outputs(857) <= not(inputs(140)) or (inputs(167));
    layer0_outputs(858) <= not(inputs(196));
    layer0_outputs(859) <= (inputs(108)) and not (inputs(159));
    layer0_outputs(860) <= inputs(104);
    layer0_outputs(861) <= not(inputs(24));
    layer0_outputs(862) <= inputs(184);
    layer0_outputs(863) <= inputs(163);
    layer0_outputs(864) <= not(inputs(85)) or (inputs(238));
    layer0_outputs(865) <= (inputs(233)) or (inputs(161));
    layer0_outputs(866) <= not(inputs(82));
    layer0_outputs(867) <= not(inputs(28)) or (inputs(239));
    layer0_outputs(868) <= '0';
    layer0_outputs(869) <= (inputs(0)) and not (inputs(124));
    layer0_outputs(870) <= not(inputs(43)) or (inputs(224));
    layer0_outputs(871) <= inputs(219);
    layer0_outputs(872) <= (inputs(34)) or (inputs(36));
    layer0_outputs(873) <= (inputs(50)) and (inputs(4));
    layer0_outputs(874) <= inputs(78);
    layer0_outputs(875) <= not(inputs(199)) or (inputs(46));
    layer0_outputs(876) <= not((inputs(240)) xor (inputs(210)));
    layer0_outputs(877) <= not(inputs(163));
    layer0_outputs(878) <= (inputs(165)) and not (inputs(37));
    layer0_outputs(879) <= not(inputs(142));
    layer0_outputs(880) <= (inputs(196)) and not (inputs(236));
    layer0_outputs(881) <= not((inputs(34)) or (inputs(4)));
    layer0_outputs(882) <= (inputs(121)) xor (inputs(91));
    layer0_outputs(883) <= not(inputs(124));
    layer0_outputs(884) <= (inputs(162)) xor (inputs(160));
    layer0_outputs(885) <= (inputs(70)) and not (inputs(190));
    layer0_outputs(886) <= not((inputs(88)) or (inputs(59)));
    layer0_outputs(887) <= (inputs(178)) and not (inputs(153));
    layer0_outputs(888) <= not(inputs(122));
    layer0_outputs(889) <= inputs(61);
    layer0_outputs(890) <= (inputs(162)) and not (inputs(62));
    layer0_outputs(891) <= not((inputs(4)) xor (inputs(182)));
    layer0_outputs(892) <= (inputs(12)) or (inputs(74));
    layer0_outputs(893) <= (inputs(116)) and (inputs(26));
    layer0_outputs(894) <= not((inputs(47)) or (inputs(252)));
    layer0_outputs(895) <= not(inputs(143)) or (inputs(48));
    layer0_outputs(896) <= inputs(211);
    layer0_outputs(897) <= not(inputs(36)) or (inputs(251));
    layer0_outputs(898) <= not((inputs(19)) xor (inputs(77)));
    layer0_outputs(899) <= (inputs(234)) xor (inputs(196));
    layer0_outputs(900) <= (inputs(228)) xor (inputs(193));
    layer0_outputs(901) <= (inputs(227)) xor (inputs(7));
    layer0_outputs(902) <= (inputs(36)) and not (inputs(237));
    layer0_outputs(903) <= (inputs(100)) xor (inputs(132));
    layer0_outputs(904) <= not(inputs(110));
    layer0_outputs(905) <= (inputs(208)) or (inputs(15));
    layer0_outputs(906) <= (inputs(125)) or (inputs(17));
    layer0_outputs(907) <= not((inputs(79)) xor (inputs(9)));
    layer0_outputs(908) <= (inputs(175)) or (inputs(126));
    layer0_outputs(909) <= (inputs(85)) or (inputs(13));
    layer0_outputs(910) <= not((inputs(226)) xor (inputs(20)));
    layer0_outputs(911) <= (inputs(15)) or (inputs(57));
    layer0_outputs(912) <= (inputs(107)) and not (inputs(47));
    layer0_outputs(913) <= (inputs(55)) and not (inputs(35));
    layer0_outputs(914) <= inputs(223);
    layer0_outputs(915) <= not(inputs(138));
    layer0_outputs(916) <= not(inputs(7)) or (inputs(16));
    layer0_outputs(917) <= (inputs(181)) and not (inputs(52));
    layer0_outputs(918) <= not((inputs(169)) and (inputs(204)));
    layer0_outputs(919) <= (inputs(109)) and not (inputs(216));
    layer0_outputs(920) <= not(inputs(38));
    layer0_outputs(921) <= (inputs(25)) or (inputs(35));
    layer0_outputs(922) <= (inputs(125)) and not (inputs(127));
    layer0_outputs(923) <= not((inputs(29)) xor (inputs(155)));
    layer0_outputs(924) <= (inputs(247)) and (inputs(20));
    layer0_outputs(925) <= not(inputs(29));
    layer0_outputs(926) <= not((inputs(244)) or (inputs(27)));
    layer0_outputs(927) <= not(inputs(122)) or (inputs(242));
    layer0_outputs(928) <= not((inputs(96)) or (inputs(134)));
    layer0_outputs(929) <= (inputs(123)) and not (inputs(235));
    layer0_outputs(930) <= inputs(128);
    layer0_outputs(931) <= inputs(113);
    layer0_outputs(932) <= inputs(16);
    layer0_outputs(933) <= (inputs(78)) xor (inputs(252));
    layer0_outputs(934) <= not((inputs(228)) xor (inputs(73)));
    layer0_outputs(935) <= not(inputs(138)) or (inputs(73));
    layer0_outputs(936) <= inputs(90);
    layer0_outputs(937) <= (inputs(34)) or (inputs(168));
    layer0_outputs(938) <= not(inputs(199));
    layer0_outputs(939) <= (inputs(90)) or (inputs(139));
    layer0_outputs(940) <= not(inputs(83));
    layer0_outputs(941) <= (inputs(5)) or (inputs(29));
    layer0_outputs(942) <= (inputs(53)) and (inputs(92));
    layer0_outputs(943) <= not(inputs(176));
    layer0_outputs(944) <= (inputs(146)) or (inputs(123));
    layer0_outputs(945) <= inputs(138);
    layer0_outputs(946) <= (inputs(147)) and not (inputs(0));
    layer0_outputs(947) <= not(inputs(206));
    layer0_outputs(948) <= not((inputs(178)) xor (inputs(118)));
    layer0_outputs(949) <= (inputs(50)) and not (inputs(177));
    layer0_outputs(950) <= (inputs(219)) xor (inputs(85));
    layer0_outputs(951) <= not(inputs(152));
    layer0_outputs(952) <= not((inputs(221)) or (inputs(202)));
    layer0_outputs(953) <= not(inputs(23));
    layer0_outputs(954) <= (inputs(93)) and not (inputs(225));
    layer0_outputs(955) <= (inputs(91)) xor (inputs(42));
    layer0_outputs(956) <= not((inputs(170)) xor (inputs(242)));
    layer0_outputs(957) <= (inputs(101)) and not (inputs(206));
    layer0_outputs(958) <= (inputs(247)) or (inputs(97));
    layer0_outputs(959) <= not(inputs(230));
    layer0_outputs(960) <= not((inputs(84)) xor (inputs(219)));
    layer0_outputs(961) <= (inputs(174)) xor (inputs(185));
    layer0_outputs(962) <= not(inputs(227)) or (inputs(82));
    layer0_outputs(963) <= inputs(241);
    layer0_outputs(964) <= '0';
    layer0_outputs(965) <= (inputs(146)) xor (inputs(117));
    layer0_outputs(966) <= not((inputs(253)) or (inputs(123)));
    layer0_outputs(967) <= (inputs(88)) and not (inputs(50));
    layer0_outputs(968) <= inputs(45);
    layer0_outputs(969) <= not(inputs(97));
    layer0_outputs(970) <= not(inputs(119)) or (inputs(144));
    layer0_outputs(971) <= not((inputs(63)) xor (inputs(12)));
    layer0_outputs(972) <= not(inputs(70));
    layer0_outputs(973) <= not(inputs(13));
    layer0_outputs(974) <= (inputs(78)) and not (inputs(165));
    layer0_outputs(975) <= not((inputs(54)) xor (inputs(12)));
    layer0_outputs(976) <= not(inputs(171)) or (inputs(49));
    layer0_outputs(977) <= (inputs(51)) or (inputs(10));
    layer0_outputs(978) <= inputs(109);
    layer0_outputs(979) <= (inputs(164)) and not (inputs(204));
    layer0_outputs(980) <= inputs(195);
    layer0_outputs(981) <= not(inputs(112));
    layer0_outputs(982) <= not((inputs(71)) xor (inputs(51)));
    layer0_outputs(983) <= inputs(39);
    layer0_outputs(984) <= inputs(226);
    layer0_outputs(985) <= not((inputs(121)) or (inputs(138)));
    layer0_outputs(986) <= not(inputs(195));
    layer0_outputs(987) <= not(inputs(218)) or (inputs(208));
    layer0_outputs(988) <= not(inputs(235)) or (inputs(174));
    layer0_outputs(989) <= (inputs(51)) xor (inputs(245));
    layer0_outputs(990) <= not(inputs(64));
    layer0_outputs(991) <= (inputs(228)) and (inputs(249));
    layer0_outputs(992) <= not((inputs(185)) or (inputs(125)));
    layer0_outputs(993) <= not((inputs(176)) xor (inputs(202)));
    layer0_outputs(994) <= not(inputs(247));
    layer0_outputs(995) <= not(inputs(200));
    layer0_outputs(996) <= not(inputs(67));
    layer0_outputs(997) <= (inputs(10)) or (inputs(81));
    layer0_outputs(998) <= not(inputs(183));
    layer0_outputs(999) <= not(inputs(128)) or (inputs(99));
    layer0_outputs(1000) <= not(inputs(132));
    layer0_outputs(1001) <= not((inputs(197)) and (inputs(201)));
    layer0_outputs(1002) <= (inputs(230)) xor (inputs(252));
    layer0_outputs(1003) <= (inputs(60)) and not (inputs(17));
    layer0_outputs(1004) <= not(inputs(200)) or (inputs(184));
    layer0_outputs(1005) <= not(inputs(50)) or (inputs(112));
    layer0_outputs(1006) <= (inputs(241)) and (inputs(79));
    layer0_outputs(1007) <= not(inputs(102));
    layer0_outputs(1008) <= (inputs(125)) xor (inputs(152));
    layer0_outputs(1009) <= inputs(124);
    layer0_outputs(1010) <= not((inputs(190)) or (inputs(208)));
    layer0_outputs(1011) <= not((inputs(152)) or (inputs(56)));
    layer0_outputs(1012) <= not(inputs(212));
    layer0_outputs(1013) <= not(inputs(205));
    layer0_outputs(1014) <= inputs(21);
    layer0_outputs(1015) <= not(inputs(210));
    layer0_outputs(1016) <= not((inputs(34)) xor (inputs(70)));
    layer0_outputs(1017) <= '1';
    layer0_outputs(1018) <= not(inputs(84)) or (inputs(246));
    layer0_outputs(1019) <= not(inputs(118)) or (inputs(163));
    layer0_outputs(1020) <= not(inputs(43));
    layer0_outputs(1021) <= '1';
    layer0_outputs(1022) <= (inputs(21)) or (inputs(191));
    layer0_outputs(1023) <= (inputs(172)) xor (inputs(19));
    layer0_outputs(1024) <= (inputs(25)) and not (inputs(36));
    layer0_outputs(1025) <= (inputs(56)) and not (inputs(153));
    layer0_outputs(1026) <= not(inputs(55));
    layer0_outputs(1027) <= (inputs(45)) xor (inputs(147));
    layer0_outputs(1028) <= not((inputs(58)) or (inputs(63)));
    layer0_outputs(1029) <= not(inputs(243));
    layer0_outputs(1030) <= not((inputs(84)) or (inputs(177)));
    layer0_outputs(1031) <= not((inputs(4)) xor (inputs(110)));
    layer0_outputs(1032) <= not(inputs(152)) or (inputs(251));
    layer0_outputs(1033) <= inputs(72);
    layer0_outputs(1034) <= inputs(103);
    layer0_outputs(1035) <= not(inputs(159));
    layer0_outputs(1036) <= (inputs(168)) xor (inputs(136));
    layer0_outputs(1037) <= (inputs(177)) xor (inputs(218));
    layer0_outputs(1038) <= (inputs(245)) and not (inputs(38));
    layer0_outputs(1039) <= not(inputs(8));
    layer0_outputs(1040) <= not(inputs(87));
    layer0_outputs(1041) <= inputs(128);
    layer0_outputs(1042) <= not(inputs(227)) or (inputs(51));
    layer0_outputs(1043) <= not((inputs(52)) xor (inputs(53)));
    layer0_outputs(1044) <= inputs(230);
    layer0_outputs(1045) <= not((inputs(13)) xor (inputs(200)));
    layer0_outputs(1046) <= not(inputs(109));
    layer0_outputs(1047) <= not(inputs(183));
    layer0_outputs(1048) <= (inputs(6)) xor (inputs(142));
    layer0_outputs(1049) <= inputs(168);
    layer0_outputs(1050) <= not(inputs(129)) or (inputs(254));
    layer0_outputs(1051) <= not((inputs(54)) and (inputs(221)));
    layer0_outputs(1052) <= (inputs(214)) and not (inputs(128));
    layer0_outputs(1053) <= not(inputs(129));
    layer0_outputs(1054) <= (inputs(17)) and not (inputs(251));
    layer0_outputs(1055) <= (inputs(132)) and not (inputs(144));
    layer0_outputs(1056) <= not(inputs(146));
    layer0_outputs(1057) <= not(inputs(120)) or (inputs(154));
    layer0_outputs(1058) <= not(inputs(113));
    layer0_outputs(1059) <= not(inputs(111));
    layer0_outputs(1060) <= not((inputs(79)) xor (inputs(180)));
    layer0_outputs(1061) <= inputs(37);
    layer0_outputs(1062) <= not(inputs(133)) or (inputs(123));
    layer0_outputs(1063) <= not(inputs(37)) or (inputs(239));
    layer0_outputs(1064) <= (inputs(47)) or (inputs(13));
    layer0_outputs(1065) <= (inputs(240)) xor (inputs(59));
    layer0_outputs(1066) <= '1';
    layer0_outputs(1067) <= (inputs(96)) and (inputs(224));
    layer0_outputs(1068) <= inputs(74);
    layer0_outputs(1069) <= not(inputs(37)) or (inputs(209));
    layer0_outputs(1070) <= not((inputs(219)) xor (inputs(249)));
    layer0_outputs(1071) <= (inputs(162)) and not (inputs(128));
    layer0_outputs(1072) <= (inputs(147)) or (inputs(1));
    layer0_outputs(1073) <= (inputs(181)) and not (inputs(33));
    layer0_outputs(1074) <= not((inputs(62)) or (inputs(214)));
    layer0_outputs(1075) <= not((inputs(240)) xor (inputs(211)));
    layer0_outputs(1076) <= inputs(39);
    layer0_outputs(1077) <= (inputs(33)) or (inputs(34));
    layer0_outputs(1078) <= (inputs(126)) or (inputs(197));
    layer0_outputs(1079) <= not(inputs(106));
    layer0_outputs(1080) <= not((inputs(9)) xor (inputs(237)));
    layer0_outputs(1081) <= not((inputs(143)) xor (inputs(22)));
    layer0_outputs(1082) <= not((inputs(23)) xor (inputs(158)));
    layer0_outputs(1083) <= (inputs(185)) or (inputs(192));
    layer0_outputs(1084) <= inputs(75);
    layer0_outputs(1085) <= not((inputs(217)) or (inputs(18)));
    layer0_outputs(1086) <= not(inputs(121));
    layer0_outputs(1087) <= not(inputs(115)) or (inputs(2));
    layer0_outputs(1088) <= (inputs(251)) xor (inputs(222));
    layer0_outputs(1089) <= '1';
    layer0_outputs(1090) <= (inputs(81)) xor (inputs(45));
    layer0_outputs(1091) <= (inputs(215)) xor (inputs(45));
    layer0_outputs(1092) <= inputs(84);
    layer0_outputs(1093) <= (inputs(91)) or (inputs(143));
    layer0_outputs(1094) <= inputs(4);
    layer0_outputs(1095) <= inputs(172);
    layer0_outputs(1096) <= (inputs(16)) and not (inputs(236));
    layer0_outputs(1097) <= not(inputs(157)) or (inputs(127));
    layer0_outputs(1098) <= not(inputs(179));
    layer0_outputs(1099) <= not((inputs(127)) xor (inputs(156)));
    layer0_outputs(1100) <= (inputs(31)) and not (inputs(10));
    layer0_outputs(1101) <= '1';
    layer0_outputs(1102) <= not(inputs(144)) or (inputs(115));
    layer0_outputs(1103) <= not(inputs(139)) or (inputs(207));
    layer0_outputs(1104) <= not((inputs(90)) or (inputs(222)));
    layer0_outputs(1105) <= (inputs(35)) or (inputs(23));
    layer0_outputs(1106) <= (inputs(5)) and not (inputs(51));
    layer0_outputs(1107) <= not((inputs(188)) or (inputs(125)));
    layer0_outputs(1108) <= not((inputs(52)) xor (inputs(251)));
    layer0_outputs(1109) <= not(inputs(68)) or (inputs(175));
    layer0_outputs(1110) <= (inputs(136)) xor (inputs(178));
    layer0_outputs(1111) <= (inputs(0)) and not (inputs(139));
    layer0_outputs(1112) <= not(inputs(214)) or (inputs(141));
    layer0_outputs(1113) <= not((inputs(224)) or (inputs(1)));
    layer0_outputs(1114) <= (inputs(96)) and not (inputs(160));
    layer0_outputs(1115) <= inputs(47);
    layer0_outputs(1116) <= (inputs(58)) and (inputs(196));
    layer0_outputs(1117) <= not(inputs(10));
    layer0_outputs(1118) <= not((inputs(136)) or (inputs(249)));
    layer0_outputs(1119) <= '1';
    layer0_outputs(1120) <= inputs(188);
    layer0_outputs(1121) <= not((inputs(210)) or (inputs(57)));
    layer0_outputs(1122) <= (inputs(109)) xor (inputs(196));
    layer0_outputs(1123) <= inputs(213);
    layer0_outputs(1124) <= not(inputs(35)) or (inputs(98));
    layer0_outputs(1125) <= inputs(84);
    layer0_outputs(1126) <= not(inputs(71));
    layer0_outputs(1127) <= (inputs(186)) xor (inputs(157));
    layer0_outputs(1128) <= not(inputs(192));
    layer0_outputs(1129) <= (inputs(176)) xor (inputs(38));
    layer0_outputs(1130) <= not(inputs(161));
    layer0_outputs(1131) <= (inputs(133)) xor (inputs(184));
    layer0_outputs(1132) <= not(inputs(232)) or (inputs(115));
    layer0_outputs(1133) <= (inputs(205)) and not (inputs(48));
    layer0_outputs(1134) <= inputs(146);
    layer0_outputs(1135) <= '0';
    layer0_outputs(1136) <= not((inputs(225)) xor (inputs(234)));
    layer0_outputs(1137) <= not(inputs(81)) or (inputs(207));
    layer0_outputs(1138) <= not(inputs(83)) or (inputs(232));
    layer0_outputs(1139) <= inputs(123);
    layer0_outputs(1140) <= not(inputs(158));
    layer0_outputs(1141) <= (inputs(238)) or (inputs(142));
    layer0_outputs(1142) <= not((inputs(40)) xor (inputs(63)));
    layer0_outputs(1143) <= (inputs(221)) and not (inputs(239));
    layer0_outputs(1144) <= inputs(220);
    layer0_outputs(1145) <= (inputs(120)) and not (inputs(24));
    layer0_outputs(1146) <= (inputs(63)) or (inputs(29));
    layer0_outputs(1147) <= not(inputs(228));
    layer0_outputs(1148) <= inputs(93);
    layer0_outputs(1149) <= inputs(43);
    layer0_outputs(1150) <= (inputs(51)) xor (inputs(35));
    layer0_outputs(1151) <= not((inputs(1)) or (inputs(41)));
    layer0_outputs(1152) <= not((inputs(9)) xor (inputs(117)));
    layer0_outputs(1153) <= (inputs(220)) or (inputs(79));
    layer0_outputs(1154) <= not((inputs(184)) or (inputs(235)));
    layer0_outputs(1155) <= inputs(25);
    layer0_outputs(1156) <= not(inputs(247)) or (inputs(89));
    layer0_outputs(1157) <= inputs(84);
    layer0_outputs(1158) <= (inputs(33)) and not (inputs(13));
    layer0_outputs(1159) <= (inputs(30)) or (inputs(159));
    layer0_outputs(1160) <= not(inputs(142));
    layer0_outputs(1161) <= (inputs(204)) xor (inputs(173));
    layer0_outputs(1162) <= not(inputs(50));
    layer0_outputs(1163) <= (inputs(167)) or (inputs(133));
    layer0_outputs(1164) <= not(inputs(184)) or (inputs(126));
    layer0_outputs(1165) <= not((inputs(4)) or (inputs(174)));
    layer0_outputs(1166) <= not(inputs(75));
    layer0_outputs(1167) <= '1';
    layer0_outputs(1168) <= '1';
    layer0_outputs(1169) <= (inputs(238)) xor (inputs(61));
    layer0_outputs(1170) <= (inputs(254)) and (inputs(200));
    layer0_outputs(1171) <= not(inputs(212)) or (inputs(32));
    layer0_outputs(1172) <= not((inputs(64)) and (inputs(253)));
    layer0_outputs(1173) <= inputs(119);
    layer0_outputs(1174) <= (inputs(208)) and (inputs(240));
    layer0_outputs(1175) <= (inputs(247)) or (inputs(194));
    layer0_outputs(1176) <= not(inputs(113));
    layer0_outputs(1177) <= not(inputs(133));
    layer0_outputs(1178) <= not((inputs(22)) or (inputs(56)));
    layer0_outputs(1179) <= (inputs(186)) and not (inputs(207));
    layer0_outputs(1180) <= (inputs(49)) and not (inputs(158));
    layer0_outputs(1181) <= inputs(91);
    layer0_outputs(1182) <= (inputs(214)) and (inputs(160));
    layer0_outputs(1183) <= (inputs(23)) xor (inputs(223));
    layer0_outputs(1184) <= not((inputs(120)) xor (inputs(250)));
    layer0_outputs(1185) <= inputs(67);
    layer0_outputs(1186) <= (inputs(250)) xor (inputs(52));
    layer0_outputs(1187) <= (inputs(118)) or (inputs(108));
    layer0_outputs(1188) <= not((inputs(253)) or (inputs(117)));
    layer0_outputs(1189) <= '0';
    layer0_outputs(1190) <= (inputs(75)) or (inputs(67));
    layer0_outputs(1191) <= inputs(104);
    layer0_outputs(1192) <= inputs(231);
    layer0_outputs(1193) <= not(inputs(30)) or (inputs(236));
    layer0_outputs(1194) <= not((inputs(208)) or (inputs(226)));
    layer0_outputs(1195) <= (inputs(12)) and not (inputs(61));
    layer0_outputs(1196) <= not((inputs(81)) xor (inputs(68)));
    layer0_outputs(1197) <= (inputs(30)) or (inputs(2));
    layer0_outputs(1198) <= (inputs(233)) and not (inputs(198));
    layer0_outputs(1199) <= (inputs(14)) and not (inputs(184));
    layer0_outputs(1200) <= not((inputs(190)) or (inputs(143)));
    layer0_outputs(1201) <= not((inputs(242)) or (inputs(139)));
    layer0_outputs(1202) <= not((inputs(26)) xor (inputs(252)));
    layer0_outputs(1203) <= (inputs(135)) and not (inputs(41));
    layer0_outputs(1204) <= inputs(213);
    layer0_outputs(1205) <= not(inputs(100));
    layer0_outputs(1206) <= (inputs(222)) xor (inputs(5));
    layer0_outputs(1207) <= (inputs(108)) and not (inputs(235));
    layer0_outputs(1208) <= not(inputs(247)) or (inputs(12));
    layer0_outputs(1209) <= (inputs(134)) xor (inputs(189));
    layer0_outputs(1210) <= not((inputs(241)) or (inputs(199)));
    layer0_outputs(1211) <= (inputs(129)) or (inputs(197));
    layer0_outputs(1212) <= not((inputs(245)) or (inputs(87)));
    layer0_outputs(1213) <= (inputs(207)) xor (inputs(177));
    layer0_outputs(1214) <= not(inputs(188));
    layer0_outputs(1215) <= (inputs(191)) or (inputs(160));
    layer0_outputs(1216) <= not((inputs(185)) and (inputs(179)));
    layer0_outputs(1217) <= (inputs(237)) and (inputs(213));
    layer0_outputs(1218) <= not(inputs(19)) or (inputs(237));
    layer0_outputs(1219) <= not(inputs(193));
    layer0_outputs(1220) <= (inputs(70)) and not (inputs(21));
    layer0_outputs(1221) <= (inputs(37)) and (inputs(39));
    layer0_outputs(1222) <= (inputs(211)) and not (inputs(165));
    layer0_outputs(1223) <= not(inputs(77)) or (inputs(197));
    layer0_outputs(1224) <= '0';
    layer0_outputs(1225) <= not((inputs(236)) and (inputs(18)));
    layer0_outputs(1226) <= not((inputs(37)) or (inputs(20)));
    layer0_outputs(1227) <= (inputs(35)) or (inputs(4));
    layer0_outputs(1228) <= not(inputs(229)) or (inputs(62));
    layer0_outputs(1229) <= (inputs(200)) xor (inputs(165));
    layer0_outputs(1230) <= inputs(194);
    layer0_outputs(1231) <= (inputs(244)) xor (inputs(80));
    layer0_outputs(1232) <= '1';
    layer0_outputs(1233) <= not(inputs(0));
    layer0_outputs(1234) <= (inputs(83)) and not (inputs(160));
    layer0_outputs(1235) <= (inputs(70)) xor (inputs(7));
    layer0_outputs(1236) <= not(inputs(157));
    layer0_outputs(1237) <= (inputs(206)) or (inputs(190));
    layer0_outputs(1238) <= inputs(38);
    layer0_outputs(1239) <= inputs(58);
    layer0_outputs(1240) <= not((inputs(54)) or (inputs(218)));
    layer0_outputs(1241) <= not((inputs(70)) or (inputs(184)));
    layer0_outputs(1242) <= not((inputs(24)) or (inputs(38)));
    layer0_outputs(1243) <= not((inputs(73)) xor (inputs(71)));
    layer0_outputs(1244) <= (inputs(43)) xor (inputs(200));
    layer0_outputs(1245) <= not((inputs(180)) xor (inputs(173)));
    layer0_outputs(1246) <= not((inputs(255)) or (inputs(132)));
    layer0_outputs(1247) <= (inputs(73)) or (inputs(191));
    layer0_outputs(1248) <= (inputs(131)) or (inputs(237));
    layer0_outputs(1249) <= (inputs(170)) and not (inputs(192));
    layer0_outputs(1250) <= (inputs(82)) or (inputs(28));
    layer0_outputs(1251) <= (inputs(42)) and not (inputs(186));
    layer0_outputs(1252) <= not((inputs(116)) or (inputs(147)));
    layer0_outputs(1253) <= not(inputs(11));
    layer0_outputs(1254) <= (inputs(180)) and not (inputs(70));
    layer0_outputs(1255) <= inputs(175);
    layer0_outputs(1256) <= not((inputs(68)) or (inputs(129)));
    layer0_outputs(1257) <= (inputs(206)) xor (inputs(255));
    layer0_outputs(1258) <= (inputs(206)) xor (inputs(24));
    layer0_outputs(1259) <= inputs(234);
    layer0_outputs(1260) <= (inputs(172)) and not (inputs(222));
    layer0_outputs(1261) <= not((inputs(68)) xor (inputs(149)));
    layer0_outputs(1262) <= (inputs(67)) or (inputs(169));
    layer0_outputs(1263) <= (inputs(139)) and not (inputs(44));
    layer0_outputs(1264) <= not(inputs(141));
    layer0_outputs(1265) <= not(inputs(47));
    layer0_outputs(1266) <= not((inputs(131)) or (inputs(132)));
    layer0_outputs(1267) <= (inputs(35)) or (inputs(169));
    layer0_outputs(1268) <= not((inputs(113)) or (inputs(28)));
    layer0_outputs(1269) <= not(inputs(151));
    layer0_outputs(1270) <= inputs(23);
    layer0_outputs(1271) <= not(inputs(115)) or (inputs(93));
    layer0_outputs(1272) <= inputs(23);
    layer0_outputs(1273) <= not(inputs(71)) or (inputs(48));
    layer0_outputs(1274) <= inputs(239);
    layer0_outputs(1275) <= inputs(39);
    layer0_outputs(1276) <= inputs(117);
    layer0_outputs(1277) <= (inputs(153)) and not (inputs(30));
    layer0_outputs(1278) <= not((inputs(253)) xor (inputs(231)));
    layer0_outputs(1279) <= (inputs(45)) or (inputs(202));
    layer0_outputs(1280) <= not(inputs(79));
    layer0_outputs(1281) <= inputs(53);
    layer0_outputs(1282) <= not((inputs(47)) xor (inputs(59)));
    layer0_outputs(1283) <= not((inputs(153)) xor (inputs(134)));
    layer0_outputs(1284) <= not((inputs(132)) or (inputs(79)));
    layer0_outputs(1285) <= not((inputs(144)) or (inputs(143)));
    layer0_outputs(1286) <= inputs(129);
    layer0_outputs(1287) <= not(inputs(203));
    layer0_outputs(1288) <= inputs(8);
    layer0_outputs(1289) <= (inputs(212)) and not (inputs(120));
    layer0_outputs(1290) <= not((inputs(225)) or (inputs(253)));
    layer0_outputs(1291) <= not(inputs(221)) or (inputs(240));
    layer0_outputs(1292) <= inputs(132);
    layer0_outputs(1293) <= inputs(168);
    layer0_outputs(1294) <= not((inputs(139)) or (inputs(28)));
    layer0_outputs(1295) <= inputs(23);
    layer0_outputs(1296) <= not((inputs(203)) xor (inputs(187)));
    layer0_outputs(1297) <= not((inputs(19)) or (inputs(46)));
    layer0_outputs(1298) <= not(inputs(232));
    layer0_outputs(1299) <= inputs(42);
    layer0_outputs(1300) <= (inputs(150)) xor (inputs(251));
    layer0_outputs(1301) <= not((inputs(170)) and (inputs(184)));
    layer0_outputs(1302) <= '0';
    layer0_outputs(1303) <= (inputs(210)) or (inputs(240));
    layer0_outputs(1304) <= (inputs(212)) and not (inputs(197));
    layer0_outputs(1305) <= not(inputs(90));
    layer0_outputs(1306) <= not(inputs(215));
    layer0_outputs(1307) <= inputs(251);
    layer0_outputs(1308) <= not(inputs(199));
    layer0_outputs(1309) <= not((inputs(121)) or (inputs(19)));
    layer0_outputs(1310) <= inputs(146);
    layer0_outputs(1311) <= (inputs(143)) xor (inputs(116));
    layer0_outputs(1312) <= (inputs(103)) xor (inputs(138));
    layer0_outputs(1313) <= not(inputs(12));
    layer0_outputs(1314) <= (inputs(86)) and not (inputs(251));
    layer0_outputs(1315) <= inputs(228);
    layer0_outputs(1316) <= not(inputs(100));
    layer0_outputs(1317) <= not(inputs(111));
    layer0_outputs(1318) <= (inputs(204)) and not (inputs(145));
    layer0_outputs(1319) <= not((inputs(13)) or (inputs(84)));
    layer0_outputs(1320) <= (inputs(64)) or (inputs(49));
    layer0_outputs(1321) <= not((inputs(67)) or (inputs(255)));
    layer0_outputs(1322) <= '0';
    layer0_outputs(1323) <= not(inputs(206));
    layer0_outputs(1324) <= not(inputs(55)) or (inputs(230));
    layer0_outputs(1325) <= not(inputs(76));
    layer0_outputs(1326) <= (inputs(174)) xor (inputs(79));
    layer0_outputs(1327) <= (inputs(190)) and not (inputs(7));
    layer0_outputs(1328) <= not(inputs(19)) or (inputs(100));
    layer0_outputs(1329) <= not(inputs(236)) or (inputs(82));
    layer0_outputs(1330) <= not((inputs(144)) or (inputs(55)));
    layer0_outputs(1331) <= not(inputs(117)) or (inputs(21));
    layer0_outputs(1332) <= not(inputs(181)) or (inputs(61));
    layer0_outputs(1333) <= (inputs(44)) and not (inputs(183));
    layer0_outputs(1334) <= (inputs(104)) or (inputs(137));
    layer0_outputs(1335) <= not((inputs(159)) or (inputs(43)));
    layer0_outputs(1336) <= not(inputs(181)) or (inputs(15));
    layer0_outputs(1337) <= (inputs(40)) and not (inputs(156));
    layer0_outputs(1338) <= not(inputs(24)) or (inputs(161));
    layer0_outputs(1339) <= inputs(9);
    layer0_outputs(1340) <= not(inputs(167)) or (inputs(27));
    layer0_outputs(1341) <= not(inputs(35)) or (inputs(225));
    layer0_outputs(1342) <= not(inputs(177));
    layer0_outputs(1343) <= not(inputs(124));
    layer0_outputs(1344) <= (inputs(19)) or (inputs(41));
    layer0_outputs(1345) <= not(inputs(151));
    layer0_outputs(1346) <= inputs(190);
    layer0_outputs(1347) <= (inputs(227)) and not (inputs(255));
    layer0_outputs(1348) <= (inputs(179)) xor (inputs(105));
    layer0_outputs(1349) <= (inputs(230)) and (inputs(74));
    layer0_outputs(1350) <= inputs(50);
    layer0_outputs(1351) <= not(inputs(84));
    layer0_outputs(1352) <= not(inputs(151)) or (inputs(110));
    layer0_outputs(1353) <= '1';
    layer0_outputs(1354) <= not((inputs(217)) or (inputs(222)));
    layer0_outputs(1355) <= not((inputs(7)) xor (inputs(182)));
    layer0_outputs(1356) <= not(inputs(150)) or (inputs(208));
    layer0_outputs(1357) <= not(inputs(228)) or (inputs(69));
    layer0_outputs(1358) <= '1';
    layer0_outputs(1359) <= not(inputs(165));
    layer0_outputs(1360) <= not((inputs(89)) xor (inputs(148)));
    layer0_outputs(1361) <= inputs(72);
    layer0_outputs(1362) <= not(inputs(131));
    layer0_outputs(1363) <= not(inputs(14));
    layer0_outputs(1364) <= (inputs(234)) xor (inputs(160));
    layer0_outputs(1365) <= not((inputs(154)) and (inputs(9)));
    layer0_outputs(1366) <= (inputs(160)) xor (inputs(254));
    layer0_outputs(1367) <= not(inputs(209));
    layer0_outputs(1368) <= not(inputs(127));
    layer0_outputs(1369) <= (inputs(176)) xor (inputs(58));
    layer0_outputs(1370) <= not((inputs(202)) xor (inputs(178)));
    layer0_outputs(1371) <= (inputs(144)) or (inputs(45));
    layer0_outputs(1372) <= not((inputs(133)) xor (inputs(218)));
    layer0_outputs(1373) <= (inputs(190)) or (inputs(229));
    layer0_outputs(1374) <= not(inputs(170));
    layer0_outputs(1375) <= not(inputs(77)) or (inputs(96));
    layer0_outputs(1376) <= (inputs(123)) and not (inputs(204));
    layer0_outputs(1377) <= not((inputs(49)) or (inputs(162)));
    layer0_outputs(1378) <= not(inputs(134));
    layer0_outputs(1379) <= (inputs(158)) and not (inputs(51));
    layer0_outputs(1380) <= not(inputs(182)) or (inputs(62));
    layer0_outputs(1381) <= (inputs(226)) or (inputs(135));
    layer0_outputs(1382) <= not(inputs(229)) or (inputs(126));
    layer0_outputs(1383) <= inputs(179);
    layer0_outputs(1384) <= inputs(121);
    layer0_outputs(1385) <= not((inputs(3)) xor (inputs(195)));
    layer0_outputs(1386) <= not(inputs(252)) or (inputs(17));
    layer0_outputs(1387) <= not(inputs(99)) or (inputs(125));
    layer0_outputs(1388) <= not((inputs(228)) and (inputs(199)));
    layer0_outputs(1389) <= not((inputs(138)) and (inputs(233)));
    layer0_outputs(1390) <= (inputs(140)) and not (inputs(140));
    layer0_outputs(1391) <= not(inputs(121)) or (inputs(41));
    layer0_outputs(1392) <= (inputs(101)) xor (inputs(80));
    layer0_outputs(1393) <= not(inputs(248));
    layer0_outputs(1394) <= inputs(26);
    layer0_outputs(1395) <= not((inputs(23)) or (inputs(16)));
    layer0_outputs(1396) <= not(inputs(39)) or (inputs(181));
    layer0_outputs(1397) <= (inputs(212)) and (inputs(209));
    layer0_outputs(1398) <= (inputs(222)) or (inputs(126));
    layer0_outputs(1399) <= (inputs(11)) or (inputs(27));
    layer0_outputs(1400) <= not(inputs(103));
    layer0_outputs(1401) <= inputs(214);
    layer0_outputs(1402) <= inputs(126);
    layer0_outputs(1403) <= (inputs(26)) and (inputs(92));
    layer0_outputs(1404) <= not((inputs(197)) xor (inputs(250)));
    layer0_outputs(1405) <= not(inputs(95)) or (inputs(31));
    layer0_outputs(1406) <= not((inputs(104)) xor (inputs(224)));
    layer0_outputs(1407) <= not(inputs(200));
    layer0_outputs(1408) <= not(inputs(105));
    layer0_outputs(1409) <= (inputs(181)) or (inputs(97));
    layer0_outputs(1410) <= '0';
    layer0_outputs(1411) <= (inputs(57)) or (inputs(254));
    layer0_outputs(1412) <= not(inputs(185));
    layer0_outputs(1413) <= not((inputs(108)) xor (inputs(143)));
    layer0_outputs(1414) <= inputs(205);
    layer0_outputs(1415) <= not(inputs(187));
    layer0_outputs(1416) <= (inputs(9)) xor (inputs(109));
    layer0_outputs(1417) <= not(inputs(89)) or (inputs(128));
    layer0_outputs(1418) <= inputs(25);
    layer0_outputs(1419) <= (inputs(233)) xor (inputs(93));
    layer0_outputs(1420) <= (inputs(188)) and not (inputs(30));
    layer0_outputs(1421) <= not(inputs(140)) or (inputs(66));
    layer0_outputs(1422) <= not(inputs(103));
    layer0_outputs(1423) <= (inputs(12)) xor (inputs(177));
    layer0_outputs(1424) <= inputs(213);
    layer0_outputs(1425) <= not((inputs(143)) or (inputs(21)));
    layer0_outputs(1426) <= not((inputs(25)) xor (inputs(111)));
    layer0_outputs(1427) <= (inputs(125)) or (inputs(117));
    layer0_outputs(1428) <= (inputs(31)) xor (inputs(246));
    layer0_outputs(1429) <= not(inputs(44)) or (inputs(129));
    layer0_outputs(1430) <= not((inputs(149)) or (inputs(177)));
    layer0_outputs(1431) <= not((inputs(240)) xor (inputs(45)));
    layer0_outputs(1432) <= not(inputs(107));
    layer0_outputs(1433) <= (inputs(59)) or (inputs(166));
    layer0_outputs(1434) <= not((inputs(112)) or (inputs(172)));
    layer0_outputs(1435) <= (inputs(116)) and not (inputs(186));
    layer0_outputs(1436) <= (inputs(225)) and (inputs(22));
    layer0_outputs(1437) <= (inputs(18)) and not (inputs(34));
    layer0_outputs(1438) <= (inputs(104)) or (inputs(49));
    layer0_outputs(1439) <= not(inputs(96));
    layer0_outputs(1440) <= not(inputs(124)) or (inputs(129));
    layer0_outputs(1441) <= inputs(220);
    layer0_outputs(1442) <= not((inputs(52)) xor (inputs(101)));
    layer0_outputs(1443) <= not(inputs(168));
    layer0_outputs(1444) <= not(inputs(123));
    layer0_outputs(1445) <= (inputs(195)) or (inputs(211));
    layer0_outputs(1446) <= not((inputs(123)) and (inputs(224)));
    layer0_outputs(1447) <= (inputs(204)) and not (inputs(114));
    layer0_outputs(1448) <= inputs(124);
    layer0_outputs(1449) <= (inputs(201)) or (inputs(214));
    layer0_outputs(1450) <= not(inputs(107)) or (inputs(40));
    layer0_outputs(1451) <= (inputs(195)) or (inputs(171));
    layer0_outputs(1452) <= not((inputs(180)) or (inputs(176)));
    layer0_outputs(1453) <= not(inputs(52)) or (inputs(208));
    layer0_outputs(1454) <= (inputs(73)) and not (inputs(210));
    layer0_outputs(1455) <= (inputs(25)) or (inputs(144));
    layer0_outputs(1456) <= (inputs(41)) and (inputs(73));
    layer0_outputs(1457) <= not(inputs(177)) or (inputs(160));
    layer0_outputs(1458) <= (inputs(242)) xor (inputs(153));
    layer0_outputs(1459) <= inputs(49);
    layer0_outputs(1460) <= (inputs(114)) and (inputs(12));
    layer0_outputs(1461) <= not(inputs(199)) or (inputs(93));
    layer0_outputs(1462) <= (inputs(5)) or (inputs(121));
    layer0_outputs(1463) <= (inputs(247)) and not (inputs(2));
    layer0_outputs(1464) <= inputs(233);
    layer0_outputs(1465) <= not(inputs(10));
    layer0_outputs(1466) <= not(inputs(58)) or (inputs(27));
    layer0_outputs(1467) <= (inputs(203)) or (inputs(113));
    layer0_outputs(1468) <= (inputs(65)) and (inputs(247));
    layer0_outputs(1469) <= not((inputs(144)) or (inputs(25)));
    layer0_outputs(1470) <= '1';
    layer0_outputs(1471) <= inputs(99);
    layer0_outputs(1472) <= (inputs(194)) or (inputs(190));
    layer0_outputs(1473) <= not((inputs(95)) xor (inputs(17)));
    layer0_outputs(1474) <= (inputs(42)) or (inputs(174));
    layer0_outputs(1475) <= not((inputs(191)) or (inputs(121)));
    layer0_outputs(1476) <= not(inputs(144)) or (inputs(149));
    layer0_outputs(1477) <= (inputs(2)) and not (inputs(47));
    layer0_outputs(1478) <= not((inputs(210)) xor (inputs(99)));
    layer0_outputs(1479) <= (inputs(26)) and not (inputs(143));
    layer0_outputs(1480) <= inputs(187);
    layer0_outputs(1481) <= (inputs(243)) and (inputs(128));
    layer0_outputs(1482) <= not((inputs(166)) or (inputs(252)));
    layer0_outputs(1483) <= not((inputs(44)) or (inputs(128)));
    layer0_outputs(1484) <= inputs(219);
    layer0_outputs(1485) <= (inputs(249)) or (inputs(112));
    layer0_outputs(1486) <= (inputs(133)) and not (inputs(230));
    layer0_outputs(1487) <= not(inputs(233));
    layer0_outputs(1488) <= (inputs(6)) and not (inputs(35));
    layer0_outputs(1489) <= not(inputs(197)) or (inputs(45));
    layer0_outputs(1490) <= (inputs(231)) xor (inputs(210));
    layer0_outputs(1491) <= not(inputs(118)) or (inputs(59));
    layer0_outputs(1492) <= (inputs(115)) xor (inputs(102));
    layer0_outputs(1493) <= (inputs(182)) and not (inputs(132));
    layer0_outputs(1494) <= (inputs(48)) or (inputs(135));
    layer0_outputs(1495) <= not(inputs(64));
    layer0_outputs(1496) <= not((inputs(150)) xor (inputs(69)));
    layer0_outputs(1497) <= '0';
    layer0_outputs(1498) <= not((inputs(72)) xor (inputs(244)));
    layer0_outputs(1499) <= not(inputs(77));
    layer0_outputs(1500) <= not(inputs(135));
    layer0_outputs(1501) <= inputs(75);
    layer0_outputs(1502) <= (inputs(56)) or (inputs(12));
    layer0_outputs(1503) <= not(inputs(19));
    layer0_outputs(1504) <= not(inputs(117));
    layer0_outputs(1505) <= (inputs(21)) or (inputs(141));
    layer0_outputs(1506) <= not(inputs(201));
    layer0_outputs(1507) <= inputs(228);
    layer0_outputs(1508) <= not(inputs(25)) or (inputs(248));
    layer0_outputs(1509) <= (inputs(234)) and (inputs(229));
    layer0_outputs(1510) <= '0';
    layer0_outputs(1511) <= (inputs(185)) and not (inputs(242));
    layer0_outputs(1512) <= not(inputs(169)) or (inputs(65));
    layer0_outputs(1513) <= (inputs(175)) or (inputs(159));
    layer0_outputs(1514) <= not(inputs(172)) or (inputs(19));
    layer0_outputs(1515) <= not(inputs(198)) or (inputs(140));
    layer0_outputs(1516) <= not((inputs(85)) or (inputs(19)));
    layer0_outputs(1517) <= not(inputs(21));
    layer0_outputs(1518) <= not((inputs(61)) or (inputs(228)));
    layer0_outputs(1519) <= inputs(171);
    layer0_outputs(1520) <= not((inputs(89)) or (inputs(238)));
    layer0_outputs(1521) <= (inputs(75)) and not (inputs(146));
    layer0_outputs(1522) <= not((inputs(141)) xor (inputs(244)));
    layer0_outputs(1523) <= not((inputs(172)) xor (inputs(39)));
    layer0_outputs(1524) <= not((inputs(149)) or (inputs(162)));
    layer0_outputs(1525) <= inputs(134);
    layer0_outputs(1526) <= not((inputs(2)) xor (inputs(153)));
    layer0_outputs(1527) <= (inputs(145)) xor (inputs(22));
    layer0_outputs(1528) <= not((inputs(76)) or (inputs(24)));
    layer0_outputs(1529) <= (inputs(15)) or (inputs(147));
    layer0_outputs(1530) <= not(inputs(5));
    layer0_outputs(1531) <= not((inputs(74)) xor (inputs(169)));
    layer0_outputs(1532) <= not((inputs(65)) xor (inputs(42)));
    layer0_outputs(1533) <= (inputs(77)) and not (inputs(39));
    layer0_outputs(1534) <= not(inputs(76)) or (inputs(254));
    layer0_outputs(1535) <= (inputs(40)) xor (inputs(76));
    layer0_outputs(1536) <= (inputs(95)) or (inputs(145));
    layer0_outputs(1537) <= (inputs(188)) xor (inputs(123));
    layer0_outputs(1538) <= not((inputs(114)) xor (inputs(151)));
    layer0_outputs(1539) <= inputs(19);
    layer0_outputs(1540) <= (inputs(230)) and not (inputs(88));
    layer0_outputs(1541) <= not((inputs(93)) or (inputs(174)));
    layer0_outputs(1542) <= (inputs(124)) and (inputs(153));
    layer0_outputs(1543) <= (inputs(133)) or (inputs(8));
    layer0_outputs(1544) <= not(inputs(145));
    layer0_outputs(1545) <= not(inputs(24)) or (inputs(181));
    layer0_outputs(1546) <= inputs(200);
    layer0_outputs(1547) <= not((inputs(121)) or (inputs(123)));
    layer0_outputs(1548) <= not(inputs(238));
    layer0_outputs(1549) <= not((inputs(213)) or (inputs(226)));
    layer0_outputs(1550) <= not((inputs(121)) xor (inputs(48)));
    layer0_outputs(1551) <= not(inputs(110));
    layer0_outputs(1552) <= inputs(82);
    layer0_outputs(1553) <= not(inputs(92));
    layer0_outputs(1554) <= inputs(234);
    layer0_outputs(1555) <= (inputs(4)) and not (inputs(58));
    layer0_outputs(1556) <= not((inputs(53)) xor (inputs(42)));
    layer0_outputs(1557) <= not(inputs(196)) or (inputs(40));
    layer0_outputs(1558) <= not(inputs(119));
    layer0_outputs(1559) <= not(inputs(108)) or (inputs(88));
    layer0_outputs(1560) <= not(inputs(118)) or (inputs(88));
    layer0_outputs(1561) <= not((inputs(24)) xor (inputs(21)));
    layer0_outputs(1562) <= inputs(94);
    layer0_outputs(1563) <= not(inputs(75));
    layer0_outputs(1564) <= not(inputs(163));
    layer0_outputs(1565) <= not(inputs(68)) or (inputs(93));
    layer0_outputs(1566) <= inputs(79);
    layer0_outputs(1567) <= inputs(11);
    layer0_outputs(1568) <= not((inputs(154)) or (inputs(25)));
    layer0_outputs(1569) <= (inputs(1)) and not (inputs(241));
    layer0_outputs(1570) <= (inputs(133)) xor (inputs(98));
    layer0_outputs(1571) <= inputs(102);
    layer0_outputs(1572) <= not((inputs(64)) xor (inputs(10)));
    layer0_outputs(1573) <= (inputs(44)) and (inputs(14));
    layer0_outputs(1574) <= (inputs(185)) or (inputs(238));
    layer0_outputs(1575) <= not(inputs(215));
    layer0_outputs(1576) <= not((inputs(67)) or (inputs(68)));
    layer0_outputs(1577) <= (inputs(156)) xor (inputs(207));
    layer0_outputs(1578) <= not((inputs(194)) or (inputs(124)));
    layer0_outputs(1579) <= not(inputs(202));
    layer0_outputs(1580) <= not(inputs(157)) or (inputs(15));
    layer0_outputs(1581) <= not((inputs(30)) xor (inputs(103)));
    layer0_outputs(1582) <= inputs(178);
    layer0_outputs(1583) <= not(inputs(26)) or (inputs(97));
    layer0_outputs(1584) <= (inputs(102)) and not (inputs(235));
    layer0_outputs(1585) <= (inputs(146)) and not (inputs(187));
    layer0_outputs(1586) <= not(inputs(237));
    layer0_outputs(1587) <= (inputs(197)) xor (inputs(185));
    layer0_outputs(1588) <= not(inputs(29)) or (inputs(93));
    layer0_outputs(1589) <= (inputs(20)) xor (inputs(127));
    layer0_outputs(1590) <= inputs(88);
    layer0_outputs(1591) <= (inputs(187)) and not (inputs(83));
    layer0_outputs(1592) <= not(inputs(209)) or (inputs(203));
    layer0_outputs(1593) <= not(inputs(47)) or (inputs(1));
    layer0_outputs(1594) <= not((inputs(121)) xor (inputs(19)));
    layer0_outputs(1595) <= inputs(66);
    layer0_outputs(1596) <= not((inputs(15)) xor (inputs(83)));
    layer0_outputs(1597) <= '0';
    layer0_outputs(1598) <= (inputs(174)) or (inputs(85));
    layer0_outputs(1599) <= (inputs(39)) and not (inputs(17));
    layer0_outputs(1600) <= (inputs(243)) xor (inputs(177));
    layer0_outputs(1601) <= not(inputs(137));
    layer0_outputs(1602) <= not((inputs(30)) or (inputs(83)));
    layer0_outputs(1603) <= not((inputs(4)) xor (inputs(135)));
    layer0_outputs(1604) <= (inputs(56)) and not (inputs(202));
    layer0_outputs(1605) <= not(inputs(133));
    layer0_outputs(1606) <= not(inputs(179)) or (inputs(96));
    layer0_outputs(1607) <= not(inputs(170));
    layer0_outputs(1608) <= (inputs(182)) or (inputs(207));
    layer0_outputs(1609) <= not(inputs(74)) or (inputs(208));
    layer0_outputs(1610) <= inputs(111);
    layer0_outputs(1611) <= not((inputs(59)) or (inputs(242)));
    layer0_outputs(1612) <= not(inputs(116)) or (inputs(76));
    layer0_outputs(1613) <= inputs(108);
    layer0_outputs(1614) <= not((inputs(188)) xor (inputs(180)));
    layer0_outputs(1615) <= not(inputs(182)) or (inputs(222));
    layer0_outputs(1616) <= inputs(216);
    layer0_outputs(1617) <= not((inputs(14)) or (inputs(187)));
    layer0_outputs(1618) <= (inputs(205)) or (inputs(149));
    layer0_outputs(1619) <= not((inputs(252)) or (inputs(34)));
    layer0_outputs(1620) <= (inputs(228)) and not (inputs(104));
    layer0_outputs(1621) <= not((inputs(157)) or (inputs(234)));
    layer0_outputs(1622) <= not(inputs(82));
    layer0_outputs(1623) <= (inputs(203)) and not (inputs(149));
    layer0_outputs(1624) <= (inputs(87)) or (inputs(34));
    layer0_outputs(1625) <= inputs(203);
    layer0_outputs(1626) <= (inputs(235)) and not (inputs(78));
    layer0_outputs(1627) <= (inputs(43)) and not (inputs(188));
    layer0_outputs(1628) <= not(inputs(88));
    layer0_outputs(1629) <= '0';
    layer0_outputs(1630) <= (inputs(153)) xor (inputs(156));
    layer0_outputs(1631) <= not(inputs(89)) or (inputs(128));
    layer0_outputs(1632) <= (inputs(197)) or (inputs(111));
    layer0_outputs(1633) <= (inputs(232)) or (inputs(233));
    layer0_outputs(1634) <= not(inputs(38));
    layer0_outputs(1635) <= (inputs(69)) and not (inputs(80));
    layer0_outputs(1636) <= (inputs(197)) or (inputs(19));
    layer0_outputs(1637) <= inputs(107);
    layer0_outputs(1638) <= inputs(100);
    layer0_outputs(1639) <= not(inputs(241)) or (inputs(33));
    layer0_outputs(1640) <= (inputs(157)) or (inputs(16));
    layer0_outputs(1641) <= (inputs(245)) or (inputs(190));
    layer0_outputs(1642) <= (inputs(142)) and not (inputs(253));
    layer0_outputs(1643) <= (inputs(222)) xor (inputs(60));
    layer0_outputs(1644) <= not((inputs(0)) and (inputs(149)));
    layer0_outputs(1645) <= (inputs(2)) or (inputs(21));
    layer0_outputs(1646) <= (inputs(241)) and not (inputs(103));
    layer0_outputs(1647) <= inputs(152);
    layer0_outputs(1648) <= (inputs(49)) xor (inputs(21));
    layer0_outputs(1649) <= not((inputs(109)) xor (inputs(104)));
    layer0_outputs(1650) <= not((inputs(157)) xor (inputs(169)));
    layer0_outputs(1651) <= (inputs(160)) xor (inputs(160));
    layer0_outputs(1652) <= inputs(62);
    layer0_outputs(1653) <= (inputs(184)) or (inputs(150));
    layer0_outputs(1654) <= inputs(88);
    layer0_outputs(1655) <= not((inputs(213)) and (inputs(248)));
    layer0_outputs(1656) <= not((inputs(15)) xor (inputs(50)));
    layer0_outputs(1657) <= not(inputs(84)) or (inputs(57));
    layer0_outputs(1658) <= (inputs(232)) xor (inputs(218));
    layer0_outputs(1659) <= (inputs(77)) and not (inputs(198));
    layer0_outputs(1660) <= not(inputs(91));
    layer0_outputs(1661) <= not(inputs(255));
    layer0_outputs(1662) <= (inputs(164)) and (inputs(230));
    layer0_outputs(1663) <= not(inputs(186));
    layer0_outputs(1664) <= (inputs(121)) and not (inputs(222));
    layer0_outputs(1665) <= not(inputs(139));
    layer0_outputs(1666) <= not(inputs(148));
    layer0_outputs(1667) <= not(inputs(50)) or (inputs(124));
    layer0_outputs(1668) <= not(inputs(120)) or (inputs(145));
    layer0_outputs(1669) <= (inputs(218)) xor (inputs(192));
    layer0_outputs(1670) <= (inputs(189)) xor (inputs(19));
    layer0_outputs(1671) <= not(inputs(61)) or (inputs(100));
    layer0_outputs(1672) <= (inputs(200)) xor (inputs(197));
    layer0_outputs(1673) <= not(inputs(126)) or (inputs(224));
    layer0_outputs(1674) <= not(inputs(135)) or (inputs(105));
    layer0_outputs(1675) <= (inputs(36)) and not (inputs(158));
    layer0_outputs(1676) <= not(inputs(213));
    layer0_outputs(1677) <= not((inputs(178)) xor (inputs(92)));
    layer0_outputs(1678) <= not(inputs(137)) or (inputs(12));
    layer0_outputs(1679) <= not((inputs(158)) xor (inputs(161)));
    layer0_outputs(1680) <= (inputs(212)) xor (inputs(55));
    layer0_outputs(1681) <= '0';
    layer0_outputs(1682) <= not((inputs(108)) xor (inputs(189)));
    layer0_outputs(1683) <= not((inputs(253)) or (inputs(238)));
    layer0_outputs(1684) <= (inputs(72)) or (inputs(226));
    layer0_outputs(1685) <= not((inputs(227)) or (inputs(209)));
    layer0_outputs(1686) <= inputs(234);
    layer0_outputs(1687) <= inputs(55);
    layer0_outputs(1688) <= (inputs(127)) xor (inputs(219));
    layer0_outputs(1689) <= inputs(207);
    layer0_outputs(1690) <= not(inputs(124));
    layer0_outputs(1691) <= (inputs(69)) and not (inputs(220));
    layer0_outputs(1692) <= (inputs(227)) xor (inputs(80));
    layer0_outputs(1693) <= (inputs(254)) xor (inputs(57));
    layer0_outputs(1694) <= (inputs(229)) and not (inputs(27));
    layer0_outputs(1695) <= not(inputs(184)) or (inputs(100));
    layer0_outputs(1696) <= (inputs(152)) and not (inputs(112));
    layer0_outputs(1697) <= not(inputs(75));
    layer0_outputs(1698) <= inputs(204);
    layer0_outputs(1699) <= not(inputs(205));
    layer0_outputs(1700) <= not((inputs(132)) xor (inputs(145)));
    layer0_outputs(1701) <= '1';
    layer0_outputs(1702) <= not(inputs(166));
    layer0_outputs(1703) <= '1';
    layer0_outputs(1704) <= not(inputs(220));
    layer0_outputs(1705) <= inputs(119);
    layer0_outputs(1706) <= (inputs(50)) or (inputs(243));
    layer0_outputs(1707) <= (inputs(123)) and not (inputs(239));
    layer0_outputs(1708) <= inputs(28);
    layer0_outputs(1709) <= not(inputs(25)) or (inputs(83));
    layer0_outputs(1710) <= not(inputs(185)) or (inputs(72));
    layer0_outputs(1711) <= not((inputs(83)) or (inputs(255)));
    layer0_outputs(1712) <= inputs(7);
    layer0_outputs(1713) <= not((inputs(219)) xor (inputs(64)));
    layer0_outputs(1714) <= not(inputs(167));
    layer0_outputs(1715) <= not((inputs(67)) or (inputs(80)));
    layer0_outputs(1716) <= inputs(117);
    layer0_outputs(1717) <= not((inputs(10)) xor (inputs(30)));
    layer0_outputs(1718) <= inputs(244);
    layer0_outputs(1719) <= not(inputs(246)) or (inputs(81));
    layer0_outputs(1720) <= not((inputs(51)) or (inputs(212)));
    layer0_outputs(1721) <= (inputs(39)) xor (inputs(70));
    layer0_outputs(1722) <= not((inputs(32)) xor (inputs(117)));
    layer0_outputs(1723) <= '1';
    layer0_outputs(1724) <= not((inputs(184)) or (inputs(116)));
    layer0_outputs(1725) <= inputs(131);
    layer0_outputs(1726) <= not(inputs(88));
    layer0_outputs(1727) <= not(inputs(8));
    layer0_outputs(1728) <= (inputs(126)) or (inputs(81));
    layer0_outputs(1729) <= (inputs(229)) and not (inputs(253));
    layer0_outputs(1730) <= (inputs(208)) or (inputs(16));
    layer0_outputs(1731) <= not(inputs(246)) or (inputs(98));
    layer0_outputs(1732) <= not(inputs(150)) or (inputs(113));
    layer0_outputs(1733) <= (inputs(90)) xor (inputs(92));
    layer0_outputs(1734) <= not(inputs(122)) or (inputs(190));
    layer0_outputs(1735) <= not(inputs(179));
    layer0_outputs(1736) <= (inputs(22)) and (inputs(197));
    layer0_outputs(1737) <= inputs(153);
    layer0_outputs(1738) <= (inputs(214)) xor (inputs(213));
    layer0_outputs(1739) <= not((inputs(94)) xor (inputs(112)));
    layer0_outputs(1740) <= not((inputs(251)) and (inputs(159)));
    layer0_outputs(1741) <= inputs(144);
    layer0_outputs(1742) <= not(inputs(23));
    layer0_outputs(1743) <= not(inputs(178)) or (inputs(219));
    layer0_outputs(1744) <= not(inputs(2));
    layer0_outputs(1745) <= (inputs(7)) or (inputs(0));
    layer0_outputs(1746) <= not(inputs(64)) or (inputs(252));
    layer0_outputs(1747) <= not(inputs(161));
    layer0_outputs(1748) <= (inputs(175)) or (inputs(252));
    layer0_outputs(1749) <= '1';
    layer0_outputs(1750) <= not((inputs(179)) and (inputs(247)));
    layer0_outputs(1751) <= (inputs(226)) or (inputs(234));
    layer0_outputs(1752) <= (inputs(169)) and not (inputs(79));
    layer0_outputs(1753) <= not(inputs(9));
    layer0_outputs(1754) <= not(inputs(242)) or (inputs(4));
    layer0_outputs(1755) <= not(inputs(219));
    layer0_outputs(1756) <= not(inputs(14));
    layer0_outputs(1757) <= not(inputs(200)) or (inputs(8));
    layer0_outputs(1758) <= inputs(65);
    layer0_outputs(1759) <= (inputs(7)) xor (inputs(160));
    layer0_outputs(1760) <= not(inputs(136)) or (inputs(23));
    layer0_outputs(1761) <= (inputs(2)) xor (inputs(213));
    layer0_outputs(1762) <= inputs(70);
    layer0_outputs(1763) <= not(inputs(95));
    layer0_outputs(1764) <= (inputs(102)) xor (inputs(62));
    layer0_outputs(1765) <= (inputs(186)) and not (inputs(226));
    layer0_outputs(1766) <= not((inputs(178)) or (inputs(156)));
    layer0_outputs(1767) <= (inputs(199)) or (inputs(19));
    layer0_outputs(1768) <= (inputs(169)) or (inputs(236));
    layer0_outputs(1769) <= (inputs(94)) or (inputs(55));
    layer0_outputs(1770) <= (inputs(133)) and not (inputs(158));
    layer0_outputs(1771) <= (inputs(60)) or (inputs(14));
    layer0_outputs(1772) <= (inputs(5)) xor (inputs(174));
    layer0_outputs(1773) <= (inputs(89)) or (inputs(104));
    layer0_outputs(1774) <= (inputs(66)) and not (inputs(97));
    layer0_outputs(1775) <= inputs(164);
    layer0_outputs(1776) <= not(inputs(212)) or (inputs(109));
    layer0_outputs(1777) <= not(inputs(95));
    layer0_outputs(1778) <= inputs(73);
    layer0_outputs(1779) <= inputs(200);
    layer0_outputs(1780) <= (inputs(104)) and not (inputs(235));
    layer0_outputs(1781) <= not((inputs(14)) and (inputs(121)));
    layer0_outputs(1782) <= (inputs(4)) xor (inputs(49));
    layer0_outputs(1783) <= not(inputs(110));
    layer0_outputs(1784) <= not(inputs(231)) or (inputs(128));
    layer0_outputs(1785) <= not(inputs(19)) or (inputs(223));
    layer0_outputs(1786) <= not((inputs(164)) or (inputs(148)));
    layer0_outputs(1787) <= not((inputs(84)) xor (inputs(147)));
    layer0_outputs(1788) <= not((inputs(177)) xor (inputs(185)));
    layer0_outputs(1789) <= '1';
    layer0_outputs(1790) <= not((inputs(101)) or (inputs(35)));
    layer0_outputs(1791) <= inputs(95);
    layer0_outputs(1792) <= inputs(141);
    layer0_outputs(1793) <= inputs(80);
    layer0_outputs(1794) <= not((inputs(10)) xor (inputs(15)));
    layer0_outputs(1795) <= inputs(122);
    layer0_outputs(1796) <= (inputs(130)) or (inputs(217));
    layer0_outputs(1797) <= (inputs(151)) and not (inputs(154));
    layer0_outputs(1798) <= '0';
    layer0_outputs(1799) <= not(inputs(89)) or (inputs(255));
    layer0_outputs(1800) <= inputs(132);
    layer0_outputs(1801) <= not(inputs(221));
    layer0_outputs(1802) <= inputs(178);
    layer0_outputs(1803) <= not(inputs(231)) or (inputs(252));
    layer0_outputs(1804) <= not((inputs(184)) xor (inputs(174)));
    layer0_outputs(1805) <= not(inputs(132));
    layer0_outputs(1806) <= not((inputs(139)) xor (inputs(76)));
    layer0_outputs(1807) <= (inputs(74)) or (inputs(111));
    layer0_outputs(1808) <= (inputs(248)) and not (inputs(31));
    layer0_outputs(1809) <= inputs(26);
    layer0_outputs(1810) <= (inputs(146)) and (inputs(162));
    layer0_outputs(1811) <= inputs(152);
    layer0_outputs(1812) <= inputs(53);
    layer0_outputs(1813) <= (inputs(70)) or (inputs(129));
    layer0_outputs(1814) <= (inputs(179)) and not (inputs(71));
    layer0_outputs(1815) <= (inputs(98)) or (inputs(54));
    layer0_outputs(1816) <= (inputs(132)) or (inputs(14));
    layer0_outputs(1817) <= not((inputs(37)) and (inputs(156)));
    layer0_outputs(1818) <= (inputs(99)) and not (inputs(134));
    layer0_outputs(1819) <= inputs(249);
    layer0_outputs(1820) <= inputs(120);
    layer0_outputs(1821) <= inputs(151);
    layer0_outputs(1822) <= inputs(230);
    layer0_outputs(1823) <= not(inputs(53)) or (inputs(127));
    layer0_outputs(1824) <= not(inputs(163));
    layer0_outputs(1825) <= inputs(184);
    layer0_outputs(1826) <= not(inputs(75));
    layer0_outputs(1827) <= not(inputs(239)) or (inputs(72));
    layer0_outputs(1828) <= (inputs(234)) or (inputs(176));
    layer0_outputs(1829) <= (inputs(209)) xor (inputs(160));
    layer0_outputs(1830) <= not(inputs(81));
    layer0_outputs(1831) <= inputs(49);
    layer0_outputs(1832) <= (inputs(239)) or (inputs(160));
    layer0_outputs(1833) <= inputs(247);
    layer0_outputs(1834) <= (inputs(178)) xor (inputs(235));
    layer0_outputs(1835) <= (inputs(83)) and not (inputs(15));
    layer0_outputs(1836) <= not((inputs(71)) xor (inputs(41)));
    layer0_outputs(1837) <= inputs(184);
    layer0_outputs(1838) <= inputs(148);
    layer0_outputs(1839) <= (inputs(73)) and not (inputs(140));
    layer0_outputs(1840) <= (inputs(183)) or (inputs(113));
    layer0_outputs(1841) <= not(inputs(186));
    layer0_outputs(1842) <= inputs(115);
    layer0_outputs(1843) <= inputs(77);
    layer0_outputs(1844) <= not((inputs(42)) and (inputs(150)));
    layer0_outputs(1845) <= inputs(78);
    layer0_outputs(1846) <= not((inputs(197)) or (inputs(112)));
    layer0_outputs(1847) <= not((inputs(57)) or (inputs(209)));
    layer0_outputs(1848) <= (inputs(173)) or (inputs(174));
    layer0_outputs(1849) <= (inputs(194)) and not (inputs(102));
    layer0_outputs(1850) <= not((inputs(28)) xor (inputs(9)));
    layer0_outputs(1851) <= not((inputs(120)) or (inputs(225)));
    layer0_outputs(1852) <= not(inputs(22));
    layer0_outputs(1853) <= (inputs(181)) or (inputs(73));
    layer0_outputs(1854) <= not((inputs(18)) and (inputs(89)));
    layer0_outputs(1855) <= inputs(147);
    layer0_outputs(1856) <= inputs(26);
    layer0_outputs(1857) <= not(inputs(55)) or (inputs(175));
    layer0_outputs(1858) <= not(inputs(120));
    layer0_outputs(1859) <= '0';
    layer0_outputs(1860) <= (inputs(213)) and not (inputs(85));
    layer0_outputs(1861) <= (inputs(151)) or (inputs(135));
    layer0_outputs(1862) <= not((inputs(194)) or (inputs(158)));
    layer0_outputs(1863) <= (inputs(95)) or (inputs(179));
    layer0_outputs(1864) <= inputs(78);
    layer0_outputs(1865) <= not(inputs(62)) or (inputs(41));
    layer0_outputs(1866) <= not((inputs(154)) or (inputs(125)));
    layer0_outputs(1867) <= not((inputs(14)) xor (inputs(184)));
    layer0_outputs(1868) <= not((inputs(13)) or (inputs(83)));
    layer0_outputs(1869) <= not((inputs(113)) or (inputs(175)));
    layer0_outputs(1870) <= (inputs(165)) xor (inputs(56));
    layer0_outputs(1871) <= not((inputs(228)) and (inputs(96)));
    layer0_outputs(1872) <= (inputs(48)) and not (inputs(21));
    layer0_outputs(1873) <= (inputs(80)) xor (inputs(66));
    layer0_outputs(1874) <= inputs(94);
    layer0_outputs(1875) <= inputs(136);
    layer0_outputs(1876) <= inputs(85);
    layer0_outputs(1877) <= not(inputs(134));
    layer0_outputs(1878) <= inputs(234);
    layer0_outputs(1879) <= inputs(204);
    layer0_outputs(1880) <= inputs(72);
    layer0_outputs(1881) <= inputs(14);
    layer0_outputs(1882) <= (inputs(101)) and not (inputs(233));
    layer0_outputs(1883) <= not((inputs(222)) or (inputs(50)));
    layer0_outputs(1884) <= inputs(234);
    layer0_outputs(1885) <= not(inputs(80));
    layer0_outputs(1886) <= inputs(60);
    layer0_outputs(1887) <= not(inputs(186));
    layer0_outputs(1888) <= not(inputs(135)) or (inputs(57));
    layer0_outputs(1889) <= inputs(170);
    layer0_outputs(1890) <= (inputs(143)) or (inputs(197));
    layer0_outputs(1891) <= (inputs(198)) xor (inputs(135));
    layer0_outputs(1892) <= (inputs(5)) or (inputs(185));
    layer0_outputs(1893) <= not((inputs(14)) or (inputs(221)));
    layer0_outputs(1894) <= not((inputs(78)) or (inputs(13)));
    layer0_outputs(1895) <= not((inputs(163)) or (inputs(176)));
    layer0_outputs(1896) <= not(inputs(187)) or (inputs(224));
    layer0_outputs(1897) <= inputs(56);
    layer0_outputs(1898) <= not(inputs(182)) or (inputs(139));
    layer0_outputs(1899) <= not(inputs(25)) or (inputs(0));
    layer0_outputs(1900) <= (inputs(61)) or (inputs(141));
    layer0_outputs(1901) <= not(inputs(117));
    layer0_outputs(1902) <= not(inputs(147)) or (inputs(137));
    layer0_outputs(1903) <= not(inputs(70));
    layer0_outputs(1904) <= not((inputs(217)) xor (inputs(250)));
    layer0_outputs(1905) <= not((inputs(91)) xor (inputs(176)));
    layer0_outputs(1906) <= not((inputs(8)) xor (inputs(179)));
    layer0_outputs(1907) <= (inputs(18)) or (inputs(37));
    layer0_outputs(1908) <= not(inputs(157)) or (inputs(241));
    layer0_outputs(1909) <= inputs(237);
    layer0_outputs(1910) <= (inputs(167)) and not (inputs(93));
    layer0_outputs(1911) <= inputs(252);
    layer0_outputs(1912) <= inputs(102);
    layer0_outputs(1913) <= not(inputs(56));
    layer0_outputs(1914) <= inputs(150);
    layer0_outputs(1915) <= inputs(60);
    layer0_outputs(1916) <= inputs(15);
    layer0_outputs(1917) <= not((inputs(131)) or (inputs(72)));
    layer0_outputs(1918) <= inputs(218);
    layer0_outputs(1919) <= (inputs(141)) xor (inputs(160));
    layer0_outputs(1920) <= inputs(209);
    layer0_outputs(1921) <= not(inputs(130));
    layer0_outputs(1922) <= not((inputs(242)) xor (inputs(143)));
    layer0_outputs(1923) <= (inputs(163)) and not (inputs(33));
    layer0_outputs(1924) <= (inputs(244)) and not (inputs(182));
    layer0_outputs(1925) <= not(inputs(78));
    layer0_outputs(1926) <= not(inputs(186));
    layer0_outputs(1927) <= (inputs(140)) xor (inputs(223));
    layer0_outputs(1928) <= '0';
    layer0_outputs(1929) <= not((inputs(210)) or (inputs(94)));
    layer0_outputs(1930) <= inputs(172);
    layer0_outputs(1931) <= (inputs(122)) xor (inputs(179));
    layer0_outputs(1932) <= (inputs(207)) and not (inputs(48));
    layer0_outputs(1933) <= inputs(60);
    layer0_outputs(1934) <= not(inputs(120));
    layer0_outputs(1935) <= inputs(234);
    layer0_outputs(1936) <= (inputs(44)) and not (inputs(232));
    layer0_outputs(1937) <= not((inputs(243)) xor (inputs(43)));
    layer0_outputs(1938) <= inputs(67);
    layer0_outputs(1939) <= not((inputs(238)) or (inputs(222)));
    layer0_outputs(1940) <= not((inputs(98)) xor (inputs(21)));
    layer0_outputs(1941) <= not(inputs(160));
    layer0_outputs(1942) <= inputs(86);
    layer0_outputs(1943) <= not(inputs(94));
    layer0_outputs(1944) <= not((inputs(98)) or (inputs(46)));
    layer0_outputs(1945) <= (inputs(184)) xor (inputs(139));
    layer0_outputs(1946) <= (inputs(1)) xor (inputs(210));
    layer0_outputs(1947) <= not(inputs(84));
    layer0_outputs(1948) <= inputs(167);
    layer0_outputs(1949) <= not(inputs(189));
    layer0_outputs(1950) <= not(inputs(185));
    layer0_outputs(1951) <= not((inputs(211)) xor (inputs(44)));
    layer0_outputs(1952) <= not(inputs(3)) or (inputs(239));
    layer0_outputs(1953) <= not(inputs(224));
    layer0_outputs(1954) <= (inputs(123)) and not (inputs(162));
    layer0_outputs(1955) <= not(inputs(97));
    layer0_outputs(1956) <= not((inputs(110)) or (inputs(160)));
    layer0_outputs(1957) <= (inputs(64)) xor (inputs(156));
    layer0_outputs(1958) <= (inputs(194)) xor (inputs(180));
    layer0_outputs(1959) <= (inputs(116)) xor (inputs(136));
    layer0_outputs(1960) <= not(inputs(86));
    layer0_outputs(1961) <= (inputs(177)) and not (inputs(134));
    layer0_outputs(1962) <= (inputs(197)) xor (inputs(231));
    layer0_outputs(1963) <= not((inputs(189)) xor (inputs(174)));
    layer0_outputs(1964) <= not((inputs(125)) or (inputs(112)));
    layer0_outputs(1965) <= (inputs(14)) and not (inputs(142));
    layer0_outputs(1966) <= (inputs(48)) and (inputs(125));
    layer0_outputs(1967) <= inputs(103);
    layer0_outputs(1968) <= not(inputs(42));
    layer0_outputs(1969) <= inputs(84);
    layer0_outputs(1970) <= inputs(0);
    layer0_outputs(1971) <= (inputs(158)) xor (inputs(18));
    layer0_outputs(1972) <= (inputs(197)) and not (inputs(15));
    layer0_outputs(1973) <= not(inputs(232));
    layer0_outputs(1974) <= not(inputs(85));
    layer0_outputs(1975) <= not((inputs(216)) or (inputs(190)));
    layer0_outputs(1976) <= not((inputs(22)) and (inputs(39)));
    layer0_outputs(1977) <= not((inputs(236)) or (inputs(234)));
    layer0_outputs(1978) <= not(inputs(214));
    layer0_outputs(1979) <= not((inputs(251)) or (inputs(162)));
    layer0_outputs(1980) <= '0';
    layer0_outputs(1981) <= not(inputs(123));
    layer0_outputs(1982) <= not((inputs(129)) xor (inputs(39)));
    layer0_outputs(1983) <= not((inputs(172)) or (inputs(115)));
    layer0_outputs(1984) <= inputs(180);
    layer0_outputs(1985) <= not((inputs(182)) or (inputs(221)));
    layer0_outputs(1986) <= inputs(168);
    layer0_outputs(1987) <= not(inputs(143)) or (inputs(185));
    layer0_outputs(1988) <= (inputs(3)) and (inputs(53));
    layer0_outputs(1989) <= not(inputs(140)) or (inputs(19));
    layer0_outputs(1990) <= (inputs(53)) xor (inputs(168));
    layer0_outputs(1991) <= not(inputs(194));
    layer0_outputs(1992) <= (inputs(158)) and not (inputs(15));
    layer0_outputs(1993) <= not(inputs(58));
    layer0_outputs(1994) <= inputs(198);
    layer0_outputs(1995) <= not(inputs(19)) or (inputs(128));
    layer0_outputs(1996) <= (inputs(194)) or (inputs(147));
    layer0_outputs(1997) <= (inputs(71)) and not (inputs(97));
    layer0_outputs(1998) <= not(inputs(155));
    layer0_outputs(1999) <= inputs(178);
    layer0_outputs(2000) <= not((inputs(152)) and (inputs(145)));
    layer0_outputs(2001) <= not(inputs(234));
    layer0_outputs(2002) <= not((inputs(44)) or (inputs(5)));
    layer0_outputs(2003) <= (inputs(254)) or (inputs(98));
    layer0_outputs(2004) <= inputs(168);
    layer0_outputs(2005) <= inputs(21);
    layer0_outputs(2006) <= not((inputs(143)) or (inputs(157)));
    layer0_outputs(2007) <= inputs(89);
    layer0_outputs(2008) <= inputs(42);
    layer0_outputs(2009) <= (inputs(6)) or (inputs(110));
    layer0_outputs(2010) <= not(inputs(231)) or (inputs(110));
    layer0_outputs(2011) <= not(inputs(27));
    layer0_outputs(2012) <= not(inputs(89)) or (inputs(113));
    layer0_outputs(2013) <= (inputs(60)) or (inputs(11));
    layer0_outputs(2014) <= (inputs(153)) or (inputs(152));
    layer0_outputs(2015) <= not(inputs(37)) or (inputs(187));
    layer0_outputs(2016) <= not((inputs(231)) xor (inputs(184)));
    layer0_outputs(2017) <= not((inputs(193)) and (inputs(131)));
    layer0_outputs(2018) <= not(inputs(108));
    layer0_outputs(2019) <= inputs(55);
    layer0_outputs(2020) <= (inputs(37)) and not (inputs(213));
    layer0_outputs(2021) <= (inputs(175)) or (inputs(112));
    layer0_outputs(2022) <= not((inputs(203)) xor (inputs(108)));
    layer0_outputs(2023) <= not(inputs(97)) or (inputs(241));
    layer0_outputs(2024) <= not(inputs(165));
    layer0_outputs(2025) <= not((inputs(189)) xor (inputs(109)));
    layer0_outputs(2026) <= (inputs(231)) xor (inputs(198));
    layer0_outputs(2027) <= (inputs(8)) or (inputs(84));
    layer0_outputs(2028) <= (inputs(74)) and (inputs(140));
    layer0_outputs(2029) <= inputs(40);
    layer0_outputs(2030) <= (inputs(23)) xor (inputs(96));
    layer0_outputs(2031) <= (inputs(202)) and (inputs(167));
    layer0_outputs(2032) <= (inputs(124)) and (inputs(230));
    layer0_outputs(2033) <= not((inputs(95)) or (inputs(241)));
    layer0_outputs(2034) <= (inputs(68)) xor (inputs(141));
    layer0_outputs(2035) <= not(inputs(21)) or (inputs(147));
    layer0_outputs(2036) <= (inputs(40)) and not (inputs(84));
    layer0_outputs(2037) <= (inputs(100)) and not (inputs(239));
    layer0_outputs(2038) <= inputs(103);
    layer0_outputs(2039) <= (inputs(179)) and not (inputs(31));
    layer0_outputs(2040) <= not(inputs(217));
    layer0_outputs(2041) <= (inputs(184)) and not (inputs(117));
    layer0_outputs(2042) <= inputs(107);
    layer0_outputs(2043) <= not((inputs(225)) xor (inputs(180)));
    layer0_outputs(2044) <= not((inputs(80)) xor (inputs(84)));
    layer0_outputs(2045) <= not((inputs(182)) or (inputs(14)));
    layer0_outputs(2046) <= not(inputs(17)) or (inputs(18));
    layer0_outputs(2047) <= inputs(117);
    layer0_outputs(2048) <= (inputs(185)) xor (inputs(216));
    layer0_outputs(2049) <= not(inputs(246));
    layer0_outputs(2050) <= (inputs(52)) and not (inputs(17));
    layer0_outputs(2051) <= (inputs(209)) or (inputs(110));
    layer0_outputs(2052) <= not(inputs(196));
    layer0_outputs(2053) <= (inputs(200)) or (inputs(65));
    layer0_outputs(2054) <= not(inputs(115));
    layer0_outputs(2055) <= (inputs(37)) and not (inputs(129));
    layer0_outputs(2056) <= (inputs(132)) and not (inputs(151));
    layer0_outputs(2057) <= (inputs(200)) xor (inputs(250));
    layer0_outputs(2058) <= not(inputs(203));
    layer0_outputs(2059) <= not(inputs(58));
    layer0_outputs(2060) <= inputs(118);
    layer0_outputs(2061) <= not(inputs(140)) or (inputs(152));
    layer0_outputs(2062) <= '0';
    layer0_outputs(2063) <= inputs(35);
    layer0_outputs(2064) <= not(inputs(108));
    layer0_outputs(2065) <= (inputs(158)) or (inputs(19));
    layer0_outputs(2066) <= not(inputs(206)) or (inputs(129));
    layer0_outputs(2067) <= (inputs(212)) and not (inputs(98));
    layer0_outputs(2068) <= not((inputs(197)) or (inputs(245)));
    layer0_outputs(2069) <= (inputs(111)) and not (inputs(252));
    layer0_outputs(2070) <= not((inputs(1)) or (inputs(79)));
    layer0_outputs(2071) <= not(inputs(100)) or (inputs(190));
    layer0_outputs(2072) <= (inputs(43)) or (inputs(224));
    layer0_outputs(2073) <= (inputs(131)) or (inputs(129));
    layer0_outputs(2074) <= (inputs(15)) xor (inputs(12));
    layer0_outputs(2075) <= not(inputs(56));
    layer0_outputs(2076) <= not((inputs(94)) xor (inputs(103)));
    layer0_outputs(2077) <= not((inputs(13)) xor (inputs(144)));
    layer0_outputs(2078) <= not(inputs(103)) or (inputs(139));
    layer0_outputs(2079) <= (inputs(60)) xor (inputs(91));
    layer0_outputs(2080) <= inputs(118);
    layer0_outputs(2081) <= (inputs(219)) and not (inputs(124));
    layer0_outputs(2082) <= inputs(99);
    layer0_outputs(2083) <= not(inputs(177));
    layer0_outputs(2084) <= (inputs(106)) xor (inputs(79));
    layer0_outputs(2085) <= not(inputs(228)) or (inputs(30));
    layer0_outputs(2086) <= not((inputs(3)) and (inputs(114)));
    layer0_outputs(2087) <= (inputs(84)) or (inputs(69));
    layer0_outputs(2088) <= inputs(109);
    layer0_outputs(2089) <= (inputs(227)) and not (inputs(80));
    layer0_outputs(2090) <= (inputs(170)) and not (inputs(98));
    layer0_outputs(2091) <= not((inputs(126)) or (inputs(36)));
    layer0_outputs(2092) <= (inputs(242)) or (inputs(129));
    layer0_outputs(2093) <= not(inputs(95));
    layer0_outputs(2094) <= (inputs(224)) or (inputs(78));
    layer0_outputs(2095) <= not(inputs(211));
    layer0_outputs(2096) <= (inputs(174)) xor (inputs(132));
    layer0_outputs(2097) <= '1';
    layer0_outputs(2098) <= inputs(226);
    layer0_outputs(2099) <= (inputs(105)) xor (inputs(178));
    layer0_outputs(2100) <= not((inputs(5)) or (inputs(80)));
    layer0_outputs(2101) <= inputs(124);
    layer0_outputs(2102) <= (inputs(44)) and not (inputs(200));
    layer0_outputs(2103) <= (inputs(213)) or (inputs(153));
    layer0_outputs(2104) <= not((inputs(206)) or (inputs(71)));
    layer0_outputs(2105) <= (inputs(165)) and (inputs(10));
    layer0_outputs(2106) <= inputs(160);
    layer0_outputs(2107) <= not((inputs(214)) xor (inputs(161)));
    layer0_outputs(2108) <= not((inputs(214)) or (inputs(63)));
    layer0_outputs(2109) <= not((inputs(159)) or (inputs(242)));
    layer0_outputs(2110) <= inputs(84);
    layer0_outputs(2111) <= (inputs(152)) and not (inputs(204));
    layer0_outputs(2112) <= not(inputs(181));
    layer0_outputs(2113) <= (inputs(103)) and not (inputs(222));
    layer0_outputs(2114) <= inputs(106);
    layer0_outputs(2115) <= (inputs(195)) xor (inputs(206));
    layer0_outputs(2116) <= not((inputs(200)) xor (inputs(191)));
    layer0_outputs(2117) <= not(inputs(26)) or (inputs(193));
    layer0_outputs(2118) <= not(inputs(53));
    layer0_outputs(2119) <= (inputs(132)) xor (inputs(167));
    layer0_outputs(2120) <= not(inputs(149));
    layer0_outputs(2121) <= inputs(70);
    layer0_outputs(2122) <= inputs(13);
    layer0_outputs(2123) <= (inputs(160)) and not (inputs(49));
    layer0_outputs(2124) <= (inputs(54)) and not (inputs(11));
    layer0_outputs(2125) <= not(inputs(80));
    layer0_outputs(2126) <= not(inputs(67)) or (inputs(63));
    layer0_outputs(2127) <= not(inputs(92)) or (inputs(2));
    layer0_outputs(2128) <= not(inputs(69)) or (inputs(0));
    layer0_outputs(2129) <= (inputs(215)) xor (inputs(77));
    layer0_outputs(2130) <= (inputs(143)) xor (inputs(108));
    layer0_outputs(2131) <= not((inputs(41)) or (inputs(137)));
    layer0_outputs(2132) <= (inputs(24)) or (inputs(16));
    layer0_outputs(2133) <= not(inputs(67));
    layer0_outputs(2134) <= inputs(246);
    layer0_outputs(2135) <= not((inputs(154)) and (inputs(136)));
    layer0_outputs(2136) <= not((inputs(106)) or (inputs(31)));
    layer0_outputs(2137) <= not(inputs(158));
    layer0_outputs(2138) <= inputs(75);
    layer0_outputs(2139) <= (inputs(214)) and (inputs(39));
    layer0_outputs(2140) <= (inputs(236)) or (inputs(33));
    layer0_outputs(2141) <= inputs(188);
    layer0_outputs(2142) <= not((inputs(243)) xor (inputs(247)));
    layer0_outputs(2143) <= (inputs(191)) or (inputs(115));
    layer0_outputs(2144) <= (inputs(8)) or (inputs(23));
    layer0_outputs(2145) <= inputs(238);
    layer0_outputs(2146) <= not((inputs(5)) xor (inputs(168)));
    layer0_outputs(2147) <= not(inputs(24)) or (inputs(191));
    layer0_outputs(2148) <= inputs(101);
    layer0_outputs(2149) <= not(inputs(122));
    layer0_outputs(2150) <= (inputs(105)) or (inputs(139));
    layer0_outputs(2151) <= not((inputs(245)) or (inputs(220)));
    layer0_outputs(2152) <= not((inputs(41)) or (inputs(92)));
    layer0_outputs(2153) <= not(inputs(108)) or (inputs(232));
    layer0_outputs(2154) <= (inputs(4)) and not (inputs(178));
    layer0_outputs(2155) <= not((inputs(253)) or (inputs(197)));
    layer0_outputs(2156) <= (inputs(12)) or (inputs(132));
    layer0_outputs(2157) <= not((inputs(129)) xor (inputs(101)));
    layer0_outputs(2158) <= (inputs(5)) or (inputs(236));
    layer0_outputs(2159) <= (inputs(185)) and (inputs(243));
    layer0_outputs(2160) <= not(inputs(155)) or (inputs(80));
    layer0_outputs(2161) <= (inputs(146)) or (inputs(174));
    layer0_outputs(2162) <= not((inputs(79)) xor (inputs(188)));
    layer0_outputs(2163) <= not(inputs(42)) or (inputs(65));
    layer0_outputs(2164) <= (inputs(113)) or (inputs(0));
    layer0_outputs(2165) <= (inputs(107)) and not (inputs(57));
    layer0_outputs(2166) <= not((inputs(210)) or (inputs(223)));
    layer0_outputs(2167) <= not((inputs(146)) and (inputs(67)));
    layer0_outputs(2168) <= (inputs(185)) or (inputs(51));
    layer0_outputs(2169) <= not(inputs(10));
    layer0_outputs(2170) <= not((inputs(42)) xor (inputs(59)));
    layer0_outputs(2171) <= inputs(29);
    layer0_outputs(2172) <= (inputs(107)) and not (inputs(6));
    layer0_outputs(2173) <= not(inputs(141));
    layer0_outputs(2174) <= (inputs(95)) and not (inputs(236));
    layer0_outputs(2175) <= (inputs(145)) or (inputs(60));
    layer0_outputs(2176) <= not(inputs(242)) or (inputs(169));
    layer0_outputs(2177) <= (inputs(29)) and (inputs(11));
    layer0_outputs(2178) <= inputs(162);
    layer0_outputs(2179) <= not((inputs(144)) or (inputs(175)));
    layer0_outputs(2180) <= '0';
    layer0_outputs(2181) <= (inputs(52)) xor (inputs(120));
    layer0_outputs(2182) <= not((inputs(130)) or (inputs(146)));
    layer0_outputs(2183) <= (inputs(250)) or (inputs(81));
    layer0_outputs(2184) <= (inputs(88)) xor (inputs(102));
    layer0_outputs(2185) <= (inputs(200)) or (inputs(245));
    layer0_outputs(2186) <= inputs(31);
    layer0_outputs(2187) <= inputs(113);
    layer0_outputs(2188) <= (inputs(121)) and not (inputs(77));
    layer0_outputs(2189) <= inputs(81);
    layer0_outputs(2190) <= not((inputs(57)) or (inputs(143)));
    layer0_outputs(2191) <= not(inputs(153));
    layer0_outputs(2192) <= inputs(72);
    layer0_outputs(2193) <= not(inputs(125));
    layer0_outputs(2194) <= inputs(181);
    layer0_outputs(2195) <= inputs(8);
    layer0_outputs(2196) <= not(inputs(122)) or (inputs(242));
    layer0_outputs(2197) <= not((inputs(213)) and (inputs(137)));
    layer0_outputs(2198) <= not(inputs(73));
    layer0_outputs(2199) <= (inputs(10)) xor (inputs(52));
    layer0_outputs(2200) <= not((inputs(126)) or (inputs(62)));
    layer0_outputs(2201) <= (inputs(9)) and not (inputs(72));
    layer0_outputs(2202) <= inputs(142);
    layer0_outputs(2203) <= not(inputs(230));
    layer0_outputs(2204) <= (inputs(96)) and (inputs(44));
    layer0_outputs(2205) <= not((inputs(219)) xor (inputs(71)));
    layer0_outputs(2206) <= not(inputs(183));
    layer0_outputs(2207) <= (inputs(72)) or (inputs(16));
    layer0_outputs(2208) <= (inputs(14)) or (inputs(30));
    layer0_outputs(2209) <= (inputs(138)) and (inputs(167));
    layer0_outputs(2210) <= (inputs(225)) xor (inputs(56));
    layer0_outputs(2211) <= (inputs(115)) and not (inputs(63));
    layer0_outputs(2212) <= not(inputs(193));
    layer0_outputs(2213) <= not(inputs(53));
    layer0_outputs(2214) <= inputs(109);
    layer0_outputs(2215) <= not(inputs(76)) or (inputs(71));
    layer0_outputs(2216) <= (inputs(48)) xor (inputs(160));
    layer0_outputs(2217) <= (inputs(52)) or (inputs(98));
    layer0_outputs(2218) <= (inputs(78)) xor (inputs(190));
    layer0_outputs(2219) <= not((inputs(211)) or (inputs(199)));
    layer0_outputs(2220) <= inputs(241);
    layer0_outputs(2221) <= not(inputs(84)) or (inputs(215));
    layer0_outputs(2222) <= not(inputs(206));
    layer0_outputs(2223) <= not(inputs(82));
    layer0_outputs(2224) <= not(inputs(27));
    layer0_outputs(2225) <= (inputs(63)) or (inputs(170));
    layer0_outputs(2226) <= (inputs(47)) and (inputs(126));
    layer0_outputs(2227) <= inputs(151);
    layer0_outputs(2228) <= inputs(131);
    layer0_outputs(2229) <= (inputs(142)) or (inputs(39));
    layer0_outputs(2230) <= not((inputs(218)) or (inputs(202)));
    layer0_outputs(2231) <= not((inputs(180)) or (inputs(115)));
    layer0_outputs(2232) <= inputs(183);
    layer0_outputs(2233) <= (inputs(71)) and not (inputs(64));
    layer0_outputs(2234) <= not(inputs(112)) or (inputs(165));
    layer0_outputs(2235) <= not(inputs(164));
    layer0_outputs(2236) <= not(inputs(142)) or (inputs(238));
    layer0_outputs(2237) <= not(inputs(82));
    layer0_outputs(2238) <= (inputs(234)) xor (inputs(80));
    layer0_outputs(2239) <= '1';
    layer0_outputs(2240) <= not((inputs(71)) and (inputs(71)));
    layer0_outputs(2241) <= (inputs(46)) xor (inputs(213));
    layer0_outputs(2242) <= (inputs(67)) and not (inputs(150));
    layer0_outputs(2243) <= not(inputs(132));
    layer0_outputs(2244) <= inputs(151);
    layer0_outputs(2245) <= not(inputs(230));
    layer0_outputs(2246) <= inputs(233);
    layer0_outputs(2247) <= not(inputs(248)) or (inputs(126));
    layer0_outputs(2248) <= inputs(101);
    layer0_outputs(2249) <= inputs(163);
    layer0_outputs(2250) <= not(inputs(92));
    layer0_outputs(2251) <= '0';
    layer0_outputs(2252) <= not((inputs(234)) or (inputs(123)));
    layer0_outputs(2253) <= (inputs(99)) xor (inputs(131));
    layer0_outputs(2254) <= not(inputs(233)) or (inputs(149));
    layer0_outputs(2255) <= (inputs(195)) xor (inputs(145));
    layer0_outputs(2256) <= not(inputs(154));
    layer0_outputs(2257) <= (inputs(185)) and not (inputs(247));
    layer0_outputs(2258) <= not((inputs(87)) or (inputs(208)));
    layer0_outputs(2259) <= (inputs(179)) or (inputs(131));
    layer0_outputs(2260) <= not((inputs(105)) xor (inputs(196)));
    layer0_outputs(2261) <= not(inputs(120)) or (inputs(158));
    layer0_outputs(2262) <= not((inputs(24)) and (inputs(229)));
    layer0_outputs(2263) <= (inputs(4)) and not (inputs(94));
    layer0_outputs(2264) <= (inputs(58)) xor (inputs(62));
    layer0_outputs(2265) <= '1';
    layer0_outputs(2266) <= not((inputs(64)) xor (inputs(197)));
    layer0_outputs(2267) <= not((inputs(27)) or (inputs(110)));
    layer0_outputs(2268) <= not(inputs(232));
    layer0_outputs(2269) <= '0';
    layer0_outputs(2270) <= not(inputs(193));
    layer0_outputs(2271) <= (inputs(49)) or (inputs(66));
    layer0_outputs(2272) <= (inputs(73)) xor (inputs(61));
    layer0_outputs(2273) <= not((inputs(142)) or (inputs(39)));
    layer0_outputs(2274) <= (inputs(90)) and not (inputs(205));
    layer0_outputs(2275) <= (inputs(104)) xor (inputs(95));
    layer0_outputs(2276) <= not((inputs(235)) xor (inputs(230)));
    layer0_outputs(2277) <= not((inputs(156)) xor (inputs(99)));
    layer0_outputs(2278) <= inputs(90);
    layer0_outputs(2279) <= not((inputs(62)) or (inputs(100)));
    layer0_outputs(2280) <= not(inputs(215)) or (inputs(192));
    layer0_outputs(2281) <= (inputs(146)) xor (inputs(220));
    layer0_outputs(2282) <= (inputs(174)) or (inputs(198));
    layer0_outputs(2283) <= not((inputs(161)) and (inputs(207)));
    layer0_outputs(2284) <= (inputs(234)) and not (inputs(16));
    layer0_outputs(2285) <= (inputs(195)) xor (inputs(207));
    layer0_outputs(2286) <= not((inputs(223)) or (inputs(237)));
    layer0_outputs(2287) <= '1';
    layer0_outputs(2288) <= (inputs(61)) and not (inputs(212));
    layer0_outputs(2289) <= (inputs(22)) xor (inputs(197));
    layer0_outputs(2290) <= (inputs(37)) xor (inputs(131));
    layer0_outputs(2291) <= not(inputs(232));
    layer0_outputs(2292) <= not(inputs(182));
    layer0_outputs(2293) <= not(inputs(240));
    layer0_outputs(2294) <= not(inputs(42)) or (inputs(238));
    layer0_outputs(2295) <= not(inputs(202)) or (inputs(255));
    layer0_outputs(2296) <= not((inputs(205)) xor (inputs(132)));
    layer0_outputs(2297) <= not((inputs(231)) and (inputs(76)));
    layer0_outputs(2298) <= not(inputs(97));
    layer0_outputs(2299) <= not(inputs(242)) or (inputs(133));
    layer0_outputs(2300) <= (inputs(85)) and not (inputs(247));
    layer0_outputs(2301) <= not((inputs(166)) or (inputs(4)));
    layer0_outputs(2302) <= (inputs(100)) and not (inputs(179));
    layer0_outputs(2303) <= (inputs(232)) or (inputs(116));
    layer0_outputs(2304) <= (inputs(12)) and not (inputs(127));
    layer0_outputs(2305) <= '0';
    layer0_outputs(2306) <= not(inputs(55));
    layer0_outputs(2307) <= (inputs(57)) and (inputs(231));
    layer0_outputs(2308) <= not((inputs(36)) xor (inputs(27)));
    layer0_outputs(2309) <= inputs(121);
    layer0_outputs(2310) <= not(inputs(57));
    layer0_outputs(2311) <= (inputs(7)) xor (inputs(226));
    layer0_outputs(2312) <= not(inputs(77)) or (inputs(168));
    layer0_outputs(2313) <= (inputs(66)) or (inputs(185));
    layer0_outputs(2314) <= (inputs(73)) xor (inputs(160));
    layer0_outputs(2315) <= (inputs(44)) or (inputs(120));
    layer0_outputs(2316) <= not((inputs(31)) or (inputs(139)));
    layer0_outputs(2317) <= (inputs(174)) or (inputs(32));
    layer0_outputs(2318) <= (inputs(202)) xor (inputs(104));
    layer0_outputs(2319) <= not((inputs(251)) xor (inputs(80)));
    layer0_outputs(2320) <= not(inputs(170)) or (inputs(5));
    layer0_outputs(2321) <= not((inputs(49)) xor (inputs(31)));
    layer0_outputs(2322) <= '1';
    layer0_outputs(2323) <= (inputs(113)) xor (inputs(132));
    layer0_outputs(2324) <= not(inputs(133));
    layer0_outputs(2325) <= not(inputs(42));
    layer0_outputs(2326) <= not(inputs(63)) or (inputs(242));
    layer0_outputs(2327) <= not(inputs(7));
    layer0_outputs(2328) <= not(inputs(167));
    layer0_outputs(2329) <= (inputs(107)) and not (inputs(110));
    layer0_outputs(2330) <= (inputs(186)) and (inputs(143));
    layer0_outputs(2331) <= not(inputs(193)) or (inputs(174));
    layer0_outputs(2332) <= (inputs(228)) and (inputs(79));
    layer0_outputs(2333) <= (inputs(248)) and not (inputs(180));
    layer0_outputs(2334) <= not(inputs(84)) or (inputs(126));
    layer0_outputs(2335) <= '1';
    layer0_outputs(2336) <= inputs(169);
    layer0_outputs(2337) <= not((inputs(141)) xor (inputs(106)));
    layer0_outputs(2338) <= (inputs(72)) and not (inputs(158));
    layer0_outputs(2339) <= '1';
    layer0_outputs(2340) <= (inputs(187)) or (inputs(164));
    layer0_outputs(2341) <= not(inputs(8));
    layer0_outputs(2342) <= (inputs(191)) xor (inputs(255));
    layer0_outputs(2343) <= (inputs(104)) xor (inputs(204));
    layer0_outputs(2344) <= inputs(234);
    layer0_outputs(2345) <= (inputs(98)) and not (inputs(217));
    layer0_outputs(2346) <= (inputs(68)) and not (inputs(115));
    layer0_outputs(2347) <= not((inputs(253)) or (inputs(211)));
    layer0_outputs(2348) <= (inputs(53)) xor (inputs(13));
    layer0_outputs(2349) <= (inputs(63)) or (inputs(250));
    layer0_outputs(2350) <= inputs(57);
    layer0_outputs(2351) <= (inputs(132)) and not (inputs(143));
    layer0_outputs(2352) <= not(inputs(150)) or (inputs(27));
    layer0_outputs(2353) <= inputs(13);
    layer0_outputs(2354) <= (inputs(237)) and not (inputs(255));
    layer0_outputs(2355) <= (inputs(65)) and not (inputs(242));
    layer0_outputs(2356) <= not((inputs(215)) xor (inputs(183)));
    layer0_outputs(2357) <= (inputs(204)) xor (inputs(222));
    layer0_outputs(2358) <= (inputs(124)) and (inputs(41));
    layer0_outputs(2359) <= (inputs(242)) or (inputs(110));
    layer0_outputs(2360) <= (inputs(81)) xor (inputs(50));
    layer0_outputs(2361) <= (inputs(252)) and (inputs(95));
    layer0_outputs(2362) <= (inputs(42)) and not (inputs(233));
    layer0_outputs(2363) <= '1';
    layer0_outputs(2364) <= (inputs(206)) xor (inputs(252));
    layer0_outputs(2365) <= not((inputs(130)) xor (inputs(80)));
    layer0_outputs(2366) <= (inputs(124)) xor (inputs(113));
    layer0_outputs(2367) <= (inputs(9)) and not (inputs(175));
    layer0_outputs(2368) <= not(inputs(45)) or (inputs(176));
    layer0_outputs(2369) <= inputs(25);
    layer0_outputs(2370) <= (inputs(153)) xor (inputs(58));
    layer0_outputs(2371) <= not((inputs(197)) xor (inputs(155)));
    layer0_outputs(2372) <= not(inputs(71));
    layer0_outputs(2373) <= inputs(99);
    layer0_outputs(2374) <= not(inputs(8)) or (inputs(132));
    layer0_outputs(2375) <= inputs(148);
    layer0_outputs(2376) <= not(inputs(145)) or (inputs(12));
    layer0_outputs(2377) <= (inputs(242)) or (inputs(16));
    layer0_outputs(2378) <= (inputs(62)) or (inputs(67));
    layer0_outputs(2379) <= (inputs(162)) or (inputs(160));
    layer0_outputs(2380) <= not(inputs(175));
    layer0_outputs(2381) <= not((inputs(35)) xor (inputs(143)));
    layer0_outputs(2382) <= inputs(195);
    layer0_outputs(2383) <= not(inputs(75)) or (inputs(15));
    layer0_outputs(2384) <= (inputs(11)) and not (inputs(203));
    layer0_outputs(2385) <= not((inputs(113)) or (inputs(216)));
    layer0_outputs(2386) <= (inputs(135)) and not (inputs(3));
    layer0_outputs(2387) <= not(inputs(212)) or (inputs(207));
    layer0_outputs(2388) <= not((inputs(253)) or (inputs(5)));
    layer0_outputs(2389) <= inputs(102);
    layer0_outputs(2390) <= not(inputs(233));
    layer0_outputs(2391) <= not(inputs(195));
    layer0_outputs(2392) <= (inputs(248)) and (inputs(181));
    layer0_outputs(2393) <= (inputs(41)) xor (inputs(158));
    layer0_outputs(2394) <= not(inputs(143)) or (inputs(38));
    layer0_outputs(2395) <= inputs(137);
    layer0_outputs(2396) <= not((inputs(241)) or (inputs(9)));
    layer0_outputs(2397) <= not((inputs(75)) or (inputs(19)));
    layer0_outputs(2398) <= (inputs(89)) and not (inputs(63));
    layer0_outputs(2399) <= not(inputs(94));
    layer0_outputs(2400) <= (inputs(223)) xor (inputs(191));
    layer0_outputs(2401) <= not(inputs(236));
    layer0_outputs(2402) <= inputs(55);
    layer0_outputs(2403) <= not((inputs(159)) or (inputs(194)));
    layer0_outputs(2404) <= (inputs(90)) or (inputs(49));
    layer0_outputs(2405) <= '1';
    layer0_outputs(2406) <= (inputs(217)) and not (inputs(255));
    layer0_outputs(2407) <= not(inputs(189)) or (inputs(108));
    layer0_outputs(2408) <= inputs(4);
    layer0_outputs(2409) <= not(inputs(99));
    layer0_outputs(2410) <= (inputs(96)) or (inputs(250));
    layer0_outputs(2411) <= (inputs(27)) and not (inputs(161));
    layer0_outputs(2412) <= inputs(68);
    layer0_outputs(2413) <= (inputs(66)) xor (inputs(67));
    layer0_outputs(2414) <= not((inputs(65)) xor (inputs(62)));
    layer0_outputs(2415) <= not(inputs(214));
    layer0_outputs(2416) <= not((inputs(200)) or (inputs(143)));
    layer0_outputs(2417) <= (inputs(212)) xor (inputs(243));
    layer0_outputs(2418) <= (inputs(111)) and not (inputs(191));
    layer0_outputs(2419) <= (inputs(145)) or (inputs(189));
    layer0_outputs(2420) <= '1';
    layer0_outputs(2421) <= not((inputs(210)) and (inputs(99)));
    layer0_outputs(2422) <= not(inputs(131)) or (inputs(53));
    layer0_outputs(2423) <= (inputs(85)) and not (inputs(88));
    layer0_outputs(2424) <= not(inputs(152));
    layer0_outputs(2425) <= not(inputs(116)) or (inputs(71));
    layer0_outputs(2426) <= (inputs(118)) or (inputs(10));
    layer0_outputs(2427) <= inputs(9);
    layer0_outputs(2428) <= not(inputs(73));
    layer0_outputs(2429) <= not(inputs(105));
    layer0_outputs(2430) <= not(inputs(36));
    layer0_outputs(2431) <= not((inputs(10)) xor (inputs(1)));
    layer0_outputs(2432) <= not(inputs(7));
    layer0_outputs(2433) <= not(inputs(89)) or (inputs(19));
    layer0_outputs(2434) <= (inputs(76)) and not (inputs(14));
    layer0_outputs(2435) <= (inputs(87)) xor (inputs(177));
    layer0_outputs(2436) <= not((inputs(68)) xor (inputs(133)));
    layer0_outputs(2437) <= inputs(78);
    layer0_outputs(2438) <= not(inputs(158)) or (inputs(183));
    layer0_outputs(2439) <= (inputs(187)) xor (inputs(236));
    layer0_outputs(2440) <= not(inputs(83)) or (inputs(78));
    layer0_outputs(2441) <= not((inputs(121)) xor (inputs(16)));
    layer0_outputs(2442) <= '0';
    layer0_outputs(2443) <= not(inputs(138)) or (inputs(137));
    layer0_outputs(2444) <= inputs(194);
    layer0_outputs(2445) <= (inputs(252)) or (inputs(239));
    layer0_outputs(2446) <= not((inputs(222)) and (inputs(17)));
    layer0_outputs(2447) <= not((inputs(143)) xor (inputs(79)));
    layer0_outputs(2448) <= not(inputs(212)) or (inputs(124));
    layer0_outputs(2449) <= not((inputs(68)) or (inputs(18)));
    layer0_outputs(2450) <= not(inputs(164)) or (inputs(47));
    layer0_outputs(2451) <= not(inputs(185));
    layer0_outputs(2452) <= not(inputs(212));
    layer0_outputs(2453) <= inputs(86);
    layer0_outputs(2454) <= not((inputs(217)) or (inputs(172)));
    layer0_outputs(2455) <= (inputs(157)) or (inputs(160));
    layer0_outputs(2456) <= not((inputs(15)) xor (inputs(172)));
    layer0_outputs(2457) <= not((inputs(112)) or (inputs(69)));
    layer0_outputs(2458) <= not(inputs(250)) or (inputs(60));
    layer0_outputs(2459) <= inputs(18);
    layer0_outputs(2460) <= (inputs(55)) xor (inputs(88));
    layer0_outputs(2461) <= (inputs(2)) or (inputs(142));
    layer0_outputs(2462) <= inputs(103);
    layer0_outputs(2463) <= not(inputs(106));
    layer0_outputs(2464) <= not(inputs(133)) or (inputs(50));
    layer0_outputs(2465) <= (inputs(250)) and not (inputs(62));
    layer0_outputs(2466) <= (inputs(206)) xor (inputs(109));
    layer0_outputs(2467) <= not((inputs(148)) or (inputs(85)));
    layer0_outputs(2468) <= (inputs(133)) xor (inputs(180));
    layer0_outputs(2469) <= (inputs(194)) and not (inputs(15));
    layer0_outputs(2470) <= not(inputs(23)) or (inputs(214));
    layer0_outputs(2471) <= not(inputs(8)) or (inputs(240));
    layer0_outputs(2472) <= (inputs(88)) and not (inputs(225));
    layer0_outputs(2473) <= (inputs(144)) or (inputs(211));
    layer0_outputs(2474) <= inputs(69);
    layer0_outputs(2475) <= not(inputs(45));
    layer0_outputs(2476) <= '1';
    layer0_outputs(2477) <= (inputs(208)) and not (inputs(244));
    layer0_outputs(2478) <= inputs(21);
    layer0_outputs(2479) <= (inputs(49)) or (inputs(225));
    layer0_outputs(2480) <= inputs(227);
    layer0_outputs(2481) <= not((inputs(27)) or (inputs(216)));
    layer0_outputs(2482) <= not(inputs(51)) or (inputs(137));
    layer0_outputs(2483) <= not(inputs(226)) or (inputs(52));
    layer0_outputs(2484) <= (inputs(126)) or (inputs(160));
    layer0_outputs(2485) <= inputs(145);
    layer0_outputs(2486) <= not(inputs(21)) or (inputs(13));
    layer0_outputs(2487) <= inputs(74);
    layer0_outputs(2488) <= inputs(5);
    layer0_outputs(2489) <= not(inputs(59));
    layer0_outputs(2490) <= not((inputs(77)) and (inputs(71)));
    layer0_outputs(2491) <= not(inputs(62));
    layer0_outputs(2492) <= not(inputs(101)) or (inputs(64));
    layer0_outputs(2493) <= not((inputs(72)) or (inputs(159)));
    layer0_outputs(2494) <= not(inputs(166));
    layer0_outputs(2495) <= inputs(159);
    layer0_outputs(2496) <= not(inputs(149));
    layer0_outputs(2497) <= (inputs(104)) and not (inputs(130));
    layer0_outputs(2498) <= not(inputs(74)) or (inputs(145));
    layer0_outputs(2499) <= (inputs(128)) and not (inputs(125));
    layer0_outputs(2500) <= not(inputs(136));
    layer0_outputs(2501) <= (inputs(77)) and not (inputs(127));
    layer0_outputs(2502) <= not(inputs(97));
    layer0_outputs(2503) <= inputs(62);
    layer0_outputs(2504) <= not((inputs(249)) or (inputs(248)));
    layer0_outputs(2505) <= not(inputs(7));
    layer0_outputs(2506) <= (inputs(190)) xor (inputs(149));
    layer0_outputs(2507) <= inputs(130);
    layer0_outputs(2508) <= not(inputs(115)) or (inputs(215));
    layer0_outputs(2509) <= not((inputs(1)) xor (inputs(207)));
    layer0_outputs(2510) <= (inputs(25)) and not (inputs(206));
    layer0_outputs(2511) <= not((inputs(185)) or (inputs(140)));
    layer0_outputs(2512) <= not(inputs(211)) or (inputs(49));
    layer0_outputs(2513) <= not(inputs(103));
    layer0_outputs(2514) <= not((inputs(17)) or (inputs(195)));
    layer0_outputs(2515) <= inputs(85);
    layer0_outputs(2516) <= inputs(165);
    layer0_outputs(2517) <= inputs(163);
    layer0_outputs(2518) <= not((inputs(129)) xor (inputs(95)));
    layer0_outputs(2519) <= (inputs(55)) and not (inputs(86));
    layer0_outputs(2520) <= (inputs(205)) or (inputs(90));
    layer0_outputs(2521) <= (inputs(27)) xor (inputs(122));
    layer0_outputs(2522) <= not((inputs(79)) or (inputs(94)));
    layer0_outputs(2523) <= (inputs(59)) and not (inputs(86));
    layer0_outputs(2524) <= not((inputs(124)) xor (inputs(122)));
    layer0_outputs(2525) <= (inputs(173)) xor (inputs(88));
    layer0_outputs(2526) <= not(inputs(184)) or (inputs(175));
    layer0_outputs(2527) <= (inputs(205)) xor (inputs(125));
    layer0_outputs(2528) <= not(inputs(182)) or (inputs(17));
    layer0_outputs(2529) <= not(inputs(202)) or (inputs(68));
    layer0_outputs(2530) <= not((inputs(16)) or (inputs(54)));
    layer0_outputs(2531) <= (inputs(193)) and not (inputs(143));
    layer0_outputs(2532) <= (inputs(207)) and not (inputs(52));
    layer0_outputs(2533) <= not(inputs(114)) or (inputs(191));
    layer0_outputs(2534) <= inputs(103);
    layer0_outputs(2535) <= inputs(29);
    layer0_outputs(2536) <= not(inputs(100));
    layer0_outputs(2537) <= (inputs(93)) xor (inputs(91));
    layer0_outputs(2538) <= not(inputs(183)) or (inputs(52));
    layer0_outputs(2539) <= not((inputs(21)) xor (inputs(69)));
    layer0_outputs(2540) <= (inputs(162)) or (inputs(214));
    layer0_outputs(2541) <= not(inputs(68));
    layer0_outputs(2542) <= not((inputs(145)) xor (inputs(87)));
    layer0_outputs(2543) <= not((inputs(18)) or (inputs(213)));
    layer0_outputs(2544) <= (inputs(14)) or (inputs(79));
    layer0_outputs(2545) <= '1';
    layer0_outputs(2546) <= (inputs(32)) or (inputs(113));
    layer0_outputs(2547) <= not(inputs(223));
    layer0_outputs(2548) <= not(inputs(102));
    layer0_outputs(2549) <= (inputs(245)) or (inputs(55));
    layer0_outputs(2550) <= not(inputs(43)) or (inputs(2));
    layer0_outputs(2551) <= not((inputs(166)) or (inputs(122)));
    layer0_outputs(2552) <= not(inputs(104));
    layer0_outputs(2553) <= not(inputs(73));
    layer0_outputs(2554) <= not(inputs(221)) or (inputs(3));
    layer0_outputs(2555) <= inputs(72);
    layer0_outputs(2556) <= (inputs(77)) xor (inputs(232));
    layer0_outputs(2557) <= (inputs(223)) xor (inputs(49));
    layer0_outputs(2558) <= not((inputs(8)) or (inputs(161)));
    layer0_outputs(2559) <= not((inputs(12)) or (inputs(89)));
    layer0_outputs(2560) <= (inputs(187)) xor (inputs(146));
    layer0_outputs(2561) <= not(inputs(168));
    layer0_outputs(2562) <= (inputs(98)) xor (inputs(235));
    layer0_outputs(2563) <= not(inputs(238)) or (inputs(198));
    layer0_outputs(2564) <= (inputs(31)) xor (inputs(122));
    layer0_outputs(2565) <= (inputs(95)) xor (inputs(108));
    layer0_outputs(2566) <= (inputs(48)) or (inputs(111));
    layer0_outputs(2567) <= (inputs(155)) xor (inputs(108));
    layer0_outputs(2568) <= not(inputs(60)) or (inputs(37));
    layer0_outputs(2569) <= inputs(72);
    layer0_outputs(2570) <= inputs(16);
    layer0_outputs(2571) <= inputs(234);
    layer0_outputs(2572) <= (inputs(229)) and not (inputs(76));
    layer0_outputs(2573) <= inputs(18);
    layer0_outputs(2574) <= inputs(148);
    layer0_outputs(2575) <= inputs(83);
    layer0_outputs(2576) <= inputs(104);
    layer0_outputs(2577) <= (inputs(111)) or (inputs(162));
    layer0_outputs(2578) <= not((inputs(91)) xor (inputs(138)));
    layer0_outputs(2579) <= not((inputs(202)) or (inputs(0)));
    layer0_outputs(2580) <= not(inputs(100)) or (inputs(158));
    layer0_outputs(2581) <= (inputs(175)) or (inputs(190));
    layer0_outputs(2582) <= inputs(3);
    layer0_outputs(2583) <= not(inputs(247)) or (inputs(15));
    layer0_outputs(2584) <= inputs(97);
    layer0_outputs(2585) <= not(inputs(3));
    layer0_outputs(2586) <= not((inputs(206)) xor (inputs(238)));
    layer0_outputs(2587) <= not((inputs(55)) or (inputs(185)));
    layer0_outputs(2588) <= inputs(212);
    layer0_outputs(2589) <= not(inputs(164));
    layer0_outputs(2590) <= (inputs(6)) and not (inputs(247));
    layer0_outputs(2591) <= (inputs(125)) or (inputs(71));
    layer0_outputs(2592) <= not(inputs(155));
    layer0_outputs(2593) <= inputs(60);
    layer0_outputs(2594) <= not(inputs(119)) or (inputs(97));
    layer0_outputs(2595) <= (inputs(174)) and (inputs(202));
    layer0_outputs(2596) <= not(inputs(202)) or (inputs(220));
    layer0_outputs(2597) <= not((inputs(53)) xor (inputs(253)));
    layer0_outputs(2598) <= not(inputs(66));
    layer0_outputs(2599) <= (inputs(246)) and not (inputs(166));
    layer0_outputs(2600) <= inputs(189);
    layer0_outputs(2601) <= (inputs(57)) and not (inputs(13));
    layer0_outputs(2602) <= not(inputs(163));
    layer0_outputs(2603) <= inputs(226);
    layer0_outputs(2604) <= not((inputs(205)) or (inputs(155)));
    layer0_outputs(2605) <= not((inputs(81)) or (inputs(176)));
    layer0_outputs(2606) <= (inputs(169)) xor (inputs(0));
    layer0_outputs(2607) <= (inputs(33)) xor (inputs(121));
    layer0_outputs(2608) <= not(inputs(121));
    layer0_outputs(2609) <= inputs(26);
    layer0_outputs(2610) <= (inputs(190)) and not (inputs(2));
    layer0_outputs(2611) <= inputs(125);
    layer0_outputs(2612) <= not((inputs(201)) xor (inputs(157)));
    layer0_outputs(2613) <= not((inputs(184)) or (inputs(36)));
    layer0_outputs(2614) <= '1';
    layer0_outputs(2615) <= inputs(101);
    layer0_outputs(2616) <= (inputs(243)) xor (inputs(242));
    layer0_outputs(2617) <= not((inputs(215)) xor (inputs(228)));
    layer0_outputs(2618) <= inputs(218);
    layer0_outputs(2619) <= not(inputs(156));
    layer0_outputs(2620) <= not(inputs(148));
    layer0_outputs(2621) <= (inputs(6)) or (inputs(101));
    layer0_outputs(2622) <= not((inputs(237)) xor (inputs(138)));
    layer0_outputs(2623) <= not(inputs(34)) or (inputs(228));
    layer0_outputs(2624) <= not((inputs(136)) and (inputs(119)));
    layer0_outputs(2625) <= not((inputs(78)) or (inputs(228)));
    layer0_outputs(2626) <= not(inputs(242));
    layer0_outputs(2627) <= inputs(166);
    layer0_outputs(2628) <= not(inputs(123)) or (inputs(103));
    layer0_outputs(2629) <= (inputs(77)) or (inputs(76));
    layer0_outputs(2630) <= not(inputs(213)) or (inputs(43));
    layer0_outputs(2631) <= (inputs(186)) xor (inputs(1));
    layer0_outputs(2632) <= not(inputs(213)) or (inputs(0));
    layer0_outputs(2633) <= (inputs(7)) and not (inputs(253));
    layer0_outputs(2634) <= not(inputs(142));
    layer0_outputs(2635) <= not(inputs(80));
    layer0_outputs(2636) <= not((inputs(65)) xor (inputs(19)));
    layer0_outputs(2637) <= '0';
    layer0_outputs(2638) <= inputs(183);
    layer0_outputs(2639) <= (inputs(210)) and (inputs(77));
    layer0_outputs(2640) <= (inputs(60)) or (inputs(36));
    layer0_outputs(2641) <= (inputs(186)) and not (inputs(30));
    layer0_outputs(2642) <= not(inputs(252)) or (inputs(81));
    layer0_outputs(2643) <= inputs(242);
    layer0_outputs(2644) <= inputs(83);
    layer0_outputs(2645) <= not(inputs(152)) or (inputs(7));
    layer0_outputs(2646) <= inputs(70);
    layer0_outputs(2647) <= not(inputs(9));
    layer0_outputs(2648) <= (inputs(248)) xor (inputs(192));
    layer0_outputs(2649) <= not(inputs(194));
    layer0_outputs(2650) <= not(inputs(169)) or (inputs(26));
    layer0_outputs(2651) <= not((inputs(1)) or (inputs(49)));
    layer0_outputs(2652) <= (inputs(156)) and not (inputs(73));
    layer0_outputs(2653) <= not(inputs(81)) or (inputs(167));
    layer0_outputs(2654) <= not(inputs(209)) or (inputs(2));
    layer0_outputs(2655) <= (inputs(215)) and not (inputs(92));
    layer0_outputs(2656) <= (inputs(117)) and not (inputs(166));
    layer0_outputs(2657) <= not((inputs(21)) xor (inputs(11)));
    layer0_outputs(2658) <= not((inputs(214)) or (inputs(209)));
    layer0_outputs(2659) <= '1';
    layer0_outputs(2660) <= (inputs(170)) or (inputs(102));
    layer0_outputs(2661) <= (inputs(122)) and not (inputs(207));
    layer0_outputs(2662) <= not(inputs(38)) or (inputs(146));
    layer0_outputs(2663) <= (inputs(228)) and not (inputs(82));
    layer0_outputs(2664) <= not((inputs(191)) or (inputs(229)));
    layer0_outputs(2665) <= not(inputs(23)) or (inputs(97));
    layer0_outputs(2666) <= (inputs(148)) and not (inputs(96));
    layer0_outputs(2667) <= not((inputs(241)) xor (inputs(150)));
    layer0_outputs(2668) <= inputs(153);
    layer0_outputs(2669) <= '1';
    layer0_outputs(2670) <= not(inputs(142)) or (inputs(94));
    layer0_outputs(2671) <= inputs(164);
    layer0_outputs(2672) <= (inputs(66)) and not (inputs(97));
    layer0_outputs(2673) <= not(inputs(98));
    layer0_outputs(2674) <= (inputs(106)) and not (inputs(12));
    layer0_outputs(2675) <= not((inputs(12)) and (inputs(41)));
    layer0_outputs(2676) <= (inputs(213)) and (inputs(2));
    layer0_outputs(2677) <= not(inputs(105)) or (inputs(63));
    layer0_outputs(2678) <= inputs(107);
    layer0_outputs(2679) <= (inputs(20)) or (inputs(32));
    layer0_outputs(2680) <= not((inputs(118)) or (inputs(255)));
    layer0_outputs(2681) <= (inputs(230)) and not (inputs(90));
    layer0_outputs(2682) <= not(inputs(106));
    layer0_outputs(2683) <= not(inputs(211)) or (inputs(33));
    layer0_outputs(2684) <= not(inputs(211));
    layer0_outputs(2685) <= not(inputs(88)) or (inputs(4));
    layer0_outputs(2686) <= inputs(200);
    layer0_outputs(2687) <= (inputs(187)) and (inputs(93));
    layer0_outputs(2688) <= not(inputs(98)) or (inputs(210));
    layer0_outputs(2689) <= (inputs(213)) or (inputs(129));
    layer0_outputs(2690) <= (inputs(77)) xor (inputs(171));
    layer0_outputs(2691) <= (inputs(179)) or (inputs(187));
    layer0_outputs(2692) <= (inputs(136)) xor (inputs(226));
    layer0_outputs(2693) <= (inputs(48)) or (inputs(44));
    layer0_outputs(2694) <= (inputs(255)) xor (inputs(247));
    layer0_outputs(2695) <= (inputs(90)) and not (inputs(142));
    layer0_outputs(2696) <= (inputs(113)) or (inputs(158));
    layer0_outputs(2697) <= not(inputs(16));
    layer0_outputs(2698) <= not(inputs(125));
    layer0_outputs(2699) <= not(inputs(56));
    layer0_outputs(2700) <= not(inputs(115)) or (inputs(91));
    layer0_outputs(2701) <= inputs(61);
    layer0_outputs(2702) <= inputs(229);
    layer0_outputs(2703) <= (inputs(23)) or (inputs(111));
    layer0_outputs(2704) <= inputs(37);
    layer0_outputs(2705) <= '0';
    layer0_outputs(2706) <= not(inputs(4));
    layer0_outputs(2707) <= not((inputs(180)) and (inputs(207)));
    layer0_outputs(2708) <= (inputs(71)) or (inputs(110));
    layer0_outputs(2709) <= not((inputs(85)) or (inputs(96)));
    layer0_outputs(2710) <= (inputs(24)) and not (inputs(129));
    layer0_outputs(2711) <= not(inputs(119));
    layer0_outputs(2712) <= inputs(52);
    layer0_outputs(2713) <= (inputs(98)) and (inputs(74));
    layer0_outputs(2714) <= not(inputs(102)) or (inputs(203));
    layer0_outputs(2715) <= not((inputs(123)) xor (inputs(247)));
    layer0_outputs(2716) <= (inputs(93)) xor (inputs(6));
    layer0_outputs(2717) <= (inputs(107)) and not (inputs(234));
    layer0_outputs(2718) <= (inputs(241)) and not (inputs(248));
    layer0_outputs(2719) <= inputs(233);
    layer0_outputs(2720) <= not(inputs(146));
    layer0_outputs(2721) <= not((inputs(2)) or (inputs(159)));
    layer0_outputs(2722) <= not((inputs(177)) or (inputs(177)));
    layer0_outputs(2723) <= inputs(102);
    layer0_outputs(2724) <= inputs(222);
    layer0_outputs(2725) <= inputs(179);
    layer0_outputs(2726) <= not(inputs(43));
    layer0_outputs(2727) <= not(inputs(175)) or (inputs(15));
    layer0_outputs(2728) <= not(inputs(228));
    layer0_outputs(2729) <= not((inputs(187)) or (inputs(134)));
    layer0_outputs(2730) <= inputs(124);
    layer0_outputs(2731) <= not(inputs(237)) or (inputs(207));
    layer0_outputs(2732) <= (inputs(245)) and not (inputs(32));
    layer0_outputs(2733) <= (inputs(5)) and not (inputs(240));
    layer0_outputs(2734) <= not(inputs(156));
    layer0_outputs(2735) <= (inputs(71)) and not (inputs(2));
    layer0_outputs(2736) <= not(inputs(166)) or (inputs(250));
    layer0_outputs(2737) <= (inputs(122)) and not (inputs(8));
    layer0_outputs(2738) <= inputs(75);
    layer0_outputs(2739) <= not((inputs(37)) xor (inputs(120)));
    layer0_outputs(2740) <= not((inputs(122)) and (inputs(123)));
    layer0_outputs(2741) <= not(inputs(100));
    layer0_outputs(2742) <= not(inputs(229));
    layer0_outputs(2743) <= not(inputs(101));
    layer0_outputs(2744) <= not(inputs(177));
    layer0_outputs(2745) <= inputs(188);
    layer0_outputs(2746) <= not(inputs(149));
    layer0_outputs(2747) <= not(inputs(201));
    layer0_outputs(2748) <= (inputs(62)) xor (inputs(11));
    layer0_outputs(2749) <= not((inputs(11)) or (inputs(250)));
    layer0_outputs(2750) <= not((inputs(88)) or (inputs(35)));
    layer0_outputs(2751) <= (inputs(106)) and not (inputs(97));
    layer0_outputs(2752) <= not(inputs(90));
    layer0_outputs(2753) <= (inputs(87)) and (inputs(207));
    layer0_outputs(2754) <= inputs(23);
    layer0_outputs(2755) <= not((inputs(188)) xor (inputs(211)));
    layer0_outputs(2756) <= not((inputs(248)) xor (inputs(213)));
    layer0_outputs(2757) <= not((inputs(37)) xor (inputs(213)));
    layer0_outputs(2758) <= (inputs(252)) and (inputs(49));
    layer0_outputs(2759) <= inputs(50);
    layer0_outputs(2760) <= not((inputs(237)) xor (inputs(190)));
    layer0_outputs(2761) <= not(inputs(163));
    layer0_outputs(2762) <= not((inputs(146)) or (inputs(105)));
    layer0_outputs(2763) <= (inputs(146)) and not (inputs(242));
    layer0_outputs(2764) <= not((inputs(130)) or (inputs(82)));
    layer0_outputs(2765) <= (inputs(92)) xor (inputs(27));
    layer0_outputs(2766) <= not(inputs(182));
    layer0_outputs(2767) <= (inputs(19)) or (inputs(157));
    layer0_outputs(2768) <= (inputs(226)) and not (inputs(29));
    layer0_outputs(2769) <= not(inputs(247)) or (inputs(251));
    layer0_outputs(2770) <= not((inputs(77)) or (inputs(150)));
    layer0_outputs(2771) <= inputs(157);
    layer0_outputs(2772) <= not(inputs(111));
    layer0_outputs(2773) <= not((inputs(245)) or (inputs(43)));
    layer0_outputs(2774) <= not((inputs(97)) or (inputs(191)));
    layer0_outputs(2775) <= not((inputs(169)) and (inputs(58)));
    layer0_outputs(2776) <= inputs(89);
    layer0_outputs(2777) <= not((inputs(116)) or (inputs(248)));
    layer0_outputs(2778) <= (inputs(173)) or (inputs(220));
    layer0_outputs(2779) <= inputs(64);
    layer0_outputs(2780) <= not((inputs(117)) xor (inputs(66)));
    layer0_outputs(2781) <= not((inputs(143)) xor (inputs(45)));
    layer0_outputs(2782) <= (inputs(101)) xor (inputs(123));
    layer0_outputs(2783) <= not((inputs(216)) or (inputs(138)));
    layer0_outputs(2784) <= inputs(178);
    layer0_outputs(2785) <= not(inputs(121));
    layer0_outputs(2786) <= not(inputs(181)) or (inputs(0));
    layer0_outputs(2787) <= not((inputs(226)) or (inputs(177)));
    layer0_outputs(2788) <= not((inputs(200)) xor (inputs(252)));
    layer0_outputs(2789) <= not((inputs(253)) or (inputs(160)));
    layer0_outputs(2790) <= (inputs(81)) xor (inputs(33));
    layer0_outputs(2791) <= inputs(189);
    layer0_outputs(2792) <= (inputs(144)) xor (inputs(8));
    layer0_outputs(2793) <= not(inputs(46));
    layer0_outputs(2794) <= not((inputs(136)) xor (inputs(218)));
    layer0_outputs(2795) <= not(inputs(121));
    layer0_outputs(2796) <= (inputs(100)) or (inputs(78));
    layer0_outputs(2797) <= not((inputs(109)) xor (inputs(245)));
    layer0_outputs(2798) <= inputs(194);
    layer0_outputs(2799) <= (inputs(229)) and not (inputs(60));
    layer0_outputs(2800) <= (inputs(240)) and not (inputs(53));
    layer0_outputs(2801) <= not(inputs(58)) or (inputs(234));
    layer0_outputs(2802) <= inputs(193);
    layer0_outputs(2803) <= (inputs(68)) and not (inputs(87));
    layer0_outputs(2804) <= inputs(210);
    layer0_outputs(2805) <= (inputs(154)) xor (inputs(203));
    layer0_outputs(2806) <= not(inputs(38));
    layer0_outputs(2807) <= not(inputs(166));
    layer0_outputs(2808) <= (inputs(109)) xor (inputs(204));
    layer0_outputs(2809) <= not(inputs(58));
    layer0_outputs(2810) <= inputs(194);
    layer0_outputs(2811) <= not(inputs(129));
    layer0_outputs(2812) <= not(inputs(197)) or (inputs(17));
    layer0_outputs(2813) <= not((inputs(156)) or (inputs(84)));
    layer0_outputs(2814) <= not((inputs(164)) or (inputs(237)));
    layer0_outputs(2815) <= inputs(84);
    layer0_outputs(2816) <= not(inputs(106)) or (inputs(172));
    layer0_outputs(2817) <= not(inputs(59));
    layer0_outputs(2818) <= inputs(58);
    layer0_outputs(2819) <= not((inputs(232)) or (inputs(243)));
    layer0_outputs(2820) <= not((inputs(221)) xor (inputs(250)));
    layer0_outputs(2821) <= (inputs(10)) xor (inputs(22));
    layer0_outputs(2822) <= inputs(180);
    layer0_outputs(2823) <= not(inputs(249));
    layer0_outputs(2824) <= not(inputs(210));
    layer0_outputs(2825) <= not(inputs(206));
    layer0_outputs(2826) <= not(inputs(172));
    layer0_outputs(2827) <= inputs(101);
    layer0_outputs(2828) <= (inputs(108)) and not (inputs(144));
    layer0_outputs(2829) <= not(inputs(209));
    layer0_outputs(2830) <= not(inputs(236));
    layer0_outputs(2831) <= '0';
    layer0_outputs(2832) <= not(inputs(230));
    layer0_outputs(2833) <= not(inputs(90));
    layer0_outputs(2834) <= inputs(245);
    layer0_outputs(2835) <= not(inputs(99));
    layer0_outputs(2836) <= not(inputs(87));
    layer0_outputs(2837) <= not(inputs(129));
    layer0_outputs(2838) <= (inputs(128)) and not (inputs(250));
    layer0_outputs(2839) <= not((inputs(28)) xor (inputs(108)));
    layer0_outputs(2840) <= not(inputs(8));
    layer0_outputs(2841) <= (inputs(135)) and not (inputs(127));
    layer0_outputs(2842) <= not((inputs(23)) or (inputs(6)));
    layer0_outputs(2843) <= inputs(101);
    layer0_outputs(2844) <= (inputs(174)) and not (inputs(209));
    layer0_outputs(2845) <= not(inputs(102));
    layer0_outputs(2846) <= inputs(68);
    layer0_outputs(2847) <= (inputs(131)) and not (inputs(51));
    layer0_outputs(2848) <= not((inputs(15)) or (inputs(100)));
    layer0_outputs(2849) <= inputs(228);
    layer0_outputs(2850) <= not(inputs(109)) or (inputs(16));
    layer0_outputs(2851) <= not((inputs(100)) xor (inputs(255)));
    layer0_outputs(2852) <= not(inputs(13)) or (inputs(51));
    layer0_outputs(2853) <= not((inputs(52)) xor (inputs(53)));
    layer0_outputs(2854) <= not((inputs(16)) xor (inputs(134)));
    layer0_outputs(2855) <= inputs(121);
    layer0_outputs(2856) <= inputs(146);
    layer0_outputs(2857) <= (inputs(213)) and not (inputs(131));
    layer0_outputs(2858) <= not((inputs(58)) xor (inputs(77)));
    layer0_outputs(2859) <= (inputs(1)) and not (inputs(13));
    layer0_outputs(2860) <= not((inputs(118)) or (inputs(196)));
    layer0_outputs(2861) <= inputs(255);
    layer0_outputs(2862) <= not((inputs(11)) xor (inputs(97)));
    layer0_outputs(2863) <= (inputs(24)) or (inputs(77));
    layer0_outputs(2864) <= (inputs(188)) xor (inputs(23));
    layer0_outputs(2865) <= inputs(8);
    layer0_outputs(2866) <= not((inputs(158)) or (inputs(153)));
    layer0_outputs(2867) <= not(inputs(70));
    layer0_outputs(2868) <= not((inputs(149)) xor (inputs(5)));
    layer0_outputs(2869) <= not((inputs(176)) and (inputs(57)));
    layer0_outputs(2870) <= (inputs(136)) and not (inputs(26));
    layer0_outputs(2871) <= inputs(111);
    layer0_outputs(2872) <= not((inputs(23)) or (inputs(122)));
    layer0_outputs(2873) <= not((inputs(123)) xor (inputs(130)));
    layer0_outputs(2874) <= (inputs(247)) xor (inputs(46));
    layer0_outputs(2875) <= inputs(164);
    layer0_outputs(2876) <= '0';
    layer0_outputs(2877) <= not(inputs(162));
    layer0_outputs(2878) <= not(inputs(214)) or (inputs(164));
    layer0_outputs(2879) <= (inputs(230)) and not (inputs(231));
    layer0_outputs(2880) <= inputs(117);
    layer0_outputs(2881) <= inputs(142);
    layer0_outputs(2882) <= not((inputs(76)) xor (inputs(141)));
    layer0_outputs(2883) <= (inputs(206)) xor (inputs(89));
    layer0_outputs(2884) <= not(inputs(162));
    layer0_outputs(2885) <= (inputs(126)) and (inputs(242));
    layer0_outputs(2886) <= (inputs(89)) xor (inputs(122));
    layer0_outputs(2887) <= (inputs(193)) xor (inputs(51));
    layer0_outputs(2888) <= not(inputs(130));
    layer0_outputs(2889) <= (inputs(82)) or (inputs(149));
    layer0_outputs(2890) <= not(inputs(89));
    layer0_outputs(2891) <= (inputs(87)) xor (inputs(99));
    layer0_outputs(2892) <= '0';
    layer0_outputs(2893) <= (inputs(100)) and not (inputs(172));
    layer0_outputs(2894) <= not((inputs(80)) or (inputs(156)));
    layer0_outputs(2895) <= not(inputs(180));
    layer0_outputs(2896) <= '1';
    layer0_outputs(2897) <= not(inputs(210));
    layer0_outputs(2898) <= not(inputs(232)) or (inputs(128));
    layer0_outputs(2899) <= '1';
    layer0_outputs(2900) <= not(inputs(96));
    layer0_outputs(2901) <= (inputs(82)) or (inputs(156));
    layer0_outputs(2902) <= (inputs(57)) and (inputs(70));
    layer0_outputs(2903) <= inputs(86);
    layer0_outputs(2904) <= not((inputs(215)) or (inputs(159)));
    layer0_outputs(2905) <= not(inputs(251)) or (inputs(73));
    layer0_outputs(2906) <= not((inputs(70)) or (inputs(119)));
    layer0_outputs(2907) <= not(inputs(229)) or (inputs(89));
    layer0_outputs(2908) <= (inputs(1)) xor (inputs(189));
    layer0_outputs(2909) <= not((inputs(211)) or (inputs(244)));
    layer0_outputs(2910) <= not((inputs(48)) or (inputs(209)));
    layer0_outputs(2911) <= inputs(92);
    layer0_outputs(2912) <= not((inputs(87)) xor (inputs(201)));
    layer0_outputs(2913) <= not((inputs(141)) xor (inputs(27)));
    layer0_outputs(2914) <= not(inputs(92));
    layer0_outputs(2915) <= (inputs(74)) and (inputs(90));
    layer0_outputs(2916) <= not((inputs(178)) or (inputs(190)));
    layer0_outputs(2917) <= (inputs(185)) and not (inputs(230));
    layer0_outputs(2918) <= (inputs(69)) xor (inputs(223));
    layer0_outputs(2919) <= (inputs(92)) and (inputs(133));
    layer0_outputs(2920) <= not(inputs(71)) or (inputs(149));
    layer0_outputs(2921) <= not((inputs(155)) xor (inputs(146)));
    layer0_outputs(2922) <= inputs(229);
    layer0_outputs(2923) <= (inputs(36)) or (inputs(156));
    layer0_outputs(2924) <= (inputs(79)) and not (inputs(94));
    layer0_outputs(2925) <= (inputs(14)) or (inputs(196));
    layer0_outputs(2926) <= not(inputs(113));
    layer0_outputs(2927) <= not((inputs(17)) and (inputs(49)));
    layer0_outputs(2928) <= (inputs(179)) or (inputs(112));
    layer0_outputs(2929) <= (inputs(219)) or (inputs(187));
    layer0_outputs(2930) <= not(inputs(204)) or (inputs(222));
    layer0_outputs(2931) <= not(inputs(138));
    layer0_outputs(2932) <= (inputs(52)) and not (inputs(116));
    layer0_outputs(2933) <= not(inputs(152)) or (inputs(62));
    layer0_outputs(2934) <= inputs(199);
    layer0_outputs(2935) <= '1';
    layer0_outputs(2936) <= not((inputs(170)) or (inputs(92)));
    layer0_outputs(2937) <= (inputs(179)) and not (inputs(66));
    layer0_outputs(2938) <= not((inputs(140)) or (inputs(252)));
    layer0_outputs(2939) <= not(inputs(201));
    layer0_outputs(2940) <= (inputs(216)) or (inputs(205));
    layer0_outputs(2941) <= not(inputs(198));
    layer0_outputs(2942) <= inputs(198);
    layer0_outputs(2943) <= (inputs(218)) or (inputs(168));
    layer0_outputs(2944) <= not(inputs(96));
    layer0_outputs(2945) <= not((inputs(148)) or (inputs(1)));
    layer0_outputs(2946) <= (inputs(41)) xor (inputs(54));
    layer0_outputs(2947) <= not(inputs(255));
    layer0_outputs(2948) <= (inputs(152)) and not (inputs(207));
    layer0_outputs(2949) <= inputs(229);
    layer0_outputs(2950) <= (inputs(155)) or (inputs(46));
    layer0_outputs(2951) <= (inputs(230)) and not (inputs(125));
    layer0_outputs(2952) <= not(inputs(37)) or (inputs(220));
    layer0_outputs(2953) <= (inputs(118)) xor (inputs(134));
    layer0_outputs(2954) <= not((inputs(14)) xor (inputs(225)));
    layer0_outputs(2955) <= not(inputs(103)) or (inputs(209));
    layer0_outputs(2956) <= not(inputs(87));
    layer0_outputs(2957) <= (inputs(108)) xor (inputs(88));
    layer0_outputs(2958) <= not((inputs(111)) or (inputs(1)));
    layer0_outputs(2959) <= not((inputs(72)) xor (inputs(9)));
    layer0_outputs(2960) <= (inputs(6)) and not (inputs(160));
    layer0_outputs(2961) <= not(inputs(159));
    layer0_outputs(2962) <= not((inputs(219)) xor (inputs(108)));
    layer0_outputs(2963) <= not((inputs(2)) or (inputs(247)));
    layer0_outputs(2964) <= not((inputs(210)) or (inputs(97)));
    layer0_outputs(2965) <= not(inputs(140)) or (inputs(226));
    layer0_outputs(2966) <= not((inputs(141)) or (inputs(30)));
    layer0_outputs(2967) <= (inputs(243)) and not (inputs(159));
    layer0_outputs(2968) <= '0';
    layer0_outputs(2969) <= inputs(6);
    layer0_outputs(2970) <= not((inputs(190)) or (inputs(150)));
    layer0_outputs(2971) <= not(inputs(107));
    layer0_outputs(2972) <= not((inputs(221)) or (inputs(88)));
    layer0_outputs(2973) <= not(inputs(11));
    layer0_outputs(2974) <= not((inputs(88)) xor (inputs(173)));
    layer0_outputs(2975) <= not(inputs(82));
    layer0_outputs(2976) <= not((inputs(244)) or (inputs(8)));
    layer0_outputs(2977) <= (inputs(179)) and (inputs(106));
    layer0_outputs(2978) <= not((inputs(38)) xor (inputs(98)));
    layer0_outputs(2979) <= inputs(142);
    layer0_outputs(2980) <= not((inputs(18)) xor (inputs(36)));
    layer0_outputs(2981) <= not(inputs(144));
    layer0_outputs(2982) <= inputs(59);
    layer0_outputs(2983) <= not((inputs(208)) xor (inputs(105)));
    layer0_outputs(2984) <= (inputs(118)) and not (inputs(94));
    layer0_outputs(2985) <= inputs(19);
    layer0_outputs(2986) <= (inputs(90)) and not (inputs(125));
    layer0_outputs(2987) <= not((inputs(222)) or (inputs(24)));
    layer0_outputs(2988) <= not(inputs(166));
    layer0_outputs(2989) <= not(inputs(158)) or (inputs(10));
    layer0_outputs(2990) <= not((inputs(229)) xor (inputs(207)));
    layer0_outputs(2991) <= (inputs(127)) or (inputs(171));
    layer0_outputs(2992) <= not((inputs(188)) xor (inputs(185)));
    layer0_outputs(2993) <= not(inputs(132)) or (inputs(151));
    layer0_outputs(2994) <= not((inputs(6)) or (inputs(45)));
    layer0_outputs(2995) <= not(inputs(248)) or (inputs(223));
    layer0_outputs(2996) <= (inputs(185)) xor (inputs(199));
    layer0_outputs(2997) <= not((inputs(103)) or (inputs(94)));
    layer0_outputs(2998) <= '0';
    layer0_outputs(2999) <= not((inputs(34)) or (inputs(27)));
    layer0_outputs(3000) <= not(inputs(151)) or (inputs(37));
    layer0_outputs(3001) <= not((inputs(189)) xor (inputs(20)));
    layer0_outputs(3002) <= '1';
    layer0_outputs(3003) <= (inputs(67)) xor (inputs(61));
    layer0_outputs(3004) <= not((inputs(64)) and (inputs(184)));
    layer0_outputs(3005) <= not((inputs(49)) and (inputs(62)));
    layer0_outputs(3006) <= (inputs(138)) and (inputs(122));
    layer0_outputs(3007) <= inputs(83);
    layer0_outputs(3008) <= (inputs(235)) and not (inputs(128));
    layer0_outputs(3009) <= not(inputs(10));
    layer0_outputs(3010) <= (inputs(253)) and not (inputs(142));
    layer0_outputs(3011) <= not((inputs(46)) xor (inputs(34)));
    layer0_outputs(3012) <= not(inputs(196));
    layer0_outputs(3013) <= (inputs(72)) or (inputs(148));
    layer0_outputs(3014) <= not(inputs(38)) or (inputs(192));
    layer0_outputs(3015) <= (inputs(244)) xor (inputs(241));
    layer0_outputs(3016) <= inputs(131);
    layer0_outputs(3017) <= (inputs(74)) and not (inputs(156));
    layer0_outputs(3018) <= not((inputs(239)) or (inputs(3)));
    layer0_outputs(3019) <= (inputs(194)) xor (inputs(227));
    layer0_outputs(3020) <= inputs(252);
    layer0_outputs(3021) <= not((inputs(95)) or (inputs(77)));
    layer0_outputs(3022) <= (inputs(95)) and not (inputs(33));
    layer0_outputs(3023) <= inputs(192);
    layer0_outputs(3024) <= (inputs(33)) or (inputs(208));
    layer0_outputs(3025) <= not(inputs(233));
    layer0_outputs(3026) <= (inputs(140)) and not (inputs(188));
    layer0_outputs(3027) <= (inputs(81)) and not (inputs(112));
    layer0_outputs(3028) <= (inputs(202)) and (inputs(180));
    layer0_outputs(3029) <= inputs(48);
    layer0_outputs(3030) <= (inputs(231)) and not (inputs(140));
    layer0_outputs(3031) <= not(inputs(9));
    layer0_outputs(3032) <= (inputs(189)) or (inputs(91));
    layer0_outputs(3033) <= (inputs(84)) and not (inputs(241));
    layer0_outputs(3034) <= not((inputs(243)) or (inputs(246)));
    layer0_outputs(3035) <= (inputs(166)) xor (inputs(167));
    layer0_outputs(3036) <= (inputs(60)) and not (inputs(147));
    layer0_outputs(3037) <= not((inputs(123)) or (inputs(32)));
    layer0_outputs(3038) <= (inputs(68)) or (inputs(14));
    layer0_outputs(3039) <= not(inputs(185));
    layer0_outputs(3040) <= inputs(232);
    layer0_outputs(3041) <= inputs(181);
    layer0_outputs(3042) <= (inputs(228)) xor (inputs(216));
    layer0_outputs(3043) <= not((inputs(83)) and (inputs(89)));
    layer0_outputs(3044) <= (inputs(142)) xor (inputs(7));
    layer0_outputs(3045) <= inputs(120);
    layer0_outputs(3046) <= (inputs(56)) and not (inputs(133));
    layer0_outputs(3047) <= not(inputs(233)) or (inputs(65));
    layer0_outputs(3048) <= not((inputs(74)) or (inputs(63)));
    layer0_outputs(3049) <= (inputs(135)) and not (inputs(57));
    layer0_outputs(3050) <= (inputs(234)) or (inputs(31));
    layer0_outputs(3051) <= not((inputs(183)) xor (inputs(215)));
    layer0_outputs(3052) <= not(inputs(66));
    layer0_outputs(3053) <= inputs(125);
    layer0_outputs(3054) <= inputs(42);
    layer0_outputs(3055) <= (inputs(48)) xor (inputs(186));
    layer0_outputs(3056) <= inputs(29);
    layer0_outputs(3057) <= not(inputs(185));
    layer0_outputs(3058) <= (inputs(178)) or (inputs(34));
    layer0_outputs(3059) <= not((inputs(174)) or (inputs(247)));
    layer0_outputs(3060) <= (inputs(76)) and not (inputs(125));
    layer0_outputs(3061) <= (inputs(218)) and not (inputs(50));
    layer0_outputs(3062) <= inputs(58);
    layer0_outputs(3063) <= (inputs(20)) and not (inputs(173));
    layer0_outputs(3064) <= inputs(170);
    layer0_outputs(3065) <= (inputs(55)) or (inputs(194));
    layer0_outputs(3066) <= inputs(182);
    layer0_outputs(3067) <= inputs(116);
    layer0_outputs(3068) <= (inputs(220)) and not (inputs(32));
    layer0_outputs(3069) <= inputs(105);
    layer0_outputs(3070) <= not(inputs(20)) or (inputs(93));
    layer0_outputs(3071) <= (inputs(255)) or (inputs(187));
    layer0_outputs(3072) <= (inputs(48)) or (inputs(58));
    layer0_outputs(3073) <= not(inputs(158));
    layer0_outputs(3074) <= not((inputs(77)) or (inputs(76)));
    layer0_outputs(3075) <= (inputs(39)) or (inputs(5));
    layer0_outputs(3076) <= not(inputs(174));
    layer0_outputs(3077) <= not(inputs(165));
    layer0_outputs(3078) <= (inputs(194)) and (inputs(192));
    layer0_outputs(3079) <= (inputs(28)) and not (inputs(114));
    layer0_outputs(3080) <= not(inputs(120));
    layer0_outputs(3081) <= (inputs(141)) or (inputs(53));
    layer0_outputs(3082) <= not(inputs(145));
    layer0_outputs(3083) <= not(inputs(117));
    layer0_outputs(3084) <= not(inputs(230));
    layer0_outputs(3085) <= not(inputs(104));
    layer0_outputs(3086) <= (inputs(220)) and (inputs(86));
    layer0_outputs(3087) <= not(inputs(57)) or (inputs(222));
    layer0_outputs(3088) <= (inputs(127)) or (inputs(147));
    layer0_outputs(3089) <= not((inputs(180)) or (inputs(177)));
    layer0_outputs(3090) <= (inputs(217)) xor (inputs(237));
    layer0_outputs(3091) <= inputs(104);
    layer0_outputs(3092) <= not((inputs(16)) or (inputs(168)));
    layer0_outputs(3093) <= (inputs(30)) or (inputs(245));
    layer0_outputs(3094) <= (inputs(238)) and (inputs(61));
    layer0_outputs(3095) <= not((inputs(50)) or (inputs(70)));
    layer0_outputs(3096) <= inputs(136);
    layer0_outputs(3097) <= not((inputs(166)) or (inputs(152)));
    layer0_outputs(3098) <= not((inputs(86)) xor (inputs(19)));
    layer0_outputs(3099) <= (inputs(82)) and not (inputs(125));
    layer0_outputs(3100) <= (inputs(149)) xor (inputs(37));
    layer0_outputs(3101) <= inputs(24);
    layer0_outputs(3102) <= (inputs(118)) and not (inputs(162));
    layer0_outputs(3103) <= (inputs(244)) and not (inputs(26));
    layer0_outputs(3104) <= not((inputs(116)) or (inputs(235)));
    layer0_outputs(3105) <= not(inputs(115)) or (inputs(49));
    layer0_outputs(3106) <= not((inputs(45)) and (inputs(227)));
    layer0_outputs(3107) <= not((inputs(117)) or (inputs(97)));
    layer0_outputs(3108) <= not(inputs(89)) or (inputs(164));
    layer0_outputs(3109) <= inputs(181);
    layer0_outputs(3110) <= (inputs(138)) and not (inputs(173));
    layer0_outputs(3111) <= (inputs(182)) and not (inputs(146));
    layer0_outputs(3112) <= not((inputs(223)) xor (inputs(197)));
    layer0_outputs(3113) <= not((inputs(67)) xor (inputs(86)));
    layer0_outputs(3114) <= (inputs(3)) or (inputs(110));
    layer0_outputs(3115) <= (inputs(176)) or (inputs(13));
    layer0_outputs(3116) <= (inputs(215)) and not (inputs(61));
    layer0_outputs(3117) <= not(inputs(183));
    layer0_outputs(3118) <= inputs(93);
    layer0_outputs(3119) <= (inputs(148)) or (inputs(139));
    layer0_outputs(3120) <= (inputs(214)) and not (inputs(60));
    layer0_outputs(3121) <= not(inputs(106)) or (inputs(117));
    layer0_outputs(3122) <= not((inputs(187)) or (inputs(232)));
    layer0_outputs(3123) <= inputs(173);
    layer0_outputs(3124) <= inputs(147);
    layer0_outputs(3125) <= not(inputs(151));
    layer0_outputs(3126) <= not(inputs(75));
    layer0_outputs(3127) <= not((inputs(10)) xor (inputs(144)));
    layer0_outputs(3128) <= (inputs(14)) or (inputs(134));
    layer0_outputs(3129) <= not((inputs(29)) or (inputs(121)));
    layer0_outputs(3130) <= (inputs(196)) xor (inputs(171));
    layer0_outputs(3131) <= (inputs(13)) or (inputs(85));
    layer0_outputs(3132) <= (inputs(137)) and not (inputs(48));
    layer0_outputs(3133) <= not(inputs(40)) or (inputs(83));
    layer0_outputs(3134) <= inputs(231);
    layer0_outputs(3135) <= (inputs(1)) or (inputs(253));
    layer0_outputs(3136) <= (inputs(143)) and not (inputs(64));
    layer0_outputs(3137) <= not(inputs(22)) or (inputs(166));
    layer0_outputs(3138) <= not((inputs(122)) or (inputs(46)));
    layer0_outputs(3139) <= not(inputs(205));
    layer0_outputs(3140) <= (inputs(116)) and (inputs(42));
    layer0_outputs(3141) <= (inputs(152)) xor (inputs(137));
    layer0_outputs(3142) <= not((inputs(89)) xor (inputs(203)));
    layer0_outputs(3143) <= (inputs(127)) xor (inputs(122));
    layer0_outputs(3144) <= (inputs(30)) xor (inputs(49));
    layer0_outputs(3145) <= not(inputs(52)) or (inputs(250));
    layer0_outputs(3146) <= (inputs(213)) and (inputs(226));
    layer0_outputs(3147) <= not((inputs(23)) or (inputs(188)));
    layer0_outputs(3148) <= not(inputs(102));
    layer0_outputs(3149) <= not(inputs(253));
    layer0_outputs(3150) <= not(inputs(190)) or (inputs(1));
    layer0_outputs(3151) <= not((inputs(65)) xor (inputs(186)));
    layer0_outputs(3152) <= inputs(167);
    layer0_outputs(3153) <= (inputs(115)) xor (inputs(1));
    layer0_outputs(3154) <= not(inputs(184)) or (inputs(17));
    layer0_outputs(3155) <= not(inputs(17));
    layer0_outputs(3156) <= not((inputs(142)) or (inputs(157)));
    layer0_outputs(3157) <= (inputs(138)) and not (inputs(225));
    layer0_outputs(3158) <= inputs(232);
    layer0_outputs(3159) <= not(inputs(132)) or (inputs(138));
    layer0_outputs(3160) <= not((inputs(6)) xor (inputs(174)));
    layer0_outputs(3161) <= not((inputs(127)) or (inputs(111)));
    layer0_outputs(3162) <= (inputs(21)) xor (inputs(81));
    layer0_outputs(3163) <= inputs(89);
    layer0_outputs(3164) <= inputs(151);
    layer0_outputs(3165) <= not(inputs(107)) or (inputs(129));
    layer0_outputs(3166) <= (inputs(29)) and (inputs(213));
    layer0_outputs(3167) <= (inputs(175)) or (inputs(155));
    layer0_outputs(3168) <= (inputs(167)) xor (inputs(25));
    layer0_outputs(3169) <= not((inputs(114)) or (inputs(83)));
    layer0_outputs(3170) <= (inputs(140)) or (inputs(91));
    layer0_outputs(3171) <= (inputs(151)) and not (inputs(35));
    layer0_outputs(3172) <= not(inputs(57)) or (inputs(250));
    layer0_outputs(3173) <= not(inputs(57)) or (inputs(82));
    layer0_outputs(3174) <= (inputs(107)) xor (inputs(60));
    layer0_outputs(3175) <= (inputs(84)) and not (inputs(161));
    layer0_outputs(3176) <= not((inputs(29)) xor (inputs(174)));
    layer0_outputs(3177) <= not((inputs(56)) and (inputs(47)));
    layer0_outputs(3178) <= not(inputs(196));
    layer0_outputs(3179) <= (inputs(96)) xor (inputs(26));
    layer0_outputs(3180) <= not((inputs(209)) or (inputs(247)));
    layer0_outputs(3181) <= not((inputs(159)) and (inputs(47)));
    layer0_outputs(3182) <= (inputs(101)) xor (inputs(182));
    layer0_outputs(3183) <= not((inputs(248)) xor (inputs(21)));
    layer0_outputs(3184) <= not((inputs(247)) and (inputs(171)));
    layer0_outputs(3185) <= '1';
    layer0_outputs(3186) <= inputs(149);
    layer0_outputs(3187) <= inputs(87);
    layer0_outputs(3188) <= inputs(101);
    layer0_outputs(3189) <= inputs(246);
    layer0_outputs(3190) <= not((inputs(109)) or (inputs(90)));
    layer0_outputs(3191) <= not(inputs(83));
    layer0_outputs(3192) <= (inputs(26)) xor (inputs(63));
    layer0_outputs(3193) <= not((inputs(11)) or (inputs(250)));
    layer0_outputs(3194) <= (inputs(76)) xor (inputs(240));
    layer0_outputs(3195) <= not(inputs(119)) or (inputs(6));
    layer0_outputs(3196) <= inputs(231);
    layer0_outputs(3197) <= (inputs(230)) and not (inputs(31));
    layer0_outputs(3198) <= not(inputs(56)) or (inputs(99));
    layer0_outputs(3199) <= not((inputs(82)) xor (inputs(30)));
    layer0_outputs(3200) <= (inputs(247)) and not (inputs(34));
    layer0_outputs(3201) <= not(inputs(252)) or (inputs(158));
    layer0_outputs(3202) <= not((inputs(199)) or (inputs(169)));
    layer0_outputs(3203) <= (inputs(248)) or (inputs(232));
    layer0_outputs(3204) <= not((inputs(106)) or (inputs(63)));
    layer0_outputs(3205) <= not((inputs(253)) or (inputs(114)));
    layer0_outputs(3206) <= (inputs(231)) and not (inputs(27));
    layer0_outputs(3207) <= (inputs(175)) and not (inputs(146));
    layer0_outputs(3208) <= not((inputs(82)) or (inputs(117)));
    layer0_outputs(3209) <= not(inputs(41)) or (inputs(152));
    layer0_outputs(3210) <= not(inputs(22));
    layer0_outputs(3211) <= not(inputs(23)) or (inputs(200));
    layer0_outputs(3212) <= inputs(129);
    layer0_outputs(3213) <= not(inputs(3));
    layer0_outputs(3214) <= inputs(106);
    layer0_outputs(3215) <= (inputs(246)) and not (inputs(5));
    layer0_outputs(3216) <= (inputs(18)) or (inputs(133));
    layer0_outputs(3217) <= (inputs(206)) or (inputs(120));
    layer0_outputs(3218) <= not(inputs(21));
    layer0_outputs(3219) <= inputs(120);
    layer0_outputs(3220) <= not(inputs(120));
    layer0_outputs(3221) <= not(inputs(100)) or (inputs(212));
    layer0_outputs(3222) <= not(inputs(45)) or (inputs(254));
    layer0_outputs(3223) <= (inputs(54)) and not (inputs(117));
    layer0_outputs(3224) <= not((inputs(55)) or (inputs(97)));
    layer0_outputs(3225) <= inputs(146);
    layer0_outputs(3226) <= (inputs(134)) xor (inputs(92));
    layer0_outputs(3227) <= inputs(87);
    layer0_outputs(3228) <= inputs(156);
    layer0_outputs(3229) <= not((inputs(46)) or (inputs(5)));
    layer0_outputs(3230) <= not((inputs(171)) or (inputs(106)));
    layer0_outputs(3231) <= inputs(201);
    layer0_outputs(3232) <= (inputs(247)) xor (inputs(135));
    layer0_outputs(3233) <= not((inputs(205)) or (inputs(9)));
    layer0_outputs(3234) <= '0';
    layer0_outputs(3235) <= not(inputs(184));
    layer0_outputs(3236) <= (inputs(164)) and (inputs(213));
    layer0_outputs(3237) <= not((inputs(153)) xor (inputs(151)));
    layer0_outputs(3238) <= (inputs(252)) or (inputs(65));
    layer0_outputs(3239) <= (inputs(39)) and not (inputs(171));
    layer0_outputs(3240) <= inputs(69);
    layer0_outputs(3241) <= not(inputs(136));
    layer0_outputs(3242) <= not(inputs(82));
    layer0_outputs(3243) <= inputs(130);
    layer0_outputs(3244) <= not(inputs(176)) or (inputs(136));
    layer0_outputs(3245) <= (inputs(36)) xor (inputs(4));
    layer0_outputs(3246) <= (inputs(248)) or (inputs(205));
    layer0_outputs(3247) <= not((inputs(252)) and (inputs(47)));
    layer0_outputs(3248) <= not((inputs(136)) or (inputs(16)));
    layer0_outputs(3249) <= not((inputs(83)) or (inputs(199)));
    layer0_outputs(3250) <= inputs(245);
    layer0_outputs(3251) <= inputs(25);
    layer0_outputs(3252) <= not((inputs(208)) or (inputs(187)));
    layer0_outputs(3253) <= inputs(146);
    layer0_outputs(3254) <= not((inputs(26)) or (inputs(45)));
    layer0_outputs(3255) <= (inputs(4)) xor (inputs(0));
    layer0_outputs(3256) <= (inputs(215)) and not (inputs(113));
    layer0_outputs(3257) <= (inputs(38)) or (inputs(125));
    layer0_outputs(3258) <= not((inputs(47)) or (inputs(52)));
    layer0_outputs(3259) <= (inputs(250)) or (inputs(80));
    layer0_outputs(3260) <= not(inputs(140));
    layer0_outputs(3261) <= (inputs(26)) and not (inputs(21));
    layer0_outputs(3262) <= (inputs(130)) and not (inputs(209));
    layer0_outputs(3263) <= not(inputs(86));
    layer0_outputs(3264) <= inputs(116);
    layer0_outputs(3265) <= not(inputs(160));
    layer0_outputs(3266) <= not((inputs(44)) or (inputs(32)));
    layer0_outputs(3267) <= (inputs(182)) and not (inputs(14));
    layer0_outputs(3268) <= (inputs(5)) xor (inputs(169));
    layer0_outputs(3269) <= not(inputs(47));
    layer0_outputs(3270) <= not(inputs(112));
    layer0_outputs(3271) <= not(inputs(194));
    layer0_outputs(3272) <= not((inputs(58)) xor (inputs(70)));
    layer0_outputs(3273) <= inputs(245);
    layer0_outputs(3274) <= inputs(151);
    layer0_outputs(3275) <= not(inputs(137));
    layer0_outputs(3276) <= not(inputs(177));
    layer0_outputs(3277) <= not(inputs(99));
    layer0_outputs(3278) <= not(inputs(180));
    layer0_outputs(3279) <= not(inputs(37)) or (inputs(65));
    layer0_outputs(3280) <= (inputs(35)) and not (inputs(68));
    layer0_outputs(3281) <= not((inputs(147)) xor (inputs(175)));
    layer0_outputs(3282) <= not(inputs(246)) or (inputs(75));
    layer0_outputs(3283) <= not((inputs(36)) xor (inputs(86)));
    layer0_outputs(3284) <= (inputs(170)) and not (inputs(94));
    layer0_outputs(3285) <= (inputs(61)) and not (inputs(210));
    layer0_outputs(3286) <= inputs(211);
    layer0_outputs(3287) <= inputs(129);
    layer0_outputs(3288) <= (inputs(79)) or (inputs(132));
    layer0_outputs(3289) <= not(inputs(92));
    layer0_outputs(3290) <= not(inputs(152)) or (inputs(83));
    layer0_outputs(3291) <= inputs(246);
    layer0_outputs(3292) <= (inputs(164)) and not (inputs(106));
    layer0_outputs(3293) <= '1';
    layer0_outputs(3294) <= (inputs(31)) or (inputs(76));
    layer0_outputs(3295) <= inputs(182);
    layer0_outputs(3296) <= not(inputs(253)) or (inputs(240));
    layer0_outputs(3297) <= (inputs(137)) or (inputs(52));
    layer0_outputs(3298) <= not(inputs(40)) or (inputs(254));
    layer0_outputs(3299) <= not((inputs(62)) or (inputs(240)));
    layer0_outputs(3300) <= not(inputs(59));
    layer0_outputs(3301) <= not(inputs(201)) or (inputs(156));
    layer0_outputs(3302) <= (inputs(97)) or (inputs(215));
    layer0_outputs(3303) <= not((inputs(20)) xor (inputs(80)));
    layer0_outputs(3304) <= (inputs(17)) xor (inputs(55));
    layer0_outputs(3305) <= not(inputs(68));
    layer0_outputs(3306) <= not((inputs(80)) xor (inputs(211)));
    layer0_outputs(3307) <= not((inputs(236)) or (inputs(13)));
    layer0_outputs(3308) <= (inputs(62)) xor (inputs(75));
    layer0_outputs(3309) <= not((inputs(252)) or (inputs(253)));
    layer0_outputs(3310) <= not(inputs(134));
    layer0_outputs(3311) <= (inputs(250)) or (inputs(75));
    layer0_outputs(3312) <= inputs(194);
    layer0_outputs(3313) <= not((inputs(48)) and (inputs(43)));
    layer0_outputs(3314) <= inputs(118);
    layer0_outputs(3315) <= inputs(42);
    layer0_outputs(3316) <= (inputs(251)) and not (inputs(212));
    layer0_outputs(3317) <= not((inputs(176)) or (inputs(88)));
    layer0_outputs(3318) <= not((inputs(6)) or (inputs(55)));
    layer0_outputs(3319) <= (inputs(133)) xor (inputs(118));
    layer0_outputs(3320) <= (inputs(99)) and not (inputs(2));
    layer0_outputs(3321) <= (inputs(201)) or (inputs(31));
    layer0_outputs(3322) <= not((inputs(61)) xor (inputs(10)));
    layer0_outputs(3323) <= (inputs(97)) or (inputs(7));
    layer0_outputs(3324) <= (inputs(244)) or (inputs(193));
    layer0_outputs(3325) <= not(inputs(7)) or (inputs(160));
    layer0_outputs(3326) <= not(inputs(215));
    layer0_outputs(3327) <= not((inputs(80)) and (inputs(13)));
    layer0_outputs(3328) <= not(inputs(227));
    layer0_outputs(3329) <= (inputs(219)) or (inputs(167));
    layer0_outputs(3330) <= (inputs(251)) and not (inputs(107));
    layer0_outputs(3331) <= not((inputs(220)) or (inputs(235)));
    layer0_outputs(3332) <= (inputs(179)) or (inputs(56));
    layer0_outputs(3333) <= (inputs(95)) xor (inputs(158));
    layer0_outputs(3334) <= not(inputs(224));
    layer0_outputs(3335) <= (inputs(97)) or (inputs(218));
    layer0_outputs(3336) <= (inputs(197)) xor (inputs(119));
    layer0_outputs(3337) <= (inputs(32)) or (inputs(115));
    layer0_outputs(3338) <= not((inputs(88)) or (inputs(57)));
    layer0_outputs(3339) <= inputs(25);
    layer0_outputs(3340) <= (inputs(248)) or (inputs(155));
    layer0_outputs(3341) <= not((inputs(187)) xor (inputs(242)));
    layer0_outputs(3342) <= not(inputs(200));
    layer0_outputs(3343) <= (inputs(232)) xor (inputs(44));
    layer0_outputs(3344) <= not((inputs(110)) or (inputs(85)));
    layer0_outputs(3345) <= (inputs(58)) or (inputs(189));
    layer0_outputs(3346) <= not((inputs(36)) xor (inputs(93)));
    layer0_outputs(3347) <= not(inputs(112)) or (inputs(194));
    layer0_outputs(3348) <= not((inputs(22)) xor (inputs(189)));
    layer0_outputs(3349) <= not(inputs(72)) or (inputs(50));
    layer0_outputs(3350) <= (inputs(152)) and not (inputs(86));
    layer0_outputs(3351) <= (inputs(167)) and not (inputs(211));
    layer0_outputs(3352) <= not(inputs(135)) or (inputs(171));
    layer0_outputs(3353) <= inputs(134);
    layer0_outputs(3354) <= (inputs(244)) or (inputs(225));
    layer0_outputs(3355) <= not((inputs(186)) and (inputs(186)));
    layer0_outputs(3356) <= (inputs(238)) or (inputs(14));
    layer0_outputs(3357) <= (inputs(201)) xor (inputs(255));
    layer0_outputs(3358) <= inputs(253);
    layer0_outputs(3359) <= not((inputs(147)) and (inputs(93)));
    layer0_outputs(3360) <= not((inputs(141)) or (inputs(43)));
    layer0_outputs(3361) <= (inputs(44)) xor (inputs(32));
    layer0_outputs(3362) <= inputs(121);
    layer0_outputs(3363) <= (inputs(224)) and (inputs(239));
    layer0_outputs(3364) <= (inputs(162)) and not (inputs(79));
    layer0_outputs(3365) <= inputs(105);
    layer0_outputs(3366) <= not((inputs(31)) or (inputs(181)));
    layer0_outputs(3367) <= (inputs(228)) or (inputs(194));
    layer0_outputs(3368) <= not(inputs(205));
    layer0_outputs(3369) <= not(inputs(42)) or (inputs(54));
    layer0_outputs(3370) <= (inputs(19)) or (inputs(181));
    layer0_outputs(3371) <= (inputs(135)) xor (inputs(120));
    layer0_outputs(3372) <= not(inputs(37)) or (inputs(40));
    layer0_outputs(3373) <= (inputs(158)) xor (inputs(118));
    layer0_outputs(3374) <= (inputs(20)) or (inputs(22));
    layer0_outputs(3375) <= (inputs(161)) or (inputs(38));
    layer0_outputs(3376) <= not((inputs(63)) or (inputs(37)));
    layer0_outputs(3377) <= (inputs(115)) or (inputs(112));
    layer0_outputs(3378) <= not((inputs(65)) xor (inputs(255)));
    layer0_outputs(3379) <= not(inputs(132));
    layer0_outputs(3380) <= (inputs(197)) and (inputs(221));
    layer0_outputs(3381) <= (inputs(189)) and (inputs(189));
    layer0_outputs(3382) <= not(inputs(77));
    layer0_outputs(3383) <= not(inputs(21)) or (inputs(203));
    layer0_outputs(3384) <= (inputs(146)) xor (inputs(211));
    layer0_outputs(3385) <= not((inputs(128)) or (inputs(196)));
    layer0_outputs(3386) <= not(inputs(123));
    layer0_outputs(3387) <= not(inputs(137)) or (inputs(153));
    layer0_outputs(3388) <= inputs(119);
    layer0_outputs(3389) <= '1';
    layer0_outputs(3390) <= not(inputs(246));
    layer0_outputs(3391) <= inputs(149);
    layer0_outputs(3392) <= not(inputs(248)) or (inputs(73));
    layer0_outputs(3393) <= (inputs(163)) or (inputs(155));
    layer0_outputs(3394) <= inputs(6);
    layer0_outputs(3395) <= (inputs(180)) xor (inputs(130));
    layer0_outputs(3396) <= not((inputs(86)) and (inputs(54)));
    layer0_outputs(3397) <= not(inputs(110));
    layer0_outputs(3398) <= (inputs(69)) or (inputs(98));
    layer0_outputs(3399) <= not((inputs(63)) or (inputs(103)));
    layer0_outputs(3400) <= not(inputs(105)) or (inputs(189));
    layer0_outputs(3401) <= inputs(164);
    layer0_outputs(3402) <= (inputs(182)) or (inputs(159));
    layer0_outputs(3403) <= not(inputs(0)) or (inputs(195));
    layer0_outputs(3404) <= (inputs(154)) or (inputs(238));
    layer0_outputs(3405) <= inputs(165);
    layer0_outputs(3406) <= (inputs(159)) and not (inputs(245));
    layer0_outputs(3407) <= (inputs(216)) or (inputs(114));
    layer0_outputs(3408) <= (inputs(64)) or (inputs(44));
    layer0_outputs(3409) <= (inputs(165)) and not (inputs(207));
    layer0_outputs(3410) <= not(inputs(93));
    layer0_outputs(3411) <= not(inputs(87)) or (inputs(10));
    layer0_outputs(3412) <= not((inputs(125)) or (inputs(84)));
    layer0_outputs(3413) <= (inputs(148)) and not (inputs(233));
    layer0_outputs(3414) <= (inputs(31)) or (inputs(123));
    layer0_outputs(3415) <= (inputs(20)) and not (inputs(82));
    layer0_outputs(3416) <= (inputs(157)) and not (inputs(64));
    layer0_outputs(3417) <= not(inputs(81));
    layer0_outputs(3418) <= not(inputs(231));
    layer0_outputs(3419) <= (inputs(0)) xor (inputs(182));
    layer0_outputs(3420) <= not(inputs(126));
    layer0_outputs(3421) <= inputs(167);
    layer0_outputs(3422) <= (inputs(47)) and not (inputs(54));
    layer0_outputs(3423) <= (inputs(193)) xor (inputs(229));
    layer0_outputs(3424) <= (inputs(215)) or (inputs(169));
    layer0_outputs(3425) <= not((inputs(167)) or (inputs(228)));
    layer0_outputs(3426) <= not(inputs(129)) or (inputs(238));
    layer0_outputs(3427) <= not(inputs(62));
    layer0_outputs(3428) <= not(inputs(108)) or (inputs(158));
    layer0_outputs(3429) <= not((inputs(63)) xor (inputs(67)));
    layer0_outputs(3430) <= (inputs(234)) and not (inputs(82));
    layer0_outputs(3431) <= not(inputs(117)) or (inputs(207));
    layer0_outputs(3432) <= not(inputs(102)) or (inputs(169));
    layer0_outputs(3433) <= not(inputs(21)) or (inputs(183));
    layer0_outputs(3434) <= not((inputs(208)) xor (inputs(235)));
    layer0_outputs(3435) <= (inputs(61)) xor (inputs(150));
    layer0_outputs(3436) <= not((inputs(54)) or (inputs(173)));
    layer0_outputs(3437) <= (inputs(173)) xor (inputs(237));
    layer0_outputs(3438) <= not((inputs(72)) and (inputs(168)));
    layer0_outputs(3439) <= (inputs(101)) and not (inputs(168));
    layer0_outputs(3440) <= inputs(201);
    layer0_outputs(3441) <= not(inputs(166)) or (inputs(155));
    layer0_outputs(3442) <= not(inputs(65)) or (inputs(215));
    layer0_outputs(3443) <= (inputs(89)) or (inputs(225));
    layer0_outputs(3444) <= not((inputs(168)) xor (inputs(188)));
    layer0_outputs(3445) <= '1';
    layer0_outputs(3446) <= not(inputs(28));
    layer0_outputs(3447) <= (inputs(250)) or (inputs(30));
    layer0_outputs(3448) <= not(inputs(89));
    layer0_outputs(3449) <= not((inputs(243)) or (inputs(73)));
    layer0_outputs(3450) <= not((inputs(89)) xor (inputs(26)));
    layer0_outputs(3451) <= not((inputs(74)) or (inputs(88)));
    layer0_outputs(3452) <= (inputs(71)) xor (inputs(21));
    layer0_outputs(3453) <= (inputs(19)) xor (inputs(117));
    layer0_outputs(3454) <= not((inputs(115)) or (inputs(46)));
    layer0_outputs(3455) <= (inputs(107)) or (inputs(15));
    layer0_outputs(3456) <= '1';
    layer0_outputs(3457) <= (inputs(186)) xor (inputs(84));
    layer0_outputs(3458) <= inputs(203);
    layer0_outputs(3459) <= (inputs(214)) xor (inputs(168));
    layer0_outputs(3460) <= '1';
    layer0_outputs(3461) <= inputs(54);
    layer0_outputs(3462) <= (inputs(190)) or (inputs(193));
    layer0_outputs(3463) <= (inputs(78)) xor (inputs(25));
    layer0_outputs(3464) <= (inputs(164)) and not (inputs(115));
    layer0_outputs(3465) <= not((inputs(247)) or (inputs(141)));
    layer0_outputs(3466) <= not((inputs(113)) xor (inputs(186)));
    layer0_outputs(3467) <= (inputs(58)) and not (inputs(177));
    layer0_outputs(3468) <= (inputs(135)) or (inputs(253));
    layer0_outputs(3469) <= not(inputs(249));
    layer0_outputs(3470) <= (inputs(95)) and not (inputs(136));
    layer0_outputs(3471) <= (inputs(195)) or (inputs(224));
    layer0_outputs(3472) <= not((inputs(116)) xor (inputs(244)));
    layer0_outputs(3473) <= not(inputs(132)) or (inputs(15));
    layer0_outputs(3474) <= not((inputs(146)) or (inputs(174)));
    layer0_outputs(3475) <= (inputs(36)) and not (inputs(239));
    layer0_outputs(3476) <= inputs(202);
    layer0_outputs(3477) <= not(inputs(88));
    layer0_outputs(3478) <= not((inputs(202)) or (inputs(25)));
    layer0_outputs(3479) <= (inputs(208)) xor (inputs(82));
    layer0_outputs(3480) <= not(inputs(89)) or (inputs(96));
    layer0_outputs(3481) <= (inputs(163)) or (inputs(107));
    layer0_outputs(3482) <= inputs(58);
    layer0_outputs(3483) <= not(inputs(231));
    layer0_outputs(3484) <= not((inputs(198)) or (inputs(5)));
    layer0_outputs(3485) <= not(inputs(198));
    layer0_outputs(3486) <= (inputs(30)) and not (inputs(122));
    layer0_outputs(3487) <= (inputs(30)) xor (inputs(234));
    layer0_outputs(3488) <= inputs(177);
    layer0_outputs(3489) <= not((inputs(50)) xor (inputs(106)));
    layer0_outputs(3490) <= not(inputs(145));
    layer0_outputs(3491) <= not((inputs(140)) or (inputs(33)));
    layer0_outputs(3492) <= inputs(7);
    layer0_outputs(3493) <= (inputs(120)) or (inputs(172));
    layer0_outputs(3494) <= not((inputs(36)) xor (inputs(254)));
    layer0_outputs(3495) <= inputs(76);
    layer0_outputs(3496) <= inputs(238);
    layer0_outputs(3497) <= (inputs(251)) and not (inputs(145));
    layer0_outputs(3498) <= inputs(28);
    layer0_outputs(3499) <= not((inputs(238)) or (inputs(17)));
    layer0_outputs(3500) <= inputs(97);
    layer0_outputs(3501) <= (inputs(37)) and (inputs(244));
    layer0_outputs(3502) <= (inputs(58)) or (inputs(61));
    layer0_outputs(3503) <= (inputs(124)) xor (inputs(156));
    layer0_outputs(3504) <= not(inputs(245)) or (inputs(223));
    layer0_outputs(3505) <= (inputs(119)) and not (inputs(124));
    layer0_outputs(3506) <= (inputs(192)) or (inputs(235));
    layer0_outputs(3507) <= not((inputs(146)) or (inputs(226)));
    layer0_outputs(3508) <= not((inputs(187)) xor (inputs(120)));
    layer0_outputs(3509) <= (inputs(182)) and not (inputs(101));
    layer0_outputs(3510) <= (inputs(234)) or (inputs(221));
    layer0_outputs(3511) <= not(inputs(56));
    layer0_outputs(3512) <= (inputs(254)) xor (inputs(179));
    layer0_outputs(3513) <= not(inputs(118));
    layer0_outputs(3514) <= (inputs(147)) and not (inputs(160));
    layer0_outputs(3515) <= (inputs(157)) and not (inputs(243));
    layer0_outputs(3516) <= not((inputs(177)) xor (inputs(221)));
    layer0_outputs(3517) <= (inputs(197)) or (inputs(67));
    layer0_outputs(3518) <= inputs(53);
    layer0_outputs(3519) <= not(inputs(9));
    layer0_outputs(3520) <= (inputs(86)) or (inputs(0));
    layer0_outputs(3521) <= not(inputs(84));
    layer0_outputs(3522) <= not(inputs(13)) or (inputs(25));
    layer0_outputs(3523) <= not(inputs(68)) or (inputs(72));
    layer0_outputs(3524) <= not(inputs(131));
    layer0_outputs(3525) <= (inputs(56)) and not (inputs(0));
    layer0_outputs(3526) <= not((inputs(237)) or (inputs(9)));
    layer0_outputs(3527) <= (inputs(244)) or (inputs(46));
    layer0_outputs(3528) <= not((inputs(218)) xor (inputs(187)));
    layer0_outputs(3529) <= not((inputs(20)) xor (inputs(32)));
    layer0_outputs(3530) <= not((inputs(22)) xor (inputs(229)));
    layer0_outputs(3531) <= (inputs(91)) or (inputs(5));
    layer0_outputs(3532) <= inputs(164);
    layer0_outputs(3533) <= not((inputs(192)) or (inputs(242)));
    layer0_outputs(3534) <= (inputs(138)) or (inputs(45));
    layer0_outputs(3535) <= not(inputs(167)) or (inputs(54));
    layer0_outputs(3536) <= (inputs(114)) or (inputs(74));
    layer0_outputs(3537) <= not((inputs(64)) xor (inputs(102)));
    layer0_outputs(3538) <= (inputs(191)) or (inputs(225));
    layer0_outputs(3539) <= (inputs(87)) xor (inputs(208));
    layer0_outputs(3540) <= (inputs(75)) xor (inputs(118));
    layer0_outputs(3541) <= not((inputs(113)) or (inputs(129)));
    layer0_outputs(3542) <= (inputs(0)) or (inputs(92));
    layer0_outputs(3543) <= (inputs(254)) and not (inputs(192));
    layer0_outputs(3544) <= not(inputs(94)) or (inputs(143));
    layer0_outputs(3545) <= (inputs(123)) and not (inputs(191));
    layer0_outputs(3546) <= '0';
    layer0_outputs(3547) <= not((inputs(210)) xor (inputs(255)));
    layer0_outputs(3548) <= inputs(88);
    layer0_outputs(3549) <= not(inputs(232));
    layer0_outputs(3550) <= not(inputs(130));
    layer0_outputs(3551) <= (inputs(36)) xor (inputs(128));
    layer0_outputs(3552) <= inputs(246);
    layer0_outputs(3553) <= not((inputs(235)) or (inputs(250)));
    layer0_outputs(3554) <= not(inputs(41));
    layer0_outputs(3555) <= inputs(97);
    layer0_outputs(3556) <= not((inputs(222)) xor (inputs(249)));
    layer0_outputs(3557) <= inputs(180);
    layer0_outputs(3558) <= not((inputs(71)) xor (inputs(8)));
    layer0_outputs(3559) <= (inputs(166)) or (inputs(167));
    layer0_outputs(3560) <= not(inputs(168));
    layer0_outputs(3561) <= not((inputs(180)) or (inputs(77)));
    layer0_outputs(3562) <= not(inputs(155));
    layer0_outputs(3563) <= (inputs(226)) and not (inputs(48));
    layer0_outputs(3564) <= not(inputs(27));
    layer0_outputs(3565) <= not((inputs(195)) or (inputs(55)));
    layer0_outputs(3566) <= inputs(59);
    layer0_outputs(3567) <= (inputs(38)) and (inputs(234));
    layer0_outputs(3568) <= (inputs(99)) or (inputs(144));
    layer0_outputs(3569) <= not(inputs(36)) or (inputs(31));
    layer0_outputs(3570) <= (inputs(203)) xor (inputs(85));
    layer0_outputs(3571) <= (inputs(102)) or (inputs(17));
    layer0_outputs(3572) <= (inputs(100)) or (inputs(4));
    layer0_outputs(3573) <= (inputs(204)) xor (inputs(124));
    layer0_outputs(3574) <= not(inputs(74)) or (inputs(247));
    layer0_outputs(3575) <= (inputs(242)) and not (inputs(95));
    layer0_outputs(3576) <= inputs(93);
    layer0_outputs(3577) <= not((inputs(76)) or (inputs(80)));
    layer0_outputs(3578) <= (inputs(36)) xor (inputs(54));
    layer0_outputs(3579) <= '1';
    layer0_outputs(3580) <= (inputs(160)) or (inputs(161));
    layer0_outputs(3581) <= not((inputs(94)) xor (inputs(244)));
    layer0_outputs(3582) <= inputs(74);
    layer0_outputs(3583) <= not((inputs(13)) or (inputs(69)));
    layer0_outputs(3584) <= not((inputs(87)) or (inputs(100)));
    layer0_outputs(3585) <= (inputs(141)) xor (inputs(123));
    layer0_outputs(3586) <= (inputs(166)) and not (inputs(12));
    layer0_outputs(3587) <= not(inputs(105));
    layer0_outputs(3588) <= inputs(244);
    layer0_outputs(3589) <= (inputs(241)) xor (inputs(221));
    layer0_outputs(3590) <= not((inputs(24)) xor (inputs(245)));
    layer0_outputs(3591) <= not(inputs(41)) or (inputs(112));
    layer0_outputs(3592) <= (inputs(200)) and (inputs(36));
    layer0_outputs(3593) <= (inputs(104)) and not (inputs(223));
    layer0_outputs(3594) <= not(inputs(237));
    layer0_outputs(3595) <= (inputs(107)) and not (inputs(239));
    layer0_outputs(3596) <= not((inputs(57)) xor (inputs(27)));
    layer0_outputs(3597) <= not(inputs(22));
    layer0_outputs(3598) <= (inputs(24)) or (inputs(30));
    layer0_outputs(3599) <= '0';
    layer0_outputs(3600) <= inputs(60);
    layer0_outputs(3601) <= not((inputs(142)) or (inputs(191)));
    layer0_outputs(3602) <= (inputs(216)) or (inputs(46));
    layer0_outputs(3603) <= not((inputs(152)) xor (inputs(99)));
    layer0_outputs(3604) <= not((inputs(26)) xor (inputs(33)));
    layer0_outputs(3605) <= inputs(37);
    layer0_outputs(3606) <= not(inputs(118));
    layer0_outputs(3607) <= not((inputs(162)) or (inputs(168)));
    layer0_outputs(3608) <= (inputs(151)) and not (inputs(4));
    layer0_outputs(3609) <= (inputs(140)) or (inputs(180));
    layer0_outputs(3610) <= inputs(116);
    layer0_outputs(3611) <= not((inputs(40)) xor (inputs(53)));
    layer0_outputs(3612) <= not(inputs(33));
    layer0_outputs(3613) <= not((inputs(139)) xor (inputs(72)));
    layer0_outputs(3614) <= inputs(101);
    layer0_outputs(3615) <= not(inputs(68)) or (inputs(182));
    layer0_outputs(3616) <= inputs(243);
    layer0_outputs(3617) <= inputs(70);
    layer0_outputs(3618) <= (inputs(185)) and not (inputs(117));
    layer0_outputs(3619) <= not(inputs(136));
    layer0_outputs(3620) <= inputs(181);
    layer0_outputs(3621) <= (inputs(2)) xor (inputs(209));
    layer0_outputs(3622) <= not((inputs(134)) or (inputs(30)));
    layer0_outputs(3623) <= not(inputs(166));
    layer0_outputs(3624) <= not((inputs(191)) or (inputs(220)));
    layer0_outputs(3625) <= not(inputs(98)) or (inputs(177));
    layer0_outputs(3626) <= inputs(219);
    layer0_outputs(3627) <= '0';
    layer0_outputs(3628) <= (inputs(12)) or (inputs(5));
    layer0_outputs(3629) <= not(inputs(131));
    layer0_outputs(3630) <= not((inputs(167)) or (inputs(103)));
    layer0_outputs(3631) <= not((inputs(112)) or (inputs(88)));
    layer0_outputs(3632) <= inputs(193);
    layer0_outputs(3633) <= not(inputs(117));
    layer0_outputs(3634) <= not(inputs(9)) or (inputs(147));
    layer0_outputs(3635) <= not((inputs(205)) xor (inputs(13)));
    layer0_outputs(3636) <= inputs(236);
    layer0_outputs(3637) <= (inputs(44)) xor (inputs(92));
    layer0_outputs(3638) <= not((inputs(242)) or (inputs(172)));
    layer0_outputs(3639) <= (inputs(87)) and not (inputs(112));
    layer0_outputs(3640) <= not((inputs(183)) xor (inputs(99)));
    layer0_outputs(3641) <= not(inputs(132)) or (inputs(243));
    layer0_outputs(3642) <= inputs(147);
    layer0_outputs(3643) <= not(inputs(38));
    layer0_outputs(3644) <= not(inputs(120));
    layer0_outputs(3645) <= (inputs(19)) and not (inputs(209));
    layer0_outputs(3646) <= (inputs(207)) or (inputs(54));
    layer0_outputs(3647) <= not((inputs(237)) xor (inputs(67)));
    layer0_outputs(3648) <= (inputs(182)) or (inputs(151));
    layer0_outputs(3649) <= not(inputs(141)) or (inputs(240));
    layer0_outputs(3650) <= inputs(209);
    layer0_outputs(3651) <= (inputs(141)) and (inputs(239));
    layer0_outputs(3652) <= not(inputs(166)) or (inputs(140));
    layer0_outputs(3653) <= (inputs(121)) and not (inputs(177));
    layer0_outputs(3654) <= not(inputs(219));
    layer0_outputs(3655) <= not((inputs(142)) xor (inputs(4)));
    layer0_outputs(3656) <= (inputs(101)) and not (inputs(218));
    layer0_outputs(3657) <= not((inputs(249)) xor (inputs(135)));
    layer0_outputs(3658) <= (inputs(194)) and not (inputs(251));
    layer0_outputs(3659) <= not((inputs(25)) or (inputs(4)));
    layer0_outputs(3660) <= inputs(85);
    layer0_outputs(3661) <= not(inputs(47)) or (inputs(191));
    layer0_outputs(3662) <= not((inputs(134)) xor (inputs(202)));
    layer0_outputs(3663) <= not((inputs(83)) or (inputs(14)));
    layer0_outputs(3664) <= inputs(50);
    layer0_outputs(3665) <= (inputs(92)) and not (inputs(212));
    layer0_outputs(3666) <= inputs(133);
    layer0_outputs(3667) <= (inputs(20)) or (inputs(17));
    layer0_outputs(3668) <= (inputs(174)) or (inputs(133));
    layer0_outputs(3669) <= not((inputs(171)) xor (inputs(202)));
    layer0_outputs(3670) <= (inputs(144)) or (inputs(74));
    layer0_outputs(3671) <= not((inputs(231)) and (inputs(233)));
    layer0_outputs(3672) <= (inputs(83)) or (inputs(96));
    layer0_outputs(3673) <= (inputs(177)) xor (inputs(240));
    layer0_outputs(3674) <= (inputs(16)) xor (inputs(159));
    layer0_outputs(3675) <= not((inputs(47)) or (inputs(173)));
    layer0_outputs(3676) <= inputs(174);
    layer0_outputs(3677) <= (inputs(178)) and not (inputs(140));
    layer0_outputs(3678) <= (inputs(254)) or (inputs(117));
    layer0_outputs(3679) <= (inputs(48)) or (inputs(18));
    layer0_outputs(3680) <= inputs(110);
    layer0_outputs(3681) <= inputs(158);
    layer0_outputs(3682) <= (inputs(220)) xor (inputs(126));
    layer0_outputs(3683) <= not((inputs(64)) or (inputs(6)));
    layer0_outputs(3684) <= not(inputs(108)) or (inputs(102));
    layer0_outputs(3685) <= inputs(234);
    layer0_outputs(3686) <= (inputs(232)) and not (inputs(40));
    layer0_outputs(3687) <= not((inputs(178)) xor (inputs(208)));
    layer0_outputs(3688) <= not(inputs(213)) or (inputs(88));
    layer0_outputs(3689) <= (inputs(139)) and not (inputs(14));
    layer0_outputs(3690) <= not(inputs(103));
    layer0_outputs(3691) <= inputs(20);
    layer0_outputs(3692) <= not((inputs(191)) xor (inputs(148)));
    layer0_outputs(3693) <= '0';
    layer0_outputs(3694) <= not(inputs(157));
    layer0_outputs(3695) <= (inputs(109)) or (inputs(31));
    layer0_outputs(3696) <= '0';
    layer0_outputs(3697) <= '0';
    layer0_outputs(3698) <= (inputs(75)) or (inputs(125));
    layer0_outputs(3699) <= not(inputs(210));
    layer0_outputs(3700) <= '1';
    layer0_outputs(3701) <= not(inputs(144));
    layer0_outputs(3702) <= (inputs(6)) and not (inputs(174));
    layer0_outputs(3703) <= not(inputs(20));
    layer0_outputs(3704) <= not(inputs(222));
    layer0_outputs(3705) <= inputs(229);
    layer0_outputs(3706) <= inputs(227);
    layer0_outputs(3707) <= inputs(88);
    layer0_outputs(3708) <= (inputs(224)) xor (inputs(158));
    layer0_outputs(3709) <= (inputs(187)) and not (inputs(138));
    layer0_outputs(3710) <= not(inputs(84)) or (inputs(252));
    layer0_outputs(3711) <= (inputs(56)) or (inputs(144));
    layer0_outputs(3712) <= not(inputs(79));
    layer0_outputs(3713) <= (inputs(12)) or (inputs(209));
    layer0_outputs(3714) <= (inputs(160)) and not (inputs(113));
    layer0_outputs(3715) <= (inputs(217)) and not (inputs(134));
    layer0_outputs(3716) <= not(inputs(45));
    layer0_outputs(3717) <= not(inputs(155)) or (inputs(5));
    layer0_outputs(3718) <= (inputs(231)) or (inputs(197));
    layer0_outputs(3719) <= not(inputs(222));
    layer0_outputs(3720) <= not(inputs(29)) or (inputs(146));
    layer0_outputs(3721) <= not(inputs(93));
    layer0_outputs(3722) <= inputs(219);
    layer0_outputs(3723) <= (inputs(137)) or (inputs(105));
    layer0_outputs(3724) <= not((inputs(156)) xor (inputs(192)));
    layer0_outputs(3725) <= not(inputs(79));
    layer0_outputs(3726) <= inputs(214);
    layer0_outputs(3727) <= inputs(43);
    layer0_outputs(3728) <= (inputs(83)) or (inputs(225));
    layer0_outputs(3729) <= not((inputs(61)) xor (inputs(19)));
    layer0_outputs(3730) <= not(inputs(24)) or (inputs(16));
    layer0_outputs(3731) <= not(inputs(71));
    layer0_outputs(3732) <= inputs(89);
    layer0_outputs(3733) <= (inputs(75)) and not (inputs(225));
    layer0_outputs(3734) <= not((inputs(67)) or (inputs(217)));
    layer0_outputs(3735) <= not(inputs(55)) or (inputs(141));
    layer0_outputs(3736) <= inputs(171);
    layer0_outputs(3737) <= not((inputs(35)) or (inputs(228)));
    layer0_outputs(3738) <= not(inputs(85)) or (inputs(216));
    layer0_outputs(3739) <= not(inputs(68)) or (inputs(103));
    layer0_outputs(3740) <= (inputs(139)) and not (inputs(161));
    layer0_outputs(3741) <= (inputs(190)) and not (inputs(254));
    layer0_outputs(3742) <= (inputs(24)) xor (inputs(163));
    layer0_outputs(3743) <= not((inputs(214)) or (inputs(127)));
    layer0_outputs(3744) <= inputs(180);
    layer0_outputs(3745) <= not(inputs(76)) or (inputs(65));
    layer0_outputs(3746) <= not(inputs(123)) or (inputs(111));
    layer0_outputs(3747) <= not(inputs(23));
    layer0_outputs(3748) <= (inputs(171)) and (inputs(160));
    layer0_outputs(3749) <= not(inputs(194));
    layer0_outputs(3750) <= (inputs(38)) or (inputs(94));
    layer0_outputs(3751) <= (inputs(255)) or (inputs(238));
    layer0_outputs(3752) <= not((inputs(84)) or (inputs(32)));
    layer0_outputs(3753) <= not(inputs(90));
    layer0_outputs(3754) <= not(inputs(250));
    layer0_outputs(3755) <= (inputs(63)) xor (inputs(231));
    layer0_outputs(3756) <= not((inputs(20)) or (inputs(55)));
    layer0_outputs(3757) <= (inputs(200)) or (inputs(137));
    layer0_outputs(3758) <= inputs(56);
    layer0_outputs(3759) <= not((inputs(188)) or (inputs(80)));
    layer0_outputs(3760) <= not(inputs(136));
    layer0_outputs(3761) <= not(inputs(49)) or (inputs(246));
    layer0_outputs(3762) <= (inputs(4)) or (inputs(198));
    layer0_outputs(3763) <= (inputs(71)) xor (inputs(134));
    layer0_outputs(3764) <= (inputs(239)) and (inputs(176));
    layer0_outputs(3765) <= inputs(152);
    layer0_outputs(3766) <= not((inputs(201)) or (inputs(4)));
    layer0_outputs(3767) <= inputs(103);
    layer0_outputs(3768) <= (inputs(120)) and not (inputs(125));
    layer0_outputs(3769) <= not((inputs(2)) xor (inputs(178)));
    layer0_outputs(3770) <= not(inputs(118)) or (inputs(212));
    layer0_outputs(3771) <= (inputs(44)) or (inputs(57));
    layer0_outputs(3772) <= (inputs(227)) or (inputs(171));
    layer0_outputs(3773) <= not(inputs(25)) or (inputs(151));
    layer0_outputs(3774) <= not((inputs(247)) and (inputs(153)));
    layer0_outputs(3775) <= (inputs(49)) or (inputs(77));
    layer0_outputs(3776) <= not(inputs(137));
    layer0_outputs(3777) <= (inputs(80)) and not (inputs(47));
    layer0_outputs(3778) <= (inputs(91)) xor (inputs(175));
    layer0_outputs(3779) <= not(inputs(70)) or (inputs(155));
    layer0_outputs(3780) <= not((inputs(228)) xor (inputs(253)));
    layer0_outputs(3781) <= inputs(229);
    layer0_outputs(3782) <= not(inputs(157)) or (inputs(246));
    layer0_outputs(3783) <= (inputs(151)) and not (inputs(26));
    layer0_outputs(3784) <= (inputs(192)) or (inputs(39));
    layer0_outputs(3785) <= (inputs(253)) or (inputs(119));
    layer0_outputs(3786) <= (inputs(73)) xor (inputs(62));
    layer0_outputs(3787) <= not((inputs(226)) or (inputs(219)));
    layer0_outputs(3788) <= not((inputs(6)) or (inputs(2)));
    layer0_outputs(3789) <= not(inputs(194)) or (inputs(92));
    layer0_outputs(3790) <= not((inputs(127)) or (inputs(233)));
    layer0_outputs(3791) <= not((inputs(199)) and (inputs(201)));
    layer0_outputs(3792) <= (inputs(52)) xor (inputs(151));
    layer0_outputs(3793) <= (inputs(204)) and not (inputs(78));
    layer0_outputs(3794) <= not((inputs(222)) xor (inputs(220)));
    layer0_outputs(3795) <= not(inputs(8));
    layer0_outputs(3796) <= not(inputs(89));
    layer0_outputs(3797) <= not((inputs(51)) or (inputs(174)));
    layer0_outputs(3798) <= '0';
    layer0_outputs(3799) <= not(inputs(195));
    layer0_outputs(3800) <= (inputs(183)) and not (inputs(104));
    layer0_outputs(3801) <= (inputs(162)) or (inputs(183));
    layer0_outputs(3802) <= (inputs(191)) xor (inputs(86));
    layer0_outputs(3803) <= not((inputs(146)) xor (inputs(111)));
    layer0_outputs(3804) <= not(inputs(124));
    layer0_outputs(3805) <= inputs(71);
    layer0_outputs(3806) <= not(inputs(37)) or (inputs(219));
    layer0_outputs(3807) <= not(inputs(28));
    layer0_outputs(3808) <= inputs(19);
    layer0_outputs(3809) <= not(inputs(230));
    layer0_outputs(3810) <= not((inputs(102)) or (inputs(103)));
    layer0_outputs(3811) <= not((inputs(201)) xor (inputs(29)));
    layer0_outputs(3812) <= not((inputs(194)) or (inputs(31)));
    layer0_outputs(3813) <= (inputs(120)) xor (inputs(93));
    layer0_outputs(3814) <= not(inputs(152));
    layer0_outputs(3815) <= not((inputs(251)) xor (inputs(84)));
    layer0_outputs(3816) <= (inputs(147)) and not (inputs(119));
    layer0_outputs(3817) <= (inputs(223)) xor (inputs(159));
    layer0_outputs(3818) <= not((inputs(254)) or (inputs(249)));
    layer0_outputs(3819) <= '1';
    layer0_outputs(3820) <= not((inputs(91)) xor (inputs(155)));
    layer0_outputs(3821) <= not((inputs(227)) xor (inputs(28)));
    layer0_outputs(3822) <= not((inputs(13)) or (inputs(169)));
    layer0_outputs(3823) <= not((inputs(130)) or (inputs(156)));
    layer0_outputs(3824) <= inputs(14);
    layer0_outputs(3825) <= (inputs(14)) xor (inputs(87));
    layer0_outputs(3826) <= (inputs(208)) xor (inputs(138));
    layer0_outputs(3827) <= (inputs(69)) or (inputs(98));
    layer0_outputs(3828) <= (inputs(140)) and not (inputs(173));
    layer0_outputs(3829) <= not((inputs(57)) and (inputs(190)));
    layer0_outputs(3830) <= inputs(232);
    layer0_outputs(3831) <= (inputs(227)) or (inputs(128));
    layer0_outputs(3832) <= not(inputs(47));
    layer0_outputs(3833) <= inputs(31);
    layer0_outputs(3834) <= not(inputs(164)) or (inputs(123));
    layer0_outputs(3835) <= not(inputs(27)) or (inputs(254));
    layer0_outputs(3836) <= (inputs(88)) or (inputs(173));
    layer0_outputs(3837) <= '1';
    layer0_outputs(3838) <= not((inputs(68)) xor (inputs(4)));
    layer0_outputs(3839) <= (inputs(152)) xor (inputs(137));
    layer0_outputs(3840) <= not((inputs(129)) or (inputs(198)));
    layer0_outputs(3841) <= inputs(250);
    layer0_outputs(3842) <= not(inputs(233)) or (inputs(206));
    layer0_outputs(3843) <= not(inputs(52)) or (inputs(195));
    layer0_outputs(3844) <= not(inputs(105));
    layer0_outputs(3845) <= not(inputs(88));
    layer0_outputs(3846) <= inputs(248);
    layer0_outputs(3847) <= not((inputs(227)) xor (inputs(161)));
    layer0_outputs(3848) <= (inputs(39)) or (inputs(19));
    layer0_outputs(3849) <= '1';
    layer0_outputs(3850) <= not(inputs(136));
    layer0_outputs(3851) <= inputs(233);
    layer0_outputs(3852) <= not(inputs(116));
    layer0_outputs(3853) <= (inputs(113)) or (inputs(168));
    layer0_outputs(3854) <= (inputs(160)) or (inputs(203));
    layer0_outputs(3855) <= not((inputs(213)) or (inputs(203)));
    layer0_outputs(3856) <= not(inputs(76));
    layer0_outputs(3857) <= (inputs(135)) or (inputs(3));
    layer0_outputs(3858) <= (inputs(29)) xor (inputs(112));
    layer0_outputs(3859) <= not(inputs(181));
    layer0_outputs(3860) <= inputs(106);
    layer0_outputs(3861) <= not((inputs(202)) or (inputs(193)));
    layer0_outputs(3862) <= not(inputs(225));
    layer0_outputs(3863) <= not((inputs(242)) xor (inputs(8)));
    layer0_outputs(3864) <= not(inputs(156)) or (inputs(133));
    layer0_outputs(3865) <= (inputs(71)) xor (inputs(233));
    layer0_outputs(3866) <= inputs(73);
    layer0_outputs(3867) <= inputs(57);
    layer0_outputs(3868) <= not((inputs(252)) xor (inputs(222)));
    layer0_outputs(3869) <= not(inputs(88));
    layer0_outputs(3870) <= (inputs(162)) or (inputs(244));
    layer0_outputs(3871) <= (inputs(135)) or (inputs(134));
    layer0_outputs(3872) <= (inputs(42)) xor (inputs(68));
    layer0_outputs(3873) <= not((inputs(34)) xor (inputs(137)));
    layer0_outputs(3874) <= inputs(55);
    layer0_outputs(3875) <= (inputs(128)) and not (inputs(241));
    layer0_outputs(3876) <= (inputs(60)) xor (inputs(121));
    layer0_outputs(3877) <= not((inputs(215)) or (inputs(221)));
    layer0_outputs(3878) <= (inputs(160)) and not (inputs(250));
    layer0_outputs(3879) <= inputs(82);
    layer0_outputs(3880) <= (inputs(212)) and not (inputs(186));
    layer0_outputs(3881) <= not((inputs(184)) xor (inputs(43)));
    layer0_outputs(3882) <= not(inputs(122));
    layer0_outputs(3883) <= not((inputs(86)) or (inputs(239)));
    layer0_outputs(3884) <= not(inputs(152));
    layer0_outputs(3885) <= inputs(60);
    layer0_outputs(3886) <= (inputs(15)) or (inputs(213));
    layer0_outputs(3887) <= (inputs(179)) and (inputs(132));
    layer0_outputs(3888) <= not(inputs(179));
    layer0_outputs(3889) <= (inputs(97)) xor (inputs(86));
    layer0_outputs(3890) <= not(inputs(214));
    layer0_outputs(3891) <= (inputs(255)) and not (inputs(169));
    layer0_outputs(3892) <= not((inputs(167)) xor (inputs(148)));
    layer0_outputs(3893) <= (inputs(244)) xor (inputs(224));
    layer0_outputs(3894) <= not(inputs(114)) or (inputs(88));
    layer0_outputs(3895) <= not(inputs(116));
    layer0_outputs(3896) <= not((inputs(61)) or (inputs(104)));
    layer0_outputs(3897) <= not((inputs(113)) or (inputs(189)));
    layer0_outputs(3898) <= not(inputs(111)) or (inputs(255));
    layer0_outputs(3899) <= not(inputs(157));
    layer0_outputs(3900) <= not((inputs(141)) or (inputs(132)));
    layer0_outputs(3901) <= (inputs(230)) and not (inputs(59));
    layer0_outputs(3902) <= inputs(118);
    layer0_outputs(3903) <= '1';
    layer0_outputs(3904) <= not(inputs(74)) or (inputs(135));
    layer0_outputs(3905) <= (inputs(55)) or (inputs(160));
    layer0_outputs(3906) <= (inputs(187)) and not (inputs(95));
    layer0_outputs(3907) <= not(inputs(92)) or (inputs(13));
    layer0_outputs(3908) <= inputs(94);
    layer0_outputs(3909) <= not(inputs(161)) or (inputs(225));
    layer0_outputs(3910) <= not((inputs(198)) xor (inputs(55)));
    layer0_outputs(3911) <= (inputs(27)) and not (inputs(132));
    layer0_outputs(3912) <= (inputs(56)) and not (inputs(210));
    layer0_outputs(3913) <= (inputs(193)) and not (inputs(5));
    layer0_outputs(3914) <= '1';
    layer0_outputs(3915) <= (inputs(71)) and (inputs(219));
    layer0_outputs(3916) <= not(inputs(148));
    layer0_outputs(3917) <= (inputs(176)) or (inputs(125));
    layer0_outputs(3918) <= inputs(23);
    layer0_outputs(3919) <= inputs(199);
    layer0_outputs(3920) <= (inputs(227)) xor (inputs(163));
    layer0_outputs(3921) <= not((inputs(28)) xor (inputs(78)));
    layer0_outputs(3922) <= not((inputs(246)) or (inputs(126)));
    layer0_outputs(3923) <= (inputs(217)) and not (inputs(125));
    layer0_outputs(3924) <= not(inputs(84)) or (inputs(125));
    layer0_outputs(3925) <= not(inputs(67));
    layer0_outputs(3926) <= inputs(203);
    layer0_outputs(3927) <= '1';
    layer0_outputs(3928) <= inputs(27);
    layer0_outputs(3929) <= not(inputs(181));
    layer0_outputs(3930) <= inputs(109);
    layer0_outputs(3931) <= (inputs(132)) xor (inputs(18));
    layer0_outputs(3932) <= not((inputs(200)) xor (inputs(1)));
    layer0_outputs(3933) <= inputs(53);
    layer0_outputs(3934) <= inputs(121);
    layer0_outputs(3935) <= (inputs(118)) and not (inputs(203));
    layer0_outputs(3936) <= not(inputs(128)) or (inputs(31));
    layer0_outputs(3937) <= (inputs(176)) and not (inputs(49));
    layer0_outputs(3938) <= (inputs(97)) or (inputs(67));
    layer0_outputs(3939) <= (inputs(185)) or (inputs(85));
    layer0_outputs(3940) <= inputs(165);
    layer0_outputs(3941) <= inputs(61);
    layer0_outputs(3942) <= not(inputs(134)) or (inputs(172));
    layer0_outputs(3943) <= inputs(87);
    layer0_outputs(3944) <= inputs(187);
    layer0_outputs(3945) <= inputs(99);
    layer0_outputs(3946) <= not((inputs(161)) xor (inputs(245)));
    layer0_outputs(3947) <= inputs(22);
    layer0_outputs(3948) <= inputs(216);
    layer0_outputs(3949) <= (inputs(145)) xor (inputs(100));
    layer0_outputs(3950) <= inputs(77);
    layer0_outputs(3951) <= (inputs(202)) xor (inputs(249));
    layer0_outputs(3952) <= inputs(115);
    layer0_outputs(3953) <= '1';
    layer0_outputs(3954) <= not(inputs(61)) or (inputs(173));
    layer0_outputs(3955) <= not((inputs(250)) or (inputs(104)));
    layer0_outputs(3956) <= (inputs(234)) and not (inputs(100));
    layer0_outputs(3957) <= not((inputs(146)) or (inputs(5)));
    layer0_outputs(3958) <= (inputs(6)) or (inputs(223));
    layer0_outputs(3959) <= inputs(93);
    layer0_outputs(3960) <= not((inputs(225)) or (inputs(217)));
    layer0_outputs(3961) <= '0';
    layer0_outputs(3962) <= not(inputs(230)) or (inputs(59));
    layer0_outputs(3963) <= not(inputs(135));
    layer0_outputs(3964) <= inputs(163);
    layer0_outputs(3965) <= (inputs(218)) and not (inputs(184));
    layer0_outputs(3966) <= not(inputs(146));
    layer0_outputs(3967) <= (inputs(241)) or (inputs(11));
    layer0_outputs(3968) <= inputs(222);
    layer0_outputs(3969) <= inputs(247);
    layer0_outputs(3970) <= not((inputs(229)) xor (inputs(250)));
    layer0_outputs(3971) <= (inputs(189)) and not (inputs(5));
    layer0_outputs(3972) <= inputs(56);
    layer0_outputs(3973) <= not((inputs(157)) xor (inputs(129)));
    layer0_outputs(3974) <= not((inputs(166)) xor (inputs(0)));
    layer0_outputs(3975) <= inputs(213);
    layer0_outputs(3976) <= not(inputs(72)) or (inputs(1));
    layer0_outputs(3977) <= (inputs(221)) xor (inputs(171));
    layer0_outputs(3978) <= (inputs(233)) xor (inputs(146));
    layer0_outputs(3979) <= not(inputs(165));
    layer0_outputs(3980) <= inputs(9);
    layer0_outputs(3981) <= not((inputs(52)) or (inputs(23)));
    layer0_outputs(3982) <= inputs(76);
    layer0_outputs(3983) <= (inputs(103)) and not (inputs(113));
    layer0_outputs(3984) <= not((inputs(245)) and (inputs(22)));
    layer0_outputs(3985) <= (inputs(112)) or (inputs(131));
    layer0_outputs(3986) <= (inputs(122)) or (inputs(118));
    layer0_outputs(3987) <= inputs(148);
    layer0_outputs(3988) <= (inputs(51)) xor (inputs(55));
    layer0_outputs(3989) <= inputs(152);
    layer0_outputs(3990) <= inputs(130);
    layer0_outputs(3991) <= (inputs(241)) and (inputs(32));
    layer0_outputs(3992) <= not(inputs(112));
    layer0_outputs(3993) <= not(inputs(98)) or (inputs(35));
    layer0_outputs(3994) <= inputs(180);
    layer0_outputs(3995) <= not(inputs(92)) or (inputs(72));
    layer0_outputs(3996) <= not((inputs(217)) xor (inputs(178)));
    layer0_outputs(3997) <= not((inputs(206)) or (inputs(186)));
    layer0_outputs(3998) <= not(inputs(58)) or (inputs(17));
    layer0_outputs(3999) <= not((inputs(65)) xor (inputs(245)));
    layer0_outputs(4000) <= (inputs(171)) and not (inputs(32));
    layer0_outputs(4001) <= inputs(198);
    layer0_outputs(4002) <= (inputs(137)) and (inputs(95));
    layer0_outputs(4003) <= not(inputs(213));
    layer0_outputs(4004) <= not(inputs(55));
    layer0_outputs(4005) <= (inputs(43)) xor (inputs(17));
    layer0_outputs(4006) <= not(inputs(30));
    layer0_outputs(4007) <= (inputs(178)) xor (inputs(10));
    layer0_outputs(4008) <= (inputs(116)) or (inputs(63));
    layer0_outputs(4009) <= (inputs(35)) or (inputs(9));
    layer0_outputs(4010) <= not(inputs(170));
    layer0_outputs(4011) <= not((inputs(49)) xor (inputs(15)));
    layer0_outputs(4012) <= (inputs(10)) xor (inputs(129));
    layer0_outputs(4013) <= (inputs(215)) and not (inputs(208));
    layer0_outputs(4014) <= inputs(255);
    layer0_outputs(4015) <= not((inputs(209)) or (inputs(237)));
    layer0_outputs(4016) <= (inputs(79)) or (inputs(193));
    layer0_outputs(4017) <= not(inputs(209)) or (inputs(111));
    layer0_outputs(4018) <= not(inputs(80));
    layer0_outputs(4019) <= not(inputs(226)) or (inputs(14));
    layer0_outputs(4020) <= (inputs(134)) and not (inputs(236));
    layer0_outputs(4021) <= (inputs(92)) xor (inputs(178));
    layer0_outputs(4022) <= not(inputs(101));
    layer0_outputs(4023) <= (inputs(68)) xor (inputs(133));
    layer0_outputs(4024) <= inputs(83);
    layer0_outputs(4025) <= not(inputs(168));
    layer0_outputs(4026) <= inputs(46);
    layer0_outputs(4027) <= inputs(141);
    layer0_outputs(4028) <= inputs(213);
    layer0_outputs(4029) <= (inputs(178)) or (inputs(83));
    layer0_outputs(4030) <= not((inputs(131)) and (inputs(172)));
    layer0_outputs(4031) <= (inputs(9)) and not (inputs(237));
    layer0_outputs(4032) <= (inputs(86)) and not (inputs(204));
    layer0_outputs(4033) <= (inputs(61)) and not (inputs(151));
    layer0_outputs(4034) <= not(inputs(184));
    layer0_outputs(4035) <= not((inputs(226)) xor (inputs(89)));
    layer0_outputs(4036) <= not((inputs(80)) or (inputs(48)));
    layer0_outputs(4037) <= not((inputs(216)) or (inputs(195)));
    layer0_outputs(4038) <= '0';
    layer0_outputs(4039) <= not((inputs(208)) or (inputs(15)));
    layer0_outputs(4040) <= not(inputs(27));
    layer0_outputs(4041) <= inputs(54);
    layer0_outputs(4042) <= not(inputs(83));
    layer0_outputs(4043) <= not((inputs(66)) xor (inputs(228)));
    layer0_outputs(4044) <= (inputs(200)) and (inputs(170));
    layer0_outputs(4045) <= inputs(100);
    layer0_outputs(4046) <= (inputs(126)) xor (inputs(100));
    layer0_outputs(4047) <= (inputs(139)) and not (inputs(243));
    layer0_outputs(4048) <= inputs(17);
    layer0_outputs(4049) <= not(inputs(232)) or (inputs(109));
    layer0_outputs(4050) <= inputs(236);
    layer0_outputs(4051) <= (inputs(49)) or (inputs(44));
    layer0_outputs(4052) <= not(inputs(186));
    layer0_outputs(4053) <= '0';
    layer0_outputs(4054) <= not((inputs(56)) or (inputs(188)));
    layer0_outputs(4055) <= (inputs(99)) and (inputs(54));
    layer0_outputs(4056) <= not(inputs(180));
    layer0_outputs(4057) <= not(inputs(52)) or (inputs(0));
    layer0_outputs(4058) <= not((inputs(95)) xor (inputs(180)));
    layer0_outputs(4059) <= not(inputs(100)) or (inputs(3));
    layer0_outputs(4060) <= not(inputs(239)) or (inputs(108));
    layer0_outputs(4061) <= not((inputs(249)) or (inputs(65)));
    layer0_outputs(4062) <= not(inputs(131));
    layer0_outputs(4063) <= not(inputs(74)) or (inputs(223));
    layer0_outputs(4064) <= (inputs(115)) or (inputs(157));
    layer0_outputs(4065) <= (inputs(211)) and not (inputs(18));
    layer0_outputs(4066) <= not(inputs(247));
    layer0_outputs(4067) <= not(inputs(63));
    layer0_outputs(4068) <= (inputs(140)) or (inputs(75));
    layer0_outputs(4069) <= inputs(6);
    layer0_outputs(4070) <= not((inputs(162)) or (inputs(128)));
    layer0_outputs(4071) <= not((inputs(111)) xor (inputs(93)));
    layer0_outputs(4072) <= (inputs(203)) or (inputs(167));
    layer0_outputs(4073) <= (inputs(227)) and not (inputs(192));
    layer0_outputs(4074) <= not(inputs(132));
    layer0_outputs(4075) <= inputs(234);
    layer0_outputs(4076) <= not(inputs(46));
    layer0_outputs(4077) <= inputs(100);
    layer0_outputs(4078) <= not((inputs(19)) xor (inputs(108)));
    layer0_outputs(4079) <= not(inputs(141));
    layer0_outputs(4080) <= (inputs(205)) or (inputs(197));
    layer0_outputs(4081) <= not(inputs(62));
    layer0_outputs(4082) <= (inputs(175)) and (inputs(31));
    layer0_outputs(4083) <= not((inputs(137)) and (inputs(187)));
    layer0_outputs(4084) <= (inputs(12)) or (inputs(34));
    layer0_outputs(4085) <= inputs(2);
    layer0_outputs(4086) <= (inputs(81)) or (inputs(131));
    layer0_outputs(4087) <= not((inputs(56)) or (inputs(1)));
    layer0_outputs(4088) <= not(inputs(83)) or (inputs(16));
    layer0_outputs(4089) <= not((inputs(182)) xor (inputs(164)));
    layer0_outputs(4090) <= inputs(209);
    layer0_outputs(4091) <= (inputs(163)) and not (inputs(224));
    layer0_outputs(4092) <= not(inputs(195));
    layer0_outputs(4093) <= not((inputs(109)) and (inputs(173)));
    layer0_outputs(4094) <= not((inputs(51)) xor (inputs(60)));
    layer0_outputs(4095) <= not(inputs(97)) or (inputs(223));
    layer0_outputs(4096) <= (inputs(192)) and not (inputs(95));
    layer0_outputs(4097) <= not((inputs(27)) xor (inputs(5)));
    layer0_outputs(4098) <= (inputs(94)) or (inputs(150));
    layer0_outputs(4099) <= not((inputs(232)) or (inputs(204)));
    layer0_outputs(4100) <= not(inputs(106));
    layer0_outputs(4101) <= (inputs(174)) xor (inputs(212));
    layer0_outputs(4102) <= (inputs(119)) and not (inputs(251));
    layer0_outputs(4103) <= (inputs(55)) and not (inputs(32));
    layer0_outputs(4104) <= (inputs(80)) xor (inputs(230));
    layer0_outputs(4105) <= not((inputs(122)) xor (inputs(99)));
    layer0_outputs(4106) <= inputs(36);
    layer0_outputs(4107) <= not(inputs(153));
    layer0_outputs(4108) <= not(inputs(122));
    layer0_outputs(4109) <= not(inputs(115));
    layer0_outputs(4110) <= (inputs(205)) or (inputs(62));
    layer0_outputs(4111) <= inputs(105);
    layer0_outputs(4112) <= not((inputs(115)) xor (inputs(71)));
    layer0_outputs(4113) <= not((inputs(48)) xor (inputs(17)));
    layer0_outputs(4114) <= not(inputs(232)) or (inputs(72));
    layer0_outputs(4115) <= not(inputs(43));
    layer0_outputs(4116) <= not((inputs(76)) xor (inputs(229)));
    layer0_outputs(4117) <= (inputs(224)) or (inputs(196));
    layer0_outputs(4118) <= (inputs(173)) or (inputs(201));
    layer0_outputs(4119) <= inputs(232);
    layer0_outputs(4120) <= (inputs(141)) xor (inputs(101));
    layer0_outputs(4121) <= not(inputs(226));
    layer0_outputs(4122) <= (inputs(164)) and not (inputs(98));
    layer0_outputs(4123) <= not(inputs(248));
    layer0_outputs(4124) <= not(inputs(162)) or (inputs(63));
    layer0_outputs(4125) <= not((inputs(87)) or (inputs(73)));
    layer0_outputs(4126) <= (inputs(96)) xor (inputs(150));
    layer0_outputs(4127) <= not((inputs(171)) or (inputs(243)));
    layer0_outputs(4128) <= not((inputs(6)) xor (inputs(156)));
    layer0_outputs(4129) <= '1';
    layer0_outputs(4130) <= not((inputs(102)) xor (inputs(115)));
    layer0_outputs(4131) <= (inputs(241)) or (inputs(241));
    layer0_outputs(4132) <= not((inputs(62)) or (inputs(34)));
    layer0_outputs(4133) <= inputs(47);
    layer0_outputs(4134) <= (inputs(103)) xor (inputs(74));
    layer0_outputs(4135) <= (inputs(58)) xor (inputs(61));
    layer0_outputs(4136) <= inputs(123);
    layer0_outputs(4137) <= not((inputs(127)) or (inputs(128)));
    layer0_outputs(4138) <= inputs(11);
    layer0_outputs(4139) <= not((inputs(14)) or (inputs(39)));
    layer0_outputs(4140) <= (inputs(253)) and not (inputs(145));
    layer0_outputs(4141) <= (inputs(32)) xor (inputs(12));
    layer0_outputs(4142) <= not((inputs(33)) xor (inputs(124)));
    layer0_outputs(4143) <= not((inputs(157)) or (inputs(191)));
    layer0_outputs(4144) <= not(inputs(66)) or (inputs(228));
    layer0_outputs(4145) <= '1';
    layer0_outputs(4146) <= (inputs(195)) or (inputs(145));
    layer0_outputs(4147) <= not(inputs(101));
    layer0_outputs(4148) <= (inputs(125)) or (inputs(108));
    layer0_outputs(4149) <= (inputs(166)) and not (inputs(242));
    layer0_outputs(4150) <= not(inputs(69)) or (inputs(18));
    layer0_outputs(4151) <= not((inputs(97)) or (inputs(146)));
    layer0_outputs(4152) <= not((inputs(63)) or (inputs(227)));
    layer0_outputs(4153) <= not((inputs(63)) or (inputs(119)));
    layer0_outputs(4154) <= not(inputs(164)) or (inputs(13));
    layer0_outputs(4155) <= (inputs(98)) or (inputs(245));
    layer0_outputs(4156) <= not((inputs(78)) xor (inputs(109)));
    layer0_outputs(4157) <= inputs(232);
    layer0_outputs(4158) <= (inputs(186)) and not (inputs(170));
    layer0_outputs(4159) <= inputs(99);
    layer0_outputs(4160) <= inputs(30);
    layer0_outputs(4161) <= (inputs(118)) and (inputs(254));
    layer0_outputs(4162) <= not((inputs(124)) or (inputs(92)));
    layer0_outputs(4163) <= (inputs(87)) xor (inputs(7));
    layer0_outputs(4164) <= (inputs(186)) or (inputs(194));
    layer0_outputs(4165) <= not((inputs(165)) or (inputs(159)));
    layer0_outputs(4166) <= (inputs(178)) xor (inputs(192));
    layer0_outputs(4167) <= not(inputs(82));
    layer0_outputs(4168) <= not((inputs(118)) xor (inputs(84)));
    layer0_outputs(4169) <= (inputs(64)) xor (inputs(208));
    layer0_outputs(4170) <= not(inputs(252)) or (inputs(67));
    layer0_outputs(4171) <= not(inputs(195));
    layer0_outputs(4172) <= not((inputs(69)) or (inputs(145)));
    layer0_outputs(4173) <= not((inputs(150)) and (inputs(245)));
    layer0_outputs(4174) <= (inputs(14)) or (inputs(162));
    layer0_outputs(4175) <= not(inputs(77));
    layer0_outputs(4176) <= not(inputs(125)) or (inputs(27));
    layer0_outputs(4177) <= not(inputs(158));
    layer0_outputs(4178) <= not((inputs(12)) and (inputs(76)));
    layer0_outputs(4179) <= (inputs(53)) xor (inputs(53));
    layer0_outputs(4180) <= inputs(201);
    layer0_outputs(4181) <= not((inputs(189)) xor (inputs(112)));
    layer0_outputs(4182) <= not(inputs(76)) or (inputs(176));
    layer0_outputs(4183) <= not((inputs(230)) xor (inputs(96)));
    layer0_outputs(4184) <= (inputs(114)) and not (inputs(37));
    layer0_outputs(4185) <= (inputs(2)) xor (inputs(32));
    layer0_outputs(4186) <= (inputs(45)) xor (inputs(218));
    layer0_outputs(4187) <= not((inputs(244)) or (inputs(219)));
    layer0_outputs(4188) <= (inputs(135)) xor (inputs(199));
    layer0_outputs(4189) <= not((inputs(143)) or (inputs(141)));
    layer0_outputs(4190) <= (inputs(204)) or (inputs(35));
    layer0_outputs(4191) <= (inputs(93)) xor (inputs(155));
    layer0_outputs(4192) <= (inputs(135)) xor (inputs(18));
    layer0_outputs(4193) <= not(inputs(137)) or (inputs(255));
    layer0_outputs(4194) <= not(inputs(214));
    layer0_outputs(4195) <= (inputs(236)) and not (inputs(141));
    layer0_outputs(4196) <= not((inputs(184)) xor (inputs(199)));
    layer0_outputs(4197) <= not(inputs(4));
    layer0_outputs(4198) <= not(inputs(195)) or (inputs(72));
    layer0_outputs(4199) <= inputs(202);
    layer0_outputs(4200) <= (inputs(44)) and (inputs(88));
    layer0_outputs(4201) <= not(inputs(91)) or (inputs(19));
    layer0_outputs(4202) <= not(inputs(57));
    layer0_outputs(4203) <= not((inputs(31)) and (inputs(31)));
    layer0_outputs(4204) <= inputs(105);
    layer0_outputs(4205) <= (inputs(117)) and not (inputs(251));
    layer0_outputs(4206) <= not(inputs(247)) or (inputs(37));
    layer0_outputs(4207) <= inputs(60);
    layer0_outputs(4208) <= (inputs(253)) or (inputs(145));
    layer0_outputs(4209) <= (inputs(205)) xor (inputs(85));
    layer0_outputs(4210) <= inputs(223);
    layer0_outputs(4211) <= (inputs(73)) and not (inputs(47));
    layer0_outputs(4212) <= not(inputs(217)) or (inputs(144));
    layer0_outputs(4213) <= (inputs(62)) and (inputs(72));
    layer0_outputs(4214) <= (inputs(66)) or (inputs(112));
    layer0_outputs(4215) <= not(inputs(229)) or (inputs(150));
    layer0_outputs(4216) <= (inputs(208)) xor (inputs(235));
    layer0_outputs(4217) <= not(inputs(145));
    layer0_outputs(4218) <= (inputs(162)) or (inputs(146));
    layer0_outputs(4219) <= (inputs(237)) or (inputs(100));
    layer0_outputs(4220) <= (inputs(121)) xor (inputs(0));
    layer0_outputs(4221) <= (inputs(164)) and not (inputs(181));
    layer0_outputs(4222) <= (inputs(169)) or (inputs(6));
    layer0_outputs(4223) <= (inputs(41)) and not (inputs(32));
    layer0_outputs(4224) <= inputs(245);
    layer0_outputs(4225) <= inputs(207);
    layer0_outputs(4226) <= (inputs(1)) or (inputs(170));
    layer0_outputs(4227) <= inputs(116);
    layer0_outputs(4228) <= not((inputs(89)) or (inputs(32)));
    layer0_outputs(4229) <= (inputs(254)) or (inputs(112));
    layer0_outputs(4230) <= '0';
    layer0_outputs(4231) <= (inputs(68)) or (inputs(176));
    layer0_outputs(4232) <= not(inputs(120));
    layer0_outputs(4233) <= not(inputs(50));
    layer0_outputs(4234) <= not((inputs(20)) or (inputs(191)));
    layer0_outputs(4235) <= '1';
    layer0_outputs(4236) <= not((inputs(243)) xor (inputs(211)));
    layer0_outputs(4237) <= (inputs(220)) xor (inputs(156));
    layer0_outputs(4238) <= inputs(84);
    layer0_outputs(4239) <= inputs(167);
    layer0_outputs(4240) <= (inputs(71)) and not (inputs(105));
    layer0_outputs(4241) <= (inputs(163)) and not (inputs(44));
    layer0_outputs(4242) <= not(inputs(74)) or (inputs(218));
    layer0_outputs(4243) <= (inputs(159)) xor (inputs(235));
    layer0_outputs(4244) <= not((inputs(44)) xor (inputs(46)));
    layer0_outputs(4245) <= not(inputs(102)) or (inputs(48));
    layer0_outputs(4246) <= (inputs(81)) and not (inputs(73));
    layer0_outputs(4247) <= inputs(132);
    layer0_outputs(4248) <= not((inputs(180)) xor (inputs(80)));
    layer0_outputs(4249) <= inputs(253);
    layer0_outputs(4250) <= not((inputs(65)) xor (inputs(188)));
    layer0_outputs(4251) <= not((inputs(20)) xor (inputs(87)));
    layer0_outputs(4252) <= inputs(39);
    layer0_outputs(4253) <= (inputs(168)) or (inputs(166));
    layer0_outputs(4254) <= not(inputs(182)) or (inputs(238));
    layer0_outputs(4255) <= (inputs(58)) or (inputs(95));
    layer0_outputs(4256) <= not(inputs(75));
    layer0_outputs(4257) <= (inputs(246)) and not (inputs(17));
    layer0_outputs(4258) <= not(inputs(74)) or (inputs(102));
    layer0_outputs(4259) <= (inputs(146)) or (inputs(250));
    layer0_outputs(4260) <= (inputs(14)) xor (inputs(87));
    layer0_outputs(4261) <= (inputs(58)) or (inputs(56));
    layer0_outputs(4262) <= not(inputs(85)) or (inputs(214));
    layer0_outputs(4263) <= (inputs(246)) or (inputs(216));
    layer0_outputs(4264) <= not(inputs(164)) or (inputs(112));
    layer0_outputs(4265) <= (inputs(90)) and not (inputs(96));
    layer0_outputs(4266) <= not(inputs(18)) or (inputs(223));
    layer0_outputs(4267) <= not((inputs(71)) or (inputs(143)));
    layer0_outputs(4268) <= inputs(147);
    layer0_outputs(4269) <= (inputs(199)) or (inputs(247));
    layer0_outputs(4270) <= inputs(20);
    layer0_outputs(4271) <= inputs(157);
    layer0_outputs(4272) <= not(inputs(214));
    layer0_outputs(4273) <= not(inputs(94)) or (inputs(149));
    layer0_outputs(4274) <= not(inputs(182));
    layer0_outputs(4275) <= not(inputs(83));
    layer0_outputs(4276) <= inputs(151);
    layer0_outputs(4277) <= (inputs(24)) and (inputs(105));
    layer0_outputs(4278) <= not(inputs(163)) or (inputs(34));
    layer0_outputs(4279) <= (inputs(86)) and not (inputs(141));
    layer0_outputs(4280) <= not(inputs(139));
    layer0_outputs(4281) <= not(inputs(150));
    layer0_outputs(4282) <= not(inputs(115)) or (inputs(190));
    layer0_outputs(4283) <= (inputs(128)) and not (inputs(127));
    layer0_outputs(4284) <= (inputs(147)) or (inputs(236));
    layer0_outputs(4285) <= (inputs(230)) or (inputs(113));
    layer0_outputs(4286) <= (inputs(109)) and (inputs(171));
    layer0_outputs(4287) <= (inputs(245)) and not (inputs(17));
    layer0_outputs(4288) <= not(inputs(254));
    layer0_outputs(4289) <= not(inputs(23));
    layer0_outputs(4290) <= not((inputs(220)) or (inputs(217)));
    layer0_outputs(4291) <= (inputs(26)) and not (inputs(129));
    layer0_outputs(4292) <= (inputs(233)) or (inputs(159));
    layer0_outputs(4293) <= not(inputs(232)) or (inputs(45));
    layer0_outputs(4294) <= not(inputs(121)) or (inputs(130));
    layer0_outputs(4295) <= not((inputs(71)) xor (inputs(199)));
    layer0_outputs(4296) <= not((inputs(159)) or (inputs(10)));
    layer0_outputs(4297) <= (inputs(21)) and not (inputs(143));
    layer0_outputs(4298) <= not((inputs(105)) or (inputs(46)));
    layer0_outputs(4299) <= not(inputs(229));
    layer0_outputs(4300) <= not(inputs(105)) or (inputs(171));
    layer0_outputs(4301) <= not(inputs(5));
    layer0_outputs(4302) <= (inputs(239)) and (inputs(13));
    layer0_outputs(4303) <= not(inputs(91)) or (inputs(230));
    layer0_outputs(4304) <= (inputs(255)) or (inputs(236));
    layer0_outputs(4305) <= (inputs(66)) and not (inputs(225));
    layer0_outputs(4306) <= not((inputs(20)) or (inputs(206)));
    layer0_outputs(4307) <= (inputs(145)) or (inputs(10));
    layer0_outputs(4308) <= inputs(192);
    layer0_outputs(4309) <= inputs(178);
    layer0_outputs(4310) <= (inputs(17)) xor (inputs(153));
    layer0_outputs(4311) <= (inputs(47)) or (inputs(155));
    layer0_outputs(4312) <= not(inputs(77));
    layer0_outputs(4313) <= not(inputs(93));
    layer0_outputs(4314) <= not(inputs(39));
    layer0_outputs(4315) <= (inputs(29)) and not (inputs(185));
    layer0_outputs(4316) <= not((inputs(191)) or (inputs(206)));
    layer0_outputs(4317) <= not((inputs(80)) or (inputs(180)));
    layer0_outputs(4318) <= not(inputs(45)) or (inputs(175));
    layer0_outputs(4319) <= not(inputs(235)) or (inputs(33));
    layer0_outputs(4320) <= not((inputs(64)) xor (inputs(91)));
    layer0_outputs(4321) <= not(inputs(235)) or (inputs(53));
    layer0_outputs(4322) <= (inputs(21)) xor (inputs(89));
    layer0_outputs(4323) <= (inputs(92)) or (inputs(170));
    layer0_outputs(4324) <= not((inputs(77)) or (inputs(185)));
    layer0_outputs(4325) <= inputs(4);
    layer0_outputs(4326) <= not(inputs(223)) or (inputs(210));
    layer0_outputs(4327) <= '1';
    layer0_outputs(4328) <= not((inputs(176)) xor (inputs(148)));
    layer0_outputs(4329) <= not(inputs(116));
    layer0_outputs(4330) <= not(inputs(87));
    layer0_outputs(4331) <= (inputs(121)) xor (inputs(125));
    layer0_outputs(4332) <= (inputs(72)) or (inputs(228));
    layer0_outputs(4333) <= not((inputs(66)) or (inputs(96)));
    layer0_outputs(4334) <= '1';
    layer0_outputs(4335) <= not(inputs(164));
    layer0_outputs(4336) <= (inputs(204)) xor (inputs(93));
    layer0_outputs(4337) <= not(inputs(199)) or (inputs(50));
    layer0_outputs(4338) <= inputs(90);
    layer0_outputs(4339) <= inputs(136);
    layer0_outputs(4340) <= inputs(163);
    layer0_outputs(4341) <= (inputs(109)) and not (inputs(20));
    layer0_outputs(4342) <= inputs(62);
    layer0_outputs(4343) <= '1';
    layer0_outputs(4344) <= not((inputs(155)) or (inputs(37)));
    layer0_outputs(4345) <= (inputs(106)) and not (inputs(2));
    layer0_outputs(4346) <= not(inputs(87));
    layer0_outputs(4347) <= (inputs(247)) or (inputs(160));
    layer0_outputs(4348) <= (inputs(212)) or (inputs(103));
    layer0_outputs(4349) <= not(inputs(136));
    layer0_outputs(4350) <= not(inputs(142));
    layer0_outputs(4351) <= not((inputs(205)) xor (inputs(237)));
    layer0_outputs(4352) <= not((inputs(50)) or (inputs(32)));
    layer0_outputs(4353) <= '1';
    layer0_outputs(4354) <= not((inputs(140)) and (inputs(215)));
    layer0_outputs(4355) <= (inputs(6)) xor (inputs(63));
    layer0_outputs(4356) <= (inputs(14)) or (inputs(168));
    layer0_outputs(4357) <= not(inputs(40));
    layer0_outputs(4358) <= inputs(229);
    layer0_outputs(4359) <= (inputs(48)) or (inputs(165));
    layer0_outputs(4360) <= (inputs(89)) or (inputs(47));
    layer0_outputs(4361) <= not(inputs(181));
    layer0_outputs(4362) <= not(inputs(5));
    layer0_outputs(4363) <= not(inputs(142)) or (inputs(15));
    layer0_outputs(4364) <= (inputs(184)) and not (inputs(127));
    layer0_outputs(4365) <= not(inputs(36));
    layer0_outputs(4366) <= inputs(110);
    layer0_outputs(4367) <= not((inputs(94)) or (inputs(195)));
    layer0_outputs(4368) <= not(inputs(120)) or (inputs(82));
    layer0_outputs(4369) <= '1';
    layer0_outputs(4370) <= (inputs(180)) xor (inputs(254));
    layer0_outputs(4371) <= (inputs(0)) or (inputs(176));
    layer0_outputs(4372) <= (inputs(33)) or (inputs(157));
    layer0_outputs(4373) <= not((inputs(205)) xor (inputs(229)));
    layer0_outputs(4374) <= not((inputs(103)) or (inputs(103)));
    layer0_outputs(4375) <= not(inputs(156));
    layer0_outputs(4376) <= not((inputs(34)) or (inputs(220)));
    layer0_outputs(4377) <= (inputs(88)) xor (inputs(222));
    layer0_outputs(4378) <= not((inputs(221)) xor (inputs(228)));
    layer0_outputs(4379) <= (inputs(97)) or (inputs(237));
    layer0_outputs(4380) <= inputs(125);
    layer0_outputs(4381) <= (inputs(36)) and not (inputs(73));
    layer0_outputs(4382) <= (inputs(156)) or (inputs(173));
    layer0_outputs(4383) <= (inputs(65)) xor (inputs(17));
    layer0_outputs(4384) <= (inputs(234)) and not (inputs(29));
    layer0_outputs(4385) <= inputs(201);
    layer0_outputs(4386) <= inputs(137);
    layer0_outputs(4387) <= (inputs(84)) xor (inputs(196));
    layer0_outputs(4388) <= (inputs(69)) and not (inputs(134));
    layer0_outputs(4389) <= (inputs(166)) or (inputs(130));
    layer0_outputs(4390) <= not((inputs(238)) or (inputs(53)));
    layer0_outputs(4391) <= not((inputs(142)) or (inputs(116)));
    layer0_outputs(4392) <= not((inputs(18)) xor (inputs(81)));
    layer0_outputs(4393) <= not(inputs(120)) or (inputs(65));
    layer0_outputs(4394) <= not(inputs(121));
    layer0_outputs(4395) <= inputs(202);
    layer0_outputs(4396) <= not((inputs(202)) xor (inputs(126)));
    layer0_outputs(4397) <= not((inputs(42)) or (inputs(242)));
    layer0_outputs(4398) <= not(inputs(173)) or (inputs(98));
    layer0_outputs(4399) <= not(inputs(128));
    layer0_outputs(4400) <= inputs(132);
    layer0_outputs(4401) <= (inputs(150)) and (inputs(196));
    layer0_outputs(4402) <= not(inputs(117)) or (inputs(233));
    layer0_outputs(4403) <= (inputs(99)) or (inputs(59));
    layer0_outputs(4404) <= not(inputs(178));
    layer0_outputs(4405) <= not(inputs(183));
    layer0_outputs(4406) <= not(inputs(40));
    layer0_outputs(4407) <= not(inputs(8)) or (inputs(58));
    layer0_outputs(4408) <= (inputs(253)) or (inputs(216));
    layer0_outputs(4409) <= (inputs(18)) or (inputs(188));
    layer0_outputs(4410) <= (inputs(246)) xor (inputs(184));
    layer0_outputs(4411) <= not((inputs(104)) xor (inputs(171)));
    layer0_outputs(4412) <= not((inputs(229)) xor (inputs(215)));
    layer0_outputs(4413) <= not(inputs(173)) or (inputs(66));
    layer0_outputs(4414) <= (inputs(94)) xor (inputs(37));
    layer0_outputs(4415) <= (inputs(118)) or (inputs(238));
    layer0_outputs(4416) <= inputs(211);
    layer0_outputs(4417) <= inputs(9);
    layer0_outputs(4418) <= not((inputs(154)) or (inputs(234)));
    layer0_outputs(4419) <= (inputs(180)) xor (inputs(145));
    layer0_outputs(4420) <= (inputs(27)) xor (inputs(70));
    layer0_outputs(4421) <= '1';
    layer0_outputs(4422) <= (inputs(139)) and (inputs(116));
    layer0_outputs(4423) <= (inputs(47)) and (inputs(200));
    layer0_outputs(4424) <= not(inputs(123)) or (inputs(219));
    layer0_outputs(4425) <= inputs(248);
    layer0_outputs(4426) <= not(inputs(19)) or (inputs(82));
    layer0_outputs(4427) <= inputs(182);
    layer0_outputs(4428) <= not(inputs(249));
    layer0_outputs(4429) <= (inputs(25)) or (inputs(2));
    layer0_outputs(4430) <= not((inputs(161)) or (inputs(143)));
    layer0_outputs(4431) <= (inputs(79)) or (inputs(6));
    layer0_outputs(4432) <= not(inputs(66));
    layer0_outputs(4433) <= (inputs(111)) and not (inputs(60));
    layer0_outputs(4434) <= (inputs(162)) and not (inputs(81));
    layer0_outputs(4435) <= not((inputs(137)) and (inputs(123)));
    layer0_outputs(4436) <= (inputs(86)) xor (inputs(254));
    layer0_outputs(4437) <= not(inputs(58)) or (inputs(239));
    layer0_outputs(4438) <= (inputs(231)) and (inputs(213));
    layer0_outputs(4439) <= not((inputs(119)) xor (inputs(148)));
    layer0_outputs(4440) <= not((inputs(32)) and (inputs(254)));
    layer0_outputs(4441) <= not(inputs(215)) or (inputs(147));
    layer0_outputs(4442) <= not((inputs(227)) xor (inputs(250)));
    layer0_outputs(4443) <= (inputs(138)) xor (inputs(169));
    layer0_outputs(4444) <= not((inputs(200)) or (inputs(4)));
    layer0_outputs(4445) <= (inputs(13)) or (inputs(65));
    layer0_outputs(4446) <= not(inputs(216));
    layer0_outputs(4447) <= not(inputs(153)) or (inputs(3));
    layer0_outputs(4448) <= inputs(22);
    layer0_outputs(4449) <= inputs(163);
    layer0_outputs(4450) <= not((inputs(172)) or (inputs(246)));
    layer0_outputs(4451) <= (inputs(32)) and not (inputs(200));
    layer0_outputs(4452) <= not((inputs(71)) or (inputs(91)));
    layer0_outputs(4453) <= not(inputs(199));
    layer0_outputs(4454) <= not(inputs(161)) or (inputs(255));
    layer0_outputs(4455) <= (inputs(86)) xor (inputs(116));
    layer0_outputs(4456) <= not(inputs(43));
    layer0_outputs(4457) <= not(inputs(3));
    layer0_outputs(4458) <= (inputs(247)) or (inputs(206));
    layer0_outputs(4459) <= (inputs(105)) and not (inputs(224));
    layer0_outputs(4460) <= (inputs(170)) and not (inputs(216));
    layer0_outputs(4461) <= not(inputs(157)) or (inputs(64));
    layer0_outputs(4462) <= (inputs(148)) xor (inputs(67));
    layer0_outputs(4463) <= not(inputs(84)) or (inputs(149));
    layer0_outputs(4464) <= not(inputs(213));
    layer0_outputs(4465) <= not(inputs(114));
    layer0_outputs(4466) <= inputs(26);
    layer0_outputs(4467) <= inputs(148);
    layer0_outputs(4468) <= not((inputs(199)) xor (inputs(18)));
    layer0_outputs(4469) <= (inputs(118)) and not (inputs(5));
    layer0_outputs(4470) <= not(inputs(83)) or (inputs(155));
    layer0_outputs(4471) <= not((inputs(244)) xor (inputs(157)));
    layer0_outputs(4472) <= not(inputs(82)) or (inputs(230));
    layer0_outputs(4473) <= not((inputs(18)) xor (inputs(86)));
    layer0_outputs(4474) <= not(inputs(164));
    layer0_outputs(4475) <= not((inputs(239)) xor (inputs(170)));
    layer0_outputs(4476) <= not((inputs(120)) or (inputs(158)));
    layer0_outputs(4477) <= (inputs(17)) and (inputs(159));
    layer0_outputs(4478) <= (inputs(200)) or (inputs(222));
    layer0_outputs(4479) <= (inputs(152)) and not (inputs(63));
    layer0_outputs(4480) <= not((inputs(161)) xor (inputs(220)));
    layer0_outputs(4481) <= not((inputs(244)) or (inputs(199)));
    layer0_outputs(4482) <= not(inputs(186));
    layer0_outputs(4483) <= (inputs(23)) and not (inputs(129));
    layer0_outputs(4484) <= not(inputs(180));
    layer0_outputs(4485) <= (inputs(81)) xor (inputs(132));
    layer0_outputs(4486) <= not(inputs(210));
    layer0_outputs(4487) <= (inputs(26)) xor (inputs(237));
    layer0_outputs(4488) <= (inputs(213)) and not (inputs(100));
    layer0_outputs(4489) <= inputs(13);
    layer0_outputs(4490) <= not((inputs(69)) or (inputs(76)));
    layer0_outputs(4491) <= not((inputs(213)) xor (inputs(225)));
    layer0_outputs(4492) <= not(inputs(215));
    layer0_outputs(4493) <= not((inputs(168)) xor (inputs(230)));
    layer0_outputs(4494) <= (inputs(116)) and not (inputs(48));
    layer0_outputs(4495) <= (inputs(157)) and not (inputs(226));
    layer0_outputs(4496) <= not((inputs(199)) xor (inputs(220)));
    layer0_outputs(4497) <= (inputs(215)) xor (inputs(36));
    layer0_outputs(4498) <= (inputs(248)) or (inputs(193));
    layer0_outputs(4499) <= (inputs(31)) or (inputs(116));
    layer0_outputs(4500) <= not((inputs(238)) or (inputs(237)));
    layer0_outputs(4501) <= inputs(230);
    layer0_outputs(4502) <= inputs(156);
    layer0_outputs(4503) <= (inputs(109)) and (inputs(143));
    layer0_outputs(4504) <= inputs(139);
    layer0_outputs(4505) <= not(inputs(226));
    layer0_outputs(4506) <= (inputs(210)) or (inputs(174));
    layer0_outputs(4507) <= not((inputs(75)) xor (inputs(119)));
    layer0_outputs(4508) <= (inputs(65)) xor (inputs(245));
    layer0_outputs(4509) <= not((inputs(105)) xor (inputs(207)));
    layer0_outputs(4510) <= not((inputs(232)) xor (inputs(193)));
    layer0_outputs(4511) <= not(inputs(130));
    layer0_outputs(4512) <= not(inputs(98));
    layer0_outputs(4513) <= not(inputs(107));
    layer0_outputs(4514) <= (inputs(118)) and (inputs(208));
    layer0_outputs(4515) <= (inputs(96)) and not (inputs(89));
    layer0_outputs(4516) <= not((inputs(177)) or (inputs(140)));
    layer0_outputs(4517) <= (inputs(112)) or (inputs(35));
    layer0_outputs(4518) <= not(inputs(121));
    layer0_outputs(4519) <= inputs(246);
    layer0_outputs(4520) <= not(inputs(137)) or (inputs(143));
    layer0_outputs(4521) <= (inputs(66)) and not (inputs(13));
    layer0_outputs(4522) <= (inputs(75)) and not (inputs(202));
    layer0_outputs(4523) <= not((inputs(160)) and (inputs(164)));
    layer0_outputs(4524) <= not((inputs(45)) or (inputs(62)));
    layer0_outputs(4525) <= not((inputs(45)) or (inputs(154)));
    layer0_outputs(4526) <= '0';
    layer0_outputs(4527) <= (inputs(126)) and (inputs(107));
    layer0_outputs(4528) <= (inputs(241)) and not (inputs(79));
    layer0_outputs(4529) <= (inputs(232)) and not (inputs(123));
    layer0_outputs(4530) <= not(inputs(102));
    layer0_outputs(4531) <= inputs(77);
    layer0_outputs(4532) <= inputs(71);
    layer0_outputs(4533) <= inputs(189);
    layer0_outputs(4534) <= not((inputs(72)) or (inputs(139)));
    layer0_outputs(4535) <= not((inputs(55)) or (inputs(42)));
    layer0_outputs(4536) <= (inputs(228)) xor (inputs(102));
    layer0_outputs(4537) <= not(inputs(28)) or (inputs(16));
    layer0_outputs(4538) <= inputs(135);
    layer0_outputs(4539) <= (inputs(217)) and not (inputs(108));
    layer0_outputs(4540) <= (inputs(18)) or (inputs(147));
    layer0_outputs(4541) <= inputs(98);
    layer0_outputs(4542) <= (inputs(107)) and (inputs(167));
    layer0_outputs(4543) <= (inputs(8)) or (inputs(245));
    layer0_outputs(4544) <= not(inputs(208)) or (inputs(34));
    layer0_outputs(4545) <= not(inputs(104));
    layer0_outputs(4546) <= inputs(255);
    layer0_outputs(4547) <= (inputs(104)) and not (inputs(223));
    layer0_outputs(4548) <= not(inputs(126));
    layer0_outputs(4549) <= (inputs(92)) xor (inputs(124));
    layer0_outputs(4550) <= not(inputs(30));
    layer0_outputs(4551) <= (inputs(27)) and not (inputs(135));
    layer0_outputs(4552) <= inputs(171);
    layer0_outputs(4553) <= not((inputs(54)) or (inputs(130)));
    layer0_outputs(4554) <= (inputs(69)) and not (inputs(56));
    layer0_outputs(4555) <= not((inputs(18)) or (inputs(152)));
    layer0_outputs(4556) <= (inputs(158)) or (inputs(161));
    layer0_outputs(4557) <= not(inputs(133)) or (inputs(57));
    layer0_outputs(4558) <= (inputs(172)) and not (inputs(232));
    layer0_outputs(4559) <= (inputs(237)) or (inputs(112));
    layer0_outputs(4560) <= not(inputs(210));
    layer0_outputs(4561) <= (inputs(61)) and not (inputs(236));
    layer0_outputs(4562) <= not(inputs(177));
    layer0_outputs(4563) <= (inputs(27)) and not (inputs(173));
    layer0_outputs(4564) <= not((inputs(204)) and (inputs(214)));
    layer0_outputs(4565) <= (inputs(159)) xor (inputs(16));
    layer0_outputs(4566) <= not(inputs(155));
    layer0_outputs(4567) <= not((inputs(181)) xor (inputs(78)));
    layer0_outputs(4568) <= (inputs(222)) or (inputs(230));
    layer0_outputs(4569) <= not(inputs(143)) or (inputs(49));
    layer0_outputs(4570) <= not(inputs(209));
    layer0_outputs(4571) <= inputs(141);
    layer0_outputs(4572) <= not(inputs(155));
    layer0_outputs(4573) <= inputs(220);
    layer0_outputs(4574) <= not((inputs(61)) xor (inputs(36)));
    layer0_outputs(4575) <= inputs(158);
    layer0_outputs(4576) <= not(inputs(123)) or (inputs(227));
    layer0_outputs(4577) <= not(inputs(60)) or (inputs(235));
    layer0_outputs(4578) <= not((inputs(147)) xor (inputs(91)));
    layer0_outputs(4579) <= (inputs(169)) or (inputs(186));
    layer0_outputs(4580) <= not(inputs(44)) or (inputs(251));
    layer0_outputs(4581) <= (inputs(163)) and not (inputs(201));
    layer0_outputs(4582) <= not((inputs(198)) and (inputs(150)));
    layer0_outputs(4583) <= inputs(235);
    layer0_outputs(4584) <= not(inputs(162));
    layer0_outputs(4585) <= (inputs(109)) or (inputs(61));
    layer0_outputs(4586) <= (inputs(33)) xor (inputs(60));
    layer0_outputs(4587) <= not(inputs(138));
    layer0_outputs(4588) <= not(inputs(52));
    layer0_outputs(4589) <= not((inputs(48)) xor (inputs(187)));
    layer0_outputs(4590) <= not((inputs(173)) or (inputs(89)));
    layer0_outputs(4591) <= (inputs(55)) or (inputs(4));
    layer0_outputs(4592) <= (inputs(96)) and not (inputs(155));
    layer0_outputs(4593) <= (inputs(123)) xor (inputs(131));
    layer0_outputs(4594) <= not((inputs(24)) and (inputs(135)));
    layer0_outputs(4595) <= (inputs(215)) and not (inputs(219));
    layer0_outputs(4596) <= (inputs(27)) and not (inputs(146));
    layer0_outputs(4597) <= (inputs(234)) and (inputs(205));
    layer0_outputs(4598) <= not(inputs(118));
    layer0_outputs(4599) <= not(inputs(99)) or (inputs(118));
    layer0_outputs(4600) <= not(inputs(23));
    layer0_outputs(4601) <= inputs(115);
    layer0_outputs(4602) <= not(inputs(83)) or (inputs(29));
    layer0_outputs(4603) <= not((inputs(17)) xor (inputs(39)));
    layer0_outputs(4604) <= '1';
    layer0_outputs(4605) <= not(inputs(7));
    layer0_outputs(4606) <= not(inputs(131)) or (inputs(223));
    layer0_outputs(4607) <= not(inputs(181));
    layer0_outputs(4608) <= (inputs(86)) xor (inputs(225));
    layer0_outputs(4609) <= (inputs(13)) or (inputs(32));
    layer0_outputs(4610) <= '1';
    layer0_outputs(4611) <= not((inputs(170)) or (inputs(204)));
    layer0_outputs(4612) <= not((inputs(43)) xor (inputs(189)));
    layer0_outputs(4613) <= (inputs(11)) or (inputs(176));
    layer0_outputs(4614) <= (inputs(119)) and not (inputs(205));
    layer0_outputs(4615) <= not((inputs(134)) xor (inputs(47)));
    layer0_outputs(4616) <= (inputs(27)) xor (inputs(41));
    layer0_outputs(4617) <= (inputs(187)) and not (inputs(118));
    layer0_outputs(4618) <= not(inputs(85)) or (inputs(255));
    layer0_outputs(4619) <= inputs(118);
    layer0_outputs(4620) <= (inputs(83)) and not (inputs(195));
    layer0_outputs(4621) <= '0';
    layer0_outputs(4622) <= not(inputs(227));
    layer0_outputs(4623) <= (inputs(161)) or (inputs(216));
    layer0_outputs(4624) <= inputs(69);
    layer0_outputs(4625) <= inputs(16);
    layer0_outputs(4626) <= not(inputs(204));
    layer0_outputs(4627) <= (inputs(178)) xor (inputs(87));
    layer0_outputs(4628) <= not((inputs(109)) and (inputs(254)));
    layer0_outputs(4629) <= not((inputs(230)) or (inputs(208)));
    layer0_outputs(4630) <= not((inputs(18)) or (inputs(255)));
    layer0_outputs(4631) <= not(inputs(69));
    layer0_outputs(4632) <= (inputs(246)) or (inputs(160));
    layer0_outputs(4633) <= inputs(72);
    layer0_outputs(4634) <= (inputs(92)) xor (inputs(17));
    layer0_outputs(4635) <= inputs(41);
    layer0_outputs(4636) <= inputs(83);
    layer0_outputs(4637) <= not((inputs(63)) or (inputs(1)));
    layer0_outputs(4638) <= (inputs(217)) or (inputs(6));
    layer0_outputs(4639) <= inputs(62);
    layer0_outputs(4640) <= not(inputs(27)) or (inputs(150));
    layer0_outputs(4641) <= (inputs(159)) or (inputs(179));
    layer0_outputs(4642) <= (inputs(119)) and not (inputs(4));
    layer0_outputs(4643) <= (inputs(47)) or (inputs(50));
    layer0_outputs(4644) <= not((inputs(134)) or (inputs(97)));
    layer0_outputs(4645) <= not((inputs(186)) xor (inputs(139)));
    layer0_outputs(4646) <= inputs(210);
    layer0_outputs(4647) <= not(inputs(131)) or (inputs(220));
    layer0_outputs(4648) <= not((inputs(122)) xor (inputs(210)));
    layer0_outputs(4649) <= not(inputs(248));
    layer0_outputs(4650) <= inputs(212);
    layer0_outputs(4651) <= (inputs(59)) and not (inputs(95));
    layer0_outputs(4652) <= not((inputs(51)) xor (inputs(68)));
    layer0_outputs(4653) <= not((inputs(99)) and (inputs(212)));
    layer0_outputs(4654) <= not(inputs(234));
    layer0_outputs(4655) <= inputs(152);
    layer0_outputs(4656) <= not(inputs(74));
    layer0_outputs(4657) <= (inputs(70)) xor (inputs(129));
    layer0_outputs(4658) <= not((inputs(106)) xor (inputs(156)));
    layer0_outputs(4659) <= '1';
    layer0_outputs(4660) <= not(inputs(11)) or (inputs(210));
    layer0_outputs(4661) <= not((inputs(164)) xor (inputs(112)));
    layer0_outputs(4662) <= (inputs(112)) xor (inputs(98));
    layer0_outputs(4663) <= not(inputs(26)) or (inputs(208));
    layer0_outputs(4664) <= not((inputs(148)) and (inputs(164)));
    layer0_outputs(4665) <= not((inputs(239)) or (inputs(107)));
    layer0_outputs(4666) <= not(inputs(230));
    layer0_outputs(4667) <= '1';
    layer0_outputs(4668) <= not(inputs(191));
    layer0_outputs(4669) <= not((inputs(90)) and (inputs(53)));
    layer0_outputs(4670) <= (inputs(36)) and not (inputs(179));
    layer0_outputs(4671) <= (inputs(132)) and not (inputs(178));
    layer0_outputs(4672) <= not((inputs(45)) or (inputs(19)));
    layer0_outputs(4673) <= (inputs(171)) and not (inputs(49));
    layer0_outputs(4674) <= (inputs(219)) and not (inputs(130));
    layer0_outputs(4675) <= (inputs(190)) and not (inputs(79));
    layer0_outputs(4676) <= not(inputs(83));
    layer0_outputs(4677) <= not(inputs(119)) or (inputs(48));
    layer0_outputs(4678) <= inputs(165);
    layer0_outputs(4679) <= inputs(74);
    layer0_outputs(4680) <= not(inputs(214));
    layer0_outputs(4681) <= (inputs(238)) or (inputs(124));
    layer0_outputs(4682) <= (inputs(62)) and not (inputs(112));
    layer0_outputs(4683) <= inputs(189);
    layer0_outputs(4684) <= not(inputs(129));
    layer0_outputs(4685) <= (inputs(225)) or (inputs(187));
    layer0_outputs(4686) <= (inputs(132)) and not (inputs(17));
    layer0_outputs(4687) <= not((inputs(209)) or (inputs(30)));
    layer0_outputs(4688) <= (inputs(141)) xor (inputs(38));
    layer0_outputs(4689) <= not((inputs(136)) and (inputs(41)));
    layer0_outputs(4690) <= (inputs(152)) or (inputs(206));
    layer0_outputs(4691) <= not(inputs(214)) or (inputs(1));
    layer0_outputs(4692) <= not(inputs(212));
    layer0_outputs(4693) <= inputs(31);
    layer0_outputs(4694) <= (inputs(233)) and not (inputs(134));
    layer0_outputs(4695) <= inputs(217);
    layer0_outputs(4696) <= not(inputs(25));
    layer0_outputs(4697) <= inputs(54);
    layer0_outputs(4698) <= (inputs(29)) and not (inputs(200));
    layer0_outputs(4699) <= not(inputs(43)) or (inputs(64));
    layer0_outputs(4700) <= inputs(100);
    layer0_outputs(4701) <= (inputs(107)) and not (inputs(239));
    layer0_outputs(4702) <= inputs(218);
    layer0_outputs(4703) <= not(inputs(241)) or (inputs(1));
    layer0_outputs(4704) <= not((inputs(41)) xor (inputs(245)));
    layer0_outputs(4705) <= not(inputs(22));
    layer0_outputs(4706) <= (inputs(74)) xor (inputs(217));
    layer0_outputs(4707) <= inputs(146);
    layer0_outputs(4708) <= inputs(57);
    layer0_outputs(4709) <= not(inputs(105)) or (inputs(16));
    layer0_outputs(4710) <= inputs(230);
    layer0_outputs(4711) <= inputs(192);
    layer0_outputs(4712) <= (inputs(133)) or (inputs(50));
    layer0_outputs(4713) <= not((inputs(172)) or (inputs(131)));
    layer0_outputs(4714) <= (inputs(186)) and (inputs(241));
    layer0_outputs(4715) <= not((inputs(137)) or (inputs(121)));
    layer0_outputs(4716) <= (inputs(132)) and not (inputs(22));
    layer0_outputs(4717) <= (inputs(254)) or (inputs(195));
    layer0_outputs(4718) <= not((inputs(249)) or (inputs(111)));
    layer0_outputs(4719) <= not(inputs(211));
    layer0_outputs(4720) <= (inputs(31)) xor (inputs(221));
    layer0_outputs(4721) <= not((inputs(5)) and (inputs(161)));
    layer0_outputs(4722) <= not(inputs(120)) or (inputs(198));
    layer0_outputs(4723) <= (inputs(18)) and not (inputs(142));
    layer0_outputs(4724) <= not(inputs(211));
    layer0_outputs(4725) <= not((inputs(94)) or (inputs(2)));
    layer0_outputs(4726) <= not((inputs(239)) or (inputs(52)));
    layer0_outputs(4727) <= not((inputs(185)) xor (inputs(63)));
    layer0_outputs(4728) <= not((inputs(68)) xor (inputs(251)));
    layer0_outputs(4729) <= not(inputs(196));
    layer0_outputs(4730) <= (inputs(205)) and (inputs(163));
    layer0_outputs(4731) <= inputs(166);
    layer0_outputs(4732) <= not((inputs(158)) xor (inputs(28)));
    layer0_outputs(4733) <= inputs(84);
    layer0_outputs(4734) <= not(inputs(230));
    layer0_outputs(4735) <= not(inputs(52)) or (inputs(172));
    layer0_outputs(4736) <= not((inputs(181)) or (inputs(180)));
    layer0_outputs(4737) <= inputs(47);
    layer0_outputs(4738) <= (inputs(243)) and not (inputs(78));
    layer0_outputs(4739) <= not(inputs(36));
    layer0_outputs(4740) <= (inputs(90)) and not (inputs(33));
    layer0_outputs(4741) <= not((inputs(155)) xor (inputs(62)));
    layer0_outputs(4742) <= not(inputs(23));
    layer0_outputs(4743) <= inputs(171);
    layer0_outputs(4744) <= (inputs(212)) or (inputs(53));
    layer0_outputs(4745) <= not((inputs(237)) or (inputs(232)));
    layer0_outputs(4746) <= not(inputs(205)) or (inputs(80));
    layer0_outputs(4747) <= (inputs(4)) xor (inputs(250));
    layer0_outputs(4748) <= (inputs(182)) or (inputs(86));
    layer0_outputs(4749) <= not((inputs(181)) xor (inputs(183)));
    layer0_outputs(4750) <= not(inputs(105)) or (inputs(136));
    layer0_outputs(4751) <= not(inputs(3));
    layer0_outputs(4752) <= inputs(210);
    layer0_outputs(4753) <= not((inputs(251)) and (inputs(51)));
    layer0_outputs(4754) <= (inputs(34)) xor (inputs(176));
    layer0_outputs(4755) <= (inputs(19)) xor (inputs(15));
    layer0_outputs(4756) <= (inputs(141)) or (inputs(48));
    layer0_outputs(4757) <= not(inputs(116));
    layer0_outputs(4758) <= (inputs(254)) or (inputs(210));
    layer0_outputs(4759) <= inputs(126);
    layer0_outputs(4760) <= not((inputs(150)) xor (inputs(31)));
    layer0_outputs(4761) <= '1';
    layer0_outputs(4762) <= (inputs(128)) or (inputs(129));
    layer0_outputs(4763) <= (inputs(242)) xor (inputs(205));
    layer0_outputs(4764) <= not((inputs(8)) xor (inputs(225)));
    layer0_outputs(4765) <= '1';
    layer0_outputs(4766) <= (inputs(202)) or (inputs(161));
    layer0_outputs(4767) <= not(inputs(101));
    layer0_outputs(4768) <= inputs(231);
    layer0_outputs(4769) <= not((inputs(35)) xor (inputs(25)));
    layer0_outputs(4770) <= not(inputs(9)) or (inputs(44));
    layer0_outputs(4771) <= inputs(214);
    layer0_outputs(4772) <= inputs(113);
    layer0_outputs(4773) <= not((inputs(113)) or (inputs(49)));
    layer0_outputs(4774) <= inputs(247);
    layer0_outputs(4775) <= not(inputs(28));
    layer0_outputs(4776) <= not(inputs(88)) or (inputs(95));
    layer0_outputs(4777) <= inputs(178);
    layer0_outputs(4778) <= not((inputs(193)) or (inputs(33)));
    layer0_outputs(4779) <= (inputs(114)) or (inputs(103));
    layer0_outputs(4780) <= (inputs(150)) and not (inputs(106));
    layer0_outputs(4781) <= (inputs(206)) xor (inputs(186));
    layer0_outputs(4782) <= not(inputs(41)) or (inputs(180));
    layer0_outputs(4783) <= not((inputs(210)) or (inputs(49)));
    layer0_outputs(4784) <= inputs(152);
    layer0_outputs(4785) <= inputs(23);
    layer0_outputs(4786) <= (inputs(76)) and not (inputs(217));
    layer0_outputs(4787) <= (inputs(199)) and (inputs(218));
    layer0_outputs(4788) <= inputs(126);
    layer0_outputs(4789) <= not(inputs(120));
    layer0_outputs(4790) <= (inputs(238)) and not (inputs(240));
    layer0_outputs(4791) <= (inputs(28)) and not (inputs(149));
    layer0_outputs(4792) <= (inputs(123)) or (inputs(19));
    layer0_outputs(4793) <= inputs(83);
    layer0_outputs(4794) <= not((inputs(28)) xor (inputs(54)));
    layer0_outputs(4795) <= (inputs(6)) xor (inputs(213));
    layer0_outputs(4796) <= not((inputs(218)) xor (inputs(141)));
    layer0_outputs(4797) <= inputs(140);
    layer0_outputs(4798) <= (inputs(194)) and not (inputs(186));
    layer0_outputs(4799) <= (inputs(89)) and not (inputs(33));
    layer0_outputs(4800) <= not(inputs(62)) or (inputs(223));
    layer0_outputs(4801) <= inputs(21);
    layer0_outputs(4802) <= not(inputs(38)) or (inputs(228));
    layer0_outputs(4803) <= (inputs(118)) and not (inputs(170));
    layer0_outputs(4804) <= (inputs(115)) and not (inputs(23));
    layer0_outputs(4805) <= not(inputs(103)) or (inputs(126));
    layer0_outputs(4806) <= not(inputs(99)) or (inputs(240));
    layer0_outputs(4807) <= not(inputs(175));
    layer0_outputs(4808) <= (inputs(108)) and not (inputs(207));
    layer0_outputs(4809) <= (inputs(245)) or (inputs(177));
    layer0_outputs(4810) <= (inputs(133)) xor (inputs(21));
    layer0_outputs(4811) <= inputs(184);
    layer0_outputs(4812) <= (inputs(177)) and (inputs(238));
    layer0_outputs(4813) <= inputs(117);
    layer0_outputs(4814) <= (inputs(76)) and (inputs(90));
    layer0_outputs(4815) <= inputs(150);
    layer0_outputs(4816) <= not(inputs(26));
    layer0_outputs(4817) <= not(inputs(106)) or (inputs(253));
    layer0_outputs(4818) <= (inputs(179)) or (inputs(130));
    layer0_outputs(4819) <= not((inputs(243)) or (inputs(206)));
    layer0_outputs(4820) <= not((inputs(29)) or (inputs(128)));
    layer0_outputs(4821) <= not((inputs(204)) xor (inputs(161)));
    layer0_outputs(4822) <= (inputs(143)) or (inputs(169));
    layer0_outputs(4823) <= not(inputs(136)) or (inputs(113));
    layer0_outputs(4824) <= not(inputs(230));
    layer0_outputs(4825) <= (inputs(130)) and not (inputs(50));
    layer0_outputs(4826) <= not(inputs(98));
    layer0_outputs(4827) <= not(inputs(188));
    layer0_outputs(4828) <= (inputs(93)) or (inputs(56));
    layer0_outputs(4829) <= (inputs(144)) and not (inputs(162));
    layer0_outputs(4830) <= not((inputs(109)) and (inputs(211)));
    layer0_outputs(4831) <= inputs(166);
    layer0_outputs(4832) <= (inputs(161)) xor (inputs(173));
    layer0_outputs(4833) <= (inputs(183)) xor (inputs(231));
    layer0_outputs(4834) <= (inputs(92)) xor (inputs(2));
    layer0_outputs(4835) <= not((inputs(138)) or (inputs(47)));
    layer0_outputs(4836) <= (inputs(10)) xor (inputs(155));
    layer0_outputs(4837) <= (inputs(153)) xor (inputs(151));
    layer0_outputs(4838) <= not(inputs(191));
    layer0_outputs(4839) <= (inputs(121)) or (inputs(81));
    layer0_outputs(4840) <= not((inputs(248)) and (inputs(247)));
    layer0_outputs(4841) <= not((inputs(85)) xor (inputs(180)));
    layer0_outputs(4842) <= not(inputs(103));
    layer0_outputs(4843) <= not(inputs(211)) or (inputs(9));
    layer0_outputs(4844) <= not(inputs(23));
    layer0_outputs(4845) <= not((inputs(24)) and (inputs(22)));
    layer0_outputs(4846) <= (inputs(183)) or (inputs(169));
    layer0_outputs(4847) <= not(inputs(248));
    layer0_outputs(4848) <= not(inputs(88));
    layer0_outputs(4849) <= not(inputs(220));
    layer0_outputs(4850) <= inputs(231);
    layer0_outputs(4851) <= inputs(19);
    layer0_outputs(4852) <= inputs(103);
    layer0_outputs(4853) <= (inputs(95)) or (inputs(222));
    layer0_outputs(4854) <= not(inputs(232));
    layer0_outputs(4855) <= not(inputs(104));
    layer0_outputs(4856) <= (inputs(246)) and not (inputs(237));
    layer0_outputs(4857) <= inputs(151);
    layer0_outputs(4858) <= (inputs(142)) and not (inputs(244));
    layer0_outputs(4859) <= (inputs(62)) or (inputs(25));
    layer0_outputs(4860) <= (inputs(47)) and (inputs(96));
    layer0_outputs(4861) <= not((inputs(14)) or (inputs(204)));
    layer0_outputs(4862) <= '1';
    layer0_outputs(4863) <= not(inputs(138));
    layer0_outputs(4864) <= not(inputs(163));
    layer0_outputs(4865) <= (inputs(108)) xor (inputs(113));
    layer0_outputs(4866) <= not(inputs(214));
    layer0_outputs(4867) <= inputs(121);
    layer0_outputs(4868) <= not((inputs(192)) or (inputs(102)));
    layer0_outputs(4869) <= (inputs(131)) xor (inputs(145));
    layer0_outputs(4870) <= not(inputs(51));
    layer0_outputs(4871) <= not(inputs(180));
    layer0_outputs(4872) <= inputs(130);
    layer0_outputs(4873) <= (inputs(81)) xor (inputs(188));
    layer0_outputs(4874) <= inputs(138);
    layer0_outputs(4875) <= '1';
    layer0_outputs(4876) <= not(inputs(46));
    layer0_outputs(4877) <= '0';
    layer0_outputs(4878) <= not((inputs(180)) xor (inputs(90)));
    layer0_outputs(4879) <= (inputs(199)) xor (inputs(149));
    layer0_outputs(4880) <= inputs(148);
    layer0_outputs(4881) <= (inputs(44)) or (inputs(127));
    layer0_outputs(4882) <= (inputs(82)) xor (inputs(31));
    layer0_outputs(4883) <= not((inputs(87)) xor (inputs(112)));
    layer0_outputs(4884) <= not(inputs(129)) or (inputs(154));
    layer0_outputs(4885) <= not(inputs(211)) or (inputs(45));
    layer0_outputs(4886) <= (inputs(137)) and not (inputs(65));
    layer0_outputs(4887) <= not((inputs(51)) or (inputs(167)));
    layer0_outputs(4888) <= (inputs(234)) xor (inputs(10));
    layer0_outputs(4889) <= not((inputs(98)) or (inputs(228)));
    layer0_outputs(4890) <= inputs(44);
    layer0_outputs(4891) <= not((inputs(28)) xor (inputs(2)));
    layer0_outputs(4892) <= not(inputs(110));
    layer0_outputs(4893) <= not(inputs(217));
    layer0_outputs(4894) <= not(inputs(15));
    layer0_outputs(4895) <= '0';
    layer0_outputs(4896) <= not((inputs(18)) xor (inputs(253)));
    layer0_outputs(4897) <= not(inputs(158));
    layer0_outputs(4898) <= (inputs(225)) or (inputs(26));
    layer0_outputs(4899) <= (inputs(226)) or (inputs(87));
    layer0_outputs(4900) <= not((inputs(44)) or (inputs(248)));
    layer0_outputs(4901) <= not(inputs(29)) or (inputs(85));
    layer0_outputs(4902) <= not((inputs(20)) xor (inputs(239)));
    layer0_outputs(4903) <= (inputs(127)) or (inputs(155));
    layer0_outputs(4904) <= not(inputs(122));
    layer0_outputs(4905) <= (inputs(190)) or (inputs(86));
    layer0_outputs(4906) <= (inputs(146)) or (inputs(252));
    layer0_outputs(4907) <= not(inputs(239));
    layer0_outputs(4908) <= (inputs(58)) and (inputs(177));
    layer0_outputs(4909) <= not(inputs(100));
    layer0_outputs(4910) <= (inputs(229)) xor (inputs(223));
    layer0_outputs(4911) <= inputs(57);
    layer0_outputs(4912) <= (inputs(210)) and not (inputs(236));
    layer0_outputs(4913) <= '0';
    layer0_outputs(4914) <= not((inputs(76)) or (inputs(60)));
    layer0_outputs(4915) <= (inputs(177)) xor (inputs(147));
    layer0_outputs(4916) <= (inputs(206)) or (inputs(220));
    layer0_outputs(4917) <= '0';
    layer0_outputs(4918) <= not((inputs(135)) and (inputs(83)));
    layer0_outputs(4919) <= (inputs(60)) or (inputs(7));
    layer0_outputs(4920) <= (inputs(170)) xor (inputs(32));
    layer0_outputs(4921) <= (inputs(151)) or (inputs(179));
    layer0_outputs(4922) <= not((inputs(84)) xor (inputs(21)));
    layer0_outputs(4923) <= not(inputs(214));
    layer0_outputs(4924) <= (inputs(7)) or (inputs(250));
    layer0_outputs(4925) <= inputs(42);
    layer0_outputs(4926) <= not(inputs(183));
    layer0_outputs(4927) <= inputs(221);
    layer0_outputs(4928) <= not(inputs(31));
    layer0_outputs(4929) <= not((inputs(26)) or (inputs(52)));
    layer0_outputs(4930) <= (inputs(161)) xor (inputs(1));
    layer0_outputs(4931) <= not((inputs(13)) or (inputs(240)));
    layer0_outputs(4932) <= inputs(76);
    layer0_outputs(4933) <= not((inputs(35)) and (inputs(21)));
    layer0_outputs(4934) <= not(inputs(60)) or (inputs(220));
    layer0_outputs(4935) <= (inputs(182)) xor (inputs(90));
    layer0_outputs(4936) <= (inputs(192)) xor (inputs(135));
    layer0_outputs(4937) <= not((inputs(19)) or (inputs(222)));
    layer0_outputs(4938) <= (inputs(70)) and not (inputs(161));
    layer0_outputs(4939) <= (inputs(154)) xor (inputs(86));
    layer0_outputs(4940) <= (inputs(58)) and (inputs(38));
    layer0_outputs(4941) <= not((inputs(234)) xor (inputs(224)));
    layer0_outputs(4942) <= (inputs(195)) or (inputs(6));
    layer0_outputs(4943) <= not(inputs(82));
    layer0_outputs(4944) <= not((inputs(233)) xor (inputs(47)));
    layer0_outputs(4945) <= not((inputs(170)) or (inputs(171)));
    layer0_outputs(4946) <= (inputs(120)) or (inputs(46));
    layer0_outputs(4947) <= inputs(25);
    layer0_outputs(4948) <= (inputs(40)) and not (inputs(164));
    layer0_outputs(4949) <= not(inputs(52));
    layer0_outputs(4950) <= inputs(54);
    layer0_outputs(4951) <= (inputs(46)) and (inputs(22));
    layer0_outputs(4952) <= not(inputs(209));
    layer0_outputs(4953) <= not(inputs(97));
    layer0_outputs(4954) <= not((inputs(138)) xor (inputs(193)));
    layer0_outputs(4955) <= (inputs(23)) xor (inputs(79));
    layer0_outputs(4956) <= (inputs(65)) and not (inputs(251));
    layer0_outputs(4957) <= not(inputs(163)) or (inputs(96));
    layer0_outputs(4958) <= not((inputs(222)) or (inputs(148)));
    layer0_outputs(4959) <= (inputs(17)) and not (inputs(108));
    layer0_outputs(4960) <= not(inputs(94));
    layer0_outputs(4961) <= (inputs(173)) and not (inputs(208));
    layer0_outputs(4962) <= inputs(65);
    layer0_outputs(4963) <= inputs(99);
    layer0_outputs(4964) <= not((inputs(29)) or (inputs(128)));
    layer0_outputs(4965) <= (inputs(102)) or (inputs(77));
    layer0_outputs(4966) <= not((inputs(173)) xor (inputs(202)));
    layer0_outputs(4967) <= not((inputs(0)) or (inputs(209)));
    layer0_outputs(4968) <= inputs(104);
    layer0_outputs(4969) <= not(inputs(158)) or (inputs(106));
    layer0_outputs(4970) <= inputs(69);
    layer0_outputs(4971) <= not((inputs(172)) xor (inputs(111)));
    layer0_outputs(4972) <= (inputs(233)) or (inputs(176));
    layer0_outputs(4973) <= not(inputs(93)) or (inputs(81));
    layer0_outputs(4974) <= not((inputs(216)) and (inputs(27)));
    layer0_outputs(4975) <= (inputs(177)) xor (inputs(87));
    layer0_outputs(4976) <= not(inputs(155)) or (inputs(12));
    layer0_outputs(4977) <= (inputs(121)) or (inputs(191));
    layer0_outputs(4978) <= not(inputs(182));
    layer0_outputs(4979) <= not((inputs(90)) xor (inputs(110)));
    layer0_outputs(4980) <= not(inputs(147));
    layer0_outputs(4981) <= not(inputs(158)) or (inputs(169));
    layer0_outputs(4982) <= (inputs(52)) or (inputs(95));
    layer0_outputs(4983) <= (inputs(66)) xor (inputs(101));
    layer0_outputs(4984) <= not(inputs(49)) or (inputs(145));
    layer0_outputs(4985) <= inputs(123);
    layer0_outputs(4986) <= (inputs(118)) xor (inputs(15));
    layer0_outputs(4987) <= inputs(71);
    layer0_outputs(4988) <= not(inputs(106)) or (inputs(206));
    layer0_outputs(4989) <= (inputs(133)) and not (inputs(7));
    layer0_outputs(4990) <= (inputs(59)) xor (inputs(233));
    layer0_outputs(4991) <= inputs(217);
    layer0_outputs(4992) <= (inputs(211)) xor (inputs(240));
    layer0_outputs(4993) <= inputs(70);
    layer0_outputs(4994) <= (inputs(60)) or (inputs(128));
    layer0_outputs(4995) <= not(inputs(193)) or (inputs(184));
    layer0_outputs(4996) <= (inputs(131)) or (inputs(109));
    layer0_outputs(4997) <= inputs(142);
    layer0_outputs(4998) <= inputs(97);
    layer0_outputs(4999) <= not(inputs(14)) or (inputs(66));
    layer0_outputs(5000) <= not((inputs(214)) and (inputs(102)));
    layer0_outputs(5001) <= not(inputs(27));
    layer0_outputs(5002) <= inputs(43);
    layer0_outputs(5003) <= not(inputs(4));
    layer0_outputs(5004) <= '1';
    layer0_outputs(5005) <= (inputs(217)) xor (inputs(55));
    layer0_outputs(5006) <= (inputs(95)) or (inputs(24));
    layer0_outputs(5007) <= inputs(203);
    layer0_outputs(5008) <= not((inputs(196)) xor (inputs(120)));
    layer0_outputs(5009) <= (inputs(217)) and not (inputs(18));
    layer0_outputs(5010) <= (inputs(124)) xor (inputs(165));
    layer0_outputs(5011) <= (inputs(195)) xor (inputs(122));
    layer0_outputs(5012) <= not(inputs(129));
    layer0_outputs(5013) <= inputs(151);
    layer0_outputs(5014) <= inputs(169);
    layer0_outputs(5015) <= not((inputs(86)) or (inputs(250)));
    layer0_outputs(5016) <= not((inputs(71)) xor (inputs(8)));
    layer0_outputs(5017) <= not(inputs(245));
    layer0_outputs(5018) <= inputs(77);
    layer0_outputs(5019) <= not(inputs(226)) or (inputs(44));
    layer0_outputs(5020) <= (inputs(206)) xor (inputs(188));
    layer0_outputs(5021) <= not((inputs(0)) or (inputs(198)));
    layer0_outputs(5022) <= not((inputs(12)) or (inputs(26)));
    layer0_outputs(5023) <= inputs(42);
    layer0_outputs(5024) <= not((inputs(233)) or (inputs(107)));
    layer0_outputs(5025) <= not(inputs(196));
    layer0_outputs(5026) <= (inputs(193)) xor (inputs(114));
    layer0_outputs(5027) <= not(inputs(206)) or (inputs(255));
    layer0_outputs(5028) <= not(inputs(99)) or (inputs(61));
    layer0_outputs(5029) <= not(inputs(59));
    layer0_outputs(5030) <= not((inputs(161)) or (inputs(116)));
    layer0_outputs(5031) <= not((inputs(56)) or (inputs(95)));
    layer0_outputs(5032) <= (inputs(5)) xor (inputs(88));
    layer0_outputs(5033) <= inputs(228);
    layer0_outputs(5034) <= not((inputs(45)) xor (inputs(35)));
    layer0_outputs(5035) <= not(inputs(103));
    layer0_outputs(5036) <= (inputs(141)) and (inputs(74));
    layer0_outputs(5037) <= not(inputs(131)) or (inputs(83));
    layer0_outputs(5038) <= not(inputs(156)) or (inputs(242));
    layer0_outputs(5039) <= (inputs(25)) or (inputs(64));
    layer0_outputs(5040) <= not(inputs(234)) or (inputs(47));
    layer0_outputs(5041) <= inputs(234);
    layer0_outputs(5042) <= (inputs(20)) or (inputs(7));
    layer0_outputs(5043) <= not((inputs(148)) or (inputs(75)));
    layer0_outputs(5044) <= not(inputs(233));
    layer0_outputs(5045) <= (inputs(220)) xor (inputs(38));
    layer0_outputs(5046) <= not((inputs(1)) or (inputs(209)));
    layer0_outputs(5047) <= not((inputs(121)) or (inputs(17)));
    layer0_outputs(5048) <= not(inputs(147));
    layer0_outputs(5049) <= inputs(139);
    layer0_outputs(5050) <= (inputs(227)) or (inputs(57));
    layer0_outputs(5051) <= not((inputs(217)) xor (inputs(114)));
    layer0_outputs(5052) <= not(inputs(166));
    layer0_outputs(5053) <= inputs(98);
    layer0_outputs(5054) <= (inputs(180)) or (inputs(176));
    layer0_outputs(5055) <= (inputs(202)) or (inputs(205));
    layer0_outputs(5056) <= inputs(231);
    layer0_outputs(5057) <= (inputs(139)) and not (inputs(235));
    layer0_outputs(5058) <= not(inputs(150));
    layer0_outputs(5059) <= not(inputs(76));
    layer0_outputs(5060) <= (inputs(66)) and not (inputs(135));
    layer0_outputs(5061) <= not(inputs(252));
    layer0_outputs(5062) <= not((inputs(2)) or (inputs(160)));
    layer0_outputs(5063) <= not((inputs(67)) or (inputs(177)));
    layer0_outputs(5064) <= inputs(231);
    layer0_outputs(5065) <= (inputs(17)) and (inputs(204));
    layer0_outputs(5066) <= not((inputs(53)) xor (inputs(168)));
    layer0_outputs(5067) <= not(inputs(208));
    layer0_outputs(5068) <= (inputs(46)) xor (inputs(13));
    layer0_outputs(5069) <= (inputs(223)) or (inputs(97));
    layer0_outputs(5070) <= not(inputs(90)) or (inputs(192));
    layer0_outputs(5071) <= not(inputs(168)) or (inputs(117));
    layer0_outputs(5072) <= (inputs(171)) and not (inputs(47));
    layer0_outputs(5073) <= inputs(212);
    layer0_outputs(5074) <= not(inputs(131));
    layer0_outputs(5075) <= not((inputs(226)) or (inputs(180)));
    layer0_outputs(5076) <= inputs(228);
    layer0_outputs(5077) <= not(inputs(29));
    layer0_outputs(5078) <= '0';
    layer0_outputs(5079) <= not(inputs(210));
    layer0_outputs(5080) <= not((inputs(5)) xor (inputs(238)));
    layer0_outputs(5081) <= inputs(151);
    layer0_outputs(5082) <= not(inputs(211)) or (inputs(246));
    layer0_outputs(5083) <= (inputs(174)) xor (inputs(2));
    layer0_outputs(5084) <= not(inputs(76)) or (inputs(175));
    layer0_outputs(5085) <= not(inputs(90));
    layer0_outputs(5086) <= (inputs(197)) and not (inputs(44));
    layer0_outputs(5087) <= (inputs(24)) xor (inputs(75));
    layer0_outputs(5088) <= inputs(216);
    layer0_outputs(5089) <= (inputs(22)) or (inputs(224));
    layer0_outputs(5090) <= not(inputs(22));
    layer0_outputs(5091) <= (inputs(62)) xor (inputs(198));
    layer0_outputs(5092) <= not((inputs(170)) xor (inputs(204)));
    layer0_outputs(5093) <= '1';
    layer0_outputs(5094) <= not(inputs(164));
    layer0_outputs(5095) <= (inputs(78)) or (inputs(186));
    layer0_outputs(5096) <= (inputs(234)) xor (inputs(70));
    layer0_outputs(5097) <= (inputs(50)) and not (inputs(28));
    layer0_outputs(5098) <= not(inputs(154)) or (inputs(75));
    layer0_outputs(5099) <= (inputs(117)) xor (inputs(98));
    layer0_outputs(5100) <= not(inputs(88));
    layer0_outputs(5101) <= inputs(74);
    layer0_outputs(5102) <= not(inputs(39));
    layer0_outputs(5103) <= not(inputs(177));
    layer0_outputs(5104) <= not(inputs(107)) or (inputs(201));
    layer0_outputs(5105) <= not(inputs(212));
    layer0_outputs(5106) <= (inputs(179)) and not (inputs(0));
    layer0_outputs(5107) <= inputs(212);
    layer0_outputs(5108) <= (inputs(85)) and not (inputs(192));
    layer0_outputs(5109) <= inputs(60);
    layer0_outputs(5110) <= inputs(165);
    layer0_outputs(5111) <= (inputs(99)) xor (inputs(46));
    layer0_outputs(5112) <= inputs(46);
    layer0_outputs(5113) <= not((inputs(159)) or (inputs(232)));
    layer0_outputs(5114) <= not((inputs(110)) xor (inputs(63)));
    layer0_outputs(5115) <= not((inputs(126)) or (inputs(146)));
    layer0_outputs(5116) <= inputs(180);
    layer0_outputs(5117) <= not((inputs(171)) and (inputs(0)));
    layer0_outputs(5118) <= (inputs(76)) and (inputs(103));
    layer0_outputs(5119) <= (inputs(7)) xor (inputs(79));
    layer0_outputs(5120) <= not(inputs(110)) or (inputs(106));
    layer0_outputs(5121) <= inputs(153);
    layer0_outputs(5122) <= (inputs(136)) or (inputs(183));
    layer0_outputs(5123) <= not((inputs(151)) and (inputs(190)));
    layer0_outputs(5124) <= not(inputs(233));
    layer0_outputs(5125) <= not(inputs(244));
    layer0_outputs(5126) <= (inputs(63)) or (inputs(2));
    layer0_outputs(5127) <= not(inputs(36)) or (inputs(254));
    layer0_outputs(5128) <= (inputs(225)) xor (inputs(3));
    layer0_outputs(5129) <= not(inputs(63)) or (inputs(141));
    layer0_outputs(5130) <= not(inputs(68)) or (inputs(33));
    layer0_outputs(5131) <= not(inputs(199)) or (inputs(137));
    layer0_outputs(5132) <= not(inputs(133));
    layer0_outputs(5133) <= not((inputs(113)) or (inputs(75)));
    layer0_outputs(5134) <= (inputs(251)) or (inputs(221));
    layer0_outputs(5135) <= inputs(121);
    layer0_outputs(5136) <= not(inputs(145));
    layer0_outputs(5137) <= not((inputs(179)) or (inputs(237)));
    layer0_outputs(5138) <= not(inputs(27));
    layer0_outputs(5139) <= not(inputs(13));
    layer0_outputs(5140) <= not(inputs(151)) or (inputs(47));
    layer0_outputs(5141) <= not(inputs(10));
    layer0_outputs(5142) <= (inputs(226)) or (inputs(225));
    layer0_outputs(5143) <= (inputs(98)) and not (inputs(73));
    layer0_outputs(5144) <= (inputs(26)) and not (inputs(154));
    layer0_outputs(5145) <= not(inputs(182)) or (inputs(45));
    layer0_outputs(5146) <= (inputs(195)) and not (inputs(224));
    layer0_outputs(5147) <= inputs(177);
    layer0_outputs(5148) <= (inputs(148)) or (inputs(176));
    layer0_outputs(5149) <= not((inputs(56)) or (inputs(24)));
    layer0_outputs(5150) <= not((inputs(61)) or (inputs(182)));
    layer0_outputs(5151) <= not(inputs(100)) or (inputs(224));
    layer0_outputs(5152) <= (inputs(67)) or (inputs(44));
    layer0_outputs(5153) <= not((inputs(7)) xor (inputs(158)));
    layer0_outputs(5154) <= (inputs(201)) xor (inputs(79));
    layer0_outputs(5155) <= (inputs(133)) and not (inputs(108));
    layer0_outputs(5156) <= not((inputs(168)) and (inputs(5)));
    layer0_outputs(5157) <= not((inputs(111)) and (inputs(186)));
    layer0_outputs(5158) <= (inputs(139)) and (inputs(254));
    layer0_outputs(5159) <= (inputs(64)) or (inputs(149));
    layer0_outputs(5160) <= (inputs(52)) and not (inputs(226));
    layer0_outputs(5161) <= not((inputs(242)) xor (inputs(241)));
    layer0_outputs(5162) <= not(inputs(9));
    layer0_outputs(5163) <= (inputs(136)) or (inputs(48));
    layer0_outputs(5164) <= not(inputs(62)) or (inputs(139));
    layer0_outputs(5165) <= not(inputs(68)) or (inputs(181));
    layer0_outputs(5166) <= (inputs(176)) or (inputs(195));
    layer0_outputs(5167) <= (inputs(56)) and not (inputs(175));
    layer0_outputs(5168) <= not(inputs(252));
    layer0_outputs(5169) <= not(inputs(92));
    layer0_outputs(5170) <= not((inputs(25)) and (inputs(44)));
    layer0_outputs(5171) <= '0';
    layer0_outputs(5172) <= not((inputs(224)) or (inputs(136)));
    layer0_outputs(5173) <= (inputs(248)) xor (inputs(30));
    layer0_outputs(5174) <= inputs(165);
    layer0_outputs(5175) <= inputs(108);
    layer0_outputs(5176) <= (inputs(18)) xor (inputs(187));
    layer0_outputs(5177) <= not(inputs(133)) or (inputs(33));
    layer0_outputs(5178) <= inputs(163);
    layer0_outputs(5179) <= not(inputs(211));
    layer0_outputs(5180) <= '0';
    layer0_outputs(5181) <= not((inputs(101)) xor (inputs(225)));
    layer0_outputs(5182) <= inputs(193);
    layer0_outputs(5183) <= not(inputs(135));
    layer0_outputs(5184) <= not((inputs(199)) or (inputs(86)));
    layer0_outputs(5185) <= not(inputs(229));
    layer0_outputs(5186) <= not(inputs(83));
    layer0_outputs(5187) <= inputs(93);
    layer0_outputs(5188) <= (inputs(74)) and (inputs(203));
    layer0_outputs(5189) <= not((inputs(196)) or (inputs(214)));
    layer0_outputs(5190) <= (inputs(203)) or (inputs(34));
    layer0_outputs(5191) <= not((inputs(31)) and (inputs(175)));
    layer0_outputs(5192) <= not(inputs(158)) or (inputs(198));
    layer0_outputs(5193) <= (inputs(116)) and not (inputs(0));
    layer0_outputs(5194) <= (inputs(23)) and not (inputs(128));
    layer0_outputs(5195) <= not(inputs(196));
    layer0_outputs(5196) <= (inputs(251)) xor (inputs(104));
    layer0_outputs(5197) <= not(inputs(200)) or (inputs(54));
    layer0_outputs(5198) <= not(inputs(106));
    layer0_outputs(5199) <= (inputs(106)) and not (inputs(224));
    layer0_outputs(5200) <= (inputs(240)) and not (inputs(51));
    layer0_outputs(5201) <= (inputs(130)) xor (inputs(57));
    layer0_outputs(5202) <= not(inputs(161)) or (inputs(122));
    layer0_outputs(5203) <= not((inputs(86)) or (inputs(191)));
    layer0_outputs(5204) <= inputs(230);
    layer0_outputs(5205) <= not(inputs(238));
    layer0_outputs(5206) <= (inputs(19)) xor (inputs(220));
    layer0_outputs(5207) <= (inputs(130)) xor (inputs(31));
    layer0_outputs(5208) <= inputs(148);
    layer0_outputs(5209) <= not((inputs(177)) xor (inputs(233)));
    layer0_outputs(5210) <= not((inputs(196)) and (inputs(194)));
    layer0_outputs(5211) <= (inputs(244)) and not (inputs(222));
    layer0_outputs(5212) <= '0';
    layer0_outputs(5213) <= (inputs(58)) and not (inputs(208));
    layer0_outputs(5214) <= (inputs(0)) xor (inputs(55));
    layer0_outputs(5215) <= '1';
    layer0_outputs(5216) <= inputs(180);
    layer0_outputs(5217) <= (inputs(70)) xor (inputs(5));
    layer0_outputs(5218) <= inputs(125);
    layer0_outputs(5219) <= inputs(232);
    layer0_outputs(5220) <= not((inputs(248)) or (inputs(245)));
    layer0_outputs(5221) <= (inputs(196)) xor (inputs(204));
    layer0_outputs(5222) <= (inputs(197)) xor (inputs(74));
    layer0_outputs(5223) <= inputs(224);
    layer0_outputs(5224) <= not((inputs(188)) xor (inputs(95)));
    layer0_outputs(5225) <= (inputs(190)) or (inputs(103));
    layer0_outputs(5226) <= not(inputs(86));
    layer0_outputs(5227) <= (inputs(132)) xor (inputs(227));
    layer0_outputs(5228) <= not(inputs(62)) or (inputs(198));
    layer0_outputs(5229) <= not(inputs(27));
    layer0_outputs(5230) <= inputs(247);
    layer0_outputs(5231) <= (inputs(184)) or (inputs(161));
    layer0_outputs(5232) <= (inputs(105)) and not (inputs(222));
    layer0_outputs(5233) <= not((inputs(213)) xor (inputs(245)));
    layer0_outputs(5234) <= not(inputs(193));
    layer0_outputs(5235) <= not(inputs(39)) or (inputs(154));
    layer0_outputs(5236) <= (inputs(148)) xor (inputs(73));
    layer0_outputs(5237) <= not(inputs(99));
    layer0_outputs(5238) <= inputs(154);
    layer0_outputs(5239) <= (inputs(74)) and not (inputs(136));
    layer0_outputs(5240) <= not((inputs(131)) or (inputs(198)));
    layer0_outputs(5241) <= (inputs(151)) and not (inputs(15));
    layer0_outputs(5242) <= inputs(173);
    layer0_outputs(5243) <= not(inputs(35)) or (inputs(196));
    layer0_outputs(5244) <= not(inputs(215));
    layer0_outputs(5245) <= not((inputs(150)) or (inputs(167)));
    layer0_outputs(5246) <= not((inputs(172)) xor (inputs(206)));
    layer0_outputs(5247) <= not(inputs(229));
    layer0_outputs(5248) <= (inputs(23)) and not (inputs(130));
    layer0_outputs(5249) <= not(inputs(229)) or (inputs(147));
    layer0_outputs(5250) <= not((inputs(203)) or (inputs(179)));
    layer0_outputs(5251) <= not((inputs(254)) xor (inputs(2)));
    layer0_outputs(5252) <= (inputs(87)) xor (inputs(102));
    layer0_outputs(5253) <= (inputs(162)) and not (inputs(2));
    layer0_outputs(5254) <= (inputs(50)) or (inputs(15));
    layer0_outputs(5255) <= (inputs(209)) or (inputs(211));
    layer0_outputs(5256) <= not(inputs(7)) or (inputs(113));
    layer0_outputs(5257) <= inputs(163);
    layer0_outputs(5258) <= not((inputs(177)) or (inputs(80)));
    layer0_outputs(5259) <= (inputs(55)) and not (inputs(0));
    layer0_outputs(5260) <= not((inputs(250)) or (inputs(102)));
    layer0_outputs(5261) <= inputs(83);
    layer0_outputs(5262) <= inputs(9);
    layer0_outputs(5263) <= (inputs(191)) xor (inputs(38));
    layer0_outputs(5264) <= inputs(127);
    layer0_outputs(5265) <= inputs(108);
    layer0_outputs(5266) <= not(inputs(136));
    layer0_outputs(5267) <= not((inputs(96)) xor (inputs(65)));
    layer0_outputs(5268) <= not(inputs(195));
    layer0_outputs(5269) <= not((inputs(164)) or (inputs(192)));
    layer0_outputs(5270) <= not((inputs(209)) xor (inputs(253)));
    layer0_outputs(5271) <= not((inputs(121)) or (inputs(151)));
    layer0_outputs(5272) <= not(inputs(176));
    layer0_outputs(5273) <= (inputs(155)) xor (inputs(136));
    layer0_outputs(5274) <= inputs(99);
    layer0_outputs(5275) <= (inputs(79)) or (inputs(120));
    layer0_outputs(5276) <= not((inputs(24)) xor (inputs(82)));
    layer0_outputs(5277) <= '1';
    layer0_outputs(5278) <= (inputs(208)) xor (inputs(241));
    layer0_outputs(5279) <= (inputs(243)) and not (inputs(13));
    layer0_outputs(5280) <= inputs(114);
    layer0_outputs(5281) <= (inputs(141)) or (inputs(39));
    layer0_outputs(5282) <= not((inputs(106)) and (inputs(99)));
    layer0_outputs(5283) <= not((inputs(253)) or (inputs(6)));
    layer0_outputs(5284) <= not(inputs(17));
    layer0_outputs(5285) <= not(inputs(228)) or (inputs(38));
    layer0_outputs(5286) <= (inputs(240)) xor (inputs(57));
    layer0_outputs(5287) <= not(inputs(5)) or (inputs(184));
    layer0_outputs(5288) <= not(inputs(109)) or (inputs(186));
    layer0_outputs(5289) <= (inputs(53)) or (inputs(72));
    layer0_outputs(5290) <= (inputs(236)) xor (inputs(188));
    layer0_outputs(5291) <= inputs(18);
    layer0_outputs(5292) <= inputs(246);
    layer0_outputs(5293) <= (inputs(197)) xor (inputs(247));
    layer0_outputs(5294) <= inputs(82);
    layer0_outputs(5295) <= inputs(146);
    layer0_outputs(5296) <= (inputs(8)) and not (inputs(160));
    layer0_outputs(5297) <= inputs(13);
    layer0_outputs(5298) <= (inputs(193)) or (inputs(21));
    layer0_outputs(5299) <= not((inputs(73)) or (inputs(170)));
    layer0_outputs(5300) <= inputs(229);
    layer0_outputs(5301) <= inputs(86);
    layer0_outputs(5302) <= not(inputs(41)) or (inputs(203));
    layer0_outputs(5303) <= not((inputs(163)) and (inputs(188)));
    layer0_outputs(5304) <= not(inputs(24)) or (inputs(119));
    layer0_outputs(5305) <= inputs(100);
    layer0_outputs(5306) <= inputs(203);
    layer0_outputs(5307) <= (inputs(116)) and not (inputs(191));
    layer0_outputs(5308) <= (inputs(216)) and not (inputs(74));
    layer0_outputs(5309) <= not(inputs(214)) or (inputs(238));
    layer0_outputs(5310) <= not(inputs(243));
    layer0_outputs(5311) <= not((inputs(88)) xor (inputs(52)));
    layer0_outputs(5312) <= not(inputs(243));
    layer0_outputs(5313) <= not((inputs(45)) or (inputs(121)));
    layer0_outputs(5314) <= not(inputs(178));
    layer0_outputs(5315) <= (inputs(248)) or (inputs(224));
    layer0_outputs(5316) <= (inputs(26)) and not (inputs(174));
    layer0_outputs(5317) <= not(inputs(11));
    layer0_outputs(5318) <= not((inputs(125)) and (inputs(162)));
    layer0_outputs(5319) <= (inputs(148)) or (inputs(67));
    layer0_outputs(5320) <= (inputs(126)) or (inputs(83));
    layer0_outputs(5321) <= not((inputs(235)) or (inputs(170)));
    layer0_outputs(5322) <= not(inputs(218)) or (inputs(181));
    layer0_outputs(5323) <= not(inputs(187)) or (inputs(32));
    layer0_outputs(5324) <= (inputs(248)) or (inputs(65));
    layer0_outputs(5325) <= not((inputs(197)) or (inputs(235)));
    layer0_outputs(5326) <= (inputs(166)) or (inputs(82));
    layer0_outputs(5327) <= not((inputs(239)) xor (inputs(127)));
    layer0_outputs(5328) <= (inputs(190)) and not (inputs(204));
    layer0_outputs(5329) <= not((inputs(239)) or (inputs(141)));
    layer0_outputs(5330) <= inputs(37);
    layer0_outputs(5331) <= not((inputs(82)) or (inputs(99)));
    layer0_outputs(5332) <= not((inputs(98)) xor (inputs(45)));
    layer0_outputs(5333) <= not(inputs(110)) or (inputs(251));
    layer0_outputs(5334) <= '1';
    layer0_outputs(5335) <= (inputs(86)) and (inputs(218));
    layer0_outputs(5336) <= inputs(128);
    layer0_outputs(5337) <= not(inputs(125)) or (inputs(118));
    layer0_outputs(5338) <= (inputs(105)) xor (inputs(15));
    layer0_outputs(5339) <= not(inputs(254));
    layer0_outputs(5340) <= (inputs(233)) and not (inputs(143));
    layer0_outputs(5341) <= inputs(142);
    layer0_outputs(5342) <= (inputs(64)) or (inputs(211));
    layer0_outputs(5343) <= inputs(151);
    layer0_outputs(5344) <= (inputs(92)) or (inputs(128));
    layer0_outputs(5345) <= (inputs(212)) and not (inputs(109));
    layer0_outputs(5346) <= (inputs(232)) or (inputs(220));
    layer0_outputs(5347) <= inputs(131);
    layer0_outputs(5348) <= not(inputs(193)) or (inputs(20));
    layer0_outputs(5349) <= not(inputs(82));
    layer0_outputs(5350) <= not((inputs(200)) or (inputs(234)));
    layer0_outputs(5351) <= not(inputs(83)) or (inputs(135));
    layer0_outputs(5352) <= '1';
    layer0_outputs(5353) <= inputs(229);
    layer0_outputs(5354) <= not(inputs(45));
    layer0_outputs(5355) <= not(inputs(88));
    layer0_outputs(5356) <= not(inputs(124));
    layer0_outputs(5357) <= inputs(189);
    layer0_outputs(5358) <= not((inputs(201)) xor (inputs(102)));
    layer0_outputs(5359) <= (inputs(216)) xor (inputs(132));
    layer0_outputs(5360) <= not((inputs(96)) or (inputs(46)));
    layer0_outputs(5361) <= (inputs(149)) and not (inputs(100));
    layer0_outputs(5362) <= not(inputs(13)) or (inputs(178));
    layer0_outputs(5363) <= inputs(121);
    layer0_outputs(5364) <= (inputs(168)) or (inputs(47));
    layer0_outputs(5365) <= (inputs(154)) and (inputs(147));
    layer0_outputs(5366) <= not((inputs(129)) and (inputs(10)));
    layer0_outputs(5367) <= not((inputs(184)) xor (inputs(22)));
    layer0_outputs(5368) <= not(inputs(172));
    layer0_outputs(5369) <= (inputs(105)) and not (inputs(196));
    layer0_outputs(5370) <= inputs(6);
    layer0_outputs(5371) <= not(inputs(49));
    layer0_outputs(5372) <= (inputs(74)) xor (inputs(22));
    layer0_outputs(5373) <= not(inputs(25));
    layer0_outputs(5374) <= not((inputs(169)) or (inputs(109)));
    layer0_outputs(5375) <= not(inputs(245)) or (inputs(145));
    layer0_outputs(5376) <= inputs(136);
    layer0_outputs(5377) <= not((inputs(179)) and (inputs(163)));
    layer0_outputs(5378) <= (inputs(132)) or (inputs(150));
    layer0_outputs(5379) <= (inputs(231)) and not (inputs(181));
    layer0_outputs(5380) <= (inputs(232)) xor (inputs(8));
    layer0_outputs(5381) <= not(inputs(52)) or (inputs(40));
    layer0_outputs(5382) <= not((inputs(88)) xor (inputs(97)));
    layer0_outputs(5383) <= not((inputs(92)) or (inputs(145)));
    layer0_outputs(5384) <= not((inputs(95)) xor (inputs(254)));
    layer0_outputs(5385) <= inputs(194);
    layer0_outputs(5386) <= (inputs(162)) and not (inputs(236));
    layer0_outputs(5387) <= not((inputs(197)) xor (inputs(243)));
    layer0_outputs(5388) <= not(inputs(101));
    layer0_outputs(5389) <= not(inputs(235));
    layer0_outputs(5390) <= (inputs(35)) and not (inputs(205));
    layer0_outputs(5391) <= inputs(206);
    layer0_outputs(5392) <= (inputs(81)) and not (inputs(136));
    layer0_outputs(5393) <= (inputs(125)) xor (inputs(81));
    layer0_outputs(5394) <= (inputs(65)) and not (inputs(109));
    layer0_outputs(5395) <= (inputs(210)) or (inputs(241));
    layer0_outputs(5396) <= inputs(82);
    layer0_outputs(5397) <= not(inputs(38));
    layer0_outputs(5398) <= not((inputs(61)) or (inputs(65)));
    layer0_outputs(5399) <= (inputs(165)) xor (inputs(179));
    layer0_outputs(5400) <= inputs(243);
    layer0_outputs(5401) <= not(inputs(28));
    layer0_outputs(5402) <= (inputs(212)) and not (inputs(251));
    layer0_outputs(5403) <= (inputs(72)) and not (inputs(131));
    layer0_outputs(5404) <= not(inputs(119));
    layer0_outputs(5405) <= not(inputs(151));
    layer0_outputs(5406) <= inputs(195);
    layer0_outputs(5407) <= inputs(148);
    layer0_outputs(5408) <= not(inputs(107));
    layer0_outputs(5409) <= (inputs(181)) or (inputs(43));
    layer0_outputs(5410) <= not(inputs(163)) or (inputs(170));
    layer0_outputs(5411) <= inputs(105);
    layer0_outputs(5412) <= not(inputs(182));
    layer0_outputs(5413) <= not((inputs(121)) or (inputs(103)));
    layer0_outputs(5414) <= '0';
    layer0_outputs(5415) <= (inputs(58)) or (inputs(19));
    layer0_outputs(5416) <= (inputs(5)) and not (inputs(178));
    layer0_outputs(5417) <= not(inputs(152)) or (inputs(226));
    layer0_outputs(5418) <= not(inputs(149));
    layer0_outputs(5419) <= not((inputs(198)) xor (inputs(64)));
    layer0_outputs(5420) <= (inputs(97)) xor (inputs(56));
    layer0_outputs(5421) <= not((inputs(0)) or (inputs(65)));
    layer0_outputs(5422) <= inputs(68);
    layer0_outputs(5423) <= inputs(59);
    layer0_outputs(5424) <= (inputs(48)) and not (inputs(197));
    layer0_outputs(5425) <= not(inputs(216));
    layer0_outputs(5426) <= (inputs(146)) and not (inputs(255));
    layer0_outputs(5427) <= (inputs(110)) xor (inputs(139));
    layer0_outputs(5428) <= (inputs(252)) or (inputs(207));
    layer0_outputs(5429) <= not(inputs(70)) or (inputs(61));
    layer0_outputs(5430) <= (inputs(94)) xor (inputs(29));
    layer0_outputs(5431) <= not((inputs(91)) or (inputs(65)));
    layer0_outputs(5432) <= not((inputs(0)) xor (inputs(101)));
    layer0_outputs(5433) <= (inputs(208)) or (inputs(209));
    layer0_outputs(5434) <= inputs(183);
    layer0_outputs(5435) <= not(inputs(28));
    layer0_outputs(5436) <= not((inputs(72)) or (inputs(209)));
    layer0_outputs(5437) <= not(inputs(245));
    layer0_outputs(5438) <= not(inputs(215));
    layer0_outputs(5439) <= not(inputs(34));
    layer0_outputs(5440) <= not(inputs(152));
    layer0_outputs(5441) <= not(inputs(109));
    layer0_outputs(5442) <= not((inputs(137)) or (inputs(18)));
    layer0_outputs(5443) <= not((inputs(245)) or (inputs(101)));
    layer0_outputs(5444) <= not((inputs(77)) or (inputs(94)));
    layer0_outputs(5445) <= not(inputs(200)) or (inputs(39));
    layer0_outputs(5446) <= not(inputs(38));
    layer0_outputs(5447) <= (inputs(226)) or (inputs(253));
    layer0_outputs(5448) <= not((inputs(59)) xor (inputs(9)));
    layer0_outputs(5449) <= not((inputs(41)) xor (inputs(7)));
    layer0_outputs(5450) <= not(inputs(35)) or (inputs(128));
    layer0_outputs(5451) <= inputs(214);
    layer0_outputs(5452) <= (inputs(41)) xor (inputs(31));
    layer0_outputs(5453) <= inputs(102);
    layer0_outputs(5454) <= (inputs(61)) and not (inputs(1));
    layer0_outputs(5455) <= inputs(137);
    layer0_outputs(5456) <= (inputs(9)) xor (inputs(31));
    layer0_outputs(5457) <= '0';
    layer0_outputs(5458) <= not(inputs(119));
    layer0_outputs(5459) <= not((inputs(232)) or (inputs(160)));
    layer0_outputs(5460) <= not((inputs(184)) xor (inputs(56)));
    layer0_outputs(5461) <= not(inputs(167));
    layer0_outputs(5462) <= not(inputs(37));
    layer0_outputs(5463) <= not(inputs(122));
    layer0_outputs(5464) <= (inputs(100)) or (inputs(165));
    layer0_outputs(5465) <= not((inputs(156)) xor (inputs(154)));
    layer0_outputs(5466) <= not((inputs(51)) xor (inputs(18)));
    layer0_outputs(5467) <= inputs(137);
    layer0_outputs(5468) <= (inputs(65)) xor (inputs(132));
    layer0_outputs(5469) <= inputs(95);
    layer0_outputs(5470) <= not((inputs(157)) or (inputs(200)));
    layer0_outputs(5471) <= not(inputs(184)) or (inputs(77));
    layer0_outputs(5472) <= (inputs(80)) xor (inputs(17));
    layer0_outputs(5473) <= inputs(246);
    layer0_outputs(5474) <= not(inputs(227)) or (inputs(85));
    layer0_outputs(5475) <= not(inputs(153));
    layer0_outputs(5476) <= not(inputs(233)) or (inputs(136));
    layer0_outputs(5477) <= (inputs(14)) and not (inputs(79));
    layer0_outputs(5478) <= not((inputs(57)) and (inputs(40)));
    layer0_outputs(5479) <= not((inputs(250)) or (inputs(73)));
    layer0_outputs(5480) <= inputs(65);
    layer0_outputs(5481) <= not(inputs(195)) or (inputs(22));
    layer0_outputs(5482) <= not(inputs(113));
    layer0_outputs(5483) <= not((inputs(206)) xor (inputs(159)));
    layer0_outputs(5484) <= (inputs(100)) xor (inputs(191));
    layer0_outputs(5485) <= (inputs(28)) xor (inputs(30));
    layer0_outputs(5486) <= not((inputs(25)) and (inputs(25)));
    layer0_outputs(5487) <= inputs(199);
    layer0_outputs(5488) <= (inputs(159)) and not (inputs(144));
    layer0_outputs(5489) <= (inputs(27)) and not (inputs(93));
    layer0_outputs(5490) <= not(inputs(40));
    layer0_outputs(5491) <= not(inputs(82)) or (inputs(199));
    layer0_outputs(5492) <= not((inputs(162)) or (inputs(251)));
    layer0_outputs(5493) <= (inputs(189)) xor (inputs(234));
    layer0_outputs(5494) <= (inputs(216)) xor (inputs(244));
    layer0_outputs(5495) <= (inputs(102)) xor (inputs(57));
    layer0_outputs(5496) <= not(inputs(102)) or (inputs(55));
    layer0_outputs(5497) <= not((inputs(33)) or (inputs(10)));
    layer0_outputs(5498) <= not((inputs(115)) xor (inputs(29)));
    layer0_outputs(5499) <= not(inputs(195)) or (inputs(130));
    layer0_outputs(5500) <= not(inputs(147)) or (inputs(199));
    layer0_outputs(5501) <= not(inputs(155));
    layer0_outputs(5502) <= not((inputs(174)) xor (inputs(207)));
    layer0_outputs(5503) <= (inputs(109)) xor (inputs(142));
    layer0_outputs(5504) <= inputs(218);
    layer0_outputs(5505) <= (inputs(193)) and not (inputs(246));
    layer0_outputs(5506) <= not(inputs(90));
    layer0_outputs(5507) <= not(inputs(154));
    layer0_outputs(5508) <= (inputs(172)) xor (inputs(2));
    layer0_outputs(5509) <= not(inputs(92));
    layer0_outputs(5510) <= not((inputs(94)) xor (inputs(28)));
    layer0_outputs(5511) <= not((inputs(95)) or (inputs(143)));
    layer0_outputs(5512) <= not(inputs(186));
    layer0_outputs(5513) <= not((inputs(36)) xor (inputs(195)));
    layer0_outputs(5514) <= (inputs(130)) or (inputs(253));
    layer0_outputs(5515) <= not(inputs(195));
    layer0_outputs(5516) <= (inputs(88)) and not (inputs(127));
    layer0_outputs(5517) <= inputs(52);
    layer0_outputs(5518) <= (inputs(59)) xor (inputs(15));
    layer0_outputs(5519) <= not((inputs(72)) or (inputs(191)));
    layer0_outputs(5520) <= not(inputs(52));
    layer0_outputs(5521) <= not(inputs(189));
    layer0_outputs(5522) <= inputs(24);
    layer0_outputs(5523) <= not(inputs(134));
    layer0_outputs(5524) <= (inputs(37)) xor (inputs(180));
    layer0_outputs(5525) <= not(inputs(130));
    layer0_outputs(5526) <= (inputs(182)) or (inputs(64));
    layer0_outputs(5527) <= not((inputs(118)) or (inputs(47)));
    layer0_outputs(5528) <= (inputs(226)) or (inputs(17));
    layer0_outputs(5529) <= not((inputs(21)) or (inputs(245)));
    layer0_outputs(5530) <= not(inputs(204));
    layer0_outputs(5531) <= inputs(30);
    layer0_outputs(5532) <= inputs(193);
    layer0_outputs(5533) <= not(inputs(213));
    layer0_outputs(5534) <= not((inputs(161)) or (inputs(94)));
    layer0_outputs(5535) <= inputs(142);
    layer0_outputs(5536) <= inputs(77);
    layer0_outputs(5537) <= not((inputs(230)) xor (inputs(232)));
    layer0_outputs(5538) <= (inputs(227)) and not (inputs(159));
    layer0_outputs(5539) <= not((inputs(118)) or (inputs(111)));
    layer0_outputs(5540) <= inputs(51);
    layer0_outputs(5541) <= (inputs(12)) xor (inputs(43));
    layer0_outputs(5542) <= inputs(228);
    layer0_outputs(5543) <= (inputs(125)) xor (inputs(61));
    layer0_outputs(5544) <= not(inputs(63)) or (inputs(139));
    layer0_outputs(5545) <= not(inputs(206));
    layer0_outputs(5546) <= (inputs(196)) and not (inputs(45));
    layer0_outputs(5547) <= (inputs(214)) or (inputs(247));
    layer0_outputs(5548) <= not((inputs(193)) or (inputs(40)));
    layer0_outputs(5549) <= not((inputs(33)) xor (inputs(210)));
    layer0_outputs(5550) <= inputs(78);
    layer0_outputs(5551) <= (inputs(95)) xor (inputs(122));
    layer0_outputs(5552) <= inputs(182);
    layer0_outputs(5553) <= not(inputs(228));
    layer0_outputs(5554) <= not((inputs(213)) xor (inputs(244)));
    layer0_outputs(5555) <= (inputs(226)) and not (inputs(48));
    layer0_outputs(5556) <= (inputs(69)) and not (inputs(198));
    layer0_outputs(5557) <= not((inputs(24)) xor (inputs(81)));
    layer0_outputs(5558) <= not(inputs(25));
    layer0_outputs(5559) <= inputs(135);
    layer0_outputs(5560) <= inputs(70);
    layer0_outputs(5561) <= not((inputs(45)) and (inputs(122)));
    layer0_outputs(5562) <= not((inputs(91)) or (inputs(109)));
    layer0_outputs(5563) <= (inputs(121)) xor (inputs(237));
    layer0_outputs(5564) <= inputs(39);
    layer0_outputs(5565) <= not((inputs(198)) xor (inputs(46)));
    layer0_outputs(5566) <= (inputs(186)) or (inputs(237));
    layer0_outputs(5567) <= (inputs(60)) and not (inputs(0));
    layer0_outputs(5568) <= (inputs(15)) and (inputs(151));
    layer0_outputs(5569) <= not((inputs(230)) or (inputs(145)));
    layer0_outputs(5570) <= (inputs(173)) xor (inputs(78));
    layer0_outputs(5571) <= (inputs(137)) or (inputs(21));
    layer0_outputs(5572) <= not((inputs(137)) or (inputs(2)));
    layer0_outputs(5573) <= '0';
    layer0_outputs(5574) <= not(inputs(124)) or (inputs(177));
    layer0_outputs(5575) <= (inputs(170)) xor (inputs(138));
    layer0_outputs(5576) <= not((inputs(159)) and (inputs(33)));
    layer0_outputs(5577) <= not(inputs(12));
    layer0_outputs(5578) <= (inputs(122)) or (inputs(224));
    layer0_outputs(5579) <= inputs(51);
    layer0_outputs(5580) <= inputs(164);
    layer0_outputs(5581) <= not((inputs(190)) or (inputs(214)));
    layer0_outputs(5582) <= not(inputs(223)) or (inputs(126));
    layer0_outputs(5583) <= not((inputs(249)) or (inputs(155)));
    layer0_outputs(5584) <= (inputs(82)) or (inputs(217));
    layer0_outputs(5585) <= inputs(102);
    layer0_outputs(5586) <= (inputs(81)) and (inputs(1));
    layer0_outputs(5587) <= not((inputs(233)) xor (inputs(169)));
    layer0_outputs(5588) <= inputs(26);
    layer0_outputs(5589) <= (inputs(111)) and not (inputs(192));
    layer0_outputs(5590) <= not(inputs(56));
    layer0_outputs(5591) <= not((inputs(161)) xor (inputs(162)));
    layer0_outputs(5592) <= (inputs(140)) or (inputs(11));
    layer0_outputs(5593) <= (inputs(216)) and not (inputs(181));
    layer0_outputs(5594) <= not(inputs(9));
    layer0_outputs(5595) <= (inputs(75)) and not (inputs(191));
    layer0_outputs(5596) <= not(inputs(43));
    layer0_outputs(5597) <= inputs(225);
    layer0_outputs(5598) <= (inputs(103)) and (inputs(102));
    layer0_outputs(5599) <= inputs(99);
    layer0_outputs(5600) <= (inputs(71)) xor (inputs(219));
    layer0_outputs(5601) <= (inputs(114)) xor (inputs(128));
    layer0_outputs(5602) <= inputs(174);
    layer0_outputs(5603) <= not(inputs(102));
    layer0_outputs(5604) <= (inputs(245)) and not (inputs(106));
    layer0_outputs(5605) <= not(inputs(234)) or (inputs(83));
    layer0_outputs(5606) <= not(inputs(78)) or (inputs(32));
    layer0_outputs(5607) <= not(inputs(28));
    layer0_outputs(5608) <= not(inputs(108));
    layer0_outputs(5609) <= not(inputs(147));
    layer0_outputs(5610) <= not((inputs(4)) and (inputs(69)));
    layer0_outputs(5611) <= (inputs(199)) and not (inputs(22));
    layer0_outputs(5612) <= not((inputs(158)) xor (inputs(127)));
    layer0_outputs(5613) <= (inputs(248)) xor (inputs(5));
    layer0_outputs(5614) <= not((inputs(95)) xor (inputs(81)));
    layer0_outputs(5615) <= (inputs(6)) xor (inputs(197));
    layer0_outputs(5616) <= not(inputs(122));
    layer0_outputs(5617) <= inputs(209);
    layer0_outputs(5618) <= (inputs(166)) or (inputs(219));
    layer0_outputs(5619) <= (inputs(12)) and not (inputs(87));
    layer0_outputs(5620) <= not(inputs(43));
    layer0_outputs(5621) <= inputs(150);
    layer0_outputs(5622) <= (inputs(30)) or (inputs(152));
    layer0_outputs(5623) <= not(inputs(241));
    layer0_outputs(5624) <= (inputs(177)) xor (inputs(75));
    layer0_outputs(5625) <= not(inputs(113));
    layer0_outputs(5626) <= inputs(141);
    layer0_outputs(5627) <= not(inputs(141));
    layer0_outputs(5628) <= not((inputs(43)) xor (inputs(228)));
    layer0_outputs(5629) <= not(inputs(168));
    layer0_outputs(5630) <= not(inputs(58));
    layer0_outputs(5631) <= inputs(217);
    layer0_outputs(5632) <= (inputs(225)) or (inputs(251));
    layer0_outputs(5633) <= (inputs(245)) or (inputs(161));
    layer0_outputs(5634) <= (inputs(65)) xor (inputs(35));
    layer0_outputs(5635) <= not((inputs(133)) xor (inputs(130)));
    layer0_outputs(5636) <= not((inputs(139)) or (inputs(30)));
    layer0_outputs(5637) <= not(inputs(116)) or (inputs(242));
    layer0_outputs(5638) <= not((inputs(33)) xor (inputs(238)));
    layer0_outputs(5639) <= (inputs(50)) xor (inputs(75));
    layer0_outputs(5640) <= not((inputs(75)) xor (inputs(44)));
    layer0_outputs(5641) <= (inputs(220)) and (inputs(6));
    layer0_outputs(5642) <= (inputs(111)) and not (inputs(95));
    layer0_outputs(5643) <= not(inputs(104));
    layer0_outputs(5644) <= not(inputs(83)) or (inputs(118));
    layer0_outputs(5645) <= (inputs(59)) and not (inputs(21));
    layer0_outputs(5646) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(5647) <= not((inputs(163)) xor (inputs(70)));
    layer0_outputs(5648) <= not(inputs(206));
    layer0_outputs(5649) <= (inputs(8)) and not (inputs(177));
    layer0_outputs(5650) <= inputs(168);
    layer0_outputs(5651) <= (inputs(94)) and not (inputs(47));
    layer0_outputs(5652) <= (inputs(7)) or (inputs(116));
    layer0_outputs(5653) <= not((inputs(221)) or (inputs(65)));
    layer0_outputs(5654) <= not((inputs(12)) or (inputs(251)));
    layer0_outputs(5655) <= not(inputs(30));
    layer0_outputs(5656) <= inputs(32);
    layer0_outputs(5657) <= not((inputs(223)) or (inputs(247)));
    layer0_outputs(5658) <= not((inputs(111)) xor (inputs(69)));
    layer0_outputs(5659) <= not(inputs(169));
    layer0_outputs(5660) <= (inputs(210)) and not (inputs(170));
    layer0_outputs(5661) <= not((inputs(205)) xor (inputs(78)));
    layer0_outputs(5662) <= not(inputs(245)) or (inputs(152));
    layer0_outputs(5663) <= not(inputs(10)) or (inputs(239));
    layer0_outputs(5664) <= (inputs(163)) and (inputs(216));
    layer0_outputs(5665) <= not((inputs(243)) or (inputs(238)));
    layer0_outputs(5666) <= not((inputs(125)) and (inputs(32)));
    layer0_outputs(5667) <= inputs(120);
    layer0_outputs(5668) <= not(inputs(24)) or (inputs(24));
    layer0_outputs(5669) <= not(inputs(192));
    layer0_outputs(5670) <= not(inputs(129));
    layer0_outputs(5671) <= (inputs(169)) or (inputs(218));
    layer0_outputs(5672) <= not((inputs(136)) or (inputs(152)));
    layer0_outputs(5673) <= not(inputs(50));
    layer0_outputs(5674) <= not(inputs(68));
    layer0_outputs(5675) <= (inputs(18)) xor (inputs(177));
    layer0_outputs(5676) <= not(inputs(125));
    layer0_outputs(5677) <= (inputs(74)) and (inputs(84));
    layer0_outputs(5678) <= (inputs(154)) or (inputs(173));
    layer0_outputs(5679) <= (inputs(23)) and not (inputs(206));
    layer0_outputs(5680) <= not(inputs(218)) or (inputs(237));
    layer0_outputs(5681) <= not((inputs(25)) xor (inputs(207)));
    layer0_outputs(5682) <= inputs(242);
    layer0_outputs(5683) <= not(inputs(98));
    layer0_outputs(5684) <= (inputs(197)) xor (inputs(243));
    layer0_outputs(5685) <= (inputs(133)) and not (inputs(161));
    layer0_outputs(5686) <= (inputs(245)) xor (inputs(51));
    layer0_outputs(5687) <= '0';
    layer0_outputs(5688) <= not((inputs(188)) xor (inputs(195)));
    layer0_outputs(5689) <= (inputs(53)) and (inputs(59));
    layer0_outputs(5690) <= not(inputs(45)) or (inputs(254));
    layer0_outputs(5691) <= not(inputs(248)) or (inputs(10));
    layer0_outputs(5692) <= inputs(82);
    layer0_outputs(5693) <= not((inputs(157)) or (inputs(232)));
    layer0_outputs(5694) <= not((inputs(181)) xor (inputs(31)));
    layer0_outputs(5695) <= not((inputs(51)) and (inputs(233)));
    layer0_outputs(5696) <= (inputs(255)) and (inputs(71));
    layer0_outputs(5697) <= not(inputs(220));
    layer0_outputs(5698) <= not(inputs(100));
    layer0_outputs(5699) <= not(inputs(245));
    layer0_outputs(5700) <= not(inputs(189)) or (inputs(36));
    layer0_outputs(5701) <= (inputs(88)) xor (inputs(145));
    layer0_outputs(5702) <= (inputs(124)) and not (inputs(13));
    layer0_outputs(5703) <= not(inputs(172));
    layer0_outputs(5704) <= not(inputs(227)) or (inputs(252));
    layer0_outputs(5705) <= '0';
    layer0_outputs(5706) <= not(inputs(23));
    layer0_outputs(5707) <= (inputs(28)) xor (inputs(79));
    layer0_outputs(5708) <= (inputs(173)) and not (inputs(217));
    layer0_outputs(5709) <= not((inputs(18)) xor (inputs(6)));
    layer0_outputs(5710) <= (inputs(230)) and (inputs(214));
    layer0_outputs(5711) <= not(inputs(75));
    layer0_outputs(5712) <= (inputs(24)) and not (inputs(217));
    layer0_outputs(5713) <= inputs(31);
    layer0_outputs(5714) <= not(inputs(99)) or (inputs(217));
    layer0_outputs(5715) <= inputs(246);
    layer0_outputs(5716) <= inputs(85);
    layer0_outputs(5717) <= not((inputs(207)) or (inputs(2)));
    layer0_outputs(5718) <= not((inputs(3)) or (inputs(162)));
    layer0_outputs(5719) <= (inputs(97)) and not (inputs(68));
    layer0_outputs(5720) <= not((inputs(98)) xor (inputs(153)));
    layer0_outputs(5721) <= not((inputs(32)) xor (inputs(121)));
    layer0_outputs(5722) <= (inputs(127)) and not (inputs(154));
    layer0_outputs(5723) <= not(inputs(13));
    layer0_outputs(5724) <= (inputs(34)) xor (inputs(36));
    layer0_outputs(5725) <= (inputs(139)) or (inputs(118));
    layer0_outputs(5726) <= inputs(247);
    layer0_outputs(5727) <= (inputs(64)) or (inputs(249));
    layer0_outputs(5728) <= not((inputs(229)) or (inputs(2)));
    layer0_outputs(5729) <= inputs(102);
    layer0_outputs(5730) <= not(inputs(14));
    layer0_outputs(5731) <= inputs(99);
    layer0_outputs(5732) <= not(inputs(51)) or (inputs(192));
    layer0_outputs(5733) <= not((inputs(16)) or (inputs(154)));
    layer0_outputs(5734) <= not((inputs(30)) or (inputs(19)));
    layer0_outputs(5735) <= inputs(248);
    layer0_outputs(5736) <= (inputs(110)) or (inputs(109));
    layer0_outputs(5737) <= not(inputs(74)) or (inputs(162));
    layer0_outputs(5738) <= not(inputs(122));
    layer0_outputs(5739) <= not((inputs(119)) or (inputs(231)));
    layer0_outputs(5740) <= not((inputs(177)) or (inputs(6)));
    layer0_outputs(5741) <= inputs(118);
    layer0_outputs(5742) <= not(inputs(70));
    layer0_outputs(5743) <= (inputs(92)) or (inputs(223));
    layer0_outputs(5744) <= not((inputs(34)) or (inputs(244)));
    layer0_outputs(5745) <= not(inputs(54));
    layer0_outputs(5746) <= not(inputs(249));
    layer0_outputs(5747) <= inputs(40);
    layer0_outputs(5748) <= not(inputs(163)) or (inputs(46));
    layer0_outputs(5749) <= not(inputs(188)) or (inputs(27));
    layer0_outputs(5750) <= (inputs(70)) or (inputs(182));
    layer0_outputs(5751) <= not(inputs(139));
    layer0_outputs(5752) <= inputs(87);
    layer0_outputs(5753) <= not((inputs(80)) xor (inputs(202)));
    layer0_outputs(5754) <= (inputs(108)) and not (inputs(207));
    layer0_outputs(5755) <= (inputs(161)) xor (inputs(180));
    layer0_outputs(5756) <= (inputs(236)) and (inputs(234));
    layer0_outputs(5757) <= (inputs(150)) and not (inputs(223));
    layer0_outputs(5758) <= not((inputs(131)) xor (inputs(32)));
    layer0_outputs(5759) <= not((inputs(245)) xor (inputs(225)));
    layer0_outputs(5760) <= (inputs(114)) or (inputs(217));
    layer0_outputs(5761) <= not((inputs(245)) or (inputs(29)));
    layer0_outputs(5762) <= (inputs(137)) and not (inputs(39));
    layer0_outputs(5763) <= (inputs(232)) or (inputs(191));
    layer0_outputs(5764) <= inputs(119);
    layer0_outputs(5765) <= not(inputs(184)) or (inputs(30));
    layer0_outputs(5766) <= not((inputs(42)) and (inputs(242)));
    layer0_outputs(5767) <= not(inputs(193));
    layer0_outputs(5768) <= not(inputs(42));
    layer0_outputs(5769) <= not((inputs(166)) xor (inputs(123)));
    layer0_outputs(5770) <= not((inputs(50)) xor (inputs(116)));
    layer0_outputs(5771) <= not(inputs(215));
    layer0_outputs(5772) <= inputs(228);
    layer0_outputs(5773) <= not(inputs(136)) or (inputs(126));
    layer0_outputs(5774) <= (inputs(46)) or (inputs(0));
    layer0_outputs(5775) <= inputs(184);
    layer0_outputs(5776) <= (inputs(219)) xor (inputs(121));
    layer0_outputs(5777) <= not(inputs(82));
    layer0_outputs(5778) <= not((inputs(251)) and (inputs(1)));
    layer0_outputs(5779) <= not(inputs(182)) or (inputs(70));
    layer0_outputs(5780) <= not(inputs(182));
    layer0_outputs(5781) <= (inputs(93)) or (inputs(88));
    layer0_outputs(5782) <= not((inputs(240)) xor (inputs(5)));
    layer0_outputs(5783) <= (inputs(134)) and (inputs(39));
    layer0_outputs(5784) <= not((inputs(143)) xor (inputs(239)));
    layer0_outputs(5785) <= not(inputs(104)) or (inputs(144));
    layer0_outputs(5786) <= not((inputs(33)) or (inputs(207)));
    layer0_outputs(5787) <= (inputs(110)) or (inputs(16));
    layer0_outputs(5788) <= not(inputs(231));
    layer0_outputs(5789) <= not((inputs(7)) or (inputs(59)));
    layer0_outputs(5790) <= not((inputs(101)) or (inputs(159)));
    layer0_outputs(5791) <= inputs(145);
    layer0_outputs(5792) <= (inputs(251)) xor (inputs(202));
    layer0_outputs(5793) <= not(inputs(159));
    layer0_outputs(5794) <= (inputs(7)) xor (inputs(170));
    layer0_outputs(5795) <= not(inputs(217)) or (inputs(61));
    layer0_outputs(5796) <= (inputs(152)) or (inputs(142));
    layer0_outputs(5797) <= inputs(221);
    layer0_outputs(5798) <= not(inputs(60)) or (inputs(164));
    layer0_outputs(5799) <= not(inputs(59)) or (inputs(189));
    layer0_outputs(5800) <= (inputs(117)) and not (inputs(123));
    layer0_outputs(5801) <= not((inputs(31)) or (inputs(191)));
    layer0_outputs(5802) <= (inputs(113)) or (inputs(112));
    layer0_outputs(5803) <= (inputs(59)) xor (inputs(27));
    layer0_outputs(5804) <= not((inputs(198)) xor (inputs(182)));
    layer0_outputs(5805) <= (inputs(150)) or (inputs(192));
    layer0_outputs(5806) <= (inputs(57)) or (inputs(48));
    layer0_outputs(5807) <= inputs(167);
    layer0_outputs(5808) <= not((inputs(186)) or (inputs(155)));
    layer0_outputs(5809) <= not((inputs(127)) or (inputs(212)));
    layer0_outputs(5810) <= not(inputs(210));
    layer0_outputs(5811) <= inputs(73);
    layer0_outputs(5812) <= (inputs(122)) or (inputs(11));
    layer0_outputs(5813) <= (inputs(196)) and not (inputs(208));
    layer0_outputs(5814) <= '0';
    layer0_outputs(5815) <= inputs(147);
    layer0_outputs(5816) <= not((inputs(115)) or (inputs(177)));
    layer0_outputs(5817) <= not(inputs(107)) or (inputs(130));
    layer0_outputs(5818) <= not((inputs(64)) xor (inputs(21)));
    layer0_outputs(5819) <= not((inputs(51)) xor (inputs(198)));
    layer0_outputs(5820) <= (inputs(100)) and not (inputs(227));
    layer0_outputs(5821) <= not((inputs(5)) or (inputs(181)));
    layer0_outputs(5822) <= (inputs(69)) or (inputs(11));
    layer0_outputs(5823) <= (inputs(103)) and not (inputs(96));
    layer0_outputs(5824) <= not(inputs(152)) or (inputs(63));
    layer0_outputs(5825) <= '0';
    layer0_outputs(5826) <= (inputs(146)) and not (inputs(254));
    layer0_outputs(5827) <= inputs(180);
    layer0_outputs(5828) <= not((inputs(201)) or (inputs(227)));
    layer0_outputs(5829) <= inputs(11);
    layer0_outputs(5830) <= inputs(89);
    layer0_outputs(5831) <= inputs(229);
    layer0_outputs(5832) <= not((inputs(149)) and (inputs(130)));
    layer0_outputs(5833) <= not(inputs(250)) or (inputs(56));
    layer0_outputs(5834) <= not(inputs(125));
    layer0_outputs(5835) <= (inputs(248)) and not (inputs(149));
    layer0_outputs(5836) <= not((inputs(24)) and (inputs(90)));
    layer0_outputs(5837) <= '1';
    layer0_outputs(5838) <= (inputs(34)) xor (inputs(227));
    layer0_outputs(5839) <= not(inputs(58)) or (inputs(238));
    layer0_outputs(5840) <= inputs(59);
    layer0_outputs(5841) <= (inputs(181)) and not (inputs(125));
    layer0_outputs(5842) <= not((inputs(1)) xor (inputs(247)));
    layer0_outputs(5843) <= inputs(89);
    layer0_outputs(5844) <= '1';
    layer0_outputs(5845) <= not(inputs(219));
    layer0_outputs(5846) <= not(inputs(191)) or (inputs(73));
    layer0_outputs(5847) <= inputs(238);
    layer0_outputs(5848) <= not((inputs(177)) xor (inputs(147)));
    layer0_outputs(5849) <= not((inputs(69)) or (inputs(166)));
    layer0_outputs(5850) <= not(inputs(236));
    layer0_outputs(5851) <= inputs(58);
    layer0_outputs(5852) <= not(inputs(44));
    layer0_outputs(5853) <= inputs(70);
    layer0_outputs(5854) <= not((inputs(31)) xor (inputs(96)));
    layer0_outputs(5855) <= (inputs(91)) or (inputs(220));
    layer0_outputs(5856) <= not(inputs(37));
    layer0_outputs(5857) <= not((inputs(47)) or (inputs(221)));
    layer0_outputs(5858) <= not(inputs(218));
    layer0_outputs(5859) <= not(inputs(61)) or (inputs(96));
    layer0_outputs(5860) <= not(inputs(255));
    layer0_outputs(5861) <= not(inputs(180));
    layer0_outputs(5862) <= not(inputs(209));
    layer0_outputs(5863) <= (inputs(197)) or (inputs(141));
    layer0_outputs(5864) <= not((inputs(131)) or (inputs(253)));
    layer0_outputs(5865) <= inputs(213);
    layer0_outputs(5866) <= (inputs(7)) and not (inputs(110));
    layer0_outputs(5867) <= not(inputs(162));
    layer0_outputs(5868) <= (inputs(141)) xor (inputs(171));
    layer0_outputs(5869) <= (inputs(52)) xor (inputs(22));
    layer0_outputs(5870) <= not(inputs(14));
    layer0_outputs(5871) <= (inputs(187)) and not (inputs(2));
    layer0_outputs(5872) <= not((inputs(178)) and (inputs(172)));
    layer0_outputs(5873) <= not((inputs(90)) xor (inputs(10)));
    layer0_outputs(5874) <= (inputs(123)) xor (inputs(132));
    layer0_outputs(5875) <= not(inputs(73));
    layer0_outputs(5876) <= (inputs(4)) xor (inputs(145));
    layer0_outputs(5877) <= (inputs(174)) and not (inputs(3));
    layer0_outputs(5878) <= (inputs(81)) xor (inputs(235));
    layer0_outputs(5879) <= (inputs(173)) or (inputs(248));
    layer0_outputs(5880) <= (inputs(183)) and not (inputs(69));
    layer0_outputs(5881) <= (inputs(206)) or (inputs(214));
    layer0_outputs(5882) <= (inputs(210)) and (inputs(148));
    layer0_outputs(5883) <= (inputs(206)) or (inputs(135));
    layer0_outputs(5884) <= (inputs(95)) or (inputs(225));
    layer0_outputs(5885) <= inputs(94);
    layer0_outputs(5886) <= (inputs(77)) and not (inputs(223));
    layer0_outputs(5887) <= not((inputs(32)) or (inputs(243)));
    layer0_outputs(5888) <= inputs(136);
    layer0_outputs(5889) <= (inputs(20)) and not (inputs(141));
    layer0_outputs(5890) <= inputs(178);
    layer0_outputs(5891) <= (inputs(100)) xor (inputs(70));
    layer0_outputs(5892) <= not(inputs(248)) or (inputs(1));
    layer0_outputs(5893) <= not(inputs(59));
    layer0_outputs(5894) <= (inputs(74)) and not (inputs(142));
    layer0_outputs(5895) <= (inputs(102)) and not (inputs(232));
    layer0_outputs(5896) <= (inputs(32)) or (inputs(55));
    layer0_outputs(5897) <= (inputs(150)) or (inputs(49));
    layer0_outputs(5898) <= (inputs(116)) and not (inputs(4));
    layer0_outputs(5899) <= inputs(226);
    layer0_outputs(5900) <= inputs(147);
    layer0_outputs(5901) <= (inputs(119)) and not (inputs(20));
    layer0_outputs(5902) <= (inputs(5)) or (inputs(236));
    layer0_outputs(5903) <= inputs(193);
    layer0_outputs(5904) <= (inputs(23)) and not (inputs(149));
    layer0_outputs(5905) <= (inputs(85)) or (inputs(162));
    layer0_outputs(5906) <= not(inputs(22)) or (inputs(254));
    layer0_outputs(5907) <= inputs(10);
    layer0_outputs(5908) <= not(inputs(20));
    layer0_outputs(5909) <= not(inputs(45));
    layer0_outputs(5910) <= not((inputs(157)) or (inputs(193)));
    layer0_outputs(5911) <= (inputs(36)) xor (inputs(185));
    layer0_outputs(5912) <= inputs(123);
    layer0_outputs(5913) <= (inputs(20)) xor (inputs(249));
    layer0_outputs(5914) <= inputs(79);
    layer0_outputs(5915) <= not(inputs(26));
    layer0_outputs(5916) <= not((inputs(6)) or (inputs(138)));
    layer0_outputs(5917) <= inputs(130);
    layer0_outputs(5918) <= not((inputs(40)) and (inputs(215)));
    layer0_outputs(5919) <= (inputs(140)) xor (inputs(117));
    layer0_outputs(5920) <= not(inputs(227));
    layer0_outputs(5921) <= not((inputs(123)) or (inputs(149)));
    layer0_outputs(5922) <= (inputs(225)) and not (inputs(48));
    layer0_outputs(5923) <= not((inputs(139)) or (inputs(51)));
    layer0_outputs(5924) <= (inputs(84)) and not (inputs(150));
    layer0_outputs(5925) <= (inputs(47)) and (inputs(42));
    layer0_outputs(5926) <= inputs(27);
    layer0_outputs(5927) <= (inputs(147)) and not (inputs(0));
    layer0_outputs(5928) <= not((inputs(148)) or (inputs(95)));
    layer0_outputs(5929) <= not(inputs(22)) or (inputs(118));
    layer0_outputs(5930) <= not((inputs(69)) xor (inputs(38)));
    layer0_outputs(5931) <= (inputs(53)) xor (inputs(9));
    layer0_outputs(5932) <= (inputs(6)) and (inputs(151));
    layer0_outputs(5933) <= not(inputs(137));
    layer0_outputs(5934) <= (inputs(207)) and not (inputs(63));
    layer0_outputs(5935) <= (inputs(88)) xor (inputs(238));
    layer0_outputs(5936) <= '0';
    layer0_outputs(5937) <= not((inputs(231)) or (inputs(243)));
    layer0_outputs(5938) <= not((inputs(21)) or (inputs(12)));
    layer0_outputs(5939) <= not((inputs(116)) or (inputs(232)));
    layer0_outputs(5940) <= (inputs(215)) xor (inputs(248));
    layer0_outputs(5941) <= not((inputs(87)) xor (inputs(113)));
    layer0_outputs(5942) <= not((inputs(105)) or (inputs(0)));
    layer0_outputs(5943) <= (inputs(26)) xor (inputs(179));
    layer0_outputs(5944) <= (inputs(183)) and not (inputs(70));
    layer0_outputs(5945) <= not(inputs(163));
    layer0_outputs(5946) <= (inputs(139)) or (inputs(125));
    layer0_outputs(5947) <= (inputs(188)) xor (inputs(205));
    layer0_outputs(5948) <= not(inputs(139));
    layer0_outputs(5949) <= inputs(226);
    layer0_outputs(5950) <= inputs(161);
    layer0_outputs(5951) <= not(inputs(247));
    layer0_outputs(5952) <= (inputs(219)) xor (inputs(154));
    layer0_outputs(5953) <= not((inputs(97)) or (inputs(173)));
    layer0_outputs(5954) <= not(inputs(161));
    layer0_outputs(5955) <= (inputs(52)) and not (inputs(199));
    layer0_outputs(5956) <= (inputs(161)) or (inputs(162));
    layer0_outputs(5957) <= (inputs(218)) and not (inputs(50));
    layer0_outputs(5958) <= (inputs(163)) xor (inputs(74));
    layer0_outputs(5959) <= not((inputs(230)) or (inputs(209)));
    layer0_outputs(5960) <= not(inputs(130));
    layer0_outputs(5961) <= (inputs(223)) xor (inputs(47));
    layer0_outputs(5962) <= not((inputs(152)) or (inputs(149)));
    layer0_outputs(5963) <= '1';
    layer0_outputs(5964) <= (inputs(42)) and not (inputs(33));
    layer0_outputs(5965) <= not((inputs(38)) or (inputs(167)));
    layer0_outputs(5966) <= inputs(176);
    layer0_outputs(5967) <= (inputs(174)) and not (inputs(227));
    layer0_outputs(5968) <= inputs(115);
    layer0_outputs(5969) <= not(inputs(238));
    layer0_outputs(5970) <= not(inputs(160));
    layer0_outputs(5971) <= inputs(66);
    layer0_outputs(5972) <= not(inputs(159)) or (inputs(163));
    layer0_outputs(5973) <= (inputs(39)) or (inputs(183));
    layer0_outputs(5974) <= not(inputs(120));
    layer0_outputs(5975) <= not((inputs(12)) or (inputs(197)));
    layer0_outputs(5976) <= not((inputs(253)) xor (inputs(222)));
    layer0_outputs(5977) <= '0';
    layer0_outputs(5978) <= (inputs(240)) and not (inputs(15));
    layer0_outputs(5979) <= inputs(169);
    layer0_outputs(5980) <= '1';
    layer0_outputs(5981) <= (inputs(176)) xor (inputs(74));
    layer0_outputs(5982) <= not(inputs(59)) or (inputs(35));
    layer0_outputs(5983) <= (inputs(74)) xor (inputs(203));
    layer0_outputs(5984) <= not(inputs(155));
    layer0_outputs(5985) <= (inputs(65)) xor (inputs(71));
    layer0_outputs(5986) <= (inputs(222)) or (inputs(169));
    layer0_outputs(5987) <= inputs(4);
    layer0_outputs(5988) <= not((inputs(242)) xor (inputs(238)));
    layer0_outputs(5989) <= not((inputs(217)) xor (inputs(171)));
    layer0_outputs(5990) <= not((inputs(202)) xor (inputs(85)));
    layer0_outputs(5991) <= not(inputs(119)) or (inputs(127));
    layer0_outputs(5992) <= not((inputs(15)) xor (inputs(227)));
    layer0_outputs(5993) <= (inputs(0)) or (inputs(129));
    layer0_outputs(5994) <= (inputs(243)) and (inputs(119));
    layer0_outputs(5995) <= not(inputs(152)) or (inputs(190));
    layer0_outputs(5996) <= not((inputs(120)) or (inputs(129)));
    layer0_outputs(5997) <= (inputs(0)) xor (inputs(170));
    layer0_outputs(5998) <= not((inputs(117)) xor (inputs(3)));
    layer0_outputs(5999) <= not(inputs(242)) or (inputs(94));
    layer0_outputs(6000) <= (inputs(142)) and not (inputs(254));
    layer0_outputs(6001) <= (inputs(240)) and (inputs(66));
    layer0_outputs(6002) <= not((inputs(198)) xor (inputs(176)));
    layer0_outputs(6003) <= not((inputs(58)) or (inputs(249)));
    layer0_outputs(6004) <= (inputs(215)) and not (inputs(107));
    layer0_outputs(6005) <= (inputs(114)) and not (inputs(49));
    layer0_outputs(6006) <= (inputs(19)) or (inputs(4));
    layer0_outputs(6007) <= not((inputs(134)) xor (inputs(86)));
    layer0_outputs(6008) <= not(inputs(252)) or (inputs(152));
    layer0_outputs(6009) <= (inputs(28)) and not (inputs(139));
    layer0_outputs(6010) <= not(inputs(123));
    layer0_outputs(6011) <= inputs(213);
    layer0_outputs(6012) <= not((inputs(80)) or (inputs(121)));
    layer0_outputs(6013) <= not((inputs(144)) xor (inputs(96)));
    layer0_outputs(6014) <= inputs(180);
    layer0_outputs(6015) <= (inputs(96)) and not (inputs(253));
    layer0_outputs(6016) <= inputs(233);
    layer0_outputs(6017) <= (inputs(157)) and not (inputs(169));
    layer0_outputs(6018) <= inputs(91);
    layer0_outputs(6019) <= inputs(59);
    layer0_outputs(6020) <= (inputs(248)) or (inputs(10));
    layer0_outputs(6021) <= (inputs(187)) or (inputs(9));
    layer0_outputs(6022) <= (inputs(252)) and not (inputs(96));
    layer0_outputs(6023) <= not(inputs(37)) or (inputs(207));
    layer0_outputs(6024) <= not(inputs(233));
    layer0_outputs(6025) <= not(inputs(53));
    layer0_outputs(6026) <= inputs(141);
    layer0_outputs(6027) <= not(inputs(90));
    layer0_outputs(6028) <= not(inputs(146));
    layer0_outputs(6029) <= not((inputs(32)) or (inputs(55)));
    layer0_outputs(6030) <= (inputs(105)) or (inputs(121));
    layer0_outputs(6031) <= not(inputs(166));
    layer0_outputs(6032) <= not((inputs(173)) or (inputs(20)));
    layer0_outputs(6033) <= (inputs(2)) and not (inputs(240));
    layer0_outputs(6034) <= not((inputs(38)) or (inputs(49)));
    layer0_outputs(6035) <= (inputs(20)) and not (inputs(179));
    layer0_outputs(6036) <= (inputs(5)) and not (inputs(220));
    layer0_outputs(6037) <= inputs(40);
    layer0_outputs(6038) <= inputs(34);
    layer0_outputs(6039) <= (inputs(132)) xor (inputs(206));
    layer0_outputs(6040) <= (inputs(145)) xor (inputs(71));
    layer0_outputs(6041) <= not(inputs(196));
    layer0_outputs(6042) <= not((inputs(163)) or (inputs(3)));
    layer0_outputs(6043) <= (inputs(227)) xor (inputs(159));
    layer0_outputs(6044) <= inputs(188);
    layer0_outputs(6045) <= not(inputs(177));
    layer0_outputs(6046) <= not(inputs(11)) or (inputs(156));
    layer0_outputs(6047) <= (inputs(68)) or (inputs(141));
    layer0_outputs(6048) <= not((inputs(76)) xor (inputs(209)));
    layer0_outputs(6049) <= not(inputs(6));
    layer0_outputs(6050) <= inputs(150);
    layer0_outputs(6051) <= not(inputs(41)) or (inputs(94));
    layer0_outputs(6052) <= not(inputs(66)) or (inputs(48));
    layer0_outputs(6053) <= not(inputs(147));
    layer0_outputs(6054) <= not((inputs(113)) or (inputs(201)));
    layer0_outputs(6055) <= inputs(230);
    layer0_outputs(6056) <= not(inputs(171)) or (inputs(26));
    layer0_outputs(6057) <= (inputs(224)) or (inputs(156));
    layer0_outputs(6058) <= (inputs(123)) or (inputs(132));
    layer0_outputs(6059) <= not((inputs(250)) xor (inputs(155)));
    layer0_outputs(6060) <= not(inputs(245));
    layer0_outputs(6061) <= not((inputs(102)) xor (inputs(54)));
    layer0_outputs(6062) <= (inputs(79)) or (inputs(54));
    layer0_outputs(6063) <= not(inputs(182)) or (inputs(81));
    layer0_outputs(6064) <= (inputs(186)) xor (inputs(1));
    layer0_outputs(6065) <= not(inputs(234));
    layer0_outputs(6066) <= not((inputs(125)) xor (inputs(50)));
    layer0_outputs(6067) <= (inputs(174)) and not (inputs(204));
    layer0_outputs(6068) <= not(inputs(198));
    layer0_outputs(6069) <= not(inputs(19));
    layer0_outputs(6070) <= '0';
    layer0_outputs(6071) <= (inputs(115)) and not (inputs(238));
    layer0_outputs(6072) <= not((inputs(190)) or (inputs(195)));
    layer0_outputs(6073) <= (inputs(96)) and not (inputs(193));
    layer0_outputs(6074) <= not((inputs(205)) and (inputs(138)));
    layer0_outputs(6075) <= inputs(146);
    layer0_outputs(6076) <= not(inputs(211)) or (inputs(136));
    layer0_outputs(6077) <= not((inputs(44)) xor (inputs(121)));
    layer0_outputs(6078) <= not((inputs(131)) xor (inputs(100)));
    layer0_outputs(6079) <= (inputs(203)) and not (inputs(95));
    layer0_outputs(6080) <= (inputs(78)) or (inputs(55));
    layer0_outputs(6081) <= (inputs(172)) xor (inputs(152));
    layer0_outputs(6082) <= (inputs(51)) and not (inputs(162));
    layer0_outputs(6083) <= (inputs(236)) xor (inputs(186));
    layer0_outputs(6084) <= inputs(249);
    layer0_outputs(6085) <= (inputs(7)) xor (inputs(10));
    layer0_outputs(6086) <= not(inputs(210));
    layer0_outputs(6087) <= inputs(232);
    layer0_outputs(6088) <= not(inputs(183));
    layer0_outputs(6089) <= not(inputs(89)) or (inputs(67));
    layer0_outputs(6090) <= not((inputs(249)) or (inputs(215)));
    layer0_outputs(6091) <= not(inputs(56));
    layer0_outputs(6092) <= not(inputs(178)) or (inputs(69));
    layer0_outputs(6093) <= not(inputs(115)) or (inputs(78));
    layer0_outputs(6094) <= not((inputs(12)) or (inputs(124)));
    layer0_outputs(6095) <= not(inputs(219)) or (inputs(109));
    layer0_outputs(6096) <= inputs(201);
    layer0_outputs(6097) <= (inputs(45)) xor (inputs(183));
    layer0_outputs(6098) <= not(inputs(113));
    layer0_outputs(6099) <= (inputs(95)) and not (inputs(26));
    layer0_outputs(6100) <= not(inputs(7)) or (inputs(237));
    layer0_outputs(6101) <= not(inputs(235)) or (inputs(94));
    layer0_outputs(6102) <= not(inputs(157));
    layer0_outputs(6103) <= (inputs(165)) and not (inputs(81));
    layer0_outputs(6104) <= not((inputs(98)) or (inputs(86)));
    layer0_outputs(6105) <= not(inputs(154)) or (inputs(52));
    layer0_outputs(6106) <= not(inputs(165)) or (inputs(112));
    layer0_outputs(6107) <= (inputs(33)) or (inputs(227));
    layer0_outputs(6108) <= not((inputs(43)) or (inputs(124)));
    layer0_outputs(6109) <= not(inputs(146));
    layer0_outputs(6110) <= not(inputs(147));
    layer0_outputs(6111) <= not((inputs(40)) and (inputs(42)));
    layer0_outputs(6112) <= '0';
    layer0_outputs(6113) <= not(inputs(235)) or (inputs(114));
    layer0_outputs(6114) <= not((inputs(225)) xor (inputs(148)));
    layer0_outputs(6115) <= (inputs(248)) or (inputs(163));
    layer0_outputs(6116) <= inputs(72);
    layer0_outputs(6117) <= (inputs(212)) and not (inputs(142));
    layer0_outputs(6118) <= (inputs(178)) and not (inputs(72));
    layer0_outputs(6119) <= inputs(188);
    layer0_outputs(6120) <= not(inputs(219));
    layer0_outputs(6121) <= not((inputs(33)) or (inputs(42)));
    layer0_outputs(6122) <= inputs(139);
    layer0_outputs(6123) <= not((inputs(204)) or (inputs(181)));
    layer0_outputs(6124) <= inputs(41);
    layer0_outputs(6125) <= not(inputs(94)) or (inputs(69));
    layer0_outputs(6126) <= not((inputs(56)) or (inputs(122)));
    layer0_outputs(6127) <= (inputs(140)) or (inputs(36));
    layer0_outputs(6128) <= (inputs(175)) and not (inputs(252));
    layer0_outputs(6129) <= not((inputs(226)) or (inputs(35)));
    layer0_outputs(6130) <= not((inputs(124)) xor (inputs(212)));
    layer0_outputs(6131) <= not((inputs(133)) and (inputs(31)));
    layer0_outputs(6132) <= (inputs(23)) and not (inputs(209));
    layer0_outputs(6133) <= (inputs(136)) xor (inputs(167));
    layer0_outputs(6134) <= not(inputs(76));
    layer0_outputs(6135) <= (inputs(67)) or (inputs(179));
    layer0_outputs(6136) <= (inputs(248)) or (inputs(10));
    layer0_outputs(6137) <= not(inputs(189));
    layer0_outputs(6138) <= not(inputs(114));
    layer0_outputs(6139) <= (inputs(207)) xor (inputs(100));
    layer0_outputs(6140) <= not((inputs(223)) xor (inputs(245)));
    layer0_outputs(6141) <= (inputs(93)) and not (inputs(157));
    layer0_outputs(6142) <= not((inputs(254)) and (inputs(69)));
    layer0_outputs(6143) <= not((inputs(55)) or (inputs(17)));
    layer0_outputs(6144) <= (inputs(131)) and not (inputs(207));
    layer0_outputs(6145) <= not(inputs(160)) or (inputs(251));
    layer0_outputs(6146) <= not((inputs(144)) xor (inputs(147)));
    layer0_outputs(6147) <= not((inputs(239)) or (inputs(99)));
    layer0_outputs(6148) <= not((inputs(196)) and (inputs(1)));
    layer0_outputs(6149) <= not(inputs(160));
    layer0_outputs(6150) <= '0';
    layer0_outputs(6151) <= (inputs(30)) or (inputs(104));
    layer0_outputs(6152) <= (inputs(229)) or (inputs(194));
    layer0_outputs(6153) <= (inputs(120)) or (inputs(158));
    layer0_outputs(6154) <= (inputs(2)) and (inputs(237));
    layer0_outputs(6155) <= not(inputs(36)) or (inputs(202));
    layer0_outputs(6156) <= not((inputs(45)) xor (inputs(58)));
    layer0_outputs(6157) <= not((inputs(161)) or (inputs(59)));
    layer0_outputs(6158) <= inputs(204);
    layer0_outputs(6159) <= not(inputs(114));
    layer0_outputs(6160) <= not((inputs(193)) xor (inputs(181)));
    layer0_outputs(6161) <= not((inputs(91)) or (inputs(31)));
    layer0_outputs(6162) <= not((inputs(5)) or (inputs(144)));
    layer0_outputs(6163) <= inputs(170);
    layer0_outputs(6164) <= (inputs(128)) xor (inputs(208));
    layer0_outputs(6165) <= (inputs(146)) and not (inputs(251));
    layer0_outputs(6166) <= (inputs(54)) xor (inputs(225));
    layer0_outputs(6167) <= (inputs(96)) and (inputs(30));
    layer0_outputs(6168) <= (inputs(29)) and not (inputs(224));
    layer0_outputs(6169) <= (inputs(59)) xor (inputs(47));
    layer0_outputs(6170) <= inputs(248);
    layer0_outputs(6171) <= (inputs(94)) and not (inputs(231));
    layer0_outputs(6172) <= not(inputs(232)) or (inputs(95));
    layer0_outputs(6173) <= (inputs(116)) and not (inputs(220));
    layer0_outputs(6174) <= not((inputs(197)) or (inputs(213)));
    layer0_outputs(6175) <= not((inputs(183)) or (inputs(201)));
    layer0_outputs(6176) <= not(inputs(0)) or (inputs(37));
    layer0_outputs(6177) <= not((inputs(219)) xor (inputs(225)));
    layer0_outputs(6178) <= not((inputs(252)) or (inputs(252)));
    layer0_outputs(6179) <= (inputs(164)) and not (inputs(105));
    layer0_outputs(6180) <= (inputs(143)) or (inputs(40));
    layer0_outputs(6181) <= not(inputs(189));
    layer0_outputs(6182) <= not(inputs(237));
    layer0_outputs(6183) <= not((inputs(104)) or (inputs(50)));
    layer0_outputs(6184) <= inputs(122);
    layer0_outputs(6185) <= not((inputs(190)) or (inputs(38)));
    layer0_outputs(6186) <= not((inputs(254)) xor (inputs(142)));
    layer0_outputs(6187) <= not(inputs(154)) or (inputs(174));
    layer0_outputs(6188) <= inputs(145);
    layer0_outputs(6189) <= (inputs(179)) and not (inputs(175));
    layer0_outputs(6190) <= (inputs(250)) or (inputs(252));
    layer0_outputs(6191) <= inputs(190);
    layer0_outputs(6192) <= not(inputs(163));
    layer0_outputs(6193) <= (inputs(180)) and not (inputs(223));
    layer0_outputs(6194) <= not(inputs(198)) or (inputs(158));
    layer0_outputs(6195) <= not((inputs(152)) xor (inputs(105)));
    layer0_outputs(6196) <= (inputs(182)) or (inputs(160));
    layer0_outputs(6197) <= not(inputs(174)) or (inputs(11));
    layer0_outputs(6198) <= (inputs(126)) and (inputs(123));
    layer0_outputs(6199) <= not(inputs(81));
    layer0_outputs(6200) <= not((inputs(155)) or (inputs(54)));
    layer0_outputs(6201) <= not(inputs(236));
    layer0_outputs(6202) <= not((inputs(170)) or (inputs(211)));
    layer0_outputs(6203) <= (inputs(117)) and not (inputs(53));
    layer0_outputs(6204) <= not(inputs(189)) or (inputs(150));
    layer0_outputs(6205) <= not(inputs(192));
    layer0_outputs(6206) <= '0';
    layer0_outputs(6207) <= inputs(220);
    layer0_outputs(6208) <= not(inputs(229));
    layer0_outputs(6209) <= not(inputs(221));
    layer0_outputs(6210) <= (inputs(242)) and (inputs(96));
    layer0_outputs(6211) <= not(inputs(27)) or (inputs(156));
    layer0_outputs(6212) <= not(inputs(60));
    layer0_outputs(6213) <= not(inputs(67)) or (inputs(199));
    layer0_outputs(6214) <= not(inputs(42));
    layer0_outputs(6215) <= not(inputs(38)) or (inputs(129));
    layer0_outputs(6216) <= (inputs(170)) and not (inputs(31));
    layer0_outputs(6217) <= not(inputs(249));
    layer0_outputs(6218) <= not((inputs(222)) xor (inputs(88)));
    layer0_outputs(6219) <= (inputs(179)) or (inputs(219));
    layer0_outputs(6220) <= not(inputs(141));
    layer0_outputs(6221) <= inputs(246);
    layer0_outputs(6222) <= (inputs(129)) and (inputs(65));
    layer0_outputs(6223) <= (inputs(170)) xor (inputs(81));
    layer0_outputs(6224) <= not(inputs(48));
    layer0_outputs(6225) <= not((inputs(235)) xor (inputs(141)));
    layer0_outputs(6226) <= (inputs(41)) and not (inputs(122));
    layer0_outputs(6227) <= (inputs(122)) and (inputs(9));
    layer0_outputs(6228) <= not(inputs(246));
    layer0_outputs(6229) <= (inputs(109)) xor (inputs(108));
    layer0_outputs(6230) <= not((inputs(58)) or (inputs(94)));
    layer0_outputs(6231) <= not((inputs(173)) or (inputs(205)));
    layer0_outputs(6232) <= inputs(87);
    layer0_outputs(6233) <= (inputs(192)) xor (inputs(35));
    layer0_outputs(6234) <= not((inputs(63)) xor (inputs(156)));
    layer0_outputs(6235) <= not((inputs(129)) or (inputs(246)));
    layer0_outputs(6236) <= (inputs(15)) or (inputs(252));
    layer0_outputs(6237) <= (inputs(149)) xor (inputs(38));
    layer0_outputs(6238) <= not(inputs(87));
    layer0_outputs(6239) <= not(inputs(108));
    layer0_outputs(6240) <= not((inputs(224)) or (inputs(24)));
    layer0_outputs(6241) <= not((inputs(185)) or (inputs(111)));
    layer0_outputs(6242) <= not((inputs(54)) or (inputs(79)));
    layer0_outputs(6243) <= (inputs(157)) or (inputs(197));
    layer0_outputs(6244) <= (inputs(253)) or (inputs(150));
    layer0_outputs(6245) <= not((inputs(170)) or (inputs(94)));
    layer0_outputs(6246) <= (inputs(166)) and not (inputs(16));
    layer0_outputs(6247) <= not(inputs(115));
    layer0_outputs(6248) <= not(inputs(57)) or (inputs(198));
    layer0_outputs(6249) <= not(inputs(56));
    layer0_outputs(6250) <= (inputs(137)) xor (inputs(254));
    layer0_outputs(6251) <= not(inputs(249)) or (inputs(66));
    layer0_outputs(6252) <= not(inputs(187)) or (inputs(93));
    layer0_outputs(6253) <= not((inputs(206)) or (inputs(132)));
    layer0_outputs(6254) <= inputs(222);
    layer0_outputs(6255) <= not(inputs(60)) or (inputs(216));
    layer0_outputs(6256) <= (inputs(185)) xor (inputs(232));
    layer0_outputs(6257) <= not((inputs(98)) xor (inputs(47)));
    layer0_outputs(6258) <= (inputs(184)) and not (inputs(134));
    layer0_outputs(6259) <= (inputs(215)) and not (inputs(166));
    layer0_outputs(6260) <= inputs(38);
    layer0_outputs(6261) <= (inputs(253)) or (inputs(199));
    layer0_outputs(6262) <= not(inputs(149)) or (inputs(160));
    layer0_outputs(6263) <= (inputs(211)) and not (inputs(49));
    layer0_outputs(6264) <= (inputs(53)) and not (inputs(207));
    layer0_outputs(6265) <= (inputs(174)) or (inputs(154));
    layer0_outputs(6266) <= not(inputs(174));
    layer0_outputs(6267) <= not((inputs(193)) or (inputs(93)));
    layer0_outputs(6268) <= (inputs(227)) and not (inputs(65));
    layer0_outputs(6269) <= (inputs(113)) or (inputs(30));
    layer0_outputs(6270) <= not(inputs(46));
    layer0_outputs(6271) <= not((inputs(72)) xor (inputs(62)));
    layer0_outputs(6272) <= (inputs(40)) or (inputs(45));
    layer0_outputs(6273) <= not((inputs(20)) xor (inputs(176)));
    layer0_outputs(6274) <= not((inputs(100)) and (inputs(114)));
    layer0_outputs(6275) <= inputs(181);
    layer0_outputs(6276) <= not(inputs(222));
    layer0_outputs(6277) <= not((inputs(214)) or (inputs(130)));
    layer0_outputs(6278) <= inputs(11);
    layer0_outputs(6279) <= (inputs(27)) or (inputs(174));
    layer0_outputs(6280) <= not(inputs(131)) or (inputs(15));
    layer0_outputs(6281) <= inputs(117);
    layer0_outputs(6282) <= (inputs(8)) xor (inputs(100));
    layer0_outputs(6283) <= not(inputs(216));
    layer0_outputs(6284) <= not(inputs(123)) or (inputs(123));
    layer0_outputs(6285) <= not((inputs(23)) xor (inputs(119)));
    layer0_outputs(6286) <= inputs(95);
    layer0_outputs(6287) <= not((inputs(12)) or (inputs(202)));
    layer0_outputs(6288) <= (inputs(249)) and not (inputs(109));
    layer0_outputs(6289) <= not((inputs(215)) or (inputs(10)));
    layer0_outputs(6290) <= not(inputs(39));
    layer0_outputs(6291) <= not(inputs(198));
    layer0_outputs(6292) <= (inputs(147)) or (inputs(172));
    layer0_outputs(6293) <= not((inputs(238)) xor (inputs(120)));
    layer0_outputs(6294) <= (inputs(163)) xor (inputs(165));
    layer0_outputs(6295) <= not(inputs(73));
    layer0_outputs(6296) <= not(inputs(167)) or (inputs(65));
    layer0_outputs(6297) <= not(inputs(132)) or (inputs(174));
    layer0_outputs(6298) <= not((inputs(77)) or (inputs(206)));
    layer0_outputs(6299) <= not(inputs(249)) or (inputs(30));
    layer0_outputs(6300) <= not((inputs(49)) xor (inputs(91)));
    layer0_outputs(6301) <= (inputs(210)) xor (inputs(218));
    layer0_outputs(6302) <= (inputs(15)) or (inputs(158));
    layer0_outputs(6303) <= not(inputs(98));
    layer0_outputs(6304) <= not(inputs(45));
    layer0_outputs(6305) <= not(inputs(255)) or (inputs(190));
    layer0_outputs(6306) <= (inputs(115)) or (inputs(124));
    layer0_outputs(6307) <= (inputs(141)) xor (inputs(0));
    layer0_outputs(6308) <= (inputs(48)) and not (inputs(237));
    layer0_outputs(6309) <= (inputs(105)) or (inputs(108));
    layer0_outputs(6310) <= (inputs(225)) and not (inputs(3));
    layer0_outputs(6311) <= not(inputs(71)) or (inputs(14));
    layer0_outputs(6312) <= not((inputs(245)) xor (inputs(101)));
    layer0_outputs(6313) <= inputs(110);
    layer0_outputs(6314) <= not((inputs(160)) or (inputs(196)));
    layer0_outputs(6315) <= (inputs(42)) or (inputs(101));
    layer0_outputs(6316) <= not((inputs(247)) xor (inputs(184)));
    layer0_outputs(6317) <= not(inputs(100));
    layer0_outputs(6318) <= not(inputs(147)) or (inputs(130));
    layer0_outputs(6319) <= not(inputs(147));
    layer0_outputs(6320) <= not(inputs(133));
    layer0_outputs(6321) <= not((inputs(246)) xor (inputs(233)));
    layer0_outputs(6322) <= not(inputs(242));
    layer0_outputs(6323) <= (inputs(203)) and not (inputs(127));
    layer0_outputs(6324) <= (inputs(183)) or (inputs(237));
    layer0_outputs(6325) <= not(inputs(239));
    layer0_outputs(6326) <= inputs(44);
    layer0_outputs(6327) <= inputs(14);
    layer0_outputs(6328) <= (inputs(191)) and not (inputs(176));
    layer0_outputs(6329) <= not(inputs(116));
    layer0_outputs(6330) <= not(inputs(78));
    layer0_outputs(6331) <= not(inputs(87)) or (inputs(207));
    layer0_outputs(6332) <= not(inputs(59)) or (inputs(12));
    layer0_outputs(6333) <= not((inputs(112)) xor (inputs(86)));
    layer0_outputs(6334) <= not((inputs(169)) or (inputs(104)));
    layer0_outputs(6335) <= not(inputs(189));
    layer0_outputs(6336) <= not((inputs(202)) or (inputs(143)));
    layer0_outputs(6337) <= not(inputs(162));
    layer0_outputs(6338) <= not((inputs(112)) or (inputs(187)));
    layer0_outputs(6339) <= not((inputs(124)) and (inputs(139)));
    layer0_outputs(6340) <= not((inputs(95)) xor (inputs(7)));
    layer0_outputs(6341) <= inputs(211);
    layer0_outputs(6342) <= not(inputs(87)) or (inputs(98));
    layer0_outputs(6343) <= inputs(143);
    layer0_outputs(6344) <= (inputs(240)) or (inputs(211));
    layer0_outputs(6345) <= not(inputs(166));
    layer0_outputs(6346) <= not(inputs(37)) or (inputs(173));
    layer0_outputs(6347) <= (inputs(161)) or (inputs(47));
    layer0_outputs(6348) <= (inputs(42)) and not (inputs(118));
    layer0_outputs(6349) <= (inputs(167)) or (inputs(102));
    layer0_outputs(6350) <= '1';
    layer0_outputs(6351) <= '1';
    layer0_outputs(6352) <= inputs(197);
    layer0_outputs(6353) <= not((inputs(225)) xor (inputs(130)));
    layer0_outputs(6354) <= (inputs(145)) xor (inputs(100));
    layer0_outputs(6355) <= not((inputs(213)) xor (inputs(132)));
    layer0_outputs(6356) <= not((inputs(53)) or (inputs(161)));
    layer0_outputs(6357) <= not((inputs(147)) or (inputs(146)));
    layer0_outputs(6358) <= not((inputs(57)) and (inputs(226)));
    layer0_outputs(6359) <= '0';
    layer0_outputs(6360) <= (inputs(40)) or (inputs(127));
    layer0_outputs(6361) <= inputs(88);
    layer0_outputs(6362) <= inputs(27);
    layer0_outputs(6363) <= not(inputs(67)) or (inputs(47));
    layer0_outputs(6364) <= (inputs(114)) or (inputs(188));
    layer0_outputs(6365) <= not(inputs(238));
    layer0_outputs(6366) <= (inputs(169)) xor (inputs(177));
    layer0_outputs(6367) <= (inputs(38)) and (inputs(172));
    layer0_outputs(6368) <= not((inputs(33)) xor (inputs(238)));
    layer0_outputs(6369) <= not(inputs(147)) or (inputs(20));
    layer0_outputs(6370) <= (inputs(155)) xor (inputs(223));
    layer0_outputs(6371) <= not((inputs(211)) or (inputs(250)));
    layer0_outputs(6372) <= (inputs(118)) xor (inputs(57));
    layer0_outputs(6373) <= not((inputs(145)) or (inputs(212)));
    layer0_outputs(6374) <= (inputs(247)) or (inputs(26));
    layer0_outputs(6375) <= (inputs(130)) or (inputs(96));
    layer0_outputs(6376) <= not(inputs(26));
    layer0_outputs(6377) <= (inputs(126)) xor (inputs(173));
    layer0_outputs(6378) <= (inputs(70)) and not (inputs(46));
    layer0_outputs(6379) <= not((inputs(246)) xor (inputs(32)));
    layer0_outputs(6380) <= (inputs(161)) and (inputs(188));
    layer0_outputs(6381) <= (inputs(219)) and (inputs(48));
    layer0_outputs(6382) <= not(inputs(105));
    layer0_outputs(6383) <= (inputs(29)) xor (inputs(150));
    layer0_outputs(6384) <= not(inputs(237));
    layer0_outputs(6385) <= not((inputs(140)) or (inputs(100)));
    layer0_outputs(6386) <= inputs(216);
    layer0_outputs(6387) <= not(inputs(105)) or (inputs(63));
    layer0_outputs(6388) <= (inputs(23)) and not (inputs(112));
    layer0_outputs(6389) <= not((inputs(63)) xor (inputs(40)));
    layer0_outputs(6390) <= not((inputs(80)) or (inputs(134)));
    layer0_outputs(6391) <= not(inputs(41));
    layer0_outputs(6392) <= not(inputs(157));
    layer0_outputs(6393) <= (inputs(55)) xor (inputs(25));
    layer0_outputs(6394) <= not((inputs(195)) xor (inputs(196)));
    layer0_outputs(6395) <= (inputs(16)) or (inputs(114));
    layer0_outputs(6396) <= inputs(201);
    layer0_outputs(6397) <= not(inputs(239)) or (inputs(250));
    layer0_outputs(6398) <= not(inputs(233));
    layer0_outputs(6399) <= not((inputs(160)) xor (inputs(143)));
    layer0_outputs(6400) <= inputs(38);
    layer0_outputs(6401) <= (inputs(218)) and not (inputs(112));
    layer0_outputs(6402) <= not((inputs(12)) and (inputs(3)));
    layer0_outputs(6403) <= not((inputs(170)) or (inputs(39)));
    layer0_outputs(6404) <= not((inputs(162)) xor (inputs(250)));
    layer0_outputs(6405) <= not(inputs(215)) or (inputs(24));
    layer0_outputs(6406) <= not(inputs(114));
    layer0_outputs(6407) <= inputs(24);
    layer0_outputs(6408) <= not((inputs(126)) or (inputs(11)));
    layer0_outputs(6409) <= not((inputs(73)) or (inputs(145)));
    layer0_outputs(6410) <= not((inputs(187)) xor (inputs(91)));
    layer0_outputs(6411) <= (inputs(16)) or (inputs(56));
    layer0_outputs(6412) <= (inputs(78)) or (inputs(236));
    layer0_outputs(6413) <= not(inputs(118));
    layer0_outputs(6414) <= not((inputs(88)) and (inputs(73)));
    layer0_outputs(6415) <= not(inputs(138));
    layer0_outputs(6416) <= not(inputs(21)) or (inputs(162));
    layer0_outputs(6417) <= not(inputs(251)) or (inputs(110));
    layer0_outputs(6418) <= (inputs(101)) or (inputs(216));
    layer0_outputs(6419) <= not(inputs(110));
    layer0_outputs(6420) <= (inputs(182)) and not (inputs(17));
    layer0_outputs(6421) <= inputs(138);
    layer0_outputs(6422) <= not(inputs(57));
    layer0_outputs(6423) <= not((inputs(199)) xor (inputs(150)));
    layer0_outputs(6424) <= (inputs(139)) and not (inputs(57));
    layer0_outputs(6425) <= not(inputs(79));
    layer0_outputs(6426) <= not(inputs(34)) or (inputs(208));
    layer0_outputs(6427) <= not(inputs(33)) or (inputs(223));
    layer0_outputs(6428) <= (inputs(110)) or (inputs(166));
    layer0_outputs(6429) <= not(inputs(78));
    layer0_outputs(6430) <= not(inputs(74));
    layer0_outputs(6431) <= inputs(22);
    layer0_outputs(6432) <= (inputs(23)) and not (inputs(255));
    layer0_outputs(6433) <= not(inputs(180));
    layer0_outputs(6434) <= inputs(112);
    layer0_outputs(6435) <= (inputs(167)) and not (inputs(115));
    layer0_outputs(6436) <= inputs(96);
    layer0_outputs(6437) <= (inputs(244)) or (inputs(150));
    layer0_outputs(6438) <= (inputs(11)) xor (inputs(177));
    layer0_outputs(6439) <= inputs(230);
    layer0_outputs(6440) <= not(inputs(104)) or (inputs(2));
    layer0_outputs(6441) <= (inputs(7)) xor (inputs(33));
    layer0_outputs(6442) <= (inputs(198)) xor (inputs(61));
    layer0_outputs(6443) <= inputs(242);
    layer0_outputs(6444) <= (inputs(177)) or (inputs(55));
    layer0_outputs(6445) <= not((inputs(120)) and (inputs(155)));
    layer0_outputs(6446) <= (inputs(138)) or (inputs(83));
    layer0_outputs(6447) <= (inputs(140)) and not (inputs(10));
    layer0_outputs(6448) <= (inputs(181)) and not (inputs(53));
    layer0_outputs(6449) <= (inputs(182)) xor (inputs(172));
    layer0_outputs(6450) <= (inputs(192)) or (inputs(0));
    layer0_outputs(6451) <= not((inputs(125)) and (inputs(137)));
    layer0_outputs(6452) <= not(inputs(153)) or (inputs(57));
    layer0_outputs(6453) <= not(inputs(162));
    layer0_outputs(6454) <= not(inputs(243));
    layer0_outputs(6455) <= (inputs(151)) and not (inputs(117));
    layer0_outputs(6456) <= not(inputs(136));
    layer0_outputs(6457) <= (inputs(68)) and not (inputs(191));
    layer0_outputs(6458) <= inputs(1);
    layer0_outputs(6459) <= not(inputs(86));
    layer0_outputs(6460) <= (inputs(249)) or (inputs(215));
    layer0_outputs(6461) <= not(inputs(195)) or (inputs(137));
    layer0_outputs(6462) <= not((inputs(179)) and (inputs(8)));
    layer0_outputs(6463) <= not((inputs(240)) xor (inputs(56)));
    layer0_outputs(6464) <= inputs(208);
    layer0_outputs(6465) <= '0';
    layer0_outputs(6466) <= (inputs(208)) xor (inputs(58));
    layer0_outputs(6467) <= (inputs(198)) xor (inputs(44));
    layer0_outputs(6468) <= not(inputs(195));
    layer0_outputs(6469) <= inputs(149);
    layer0_outputs(6470) <= inputs(185);
    layer0_outputs(6471) <= not(inputs(210));
    layer0_outputs(6472) <= not((inputs(128)) xor (inputs(38)));
    layer0_outputs(6473) <= not((inputs(12)) xor (inputs(197)));
    layer0_outputs(6474) <= not((inputs(102)) or (inputs(215)));
    layer0_outputs(6475) <= (inputs(168)) or (inputs(183));
    layer0_outputs(6476) <= not(inputs(36));
    layer0_outputs(6477) <= not((inputs(33)) xor (inputs(46)));
    layer0_outputs(6478) <= (inputs(191)) xor (inputs(26));
    layer0_outputs(6479) <= (inputs(68)) xor (inputs(58));
    layer0_outputs(6480) <= inputs(8);
    layer0_outputs(6481) <= (inputs(233)) xor (inputs(201));
    layer0_outputs(6482) <= (inputs(40)) and (inputs(145));
    layer0_outputs(6483) <= (inputs(245)) xor (inputs(14));
    layer0_outputs(6484) <= inputs(121);
    layer0_outputs(6485) <= inputs(142);
    layer0_outputs(6486) <= not(inputs(62)) or (inputs(223));
    layer0_outputs(6487) <= not(inputs(212));
    layer0_outputs(6488) <= not(inputs(93));
    layer0_outputs(6489) <= not(inputs(203));
    layer0_outputs(6490) <= (inputs(194)) or (inputs(146));
    layer0_outputs(6491) <= not((inputs(19)) or (inputs(182)));
    layer0_outputs(6492) <= inputs(8);
    layer0_outputs(6493) <= inputs(96);
    layer0_outputs(6494) <= inputs(233);
    layer0_outputs(6495) <= (inputs(45)) and not (inputs(236));
    layer0_outputs(6496) <= not((inputs(200)) or (inputs(122)));
    layer0_outputs(6497) <= not((inputs(98)) and (inputs(178)));
    layer0_outputs(6498) <= (inputs(253)) or (inputs(197));
    layer0_outputs(6499) <= (inputs(191)) or (inputs(163));
    layer0_outputs(6500) <= (inputs(45)) or (inputs(16));
    layer0_outputs(6501) <= not(inputs(244));
    layer0_outputs(6502) <= not(inputs(174)) or (inputs(15));
    layer0_outputs(6503) <= not((inputs(49)) or (inputs(46)));
    layer0_outputs(6504) <= not(inputs(79));
    layer0_outputs(6505) <= inputs(100);
    layer0_outputs(6506) <= (inputs(74)) or (inputs(92));
    layer0_outputs(6507) <= inputs(168);
    layer0_outputs(6508) <= not(inputs(60)) or (inputs(34));
    layer0_outputs(6509) <= not(inputs(55));
    layer0_outputs(6510) <= '1';
    layer0_outputs(6511) <= not(inputs(236));
    layer0_outputs(6512) <= (inputs(0)) or (inputs(99));
    layer0_outputs(6513) <= not((inputs(106)) xor (inputs(223)));
    layer0_outputs(6514) <= (inputs(60)) or (inputs(59));
    layer0_outputs(6515) <= inputs(109);
    layer0_outputs(6516) <= not(inputs(218));
    layer0_outputs(6517) <= '1';
    layer0_outputs(6518) <= not(inputs(42)) or (inputs(241));
    layer0_outputs(6519) <= '0';
    layer0_outputs(6520) <= (inputs(133)) and not (inputs(133));
    layer0_outputs(6521) <= (inputs(74)) xor (inputs(192));
    layer0_outputs(6522) <= not(inputs(226));
    layer0_outputs(6523) <= not(inputs(9)) or (inputs(110));
    layer0_outputs(6524) <= (inputs(213)) xor (inputs(71));
    layer0_outputs(6525) <= not((inputs(203)) or (inputs(173)));
    layer0_outputs(6526) <= not((inputs(53)) or (inputs(73)));
    layer0_outputs(6527) <= (inputs(8)) or (inputs(193));
    layer0_outputs(6528) <= not((inputs(105)) xor (inputs(111)));
    layer0_outputs(6529) <= '1';
    layer0_outputs(6530) <= not(inputs(240)) or (inputs(140));
    layer0_outputs(6531) <= inputs(162);
    layer0_outputs(6532) <= (inputs(54)) or (inputs(98));
    layer0_outputs(6533) <= (inputs(168)) xor (inputs(149));
    layer0_outputs(6534) <= inputs(163);
    layer0_outputs(6535) <= inputs(144);
    layer0_outputs(6536) <= (inputs(118)) xor (inputs(0));
    layer0_outputs(6537) <= (inputs(160)) and (inputs(112));
    layer0_outputs(6538) <= (inputs(38)) and not (inputs(247));
    layer0_outputs(6539) <= not((inputs(70)) and (inputs(250)));
    layer0_outputs(6540) <= inputs(131);
    layer0_outputs(6541) <= (inputs(156)) xor (inputs(68));
    layer0_outputs(6542) <= (inputs(142)) xor (inputs(253));
    layer0_outputs(6543) <= (inputs(181)) or (inputs(226));
    layer0_outputs(6544) <= inputs(63);
    layer0_outputs(6545) <= not(inputs(165));
    layer0_outputs(6546) <= (inputs(243)) and not (inputs(5));
    layer0_outputs(6547) <= not(inputs(134)) or (inputs(197));
    layer0_outputs(6548) <= not(inputs(68)) or (inputs(78));
    layer0_outputs(6549) <= not((inputs(117)) or (inputs(48)));
    layer0_outputs(6550) <= inputs(126);
    layer0_outputs(6551) <= (inputs(103)) and not (inputs(60));
    layer0_outputs(6552) <= inputs(177);
    layer0_outputs(6553) <= inputs(8);
    layer0_outputs(6554) <= (inputs(90)) or (inputs(122));
    layer0_outputs(6555) <= not((inputs(222)) xor (inputs(151)));
    layer0_outputs(6556) <= (inputs(30)) and not (inputs(110));
    layer0_outputs(6557) <= (inputs(252)) and not (inputs(250));
    layer0_outputs(6558) <= (inputs(52)) or (inputs(42));
    layer0_outputs(6559) <= (inputs(229)) and not (inputs(7));
    layer0_outputs(6560) <= not(inputs(120));
    layer0_outputs(6561) <= (inputs(69)) or (inputs(65));
    layer0_outputs(6562) <= (inputs(203)) xor (inputs(184));
    layer0_outputs(6563) <= (inputs(2)) xor (inputs(75));
    layer0_outputs(6564) <= not((inputs(86)) xor (inputs(136)));
    layer0_outputs(6565) <= not((inputs(219)) xor (inputs(248)));
    layer0_outputs(6566) <= (inputs(28)) or (inputs(210));
    layer0_outputs(6567) <= not((inputs(196)) xor (inputs(66)));
    layer0_outputs(6568) <= inputs(85);
    layer0_outputs(6569) <= (inputs(233)) xor (inputs(96));
    layer0_outputs(6570) <= not(inputs(93));
    layer0_outputs(6571) <= inputs(236);
    layer0_outputs(6572) <= not((inputs(29)) or (inputs(191)));
    layer0_outputs(6573) <= (inputs(190)) and not (inputs(251));
    layer0_outputs(6574) <= (inputs(220)) and not (inputs(131));
    layer0_outputs(6575) <= not(inputs(111));
    layer0_outputs(6576) <= (inputs(107)) and not (inputs(249));
    layer0_outputs(6577) <= not(inputs(164));
    layer0_outputs(6578) <= not(inputs(189));
    layer0_outputs(6579) <= not(inputs(226)) or (inputs(118));
    layer0_outputs(6580) <= not((inputs(138)) xor (inputs(200)));
    layer0_outputs(6581) <= not(inputs(127));
    layer0_outputs(6582) <= inputs(219);
    layer0_outputs(6583) <= not((inputs(3)) xor (inputs(7)));
    layer0_outputs(6584) <= (inputs(255)) or (inputs(70));
    layer0_outputs(6585) <= (inputs(41)) and not (inputs(176));
    layer0_outputs(6586) <= inputs(246);
    layer0_outputs(6587) <= not((inputs(230)) or (inputs(95)));
    layer0_outputs(6588) <= not(inputs(129));
    layer0_outputs(6589) <= not((inputs(178)) xor (inputs(247)));
    layer0_outputs(6590) <= not(inputs(231)) or (inputs(156));
    layer0_outputs(6591) <= (inputs(81)) xor (inputs(166));
    layer0_outputs(6592) <= (inputs(135)) xor (inputs(225));
    layer0_outputs(6593) <= not(inputs(165)) or (inputs(158));
    layer0_outputs(6594) <= (inputs(27)) xor (inputs(92));
    layer0_outputs(6595) <= inputs(69);
    layer0_outputs(6596) <= not(inputs(69));
    layer0_outputs(6597) <= (inputs(209)) or (inputs(208));
    layer0_outputs(6598) <= not(inputs(179)) or (inputs(83));
    layer0_outputs(6599) <= inputs(158);
    layer0_outputs(6600) <= inputs(164);
    layer0_outputs(6601) <= (inputs(255)) and not (inputs(234));
    layer0_outputs(6602) <= not(inputs(164));
    layer0_outputs(6603) <= not(inputs(60)) or (inputs(208));
    layer0_outputs(6604) <= not(inputs(188));
    layer0_outputs(6605) <= not((inputs(83)) or (inputs(94)));
    layer0_outputs(6606) <= (inputs(163)) or (inputs(70));
    layer0_outputs(6607) <= not((inputs(13)) or (inputs(18)));
    layer0_outputs(6608) <= (inputs(25)) and (inputs(194));
    layer0_outputs(6609) <= not(inputs(216));
    layer0_outputs(6610) <= (inputs(27)) xor (inputs(199));
    layer0_outputs(6611) <= not(inputs(142)) or (inputs(132));
    layer0_outputs(6612) <= not(inputs(166));
    layer0_outputs(6613) <= not((inputs(68)) or (inputs(183)));
    layer0_outputs(6614) <= not((inputs(176)) xor (inputs(196)));
    layer0_outputs(6615) <= not((inputs(68)) xor (inputs(150)));
    layer0_outputs(6616) <= (inputs(159)) or (inputs(73));
    layer0_outputs(6617) <= not(inputs(3)) or (inputs(132));
    layer0_outputs(6618) <= (inputs(234)) or (inputs(246));
    layer0_outputs(6619) <= (inputs(38)) and not (inputs(158));
    layer0_outputs(6620) <= not(inputs(131)) or (inputs(76));
    layer0_outputs(6621) <= not((inputs(211)) or (inputs(71)));
    layer0_outputs(6622) <= not((inputs(19)) xor (inputs(102)));
    layer0_outputs(6623) <= not((inputs(143)) or (inputs(89)));
    layer0_outputs(6624) <= inputs(218);
    layer0_outputs(6625) <= (inputs(106)) or (inputs(57));
    layer0_outputs(6626) <= not(inputs(42));
    layer0_outputs(6627) <= (inputs(28)) or (inputs(94));
    layer0_outputs(6628) <= not(inputs(14));
    layer0_outputs(6629) <= (inputs(85)) and not (inputs(251));
    layer0_outputs(6630) <= inputs(146);
    layer0_outputs(6631) <= not(inputs(37)) or (inputs(238));
    layer0_outputs(6632) <= (inputs(222)) and not (inputs(2));
    layer0_outputs(6633) <= not(inputs(85)) or (inputs(32));
    layer0_outputs(6634) <= not(inputs(171)) or (inputs(35));
    layer0_outputs(6635) <= (inputs(237)) and not (inputs(15));
    layer0_outputs(6636) <= inputs(212);
    layer0_outputs(6637) <= inputs(151);
    layer0_outputs(6638) <= (inputs(174)) xor (inputs(195));
    layer0_outputs(6639) <= (inputs(116)) xor (inputs(113));
    layer0_outputs(6640) <= inputs(180);
    layer0_outputs(6641) <= not((inputs(3)) or (inputs(211)));
    layer0_outputs(6642) <= not((inputs(182)) xor (inputs(94)));
    layer0_outputs(6643) <= inputs(129);
    layer0_outputs(6644) <= not(inputs(101)) or (inputs(15));
    layer0_outputs(6645) <= inputs(58);
    layer0_outputs(6646) <= not(inputs(149)) or (inputs(21));
    layer0_outputs(6647) <= '1';
    layer0_outputs(6648) <= not(inputs(159));
    layer0_outputs(6649) <= inputs(238);
    layer0_outputs(6650) <= not(inputs(8));
    layer0_outputs(6651) <= not(inputs(237)) or (inputs(156));
    layer0_outputs(6652) <= inputs(220);
    layer0_outputs(6653) <= not((inputs(184)) xor (inputs(180)));
    layer0_outputs(6654) <= (inputs(35)) and not (inputs(227));
    layer0_outputs(6655) <= inputs(130);
    layer0_outputs(6656) <= inputs(253);
    layer0_outputs(6657) <= (inputs(207)) or (inputs(137));
    layer0_outputs(6658) <= inputs(0);
    layer0_outputs(6659) <= not((inputs(58)) or (inputs(64)));
    layer0_outputs(6660) <= not(inputs(87));
    layer0_outputs(6661) <= (inputs(204)) xor (inputs(195));
    layer0_outputs(6662) <= not(inputs(179));
    layer0_outputs(6663) <= inputs(110);
    layer0_outputs(6664) <= not((inputs(218)) xor (inputs(24)));
    layer0_outputs(6665) <= (inputs(75)) xor (inputs(118));
    layer0_outputs(6666) <= inputs(217);
    layer0_outputs(6667) <= (inputs(49)) xor (inputs(80));
    layer0_outputs(6668) <= (inputs(36)) or (inputs(213));
    layer0_outputs(6669) <= not((inputs(155)) or (inputs(16)));
    layer0_outputs(6670) <= (inputs(79)) and (inputs(200));
    layer0_outputs(6671) <= (inputs(58)) or (inputs(114));
    layer0_outputs(6672) <= inputs(35);
    layer0_outputs(6673) <= inputs(108);
    layer0_outputs(6674) <= (inputs(244)) or (inputs(10));
    layer0_outputs(6675) <= not(inputs(137)) or (inputs(20));
    layer0_outputs(6676) <= not(inputs(164));
    layer0_outputs(6677) <= inputs(123);
    layer0_outputs(6678) <= not(inputs(58));
    layer0_outputs(6679) <= '1';
    layer0_outputs(6680) <= not((inputs(199)) xor (inputs(244)));
    layer0_outputs(6681) <= (inputs(164)) or (inputs(61));
    layer0_outputs(6682) <= not((inputs(8)) xor (inputs(210)));
    layer0_outputs(6683) <= not((inputs(202)) or (inputs(47)));
    layer0_outputs(6684) <= (inputs(56)) and not (inputs(160));
    layer0_outputs(6685) <= not(inputs(166)) or (inputs(133));
    layer0_outputs(6686) <= not(inputs(66)) or (inputs(194));
    layer0_outputs(6687) <= not(inputs(133));
    layer0_outputs(6688) <= not((inputs(145)) or (inputs(68)));
    layer0_outputs(6689) <= not(inputs(3));
    layer0_outputs(6690) <= not((inputs(30)) and (inputs(58)));
    layer0_outputs(6691) <= (inputs(131)) and not (inputs(233));
    layer0_outputs(6692) <= (inputs(16)) or (inputs(34));
    layer0_outputs(6693) <= inputs(223);
    layer0_outputs(6694) <= (inputs(197)) and (inputs(169));
    layer0_outputs(6695) <= inputs(100);
    layer0_outputs(6696) <= not(inputs(23));
    layer0_outputs(6697) <= (inputs(48)) and not (inputs(6));
    layer0_outputs(6698) <= not(inputs(230)) or (inputs(133));
    layer0_outputs(6699) <= (inputs(180)) xor (inputs(30));
    layer0_outputs(6700) <= not((inputs(246)) or (inputs(211)));
    layer0_outputs(6701) <= not(inputs(129));
    layer0_outputs(6702) <= (inputs(56)) and not (inputs(47));
    layer0_outputs(6703) <= not((inputs(10)) or (inputs(59)));
    layer0_outputs(6704) <= (inputs(143)) xor (inputs(142));
    layer0_outputs(6705) <= not(inputs(97));
    layer0_outputs(6706) <= not(inputs(181));
    layer0_outputs(6707) <= (inputs(115)) or (inputs(29));
    layer0_outputs(6708) <= (inputs(123)) and not (inputs(144));
    layer0_outputs(6709) <= not(inputs(182));
    layer0_outputs(6710) <= (inputs(136)) or (inputs(151));
    layer0_outputs(6711) <= (inputs(204)) and not (inputs(194));
    layer0_outputs(6712) <= '1';
    layer0_outputs(6713) <= (inputs(115)) or (inputs(131));
    layer0_outputs(6714) <= not(inputs(35));
    layer0_outputs(6715) <= (inputs(100)) xor (inputs(96));
    layer0_outputs(6716) <= (inputs(180)) xor (inputs(135));
    layer0_outputs(6717) <= not(inputs(113)) or (inputs(235));
    layer0_outputs(6718) <= inputs(151);
    layer0_outputs(6719) <= not(inputs(221)) or (inputs(73));
    layer0_outputs(6720) <= (inputs(198)) xor (inputs(63));
    layer0_outputs(6721) <= inputs(89);
    layer0_outputs(6722) <= (inputs(53)) and (inputs(207));
    layer0_outputs(6723) <= (inputs(213)) and not (inputs(130));
    layer0_outputs(6724) <= (inputs(188)) and not (inputs(0));
    layer0_outputs(6725) <= not((inputs(214)) xor (inputs(216)));
    layer0_outputs(6726) <= (inputs(39)) and not (inputs(160));
    layer0_outputs(6727) <= (inputs(248)) and not (inputs(115));
    layer0_outputs(6728) <= not(inputs(25));
    layer0_outputs(6729) <= (inputs(59)) and not (inputs(224));
    layer0_outputs(6730) <= (inputs(117)) xor (inputs(35));
    layer0_outputs(6731) <= not((inputs(125)) or (inputs(127)));
    layer0_outputs(6732) <= not((inputs(123)) xor (inputs(242)));
    layer0_outputs(6733) <= not(inputs(48));
    layer0_outputs(6734) <= inputs(245);
    layer0_outputs(6735) <= (inputs(37)) and (inputs(86));
    layer0_outputs(6736) <= not((inputs(7)) or (inputs(176)));
    layer0_outputs(6737) <= (inputs(208)) and not (inputs(187));
    layer0_outputs(6738) <= not((inputs(132)) xor (inputs(106)));
    layer0_outputs(6739) <= not(inputs(26));
    layer0_outputs(6740) <= (inputs(250)) and not (inputs(141));
    layer0_outputs(6741) <= not((inputs(36)) or (inputs(221)));
    layer0_outputs(6742) <= not((inputs(111)) or (inputs(167)));
    layer0_outputs(6743) <= not((inputs(231)) and (inputs(103)));
    layer0_outputs(6744) <= not(inputs(121));
    layer0_outputs(6745) <= (inputs(108)) xor (inputs(104));
    layer0_outputs(6746) <= not(inputs(14));
    layer0_outputs(6747) <= not(inputs(249));
    layer0_outputs(6748) <= (inputs(195)) and not (inputs(139));
    layer0_outputs(6749) <= (inputs(69)) and (inputs(103));
    layer0_outputs(6750) <= not((inputs(252)) and (inputs(140)));
    layer0_outputs(6751) <= not((inputs(106)) xor (inputs(61)));
    layer0_outputs(6752) <= not((inputs(232)) xor (inputs(204)));
    layer0_outputs(6753) <= (inputs(221)) xor (inputs(190));
    layer0_outputs(6754) <= '1';
    layer0_outputs(6755) <= inputs(166);
    layer0_outputs(6756) <= inputs(243);
    layer0_outputs(6757) <= not(inputs(180));
    layer0_outputs(6758) <= not(inputs(36)) or (inputs(186));
    layer0_outputs(6759) <= not(inputs(82)) or (inputs(215));
    layer0_outputs(6760) <= not(inputs(75));
    layer0_outputs(6761) <= (inputs(112)) or (inputs(171));
    layer0_outputs(6762) <= (inputs(97)) or (inputs(99));
    layer0_outputs(6763) <= (inputs(235)) xor (inputs(101));
    layer0_outputs(6764) <= not((inputs(23)) and (inputs(22)));
    layer0_outputs(6765) <= not((inputs(222)) xor (inputs(154)));
    layer0_outputs(6766) <= '1';
    layer0_outputs(6767) <= (inputs(116)) or (inputs(48));
    layer0_outputs(6768) <= not(inputs(230));
    layer0_outputs(6769) <= inputs(16);
    layer0_outputs(6770) <= (inputs(11)) or (inputs(84));
    layer0_outputs(6771) <= (inputs(110)) and (inputs(30));
    layer0_outputs(6772) <= not(inputs(250)) or (inputs(112));
    layer0_outputs(6773) <= not(inputs(177));
    layer0_outputs(6774) <= (inputs(57)) or (inputs(176));
    layer0_outputs(6775) <= not(inputs(41));
    layer0_outputs(6776) <= not(inputs(173)) or (inputs(8));
    layer0_outputs(6777) <= (inputs(63)) or (inputs(119));
    layer0_outputs(6778) <= not((inputs(47)) xor (inputs(57)));
    layer0_outputs(6779) <= (inputs(140)) and not (inputs(175));
    layer0_outputs(6780) <= not((inputs(178)) xor (inputs(230)));
    layer0_outputs(6781) <= (inputs(193)) and not (inputs(82));
    layer0_outputs(6782) <= not((inputs(160)) or (inputs(242)));
    layer0_outputs(6783) <= (inputs(11)) or (inputs(19));
    layer0_outputs(6784) <= not((inputs(153)) xor (inputs(247)));
    layer0_outputs(6785) <= inputs(227);
    layer0_outputs(6786) <= not((inputs(235)) or (inputs(208)));
    layer0_outputs(6787) <= not(inputs(134)) or (inputs(202));
    layer0_outputs(6788) <= not(inputs(249)) or (inputs(155));
    layer0_outputs(6789) <= (inputs(40)) xor (inputs(38));
    layer0_outputs(6790) <= not((inputs(255)) or (inputs(22)));
    layer0_outputs(6791) <= inputs(206);
    layer0_outputs(6792) <= (inputs(70)) xor (inputs(70));
    layer0_outputs(6793) <= not(inputs(193)) or (inputs(95));
    layer0_outputs(6794) <= not(inputs(228)) or (inputs(28));
    layer0_outputs(6795) <= (inputs(20)) or (inputs(43));
    layer0_outputs(6796) <= not(inputs(167));
    layer0_outputs(6797) <= (inputs(70)) or (inputs(249));
    layer0_outputs(6798) <= inputs(144);
    layer0_outputs(6799) <= not(inputs(194));
    layer0_outputs(6800) <= not((inputs(62)) or (inputs(236)));
    layer0_outputs(6801) <= not(inputs(148));
    layer0_outputs(6802) <= not(inputs(141));
    layer0_outputs(6803) <= not((inputs(114)) and (inputs(15)));
    layer0_outputs(6804) <= not((inputs(240)) or (inputs(123)));
    layer0_outputs(6805) <= (inputs(8)) or (inputs(163));
    layer0_outputs(6806) <= (inputs(162)) and not (inputs(206));
    layer0_outputs(6807) <= (inputs(174)) xor (inputs(225));
    layer0_outputs(6808) <= not(inputs(25));
    layer0_outputs(6809) <= (inputs(202)) or (inputs(76));
    layer0_outputs(6810) <= inputs(167);
    layer0_outputs(6811) <= inputs(197);
    layer0_outputs(6812) <= not(inputs(178));
    layer0_outputs(6813) <= inputs(203);
    layer0_outputs(6814) <= not((inputs(176)) or (inputs(213)));
    layer0_outputs(6815) <= not(inputs(25));
    layer0_outputs(6816) <= (inputs(21)) and (inputs(119));
    layer0_outputs(6817) <= inputs(176);
    layer0_outputs(6818) <= not(inputs(212));
    layer0_outputs(6819) <= not((inputs(42)) or (inputs(248)));
    layer0_outputs(6820) <= (inputs(95)) xor (inputs(250));
    layer0_outputs(6821) <= not(inputs(170)) or (inputs(206));
    layer0_outputs(6822) <= inputs(248);
    layer0_outputs(6823) <= inputs(29);
    layer0_outputs(6824) <= (inputs(105)) and not (inputs(34));
    layer0_outputs(6825) <= not(inputs(25)) or (inputs(120));
    layer0_outputs(6826) <= inputs(164);
    layer0_outputs(6827) <= not((inputs(192)) or (inputs(22)));
    layer0_outputs(6828) <= inputs(244);
    layer0_outputs(6829) <= inputs(211);
    layer0_outputs(6830) <= not(inputs(166));
    layer0_outputs(6831) <= (inputs(148)) and (inputs(21));
    layer0_outputs(6832) <= not(inputs(148));
    layer0_outputs(6833) <= (inputs(74)) and not (inputs(144));
    layer0_outputs(6834) <= not(inputs(247));
    layer0_outputs(6835) <= inputs(115);
    layer0_outputs(6836) <= (inputs(139)) and not (inputs(177));
    layer0_outputs(6837) <= not((inputs(197)) or (inputs(209)));
    layer0_outputs(6838) <= not((inputs(134)) xor (inputs(234)));
    layer0_outputs(6839) <= (inputs(38)) xor (inputs(35));
    layer0_outputs(6840) <= (inputs(121)) and not (inputs(177));
    layer0_outputs(6841) <= (inputs(126)) or (inputs(2));
    layer0_outputs(6842) <= not((inputs(132)) xor (inputs(181)));
    layer0_outputs(6843) <= inputs(0);
    layer0_outputs(6844) <= not(inputs(232)) or (inputs(65));
    layer0_outputs(6845) <= '1';
    layer0_outputs(6846) <= inputs(60);
    layer0_outputs(6847) <= not((inputs(159)) xor (inputs(254)));
    layer0_outputs(6848) <= (inputs(190)) or (inputs(15));
    layer0_outputs(6849) <= not(inputs(203)) or (inputs(15));
    layer0_outputs(6850) <= not(inputs(94)) or (inputs(198));
    layer0_outputs(6851) <= not((inputs(170)) xor (inputs(243)));
    layer0_outputs(6852) <= not((inputs(40)) or (inputs(162)));
    layer0_outputs(6853) <= not(inputs(246));
    layer0_outputs(6854) <= (inputs(209)) or (inputs(159));
    layer0_outputs(6855) <= inputs(166);
    layer0_outputs(6856) <= (inputs(231)) and not (inputs(242));
    layer0_outputs(6857) <= not(inputs(108));
    layer0_outputs(6858) <= not((inputs(158)) xor (inputs(115)));
    layer0_outputs(6859) <= (inputs(63)) and (inputs(111));
    layer0_outputs(6860) <= (inputs(242)) or (inputs(131));
    layer0_outputs(6861) <= not(inputs(98)) or (inputs(159));
    layer0_outputs(6862) <= not((inputs(156)) xor (inputs(46)));
    layer0_outputs(6863) <= not((inputs(8)) xor (inputs(191)));
    layer0_outputs(6864) <= (inputs(87)) and not (inputs(127));
    layer0_outputs(6865) <= not((inputs(250)) xor (inputs(249)));
    layer0_outputs(6866) <= not(inputs(101));
    layer0_outputs(6867) <= (inputs(204)) and not (inputs(6));
    layer0_outputs(6868) <= not((inputs(91)) or (inputs(92)));
    layer0_outputs(6869) <= (inputs(73)) or (inputs(169));
    layer0_outputs(6870) <= not(inputs(229)) or (inputs(78));
    layer0_outputs(6871) <= (inputs(4)) xor (inputs(44));
    layer0_outputs(6872) <= (inputs(10)) or (inputs(255));
    layer0_outputs(6873) <= (inputs(138)) and not (inputs(24));
    layer0_outputs(6874) <= inputs(148);
    layer0_outputs(6875) <= not(inputs(103));
    layer0_outputs(6876) <= not(inputs(231)) or (inputs(110));
    layer0_outputs(6877) <= (inputs(197)) xor (inputs(50));
    layer0_outputs(6878) <= not(inputs(156));
    layer0_outputs(6879) <= not((inputs(122)) or (inputs(254)));
    layer0_outputs(6880) <= not((inputs(195)) or (inputs(55)));
    layer0_outputs(6881) <= not((inputs(156)) or (inputs(107)));
    layer0_outputs(6882) <= (inputs(65)) or (inputs(57));
    layer0_outputs(6883) <= not(inputs(82));
    layer0_outputs(6884) <= (inputs(190)) xor (inputs(22));
    layer0_outputs(6885) <= (inputs(62)) and not (inputs(87));
    layer0_outputs(6886) <= inputs(120);
    layer0_outputs(6887) <= not(inputs(148)) or (inputs(80));
    layer0_outputs(6888) <= not(inputs(41));
    layer0_outputs(6889) <= not((inputs(148)) and (inputs(134)));
    layer0_outputs(6890) <= not(inputs(110));
    layer0_outputs(6891) <= (inputs(126)) or (inputs(172));
    layer0_outputs(6892) <= not(inputs(153));
    layer0_outputs(6893) <= inputs(102);
    layer0_outputs(6894) <= not((inputs(37)) and (inputs(75)));
    layer0_outputs(6895) <= not((inputs(60)) and (inputs(62)));
    layer0_outputs(6896) <= not((inputs(183)) xor (inputs(106)));
    layer0_outputs(6897) <= not((inputs(215)) or (inputs(32)));
    layer0_outputs(6898) <= not((inputs(127)) xor (inputs(92)));
    layer0_outputs(6899) <= not(inputs(241)) or (inputs(36));
    layer0_outputs(6900) <= inputs(99);
    layer0_outputs(6901) <= not(inputs(186)) or (inputs(30));
    layer0_outputs(6902) <= (inputs(160)) and not (inputs(131));
    layer0_outputs(6903) <= not(inputs(7));
    layer0_outputs(6904) <= '0';
    layer0_outputs(6905) <= not((inputs(120)) or (inputs(74)));
    layer0_outputs(6906) <= not(inputs(81));
    layer0_outputs(6907) <= (inputs(107)) xor (inputs(183));
    layer0_outputs(6908) <= (inputs(254)) and not (inputs(242));
    layer0_outputs(6909) <= (inputs(172)) and not (inputs(236));
    layer0_outputs(6910) <= not((inputs(156)) and (inputs(64)));
    layer0_outputs(6911) <= (inputs(109)) xor (inputs(75));
    layer0_outputs(6912) <= '1';
    layer0_outputs(6913) <= inputs(107);
    layer0_outputs(6914) <= (inputs(58)) and (inputs(206));
    layer0_outputs(6915) <= not(inputs(210)) or (inputs(252));
    layer0_outputs(6916) <= (inputs(234)) or (inputs(128));
    layer0_outputs(6917) <= (inputs(59)) xor (inputs(197));
    layer0_outputs(6918) <= (inputs(7)) and not (inputs(146));
    layer0_outputs(6919) <= not(inputs(101));
    layer0_outputs(6920) <= not(inputs(34));
    layer0_outputs(6921) <= not((inputs(46)) or (inputs(224)));
    layer0_outputs(6922) <= not(inputs(49)) or (inputs(119));
    layer0_outputs(6923) <= (inputs(170)) or (inputs(194));
    layer0_outputs(6924) <= (inputs(12)) or (inputs(225));
    layer0_outputs(6925) <= inputs(213);
    layer0_outputs(6926) <= (inputs(9)) or (inputs(219));
    layer0_outputs(6927) <= (inputs(190)) xor (inputs(121));
    layer0_outputs(6928) <= not(inputs(190));
    layer0_outputs(6929) <= (inputs(182)) and not (inputs(8));
    layer0_outputs(6930) <= (inputs(108)) xor (inputs(111));
    layer0_outputs(6931) <= (inputs(140)) and not (inputs(86));
    layer0_outputs(6932) <= inputs(229);
    layer0_outputs(6933) <= not(inputs(70)) or (inputs(180));
    layer0_outputs(6934) <= not((inputs(233)) xor (inputs(101)));
    layer0_outputs(6935) <= not(inputs(217)) or (inputs(40));
    layer0_outputs(6936) <= inputs(86);
    layer0_outputs(6937) <= inputs(9);
    layer0_outputs(6938) <= not((inputs(18)) or (inputs(192)));
    layer0_outputs(6939) <= (inputs(173)) or (inputs(193));
    layer0_outputs(6940) <= not((inputs(239)) or (inputs(220)));
    layer0_outputs(6941) <= not((inputs(154)) or (inputs(163)));
    layer0_outputs(6942) <= not(inputs(128));
    layer0_outputs(6943) <= (inputs(91)) or (inputs(87));
    layer0_outputs(6944) <= inputs(205);
    layer0_outputs(6945) <= not((inputs(187)) or (inputs(253)));
    layer0_outputs(6946) <= not((inputs(74)) or (inputs(18)));
    layer0_outputs(6947) <= not(inputs(144));
    layer0_outputs(6948) <= not(inputs(185)) or (inputs(164));
    layer0_outputs(6949) <= not((inputs(194)) or (inputs(41)));
    layer0_outputs(6950) <= (inputs(59)) and not (inputs(134));
    layer0_outputs(6951) <= (inputs(184)) and not (inputs(57));
    layer0_outputs(6952) <= not((inputs(213)) xor (inputs(212)));
    layer0_outputs(6953) <= (inputs(104)) and not (inputs(149));
    layer0_outputs(6954) <= not(inputs(194));
    layer0_outputs(6955) <= not((inputs(110)) or (inputs(141)));
    layer0_outputs(6956) <= (inputs(219)) xor (inputs(6));
    layer0_outputs(6957) <= inputs(105);
    layer0_outputs(6958) <= not((inputs(175)) or (inputs(134)));
    layer0_outputs(6959) <= not(inputs(117));
    layer0_outputs(6960) <= inputs(216);
    layer0_outputs(6961) <= (inputs(57)) and not (inputs(211));
    layer0_outputs(6962) <= (inputs(245)) xor (inputs(210));
    layer0_outputs(6963) <= not((inputs(19)) xor (inputs(89)));
    layer0_outputs(6964) <= not((inputs(144)) and (inputs(222)));
    layer0_outputs(6965) <= not(inputs(194)) or (inputs(93));
    layer0_outputs(6966) <= inputs(49);
    layer0_outputs(6967) <= not((inputs(251)) or (inputs(56)));
    layer0_outputs(6968) <= not((inputs(203)) or (inputs(131)));
    layer0_outputs(6969) <= '1';
    layer0_outputs(6970) <= not((inputs(169)) or (inputs(128)));
    layer0_outputs(6971) <= not((inputs(90)) and (inputs(99)));
    layer0_outputs(6972) <= not(inputs(90));
    layer0_outputs(6973) <= not(inputs(166));
    layer0_outputs(6974) <= (inputs(50)) or (inputs(119));
    layer0_outputs(6975) <= not((inputs(67)) xor (inputs(85)));
    layer0_outputs(6976) <= not((inputs(12)) or (inputs(242)));
    layer0_outputs(6977) <= not(inputs(199));
    layer0_outputs(6978) <= (inputs(66)) and not (inputs(0));
    layer0_outputs(6979) <= not(inputs(175)) or (inputs(32));
    layer0_outputs(6980) <= not(inputs(69)) or (inputs(175));
    layer0_outputs(6981) <= inputs(251);
    layer0_outputs(6982) <= (inputs(181)) xor (inputs(21));
    layer0_outputs(6983) <= inputs(102);
    layer0_outputs(6984) <= not(inputs(251)) or (inputs(196));
    layer0_outputs(6985) <= not(inputs(1)) or (inputs(113));
    layer0_outputs(6986) <= (inputs(218)) xor (inputs(203));
    layer0_outputs(6987) <= not((inputs(104)) xor (inputs(13)));
    layer0_outputs(6988) <= (inputs(13)) and not (inputs(49));
    layer0_outputs(6989) <= inputs(163);
    layer0_outputs(6990) <= (inputs(34)) xor (inputs(19));
    layer0_outputs(6991) <= inputs(105);
    layer0_outputs(6992) <= not((inputs(176)) and (inputs(161)));
    layer0_outputs(6993) <= (inputs(123)) and (inputs(147));
    layer0_outputs(6994) <= not(inputs(140));
    layer0_outputs(6995) <= not((inputs(124)) xor (inputs(13)));
    layer0_outputs(6996) <= not((inputs(219)) and (inputs(6)));
    layer0_outputs(6997) <= not(inputs(18)) or (inputs(255));
    layer0_outputs(6998) <= not(inputs(233)) or (inputs(129));
    layer0_outputs(6999) <= not((inputs(57)) or (inputs(246)));
    layer0_outputs(7000) <= (inputs(127)) xor (inputs(79));
    layer0_outputs(7001) <= not(inputs(54));
    layer0_outputs(7002) <= (inputs(98)) or (inputs(69));
    layer0_outputs(7003) <= (inputs(155)) or (inputs(2));
    layer0_outputs(7004) <= not((inputs(40)) xor (inputs(213)));
    layer0_outputs(7005) <= inputs(159);
    layer0_outputs(7006) <= (inputs(210)) and not (inputs(16));
    layer0_outputs(7007) <= inputs(122);
    layer0_outputs(7008) <= not(inputs(152));
    layer0_outputs(7009) <= not((inputs(57)) or (inputs(15)));
    layer0_outputs(7010) <= not((inputs(213)) xor (inputs(238)));
    layer0_outputs(7011) <= (inputs(184)) or (inputs(143));
    layer0_outputs(7012) <= not(inputs(185));
    layer0_outputs(7013) <= (inputs(225)) xor (inputs(249));
    layer0_outputs(7014) <= not((inputs(206)) or (inputs(212)));
    layer0_outputs(7015) <= not((inputs(182)) or (inputs(191)));
    layer0_outputs(7016) <= not(inputs(105)) or (inputs(239));
    layer0_outputs(7017) <= not((inputs(51)) xor (inputs(139)));
    layer0_outputs(7018) <= not(inputs(0));
    layer0_outputs(7019) <= not((inputs(192)) xor (inputs(96)));
    layer0_outputs(7020) <= (inputs(225)) xor (inputs(124));
    layer0_outputs(7021) <= not(inputs(116));
    layer0_outputs(7022) <= not(inputs(232));
    layer0_outputs(7023) <= inputs(165);
    layer0_outputs(7024) <= (inputs(6)) or (inputs(166));
    layer0_outputs(7025) <= not(inputs(107)) or (inputs(158));
    layer0_outputs(7026) <= not(inputs(106));
    layer0_outputs(7027) <= not((inputs(218)) and (inputs(34)));
    layer0_outputs(7028) <= inputs(92);
    layer0_outputs(7029) <= inputs(149);
    layer0_outputs(7030) <= not(inputs(133));
    layer0_outputs(7031) <= inputs(140);
    layer0_outputs(7032) <= not((inputs(129)) or (inputs(128)));
    layer0_outputs(7033) <= not(inputs(238)) or (inputs(2));
    layer0_outputs(7034) <= not((inputs(228)) xor (inputs(62)));
    layer0_outputs(7035) <= not(inputs(132));
    layer0_outputs(7036) <= (inputs(173)) or (inputs(6));
    layer0_outputs(7037) <= not((inputs(43)) or (inputs(50)));
    layer0_outputs(7038) <= not(inputs(89));
    layer0_outputs(7039) <= not((inputs(201)) and (inputs(69)));
    layer0_outputs(7040) <= (inputs(60)) and not (inputs(55));
    layer0_outputs(7041) <= (inputs(144)) xor (inputs(205));
    layer0_outputs(7042) <= not(inputs(228)) or (inputs(152));
    layer0_outputs(7043) <= (inputs(124)) or (inputs(15));
    layer0_outputs(7044) <= not(inputs(8));
    layer0_outputs(7045) <= (inputs(6)) or (inputs(1));
    layer0_outputs(7046) <= inputs(104);
    layer0_outputs(7047) <= not((inputs(235)) or (inputs(4)));
    layer0_outputs(7048) <= not((inputs(220)) xor (inputs(252)));
    layer0_outputs(7049) <= (inputs(226)) and not (inputs(174));
    layer0_outputs(7050) <= '1';
    layer0_outputs(7051) <= not(inputs(39));
    layer0_outputs(7052) <= not(inputs(59)) or (inputs(145));
    layer0_outputs(7053) <= not((inputs(73)) xor (inputs(107)));
    layer0_outputs(7054) <= not((inputs(64)) xor (inputs(71)));
    layer0_outputs(7055) <= not((inputs(152)) xor (inputs(169)));
    layer0_outputs(7056) <= not(inputs(231));
    layer0_outputs(7057) <= (inputs(243)) and not (inputs(119));
    layer0_outputs(7058) <= not((inputs(200)) or (inputs(7)));
    layer0_outputs(7059) <= (inputs(251)) and not (inputs(20));
    layer0_outputs(7060) <= '0';
    layer0_outputs(7061) <= not(inputs(228)) or (inputs(1));
    layer0_outputs(7062) <= not(inputs(114));
    layer0_outputs(7063) <= inputs(31);
    layer0_outputs(7064) <= inputs(190);
    layer0_outputs(7065) <= (inputs(211)) and not (inputs(81));
    layer0_outputs(7066) <= '1';
    layer0_outputs(7067) <= (inputs(76)) or (inputs(202));
    layer0_outputs(7068) <= not(inputs(209));
    layer0_outputs(7069) <= (inputs(50)) and not (inputs(180));
    layer0_outputs(7070) <= not(inputs(132)) or (inputs(2));
    layer0_outputs(7071) <= not(inputs(164)) or (inputs(78));
    layer0_outputs(7072) <= '0';
    layer0_outputs(7073) <= inputs(125);
    layer0_outputs(7074) <= not((inputs(70)) or (inputs(222)));
    layer0_outputs(7075) <= inputs(225);
    layer0_outputs(7076) <= (inputs(85)) or (inputs(84));
    layer0_outputs(7077) <= not((inputs(134)) or (inputs(32)));
    layer0_outputs(7078) <= not(inputs(130)) or (inputs(186));
    layer0_outputs(7079) <= not((inputs(225)) or (inputs(151)));
    layer0_outputs(7080) <= not((inputs(73)) xor (inputs(212)));
    layer0_outputs(7081) <= (inputs(22)) and not (inputs(113));
    layer0_outputs(7082) <= inputs(134);
    layer0_outputs(7083) <= (inputs(180)) and not (inputs(224));
    layer0_outputs(7084) <= not(inputs(37)) or (inputs(176));
    layer0_outputs(7085) <= (inputs(144)) xor (inputs(165));
    layer0_outputs(7086) <= (inputs(215)) and not (inputs(46));
    layer0_outputs(7087) <= inputs(129);
    layer0_outputs(7088) <= (inputs(220)) or (inputs(105));
    layer0_outputs(7089) <= not((inputs(17)) or (inputs(147)));
    layer0_outputs(7090) <= (inputs(51)) xor (inputs(234));
    layer0_outputs(7091) <= not(inputs(212));
    layer0_outputs(7092) <= not(inputs(112));
    layer0_outputs(7093) <= (inputs(119)) or (inputs(226));
    layer0_outputs(7094) <= (inputs(76)) and not (inputs(254));
    layer0_outputs(7095) <= not((inputs(32)) xor (inputs(74)));
    layer0_outputs(7096) <= not(inputs(216)) or (inputs(64));
    layer0_outputs(7097) <= (inputs(99)) and not (inputs(180));
    layer0_outputs(7098) <= (inputs(221)) xor (inputs(64));
    layer0_outputs(7099) <= not(inputs(25));
    layer0_outputs(7100) <= not((inputs(179)) or (inputs(162)));
    layer0_outputs(7101) <= not((inputs(186)) or (inputs(3)));
    layer0_outputs(7102) <= (inputs(0)) or (inputs(149));
    layer0_outputs(7103) <= (inputs(201)) xor (inputs(177));
    layer0_outputs(7104) <= not((inputs(196)) xor (inputs(40)));
    layer0_outputs(7105) <= not((inputs(60)) or (inputs(92)));
    layer0_outputs(7106) <= '0';
    layer0_outputs(7107) <= '1';
    layer0_outputs(7108) <= not(inputs(147)) or (inputs(113));
    layer0_outputs(7109) <= (inputs(12)) xor (inputs(220));
    layer0_outputs(7110) <= not((inputs(183)) xor (inputs(130)));
    layer0_outputs(7111) <= not((inputs(99)) and (inputs(62)));
    layer0_outputs(7112) <= inputs(89);
    layer0_outputs(7113) <= inputs(78);
    layer0_outputs(7114) <= '1';
    layer0_outputs(7115) <= (inputs(119)) or (inputs(105));
    layer0_outputs(7116) <= not(inputs(122));
    layer0_outputs(7117) <= (inputs(198)) xor (inputs(199));
    layer0_outputs(7118) <= inputs(137);
    layer0_outputs(7119) <= (inputs(121)) or (inputs(189));
    layer0_outputs(7120) <= (inputs(224)) and not (inputs(50));
    layer0_outputs(7121) <= not((inputs(180)) xor (inputs(93)));
    layer0_outputs(7122) <= not(inputs(45));
    layer0_outputs(7123) <= not((inputs(51)) and (inputs(105)));
    layer0_outputs(7124) <= not((inputs(169)) and (inputs(187)));
    layer0_outputs(7125) <= inputs(249);
    layer0_outputs(7126) <= (inputs(253)) and not (inputs(175));
    layer0_outputs(7127) <= (inputs(242)) or (inputs(195));
    layer0_outputs(7128) <= inputs(178);
    layer0_outputs(7129) <= (inputs(155)) and not (inputs(208));
    layer0_outputs(7130) <= (inputs(131)) or (inputs(87));
    layer0_outputs(7131) <= inputs(192);
    layer0_outputs(7132) <= not((inputs(239)) or (inputs(40)));
    layer0_outputs(7133) <= (inputs(24)) xor (inputs(177));
    layer0_outputs(7134) <= not(inputs(152));
    layer0_outputs(7135) <= not((inputs(230)) or (inputs(175)));
    layer0_outputs(7136) <= not(inputs(246)) or (inputs(134));
    layer0_outputs(7137) <= (inputs(66)) and not (inputs(95));
    layer0_outputs(7138) <= (inputs(205)) xor (inputs(33));
    layer0_outputs(7139) <= '0';
    layer0_outputs(7140) <= not((inputs(249)) or (inputs(228)));
    layer0_outputs(7141) <= (inputs(239)) or (inputs(173));
    layer0_outputs(7142) <= not((inputs(239)) xor (inputs(175)));
    layer0_outputs(7143) <= inputs(180);
    layer0_outputs(7144) <= not(inputs(130)) or (inputs(132));
    layer0_outputs(7145) <= inputs(21);
    layer0_outputs(7146) <= (inputs(246)) or (inputs(68));
    layer0_outputs(7147) <= (inputs(23)) and (inputs(151));
    layer0_outputs(7148) <= not(inputs(76)) or (inputs(4));
    layer0_outputs(7149) <= (inputs(211)) and not (inputs(110));
    layer0_outputs(7150) <= not(inputs(99)) or (inputs(54));
    layer0_outputs(7151) <= not(inputs(233));
    layer0_outputs(7152) <= not(inputs(153)) or (inputs(235));
    layer0_outputs(7153) <= inputs(197);
    layer0_outputs(7154) <= (inputs(115)) or (inputs(126));
    layer0_outputs(7155) <= not(inputs(170)) or (inputs(217));
    layer0_outputs(7156) <= not((inputs(166)) xor (inputs(136)));
    layer0_outputs(7157) <= not(inputs(188));
    layer0_outputs(7158) <= inputs(212);
    layer0_outputs(7159) <= inputs(77);
    layer0_outputs(7160) <= not((inputs(157)) or (inputs(154)));
    layer0_outputs(7161) <= (inputs(162)) xor (inputs(0));
    layer0_outputs(7162) <= (inputs(148)) xor (inputs(63));
    layer0_outputs(7163) <= (inputs(154)) or (inputs(179));
    layer0_outputs(7164) <= not(inputs(76));
    layer0_outputs(7165) <= (inputs(106)) or (inputs(129));
    layer0_outputs(7166) <= not(inputs(230)) or (inputs(70));
    layer0_outputs(7167) <= (inputs(88)) and not (inputs(52));
    layer0_outputs(7168) <= not(inputs(40));
    layer0_outputs(7169) <= '0';
    layer0_outputs(7170) <= not(inputs(110));
    layer0_outputs(7171) <= not(inputs(219));
    layer0_outputs(7172) <= not((inputs(50)) or (inputs(24)));
    layer0_outputs(7173) <= not((inputs(35)) or (inputs(43)));
    layer0_outputs(7174) <= not((inputs(207)) or (inputs(37)));
    layer0_outputs(7175) <= not(inputs(50));
    layer0_outputs(7176) <= not(inputs(151)) or (inputs(223));
    layer0_outputs(7177) <= not(inputs(83));
    layer0_outputs(7178) <= not(inputs(51)) or (inputs(58));
    layer0_outputs(7179) <= inputs(26);
    layer0_outputs(7180) <= not(inputs(105)) or (inputs(157));
    layer0_outputs(7181) <= '1';
    layer0_outputs(7182) <= inputs(168);
    layer0_outputs(7183) <= not(inputs(162));
    layer0_outputs(7184) <= not(inputs(245)) or (inputs(91));
    layer0_outputs(7185) <= not((inputs(6)) or (inputs(62)));
    layer0_outputs(7186) <= (inputs(86)) xor (inputs(116));
    layer0_outputs(7187) <= inputs(165);
    layer0_outputs(7188) <= inputs(236);
    layer0_outputs(7189) <= inputs(210);
    layer0_outputs(7190) <= (inputs(55)) and not (inputs(49));
    layer0_outputs(7191) <= inputs(186);
    layer0_outputs(7192) <= not((inputs(100)) xor (inputs(147)));
    layer0_outputs(7193) <= not(inputs(22));
    layer0_outputs(7194) <= not(inputs(92)) or (inputs(241));
    layer0_outputs(7195) <= (inputs(104)) or (inputs(227));
    layer0_outputs(7196) <= inputs(27);
    layer0_outputs(7197) <= inputs(104);
    layer0_outputs(7198) <= (inputs(247)) and not (inputs(18));
    layer0_outputs(7199) <= inputs(128);
    layer0_outputs(7200) <= (inputs(219)) or (inputs(4));
    layer0_outputs(7201) <= not(inputs(27));
    layer0_outputs(7202) <= (inputs(135)) and not (inputs(163));
    layer0_outputs(7203) <= (inputs(22)) and not (inputs(63));
    layer0_outputs(7204) <= not(inputs(14)) or (inputs(127));
    layer0_outputs(7205) <= not((inputs(235)) xor (inputs(229)));
    layer0_outputs(7206) <= not(inputs(166));
    layer0_outputs(7207) <= (inputs(64)) or (inputs(159));
    layer0_outputs(7208) <= not((inputs(13)) or (inputs(218)));
    layer0_outputs(7209) <= not((inputs(171)) or (inputs(85)));
    layer0_outputs(7210) <= not((inputs(7)) or (inputs(51)));
    layer0_outputs(7211) <= (inputs(90)) and not (inputs(252));
    layer0_outputs(7212) <= (inputs(46)) xor (inputs(68));
    layer0_outputs(7213) <= (inputs(26)) xor (inputs(23));
    layer0_outputs(7214) <= (inputs(121)) and (inputs(246));
    layer0_outputs(7215) <= inputs(78);
    layer0_outputs(7216) <= not((inputs(252)) xor (inputs(187)));
    layer0_outputs(7217) <= (inputs(189)) and not (inputs(34));
    layer0_outputs(7218) <= '1';
    layer0_outputs(7219) <= not(inputs(209));
    layer0_outputs(7220) <= not(inputs(23)) or (inputs(173));
    layer0_outputs(7221) <= (inputs(250)) xor (inputs(138));
    layer0_outputs(7222) <= (inputs(63)) and not (inputs(216));
    layer0_outputs(7223) <= inputs(82);
    layer0_outputs(7224) <= '1';
    layer0_outputs(7225) <= not((inputs(81)) or (inputs(46)));
    layer0_outputs(7226) <= inputs(244);
    layer0_outputs(7227) <= '0';
    layer0_outputs(7228) <= not((inputs(150)) xor (inputs(62)));
    layer0_outputs(7229) <= (inputs(124)) or (inputs(124));
    layer0_outputs(7230) <= (inputs(148)) xor (inputs(142));
    layer0_outputs(7231) <= inputs(89);
    layer0_outputs(7232) <= (inputs(108)) and (inputs(171));
    layer0_outputs(7233) <= not(inputs(44)) or (inputs(160));
    layer0_outputs(7234) <= inputs(55);
    layer0_outputs(7235) <= not((inputs(104)) or (inputs(118)));
    layer0_outputs(7236) <= not(inputs(170)) or (inputs(241));
    layer0_outputs(7237) <= not((inputs(28)) xor (inputs(70)));
    layer0_outputs(7238) <= inputs(23);
    layer0_outputs(7239) <= (inputs(88)) and not (inputs(34));
    layer0_outputs(7240) <= not((inputs(135)) xor (inputs(110)));
    layer0_outputs(7241) <= inputs(239);
    layer0_outputs(7242) <= '1';
    layer0_outputs(7243) <= not((inputs(76)) or (inputs(62)));
    layer0_outputs(7244) <= not((inputs(161)) or (inputs(196)));
    layer0_outputs(7245) <= (inputs(162)) or (inputs(192));
    layer0_outputs(7246) <= not((inputs(88)) xor (inputs(186)));
    layer0_outputs(7247) <= (inputs(54)) or (inputs(148));
    layer0_outputs(7248) <= (inputs(86)) xor (inputs(255));
    layer0_outputs(7249) <= not(inputs(254));
    layer0_outputs(7250) <= (inputs(235)) and not (inputs(112));
    layer0_outputs(7251) <= not((inputs(172)) or (inputs(219)));
    layer0_outputs(7252) <= inputs(43);
    layer0_outputs(7253) <= not(inputs(71)) or (inputs(107));
    layer0_outputs(7254) <= inputs(145);
    layer0_outputs(7255) <= (inputs(181)) and not (inputs(65));
    layer0_outputs(7256) <= not(inputs(25));
    layer0_outputs(7257) <= '0';
    layer0_outputs(7258) <= inputs(40);
    layer0_outputs(7259) <= (inputs(70)) and not (inputs(1));
    layer0_outputs(7260) <= (inputs(190)) or (inputs(76));
    layer0_outputs(7261) <= (inputs(69)) and not (inputs(15));
    layer0_outputs(7262) <= (inputs(138)) and not (inputs(52));
    layer0_outputs(7263) <= inputs(210);
    layer0_outputs(7264) <= inputs(117);
    layer0_outputs(7265) <= inputs(233);
    layer0_outputs(7266) <= not(inputs(178));
    layer0_outputs(7267) <= inputs(83);
    layer0_outputs(7268) <= inputs(110);
    layer0_outputs(7269) <= inputs(19);
    layer0_outputs(7270) <= (inputs(194)) or (inputs(224));
    layer0_outputs(7271) <= (inputs(8)) and not (inputs(147));
    layer0_outputs(7272) <= (inputs(45)) and not (inputs(17));
    layer0_outputs(7273) <= not(inputs(38)) or (inputs(185));
    layer0_outputs(7274) <= not((inputs(219)) or (inputs(175)));
    layer0_outputs(7275) <= not(inputs(238));
    layer0_outputs(7276) <= inputs(113);
    layer0_outputs(7277) <= (inputs(177)) or (inputs(170));
    layer0_outputs(7278) <= not(inputs(199)) or (inputs(29));
    layer0_outputs(7279) <= (inputs(216)) and not (inputs(49));
    layer0_outputs(7280) <= (inputs(48)) and not (inputs(3));
    layer0_outputs(7281) <= (inputs(140)) and not (inputs(49));
    layer0_outputs(7282) <= inputs(244);
    layer0_outputs(7283) <= inputs(34);
    layer0_outputs(7284) <= inputs(145);
    layer0_outputs(7285) <= not((inputs(28)) xor (inputs(176)));
    layer0_outputs(7286) <= not(inputs(60));
    layer0_outputs(7287) <= inputs(41);
    layer0_outputs(7288) <= not((inputs(199)) or (inputs(17)));
    layer0_outputs(7289) <= not(inputs(48));
    layer0_outputs(7290) <= not((inputs(174)) or (inputs(156)));
    layer0_outputs(7291) <= not(inputs(102));
    layer0_outputs(7292) <= (inputs(82)) and not (inputs(40));
    layer0_outputs(7293) <= not((inputs(14)) or (inputs(236)));
    layer0_outputs(7294) <= not(inputs(230));
    layer0_outputs(7295) <= (inputs(210)) and not (inputs(252));
    layer0_outputs(7296) <= not((inputs(152)) or (inputs(211)));
    layer0_outputs(7297) <= not(inputs(100));
    layer0_outputs(7298) <= not(inputs(114));
    layer0_outputs(7299) <= (inputs(154)) xor (inputs(201));
    layer0_outputs(7300) <= not(inputs(135));
    layer0_outputs(7301) <= inputs(56);
    layer0_outputs(7302) <= (inputs(16)) or (inputs(212));
    layer0_outputs(7303) <= (inputs(75)) or (inputs(95));
    layer0_outputs(7304) <= (inputs(153)) and not (inputs(195));
    layer0_outputs(7305) <= (inputs(157)) and not (inputs(28));
    layer0_outputs(7306) <= not((inputs(30)) or (inputs(29)));
    layer0_outputs(7307) <= not((inputs(33)) or (inputs(19)));
    layer0_outputs(7308) <= (inputs(54)) and not (inputs(148));
    layer0_outputs(7309) <= not((inputs(93)) xor (inputs(189)));
    layer0_outputs(7310) <= not((inputs(80)) xor (inputs(20)));
    layer0_outputs(7311) <= (inputs(35)) xor (inputs(39));
    layer0_outputs(7312) <= not(inputs(21));
    layer0_outputs(7313) <= (inputs(130)) or (inputs(6));
    layer0_outputs(7314) <= inputs(39);
    layer0_outputs(7315) <= '1';
    layer0_outputs(7316) <= not(inputs(251));
    layer0_outputs(7317) <= not(inputs(57)) or (inputs(222));
    layer0_outputs(7318) <= not(inputs(137)) or (inputs(80));
    layer0_outputs(7319) <= inputs(105);
    layer0_outputs(7320) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(7321) <= not(inputs(229));
    layer0_outputs(7322) <= not(inputs(36)) or (inputs(196));
    layer0_outputs(7323) <= (inputs(43)) xor (inputs(71));
    layer0_outputs(7324) <= not((inputs(153)) xor (inputs(144)));
    layer0_outputs(7325) <= (inputs(180)) and not (inputs(216));
    layer0_outputs(7326) <= (inputs(101)) and not (inputs(3));
    layer0_outputs(7327) <= not(inputs(145));
    layer0_outputs(7328) <= not((inputs(35)) or (inputs(101)));
    layer0_outputs(7329) <= not((inputs(35)) or (inputs(21)));
    layer0_outputs(7330) <= (inputs(74)) and not (inputs(230));
    layer0_outputs(7331) <= not((inputs(79)) or (inputs(73)));
    layer0_outputs(7332) <= (inputs(99)) and not (inputs(241));
    layer0_outputs(7333) <= '1';
    layer0_outputs(7334) <= not(inputs(229));
    layer0_outputs(7335) <= not(inputs(107)) or (inputs(212));
    layer0_outputs(7336) <= not((inputs(69)) xor (inputs(170)));
    layer0_outputs(7337) <= not((inputs(213)) or (inputs(36)));
    layer0_outputs(7338) <= not((inputs(237)) or (inputs(47)));
    layer0_outputs(7339) <= not((inputs(161)) or (inputs(82)));
    layer0_outputs(7340) <= not((inputs(203)) and (inputs(241)));
    layer0_outputs(7341) <= not((inputs(171)) xor (inputs(97)));
    layer0_outputs(7342) <= (inputs(49)) xor (inputs(7));
    layer0_outputs(7343) <= inputs(190);
    layer0_outputs(7344) <= inputs(110);
    layer0_outputs(7345) <= not((inputs(175)) or (inputs(115)));
    layer0_outputs(7346) <= not((inputs(94)) or (inputs(191)));
    layer0_outputs(7347) <= inputs(167);
    layer0_outputs(7348) <= not((inputs(83)) or (inputs(191)));
    layer0_outputs(7349) <= inputs(174);
    layer0_outputs(7350) <= inputs(206);
    layer0_outputs(7351) <= not((inputs(126)) or (inputs(197)));
    layer0_outputs(7352) <= (inputs(75)) and not (inputs(185));
    layer0_outputs(7353) <= inputs(85);
    layer0_outputs(7354) <= not((inputs(224)) or (inputs(149)));
    layer0_outputs(7355) <= not(inputs(182));
    layer0_outputs(7356) <= not((inputs(41)) xor (inputs(43)));
    layer0_outputs(7357) <= not((inputs(4)) xor (inputs(42)));
    layer0_outputs(7358) <= not(inputs(231)) or (inputs(4));
    layer0_outputs(7359) <= not(inputs(130));
    layer0_outputs(7360) <= not((inputs(74)) or (inputs(66)));
    layer0_outputs(7361) <= (inputs(172)) xor (inputs(197));
    layer0_outputs(7362) <= not((inputs(6)) xor (inputs(58)));
    layer0_outputs(7363) <= not((inputs(93)) and (inputs(200)));
    layer0_outputs(7364) <= '0';
    layer0_outputs(7365) <= (inputs(78)) or (inputs(51));
    layer0_outputs(7366) <= (inputs(93)) and not (inputs(121));
    layer0_outputs(7367) <= inputs(218);
    layer0_outputs(7368) <= inputs(169);
    layer0_outputs(7369) <= not(inputs(217));
    layer0_outputs(7370) <= not(inputs(119));
    layer0_outputs(7371) <= (inputs(166)) xor (inputs(176));
    layer0_outputs(7372) <= not(inputs(145)) or (inputs(196));
    layer0_outputs(7373) <= (inputs(226)) xor (inputs(170));
    layer0_outputs(7374) <= (inputs(165)) and not (inputs(78));
    layer0_outputs(7375) <= inputs(128);
    layer0_outputs(7376) <= (inputs(243)) and not (inputs(69));
    layer0_outputs(7377) <= inputs(102);
    layer0_outputs(7378) <= not((inputs(206)) xor (inputs(146)));
    layer0_outputs(7379) <= not(inputs(99));
    layer0_outputs(7380) <= not((inputs(36)) and (inputs(35)));
    layer0_outputs(7381) <= (inputs(181)) and (inputs(22));
    layer0_outputs(7382) <= not((inputs(101)) or (inputs(122)));
    layer0_outputs(7383) <= (inputs(101)) and not (inputs(163));
    layer0_outputs(7384) <= '1';
    layer0_outputs(7385) <= (inputs(87)) xor (inputs(84));
    layer0_outputs(7386) <= not((inputs(71)) or (inputs(72)));
    layer0_outputs(7387) <= not(inputs(126)) or (inputs(15));
    layer0_outputs(7388) <= not((inputs(44)) xor (inputs(247)));
    layer0_outputs(7389) <= not(inputs(58)) or (inputs(254));
    layer0_outputs(7390) <= (inputs(145)) or (inputs(13));
    layer0_outputs(7391) <= not((inputs(16)) xor (inputs(84)));
    layer0_outputs(7392) <= not((inputs(168)) or (inputs(222)));
    layer0_outputs(7393) <= not(inputs(146)) or (inputs(124));
    layer0_outputs(7394) <= not((inputs(31)) or (inputs(92)));
    layer0_outputs(7395) <= not(inputs(163));
    layer0_outputs(7396) <= (inputs(98)) or (inputs(140));
    layer0_outputs(7397) <= (inputs(74)) or (inputs(43));
    layer0_outputs(7398) <= (inputs(197)) xor (inputs(193));
    layer0_outputs(7399) <= inputs(98);
    layer0_outputs(7400) <= not(inputs(200));
    layer0_outputs(7401) <= (inputs(247)) or (inputs(230));
    layer0_outputs(7402) <= (inputs(189)) and not (inputs(103));
    layer0_outputs(7403) <= not(inputs(236)) or (inputs(185));
    layer0_outputs(7404) <= not(inputs(153));
    layer0_outputs(7405) <= inputs(81);
    layer0_outputs(7406) <= (inputs(44)) and not (inputs(190));
    layer0_outputs(7407) <= not(inputs(150));
    layer0_outputs(7408) <= (inputs(108)) and not (inputs(191));
    layer0_outputs(7409) <= inputs(128);
    layer0_outputs(7410) <= inputs(25);
    layer0_outputs(7411) <= not((inputs(180)) or (inputs(208)));
    layer0_outputs(7412) <= (inputs(187)) and not (inputs(129));
    layer0_outputs(7413) <= (inputs(158)) or (inputs(37));
    layer0_outputs(7414) <= '0';
    layer0_outputs(7415) <= not(inputs(213));
    layer0_outputs(7416) <= (inputs(45)) xor (inputs(73));
    layer0_outputs(7417) <= '1';
    layer0_outputs(7418) <= not(inputs(30)) or (inputs(225));
    layer0_outputs(7419) <= not(inputs(170));
    layer0_outputs(7420) <= not((inputs(3)) or (inputs(1)));
    layer0_outputs(7421) <= not(inputs(134)) or (inputs(156));
    layer0_outputs(7422) <= not(inputs(164));
    layer0_outputs(7423) <= not((inputs(8)) xor (inputs(45)));
    layer0_outputs(7424) <= (inputs(44)) and not (inputs(216));
    layer0_outputs(7425) <= (inputs(30)) or (inputs(10));
    layer0_outputs(7426) <= (inputs(235)) and not (inputs(130));
    layer0_outputs(7427) <= (inputs(28)) xor (inputs(23));
    layer0_outputs(7428) <= (inputs(181)) and not (inputs(188));
    layer0_outputs(7429) <= (inputs(205)) xor (inputs(192));
    layer0_outputs(7430) <= not((inputs(248)) or (inputs(22)));
    layer0_outputs(7431) <= (inputs(144)) or (inputs(57));
    layer0_outputs(7432) <= not((inputs(243)) or (inputs(150)));
    layer0_outputs(7433) <= (inputs(17)) and not (inputs(144));
    layer0_outputs(7434) <= (inputs(33)) and (inputs(209));
    layer0_outputs(7435) <= not(inputs(171));
    layer0_outputs(7436) <= (inputs(78)) xor (inputs(34));
    layer0_outputs(7437) <= not(inputs(43)) or (inputs(86));
    layer0_outputs(7438) <= not(inputs(15)) or (inputs(222));
    layer0_outputs(7439) <= not((inputs(1)) xor (inputs(16)));
    layer0_outputs(7440) <= not(inputs(113));
    layer0_outputs(7441) <= not(inputs(67)) or (inputs(137));
    layer0_outputs(7442) <= (inputs(60)) xor (inputs(67));
    layer0_outputs(7443) <= not(inputs(117)) or (inputs(197));
    layer0_outputs(7444) <= (inputs(19)) xor (inputs(63));
    layer0_outputs(7445) <= (inputs(54)) and not (inputs(254));
    layer0_outputs(7446) <= not((inputs(239)) xor (inputs(81)));
    layer0_outputs(7447) <= not(inputs(203));
    layer0_outputs(7448) <= '0';
    layer0_outputs(7449) <= not(inputs(219));
    layer0_outputs(7450) <= not(inputs(134));
    layer0_outputs(7451) <= not(inputs(10));
    layer0_outputs(7452) <= not(inputs(84));
    layer0_outputs(7453) <= not(inputs(86));
    layer0_outputs(7454) <= not((inputs(171)) or (inputs(155)));
    layer0_outputs(7455) <= not(inputs(111));
    layer0_outputs(7456) <= not((inputs(229)) and (inputs(102)));
    layer0_outputs(7457) <= not(inputs(103));
    layer0_outputs(7458) <= inputs(26);
    layer0_outputs(7459) <= inputs(35);
    layer0_outputs(7460) <= inputs(168);
    layer0_outputs(7461) <= '1';
    layer0_outputs(7462) <= (inputs(149)) xor (inputs(89));
    layer0_outputs(7463) <= (inputs(54)) or (inputs(7));
    layer0_outputs(7464) <= inputs(86);
    layer0_outputs(7465) <= inputs(227);
    layer0_outputs(7466) <= not((inputs(73)) xor (inputs(70)));
    layer0_outputs(7467) <= (inputs(107)) xor (inputs(93));
    layer0_outputs(7468) <= not(inputs(158));
    layer0_outputs(7469) <= not((inputs(10)) and (inputs(155)));
    layer0_outputs(7470) <= (inputs(195)) and not (inputs(81));
    layer0_outputs(7471) <= not((inputs(8)) or (inputs(82)));
    layer0_outputs(7472) <= not((inputs(223)) xor (inputs(209)));
    layer0_outputs(7473) <= not((inputs(22)) and (inputs(22)));
    layer0_outputs(7474) <= not(inputs(254)) or (inputs(1));
    layer0_outputs(7475) <= (inputs(193)) xor (inputs(12));
    layer0_outputs(7476) <= (inputs(140)) xor (inputs(159));
    layer0_outputs(7477) <= not((inputs(150)) or (inputs(206)));
    layer0_outputs(7478) <= not(inputs(6)) or (inputs(146));
    layer0_outputs(7479) <= (inputs(40)) and not (inputs(165));
    layer0_outputs(7480) <= not(inputs(31)) or (inputs(70));
    layer0_outputs(7481) <= '0';
    layer0_outputs(7482) <= '1';
    layer0_outputs(7483) <= (inputs(108)) and not (inputs(237));
    layer0_outputs(7484) <= inputs(249);
    layer0_outputs(7485) <= (inputs(127)) and not (inputs(201));
    layer0_outputs(7486) <= not(inputs(202)) or (inputs(114));
    layer0_outputs(7487) <= not(inputs(11));
    layer0_outputs(7488) <= (inputs(33)) or (inputs(246));
    layer0_outputs(7489) <= (inputs(139)) and not (inputs(60));
    layer0_outputs(7490) <= not(inputs(12));
    layer0_outputs(7491) <= (inputs(16)) and (inputs(153));
    layer0_outputs(7492) <= (inputs(227)) or (inputs(189));
    layer0_outputs(7493) <= not(inputs(134));
    layer0_outputs(7494) <= (inputs(204)) or (inputs(169));
    layer0_outputs(7495) <= inputs(84);
    layer0_outputs(7496) <= (inputs(126)) or (inputs(27));
    layer0_outputs(7497) <= inputs(210);
    layer0_outputs(7498) <= not(inputs(26));
    layer0_outputs(7499) <= inputs(122);
    layer0_outputs(7500) <= not((inputs(109)) or (inputs(205)));
    layer0_outputs(7501) <= not(inputs(221));
    layer0_outputs(7502) <= not(inputs(247)) or (inputs(27));
    layer0_outputs(7503) <= (inputs(105)) or (inputs(49));
    layer0_outputs(7504) <= not((inputs(125)) xor (inputs(55)));
    layer0_outputs(7505) <= not(inputs(22));
    layer0_outputs(7506) <= not(inputs(194)) or (inputs(123));
    layer0_outputs(7507) <= (inputs(184)) or (inputs(240));
    layer0_outputs(7508) <= not(inputs(82));
    layer0_outputs(7509) <= (inputs(154)) xor (inputs(149));
    layer0_outputs(7510) <= (inputs(90)) xor (inputs(11));
    layer0_outputs(7511) <= not((inputs(77)) or (inputs(233)));
    layer0_outputs(7512) <= (inputs(55)) xor (inputs(55));
    layer0_outputs(7513) <= not((inputs(61)) xor (inputs(200)));
    layer0_outputs(7514) <= (inputs(82)) xor (inputs(118));
    layer0_outputs(7515) <= not((inputs(189)) xor (inputs(26)));
    layer0_outputs(7516) <= not(inputs(135)) or (inputs(61));
    layer0_outputs(7517) <= not(inputs(25)) or (inputs(237));
    layer0_outputs(7518) <= (inputs(104)) and (inputs(147));
    layer0_outputs(7519) <= not(inputs(14));
    layer0_outputs(7520) <= not(inputs(187));
    layer0_outputs(7521) <= not(inputs(182));
    layer0_outputs(7522) <= inputs(20);
    layer0_outputs(7523) <= not((inputs(223)) xor (inputs(35)));
    layer0_outputs(7524) <= (inputs(130)) and not (inputs(49));
    layer0_outputs(7525) <= '0';
    layer0_outputs(7526) <= (inputs(142)) and not (inputs(141));
    layer0_outputs(7527) <= not((inputs(97)) xor (inputs(136)));
    layer0_outputs(7528) <= not(inputs(209)) or (inputs(117));
    layer0_outputs(7529) <= (inputs(29)) xor (inputs(196));
    layer0_outputs(7530) <= (inputs(87)) or (inputs(211));
    layer0_outputs(7531) <= inputs(213);
    layer0_outputs(7532) <= inputs(96);
    layer0_outputs(7533) <= inputs(2);
    layer0_outputs(7534) <= not(inputs(58));
    layer0_outputs(7535) <= not(inputs(97)) or (inputs(38));
    layer0_outputs(7536) <= inputs(37);
    layer0_outputs(7537) <= not(inputs(9));
    layer0_outputs(7538) <= (inputs(60)) or (inputs(69));
    layer0_outputs(7539) <= not(inputs(64));
    layer0_outputs(7540) <= (inputs(21)) or (inputs(80));
    layer0_outputs(7541) <= not((inputs(207)) or (inputs(111)));
    layer0_outputs(7542) <= not((inputs(37)) xor (inputs(174)));
    layer0_outputs(7543) <= not(inputs(246));
    layer0_outputs(7544) <= (inputs(50)) and not (inputs(139));
    layer0_outputs(7545) <= (inputs(244)) xor (inputs(209));
    layer0_outputs(7546) <= not((inputs(121)) or (inputs(55)));
    layer0_outputs(7547) <= (inputs(36)) xor (inputs(21));
    layer0_outputs(7548) <= inputs(122);
    layer0_outputs(7549) <= not((inputs(5)) or (inputs(141)));
    layer0_outputs(7550) <= not(inputs(115));
    layer0_outputs(7551) <= not(inputs(86)) or (inputs(252));
    layer0_outputs(7552) <= (inputs(230)) or (inputs(243));
    layer0_outputs(7553) <= inputs(243);
    layer0_outputs(7554) <= not(inputs(218)) or (inputs(83));
    layer0_outputs(7555) <= inputs(6);
    layer0_outputs(7556) <= (inputs(24)) and not (inputs(203));
    layer0_outputs(7557) <= (inputs(221)) or (inputs(43));
    layer0_outputs(7558) <= (inputs(35)) or (inputs(25));
    layer0_outputs(7559) <= not((inputs(126)) or (inputs(218)));
    layer0_outputs(7560) <= not(inputs(148)) or (inputs(160));
    layer0_outputs(7561) <= (inputs(89)) and not (inputs(180));
    layer0_outputs(7562) <= not(inputs(233));
    layer0_outputs(7563) <= not((inputs(180)) or (inputs(191)));
    layer0_outputs(7564) <= not(inputs(152)) or (inputs(196));
    layer0_outputs(7565) <= (inputs(90)) xor (inputs(79));
    layer0_outputs(7566) <= not((inputs(209)) xor (inputs(215)));
    layer0_outputs(7567) <= not(inputs(195));
    layer0_outputs(7568) <= (inputs(13)) and not (inputs(78));
    layer0_outputs(7569) <= (inputs(50)) xor (inputs(88));
    layer0_outputs(7570) <= not((inputs(13)) xor (inputs(7)));
    layer0_outputs(7571) <= not(inputs(150));
    layer0_outputs(7572) <= not(inputs(150)) or (inputs(186));
    layer0_outputs(7573) <= (inputs(3)) or (inputs(114));
    layer0_outputs(7574) <= not(inputs(113));
    layer0_outputs(7575) <= inputs(246);
    layer0_outputs(7576) <= not(inputs(216));
    layer0_outputs(7577) <= not(inputs(85)) or (inputs(57));
    layer0_outputs(7578) <= (inputs(11)) or (inputs(237));
    layer0_outputs(7579) <= not(inputs(75));
    layer0_outputs(7580) <= not(inputs(176));
    layer0_outputs(7581) <= inputs(149);
    layer0_outputs(7582) <= (inputs(181)) and not (inputs(36));
    layer0_outputs(7583) <= not((inputs(174)) xor (inputs(225)));
    layer0_outputs(7584) <= not((inputs(128)) xor (inputs(95)));
    layer0_outputs(7585) <= inputs(141);
    layer0_outputs(7586) <= not((inputs(170)) xor (inputs(19)));
    layer0_outputs(7587) <= (inputs(246)) xor (inputs(105));
    layer0_outputs(7588) <= (inputs(87)) or (inputs(214));
    layer0_outputs(7589) <= inputs(110);
    layer0_outputs(7590) <= (inputs(96)) xor (inputs(245));
    layer0_outputs(7591) <= not((inputs(10)) xor (inputs(41)));
    layer0_outputs(7592) <= not(inputs(237));
    layer0_outputs(7593) <= inputs(9);
    layer0_outputs(7594) <= not((inputs(210)) xor (inputs(224)));
    layer0_outputs(7595) <= not((inputs(202)) or (inputs(86)));
    layer0_outputs(7596) <= (inputs(249)) and not (inputs(94));
    layer0_outputs(7597) <= not((inputs(115)) and (inputs(13)));
    layer0_outputs(7598) <= not(inputs(129));
    layer0_outputs(7599) <= not((inputs(79)) or (inputs(137)));
    layer0_outputs(7600) <= (inputs(174)) and not (inputs(153));
    layer0_outputs(7601) <= not((inputs(134)) and (inputs(231)));
    layer0_outputs(7602) <= inputs(5);
    layer0_outputs(7603) <= not(inputs(87));
    layer0_outputs(7604) <= not(inputs(40));
    layer0_outputs(7605) <= not((inputs(131)) or (inputs(160)));
    layer0_outputs(7606) <= not(inputs(89));
    layer0_outputs(7607) <= (inputs(147)) and not (inputs(4));
    layer0_outputs(7608) <= not((inputs(249)) or (inputs(20)));
    layer0_outputs(7609) <= not(inputs(142));
    layer0_outputs(7610) <= not(inputs(26)) or (inputs(161));
    layer0_outputs(7611) <= (inputs(24)) and not (inputs(128));
    layer0_outputs(7612) <= not(inputs(30));
    layer0_outputs(7613) <= inputs(146);
    layer0_outputs(7614) <= inputs(173);
    layer0_outputs(7615) <= (inputs(220)) and not (inputs(185));
    layer0_outputs(7616) <= not((inputs(190)) or (inputs(164)));
    layer0_outputs(7617) <= inputs(63);
    layer0_outputs(7618) <= inputs(249);
    layer0_outputs(7619) <= inputs(226);
    layer0_outputs(7620) <= not(inputs(214));
    layer0_outputs(7621) <= '1';
    layer0_outputs(7622) <= not(inputs(210));
    layer0_outputs(7623) <= not(inputs(173));
    layer0_outputs(7624) <= not((inputs(174)) and (inputs(27)));
    layer0_outputs(7625) <= not((inputs(39)) and (inputs(249)));
    layer0_outputs(7626) <= not((inputs(214)) xor (inputs(32)));
    layer0_outputs(7627) <= not(inputs(67)) or (inputs(111));
    layer0_outputs(7628) <= not((inputs(120)) and (inputs(75)));
    layer0_outputs(7629) <= inputs(123);
    layer0_outputs(7630) <= inputs(233);
    layer0_outputs(7631) <= not(inputs(232));
    layer0_outputs(7632) <= inputs(8);
    layer0_outputs(7633) <= (inputs(97)) and not (inputs(73));
    layer0_outputs(7634) <= not((inputs(78)) or (inputs(69)));
    layer0_outputs(7635) <= not((inputs(221)) or (inputs(6)));
    layer0_outputs(7636) <= not((inputs(25)) xor (inputs(117)));
    layer0_outputs(7637) <= (inputs(133)) and not (inputs(111));
    layer0_outputs(7638) <= inputs(158);
    layer0_outputs(7639) <= not((inputs(179)) or (inputs(218)));
    layer0_outputs(7640) <= inputs(252);
    layer0_outputs(7641) <= not((inputs(194)) xor (inputs(11)));
    layer0_outputs(7642) <= not((inputs(78)) or (inputs(43)));
    layer0_outputs(7643) <= not(inputs(3));
    layer0_outputs(7644) <= not(inputs(109));
    layer0_outputs(7645) <= (inputs(181)) and not (inputs(192));
    layer0_outputs(7646) <= not(inputs(186)) or (inputs(222));
    layer0_outputs(7647) <= not((inputs(85)) or (inputs(146)));
    layer0_outputs(7648) <= '0';
    layer0_outputs(7649) <= not(inputs(188)) or (inputs(29));
    layer0_outputs(7650) <= not((inputs(30)) or (inputs(249)));
    layer0_outputs(7651) <= (inputs(254)) xor (inputs(46));
    layer0_outputs(7652) <= (inputs(229)) or (inputs(178));
    layer0_outputs(7653) <= not(inputs(249)) or (inputs(154));
    layer0_outputs(7654) <= (inputs(74)) xor (inputs(24));
    layer0_outputs(7655) <= (inputs(218)) or (inputs(2));
    layer0_outputs(7656) <= inputs(168);
    layer0_outputs(7657) <= (inputs(59)) and not (inputs(7));
    layer0_outputs(7658) <= (inputs(51)) or (inputs(157));
    layer0_outputs(7659) <= (inputs(11)) and (inputs(134));
    layer0_outputs(7660) <= not(inputs(89));
    layer0_outputs(7661) <= not(inputs(179)) or (inputs(32));
    layer0_outputs(7662) <= not(inputs(203)) or (inputs(57));
    layer0_outputs(7663) <= not(inputs(81)) or (inputs(240));
    layer0_outputs(7664) <= inputs(76);
    layer0_outputs(7665) <= (inputs(172)) or (inputs(14));
    layer0_outputs(7666) <= not(inputs(25)) or (inputs(221));
    layer0_outputs(7667) <= (inputs(78)) and not (inputs(34));
    layer0_outputs(7668) <= (inputs(34)) and (inputs(33));
    layer0_outputs(7669) <= (inputs(105)) and not (inputs(157));
    layer0_outputs(7670) <= not((inputs(55)) and (inputs(238)));
    layer0_outputs(7671) <= (inputs(151)) and not (inputs(163));
    layer0_outputs(7672) <= (inputs(193)) or (inputs(206));
    layer0_outputs(7673) <= not((inputs(255)) xor (inputs(241)));
    layer0_outputs(7674) <= (inputs(100)) or (inputs(196));
    layer0_outputs(7675) <= not(inputs(42));
    layer0_outputs(7676) <= inputs(248);
    layer0_outputs(7677) <= inputs(66);
    layer0_outputs(7678) <= (inputs(202)) or (inputs(77));
    layer0_outputs(7679) <= not(inputs(169));
    layer0_outputs(7680) <= (inputs(64)) xor (inputs(63));
    layer0_outputs(7681) <= inputs(108);
    layer0_outputs(7682) <= inputs(210);
    layer0_outputs(7683) <= not((inputs(76)) xor (inputs(230)));
    layer0_outputs(7684) <= (inputs(119)) and not (inputs(65));
    layer0_outputs(7685) <= (inputs(171)) or (inputs(187));
    layer0_outputs(7686) <= not(inputs(32));
    layer0_outputs(7687) <= inputs(48);
    layer0_outputs(7688) <= not((inputs(111)) or (inputs(26)));
    layer0_outputs(7689) <= (inputs(212)) and not (inputs(106));
    layer0_outputs(7690) <= '0';
    layer0_outputs(7691) <= not((inputs(149)) xor (inputs(42)));
    layer0_outputs(7692) <= not((inputs(97)) or (inputs(149)));
    layer0_outputs(7693) <= not((inputs(98)) and (inputs(112)));
    layer0_outputs(7694) <= inputs(253);
    layer0_outputs(7695) <= (inputs(228)) xor (inputs(150));
    layer0_outputs(7696) <= not((inputs(196)) and (inputs(253)));
    layer0_outputs(7697) <= (inputs(104)) and not (inputs(49));
    layer0_outputs(7698) <= not(inputs(68));
    layer0_outputs(7699) <= inputs(3);
    layer0_outputs(7700) <= (inputs(127)) xor (inputs(186));
    layer0_outputs(7701) <= (inputs(33)) and not (inputs(83));
    layer0_outputs(7702) <= not(inputs(110));
    layer0_outputs(7703) <= '0';
    layer0_outputs(7704) <= (inputs(150)) xor (inputs(55));
    layer0_outputs(7705) <= inputs(248);
    layer0_outputs(7706) <= inputs(73);
    layer0_outputs(7707) <= not((inputs(47)) or (inputs(53)));
    layer0_outputs(7708) <= (inputs(46)) xor (inputs(0));
    layer0_outputs(7709) <= not(inputs(225));
    layer0_outputs(7710) <= (inputs(91)) xor (inputs(43));
    layer0_outputs(7711) <= inputs(153);
    layer0_outputs(7712) <= inputs(128);
    layer0_outputs(7713) <= not((inputs(41)) xor (inputs(160)));
    layer0_outputs(7714) <= inputs(114);
    layer0_outputs(7715) <= not(inputs(233)) or (inputs(109));
    layer0_outputs(7716) <= not((inputs(141)) or (inputs(99)));
    layer0_outputs(7717) <= not((inputs(60)) xor (inputs(30)));
    layer0_outputs(7718) <= (inputs(126)) xor (inputs(68));
    layer0_outputs(7719) <= (inputs(137)) and not (inputs(87));
    layer0_outputs(7720) <= not((inputs(76)) or (inputs(124)));
    layer0_outputs(7721) <= not((inputs(95)) xor (inputs(233)));
    layer0_outputs(7722) <= (inputs(252)) and not (inputs(190));
    layer0_outputs(7723) <= (inputs(42)) or (inputs(241));
    layer0_outputs(7724) <= inputs(175);
    layer0_outputs(7725) <= not(inputs(235)) or (inputs(47));
    layer0_outputs(7726) <= (inputs(206)) or (inputs(54));
    layer0_outputs(7727) <= (inputs(196)) or (inputs(190));
    layer0_outputs(7728) <= (inputs(194)) or (inputs(49));
    layer0_outputs(7729) <= not((inputs(244)) xor (inputs(242)));
    layer0_outputs(7730) <= not((inputs(104)) xor (inputs(52)));
    layer0_outputs(7731) <= (inputs(153)) and not (inputs(28));
    layer0_outputs(7732) <= inputs(11);
    layer0_outputs(7733) <= not(inputs(18)) or (inputs(236));
    layer0_outputs(7734) <= (inputs(41)) xor (inputs(25));
    layer0_outputs(7735) <= not(inputs(26));
    layer0_outputs(7736) <= (inputs(137)) xor (inputs(138));
    layer0_outputs(7737) <= inputs(107);
    layer0_outputs(7738) <= (inputs(192)) or (inputs(4));
    layer0_outputs(7739) <= (inputs(40)) and not (inputs(125));
    layer0_outputs(7740) <= (inputs(46)) or (inputs(21));
    layer0_outputs(7741) <= not((inputs(6)) xor (inputs(24)));
    layer0_outputs(7742) <= not(inputs(61)) or (inputs(255));
    layer0_outputs(7743) <= (inputs(235)) xor (inputs(162));
    layer0_outputs(7744) <= inputs(65);
    layer0_outputs(7745) <= not((inputs(190)) xor (inputs(9)));
    layer0_outputs(7746) <= (inputs(204)) xor (inputs(156));
    layer0_outputs(7747) <= inputs(102);
    layer0_outputs(7748) <= not(inputs(36));
    layer0_outputs(7749) <= (inputs(75)) and not (inputs(28));
    layer0_outputs(7750) <= inputs(26);
    layer0_outputs(7751) <= not((inputs(8)) or (inputs(134)));
    layer0_outputs(7752) <= not(inputs(114));
    layer0_outputs(7753) <= '0';
    layer0_outputs(7754) <= (inputs(83)) and not (inputs(175));
    layer0_outputs(7755) <= inputs(18);
    layer0_outputs(7756) <= (inputs(59)) or (inputs(93));
    layer0_outputs(7757) <= (inputs(121)) and not (inputs(190));
    layer0_outputs(7758) <= not((inputs(23)) xor (inputs(168)));
    layer0_outputs(7759) <= not(inputs(121));
    layer0_outputs(7760) <= not((inputs(75)) or (inputs(65)));
    layer0_outputs(7761) <= not(inputs(134));
    layer0_outputs(7762) <= not(inputs(77)) or (inputs(89));
    layer0_outputs(7763) <= not((inputs(22)) or (inputs(123)));
    layer0_outputs(7764) <= not(inputs(133));
    layer0_outputs(7765) <= not(inputs(241));
    layer0_outputs(7766) <= (inputs(59)) and not (inputs(37));
    layer0_outputs(7767) <= (inputs(138)) or (inputs(246));
    layer0_outputs(7768) <= not(inputs(233)) or (inputs(5));
    layer0_outputs(7769) <= not((inputs(175)) xor (inputs(195)));
    layer0_outputs(7770) <= not((inputs(247)) xor (inputs(199)));
    layer0_outputs(7771) <= not((inputs(214)) or (inputs(189)));
    layer0_outputs(7772) <= (inputs(180)) xor (inputs(224));
    layer0_outputs(7773) <= not((inputs(154)) and (inputs(18)));
    layer0_outputs(7774) <= not(inputs(150));
    layer0_outputs(7775) <= (inputs(36)) xor (inputs(71));
    layer0_outputs(7776) <= inputs(105);
    layer0_outputs(7777) <= not((inputs(116)) or (inputs(63)));
    layer0_outputs(7778) <= not(inputs(167));
    layer0_outputs(7779) <= (inputs(181)) xor (inputs(120));
    layer0_outputs(7780) <= (inputs(188)) and not (inputs(102));
    layer0_outputs(7781) <= not(inputs(166)) or (inputs(102));
    layer0_outputs(7782) <= not((inputs(225)) and (inputs(138)));
    layer0_outputs(7783) <= inputs(92);
    layer0_outputs(7784) <= not(inputs(183)) or (inputs(188));
    layer0_outputs(7785) <= not((inputs(234)) xor (inputs(185)));
    layer0_outputs(7786) <= not(inputs(120)) or (inputs(158));
    layer0_outputs(7787) <= (inputs(192)) xor (inputs(4));
    layer0_outputs(7788) <= not((inputs(36)) or (inputs(215)));
    layer0_outputs(7789) <= '1';
    layer0_outputs(7790) <= inputs(10);
    layer0_outputs(7791) <= '1';
    layer0_outputs(7792) <= not(inputs(167));
    layer0_outputs(7793) <= (inputs(170)) or (inputs(218));
    layer0_outputs(7794) <= not(inputs(200));
    layer0_outputs(7795) <= (inputs(79)) or (inputs(85));
    layer0_outputs(7796) <= (inputs(138)) and (inputs(170));
    layer0_outputs(7797) <= inputs(196);
    layer0_outputs(7798) <= not(inputs(79));
    layer0_outputs(7799) <= not((inputs(148)) or (inputs(201)));
    layer0_outputs(7800) <= not((inputs(254)) or (inputs(17)));
    layer0_outputs(7801) <= (inputs(140)) and not (inputs(22));
    layer0_outputs(7802) <= not((inputs(201)) xor (inputs(231)));
    layer0_outputs(7803) <= inputs(189);
    layer0_outputs(7804) <= not(inputs(61));
    layer0_outputs(7805) <= not(inputs(1)) or (inputs(51));
    layer0_outputs(7806) <= not(inputs(24));
    layer0_outputs(7807) <= not(inputs(118));
    layer0_outputs(7808) <= (inputs(87)) or (inputs(34));
    layer0_outputs(7809) <= not((inputs(206)) xor (inputs(70)));
    layer0_outputs(7810) <= not(inputs(89)) or (inputs(155));
    layer0_outputs(7811) <= not(inputs(11));
    layer0_outputs(7812) <= (inputs(242)) and not (inputs(39));
    layer0_outputs(7813) <= not(inputs(122));
    layer0_outputs(7814) <= not(inputs(114)) or (inputs(250));
    layer0_outputs(7815) <= (inputs(149)) or (inputs(253));
    layer0_outputs(7816) <= (inputs(72)) or (inputs(129));
    layer0_outputs(7817) <= not(inputs(231));
    layer0_outputs(7818) <= not(inputs(87)) or (inputs(181));
    layer0_outputs(7819) <= not((inputs(72)) or (inputs(38)));
    layer0_outputs(7820) <= not((inputs(94)) or (inputs(61)));
    layer0_outputs(7821) <= not((inputs(102)) or (inputs(85)));
    layer0_outputs(7822) <= inputs(18);
    layer0_outputs(7823) <= (inputs(174)) or (inputs(55));
    layer0_outputs(7824) <= not(inputs(153)) or (inputs(71));
    layer0_outputs(7825) <= not(inputs(167));
    layer0_outputs(7826) <= (inputs(215)) and not (inputs(97));
    layer0_outputs(7827) <= inputs(241);
    layer0_outputs(7828) <= inputs(74);
    layer0_outputs(7829) <= not(inputs(220)) or (inputs(91));
    layer0_outputs(7830) <= not(inputs(19));
    layer0_outputs(7831) <= (inputs(25)) xor (inputs(56));
    layer0_outputs(7832) <= (inputs(68)) or (inputs(114));
    layer0_outputs(7833) <= not(inputs(135));
    layer0_outputs(7834) <= (inputs(110)) and not (inputs(176));
    layer0_outputs(7835) <= not(inputs(68));
    layer0_outputs(7836) <= (inputs(176)) or (inputs(63));
    layer0_outputs(7837) <= inputs(218);
    layer0_outputs(7838) <= not(inputs(182));
    layer0_outputs(7839) <= inputs(164);
    layer0_outputs(7840) <= not((inputs(55)) or (inputs(254)));
    layer0_outputs(7841) <= (inputs(203)) or (inputs(16));
    layer0_outputs(7842) <= (inputs(146)) or (inputs(175));
    layer0_outputs(7843) <= (inputs(230)) or (inputs(2));
    layer0_outputs(7844) <= not((inputs(77)) or (inputs(143)));
    layer0_outputs(7845) <= (inputs(58)) and not (inputs(101));
    layer0_outputs(7846) <= not((inputs(230)) or (inputs(110)));
    layer0_outputs(7847) <= '0';
    layer0_outputs(7848) <= (inputs(66)) or (inputs(185));
    layer0_outputs(7849) <= inputs(34);
    layer0_outputs(7850) <= inputs(22);
    layer0_outputs(7851) <= (inputs(114)) or (inputs(98));
    layer0_outputs(7852) <= (inputs(235)) or (inputs(23));
    layer0_outputs(7853) <= '1';
    layer0_outputs(7854) <= (inputs(226)) or (inputs(236));
    layer0_outputs(7855) <= (inputs(248)) or (inputs(156));
    layer0_outputs(7856) <= inputs(65);
    layer0_outputs(7857) <= (inputs(168)) or (inputs(239));
    layer0_outputs(7858) <= '0';
    layer0_outputs(7859) <= (inputs(31)) xor (inputs(6));
    layer0_outputs(7860) <= not((inputs(70)) or (inputs(194)));
    layer0_outputs(7861) <= (inputs(188)) and not (inputs(36));
    layer0_outputs(7862) <= (inputs(25)) xor (inputs(195));
    layer0_outputs(7863) <= not((inputs(244)) or (inputs(250)));
    layer0_outputs(7864) <= not((inputs(154)) and (inputs(32)));
    layer0_outputs(7865) <= not(inputs(228));
    layer0_outputs(7866) <= not(inputs(167)) or (inputs(71));
    layer0_outputs(7867) <= not((inputs(112)) xor (inputs(100)));
    layer0_outputs(7868) <= not(inputs(162));
    layer0_outputs(7869) <= inputs(139);
    layer0_outputs(7870) <= (inputs(57)) xor (inputs(103));
    layer0_outputs(7871) <= (inputs(7)) or (inputs(230));
    layer0_outputs(7872) <= not(inputs(227));
    layer0_outputs(7873) <= not((inputs(65)) or (inputs(111)));
    layer0_outputs(7874) <= not(inputs(148)) or (inputs(7));
    layer0_outputs(7875) <= inputs(245);
    layer0_outputs(7876) <= not((inputs(58)) xor (inputs(44)));
    layer0_outputs(7877) <= not(inputs(167)) or (inputs(47));
    layer0_outputs(7878) <= not(inputs(160));
    layer0_outputs(7879) <= (inputs(165)) and not (inputs(213));
    layer0_outputs(7880) <= not((inputs(151)) or (inputs(219)));
    layer0_outputs(7881) <= (inputs(97)) or (inputs(173));
    layer0_outputs(7882) <= (inputs(203)) xor (inputs(98));
    layer0_outputs(7883) <= not(inputs(57));
    layer0_outputs(7884) <= not(inputs(158));
    layer0_outputs(7885) <= not((inputs(94)) or (inputs(117)));
    layer0_outputs(7886) <= not((inputs(48)) xor (inputs(134)));
    layer0_outputs(7887) <= '1';
    layer0_outputs(7888) <= not((inputs(146)) xor (inputs(112)));
    layer0_outputs(7889) <= '0';
    layer0_outputs(7890) <= (inputs(160)) or (inputs(228));
    layer0_outputs(7891) <= (inputs(4)) and (inputs(103));
    layer0_outputs(7892) <= (inputs(196)) and (inputs(91));
    layer0_outputs(7893) <= not(inputs(220));
    layer0_outputs(7894) <= not(inputs(247)) or (inputs(81));
    layer0_outputs(7895) <= not((inputs(115)) xor (inputs(178)));
    layer0_outputs(7896) <= inputs(163);
    layer0_outputs(7897) <= not((inputs(142)) xor (inputs(109)));
    layer0_outputs(7898) <= not((inputs(81)) or (inputs(254)));
    layer0_outputs(7899) <= (inputs(238)) or (inputs(163));
    layer0_outputs(7900) <= not(inputs(196)) or (inputs(107));
    layer0_outputs(7901) <= inputs(162);
    layer0_outputs(7902) <= not(inputs(73)) or (inputs(135));
    layer0_outputs(7903) <= (inputs(202)) or (inputs(195));
    layer0_outputs(7904) <= not((inputs(205)) or (inputs(176)));
    layer0_outputs(7905) <= not(inputs(93));
    layer0_outputs(7906) <= inputs(40);
    layer0_outputs(7907) <= inputs(214);
    layer0_outputs(7908) <= not(inputs(53));
    layer0_outputs(7909) <= (inputs(112)) or (inputs(67));
    layer0_outputs(7910) <= not(inputs(58)) or (inputs(86));
    layer0_outputs(7911) <= '1';
    layer0_outputs(7912) <= not((inputs(112)) or (inputs(237)));
    layer0_outputs(7913) <= (inputs(157)) or (inputs(189));
    layer0_outputs(7914) <= inputs(62);
    layer0_outputs(7915) <= not(inputs(155)) or (inputs(224));
    layer0_outputs(7916) <= (inputs(17)) or (inputs(103));
    layer0_outputs(7917) <= not((inputs(138)) or (inputs(46)));
    layer0_outputs(7918) <= not((inputs(60)) xor (inputs(95)));
    layer0_outputs(7919) <= (inputs(244)) and not (inputs(210));
    layer0_outputs(7920) <= (inputs(104)) xor (inputs(245));
    layer0_outputs(7921) <= (inputs(163)) and not (inputs(63));
    layer0_outputs(7922) <= inputs(59);
    layer0_outputs(7923) <= (inputs(23)) and not (inputs(14));
    layer0_outputs(7924) <= inputs(69);
    layer0_outputs(7925) <= not(inputs(209));
    layer0_outputs(7926) <= not(inputs(2)) or (inputs(224));
    layer0_outputs(7927) <= not((inputs(38)) xor (inputs(111)));
    layer0_outputs(7928) <= inputs(202);
    layer0_outputs(7929) <= (inputs(175)) and not (inputs(47));
    layer0_outputs(7930) <= (inputs(83)) xor (inputs(209));
    layer0_outputs(7931) <= inputs(128);
    layer0_outputs(7932) <= inputs(113);
    layer0_outputs(7933) <= not(inputs(141)) or (inputs(253));
    layer0_outputs(7934) <= (inputs(198)) xor (inputs(202));
    layer0_outputs(7935) <= inputs(166);
    layer0_outputs(7936) <= not((inputs(243)) or (inputs(240)));
    layer0_outputs(7937) <= inputs(167);
    layer0_outputs(7938) <= not(inputs(198)) or (inputs(194));
    layer0_outputs(7939) <= inputs(41);
    layer0_outputs(7940) <= inputs(182);
    layer0_outputs(7941) <= not((inputs(106)) xor (inputs(44)));
    layer0_outputs(7942) <= (inputs(140)) or (inputs(143));
    layer0_outputs(7943) <= not((inputs(20)) or (inputs(0)));
    layer0_outputs(7944) <= not((inputs(57)) or (inputs(3)));
    layer0_outputs(7945) <= inputs(87);
    layer0_outputs(7946) <= (inputs(63)) and not (inputs(183));
    layer0_outputs(7947) <= (inputs(119)) and not (inputs(214));
    layer0_outputs(7948) <= not((inputs(23)) xor (inputs(146)));
    layer0_outputs(7949) <= (inputs(59)) and not (inputs(80));
    layer0_outputs(7950) <= (inputs(100)) or (inputs(187));
    layer0_outputs(7951) <= not((inputs(39)) or (inputs(175)));
    layer0_outputs(7952) <= (inputs(205)) xor (inputs(48));
    layer0_outputs(7953) <= not((inputs(143)) or (inputs(89)));
    layer0_outputs(7954) <= not(inputs(9)) or (inputs(129));
    layer0_outputs(7955) <= (inputs(2)) xor (inputs(201));
    layer0_outputs(7956) <= (inputs(135)) xor (inputs(163));
    layer0_outputs(7957) <= inputs(212);
    layer0_outputs(7958) <= (inputs(112)) and not (inputs(3));
    layer0_outputs(7959) <= not(inputs(201)) or (inputs(89));
    layer0_outputs(7960) <= not(inputs(8));
    layer0_outputs(7961) <= not(inputs(116));
    layer0_outputs(7962) <= inputs(233);
    layer0_outputs(7963) <= not((inputs(182)) xor (inputs(177)));
    layer0_outputs(7964) <= not(inputs(145));
    layer0_outputs(7965) <= (inputs(159)) and not (inputs(28));
    layer0_outputs(7966) <= not(inputs(135)) or (inputs(16));
    layer0_outputs(7967) <= inputs(168);
    layer0_outputs(7968) <= not((inputs(70)) xor (inputs(129)));
    layer0_outputs(7969) <= inputs(126);
    layer0_outputs(7970) <= not((inputs(87)) xor (inputs(114)));
    layer0_outputs(7971) <= not((inputs(183)) or (inputs(45)));
    layer0_outputs(7972) <= (inputs(153)) xor (inputs(239));
    layer0_outputs(7973) <= not((inputs(237)) xor (inputs(129)));
    layer0_outputs(7974) <= (inputs(37)) and not (inputs(106));
    layer0_outputs(7975) <= not((inputs(226)) and (inputs(227)));
    layer0_outputs(7976) <= not(inputs(113));
    layer0_outputs(7977) <= inputs(172);
    layer0_outputs(7978) <= (inputs(192)) or (inputs(172));
    layer0_outputs(7979) <= (inputs(16)) or (inputs(204));
    layer0_outputs(7980) <= (inputs(28)) and not (inputs(128));
    layer0_outputs(7981) <= (inputs(215)) xor (inputs(194));
    layer0_outputs(7982) <= not((inputs(7)) or (inputs(190)));
    layer0_outputs(7983) <= not((inputs(78)) or (inputs(99)));
    layer0_outputs(7984) <= not((inputs(196)) or (inputs(221)));
    layer0_outputs(7985) <= not(inputs(212)) or (inputs(3));
    layer0_outputs(7986) <= (inputs(41)) and (inputs(6));
    layer0_outputs(7987) <= (inputs(7)) or (inputs(97));
    layer0_outputs(7988) <= (inputs(52)) and not (inputs(250));
    layer0_outputs(7989) <= (inputs(102)) or (inputs(85));
    layer0_outputs(7990) <= not((inputs(240)) or (inputs(45)));
    layer0_outputs(7991) <= not(inputs(183)) or (inputs(128));
    layer0_outputs(7992) <= not(inputs(67));
    layer0_outputs(7993) <= not(inputs(44)) or (inputs(191));
    layer0_outputs(7994) <= not((inputs(253)) xor (inputs(64)));
    layer0_outputs(7995) <= (inputs(29)) and not (inputs(47));
    layer0_outputs(7996) <= not(inputs(122));
    layer0_outputs(7997) <= (inputs(206)) and not (inputs(65));
    layer0_outputs(7998) <= (inputs(223)) and not (inputs(96));
    layer0_outputs(7999) <= not((inputs(56)) or (inputs(217)));
    layer0_outputs(8000) <= not(inputs(94));
    layer0_outputs(8001) <= inputs(148);
    layer0_outputs(8002) <= (inputs(18)) or (inputs(195));
    layer0_outputs(8003) <= not(inputs(212));
    layer0_outputs(8004) <= (inputs(14)) or (inputs(129));
    layer0_outputs(8005) <= inputs(200);
    layer0_outputs(8006) <= not(inputs(7));
    layer0_outputs(8007) <= inputs(181);
    layer0_outputs(8008) <= not(inputs(168));
    layer0_outputs(8009) <= inputs(119);
    layer0_outputs(8010) <= (inputs(79)) or (inputs(249));
    layer0_outputs(8011) <= not(inputs(177));
    layer0_outputs(8012) <= inputs(76);
    layer0_outputs(8013) <= inputs(118);
    layer0_outputs(8014) <= not((inputs(140)) and (inputs(247)));
    layer0_outputs(8015) <= not(inputs(230));
    layer0_outputs(8016) <= not((inputs(180)) xor (inputs(144)));
    layer0_outputs(8017) <= not(inputs(61)) or (inputs(64));
    layer0_outputs(8018) <= not(inputs(78));
    layer0_outputs(8019) <= inputs(178);
    layer0_outputs(8020) <= (inputs(213)) xor (inputs(177));
    layer0_outputs(8021) <= not(inputs(78));
    layer0_outputs(8022) <= not((inputs(226)) xor (inputs(180)));
    layer0_outputs(8023) <= not((inputs(0)) or (inputs(133)));
    layer0_outputs(8024) <= not(inputs(216));
    layer0_outputs(8025) <= not((inputs(165)) or (inputs(166)));
    layer0_outputs(8026) <= (inputs(2)) xor (inputs(106));
    layer0_outputs(8027) <= not((inputs(115)) or (inputs(109)));
    layer0_outputs(8028) <= not((inputs(71)) and (inputs(88)));
    layer0_outputs(8029) <= (inputs(74)) and not (inputs(30));
    layer0_outputs(8030) <= (inputs(81)) or (inputs(212));
    layer0_outputs(8031) <= not((inputs(25)) and (inputs(183)));
    layer0_outputs(8032) <= not(inputs(24));
    layer0_outputs(8033) <= not(inputs(161));
    layer0_outputs(8034) <= (inputs(243)) or (inputs(87));
    layer0_outputs(8035) <= not((inputs(60)) and (inputs(186)));
    layer0_outputs(8036) <= not(inputs(162));
    layer0_outputs(8037) <= not(inputs(82));
    layer0_outputs(8038) <= (inputs(102)) xor (inputs(164));
    layer0_outputs(8039) <= not(inputs(103)) or (inputs(221));
    layer0_outputs(8040) <= (inputs(6)) xor (inputs(152));
    layer0_outputs(8041) <= inputs(51);
    layer0_outputs(8042) <= (inputs(160)) xor (inputs(129));
    layer0_outputs(8043) <= not(inputs(155));
    layer0_outputs(8044) <= not((inputs(174)) and (inputs(145)));
    layer0_outputs(8045) <= not((inputs(29)) xor (inputs(32)));
    layer0_outputs(8046) <= (inputs(236)) or (inputs(144));
    layer0_outputs(8047) <= not(inputs(174));
    layer0_outputs(8048) <= not((inputs(167)) or (inputs(193)));
    layer0_outputs(8049) <= not((inputs(153)) or (inputs(254)));
    layer0_outputs(8050) <= not(inputs(25)) or (inputs(154));
    layer0_outputs(8051) <= not(inputs(46));
    layer0_outputs(8052) <= (inputs(139)) xor (inputs(19));
    layer0_outputs(8053) <= inputs(139);
    layer0_outputs(8054) <= (inputs(0)) or (inputs(110));
    layer0_outputs(8055) <= not(inputs(100));
    layer0_outputs(8056) <= inputs(74);
    layer0_outputs(8057) <= (inputs(36)) xor (inputs(6));
    layer0_outputs(8058) <= not(inputs(221));
    layer0_outputs(8059) <= (inputs(19)) and not (inputs(183));
    layer0_outputs(8060) <= not(inputs(250));
    layer0_outputs(8061) <= not((inputs(68)) or (inputs(8)));
    layer0_outputs(8062) <= (inputs(106)) xor (inputs(187));
    layer0_outputs(8063) <= not((inputs(164)) or (inputs(222)));
    layer0_outputs(8064) <= '0';
    layer0_outputs(8065) <= (inputs(49)) and not (inputs(191));
    layer0_outputs(8066) <= inputs(55);
    layer0_outputs(8067) <= not((inputs(229)) and (inputs(167)));
    layer0_outputs(8068) <= (inputs(136)) or (inputs(64));
    layer0_outputs(8069) <= not(inputs(132));
    layer0_outputs(8070) <= not((inputs(251)) xor (inputs(69)));
    layer0_outputs(8071) <= (inputs(153)) or (inputs(110));
    layer0_outputs(8072) <= inputs(68);
    layer0_outputs(8073) <= (inputs(52)) or (inputs(181));
    layer0_outputs(8074) <= inputs(113);
    layer0_outputs(8075) <= inputs(30);
    layer0_outputs(8076) <= not((inputs(146)) or (inputs(155)));
    layer0_outputs(8077) <= not((inputs(173)) or (inputs(194)));
    layer0_outputs(8078) <= not(inputs(137));
    layer0_outputs(8079) <= (inputs(49)) xor (inputs(77));
    layer0_outputs(8080) <= not((inputs(26)) xor (inputs(227)));
    layer0_outputs(8081) <= not((inputs(27)) and (inputs(229)));
    layer0_outputs(8082) <= inputs(218);
    layer0_outputs(8083) <= not(inputs(224));
    layer0_outputs(8084) <= (inputs(131)) and not (inputs(4));
    layer0_outputs(8085) <= (inputs(95)) or (inputs(81));
    layer0_outputs(8086) <= '0';
    layer0_outputs(8087) <= (inputs(108)) or (inputs(250));
    layer0_outputs(8088) <= (inputs(172)) and (inputs(19));
    layer0_outputs(8089) <= '0';
    layer0_outputs(8090) <= inputs(142);
    layer0_outputs(8091) <= not((inputs(226)) xor (inputs(65)));
    layer0_outputs(8092) <= not((inputs(56)) xor (inputs(73)));
    layer0_outputs(8093) <= not((inputs(183)) or (inputs(8)));
    layer0_outputs(8094) <= inputs(38);
    layer0_outputs(8095) <= (inputs(174)) or (inputs(29));
    layer0_outputs(8096) <= inputs(38);
    layer0_outputs(8097) <= not(inputs(233)) or (inputs(3));
    layer0_outputs(8098) <= inputs(50);
    layer0_outputs(8099) <= (inputs(218)) xor (inputs(101));
    layer0_outputs(8100) <= not(inputs(44)) or (inputs(129));
    layer0_outputs(8101) <= not((inputs(99)) xor (inputs(29)));
    layer0_outputs(8102) <= inputs(159);
    layer0_outputs(8103) <= not((inputs(200)) or (inputs(206)));
    layer0_outputs(8104) <= (inputs(244)) and not (inputs(221));
    layer0_outputs(8105) <= (inputs(221)) xor (inputs(19));
    layer0_outputs(8106) <= not(inputs(231)) or (inputs(79));
    layer0_outputs(8107) <= not(inputs(115));
    layer0_outputs(8108) <= not((inputs(4)) or (inputs(18)));
    layer0_outputs(8109) <= (inputs(204)) xor (inputs(240));
    layer0_outputs(8110) <= not(inputs(127)) or (inputs(34));
    layer0_outputs(8111) <= inputs(179);
    layer0_outputs(8112) <= inputs(229);
    layer0_outputs(8113) <= (inputs(17)) and not (inputs(252));
    layer0_outputs(8114) <= (inputs(175)) or (inputs(211));
    layer0_outputs(8115) <= not(inputs(135));
    layer0_outputs(8116) <= not((inputs(25)) or (inputs(100)));
    layer0_outputs(8117) <= (inputs(100)) xor (inputs(19));
    layer0_outputs(8118) <= (inputs(76)) and (inputs(232));
    layer0_outputs(8119) <= (inputs(175)) or (inputs(222));
    layer0_outputs(8120) <= inputs(224);
    layer0_outputs(8121) <= not(inputs(50));
    layer0_outputs(8122) <= not((inputs(75)) or (inputs(152)));
    layer0_outputs(8123) <= inputs(187);
    layer0_outputs(8124) <= (inputs(232)) or (inputs(23));
    layer0_outputs(8125) <= (inputs(33)) xor (inputs(63));
    layer0_outputs(8126) <= (inputs(131)) or (inputs(204));
    layer0_outputs(8127) <= (inputs(214)) or (inputs(132));
    layer0_outputs(8128) <= (inputs(25)) and not (inputs(220));
    layer0_outputs(8129) <= inputs(110);
    layer0_outputs(8130) <= not((inputs(79)) or (inputs(61)));
    layer0_outputs(8131) <= inputs(38);
    layer0_outputs(8132) <= (inputs(155)) or (inputs(130));
    layer0_outputs(8133) <= inputs(114);
    layer0_outputs(8134) <= inputs(153);
    layer0_outputs(8135) <= inputs(222);
    layer0_outputs(8136) <= not((inputs(50)) or (inputs(147)));
    layer0_outputs(8137) <= not((inputs(53)) and (inputs(29)));
    layer0_outputs(8138) <= not(inputs(131));
    layer0_outputs(8139) <= (inputs(173)) or (inputs(217));
    layer0_outputs(8140) <= not((inputs(46)) xor (inputs(68)));
    layer0_outputs(8141) <= not(inputs(114)) or (inputs(216));
    layer0_outputs(8142) <= not(inputs(208)) or (inputs(169));
    layer0_outputs(8143) <= not(inputs(184)) or (inputs(95));
    layer0_outputs(8144) <= (inputs(182)) or (inputs(69));
    layer0_outputs(8145) <= (inputs(24)) xor (inputs(5));
    layer0_outputs(8146) <= not((inputs(103)) xor (inputs(41)));
    layer0_outputs(8147) <= inputs(231);
    layer0_outputs(8148) <= not((inputs(119)) or (inputs(93)));
    layer0_outputs(8149) <= (inputs(243)) and not (inputs(37));
    layer0_outputs(8150) <= not(inputs(87));
    layer0_outputs(8151) <= (inputs(251)) or (inputs(10));
    layer0_outputs(8152) <= not(inputs(105)) or (inputs(214));
    layer0_outputs(8153) <= (inputs(249)) or (inputs(105));
    layer0_outputs(8154) <= not((inputs(172)) xor (inputs(173)));
    layer0_outputs(8155) <= (inputs(24)) and not (inputs(154));
    layer0_outputs(8156) <= not(inputs(126));
    layer0_outputs(8157) <= inputs(75);
    layer0_outputs(8158) <= (inputs(144)) and not (inputs(16));
    layer0_outputs(8159) <= inputs(197);
    layer0_outputs(8160) <= (inputs(97)) and not (inputs(11));
    layer0_outputs(8161) <= not(inputs(224)) or (inputs(183));
    layer0_outputs(8162) <= (inputs(65)) xor (inputs(32));
    layer0_outputs(8163) <= '0';
    layer0_outputs(8164) <= not((inputs(58)) and (inputs(4)));
    layer0_outputs(8165) <= not((inputs(127)) xor (inputs(99)));
    layer0_outputs(8166) <= (inputs(239)) or (inputs(221));
    layer0_outputs(8167) <= not((inputs(68)) or (inputs(52)));
    layer0_outputs(8168) <= not((inputs(50)) or (inputs(166)));
    layer0_outputs(8169) <= (inputs(206)) or (inputs(142));
    layer0_outputs(8170) <= not((inputs(112)) or (inputs(131)));
    layer0_outputs(8171) <= (inputs(193)) xor (inputs(143));
    layer0_outputs(8172) <= not(inputs(193));
    layer0_outputs(8173) <= (inputs(39)) and not (inputs(171));
    layer0_outputs(8174) <= not((inputs(129)) xor (inputs(166)));
    layer0_outputs(8175) <= (inputs(35)) xor (inputs(61));
    layer0_outputs(8176) <= (inputs(85)) xor (inputs(124));
    layer0_outputs(8177) <= not((inputs(30)) xor (inputs(61)));
    layer0_outputs(8178) <= not((inputs(8)) or (inputs(97)));
    layer0_outputs(8179) <= inputs(91);
    layer0_outputs(8180) <= not(inputs(121));
    layer0_outputs(8181) <= not(inputs(110));
    layer0_outputs(8182) <= (inputs(88)) xor (inputs(13));
    layer0_outputs(8183) <= (inputs(41)) and (inputs(120));
    layer0_outputs(8184) <= not((inputs(155)) xor (inputs(47)));
    layer0_outputs(8185) <= '0';
    layer0_outputs(8186) <= (inputs(44)) or (inputs(15));
    layer0_outputs(8187) <= not((inputs(159)) and (inputs(191)));
    layer0_outputs(8188) <= not((inputs(202)) or (inputs(79)));
    layer0_outputs(8189) <= inputs(255);
    layer0_outputs(8190) <= not((inputs(253)) or (inputs(66)));
    layer0_outputs(8191) <= (inputs(252)) or (inputs(131));
    layer0_outputs(8192) <= not(inputs(212));
    layer0_outputs(8193) <= not((inputs(183)) or (inputs(221)));
    layer0_outputs(8194) <= not((inputs(96)) xor (inputs(182)));
    layer0_outputs(8195) <= inputs(71);
    layer0_outputs(8196) <= not((inputs(167)) xor (inputs(145)));
    layer0_outputs(8197) <= not(inputs(189)) or (inputs(225));
    layer0_outputs(8198) <= not((inputs(99)) or (inputs(155)));
    layer0_outputs(8199) <= not((inputs(150)) or (inputs(182)));
    layer0_outputs(8200) <= not(inputs(94));
    layer0_outputs(8201) <= (inputs(165)) or (inputs(149));
    layer0_outputs(8202) <= not(inputs(236)) or (inputs(85));
    layer0_outputs(8203) <= '0';
    layer0_outputs(8204) <= not((inputs(209)) and (inputs(126)));
    layer0_outputs(8205) <= not((inputs(252)) xor (inputs(221)));
    layer0_outputs(8206) <= not((inputs(246)) or (inputs(142)));
    layer0_outputs(8207) <= not(inputs(38));
    layer0_outputs(8208) <= inputs(23);
    layer0_outputs(8209) <= (inputs(192)) or (inputs(58));
    layer0_outputs(8210) <= (inputs(182)) and not (inputs(85));
    layer0_outputs(8211) <= not(inputs(245)) or (inputs(116));
    layer0_outputs(8212) <= not(inputs(163));
    layer0_outputs(8213) <= inputs(125);
    layer0_outputs(8214) <= (inputs(154)) or (inputs(163));
    layer0_outputs(8215) <= not(inputs(124));
    layer0_outputs(8216) <= (inputs(148)) xor (inputs(181));
    layer0_outputs(8217) <= (inputs(79)) or (inputs(93));
    layer0_outputs(8218) <= '1';
    layer0_outputs(8219) <= not(inputs(62)) or (inputs(45));
    layer0_outputs(8220) <= not((inputs(222)) or (inputs(231)));
    layer0_outputs(8221) <= not((inputs(134)) xor (inputs(241)));
    layer0_outputs(8222) <= (inputs(141)) xor (inputs(17));
    layer0_outputs(8223) <= (inputs(222)) and not (inputs(217));
    layer0_outputs(8224) <= not((inputs(71)) xor (inputs(160)));
    layer0_outputs(8225) <= not((inputs(237)) or (inputs(18)));
    layer0_outputs(8226) <= inputs(83);
    layer0_outputs(8227) <= inputs(155);
    layer0_outputs(8228) <= not(inputs(111)) or (inputs(211));
    layer0_outputs(8229) <= (inputs(210)) or (inputs(26));
    layer0_outputs(8230) <= not((inputs(91)) or (inputs(48)));
    layer0_outputs(8231) <= inputs(93);
    layer0_outputs(8232) <= not((inputs(198)) xor (inputs(92)));
    layer0_outputs(8233) <= inputs(94);
    layer0_outputs(8234) <= inputs(151);
    layer0_outputs(8235) <= (inputs(126)) and (inputs(108));
    layer0_outputs(8236) <= not((inputs(123)) xor (inputs(248)));
    layer0_outputs(8237) <= not(inputs(110));
    layer0_outputs(8238) <= not((inputs(225)) and (inputs(19)));
    layer0_outputs(8239) <= not(inputs(41));
    layer0_outputs(8240) <= (inputs(24)) and not (inputs(102));
    layer0_outputs(8241) <= inputs(21);
    layer0_outputs(8242) <= (inputs(119)) and not (inputs(193));
    layer0_outputs(8243) <= (inputs(246)) and not (inputs(254));
    layer0_outputs(8244) <= inputs(164);
    layer0_outputs(8245) <= not((inputs(131)) or (inputs(212)));
    layer0_outputs(8246) <= not((inputs(184)) xor (inputs(154)));
    layer0_outputs(8247) <= not(inputs(22));
    layer0_outputs(8248) <= not(inputs(173));
    layer0_outputs(8249) <= (inputs(96)) xor (inputs(183));
    layer0_outputs(8250) <= (inputs(27)) xor (inputs(78));
    layer0_outputs(8251) <= not((inputs(43)) or (inputs(11)));
    layer0_outputs(8252) <= not((inputs(12)) or (inputs(3)));
    layer0_outputs(8253) <= (inputs(40)) and not (inputs(149));
    layer0_outputs(8254) <= (inputs(117)) and not (inputs(233));
    layer0_outputs(8255) <= (inputs(95)) or (inputs(213));
    layer0_outputs(8256) <= not((inputs(230)) and (inputs(11)));
    layer0_outputs(8257) <= inputs(13);
    layer0_outputs(8258) <= not((inputs(2)) xor (inputs(223)));
    layer0_outputs(8259) <= not(inputs(58));
    layer0_outputs(8260) <= not(inputs(138)) or (inputs(8));
    layer0_outputs(8261) <= (inputs(25)) and not (inputs(161));
    layer0_outputs(8262) <= not(inputs(153));
    layer0_outputs(8263) <= (inputs(244)) and not (inputs(144));
    layer0_outputs(8264) <= (inputs(137)) and not (inputs(141));
    layer0_outputs(8265) <= not(inputs(229));
    layer0_outputs(8266) <= not((inputs(67)) or (inputs(98)));
    layer0_outputs(8267) <= not(inputs(14));
    layer0_outputs(8268) <= not((inputs(32)) or (inputs(37)));
    layer0_outputs(8269) <= (inputs(3)) and not (inputs(126));
    layer0_outputs(8270) <= inputs(93);
    layer0_outputs(8271) <= (inputs(167)) and (inputs(214));
    layer0_outputs(8272) <= (inputs(16)) or (inputs(12));
    layer0_outputs(8273) <= not(inputs(86)) or (inputs(236));
    layer0_outputs(8274) <= not((inputs(20)) or (inputs(155)));
    layer0_outputs(8275) <= not((inputs(69)) and (inputs(69)));
    layer0_outputs(8276) <= (inputs(194)) xor (inputs(165));
    layer0_outputs(8277) <= (inputs(22)) or (inputs(32));
    layer0_outputs(8278) <= not(inputs(126));
    layer0_outputs(8279) <= not(inputs(248)) or (inputs(131));
    layer0_outputs(8280) <= not((inputs(192)) xor (inputs(234)));
    layer0_outputs(8281) <= not(inputs(40)) or (inputs(111));
    layer0_outputs(8282) <= inputs(22);
    layer0_outputs(8283) <= '0';
    layer0_outputs(8284) <= (inputs(45)) xor (inputs(117));
    layer0_outputs(8285) <= not(inputs(41)) or (inputs(134));
    layer0_outputs(8286) <= not((inputs(246)) xor (inputs(52)));
    layer0_outputs(8287) <= (inputs(246)) and not (inputs(166));
    layer0_outputs(8288) <= not((inputs(11)) xor (inputs(152)));
    layer0_outputs(8289) <= not(inputs(228)) or (inputs(15));
    layer0_outputs(8290) <= inputs(74);
    layer0_outputs(8291) <= not(inputs(203));
    layer0_outputs(8292) <= (inputs(215)) and not (inputs(239));
    layer0_outputs(8293) <= not((inputs(52)) xor (inputs(72)));
    layer0_outputs(8294) <= (inputs(200)) or (inputs(50));
    layer0_outputs(8295) <= (inputs(216)) xor (inputs(57));
    layer0_outputs(8296) <= not(inputs(93));
    layer0_outputs(8297) <= not((inputs(186)) or (inputs(36)));
    layer0_outputs(8298) <= inputs(4);
    layer0_outputs(8299) <= not((inputs(223)) xor (inputs(219)));
    layer0_outputs(8300) <= (inputs(98)) or (inputs(74));
    layer0_outputs(8301) <= not((inputs(135)) xor (inputs(196)));
    layer0_outputs(8302) <= not(inputs(178));
    layer0_outputs(8303) <= not((inputs(199)) xor (inputs(215)));
    layer0_outputs(8304) <= not((inputs(93)) xor (inputs(199)));
    layer0_outputs(8305) <= not((inputs(227)) xor (inputs(166)));
    layer0_outputs(8306) <= not((inputs(161)) xor (inputs(66)));
    layer0_outputs(8307) <= (inputs(246)) and not (inputs(239));
    layer0_outputs(8308) <= not((inputs(189)) or (inputs(52)));
    layer0_outputs(8309) <= inputs(40);
    layer0_outputs(8310) <= (inputs(82)) and not (inputs(16));
    layer0_outputs(8311) <= not((inputs(3)) or (inputs(24)));
    layer0_outputs(8312) <= not((inputs(35)) xor (inputs(160)));
    layer0_outputs(8313) <= (inputs(93)) xor (inputs(33));
    layer0_outputs(8314) <= not(inputs(146)) or (inputs(74));
    layer0_outputs(8315) <= (inputs(202)) and (inputs(13));
    layer0_outputs(8316) <= not(inputs(42));
    layer0_outputs(8317) <= (inputs(235)) or (inputs(144));
    layer0_outputs(8318) <= (inputs(125)) xor (inputs(6));
    layer0_outputs(8319) <= (inputs(69)) or (inputs(236));
    layer0_outputs(8320) <= (inputs(159)) or (inputs(214));
    layer0_outputs(8321) <= not((inputs(151)) xor (inputs(171)));
    layer0_outputs(8322) <= not(inputs(25));
    layer0_outputs(8323) <= (inputs(232)) xor (inputs(95));
    layer0_outputs(8324) <= not((inputs(18)) or (inputs(20)));
    layer0_outputs(8325) <= not((inputs(204)) xor (inputs(158)));
    layer0_outputs(8326) <= not((inputs(173)) xor (inputs(178)));
    layer0_outputs(8327) <= not(inputs(54));
    layer0_outputs(8328) <= not((inputs(20)) xor (inputs(210)));
    layer0_outputs(8329) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(8330) <= inputs(88);
    layer0_outputs(8331) <= inputs(99);
    layer0_outputs(8332) <= (inputs(245)) xor (inputs(153));
    layer0_outputs(8333) <= not(inputs(119));
    layer0_outputs(8334) <= inputs(194);
    layer0_outputs(8335) <= (inputs(46)) xor (inputs(192));
    layer0_outputs(8336) <= (inputs(64)) or (inputs(253));
    layer0_outputs(8337) <= inputs(90);
    layer0_outputs(8338) <= (inputs(196)) and not (inputs(97));
    layer0_outputs(8339) <= not(inputs(63)) or (inputs(65));
    layer0_outputs(8340) <= not(inputs(135)) or (inputs(100));
    layer0_outputs(8341) <= (inputs(99)) and not (inputs(206));
    layer0_outputs(8342) <= not(inputs(42)) or (inputs(176));
    layer0_outputs(8343) <= (inputs(85)) and not (inputs(204));
    layer0_outputs(8344) <= not((inputs(239)) or (inputs(83)));
    layer0_outputs(8345) <= (inputs(73)) and not (inputs(237));
    layer0_outputs(8346) <= inputs(167);
    layer0_outputs(8347) <= inputs(61);
    layer0_outputs(8348) <= not(inputs(23)) or (inputs(208));
    layer0_outputs(8349) <= inputs(67);
    layer0_outputs(8350) <= not(inputs(118));
    layer0_outputs(8351) <= (inputs(161)) xor (inputs(197));
    layer0_outputs(8352) <= not(inputs(61)) or (inputs(243));
    layer0_outputs(8353) <= inputs(71);
    layer0_outputs(8354) <= not(inputs(4));
    layer0_outputs(8355) <= not(inputs(221));
    layer0_outputs(8356) <= not((inputs(146)) or (inputs(51)));
    layer0_outputs(8357) <= (inputs(20)) or (inputs(63));
    layer0_outputs(8358) <= not(inputs(67));
    layer0_outputs(8359) <= inputs(76);
    layer0_outputs(8360) <= (inputs(88)) xor (inputs(223));
    layer0_outputs(8361) <= (inputs(227)) and not (inputs(86));
    layer0_outputs(8362) <= not((inputs(253)) or (inputs(185)));
    layer0_outputs(8363) <= not(inputs(212));
    layer0_outputs(8364) <= not((inputs(203)) or (inputs(242)));
    layer0_outputs(8365) <= not(inputs(193)) or (inputs(31));
    layer0_outputs(8366) <= not((inputs(189)) xor (inputs(155)));
    layer0_outputs(8367) <= (inputs(64)) or (inputs(210));
    layer0_outputs(8368) <= inputs(230);
    layer0_outputs(8369) <= inputs(66);
    layer0_outputs(8370) <= not((inputs(148)) or (inputs(128)));
    layer0_outputs(8371) <= inputs(199);
    layer0_outputs(8372) <= not(inputs(101));
    layer0_outputs(8373) <= (inputs(91)) xor (inputs(150));
    layer0_outputs(8374) <= (inputs(199)) and not (inputs(61));
    layer0_outputs(8375) <= not(inputs(163));
    layer0_outputs(8376) <= not(inputs(86));
    layer0_outputs(8377) <= inputs(168);
    layer0_outputs(8378) <= (inputs(207)) or (inputs(26));
    layer0_outputs(8379) <= not(inputs(135));
    layer0_outputs(8380) <= not(inputs(154)) or (inputs(80));
    layer0_outputs(8381) <= not(inputs(97));
    layer0_outputs(8382) <= inputs(18);
    layer0_outputs(8383) <= not(inputs(103)) or (inputs(98));
    layer0_outputs(8384) <= not(inputs(133)) or (inputs(78));
    layer0_outputs(8385) <= not((inputs(113)) and (inputs(144)));
    layer0_outputs(8386) <= not((inputs(116)) xor (inputs(120)));
    layer0_outputs(8387) <= (inputs(30)) xor (inputs(128));
    layer0_outputs(8388) <= not((inputs(7)) or (inputs(116)));
    layer0_outputs(8389) <= not((inputs(211)) or (inputs(194)));
    layer0_outputs(8390) <= not((inputs(221)) or (inputs(103)));
    layer0_outputs(8391) <= (inputs(75)) and not (inputs(111));
    layer0_outputs(8392) <= (inputs(144)) xor (inputs(69));
    layer0_outputs(8393) <= not(inputs(227));
    layer0_outputs(8394) <= (inputs(139)) and not (inputs(62));
    layer0_outputs(8395) <= not((inputs(228)) xor (inputs(162)));
    layer0_outputs(8396) <= not((inputs(159)) or (inputs(174)));
    layer0_outputs(8397) <= not((inputs(85)) xor (inputs(82)));
    layer0_outputs(8398) <= not((inputs(35)) or (inputs(110)));
    layer0_outputs(8399) <= not((inputs(113)) xor (inputs(58)));
    layer0_outputs(8400) <= (inputs(194)) or (inputs(2));
    layer0_outputs(8401) <= (inputs(218)) or (inputs(201));
    layer0_outputs(8402) <= not(inputs(217)) or (inputs(96));
    layer0_outputs(8403) <= (inputs(255)) and not (inputs(160));
    layer0_outputs(8404) <= not((inputs(140)) or (inputs(164)));
    layer0_outputs(8405) <= (inputs(228)) and not (inputs(181));
    layer0_outputs(8406) <= (inputs(32)) or (inputs(134));
    layer0_outputs(8407) <= not((inputs(201)) or (inputs(190)));
    layer0_outputs(8408) <= (inputs(58)) xor (inputs(27));
    layer0_outputs(8409) <= inputs(32);
    layer0_outputs(8410) <= (inputs(243)) or (inputs(128));
    layer0_outputs(8411) <= not(inputs(226));
    layer0_outputs(8412) <= not(inputs(103)) or (inputs(218));
    layer0_outputs(8413) <= (inputs(161)) or (inputs(198));
    layer0_outputs(8414) <= (inputs(173)) or (inputs(176));
    layer0_outputs(8415) <= inputs(66);
    layer0_outputs(8416) <= inputs(21);
    layer0_outputs(8417) <= not(inputs(6));
    layer0_outputs(8418) <= (inputs(174)) or (inputs(208));
    layer0_outputs(8419) <= (inputs(116)) and not (inputs(31));
    layer0_outputs(8420) <= (inputs(95)) xor (inputs(181));
    layer0_outputs(8421) <= (inputs(175)) xor (inputs(238));
    layer0_outputs(8422) <= inputs(7);
    layer0_outputs(8423) <= not(inputs(100)) or (inputs(165));
    layer0_outputs(8424) <= inputs(53);
    layer0_outputs(8425) <= (inputs(14)) or (inputs(219));
    layer0_outputs(8426) <= not(inputs(160)) or (inputs(48));
    layer0_outputs(8427) <= not((inputs(44)) or (inputs(14)));
    layer0_outputs(8428) <= (inputs(195)) and (inputs(152));
    layer0_outputs(8429) <= not((inputs(153)) xor (inputs(137)));
    layer0_outputs(8430) <= (inputs(193)) or (inputs(196));
    layer0_outputs(8431) <= not((inputs(154)) xor (inputs(106)));
    layer0_outputs(8432) <= (inputs(80)) xor (inputs(27));
    layer0_outputs(8433) <= (inputs(106)) and not (inputs(255));
    layer0_outputs(8434) <= not((inputs(116)) or (inputs(154)));
    layer0_outputs(8435) <= not(inputs(84)) or (inputs(154));
    layer0_outputs(8436) <= (inputs(200)) and not (inputs(59));
    layer0_outputs(8437) <= (inputs(46)) and not (inputs(127));
    layer0_outputs(8438) <= inputs(213);
    layer0_outputs(8439) <= (inputs(10)) and not (inputs(97));
    layer0_outputs(8440) <= inputs(223);
    layer0_outputs(8441) <= not((inputs(174)) xor (inputs(161)));
    layer0_outputs(8442) <= (inputs(160)) and (inputs(14));
    layer0_outputs(8443) <= (inputs(97)) or (inputs(222));
    layer0_outputs(8444) <= (inputs(13)) or (inputs(34));
    layer0_outputs(8445) <= not((inputs(59)) or (inputs(79)));
    layer0_outputs(8446) <= not((inputs(231)) or (inputs(249)));
    layer0_outputs(8447) <= (inputs(165)) and (inputs(186));
    layer0_outputs(8448) <= (inputs(139)) or (inputs(158));
    layer0_outputs(8449) <= (inputs(130)) and (inputs(134));
    layer0_outputs(8450) <= inputs(22);
    layer0_outputs(8451) <= not((inputs(207)) or (inputs(125)));
    layer0_outputs(8452) <= not((inputs(198)) or (inputs(117)));
    layer0_outputs(8453) <= not(inputs(228));
    layer0_outputs(8454) <= not((inputs(54)) or (inputs(98)));
    layer0_outputs(8455) <= inputs(63);
    layer0_outputs(8456) <= (inputs(207)) xor (inputs(156));
    layer0_outputs(8457) <= (inputs(143)) or (inputs(221));
    layer0_outputs(8458) <= not(inputs(60)) or (inputs(32));
    layer0_outputs(8459) <= inputs(163);
    layer0_outputs(8460) <= not((inputs(80)) and (inputs(80)));
    layer0_outputs(8461) <= (inputs(25)) or (inputs(64));
    layer0_outputs(8462) <= not(inputs(7)) or (inputs(145));
    layer0_outputs(8463) <= not(inputs(81));
    layer0_outputs(8464) <= not((inputs(29)) or (inputs(113)));
    layer0_outputs(8465) <= inputs(122);
    layer0_outputs(8466) <= inputs(213);
    layer0_outputs(8467) <= (inputs(99)) and not (inputs(62));
    layer0_outputs(8468) <= not((inputs(154)) and (inputs(216)));
    layer0_outputs(8469) <= not(inputs(67));
    layer0_outputs(8470) <= not(inputs(159)) or (inputs(206));
    layer0_outputs(8471) <= not(inputs(87));
    layer0_outputs(8472) <= (inputs(186)) and not (inputs(93));
    layer0_outputs(8473) <= (inputs(104)) and not (inputs(253));
    layer0_outputs(8474) <= not((inputs(184)) xor (inputs(185)));
    layer0_outputs(8475) <= not(inputs(178));
    layer0_outputs(8476) <= (inputs(230)) and not (inputs(124));
    layer0_outputs(8477) <= not((inputs(72)) xor (inputs(130)));
    layer0_outputs(8478) <= not(inputs(245));
    layer0_outputs(8479) <= (inputs(135)) and not (inputs(125));
    layer0_outputs(8480) <= (inputs(50)) and not (inputs(150));
    layer0_outputs(8481) <= not((inputs(63)) or (inputs(61)));
    layer0_outputs(8482) <= not(inputs(31)) or (inputs(190));
    layer0_outputs(8483) <= inputs(216);
    layer0_outputs(8484) <= (inputs(70)) or (inputs(131));
    layer0_outputs(8485) <= not(inputs(90)) or (inputs(176));
    layer0_outputs(8486) <= not((inputs(181)) or (inputs(244)));
    layer0_outputs(8487) <= (inputs(50)) and not (inputs(112));
    layer0_outputs(8488) <= (inputs(58)) and not (inputs(211));
    layer0_outputs(8489) <= not((inputs(111)) or (inputs(21)));
    layer0_outputs(8490) <= (inputs(12)) xor (inputs(208));
    layer0_outputs(8491) <= not(inputs(135)) or (inputs(66));
    layer0_outputs(8492) <= (inputs(98)) and not (inputs(162));
    layer0_outputs(8493) <= inputs(114);
    layer0_outputs(8494) <= not((inputs(173)) or (inputs(148)));
    layer0_outputs(8495) <= not(inputs(98)) or (inputs(25));
    layer0_outputs(8496) <= (inputs(55)) or (inputs(179));
    layer0_outputs(8497) <= not(inputs(158)) or (inputs(224));
    layer0_outputs(8498) <= not(inputs(20));
    layer0_outputs(8499) <= (inputs(20)) and not (inputs(161));
    layer0_outputs(8500) <= not(inputs(210));
    layer0_outputs(8501) <= not((inputs(66)) xor (inputs(209)));
    layer0_outputs(8502) <= (inputs(28)) or (inputs(49));
    layer0_outputs(8503) <= inputs(168);
    layer0_outputs(8504) <= '1';
    layer0_outputs(8505) <= not((inputs(162)) xor (inputs(214)));
    layer0_outputs(8506) <= not(inputs(201));
    layer0_outputs(8507) <= (inputs(67)) or (inputs(61));
    layer0_outputs(8508) <= inputs(231);
    layer0_outputs(8509) <= inputs(209);
    layer0_outputs(8510) <= not(inputs(81));
    layer0_outputs(8511) <= inputs(89);
    layer0_outputs(8512) <= inputs(96);
    layer0_outputs(8513) <= inputs(71);
    layer0_outputs(8514) <= (inputs(78)) or (inputs(126));
    layer0_outputs(8515) <= (inputs(251)) and not (inputs(232));
    layer0_outputs(8516) <= (inputs(138)) xor (inputs(242));
    layer0_outputs(8517) <= (inputs(167)) xor (inputs(106));
    layer0_outputs(8518) <= '1';
    layer0_outputs(8519) <= (inputs(248)) or (inputs(146));
    layer0_outputs(8520) <= inputs(208);
    layer0_outputs(8521) <= inputs(54);
    layer0_outputs(8522) <= (inputs(191)) xor (inputs(119));
    layer0_outputs(8523) <= (inputs(144)) or (inputs(70));
    layer0_outputs(8524) <= '0';
    layer0_outputs(8525) <= (inputs(144)) xor (inputs(176));
    layer0_outputs(8526) <= not((inputs(117)) or (inputs(226)));
    layer0_outputs(8527) <= not((inputs(189)) or (inputs(41)));
    layer0_outputs(8528) <= not(inputs(21));
    layer0_outputs(8529) <= not(inputs(7)) or (inputs(204));
    layer0_outputs(8530) <= (inputs(132)) and not (inputs(3));
    layer0_outputs(8531) <= not(inputs(231));
    layer0_outputs(8532) <= not((inputs(6)) xor (inputs(209)));
    layer0_outputs(8533) <= (inputs(231)) and (inputs(230));
    layer0_outputs(8534) <= not(inputs(52));
    layer0_outputs(8535) <= not((inputs(220)) or (inputs(145)));
    layer0_outputs(8536) <= (inputs(240)) or (inputs(146));
    layer0_outputs(8537) <= (inputs(29)) xor (inputs(81));
    layer0_outputs(8538) <= (inputs(121)) and not (inputs(215));
    layer0_outputs(8539) <= not(inputs(24)) or (inputs(147));
    layer0_outputs(8540) <= not(inputs(122)) or (inputs(249));
    layer0_outputs(8541) <= not((inputs(114)) and (inputs(121)));
    layer0_outputs(8542) <= inputs(104);
    layer0_outputs(8543) <= not((inputs(131)) xor (inputs(99)));
    layer0_outputs(8544) <= inputs(153);
    layer0_outputs(8545) <= not((inputs(163)) xor (inputs(212)));
    layer0_outputs(8546) <= not(inputs(82)) or (inputs(93));
    layer0_outputs(8547) <= (inputs(116)) or (inputs(35));
    layer0_outputs(8548) <= (inputs(219)) and (inputs(151));
    layer0_outputs(8549) <= not(inputs(131));
    layer0_outputs(8550) <= (inputs(136)) xor (inputs(123));
    layer0_outputs(8551) <= (inputs(93)) and not (inputs(254));
    layer0_outputs(8552) <= not((inputs(187)) xor (inputs(62)));
    layer0_outputs(8553) <= not((inputs(35)) xor (inputs(142)));
    layer0_outputs(8554) <= (inputs(96)) or (inputs(201));
    layer0_outputs(8555) <= not(inputs(120)) or (inputs(200));
    layer0_outputs(8556) <= inputs(147);
    layer0_outputs(8557) <= not(inputs(199)) or (inputs(47));
    layer0_outputs(8558) <= not(inputs(138)) or (inputs(234));
    layer0_outputs(8559) <= not(inputs(69)) or (inputs(125));
    layer0_outputs(8560) <= (inputs(212)) xor (inputs(242));
    layer0_outputs(8561) <= (inputs(25)) and (inputs(122));
    layer0_outputs(8562) <= inputs(24);
    layer0_outputs(8563) <= not((inputs(12)) xor (inputs(255)));
    layer0_outputs(8564) <= (inputs(72)) xor (inputs(83));
    layer0_outputs(8565) <= inputs(167);
    layer0_outputs(8566) <= not(inputs(221));
    layer0_outputs(8567) <= (inputs(3)) xor (inputs(81));
    layer0_outputs(8568) <= (inputs(105)) and (inputs(77));
    layer0_outputs(8569) <= not(inputs(106));
    layer0_outputs(8570) <= not(inputs(202)) or (inputs(20));
    layer0_outputs(8571) <= (inputs(227)) xor (inputs(158));
    layer0_outputs(8572) <= (inputs(65)) and not (inputs(21));
    layer0_outputs(8573) <= (inputs(9)) xor (inputs(89));
    layer0_outputs(8574) <= (inputs(125)) or (inputs(83));
    layer0_outputs(8575) <= inputs(90);
    layer0_outputs(8576) <= not((inputs(33)) or (inputs(56)));
    layer0_outputs(8577) <= (inputs(166)) and not (inputs(144));
    layer0_outputs(8578) <= inputs(236);
    layer0_outputs(8579) <= not(inputs(114));
    layer0_outputs(8580) <= not(inputs(181)) or (inputs(34));
    layer0_outputs(8581) <= (inputs(114)) and not (inputs(207));
    layer0_outputs(8582) <= not((inputs(12)) or (inputs(96)));
    layer0_outputs(8583) <= inputs(254);
    layer0_outputs(8584) <= not((inputs(87)) and (inputs(39)));
    layer0_outputs(8585) <= not(inputs(11));
    layer0_outputs(8586) <= not((inputs(200)) and (inputs(184)));
    layer0_outputs(8587) <= not(inputs(75));
    layer0_outputs(8588) <= (inputs(158)) xor (inputs(137));
    layer0_outputs(8589) <= not(inputs(57));
    layer0_outputs(8590) <= (inputs(44)) and (inputs(236));
    layer0_outputs(8591) <= not((inputs(43)) or (inputs(242)));
    layer0_outputs(8592) <= (inputs(161)) and not (inputs(122));
    layer0_outputs(8593) <= (inputs(125)) or (inputs(79));
    layer0_outputs(8594) <= inputs(33);
    layer0_outputs(8595) <= (inputs(234)) xor (inputs(147));
    layer0_outputs(8596) <= (inputs(211)) and not (inputs(113));
    layer0_outputs(8597) <= (inputs(187)) xor (inputs(190));
    layer0_outputs(8598) <= (inputs(252)) or (inputs(87));
    layer0_outputs(8599) <= not(inputs(168));
    layer0_outputs(8600) <= inputs(69);
    layer0_outputs(8601) <= not((inputs(246)) or (inputs(20)));
    layer0_outputs(8602) <= inputs(13);
    layer0_outputs(8603) <= inputs(136);
    layer0_outputs(8604) <= (inputs(189)) and not (inputs(253));
    layer0_outputs(8605) <= (inputs(35)) xor (inputs(170));
    layer0_outputs(8606) <= (inputs(176)) or (inputs(79));
    layer0_outputs(8607) <= not((inputs(161)) or (inputs(127)));
    layer0_outputs(8608) <= (inputs(211)) and not (inputs(102));
    layer0_outputs(8609) <= inputs(97);
    layer0_outputs(8610) <= (inputs(183)) xor (inputs(188));
    layer0_outputs(8611) <= (inputs(173)) and not (inputs(99));
    layer0_outputs(8612) <= (inputs(73)) and not (inputs(0));
    layer0_outputs(8613) <= not((inputs(114)) xor (inputs(24)));
    layer0_outputs(8614) <= not((inputs(226)) xor (inputs(215)));
    layer0_outputs(8615) <= not(inputs(212)) or (inputs(156));
    layer0_outputs(8616) <= (inputs(3)) or (inputs(29));
    layer0_outputs(8617) <= not((inputs(159)) or (inputs(77)));
    layer0_outputs(8618) <= not(inputs(83));
    layer0_outputs(8619) <= not(inputs(151));
    layer0_outputs(8620) <= (inputs(195)) or (inputs(4));
    layer0_outputs(8621) <= not((inputs(120)) or (inputs(146)));
    layer0_outputs(8622) <= not((inputs(137)) xor (inputs(205)));
    layer0_outputs(8623) <= not(inputs(134));
    layer0_outputs(8624) <= not(inputs(13));
    layer0_outputs(8625) <= not((inputs(35)) or (inputs(241)));
    layer0_outputs(8626) <= inputs(99);
    layer0_outputs(8627) <= not(inputs(228));
    layer0_outputs(8628) <= not(inputs(75)) or (inputs(254));
    layer0_outputs(8629) <= not((inputs(52)) xor (inputs(21)));
    layer0_outputs(8630) <= inputs(71);
    layer0_outputs(8631) <= inputs(148);
    layer0_outputs(8632) <= (inputs(177)) and not (inputs(155));
    layer0_outputs(8633) <= inputs(107);
    layer0_outputs(8634) <= not(inputs(78));
    layer0_outputs(8635) <= not((inputs(208)) or (inputs(174)));
    layer0_outputs(8636) <= not((inputs(14)) or (inputs(205)));
    layer0_outputs(8637) <= not(inputs(168)) or (inputs(73));
    layer0_outputs(8638) <= (inputs(16)) or (inputs(39));
    layer0_outputs(8639) <= not(inputs(105));
    layer0_outputs(8640) <= (inputs(233)) or (inputs(116));
    layer0_outputs(8641) <= inputs(91);
    layer0_outputs(8642) <= not(inputs(87));
    layer0_outputs(8643) <= (inputs(224)) xor (inputs(27));
    layer0_outputs(8644) <= not((inputs(43)) xor (inputs(225)));
    layer0_outputs(8645) <= (inputs(79)) or (inputs(27));
    layer0_outputs(8646) <= (inputs(115)) or (inputs(42));
    layer0_outputs(8647) <= inputs(94);
    layer0_outputs(8648) <= not((inputs(203)) xor (inputs(132)));
    layer0_outputs(8649) <= inputs(111);
    layer0_outputs(8650) <= (inputs(46)) xor (inputs(103));
    layer0_outputs(8651) <= not((inputs(34)) xor (inputs(169)));
    layer0_outputs(8652) <= not(inputs(58));
    layer0_outputs(8653) <= not(inputs(157)) or (inputs(225));
    layer0_outputs(8654) <= not((inputs(106)) or (inputs(242)));
    layer0_outputs(8655) <= (inputs(229)) or (inputs(208));
    layer0_outputs(8656) <= not(inputs(88));
    layer0_outputs(8657) <= (inputs(138)) xor (inputs(185));
    layer0_outputs(8658) <= (inputs(154)) or (inputs(250));
    layer0_outputs(8659) <= (inputs(3)) and not (inputs(26));
    layer0_outputs(8660) <= (inputs(21)) and not (inputs(124));
    layer0_outputs(8661) <= not(inputs(120)) or (inputs(41));
    layer0_outputs(8662) <= inputs(253);
    layer0_outputs(8663) <= not(inputs(214));
    layer0_outputs(8664) <= not(inputs(67));
    layer0_outputs(8665) <= inputs(179);
    layer0_outputs(8666) <= inputs(34);
    layer0_outputs(8667) <= not(inputs(123)) or (inputs(205));
    layer0_outputs(8668) <= not(inputs(199)) or (inputs(43));
    layer0_outputs(8669) <= (inputs(24)) or (inputs(17));
    layer0_outputs(8670) <= inputs(32);
    layer0_outputs(8671) <= inputs(170);
    layer0_outputs(8672) <= not(inputs(160));
    layer0_outputs(8673) <= not(inputs(78)) or (inputs(249));
    layer0_outputs(8674) <= not((inputs(249)) xor (inputs(72)));
    layer0_outputs(8675) <= not((inputs(176)) xor (inputs(220)));
    layer0_outputs(8676) <= not((inputs(91)) and (inputs(135)));
    layer0_outputs(8677) <= '0';
    layer0_outputs(8678) <= (inputs(218)) or (inputs(116));
    layer0_outputs(8679) <= not((inputs(50)) xor (inputs(69)));
    layer0_outputs(8680) <= inputs(139);
    layer0_outputs(8681) <= not(inputs(157));
    layer0_outputs(8682) <= not((inputs(16)) xor (inputs(91)));
    layer0_outputs(8683) <= not(inputs(117)) or (inputs(5));
    layer0_outputs(8684) <= (inputs(12)) and not (inputs(226));
    layer0_outputs(8685) <= not(inputs(27));
    layer0_outputs(8686) <= not((inputs(127)) or (inputs(184)));
    layer0_outputs(8687) <= inputs(75);
    layer0_outputs(8688) <= not((inputs(4)) or (inputs(225)));
    layer0_outputs(8689) <= not((inputs(73)) and (inputs(67)));
    layer0_outputs(8690) <= inputs(164);
    layer0_outputs(8691) <= inputs(28);
    layer0_outputs(8692) <= (inputs(245)) xor (inputs(206));
    layer0_outputs(8693) <= not((inputs(189)) or (inputs(255)));
    layer0_outputs(8694) <= not((inputs(84)) or (inputs(205)));
    layer0_outputs(8695) <= (inputs(213)) and not (inputs(36));
    layer0_outputs(8696) <= (inputs(88)) xor (inputs(156));
    layer0_outputs(8697) <= inputs(85);
    layer0_outputs(8698) <= (inputs(109)) xor (inputs(127));
    layer0_outputs(8699) <= inputs(249);
    layer0_outputs(8700) <= not(inputs(58));
    layer0_outputs(8701) <= (inputs(66)) or (inputs(189));
    layer0_outputs(8702) <= (inputs(82)) and not (inputs(54));
    layer0_outputs(8703) <= inputs(230);
    layer0_outputs(8704) <= not((inputs(5)) or (inputs(228)));
    layer0_outputs(8705) <= (inputs(228)) and not (inputs(223));
    layer0_outputs(8706) <= not(inputs(53)) or (inputs(235));
    layer0_outputs(8707) <= not(inputs(6)) or (inputs(240));
    layer0_outputs(8708) <= not((inputs(107)) xor (inputs(91)));
    layer0_outputs(8709) <= not((inputs(28)) and (inputs(138)));
    layer0_outputs(8710) <= not((inputs(172)) or (inputs(90)));
    layer0_outputs(8711) <= inputs(181);
    layer0_outputs(8712) <= not(inputs(173));
    layer0_outputs(8713) <= (inputs(26)) or (inputs(193));
    layer0_outputs(8714) <= not((inputs(18)) or (inputs(12)));
    layer0_outputs(8715) <= not((inputs(165)) xor (inputs(47)));
    layer0_outputs(8716) <= (inputs(21)) xor (inputs(189));
    layer0_outputs(8717) <= not(inputs(241)) or (inputs(27));
    layer0_outputs(8718) <= not(inputs(215)) or (inputs(69));
    layer0_outputs(8719) <= not(inputs(106)) or (inputs(160));
    layer0_outputs(8720) <= inputs(54);
    layer0_outputs(8721) <= not(inputs(217));
    layer0_outputs(8722) <= not(inputs(50));
    layer0_outputs(8723) <= not(inputs(108)) or (inputs(89));
    layer0_outputs(8724) <= (inputs(217)) or (inputs(133));
    layer0_outputs(8725) <= not((inputs(201)) and (inputs(229)));
    layer0_outputs(8726) <= not((inputs(131)) xor (inputs(185)));
    layer0_outputs(8727) <= not(inputs(147));
    layer0_outputs(8728) <= not((inputs(55)) and (inputs(82)));
    layer0_outputs(8729) <= not((inputs(229)) xor (inputs(133)));
    layer0_outputs(8730) <= inputs(104);
    layer0_outputs(8731) <= (inputs(239)) or (inputs(220));
    layer0_outputs(8732) <= not(inputs(146)) or (inputs(152));
    layer0_outputs(8733) <= (inputs(211)) or (inputs(235));
    layer0_outputs(8734) <= (inputs(115)) and not (inputs(48));
    layer0_outputs(8735) <= (inputs(197)) and (inputs(201));
    layer0_outputs(8736) <= not(inputs(101)) or (inputs(64));
    layer0_outputs(8737) <= not(inputs(108));
    layer0_outputs(8738) <= (inputs(130)) or (inputs(131));
    layer0_outputs(8739) <= inputs(198);
    layer0_outputs(8740) <= not(inputs(222)) or (inputs(203));
    layer0_outputs(8741) <= (inputs(53)) or (inputs(59));
    layer0_outputs(8742) <= '1';
    layer0_outputs(8743) <= (inputs(133)) xor (inputs(140));
    layer0_outputs(8744) <= (inputs(130)) or (inputs(62));
    layer0_outputs(8745) <= (inputs(97)) or (inputs(145));
    layer0_outputs(8746) <= (inputs(79)) or (inputs(104));
    layer0_outputs(8747) <= (inputs(232)) and not (inputs(128));
    layer0_outputs(8748) <= not(inputs(122)) or (inputs(199));
    layer0_outputs(8749) <= not((inputs(186)) xor (inputs(98)));
    layer0_outputs(8750) <= (inputs(58)) and not (inputs(94));
    layer0_outputs(8751) <= (inputs(193)) or (inputs(216));
    layer0_outputs(8752) <= not(inputs(101)) or (inputs(215));
    layer0_outputs(8753) <= (inputs(244)) and not (inputs(53));
    layer0_outputs(8754) <= not((inputs(20)) or (inputs(180)));
    layer0_outputs(8755) <= (inputs(10)) and not (inputs(16));
    layer0_outputs(8756) <= (inputs(224)) and (inputs(16));
    layer0_outputs(8757) <= (inputs(45)) xor (inputs(166));
    layer0_outputs(8758) <= not(inputs(190));
    layer0_outputs(8759) <= not((inputs(230)) or (inputs(193)));
    layer0_outputs(8760) <= (inputs(252)) or (inputs(14));
    layer0_outputs(8761) <= (inputs(54)) and not (inputs(201));
    layer0_outputs(8762) <= inputs(189);
    layer0_outputs(8763) <= not((inputs(126)) xor (inputs(101)));
    layer0_outputs(8764) <= (inputs(213)) and not (inputs(58));
    layer0_outputs(8765) <= not(inputs(166)) or (inputs(101));
    layer0_outputs(8766) <= not(inputs(37));
    layer0_outputs(8767) <= not(inputs(24)) or (inputs(198));
    layer0_outputs(8768) <= not((inputs(49)) or (inputs(42)));
    layer0_outputs(8769) <= not((inputs(179)) or (inputs(187)));
    layer0_outputs(8770) <= not(inputs(140));
    layer0_outputs(8771) <= not(inputs(147));
    layer0_outputs(8772) <= '0';
    layer0_outputs(8773) <= not(inputs(122));
    layer0_outputs(8774) <= not(inputs(165));
    layer0_outputs(8775) <= (inputs(161)) or (inputs(146));
    layer0_outputs(8776) <= (inputs(219)) or (inputs(217));
    layer0_outputs(8777) <= (inputs(219)) and not (inputs(253));
    layer0_outputs(8778) <= not(inputs(213)) or (inputs(147));
    layer0_outputs(8779) <= (inputs(232)) or (inputs(148));
    layer0_outputs(8780) <= not(inputs(74)) or (inputs(68));
    layer0_outputs(8781) <= (inputs(7)) or (inputs(238));
    layer0_outputs(8782) <= not((inputs(93)) xor (inputs(90)));
    layer0_outputs(8783) <= not(inputs(153));
    layer0_outputs(8784) <= (inputs(237)) and not (inputs(10));
    layer0_outputs(8785) <= (inputs(253)) or (inputs(111));
    layer0_outputs(8786) <= not((inputs(17)) xor (inputs(56)));
    layer0_outputs(8787) <= (inputs(235)) and not (inputs(63));
    layer0_outputs(8788) <= not(inputs(234));
    layer0_outputs(8789) <= not(inputs(131));
    layer0_outputs(8790) <= (inputs(104)) or (inputs(251));
    layer0_outputs(8791) <= not((inputs(4)) and (inputs(237)));
    layer0_outputs(8792) <= (inputs(247)) and (inputs(118));
    layer0_outputs(8793) <= (inputs(196)) and not (inputs(33));
    layer0_outputs(8794) <= (inputs(249)) and not (inputs(17));
    layer0_outputs(8795) <= '1';
    layer0_outputs(8796) <= inputs(74);
    layer0_outputs(8797) <= not((inputs(191)) or (inputs(55)));
    layer0_outputs(8798) <= not((inputs(26)) and (inputs(85)));
    layer0_outputs(8799) <= (inputs(106)) and not (inputs(205));
    layer0_outputs(8800) <= not((inputs(142)) or (inputs(223)));
    layer0_outputs(8801) <= inputs(86);
    layer0_outputs(8802) <= (inputs(45)) and not (inputs(238));
    layer0_outputs(8803) <= (inputs(129)) or (inputs(193));
    layer0_outputs(8804) <= not(inputs(4));
    layer0_outputs(8805) <= (inputs(33)) or (inputs(21));
    layer0_outputs(8806) <= not(inputs(46));
    layer0_outputs(8807) <= not((inputs(207)) xor (inputs(94)));
    layer0_outputs(8808) <= not(inputs(28)) or (inputs(127));
    layer0_outputs(8809) <= inputs(227);
    layer0_outputs(8810) <= inputs(144);
    layer0_outputs(8811) <= (inputs(236)) and (inputs(244));
    layer0_outputs(8812) <= not(inputs(2)) or (inputs(109));
    layer0_outputs(8813) <= (inputs(154)) and not (inputs(35));
    layer0_outputs(8814) <= not(inputs(171)) or (inputs(84));
    layer0_outputs(8815) <= not((inputs(79)) or (inputs(252)));
    layer0_outputs(8816) <= not(inputs(28));
    layer0_outputs(8817) <= not(inputs(93));
    layer0_outputs(8818) <= not((inputs(15)) or (inputs(117)));
    layer0_outputs(8819) <= inputs(157);
    layer0_outputs(8820) <= inputs(85);
    layer0_outputs(8821) <= inputs(75);
    layer0_outputs(8822) <= not(inputs(124)) or (inputs(37));
    layer0_outputs(8823) <= not((inputs(201)) xor (inputs(190)));
    layer0_outputs(8824) <= (inputs(175)) or (inputs(101));
    layer0_outputs(8825) <= (inputs(39)) xor (inputs(212));
    layer0_outputs(8826) <= (inputs(8)) and not (inputs(14));
    layer0_outputs(8827) <= (inputs(85)) or (inputs(156));
    layer0_outputs(8828) <= inputs(71);
    layer0_outputs(8829) <= not(inputs(28)) or (inputs(194));
    layer0_outputs(8830) <= '1';
    layer0_outputs(8831) <= inputs(109);
    layer0_outputs(8832) <= not(inputs(102));
    layer0_outputs(8833) <= inputs(152);
    layer0_outputs(8834) <= not(inputs(242)) or (inputs(238));
    layer0_outputs(8835) <= (inputs(108)) and not (inputs(191));
    layer0_outputs(8836) <= not((inputs(43)) and (inputs(116)));
    layer0_outputs(8837) <= (inputs(205)) and not (inputs(26));
    layer0_outputs(8838) <= not((inputs(146)) xor (inputs(75)));
    layer0_outputs(8839) <= (inputs(198)) xor (inputs(197));
    layer0_outputs(8840) <= not(inputs(250)) or (inputs(36));
    layer0_outputs(8841) <= not((inputs(204)) or (inputs(1)));
    layer0_outputs(8842) <= not((inputs(154)) or (inputs(151)));
    layer0_outputs(8843) <= not((inputs(61)) xor (inputs(91)));
    layer0_outputs(8844) <= (inputs(141)) or (inputs(90));
    layer0_outputs(8845) <= not((inputs(189)) or (inputs(193)));
    layer0_outputs(8846) <= not(inputs(165));
    layer0_outputs(8847) <= not(inputs(104)) or (inputs(12));
    layer0_outputs(8848) <= not((inputs(180)) xor (inputs(77)));
    layer0_outputs(8849) <= inputs(22);
    layer0_outputs(8850) <= (inputs(163)) xor (inputs(86));
    layer0_outputs(8851) <= (inputs(216)) and not (inputs(15));
    layer0_outputs(8852) <= not((inputs(135)) or (inputs(30)));
    layer0_outputs(8853) <= not((inputs(208)) xor (inputs(70)));
    layer0_outputs(8854) <= (inputs(105)) or (inputs(209));
    layer0_outputs(8855) <= not((inputs(199)) or (inputs(186)));
    layer0_outputs(8856) <= (inputs(46)) and (inputs(195));
    layer0_outputs(8857) <= (inputs(122)) and not (inputs(15));
    layer0_outputs(8858) <= (inputs(30)) or (inputs(175));
    layer0_outputs(8859) <= not(inputs(182));
    layer0_outputs(8860) <= inputs(11);
    layer0_outputs(8861) <= inputs(60);
    layer0_outputs(8862) <= (inputs(46)) and not (inputs(71));
    layer0_outputs(8863) <= not(inputs(231)) or (inputs(126));
    layer0_outputs(8864) <= (inputs(164)) and not (inputs(64));
    layer0_outputs(8865) <= not((inputs(163)) xor (inputs(227)));
    layer0_outputs(8866) <= not(inputs(82)) or (inputs(97));
    layer0_outputs(8867) <= not((inputs(53)) or (inputs(55)));
    layer0_outputs(8868) <= not(inputs(204));
    layer0_outputs(8869) <= not(inputs(89));
    layer0_outputs(8870) <= (inputs(77)) and not (inputs(33));
    layer0_outputs(8871) <= not((inputs(16)) and (inputs(51)));
    layer0_outputs(8872) <= not((inputs(206)) and (inputs(235)));
    layer0_outputs(8873) <= not(inputs(184)) or (inputs(134));
    layer0_outputs(8874) <= not(inputs(41));
    layer0_outputs(8875) <= inputs(61);
    layer0_outputs(8876) <= (inputs(214)) and (inputs(211));
    layer0_outputs(8877) <= not(inputs(115));
    layer0_outputs(8878) <= (inputs(238)) or (inputs(150));
    layer0_outputs(8879) <= (inputs(164)) or (inputs(145));
    layer0_outputs(8880) <= inputs(67);
    layer0_outputs(8881) <= not(inputs(196)) or (inputs(15));
    layer0_outputs(8882) <= (inputs(121)) xor (inputs(151));
    layer0_outputs(8883) <= not(inputs(37));
    layer0_outputs(8884) <= not((inputs(71)) xor (inputs(10)));
    layer0_outputs(8885) <= not((inputs(255)) xor (inputs(141)));
    layer0_outputs(8886) <= (inputs(163)) or (inputs(110));
    layer0_outputs(8887) <= (inputs(233)) or (inputs(113));
    layer0_outputs(8888) <= not((inputs(94)) or (inputs(72)));
    layer0_outputs(8889) <= inputs(85);
    layer0_outputs(8890) <= (inputs(133)) or (inputs(140));
    layer0_outputs(8891) <= (inputs(140)) and not (inputs(130));
    layer0_outputs(8892) <= (inputs(147)) or (inputs(143));
    layer0_outputs(8893) <= not(inputs(3)) or (inputs(170));
    layer0_outputs(8894) <= (inputs(184)) xor (inputs(188));
    layer0_outputs(8895) <= inputs(15);
    layer0_outputs(8896) <= (inputs(119)) xor (inputs(90));
    layer0_outputs(8897) <= (inputs(44)) and not (inputs(215));
    layer0_outputs(8898) <= not(inputs(197)) or (inputs(77));
    layer0_outputs(8899) <= (inputs(5)) and not (inputs(206));
    layer0_outputs(8900) <= inputs(26);
    layer0_outputs(8901) <= not(inputs(56));
    layer0_outputs(8902) <= inputs(231);
    layer0_outputs(8903) <= not((inputs(237)) or (inputs(144)));
    layer0_outputs(8904) <= (inputs(220)) or (inputs(217));
    layer0_outputs(8905) <= (inputs(160)) xor (inputs(102));
    layer0_outputs(8906) <= not((inputs(224)) and (inputs(31)));
    layer0_outputs(8907) <= (inputs(105)) xor (inputs(139));
    layer0_outputs(8908) <= (inputs(238)) or (inputs(110));
    layer0_outputs(8909) <= (inputs(41)) and not (inputs(249));
    layer0_outputs(8910) <= '0';
    layer0_outputs(8911) <= '0';
    layer0_outputs(8912) <= not((inputs(29)) xor (inputs(151)));
    layer0_outputs(8913) <= not(inputs(187));
    layer0_outputs(8914) <= not((inputs(18)) or (inputs(37)));
    layer0_outputs(8915) <= (inputs(173)) and not (inputs(239));
    layer0_outputs(8916) <= (inputs(95)) or (inputs(145));
    layer0_outputs(8917) <= not((inputs(85)) xor (inputs(205)));
    layer0_outputs(8918) <= not(inputs(196)) or (inputs(254));
    layer0_outputs(8919) <= not(inputs(17));
    layer0_outputs(8920) <= not(inputs(20)) or (inputs(63));
    layer0_outputs(8921) <= inputs(183);
    layer0_outputs(8922) <= (inputs(171)) xor (inputs(72));
    layer0_outputs(8923) <= not((inputs(155)) xor (inputs(98)));
    layer0_outputs(8924) <= inputs(150);
    layer0_outputs(8925) <= not((inputs(193)) and (inputs(164)));
    layer0_outputs(8926) <= (inputs(49)) xor (inputs(169));
    layer0_outputs(8927) <= not(inputs(181));
    layer0_outputs(8928) <= not((inputs(210)) xor (inputs(223)));
    layer0_outputs(8929) <= not((inputs(59)) or (inputs(239)));
    layer0_outputs(8930) <= not((inputs(164)) or (inputs(110)));
    layer0_outputs(8931) <= not(inputs(234));
    layer0_outputs(8932) <= not(inputs(3)) or (inputs(101));
    layer0_outputs(8933) <= not(inputs(230));
    layer0_outputs(8934) <= not((inputs(250)) or (inputs(167)));
    layer0_outputs(8935) <= not(inputs(58)) or (inputs(20));
    layer0_outputs(8936) <= (inputs(51)) and not (inputs(142));
    layer0_outputs(8937) <= (inputs(118)) or (inputs(87));
    layer0_outputs(8938) <= inputs(215);
    layer0_outputs(8939) <= not(inputs(150));
    layer0_outputs(8940) <= not(inputs(161));
    layer0_outputs(8941) <= not(inputs(185)) or (inputs(93));
    layer0_outputs(8942) <= not((inputs(169)) and (inputs(25)));
    layer0_outputs(8943) <= not((inputs(29)) or (inputs(37)));
    layer0_outputs(8944) <= not(inputs(26));
    layer0_outputs(8945) <= inputs(78);
    layer0_outputs(8946) <= not((inputs(200)) and (inputs(88)));
    layer0_outputs(8947) <= inputs(120);
    layer0_outputs(8948) <= not((inputs(71)) xor (inputs(235)));
    layer0_outputs(8949) <= (inputs(127)) xor (inputs(148));
    layer0_outputs(8950) <= (inputs(89)) xor (inputs(181));
    layer0_outputs(8951) <= (inputs(95)) or (inputs(82));
    layer0_outputs(8952) <= not(inputs(53));
    layer0_outputs(8953) <= (inputs(64)) and not (inputs(2));
    layer0_outputs(8954) <= (inputs(159)) xor (inputs(244));
    layer0_outputs(8955) <= not((inputs(135)) or (inputs(49)));
    layer0_outputs(8956) <= not((inputs(88)) xor (inputs(117)));
    layer0_outputs(8957) <= (inputs(90)) and not (inputs(99));
    layer0_outputs(8958) <= '0';
    layer0_outputs(8959) <= not(inputs(56)) or (inputs(5));
    layer0_outputs(8960) <= not(inputs(18));
    layer0_outputs(8961) <= (inputs(240)) and not (inputs(116));
    layer0_outputs(8962) <= not(inputs(216));
    layer0_outputs(8963) <= not(inputs(246)) or (inputs(238));
    layer0_outputs(8964) <= (inputs(159)) and not (inputs(96));
    layer0_outputs(8965) <= not((inputs(90)) or (inputs(84)));
    layer0_outputs(8966) <= (inputs(232)) or (inputs(184));
    layer0_outputs(8967) <= (inputs(20)) and not (inputs(126));
    layer0_outputs(8968) <= (inputs(246)) and not (inputs(62));
    layer0_outputs(8969) <= not((inputs(10)) or (inputs(194)));
    layer0_outputs(8970) <= (inputs(149)) and not (inputs(92));
    layer0_outputs(8971) <= not(inputs(207)) or (inputs(183));
    layer0_outputs(8972) <= (inputs(137)) and not (inputs(247));
    layer0_outputs(8973) <= not(inputs(185)) or (inputs(87));
    layer0_outputs(8974) <= (inputs(144)) or (inputs(183));
    layer0_outputs(8975) <= not((inputs(72)) or (inputs(107)));
    layer0_outputs(8976) <= not((inputs(153)) xor (inputs(171)));
    layer0_outputs(8977) <= not(inputs(249));
    layer0_outputs(8978) <= (inputs(43)) and not (inputs(113));
    layer0_outputs(8979) <= not(inputs(37));
    layer0_outputs(8980) <= inputs(179);
    layer0_outputs(8981) <= (inputs(67)) or (inputs(201));
    layer0_outputs(8982) <= (inputs(253)) or (inputs(68));
    layer0_outputs(8983) <= (inputs(73)) or (inputs(179));
    layer0_outputs(8984) <= not(inputs(90));
    layer0_outputs(8985) <= not(inputs(219)) or (inputs(16));
    layer0_outputs(8986) <= (inputs(156)) or (inputs(107));
    layer0_outputs(8987) <= (inputs(119)) and not (inputs(198));
    layer0_outputs(8988) <= (inputs(93)) or (inputs(143));
    layer0_outputs(8989) <= (inputs(166)) and not (inputs(190));
    layer0_outputs(8990) <= (inputs(111)) or (inputs(35));
    layer0_outputs(8991) <= (inputs(168)) and (inputs(57));
    layer0_outputs(8992) <= inputs(18);
    layer0_outputs(8993) <= not((inputs(111)) and (inputs(187)));
    layer0_outputs(8994) <= not((inputs(109)) or (inputs(118)));
    layer0_outputs(8995) <= not(inputs(217));
    layer0_outputs(8996) <= not((inputs(28)) and (inputs(91)));
    layer0_outputs(8997) <= not(inputs(235));
    layer0_outputs(8998) <= (inputs(132)) xor (inputs(50));
    layer0_outputs(8999) <= not(inputs(88));
    layer0_outputs(9000) <= inputs(175);
    layer0_outputs(9001) <= not((inputs(3)) or (inputs(158)));
    layer0_outputs(9002) <= not((inputs(7)) or (inputs(99)));
    layer0_outputs(9003) <= (inputs(52)) and not (inputs(223));
    layer0_outputs(9004) <= not(inputs(36)) or (inputs(150));
    layer0_outputs(9005) <= inputs(23);
    layer0_outputs(9006) <= (inputs(68)) or (inputs(146));
    layer0_outputs(9007) <= (inputs(99)) xor (inputs(113));
    layer0_outputs(9008) <= inputs(136);
    layer0_outputs(9009) <= (inputs(33)) or (inputs(100));
    layer0_outputs(9010) <= inputs(152);
    layer0_outputs(9011) <= (inputs(96)) xor (inputs(107));
    layer0_outputs(9012) <= not(inputs(183));
    layer0_outputs(9013) <= inputs(127);
    layer0_outputs(9014) <= not(inputs(60));
    layer0_outputs(9015) <= inputs(229);
    layer0_outputs(9016) <= (inputs(186)) xor (inputs(54));
    layer0_outputs(9017) <= (inputs(167)) and not (inputs(102));
    layer0_outputs(9018) <= not(inputs(12)) or (inputs(114));
    layer0_outputs(9019) <= not((inputs(255)) or (inputs(250)));
    layer0_outputs(9020) <= (inputs(196)) and not (inputs(12));
    layer0_outputs(9021) <= (inputs(160)) xor (inputs(164));
    layer0_outputs(9022) <= (inputs(146)) or (inputs(22));
    layer0_outputs(9023) <= inputs(51);
    layer0_outputs(9024) <= not(inputs(18));
    layer0_outputs(9025) <= not((inputs(55)) xor (inputs(53)));
    layer0_outputs(9026) <= not((inputs(8)) xor (inputs(115)));
    layer0_outputs(9027) <= not((inputs(202)) or (inputs(18)));
    layer0_outputs(9028) <= not((inputs(134)) and (inputs(90)));
    layer0_outputs(9029) <= not((inputs(192)) or (inputs(194)));
    layer0_outputs(9030) <= (inputs(143)) or (inputs(172));
    layer0_outputs(9031) <= (inputs(22)) and not (inputs(50));
    layer0_outputs(9032) <= (inputs(233)) or (inputs(224));
    layer0_outputs(9033) <= inputs(40);
    layer0_outputs(9034) <= not((inputs(62)) or (inputs(98)));
    layer0_outputs(9035) <= not((inputs(254)) or (inputs(174)));
    layer0_outputs(9036) <= not(inputs(198));
    layer0_outputs(9037) <= inputs(245);
    layer0_outputs(9038) <= (inputs(30)) and not (inputs(3));
    layer0_outputs(9039) <= not(inputs(106));
    layer0_outputs(9040) <= not(inputs(204));
    layer0_outputs(9041) <= '0';
    layer0_outputs(9042) <= (inputs(127)) and not (inputs(141));
    layer0_outputs(9043) <= (inputs(161)) xor (inputs(165));
    layer0_outputs(9044) <= inputs(3);
    layer0_outputs(9045) <= (inputs(209)) or (inputs(244));
    layer0_outputs(9046) <= (inputs(69)) and not (inputs(250));
    layer0_outputs(9047) <= not(inputs(23)) or (inputs(249));
    layer0_outputs(9048) <= inputs(228);
    layer0_outputs(9049) <= inputs(198);
    layer0_outputs(9050) <= not(inputs(142)) or (inputs(235));
    layer0_outputs(9051) <= inputs(125);
    layer0_outputs(9052) <= not((inputs(2)) or (inputs(40)));
    layer0_outputs(9053) <= not((inputs(36)) xor (inputs(192)));
    layer0_outputs(9054) <= not((inputs(89)) xor (inputs(63)));
    layer0_outputs(9055) <= (inputs(242)) or (inputs(72));
    layer0_outputs(9056) <= not((inputs(141)) and (inputs(148)));
    layer0_outputs(9057) <= not((inputs(10)) xor (inputs(253)));
    layer0_outputs(9058) <= inputs(202);
    layer0_outputs(9059) <= not(inputs(39));
    layer0_outputs(9060) <= not(inputs(134));
    layer0_outputs(9061) <= not(inputs(83)) or (inputs(175));
    layer0_outputs(9062) <= '1';
    layer0_outputs(9063) <= not(inputs(151)) or (inputs(92));
    layer0_outputs(9064) <= inputs(164);
    layer0_outputs(9065) <= not(inputs(11)) or (inputs(251));
    layer0_outputs(9066) <= not((inputs(224)) or (inputs(56)));
    layer0_outputs(9067) <= not(inputs(82)) or (inputs(2));
    layer0_outputs(9068) <= not((inputs(186)) or (inputs(96)));
    layer0_outputs(9069) <= inputs(164);
    layer0_outputs(9070) <= not((inputs(32)) xor (inputs(100)));
    layer0_outputs(9071) <= inputs(99);
    layer0_outputs(9072) <= (inputs(67)) or (inputs(48));
    layer0_outputs(9073) <= not(inputs(183)) or (inputs(105));
    layer0_outputs(9074) <= (inputs(223)) and (inputs(173));
    layer0_outputs(9075) <= not((inputs(145)) xor (inputs(159)));
    layer0_outputs(9076) <= inputs(81);
    layer0_outputs(9077) <= (inputs(76)) and not (inputs(175));
    layer0_outputs(9078) <= (inputs(140)) and not (inputs(177));
    layer0_outputs(9079) <= not(inputs(41)) or (inputs(255));
    layer0_outputs(9080) <= not((inputs(168)) or (inputs(49)));
    layer0_outputs(9081) <= inputs(28);
    layer0_outputs(9082) <= inputs(118);
    layer0_outputs(9083) <= (inputs(234)) or (inputs(152));
    layer0_outputs(9084) <= not((inputs(174)) xor (inputs(150)));
    layer0_outputs(9085) <= not((inputs(204)) or (inputs(246)));
    layer0_outputs(9086) <= inputs(84);
    layer0_outputs(9087) <= inputs(98);
    layer0_outputs(9088) <= (inputs(150)) and not (inputs(179));
    layer0_outputs(9089) <= not(inputs(165)) or (inputs(141));
    layer0_outputs(9090) <= not(inputs(22));
    layer0_outputs(9091) <= inputs(38);
    layer0_outputs(9092) <= not(inputs(241));
    layer0_outputs(9093) <= not(inputs(23)) or (inputs(240));
    layer0_outputs(9094) <= inputs(13);
    layer0_outputs(9095) <= not(inputs(246)) or (inputs(28));
    layer0_outputs(9096) <= (inputs(154)) xor (inputs(103));
    layer0_outputs(9097) <= not(inputs(142));
    layer0_outputs(9098) <= inputs(166);
    layer0_outputs(9099) <= (inputs(81)) or (inputs(97));
    layer0_outputs(9100) <= (inputs(222)) xor (inputs(94));
    layer0_outputs(9101) <= not(inputs(174));
    layer0_outputs(9102) <= not(inputs(51));
    layer0_outputs(9103) <= inputs(135);
    layer0_outputs(9104) <= not((inputs(241)) xor (inputs(124)));
    layer0_outputs(9105) <= not(inputs(108));
    layer0_outputs(9106) <= not(inputs(204)) or (inputs(7));
    layer0_outputs(9107) <= (inputs(90)) and not (inputs(252));
    layer0_outputs(9108) <= (inputs(228)) and (inputs(248));
    layer0_outputs(9109) <= (inputs(41)) xor (inputs(147));
    layer0_outputs(9110) <= inputs(167);
    layer0_outputs(9111) <= not(inputs(246)) or (inputs(75));
    layer0_outputs(9112) <= inputs(204);
    layer0_outputs(9113) <= not((inputs(254)) and (inputs(146)));
    layer0_outputs(9114) <= inputs(167);
    layer0_outputs(9115) <= (inputs(176)) or (inputs(217));
    layer0_outputs(9116) <= (inputs(131)) or (inputs(46));
    layer0_outputs(9117) <= not(inputs(9));
    layer0_outputs(9118) <= inputs(149);
    layer0_outputs(9119) <= not((inputs(53)) or (inputs(112)));
    layer0_outputs(9120) <= (inputs(252)) and not (inputs(241));
    layer0_outputs(9121) <= (inputs(104)) and not (inputs(162));
    layer0_outputs(9122) <= (inputs(218)) or (inputs(196));
    layer0_outputs(9123) <= inputs(132);
    layer0_outputs(9124) <= (inputs(212)) or (inputs(176));
    layer0_outputs(9125) <= (inputs(154)) or (inputs(114));
    layer0_outputs(9126) <= inputs(166);
    layer0_outputs(9127) <= not((inputs(169)) xor (inputs(167)));
    layer0_outputs(9128) <= (inputs(193)) and not (inputs(155));
    layer0_outputs(9129) <= not(inputs(2)) or (inputs(98));
    layer0_outputs(9130) <= not(inputs(135));
    layer0_outputs(9131) <= not((inputs(252)) or (inputs(250)));
    layer0_outputs(9132) <= not((inputs(81)) or (inputs(249)));
    layer0_outputs(9133) <= (inputs(69)) and not (inputs(214));
    layer0_outputs(9134) <= not(inputs(80));
    layer0_outputs(9135) <= (inputs(71)) and not (inputs(116));
    layer0_outputs(9136) <= inputs(214);
    layer0_outputs(9137) <= (inputs(254)) and not (inputs(72));
    layer0_outputs(9138) <= (inputs(198)) xor (inputs(180));
    layer0_outputs(9139) <= not((inputs(44)) xor (inputs(226)));
    layer0_outputs(9140) <= not(inputs(252)) or (inputs(124));
    layer0_outputs(9141) <= not(inputs(204));
    layer0_outputs(9142) <= (inputs(5)) and not (inputs(47));
    layer0_outputs(9143) <= not((inputs(46)) or (inputs(45)));
    layer0_outputs(9144) <= (inputs(119)) and not (inputs(221));
    layer0_outputs(9145) <= inputs(61);
    layer0_outputs(9146) <= not((inputs(175)) xor (inputs(217)));
    layer0_outputs(9147) <= not((inputs(139)) or (inputs(33)));
    layer0_outputs(9148) <= not((inputs(228)) or (inputs(212)));
    layer0_outputs(9149) <= '1';
    layer0_outputs(9150) <= inputs(64);
    layer0_outputs(9151) <= (inputs(227)) or (inputs(127));
    layer0_outputs(9152) <= not(inputs(183)) or (inputs(223));
    layer0_outputs(9153) <= inputs(174);
    layer0_outputs(9154) <= not(inputs(219));
    layer0_outputs(9155) <= not(inputs(143));
    layer0_outputs(9156) <= (inputs(126)) or (inputs(153));
    layer0_outputs(9157) <= inputs(43);
    layer0_outputs(9158) <= not(inputs(120));
    layer0_outputs(9159) <= not((inputs(156)) xor (inputs(107)));
    layer0_outputs(9160) <= (inputs(226)) xor (inputs(175));
    layer0_outputs(9161) <= (inputs(14)) or (inputs(247));
    layer0_outputs(9162) <= (inputs(186)) xor (inputs(208));
    layer0_outputs(9163) <= inputs(126);
    layer0_outputs(9164) <= not(inputs(43)) or (inputs(88));
    layer0_outputs(9165) <= (inputs(75)) and (inputs(9));
    layer0_outputs(9166) <= inputs(238);
    layer0_outputs(9167) <= (inputs(60)) and (inputs(87));
    layer0_outputs(9168) <= inputs(9);
    layer0_outputs(9169) <= (inputs(136)) xor (inputs(3));
    layer0_outputs(9170) <= (inputs(73)) xor (inputs(77));
    layer0_outputs(9171) <= (inputs(41)) or (inputs(228));
    layer0_outputs(9172) <= inputs(96);
    layer0_outputs(9173) <= (inputs(187)) and not (inputs(234));
    layer0_outputs(9174) <= not((inputs(94)) or (inputs(91)));
    layer0_outputs(9175) <= not(inputs(119));
    layer0_outputs(9176) <= not((inputs(231)) or (inputs(249)));
    layer0_outputs(9177) <= (inputs(207)) and (inputs(196));
    layer0_outputs(9178) <= not(inputs(40));
    layer0_outputs(9179) <= not((inputs(251)) or (inputs(112)));
    layer0_outputs(9180) <= not((inputs(241)) or (inputs(150)));
    layer0_outputs(9181) <= not(inputs(196)) or (inputs(28));
    layer0_outputs(9182) <= inputs(199);
    layer0_outputs(9183) <= not(inputs(212)) or (inputs(100));
    layer0_outputs(9184) <= not(inputs(84)) or (inputs(16));
    layer0_outputs(9185) <= not(inputs(105)) or (inputs(190));
    layer0_outputs(9186) <= '0';
    layer0_outputs(9187) <= not(inputs(26)) or (inputs(15));
    layer0_outputs(9188) <= (inputs(76)) and not (inputs(102));
    layer0_outputs(9189) <= not(inputs(189));
    layer0_outputs(9190) <= not(inputs(144));
    layer0_outputs(9191) <= not(inputs(108)) or (inputs(65));
    layer0_outputs(9192) <= not((inputs(65)) xor (inputs(35)));
    layer0_outputs(9193) <= not((inputs(21)) xor (inputs(230)));
    layer0_outputs(9194) <= (inputs(247)) and not (inputs(40));
    layer0_outputs(9195) <= not((inputs(79)) or (inputs(97)));
    layer0_outputs(9196) <= (inputs(123)) or (inputs(43));
    layer0_outputs(9197) <= not((inputs(192)) or (inputs(174)));
    layer0_outputs(9198) <= inputs(134);
    layer0_outputs(9199) <= not((inputs(19)) or (inputs(123)));
    layer0_outputs(9200) <= (inputs(16)) or (inputs(32));
    layer0_outputs(9201) <= inputs(130);
    layer0_outputs(9202) <= not((inputs(51)) or (inputs(150)));
    layer0_outputs(9203) <= (inputs(203)) xor (inputs(238));
    layer0_outputs(9204) <= (inputs(198)) and not (inputs(205));
    layer0_outputs(9205) <= (inputs(99)) xor (inputs(21));
    layer0_outputs(9206) <= (inputs(249)) xor (inputs(48));
    layer0_outputs(9207) <= not(inputs(21));
    layer0_outputs(9208) <= not(inputs(165));
    layer0_outputs(9209) <= not(inputs(119));
    layer0_outputs(9210) <= not((inputs(201)) and (inputs(136)));
    layer0_outputs(9211) <= not((inputs(136)) or (inputs(119)));
    layer0_outputs(9212) <= (inputs(204)) and not (inputs(81));
    layer0_outputs(9213) <= inputs(214);
    layer0_outputs(9214) <= inputs(92);
    layer0_outputs(9215) <= not((inputs(182)) xor (inputs(165)));
    layer0_outputs(9216) <= not((inputs(252)) xor (inputs(77)));
    layer0_outputs(9217) <= not((inputs(61)) xor (inputs(120)));
    layer0_outputs(9218) <= (inputs(19)) xor (inputs(33));
    layer0_outputs(9219) <= (inputs(117)) and (inputs(26));
    layer0_outputs(9220) <= not(inputs(108)) or (inputs(160));
    layer0_outputs(9221) <= not((inputs(55)) xor (inputs(226)));
    layer0_outputs(9222) <= not(inputs(26)) or (inputs(179));
    layer0_outputs(9223) <= not((inputs(78)) xor (inputs(207)));
    layer0_outputs(9224) <= not(inputs(61)) or (inputs(237));
    layer0_outputs(9225) <= (inputs(33)) xor (inputs(11));
    layer0_outputs(9226) <= (inputs(56)) xor (inputs(60));
    layer0_outputs(9227) <= not((inputs(176)) xor (inputs(241)));
    layer0_outputs(9228) <= not(inputs(157)) or (inputs(242));
    layer0_outputs(9229) <= not((inputs(110)) or (inputs(0)));
    layer0_outputs(9230) <= not(inputs(114));
    layer0_outputs(9231) <= inputs(228);
    layer0_outputs(9232) <= (inputs(143)) and (inputs(183));
    layer0_outputs(9233) <= (inputs(197)) and not (inputs(18));
    layer0_outputs(9234) <= not(inputs(202)) or (inputs(109));
    layer0_outputs(9235) <= (inputs(49)) or (inputs(73));
    layer0_outputs(9236) <= not(inputs(170));
    layer0_outputs(9237) <= inputs(122);
    layer0_outputs(9238) <= (inputs(203)) or (inputs(127));
    layer0_outputs(9239) <= (inputs(172)) and not (inputs(71));
    layer0_outputs(9240) <= (inputs(233)) or (inputs(237));
    layer0_outputs(9241) <= inputs(41);
    layer0_outputs(9242) <= not(inputs(150));
    layer0_outputs(9243) <= (inputs(73)) xor (inputs(60));
    layer0_outputs(9244) <= not((inputs(4)) xor (inputs(86)));
    layer0_outputs(9245) <= (inputs(46)) or (inputs(2));
    layer0_outputs(9246) <= (inputs(183)) and not (inputs(45));
    layer0_outputs(9247) <= not(inputs(167)) or (inputs(94));
    layer0_outputs(9248) <= not(inputs(133)) or (inputs(112));
    layer0_outputs(9249) <= not(inputs(119)) or (inputs(76));
    layer0_outputs(9250) <= (inputs(18)) or (inputs(151));
    layer0_outputs(9251) <= not((inputs(29)) or (inputs(108)));
    layer0_outputs(9252) <= not((inputs(43)) or (inputs(241)));
    layer0_outputs(9253) <= not((inputs(37)) or (inputs(163)));
    layer0_outputs(9254) <= inputs(106);
    layer0_outputs(9255) <= inputs(11);
    layer0_outputs(9256) <= not((inputs(160)) or (inputs(116)));
    layer0_outputs(9257) <= not(inputs(217));
    layer0_outputs(9258) <= not(inputs(169)) or (inputs(149));
    layer0_outputs(9259) <= (inputs(60)) xor (inputs(4));
    layer0_outputs(9260) <= not((inputs(109)) or (inputs(70)));
    layer0_outputs(9261) <= not((inputs(188)) or (inputs(159)));
    layer0_outputs(9262) <= (inputs(66)) xor (inputs(42));
    layer0_outputs(9263) <= inputs(152);
    layer0_outputs(9264) <= not(inputs(106)) or (inputs(23));
    layer0_outputs(9265) <= (inputs(114)) and (inputs(67));
    layer0_outputs(9266) <= inputs(151);
    layer0_outputs(9267) <= inputs(67);
    layer0_outputs(9268) <= (inputs(161)) or (inputs(174));
    layer0_outputs(9269) <= (inputs(97)) and (inputs(104));
    layer0_outputs(9270) <= inputs(7);
    layer0_outputs(9271) <= '1';
    layer0_outputs(9272) <= not((inputs(175)) or (inputs(203)));
    layer0_outputs(9273) <= not((inputs(117)) or (inputs(251)));
    layer0_outputs(9274) <= (inputs(55)) or (inputs(6));
    layer0_outputs(9275) <= inputs(95);
    layer0_outputs(9276) <= (inputs(157)) or (inputs(143));
    layer0_outputs(9277) <= not(inputs(183)) or (inputs(41));
    layer0_outputs(9278) <= (inputs(83)) xor (inputs(53));
    layer0_outputs(9279) <= (inputs(74)) xor (inputs(165));
    layer0_outputs(9280) <= (inputs(161)) and not (inputs(46));
    layer0_outputs(9281) <= (inputs(69)) and (inputs(40));
    layer0_outputs(9282) <= (inputs(48)) or (inputs(229));
    layer0_outputs(9283) <= not((inputs(250)) or (inputs(226)));
    layer0_outputs(9284) <= not((inputs(76)) and (inputs(39)));
    layer0_outputs(9285) <= not((inputs(150)) or (inputs(190)));
    layer0_outputs(9286) <= not((inputs(170)) or (inputs(84)));
    layer0_outputs(9287) <= not(inputs(251));
    layer0_outputs(9288) <= not(inputs(208));
    layer0_outputs(9289) <= not((inputs(195)) or (inputs(35)));
    layer0_outputs(9290) <= not((inputs(104)) or (inputs(165)));
    layer0_outputs(9291) <= (inputs(190)) and not (inputs(231));
    layer0_outputs(9292) <= not(inputs(114));
    layer0_outputs(9293) <= not((inputs(57)) or (inputs(228)));
    layer0_outputs(9294) <= (inputs(13)) or (inputs(29));
    layer0_outputs(9295) <= not(inputs(90)) or (inputs(14));
    layer0_outputs(9296) <= not((inputs(171)) or (inputs(88)));
    layer0_outputs(9297) <= (inputs(72)) xor (inputs(29));
    layer0_outputs(9298) <= not(inputs(220));
    layer0_outputs(9299) <= not((inputs(5)) xor (inputs(57)));
    layer0_outputs(9300) <= not(inputs(102));
    layer0_outputs(9301) <= (inputs(188)) or (inputs(193));
    layer0_outputs(9302) <= not(inputs(23));
    layer0_outputs(9303) <= not((inputs(24)) xor (inputs(75)));
    layer0_outputs(9304) <= not(inputs(27));
    layer0_outputs(9305) <= not(inputs(245));
    layer0_outputs(9306) <= (inputs(129)) xor (inputs(169));
    layer0_outputs(9307) <= not(inputs(171)) or (inputs(163));
    layer0_outputs(9308) <= (inputs(180)) and not (inputs(15));
    layer0_outputs(9309) <= (inputs(146)) and not (inputs(190));
    layer0_outputs(9310) <= '1';
    layer0_outputs(9311) <= not((inputs(63)) xor (inputs(40)));
    layer0_outputs(9312) <= not((inputs(234)) xor (inputs(87)));
    layer0_outputs(9313) <= inputs(199);
    layer0_outputs(9314) <= not(inputs(76));
    layer0_outputs(9315) <= (inputs(64)) and not (inputs(144));
    layer0_outputs(9316) <= inputs(181);
    layer0_outputs(9317) <= '1';
    layer0_outputs(9318) <= inputs(97);
    layer0_outputs(9319) <= inputs(43);
    layer0_outputs(9320) <= not((inputs(98)) or (inputs(117)));
    layer0_outputs(9321) <= (inputs(242)) or (inputs(73));
    layer0_outputs(9322) <= (inputs(172)) or (inputs(159));
    layer0_outputs(9323) <= (inputs(27)) and (inputs(23));
    layer0_outputs(9324) <= not(inputs(245));
    layer0_outputs(9325) <= not((inputs(158)) or (inputs(239)));
    layer0_outputs(9326) <= not(inputs(93));
    layer0_outputs(9327) <= not((inputs(99)) or (inputs(65)));
    layer0_outputs(9328) <= (inputs(99)) or (inputs(199));
    layer0_outputs(9329) <= not(inputs(56));
    layer0_outputs(9330) <= not((inputs(62)) xor (inputs(237)));
    layer0_outputs(9331) <= (inputs(235)) or (inputs(221));
    layer0_outputs(9332) <= not(inputs(124)) or (inputs(255));
    layer0_outputs(9333) <= not(inputs(148));
    layer0_outputs(9334) <= (inputs(185)) and not (inputs(32));
    layer0_outputs(9335) <= not(inputs(107)) or (inputs(179));
    layer0_outputs(9336) <= (inputs(86)) and not (inputs(7));
    layer0_outputs(9337) <= (inputs(244)) and not (inputs(36));
    layer0_outputs(9338) <= not(inputs(151));
    layer0_outputs(9339) <= (inputs(108)) xor (inputs(65));
    layer0_outputs(9340) <= (inputs(231)) xor (inputs(169));
    layer0_outputs(9341) <= (inputs(164)) xor (inputs(167));
    layer0_outputs(9342) <= (inputs(38)) or (inputs(79));
    layer0_outputs(9343) <= not(inputs(12));
    layer0_outputs(9344) <= not(inputs(198));
    layer0_outputs(9345) <= (inputs(188)) and (inputs(219));
    layer0_outputs(9346) <= not(inputs(8));
    layer0_outputs(9347) <= not(inputs(230));
    layer0_outputs(9348) <= not(inputs(156)) or (inputs(109));
    layer0_outputs(9349) <= not((inputs(172)) xor (inputs(80)));
    layer0_outputs(9350) <= not((inputs(5)) or (inputs(8)));
    layer0_outputs(9351) <= not(inputs(230));
    layer0_outputs(9352) <= not(inputs(246)) or (inputs(72));
    layer0_outputs(9353) <= (inputs(30)) and not (inputs(130));
    layer0_outputs(9354) <= not(inputs(142));
    layer0_outputs(9355) <= not(inputs(168));
    layer0_outputs(9356) <= not((inputs(82)) xor (inputs(78)));
    layer0_outputs(9357) <= not(inputs(103));
    layer0_outputs(9358) <= (inputs(152)) and not (inputs(234));
    layer0_outputs(9359) <= '0';
    layer0_outputs(9360) <= not(inputs(186)) or (inputs(14));
    layer0_outputs(9361) <= not(inputs(122)) or (inputs(131));
    layer0_outputs(9362) <= not(inputs(13)) or (inputs(224));
    layer0_outputs(9363) <= not((inputs(62)) or (inputs(205)));
    layer0_outputs(9364) <= not(inputs(121));
    layer0_outputs(9365) <= (inputs(149)) or (inputs(150));
    layer0_outputs(9366) <= inputs(142);
    layer0_outputs(9367) <= (inputs(232)) or (inputs(114));
    layer0_outputs(9368) <= (inputs(134)) or (inputs(219));
    layer0_outputs(9369) <= (inputs(86)) and not (inputs(72));
    layer0_outputs(9370) <= not((inputs(111)) xor (inputs(221)));
    layer0_outputs(9371) <= not((inputs(206)) or (inputs(95)));
    layer0_outputs(9372) <= not((inputs(239)) or (inputs(142)));
    layer0_outputs(9373) <= (inputs(144)) and not (inputs(49));
    layer0_outputs(9374) <= '0';
    layer0_outputs(9375) <= not((inputs(40)) or (inputs(34)));
    layer0_outputs(9376) <= not((inputs(179)) or (inputs(238)));
    layer0_outputs(9377) <= not((inputs(153)) or (inputs(71)));
    layer0_outputs(9378) <= not(inputs(22));
    layer0_outputs(9379) <= inputs(62);
    layer0_outputs(9380) <= (inputs(33)) or (inputs(19));
    layer0_outputs(9381) <= inputs(162);
    layer0_outputs(9382) <= (inputs(40)) xor (inputs(18));
    layer0_outputs(9383) <= inputs(127);
    layer0_outputs(9384) <= (inputs(156)) or (inputs(59));
    layer0_outputs(9385) <= not((inputs(23)) or (inputs(54)));
    layer0_outputs(9386) <= inputs(136);
    layer0_outputs(9387) <= not(inputs(27));
    layer0_outputs(9388) <= (inputs(133)) xor (inputs(163));
    layer0_outputs(9389) <= not(inputs(44));
    layer0_outputs(9390) <= inputs(178);
    layer0_outputs(9391) <= not(inputs(135)) or (inputs(8));
    layer0_outputs(9392) <= (inputs(206)) and not (inputs(29));
    layer0_outputs(9393) <= not(inputs(117));
    layer0_outputs(9394) <= not(inputs(154));
    layer0_outputs(9395) <= inputs(234);
    layer0_outputs(9396) <= not((inputs(163)) or (inputs(141)));
    layer0_outputs(9397) <= not(inputs(9));
    layer0_outputs(9398) <= not(inputs(9));
    layer0_outputs(9399) <= (inputs(155)) or (inputs(62));
    layer0_outputs(9400) <= (inputs(24)) xor (inputs(193));
    layer0_outputs(9401) <= not(inputs(85));
    layer0_outputs(9402) <= inputs(242);
    layer0_outputs(9403) <= (inputs(181)) and not (inputs(243));
    layer0_outputs(9404) <= not(inputs(48));
    layer0_outputs(9405) <= not((inputs(96)) or (inputs(218)));
    layer0_outputs(9406) <= not((inputs(8)) xor (inputs(9)));
    layer0_outputs(9407) <= inputs(91);
    layer0_outputs(9408) <= not((inputs(179)) or (inputs(62)));
    layer0_outputs(9409) <= inputs(82);
    layer0_outputs(9410) <= inputs(237);
    layer0_outputs(9411) <= not(inputs(247));
    layer0_outputs(9412) <= not((inputs(41)) or (inputs(125)));
    layer0_outputs(9413) <= not(inputs(133)) or (inputs(77));
    layer0_outputs(9414) <= not(inputs(134));
    layer0_outputs(9415) <= (inputs(203)) or (inputs(2));
    layer0_outputs(9416) <= not((inputs(217)) xor (inputs(77)));
    layer0_outputs(9417) <= (inputs(253)) or (inputs(129));
    layer0_outputs(9418) <= not(inputs(92)) or (inputs(34));
    layer0_outputs(9419) <= not(inputs(188)) or (inputs(77));
    layer0_outputs(9420) <= not((inputs(188)) or (inputs(215)));
    layer0_outputs(9421) <= not((inputs(17)) or (inputs(217)));
    layer0_outputs(9422) <= (inputs(56)) and not (inputs(134));
    layer0_outputs(9423) <= not(inputs(218));
    layer0_outputs(9424) <= not((inputs(127)) or (inputs(177)));
    layer0_outputs(9425) <= inputs(65);
    layer0_outputs(9426) <= not((inputs(115)) or (inputs(158)));
    layer0_outputs(9427) <= (inputs(154)) xor (inputs(7));
    layer0_outputs(9428) <= not((inputs(44)) xor (inputs(159)));
    layer0_outputs(9429) <= not((inputs(163)) and (inputs(60)));
    layer0_outputs(9430) <= (inputs(29)) or (inputs(143));
    layer0_outputs(9431) <= inputs(165);
    layer0_outputs(9432) <= not((inputs(156)) xor (inputs(122)));
    layer0_outputs(9433) <= not((inputs(112)) and (inputs(2)));
    layer0_outputs(9434) <= not(inputs(73));
    layer0_outputs(9435) <= inputs(129);
    layer0_outputs(9436) <= not(inputs(248)) or (inputs(239));
    layer0_outputs(9437) <= inputs(97);
    layer0_outputs(9438) <= inputs(70);
    layer0_outputs(9439) <= not((inputs(31)) xor (inputs(172)));
    layer0_outputs(9440) <= not((inputs(221)) or (inputs(60)));
    layer0_outputs(9441) <= (inputs(51)) and not (inputs(113));
    layer0_outputs(9442) <= not((inputs(89)) xor (inputs(126)));
    layer0_outputs(9443) <= not(inputs(107));
    layer0_outputs(9444) <= not((inputs(186)) or (inputs(205)));
    layer0_outputs(9445) <= not((inputs(249)) xor (inputs(178)));
    layer0_outputs(9446) <= (inputs(58)) and not (inputs(110));
    layer0_outputs(9447) <= not(inputs(70)) or (inputs(157));
    layer0_outputs(9448) <= not(inputs(45)) or (inputs(136));
    layer0_outputs(9449) <= inputs(220);
    layer0_outputs(9450) <= not(inputs(116)) or (inputs(224));
    layer0_outputs(9451) <= (inputs(73)) and not (inputs(37));
    layer0_outputs(9452) <= inputs(114);
    layer0_outputs(9453) <= not(inputs(101));
    layer0_outputs(9454) <= not(inputs(59));
    layer0_outputs(9455) <= inputs(179);
    layer0_outputs(9456) <= (inputs(166)) and not (inputs(224));
    layer0_outputs(9457) <= (inputs(123)) and not (inputs(38));
    layer0_outputs(9458) <= (inputs(37)) or (inputs(79));
    layer0_outputs(9459) <= not(inputs(230));
    layer0_outputs(9460) <= inputs(118);
    layer0_outputs(9461) <= not(inputs(158));
    layer0_outputs(9462) <= inputs(193);
    layer0_outputs(9463) <= inputs(82);
    layer0_outputs(9464) <= not(inputs(92));
    layer0_outputs(9465) <= not(inputs(183)) or (inputs(32));
    layer0_outputs(9466) <= not(inputs(20));
    layer0_outputs(9467) <= not(inputs(228));
    layer0_outputs(9468) <= (inputs(231)) or (inputs(210));
    layer0_outputs(9469) <= not(inputs(132));
    layer0_outputs(9470) <= (inputs(220)) xor (inputs(115));
    layer0_outputs(9471) <= (inputs(104)) and not (inputs(238));
    layer0_outputs(9472) <= not((inputs(15)) and (inputs(224)));
    layer0_outputs(9473) <= not(inputs(136)) or (inputs(20));
    layer0_outputs(9474) <= not((inputs(136)) or (inputs(49)));
    layer0_outputs(9475) <= not(inputs(68));
    layer0_outputs(9476) <= not(inputs(99));
    layer0_outputs(9477) <= (inputs(87)) and not (inputs(96));
    layer0_outputs(9478) <= not((inputs(199)) xor (inputs(223)));
    layer0_outputs(9479) <= not(inputs(14));
    layer0_outputs(9480) <= (inputs(111)) and not (inputs(55));
    layer0_outputs(9481) <= inputs(54);
    layer0_outputs(9482) <= not(inputs(98));
    layer0_outputs(9483) <= (inputs(20)) xor (inputs(41));
    layer0_outputs(9484) <= (inputs(57)) or (inputs(239));
    layer0_outputs(9485) <= (inputs(86)) or (inputs(81));
    layer0_outputs(9486) <= (inputs(109)) and (inputs(13));
    layer0_outputs(9487) <= not(inputs(105)) or (inputs(176));
    layer0_outputs(9488) <= not(inputs(175));
    layer0_outputs(9489) <= not((inputs(223)) xor (inputs(43)));
    layer0_outputs(9490) <= not((inputs(148)) or (inputs(202)));
    layer0_outputs(9491) <= (inputs(95)) or (inputs(49));
    layer0_outputs(9492) <= (inputs(6)) xor (inputs(211));
    layer0_outputs(9493) <= not((inputs(15)) or (inputs(172)));
    layer0_outputs(9494) <= not((inputs(173)) xor (inputs(214)));
    layer0_outputs(9495) <= (inputs(249)) and not (inputs(142));
    layer0_outputs(9496) <= (inputs(169)) and not (inputs(45));
    layer0_outputs(9497) <= (inputs(56)) and not (inputs(140));
    layer0_outputs(9498) <= not((inputs(220)) or (inputs(203)));
    layer0_outputs(9499) <= (inputs(148)) xor (inputs(187));
    layer0_outputs(9500) <= (inputs(66)) or (inputs(69));
    layer0_outputs(9501) <= inputs(130);
    layer0_outputs(9502) <= inputs(178);
    layer0_outputs(9503) <= (inputs(189)) xor (inputs(29));
    layer0_outputs(9504) <= not((inputs(179)) xor (inputs(119)));
    layer0_outputs(9505) <= not(inputs(41));
    layer0_outputs(9506) <= '1';
    layer0_outputs(9507) <= not(inputs(106));
    layer0_outputs(9508) <= (inputs(120)) and not (inputs(176));
    layer0_outputs(9509) <= not(inputs(50)) or (inputs(113));
    layer0_outputs(9510) <= not((inputs(100)) xor (inputs(227)));
    layer0_outputs(9511) <= not((inputs(98)) or (inputs(165)));
    layer0_outputs(9512) <= (inputs(136)) and not (inputs(235));
    layer0_outputs(9513) <= (inputs(250)) or (inputs(213));
    layer0_outputs(9514) <= not((inputs(161)) xor (inputs(175)));
    layer0_outputs(9515) <= not(inputs(41));
    layer0_outputs(9516) <= (inputs(189)) and not (inputs(31));
    layer0_outputs(9517) <= not(inputs(11));
    layer0_outputs(9518) <= (inputs(197)) and not (inputs(93));
    layer0_outputs(9519) <= (inputs(20)) xor (inputs(66));
    layer0_outputs(9520) <= not((inputs(29)) or (inputs(47)));
    layer0_outputs(9521) <= (inputs(170)) and (inputs(188));
    layer0_outputs(9522) <= inputs(92);
    layer0_outputs(9523) <= inputs(40);
    layer0_outputs(9524) <= (inputs(142)) and not (inputs(31));
    layer0_outputs(9525) <= not((inputs(53)) and (inputs(59)));
    layer0_outputs(9526) <= not((inputs(184)) or (inputs(176)));
    layer0_outputs(9527) <= not((inputs(25)) or (inputs(78)));
    layer0_outputs(9528) <= (inputs(194)) and not (inputs(176));
    layer0_outputs(9529) <= inputs(36);
    layer0_outputs(9530) <= not((inputs(32)) or (inputs(179)));
    layer0_outputs(9531) <= inputs(231);
    layer0_outputs(9532) <= inputs(110);
    layer0_outputs(9533) <= (inputs(128)) and not (inputs(30));
    layer0_outputs(9534) <= inputs(156);
    layer0_outputs(9535) <= not((inputs(246)) xor (inputs(188)));
    layer0_outputs(9536) <= not((inputs(86)) or (inputs(195)));
    layer0_outputs(9537) <= not(inputs(63));
    layer0_outputs(9538) <= (inputs(34)) or (inputs(244));
    layer0_outputs(9539) <= not(inputs(161)) or (inputs(134));
    layer0_outputs(9540) <= not((inputs(219)) or (inputs(178)));
    layer0_outputs(9541) <= not((inputs(225)) or (inputs(6)));
    layer0_outputs(9542) <= inputs(147);
    layer0_outputs(9543) <= (inputs(231)) or (inputs(229));
    layer0_outputs(9544) <= inputs(92);
    layer0_outputs(9545) <= inputs(0);
    layer0_outputs(9546) <= not((inputs(16)) xor (inputs(64)));
    layer0_outputs(9547) <= (inputs(40)) xor (inputs(112));
    layer0_outputs(9548) <= not(inputs(100)) or (inputs(80));
    layer0_outputs(9549) <= (inputs(149)) and not (inputs(174));
    layer0_outputs(9550) <= (inputs(242)) xor (inputs(170));
    layer0_outputs(9551) <= not((inputs(124)) or (inputs(167)));
    layer0_outputs(9552) <= not((inputs(43)) xor (inputs(153)));
    layer0_outputs(9553) <= inputs(114);
    layer0_outputs(9554) <= not((inputs(210)) and (inputs(61)));
    layer0_outputs(9555) <= (inputs(46)) and not (inputs(11));
    layer0_outputs(9556) <= (inputs(195)) or (inputs(94));
    layer0_outputs(9557) <= not(inputs(148));
    layer0_outputs(9558) <= inputs(198);
    layer0_outputs(9559) <= not((inputs(17)) or (inputs(253)));
    layer0_outputs(9560) <= inputs(88);
    layer0_outputs(9561) <= not((inputs(80)) xor (inputs(50)));
    layer0_outputs(9562) <= not(inputs(102)) or (inputs(81));
    layer0_outputs(9563) <= not(inputs(53));
    layer0_outputs(9564) <= (inputs(42)) or (inputs(66));
    layer0_outputs(9565) <= inputs(239);
    layer0_outputs(9566) <= (inputs(80)) xor (inputs(20));
    layer0_outputs(9567) <= not((inputs(204)) xor (inputs(152)));
    layer0_outputs(9568) <= (inputs(167)) and not (inputs(72));
    layer0_outputs(9569) <= (inputs(22)) xor (inputs(95));
    layer0_outputs(9570) <= not(inputs(229)) or (inputs(15));
    layer0_outputs(9571) <= not((inputs(207)) or (inputs(67)));
    layer0_outputs(9572) <= not(inputs(60)) or (inputs(254));
    layer0_outputs(9573) <= inputs(68);
    layer0_outputs(9574) <= inputs(18);
    layer0_outputs(9575) <= (inputs(184)) or (inputs(14));
    layer0_outputs(9576) <= not(inputs(45));
    layer0_outputs(9577) <= (inputs(193)) or (inputs(198));
    layer0_outputs(9578) <= '0';
    layer0_outputs(9579) <= not(inputs(133));
    layer0_outputs(9580) <= '0';
    layer0_outputs(9581) <= not(inputs(69)) or (inputs(63));
    layer0_outputs(9582) <= not(inputs(81));
    layer0_outputs(9583) <= not(inputs(85)) or (inputs(215));
    layer0_outputs(9584) <= inputs(173);
    layer0_outputs(9585) <= (inputs(75)) and not (inputs(23));
    layer0_outputs(9586) <= not((inputs(88)) or (inputs(151)));
    layer0_outputs(9587) <= (inputs(100)) or (inputs(61));
    layer0_outputs(9588) <= not(inputs(53));
    layer0_outputs(9589) <= (inputs(251)) and not (inputs(241));
    layer0_outputs(9590) <= inputs(149);
    layer0_outputs(9591) <= not(inputs(67));
    layer0_outputs(9592) <= inputs(19);
    layer0_outputs(9593) <= not((inputs(128)) or (inputs(1)));
    layer0_outputs(9594) <= inputs(68);
    layer0_outputs(9595) <= not(inputs(179));
    layer0_outputs(9596) <= not((inputs(29)) xor (inputs(138)));
    layer0_outputs(9597) <= not(inputs(205));
    layer0_outputs(9598) <= not(inputs(181));
    layer0_outputs(9599) <= (inputs(115)) and not (inputs(1));
    layer0_outputs(9600) <= inputs(204);
    layer0_outputs(9601) <= not((inputs(133)) or (inputs(183)));
    layer0_outputs(9602) <= not((inputs(226)) and (inputs(136)));
    layer0_outputs(9603) <= not(inputs(168));
    layer0_outputs(9604) <= (inputs(218)) or (inputs(51));
    layer0_outputs(9605) <= inputs(173);
    layer0_outputs(9606) <= not((inputs(238)) or (inputs(183)));
    layer0_outputs(9607) <= not(inputs(85)) or (inputs(48));
    layer0_outputs(9608) <= not((inputs(122)) xor (inputs(171)));
    layer0_outputs(9609) <= not(inputs(27)) or (inputs(194));
    layer0_outputs(9610) <= (inputs(245)) or (inputs(87));
    layer0_outputs(9611) <= not(inputs(178)) or (inputs(239));
    layer0_outputs(9612) <= (inputs(216)) or (inputs(207));
    layer0_outputs(9613) <= not(inputs(245));
    layer0_outputs(9614) <= (inputs(241)) and not (inputs(234));
    layer0_outputs(9615) <= not((inputs(92)) or (inputs(39)));
    layer0_outputs(9616) <= not((inputs(179)) xor (inputs(126)));
    layer0_outputs(9617) <= not((inputs(33)) or (inputs(119)));
    layer0_outputs(9618) <= (inputs(218)) or (inputs(207));
    layer0_outputs(9619) <= (inputs(200)) xor (inputs(213));
    layer0_outputs(9620) <= not((inputs(22)) xor (inputs(162)));
    layer0_outputs(9621) <= (inputs(189)) or (inputs(63));
    layer0_outputs(9622) <= not(inputs(199));
    layer0_outputs(9623) <= not(inputs(216));
    layer0_outputs(9624) <= '0';
    layer0_outputs(9625) <= not(inputs(216));
    layer0_outputs(9626) <= not(inputs(100));
    layer0_outputs(9627) <= (inputs(164)) or (inputs(244));
    layer0_outputs(9628) <= inputs(147);
    layer0_outputs(9629) <= (inputs(44)) and not (inputs(115));
    layer0_outputs(9630) <= (inputs(38)) and not (inputs(153));
    layer0_outputs(9631) <= not((inputs(245)) xor (inputs(236)));
    layer0_outputs(9632) <= not(inputs(193));
    layer0_outputs(9633) <= not(inputs(73)) or (inputs(3));
    layer0_outputs(9634) <= not(inputs(109));
    layer0_outputs(9635) <= (inputs(155)) or (inputs(160));
    layer0_outputs(9636) <= not((inputs(185)) or (inputs(6)));
    layer0_outputs(9637) <= not((inputs(217)) xor (inputs(16)));
    layer0_outputs(9638) <= (inputs(35)) and not (inputs(108));
    layer0_outputs(9639) <= (inputs(66)) or (inputs(255));
    layer0_outputs(9640) <= not(inputs(5));
    layer0_outputs(9641) <= not(inputs(147));
    layer0_outputs(9642) <= inputs(236);
    layer0_outputs(9643) <= inputs(40);
    layer0_outputs(9644) <= (inputs(51)) and not (inputs(160));
    layer0_outputs(9645) <= inputs(183);
    layer0_outputs(9646) <= (inputs(1)) or (inputs(152));
    layer0_outputs(9647) <= inputs(120);
    layer0_outputs(9648) <= not(inputs(185)) or (inputs(69));
    layer0_outputs(9649) <= not(inputs(135)) or (inputs(237));
    layer0_outputs(9650) <= inputs(142);
    layer0_outputs(9651) <= (inputs(75)) and not (inputs(191));
    layer0_outputs(9652) <= not((inputs(31)) xor (inputs(248)));
    layer0_outputs(9653) <= inputs(114);
    layer0_outputs(9654) <= not(inputs(127));
    layer0_outputs(9655) <= not((inputs(239)) xor (inputs(182)));
    layer0_outputs(9656) <= inputs(22);
    layer0_outputs(9657) <= inputs(230);
    layer0_outputs(9658) <= not(inputs(86));
    layer0_outputs(9659) <= inputs(81);
    layer0_outputs(9660) <= not(inputs(185)) or (inputs(106));
    layer0_outputs(9661) <= not(inputs(117));
    layer0_outputs(9662) <= not(inputs(183)) or (inputs(134));
    layer0_outputs(9663) <= (inputs(125)) xor (inputs(137));
    layer0_outputs(9664) <= (inputs(129)) or (inputs(183));
    layer0_outputs(9665) <= not(inputs(148)) or (inputs(9));
    layer0_outputs(9666) <= not(inputs(213));
    layer0_outputs(9667) <= not((inputs(124)) or (inputs(110)));
    layer0_outputs(9668) <= not((inputs(92)) or (inputs(215)));
    layer0_outputs(9669) <= not(inputs(80));
    layer0_outputs(9670) <= (inputs(84)) and not (inputs(126));
    layer0_outputs(9671) <= inputs(117);
    layer0_outputs(9672) <= (inputs(193)) and not (inputs(219));
    layer0_outputs(9673) <= (inputs(22)) and not (inputs(30));
    layer0_outputs(9674) <= not((inputs(188)) xor (inputs(84)));
    layer0_outputs(9675) <= not((inputs(66)) or (inputs(126)));
    layer0_outputs(9676) <= (inputs(191)) xor (inputs(208));
    layer0_outputs(9677) <= inputs(103);
    layer0_outputs(9678) <= inputs(181);
    layer0_outputs(9679) <= (inputs(61)) and not (inputs(196));
    layer0_outputs(9680) <= not(inputs(78)) or (inputs(211));
    layer0_outputs(9681) <= not(inputs(248)) or (inputs(183));
    layer0_outputs(9682) <= not((inputs(84)) or (inputs(97)));
    layer0_outputs(9683) <= not((inputs(119)) xor (inputs(82)));
    layer0_outputs(9684) <= inputs(116);
    layer0_outputs(9685) <= (inputs(147)) and (inputs(44));
    layer0_outputs(9686) <= not((inputs(139)) xor (inputs(142)));
    layer0_outputs(9687) <= not((inputs(188)) xor (inputs(95)));
    layer0_outputs(9688) <= (inputs(11)) and not (inputs(34));
    layer0_outputs(9689) <= not(inputs(133)) or (inputs(17));
    layer0_outputs(9690) <= (inputs(33)) and not (inputs(82));
    layer0_outputs(9691) <= (inputs(124)) or (inputs(232));
    layer0_outputs(9692) <= inputs(126);
    layer0_outputs(9693) <= (inputs(134)) xor (inputs(103));
    layer0_outputs(9694) <= inputs(39);
    layer0_outputs(9695) <= (inputs(81)) xor (inputs(170));
    layer0_outputs(9696) <= (inputs(139)) and (inputs(72));
    layer0_outputs(9697) <= (inputs(129)) xor (inputs(148));
    layer0_outputs(9698) <= (inputs(188)) and not (inputs(242));
    layer0_outputs(9699) <= (inputs(243)) xor (inputs(64));
    layer0_outputs(9700) <= inputs(136);
    layer0_outputs(9701) <= not((inputs(82)) or (inputs(111)));
    layer0_outputs(9702) <= not((inputs(198)) and (inputs(219)));
    layer0_outputs(9703) <= (inputs(138)) and not (inputs(56));
    layer0_outputs(9704) <= not((inputs(176)) and (inputs(245)));
    layer0_outputs(9705) <= (inputs(84)) xor (inputs(60));
    layer0_outputs(9706) <= inputs(104);
    layer0_outputs(9707) <= not((inputs(13)) or (inputs(82)));
    layer0_outputs(9708) <= not((inputs(194)) or (inputs(234)));
    layer0_outputs(9709) <= (inputs(201)) and not (inputs(11));
    layer0_outputs(9710) <= (inputs(145)) or (inputs(52));
    layer0_outputs(9711) <= (inputs(199)) and not (inputs(151));
    layer0_outputs(9712) <= not((inputs(5)) xor (inputs(49)));
    layer0_outputs(9713) <= not((inputs(160)) or (inputs(231)));
    layer0_outputs(9714) <= not((inputs(120)) xor (inputs(10)));
    layer0_outputs(9715) <= (inputs(115)) and not (inputs(191));
    layer0_outputs(9716) <= not((inputs(24)) xor (inputs(58)));
    layer0_outputs(9717) <= inputs(111);
    layer0_outputs(9718) <= '0';
    layer0_outputs(9719) <= (inputs(75)) and not (inputs(219));
    layer0_outputs(9720) <= inputs(216);
    layer0_outputs(9721) <= (inputs(151)) and not (inputs(212));
    layer0_outputs(9722) <= (inputs(249)) xor (inputs(217));
    layer0_outputs(9723) <= not(inputs(81));
    layer0_outputs(9724) <= '1';
    layer0_outputs(9725) <= (inputs(146)) xor (inputs(117));
    layer0_outputs(9726) <= not((inputs(90)) or (inputs(218)));
    layer0_outputs(9727) <= (inputs(218)) and not (inputs(115));
    layer0_outputs(9728) <= (inputs(143)) and not (inputs(127));
    layer0_outputs(9729) <= (inputs(133)) and not (inputs(16));
    layer0_outputs(9730) <= not((inputs(244)) or (inputs(193)));
    layer0_outputs(9731) <= not((inputs(69)) xor (inputs(202)));
    layer0_outputs(9732) <= (inputs(196)) and not (inputs(33));
    layer0_outputs(9733) <= not(inputs(113));
    layer0_outputs(9734) <= not(inputs(14));
    layer0_outputs(9735) <= (inputs(146)) and (inputs(114));
    layer0_outputs(9736) <= not(inputs(43)) or (inputs(243));
    layer0_outputs(9737) <= not((inputs(215)) xor (inputs(248)));
    layer0_outputs(9738) <= (inputs(66)) xor (inputs(79));
    layer0_outputs(9739) <= (inputs(113)) and not (inputs(62));
    layer0_outputs(9740) <= not(inputs(162));
    layer0_outputs(9741) <= (inputs(160)) or (inputs(41));
    layer0_outputs(9742) <= inputs(175);
    layer0_outputs(9743) <= (inputs(21)) and not (inputs(175));
    layer0_outputs(9744) <= (inputs(85)) xor (inputs(51));
    layer0_outputs(9745) <= not((inputs(205)) and (inputs(60)));
    layer0_outputs(9746) <= inputs(180);
    layer0_outputs(9747) <= (inputs(14)) and not (inputs(207));
    layer0_outputs(9748) <= not(inputs(77));
    layer0_outputs(9749) <= not((inputs(31)) or (inputs(108)));
    layer0_outputs(9750) <= (inputs(123)) or (inputs(53));
    layer0_outputs(9751) <= not(inputs(24));
    layer0_outputs(9752) <= not(inputs(88));
    layer0_outputs(9753) <= not((inputs(104)) or (inputs(99)));
    layer0_outputs(9754) <= (inputs(144)) and (inputs(112));
    layer0_outputs(9755) <= not(inputs(173));
    layer0_outputs(9756) <= (inputs(57)) or (inputs(63));
    layer0_outputs(9757) <= (inputs(106)) and not (inputs(39));
    layer0_outputs(9758) <= not(inputs(61)) or (inputs(54));
    layer0_outputs(9759) <= not((inputs(47)) or (inputs(95)));
    layer0_outputs(9760) <= not((inputs(171)) xor (inputs(159)));
    layer0_outputs(9761) <= (inputs(102)) and not (inputs(255));
    layer0_outputs(9762) <= not(inputs(95));
    layer0_outputs(9763) <= inputs(15);
    layer0_outputs(9764) <= (inputs(2)) or (inputs(36));
    layer0_outputs(9765) <= not((inputs(90)) or (inputs(136)));
    layer0_outputs(9766) <= not(inputs(180));
    layer0_outputs(9767) <= not(inputs(50)) or (inputs(113));
    layer0_outputs(9768) <= not(inputs(136)) or (inputs(172));
    layer0_outputs(9769) <= not((inputs(77)) or (inputs(33)));
    layer0_outputs(9770) <= not(inputs(29));
    layer0_outputs(9771) <= inputs(212);
    layer0_outputs(9772) <= not((inputs(105)) or (inputs(38)));
    layer0_outputs(9773) <= not((inputs(200)) xor (inputs(5)));
    layer0_outputs(9774) <= not(inputs(141));
    layer0_outputs(9775) <= inputs(32);
    layer0_outputs(9776) <= inputs(83);
    layer0_outputs(9777) <= not(inputs(55)) or (inputs(202));
    layer0_outputs(9778) <= (inputs(102)) and not (inputs(3));
    layer0_outputs(9779) <= not(inputs(207));
    layer0_outputs(9780) <= not(inputs(136));
    layer0_outputs(9781) <= not(inputs(24));
    layer0_outputs(9782) <= (inputs(54)) or (inputs(113));
    layer0_outputs(9783) <= not(inputs(84)) or (inputs(142));
    layer0_outputs(9784) <= not((inputs(87)) xor (inputs(135)));
    layer0_outputs(9785) <= (inputs(79)) and not (inputs(11));
    layer0_outputs(9786) <= (inputs(203)) xor (inputs(128));
    layer0_outputs(9787) <= not(inputs(135));
    layer0_outputs(9788) <= (inputs(205)) xor (inputs(47));
    layer0_outputs(9789) <= (inputs(44)) xor (inputs(200));
    layer0_outputs(9790) <= not((inputs(171)) xor (inputs(84)));
    layer0_outputs(9791) <= not(inputs(152));
    layer0_outputs(9792) <= not((inputs(31)) or (inputs(37)));
    layer0_outputs(9793) <= not(inputs(165));
    layer0_outputs(9794) <= not((inputs(240)) xor (inputs(210)));
    layer0_outputs(9795) <= not((inputs(185)) or (inputs(189)));
    layer0_outputs(9796) <= not((inputs(124)) or (inputs(26)));
    layer0_outputs(9797) <= inputs(76);
    layer0_outputs(9798) <= not((inputs(247)) or (inputs(226)));
    layer0_outputs(9799) <= not((inputs(92)) xor (inputs(148)));
    layer0_outputs(9800) <= (inputs(41)) and not (inputs(144));
    layer0_outputs(9801) <= not(inputs(35));
    layer0_outputs(9802) <= not(inputs(193)) or (inputs(98));
    layer0_outputs(9803) <= not((inputs(248)) or (inputs(231)));
    layer0_outputs(9804) <= (inputs(97)) and not (inputs(201));
    layer0_outputs(9805) <= (inputs(219)) and not (inputs(172));
    layer0_outputs(9806) <= (inputs(31)) and not (inputs(205));
    layer0_outputs(9807) <= (inputs(107)) xor (inputs(199));
    layer0_outputs(9808) <= not((inputs(152)) and (inputs(187)));
    layer0_outputs(9809) <= inputs(132);
    layer0_outputs(9810) <= not((inputs(227)) xor (inputs(182)));
    layer0_outputs(9811) <= '1';
    layer0_outputs(9812) <= not(inputs(6)) or (inputs(194));
    layer0_outputs(9813) <= inputs(55);
    layer0_outputs(9814) <= not((inputs(155)) xor (inputs(255)));
    layer0_outputs(9815) <= not((inputs(142)) or (inputs(29)));
    layer0_outputs(9816) <= not(inputs(23)) or (inputs(233));
    layer0_outputs(9817) <= (inputs(145)) and not (inputs(244));
    layer0_outputs(9818) <= not(inputs(137));
    layer0_outputs(9819) <= inputs(89);
    layer0_outputs(9820) <= not((inputs(62)) or (inputs(113)));
    layer0_outputs(9821) <= not(inputs(187)) or (inputs(112));
    layer0_outputs(9822) <= not((inputs(15)) or (inputs(154)));
    layer0_outputs(9823) <= not((inputs(80)) xor (inputs(33)));
    layer0_outputs(9824) <= not(inputs(172)) or (inputs(51));
    layer0_outputs(9825) <= (inputs(193)) and not (inputs(72));
    layer0_outputs(9826) <= (inputs(154)) and not (inputs(188));
    layer0_outputs(9827) <= '0';
    layer0_outputs(9828) <= not((inputs(97)) and (inputs(55)));
    layer0_outputs(9829) <= not(inputs(46));
    layer0_outputs(9830) <= '1';
    layer0_outputs(9831) <= not((inputs(235)) or (inputs(219)));
    layer0_outputs(9832) <= not(inputs(121));
    layer0_outputs(9833) <= (inputs(32)) or (inputs(27));
    layer0_outputs(9834) <= (inputs(86)) and not (inputs(232));
    layer0_outputs(9835) <= not((inputs(229)) and (inputs(232)));
    layer0_outputs(9836) <= not(inputs(247));
    layer0_outputs(9837) <= not((inputs(225)) xor (inputs(179)));
    layer0_outputs(9838) <= not(inputs(236));
    layer0_outputs(9839) <= (inputs(205)) and not (inputs(144));
    layer0_outputs(9840) <= (inputs(216)) or (inputs(203));
    layer0_outputs(9841) <= (inputs(123)) or (inputs(7));
    layer0_outputs(9842) <= (inputs(63)) xor (inputs(86));
    layer0_outputs(9843) <= not(inputs(126)) or (inputs(151));
    layer0_outputs(9844) <= not(inputs(203));
    layer0_outputs(9845) <= not((inputs(117)) xor (inputs(37)));
    layer0_outputs(9846) <= (inputs(253)) xor (inputs(162));
    layer0_outputs(9847) <= (inputs(172)) xor (inputs(191));
    layer0_outputs(9848) <= not((inputs(196)) xor (inputs(89)));
    layer0_outputs(9849) <= '0';
    layer0_outputs(9850) <= not(inputs(4));
    layer0_outputs(9851) <= '1';
    layer0_outputs(9852) <= not((inputs(65)) or (inputs(90)));
    layer0_outputs(9853) <= (inputs(161)) xor (inputs(113));
    layer0_outputs(9854) <= (inputs(92)) xor (inputs(79));
    layer0_outputs(9855) <= not(inputs(89));
    layer0_outputs(9856) <= '1';
    layer0_outputs(9857) <= not((inputs(237)) xor (inputs(251)));
    layer0_outputs(9858) <= not(inputs(167)) or (inputs(194));
    layer0_outputs(9859) <= inputs(130);
    layer0_outputs(9860) <= (inputs(247)) and not (inputs(7));
    layer0_outputs(9861) <= inputs(196);
    layer0_outputs(9862) <= (inputs(205)) xor (inputs(103));
    layer0_outputs(9863) <= (inputs(220)) or (inputs(203));
    layer0_outputs(9864) <= (inputs(238)) and not (inputs(139));
    layer0_outputs(9865) <= not(inputs(125));
    layer0_outputs(9866) <= inputs(83);
    layer0_outputs(9867) <= inputs(74);
    layer0_outputs(9868) <= (inputs(216)) and not (inputs(163));
    layer0_outputs(9869) <= inputs(147);
    layer0_outputs(9870) <= (inputs(67)) and (inputs(119));
    layer0_outputs(9871) <= not(inputs(154));
    layer0_outputs(9872) <= (inputs(197)) xor (inputs(60));
    layer0_outputs(9873) <= inputs(75);
    layer0_outputs(9874) <= not((inputs(124)) or (inputs(129)));
    layer0_outputs(9875) <= not((inputs(192)) or (inputs(159)));
    layer0_outputs(9876) <= not(inputs(147));
    layer0_outputs(9877) <= (inputs(234)) xor (inputs(165));
    layer0_outputs(9878) <= (inputs(183)) xor (inputs(166));
    layer0_outputs(9879) <= (inputs(92)) and not (inputs(145));
    layer0_outputs(9880) <= inputs(231);
    layer0_outputs(9881) <= not((inputs(112)) or (inputs(181)));
    layer0_outputs(9882) <= not((inputs(9)) xor (inputs(73)));
    layer0_outputs(9883) <= not((inputs(168)) or (inputs(153)));
    layer0_outputs(9884) <= inputs(216);
    layer0_outputs(9885) <= (inputs(226)) or (inputs(232));
    layer0_outputs(9886) <= (inputs(149)) and not (inputs(67));
    layer0_outputs(9887) <= (inputs(95)) xor (inputs(139));
    layer0_outputs(9888) <= (inputs(171)) xor (inputs(179));
    layer0_outputs(9889) <= (inputs(188)) and not (inputs(110));
    layer0_outputs(9890) <= (inputs(126)) or (inputs(54));
    layer0_outputs(9891) <= not((inputs(49)) xor (inputs(51)));
    layer0_outputs(9892) <= not(inputs(220)) or (inputs(17));
    layer0_outputs(9893) <= not(inputs(233));
    layer0_outputs(9894) <= not((inputs(216)) xor (inputs(159)));
    layer0_outputs(9895) <= inputs(229);
    layer0_outputs(9896) <= not(inputs(192)) or (inputs(13));
    layer0_outputs(9897) <= not(inputs(198));
    layer0_outputs(9898) <= (inputs(90)) and not (inputs(146));
    layer0_outputs(9899) <= '0';
    layer0_outputs(9900) <= not((inputs(34)) or (inputs(23)));
    layer0_outputs(9901) <= (inputs(40)) xor (inputs(10));
    layer0_outputs(9902) <= (inputs(130)) and not (inputs(55));
    layer0_outputs(9903) <= not(inputs(231)) or (inputs(211));
    layer0_outputs(9904) <= not(inputs(18));
    layer0_outputs(9905) <= not((inputs(242)) or (inputs(237)));
    layer0_outputs(9906) <= not(inputs(155)) or (inputs(94));
    layer0_outputs(9907) <= inputs(134);
    layer0_outputs(9908) <= not(inputs(62));
    layer0_outputs(9909) <= (inputs(74)) or (inputs(58));
    layer0_outputs(9910) <= (inputs(210)) xor (inputs(139));
    layer0_outputs(9911) <= inputs(137);
    layer0_outputs(9912) <= inputs(59);
    layer0_outputs(9913) <= inputs(29);
    layer0_outputs(9914) <= (inputs(195)) and (inputs(134));
    layer0_outputs(9915) <= inputs(7);
    layer0_outputs(9916) <= not(inputs(89)) or (inputs(249));
    layer0_outputs(9917) <= not(inputs(84)) or (inputs(63));
    layer0_outputs(9918) <= inputs(61);
    layer0_outputs(9919) <= not(inputs(159)) or (inputs(138));
    layer0_outputs(9920) <= not(inputs(186));
    layer0_outputs(9921) <= not((inputs(5)) xor (inputs(9)));
    layer0_outputs(9922) <= not(inputs(26));
    layer0_outputs(9923) <= not(inputs(78));
    layer0_outputs(9924) <= inputs(140);
    layer0_outputs(9925) <= (inputs(237)) and (inputs(191));
    layer0_outputs(9926) <= not(inputs(152));
    layer0_outputs(9927) <= inputs(154);
    layer0_outputs(9928) <= not((inputs(231)) xor (inputs(132)));
    layer0_outputs(9929) <= not((inputs(193)) or (inputs(203)));
    layer0_outputs(9930) <= not((inputs(86)) or (inputs(163)));
    layer0_outputs(9931) <= not(inputs(99)) or (inputs(141));
    layer0_outputs(9932) <= not(inputs(78));
    layer0_outputs(9933) <= not(inputs(22)) or (inputs(232));
    layer0_outputs(9934) <= (inputs(127)) or (inputs(234));
    layer0_outputs(9935) <= (inputs(167)) or (inputs(56));
    layer0_outputs(9936) <= (inputs(196)) and not (inputs(8));
    layer0_outputs(9937) <= not((inputs(164)) and (inputs(67)));
    layer0_outputs(9938) <= (inputs(74)) and not (inputs(152));
    layer0_outputs(9939) <= inputs(68);
    layer0_outputs(9940) <= (inputs(154)) and not (inputs(51));
    layer0_outputs(9941) <= inputs(237);
    layer0_outputs(9942) <= inputs(39);
    layer0_outputs(9943) <= not((inputs(13)) or (inputs(208)));
    layer0_outputs(9944) <= not((inputs(196)) xor (inputs(9)));
    layer0_outputs(9945) <= not((inputs(81)) or (inputs(98)));
    layer0_outputs(9946) <= not(inputs(240));
    layer0_outputs(9947) <= not(inputs(72)) or (inputs(36));
    layer0_outputs(9948) <= not(inputs(171));
    layer0_outputs(9949) <= (inputs(91)) xor (inputs(95));
    layer0_outputs(9950) <= not((inputs(200)) or (inputs(206)));
    layer0_outputs(9951) <= inputs(164);
    layer0_outputs(9952) <= not((inputs(118)) or (inputs(249)));
    layer0_outputs(9953) <= (inputs(58)) and not (inputs(124));
    layer0_outputs(9954) <= not((inputs(163)) or (inputs(74)));
    layer0_outputs(9955) <= (inputs(139)) or (inputs(226));
    layer0_outputs(9956) <= (inputs(78)) and not (inputs(159));
    layer0_outputs(9957) <= not((inputs(80)) or (inputs(81)));
    layer0_outputs(9958) <= not((inputs(0)) xor (inputs(67)));
    layer0_outputs(9959) <= not(inputs(24));
    layer0_outputs(9960) <= not(inputs(59)) or (inputs(209));
    layer0_outputs(9961) <= inputs(120);
    layer0_outputs(9962) <= not((inputs(118)) and (inputs(76)));
    layer0_outputs(9963) <= not(inputs(230));
    layer0_outputs(9964) <= inputs(87);
    layer0_outputs(9965) <= not((inputs(54)) and (inputs(39)));
    layer0_outputs(9966) <= (inputs(78)) and not (inputs(204));
    layer0_outputs(9967) <= not(inputs(197)) or (inputs(89));
    layer0_outputs(9968) <= not((inputs(74)) or (inputs(2)));
    layer0_outputs(9969) <= not(inputs(153));
    layer0_outputs(9970) <= not(inputs(124)) or (inputs(33));
    layer0_outputs(9971) <= inputs(139);
    layer0_outputs(9972) <= (inputs(182)) or (inputs(192));
    layer0_outputs(9973) <= not(inputs(83));
    layer0_outputs(9974) <= (inputs(167)) and (inputs(249));
    layer0_outputs(9975) <= not(inputs(176));
    layer0_outputs(9976) <= (inputs(47)) or (inputs(237));
    layer0_outputs(9977) <= not(inputs(188));
    layer0_outputs(9978) <= inputs(221);
    layer0_outputs(9979) <= not(inputs(141)) or (inputs(252));
    layer0_outputs(9980) <= not((inputs(90)) or (inputs(162)));
    layer0_outputs(9981) <= not(inputs(121));
    layer0_outputs(9982) <= not(inputs(13));
    layer0_outputs(9983) <= inputs(93);
    layer0_outputs(9984) <= (inputs(111)) xor (inputs(77));
    layer0_outputs(9985) <= not(inputs(181));
    layer0_outputs(9986) <= '1';
    layer0_outputs(9987) <= not((inputs(191)) or (inputs(24)));
    layer0_outputs(9988) <= not((inputs(172)) or (inputs(4)));
    layer0_outputs(9989) <= (inputs(106)) or (inputs(108));
    layer0_outputs(9990) <= not(inputs(196)) or (inputs(101));
    layer0_outputs(9991) <= not(inputs(68)) or (inputs(191));
    layer0_outputs(9992) <= (inputs(20)) and not (inputs(147));
    layer0_outputs(9993) <= '1';
    layer0_outputs(9994) <= not(inputs(164));
    layer0_outputs(9995) <= inputs(169);
    layer0_outputs(9996) <= (inputs(33)) xor (inputs(87));
    layer0_outputs(9997) <= not((inputs(171)) or (inputs(177)));
    layer0_outputs(9998) <= not((inputs(22)) xor (inputs(58)));
    layer0_outputs(9999) <= (inputs(81)) and not (inputs(15));
    layer0_outputs(10000) <= inputs(91);
    layer0_outputs(10001) <= (inputs(215)) or (inputs(49));
    layer0_outputs(10002) <= not(inputs(101));
    layer0_outputs(10003) <= not((inputs(245)) xor (inputs(143)));
    layer0_outputs(10004) <= not((inputs(0)) xor (inputs(44)));
    layer0_outputs(10005) <= not(inputs(146));
    layer0_outputs(10006) <= inputs(37);
    layer0_outputs(10007) <= (inputs(229)) and (inputs(227));
    layer0_outputs(10008) <= not((inputs(206)) xor (inputs(125)));
    layer0_outputs(10009) <= not((inputs(233)) or (inputs(227)));
    layer0_outputs(10010) <= not((inputs(124)) or (inputs(105)));
    layer0_outputs(10011) <= not(inputs(99)) or (inputs(108));
    layer0_outputs(10012) <= not(inputs(213)) or (inputs(13));
    layer0_outputs(10013) <= inputs(188);
    layer0_outputs(10014) <= (inputs(92)) or (inputs(151));
    layer0_outputs(10015) <= (inputs(168)) and not (inputs(156));
    layer0_outputs(10016) <= not((inputs(64)) or (inputs(177)));
    layer0_outputs(10017) <= (inputs(60)) and not (inputs(57));
    layer0_outputs(10018) <= (inputs(227)) and not (inputs(117));
    layer0_outputs(10019) <= not(inputs(44)) or (inputs(135));
    layer0_outputs(10020) <= (inputs(150)) xor (inputs(153));
    layer0_outputs(10021) <= '1';
    layer0_outputs(10022) <= (inputs(29)) xor (inputs(72));
    layer0_outputs(10023) <= (inputs(73)) or (inputs(186));
    layer0_outputs(10024) <= (inputs(240)) or (inputs(182));
    layer0_outputs(10025) <= inputs(208);
    layer0_outputs(10026) <= (inputs(3)) or (inputs(250));
    layer0_outputs(10027) <= not(inputs(242));
    layer0_outputs(10028) <= (inputs(245)) and not (inputs(236));
    layer0_outputs(10029) <= not(inputs(245)) or (inputs(130));
    layer0_outputs(10030) <= not((inputs(102)) xor (inputs(113)));
    layer0_outputs(10031) <= inputs(228);
    layer0_outputs(10032) <= inputs(196);
    layer0_outputs(10033) <= not(inputs(84));
    layer0_outputs(10034) <= (inputs(13)) xor (inputs(44));
    layer0_outputs(10035) <= (inputs(30)) and not (inputs(130));
    layer0_outputs(10036) <= (inputs(89)) and not (inputs(220));
    layer0_outputs(10037) <= (inputs(184)) and (inputs(240));
    layer0_outputs(10038) <= not(inputs(105));
    layer0_outputs(10039) <= not(inputs(150));
    layer0_outputs(10040) <= inputs(83);
    layer0_outputs(10041) <= not((inputs(73)) or (inputs(107)));
    layer0_outputs(10042) <= not((inputs(240)) or (inputs(135)));
    layer0_outputs(10043) <= not(inputs(201));
    layer0_outputs(10044) <= (inputs(196)) xor (inputs(194));
    layer0_outputs(10045) <= (inputs(149)) and not (inputs(39));
    layer0_outputs(10046) <= inputs(135);
    layer0_outputs(10047) <= not((inputs(140)) xor (inputs(35)));
    layer0_outputs(10048) <= (inputs(164)) and (inputs(229));
    layer0_outputs(10049) <= '0';
    layer0_outputs(10050) <= (inputs(76)) xor (inputs(225));
    layer0_outputs(10051) <= inputs(23);
    layer0_outputs(10052) <= (inputs(171)) or (inputs(162));
    layer0_outputs(10053) <= not((inputs(111)) xor (inputs(90)));
    layer0_outputs(10054) <= not((inputs(26)) xor (inputs(230)));
    layer0_outputs(10055) <= (inputs(127)) xor (inputs(106));
    layer0_outputs(10056) <= not((inputs(38)) or (inputs(130)));
    layer0_outputs(10057) <= inputs(122);
    layer0_outputs(10058) <= not((inputs(187)) and (inputs(210)));
    layer0_outputs(10059) <= (inputs(230)) or (inputs(229));
    layer0_outputs(10060) <= not(inputs(173)) or (inputs(103));
    layer0_outputs(10061) <= inputs(60);
    layer0_outputs(10062) <= not(inputs(147));
    layer0_outputs(10063) <= '1';
    layer0_outputs(10064) <= not(inputs(162)) or (inputs(96));
    layer0_outputs(10065) <= not(inputs(141)) or (inputs(240));
    layer0_outputs(10066) <= not(inputs(151));
    layer0_outputs(10067) <= not((inputs(200)) or (inputs(127)));
    layer0_outputs(10068) <= not(inputs(130));
    layer0_outputs(10069) <= not(inputs(30));
    layer0_outputs(10070) <= (inputs(229)) xor (inputs(245));
    layer0_outputs(10071) <= not(inputs(227));
    layer0_outputs(10072) <= not((inputs(72)) xor (inputs(20)));
    layer0_outputs(10073) <= not((inputs(50)) xor (inputs(10)));
    layer0_outputs(10074) <= not((inputs(83)) or (inputs(145)));
    layer0_outputs(10075) <= (inputs(101)) and not (inputs(191));
    layer0_outputs(10076) <= (inputs(115)) or (inputs(64));
    layer0_outputs(10077) <= inputs(126);
    layer0_outputs(10078) <= not((inputs(195)) xor (inputs(144)));
    layer0_outputs(10079) <= not(inputs(102));
    layer0_outputs(10080) <= (inputs(149)) or (inputs(86));
    layer0_outputs(10081) <= not((inputs(1)) and (inputs(184)));
    layer0_outputs(10082) <= not((inputs(168)) xor (inputs(34)));
    layer0_outputs(10083) <= not(inputs(131)) or (inputs(25));
    layer0_outputs(10084) <= not((inputs(192)) xor (inputs(218)));
    layer0_outputs(10085) <= (inputs(185)) or (inputs(105));
    layer0_outputs(10086) <= not(inputs(89));
    layer0_outputs(10087) <= not(inputs(249)) or (inputs(101));
    layer0_outputs(10088) <= inputs(21);
    layer0_outputs(10089) <= not(inputs(82));
    layer0_outputs(10090) <= (inputs(228)) xor (inputs(198));
    layer0_outputs(10091) <= not((inputs(51)) xor (inputs(130)));
    layer0_outputs(10092) <= not(inputs(229));
    layer0_outputs(10093) <= not(inputs(240));
    layer0_outputs(10094) <= not(inputs(83)) or (inputs(99));
    layer0_outputs(10095) <= inputs(205);
    layer0_outputs(10096) <= not(inputs(234));
    layer0_outputs(10097) <= not(inputs(188));
    layer0_outputs(10098) <= inputs(146);
    layer0_outputs(10099) <= inputs(185);
    layer0_outputs(10100) <= (inputs(167)) or (inputs(34));
    layer0_outputs(10101) <= inputs(98);
    layer0_outputs(10102) <= (inputs(175)) and not (inputs(248));
    layer0_outputs(10103) <= (inputs(89)) or (inputs(135));
    layer0_outputs(10104) <= inputs(38);
    layer0_outputs(10105) <= not(inputs(236));
    layer0_outputs(10106) <= (inputs(57)) and not (inputs(145));
    layer0_outputs(10107) <= not((inputs(33)) xor (inputs(202)));
    layer0_outputs(10108) <= not((inputs(241)) or (inputs(145)));
    layer0_outputs(10109) <= not(inputs(27));
    layer0_outputs(10110) <= (inputs(201)) and (inputs(177));
    layer0_outputs(10111) <= inputs(50);
    layer0_outputs(10112) <= not(inputs(96));
    layer0_outputs(10113) <= not((inputs(223)) xor (inputs(67)));
    layer0_outputs(10114) <= inputs(177);
    layer0_outputs(10115) <= inputs(81);
    layer0_outputs(10116) <= inputs(182);
    layer0_outputs(10117) <= inputs(144);
    layer0_outputs(10118) <= not(inputs(234)) or (inputs(44));
    layer0_outputs(10119) <= not((inputs(252)) xor (inputs(140)));
    layer0_outputs(10120) <= not((inputs(21)) or (inputs(159)));
    layer0_outputs(10121) <= not(inputs(228)) or (inputs(18));
    layer0_outputs(10122) <= inputs(99);
    layer0_outputs(10123) <= (inputs(231)) and not (inputs(108));
    layer0_outputs(10124) <= inputs(46);
    layer0_outputs(10125) <= not(inputs(116));
    layer0_outputs(10126) <= not(inputs(86)) or (inputs(54));
    layer0_outputs(10127) <= (inputs(194)) or (inputs(7));
    layer0_outputs(10128) <= not((inputs(209)) or (inputs(228)));
    layer0_outputs(10129) <= not(inputs(176)) or (inputs(128));
    layer0_outputs(10130) <= not(inputs(239));
    layer0_outputs(10131) <= (inputs(228)) and not (inputs(46));
    layer0_outputs(10132) <= inputs(185);
    layer0_outputs(10133) <= not((inputs(84)) or (inputs(255)));
    layer0_outputs(10134) <= (inputs(181)) and not (inputs(81));
    layer0_outputs(10135) <= not((inputs(76)) or (inputs(80)));
    layer0_outputs(10136) <= (inputs(182)) and not (inputs(223));
    layer0_outputs(10137) <= not(inputs(33));
    layer0_outputs(10138) <= not(inputs(91)) or (inputs(229));
    layer0_outputs(10139) <= not((inputs(244)) or (inputs(228)));
    layer0_outputs(10140) <= inputs(26);
    layer0_outputs(10141) <= inputs(204);
    layer0_outputs(10142) <= (inputs(56)) and not (inputs(39));
    layer0_outputs(10143) <= not(inputs(100));
    layer0_outputs(10144) <= not((inputs(188)) xor (inputs(174)));
    layer0_outputs(10145) <= not((inputs(112)) or (inputs(218)));
    layer0_outputs(10146) <= not((inputs(172)) xor (inputs(29)));
    layer0_outputs(10147) <= (inputs(173)) xor (inputs(172));
    layer0_outputs(10148) <= (inputs(201)) xor (inputs(178));
    layer0_outputs(10149) <= not(inputs(98));
    layer0_outputs(10150) <= not((inputs(139)) xor (inputs(124)));
    layer0_outputs(10151) <= (inputs(202)) xor (inputs(41));
    layer0_outputs(10152) <= inputs(209);
    layer0_outputs(10153) <= not(inputs(140)) or (inputs(67));
    layer0_outputs(10154) <= not(inputs(190));
    layer0_outputs(10155) <= not((inputs(81)) xor (inputs(87)));
    layer0_outputs(10156) <= not(inputs(166)) or (inputs(171));
    layer0_outputs(10157) <= (inputs(162)) or (inputs(77));
    layer0_outputs(10158) <= (inputs(117)) or (inputs(29));
    layer0_outputs(10159) <= (inputs(67)) or (inputs(168));
    layer0_outputs(10160) <= not((inputs(87)) or (inputs(28)));
    layer0_outputs(10161) <= (inputs(121)) and not (inputs(35));
    layer0_outputs(10162) <= (inputs(142)) and not (inputs(30));
    layer0_outputs(10163) <= (inputs(10)) or (inputs(79));
    layer0_outputs(10164) <= not((inputs(115)) or (inputs(143)));
    layer0_outputs(10165) <= (inputs(196)) or (inputs(216));
    layer0_outputs(10166) <= not(inputs(145));
    layer0_outputs(10167) <= (inputs(238)) xor (inputs(250));
    layer0_outputs(10168) <= not(inputs(74)) or (inputs(188));
    layer0_outputs(10169) <= not(inputs(20));
    layer0_outputs(10170) <= not(inputs(206));
    layer0_outputs(10171) <= inputs(158);
    layer0_outputs(10172) <= not(inputs(24)) or (inputs(238));
    layer0_outputs(10173) <= not(inputs(102));
    layer0_outputs(10174) <= not((inputs(43)) xor (inputs(125)));
    layer0_outputs(10175) <= not(inputs(79)) or (inputs(54));
    layer0_outputs(10176) <= (inputs(233)) xor (inputs(234));
    layer0_outputs(10177) <= not((inputs(57)) xor (inputs(58)));
    layer0_outputs(10178) <= not((inputs(209)) or (inputs(171)));
    layer0_outputs(10179) <= not(inputs(214));
    layer0_outputs(10180) <= not(inputs(48));
    layer0_outputs(10181) <= (inputs(165)) or (inputs(119));
    layer0_outputs(10182) <= (inputs(210)) or (inputs(253));
    layer0_outputs(10183) <= inputs(46);
    layer0_outputs(10184) <= not((inputs(53)) xor (inputs(237)));
    layer0_outputs(10185) <= inputs(174);
    layer0_outputs(10186) <= not((inputs(5)) xor (inputs(70)));
    layer0_outputs(10187) <= (inputs(153)) and not (inputs(50));
    layer0_outputs(10188) <= not((inputs(125)) or (inputs(141)));
    layer0_outputs(10189) <= not(inputs(244)) or (inputs(224));
    layer0_outputs(10190) <= inputs(168);
    layer0_outputs(10191) <= not(inputs(25)) or (inputs(133));
    layer0_outputs(10192) <= inputs(178);
    layer0_outputs(10193) <= (inputs(119)) and not (inputs(64));
    layer0_outputs(10194) <= (inputs(49)) or (inputs(239));
    layer0_outputs(10195) <= not((inputs(218)) or (inputs(1)));
    layer0_outputs(10196) <= inputs(73);
    layer0_outputs(10197) <= not((inputs(60)) or (inputs(8)));
    layer0_outputs(10198) <= not(inputs(199));
    layer0_outputs(10199) <= not(inputs(191)) or (inputs(153));
    layer0_outputs(10200) <= not(inputs(246));
    layer0_outputs(10201) <= inputs(123);
    layer0_outputs(10202) <= not(inputs(177));
    layer0_outputs(10203) <= not(inputs(116)) or (inputs(144));
    layer0_outputs(10204) <= (inputs(91)) and not (inputs(128));
    layer0_outputs(10205) <= (inputs(31)) or (inputs(192));
    layer0_outputs(10206) <= (inputs(214)) xor (inputs(33));
    layer0_outputs(10207) <= not((inputs(82)) or (inputs(175)));
    layer0_outputs(10208) <= not(inputs(42)) or (inputs(158));
    layer0_outputs(10209) <= not(inputs(56)) or (inputs(198));
    layer0_outputs(10210) <= not((inputs(120)) and (inputs(8)));
    layer0_outputs(10211) <= inputs(164);
    layer0_outputs(10212) <= not((inputs(252)) xor (inputs(193)));
    layer0_outputs(10213) <= (inputs(122)) xor (inputs(137));
    layer0_outputs(10214) <= not(inputs(22)) or (inputs(143));
    layer0_outputs(10215) <= (inputs(90)) and not (inputs(165));
    layer0_outputs(10216) <= (inputs(124)) or (inputs(229));
    layer0_outputs(10217) <= (inputs(190)) or (inputs(54));
    layer0_outputs(10218) <= not((inputs(171)) xor (inputs(179)));
    layer0_outputs(10219) <= not((inputs(248)) or (inputs(47)));
    layer0_outputs(10220) <= inputs(233);
    layer0_outputs(10221) <= (inputs(94)) or (inputs(176));
    layer0_outputs(10222) <= inputs(150);
    layer0_outputs(10223) <= not(inputs(84)) or (inputs(155));
    layer0_outputs(10224) <= not((inputs(131)) and (inputs(211)));
    layer0_outputs(10225) <= inputs(142);
    layer0_outputs(10226) <= inputs(214);
    layer0_outputs(10227) <= not(inputs(158));
    layer0_outputs(10228) <= not(inputs(46));
    layer0_outputs(10229) <= inputs(210);
    layer0_outputs(10230) <= not((inputs(175)) or (inputs(170)));
    layer0_outputs(10231) <= not(inputs(51));
    layer0_outputs(10232) <= (inputs(218)) and not (inputs(132));
    layer0_outputs(10233) <= (inputs(234)) and (inputs(185));
    layer0_outputs(10234) <= (inputs(64)) xor (inputs(39));
    layer0_outputs(10235) <= (inputs(231)) and not (inputs(50));
    layer0_outputs(10236) <= (inputs(211)) xor (inputs(213));
    layer0_outputs(10237) <= (inputs(49)) and not (inputs(97));
    layer0_outputs(10238) <= not(inputs(235)) or (inputs(123));
    layer0_outputs(10239) <= (inputs(175)) or (inputs(11));
    layer0_outputs(10240) <= not((inputs(97)) or (inputs(119)));
    layer0_outputs(10241) <= not((inputs(155)) or (inputs(48)));
    layer0_outputs(10242) <= (inputs(202)) and not (inputs(109));
    layer0_outputs(10243) <= not(inputs(194));
    layer0_outputs(10244) <= not(inputs(214));
    layer0_outputs(10245) <= (inputs(167)) and not (inputs(208));
    layer0_outputs(10246) <= not(inputs(229));
    layer0_outputs(10247) <= (inputs(181)) or (inputs(238));
    layer0_outputs(10248) <= not(inputs(68));
    layer0_outputs(10249) <= (inputs(236)) xor (inputs(60));
    layer0_outputs(10250) <= not((inputs(96)) or (inputs(207)));
    layer0_outputs(10251) <= (inputs(4)) xor (inputs(43));
    layer0_outputs(10252) <= inputs(100);
    layer0_outputs(10253) <= inputs(168);
    layer0_outputs(10254) <= (inputs(255)) or (inputs(57));
    layer0_outputs(10255) <= (inputs(223)) xor (inputs(163));
    layer0_outputs(10256) <= not(inputs(89)) or (inputs(23));
    layer0_outputs(10257) <= not(inputs(21));
    layer0_outputs(10258) <= not((inputs(161)) or (inputs(194)));
    layer0_outputs(10259) <= not(inputs(97)) or (inputs(254));
    layer0_outputs(10260) <= '0';
    layer0_outputs(10261) <= not((inputs(148)) xor (inputs(68)));
    layer0_outputs(10262) <= not((inputs(86)) xor (inputs(113)));
    layer0_outputs(10263) <= inputs(187);
    layer0_outputs(10264) <= not(inputs(136)) or (inputs(212));
    layer0_outputs(10265) <= not(inputs(166)) or (inputs(205));
    layer0_outputs(10266) <= not(inputs(52));
    layer0_outputs(10267) <= (inputs(38)) and (inputs(59));
    layer0_outputs(10268) <= not((inputs(73)) xor (inputs(126)));
    layer0_outputs(10269) <= not(inputs(146));
    layer0_outputs(10270) <= not(inputs(162));
    layer0_outputs(10271) <= not(inputs(172)) or (inputs(120));
    layer0_outputs(10272) <= inputs(112);
    layer0_outputs(10273) <= not((inputs(240)) or (inputs(76)));
    layer0_outputs(10274) <= inputs(57);
    layer0_outputs(10275) <= (inputs(206)) or (inputs(220));
    layer0_outputs(10276) <= inputs(106);
    layer0_outputs(10277) <= inputs(91);
    layer0_outputs(10278) <= (inputs(222)) and not (inputs(31));
    layer0_outputs(10279) <= not((inputs(82)) xor (inputs(31)));
    layer0_outputs(10280) <= not((inputs(148)) xor (inputs(120)));
    layer0_outputs(10281) <= (inputs(50)) or (inputs(165));
    layer0_outputs(10282) <= (inputs(170)) or (inputs(26));
    layer0_outputs(10283) <= (inputs(95)) or (inputs(7));
    layer0_outputs(10284) <= not((inputs(243)) xor (inputs(236)));
    layer0_outputs(10285) <= not(inputs(121)) or (inputs(147));
    layer0_outputs(10286) <= (inputs(5)) xor (inputs(93));
    layer0_outputs(10287) <= not(inputs(4));
    layer0_outputs(10288) <= (inputs(7)) and (inputs(88));
    layer0_outputs(10289) <= (inputs(212)) and (inputs(210));
    layer0_outputs(10290) <= (inputs(242)) or (inputs(177));
    layer0_outputs(10291) <= not((inputs(165)) or (inputs(5)));
    layer0_outputs(10292) <= not(inputs(134)) or (inputs(114));
    layer0_outputs(10293) <= not(inputs(78));
    layer0_outputs(10294) <= not(inputs(195));
    layer0_outputs(10295) <= not(inputs(232)) or (inputs(253));
    layer0_outputs(10296) <= (inputs(28)) and (inputs(255));
    layer0_outputs(10297) <= inputs(104);
    layer0_outputs(10298) <= not((inputs(252)) or (inputs(165)));
    layer0_outputs(10299) <= (inputs(197)) or (inputs(48));
    layer0_outputs(10300) <= not((inputs(244)) or (inputs(124)));
    layer0_outputs(10301) <= not(inputs(172)) or (inputs(47));
    layer0_outputs(10302) <= not(inputs(98));
    layer0_outputs(10303) <= (inputs(128)) or (inputs(240));
    layer0_outputs(10304) <= not(inputs(233));
    layer0_outputs(10305) <= inputs(114);
    layer0_outputs(10306) <= inputs(242);
    layer0_outputs(10307) <= inputs(243);
    layer0_outputs(10308) <= not(inputs(45));
    layer0_outputs(10309) <= not((inputs(4)) or (inputs(180)));
    layer0_outputs(10310) <= not((inputs(78)) or (inputs(54)));
    layer0_outputs(10311) <= not(inputs(11));
    layer0_outputs(10312) <= (inputs(21)) or (inputs(74));
    layer0_outputs(10313) <= (inputs(160)) xor (inputs(56));
    layer0_outputs(10314) <= (inputs(110)) and not (inputs(80));
    layer0_outputs(10315) <= not(inputs(199)) or (inputs(109));
    layer0_outputs(10316) <= (inputs(46)) xor (inputs(173));
    layer0_outputs(10317) <= inputs(113);
    layer0_outputs(10318) <= (inputs(5)) xor (inputs(137));
    layer0_outputs(10319) <= (inputs(67)) or (inputs(212));
    layer0_outputs(10320) <= (inputs(146)) or (inputs(109));
    layer0_outputs(10321) <= (inputs(112)) and (inputs(17));
    layer0_outputs(10322) <= (inputs(184)) and not (inputs(195));
    layer0_outputs(10323) <= not((inputs(243)) or (inputs(116)));
    layer0_outputs(10324) <= not((inputs(253)) or (inputs(219)));
    layer0_outputs(10325) <= (inputs(213)) or (inputs(68));
    layer0_outputs(10326) <= not((inputs(43)) xor (inputs(197)));
    layer0_outputs(10327) <= not(inputs(41)) or (inputs(166));
    layer0_outputs(10328) <= not(inputs(61)) or (inputs(98));
    layer0_outputs(10329) <= not(inputs(214)) or (inputs(136));
    layer0_outputs(10330) <= inputs(25);
    layer0_outputs(10331) <= not(inputs(127));
    layer0_outputs(10332) <= not((inputs(235)) xor (inputs(98)));
    layer0_outputs(10333) <= inputs(58);
    layer0_outputs(10334) <= not((inputs(83)) xor (inputs(108)));
    layer0_outputs(10335) <= not(inputs(254));
    layer0_outputs(10336) <= not(inputs(130));
    layer0_outputs(10337) <= (inputs(86)) or (inputs(31));
    layer0_outputs(10338) <= not(inputs(232)) or (inputs(206));
    layer0_outputs(10339) <= not(inputs(61));
    layer0_outputs(10340) <= '1';
    layer0_outputs(10341) <= inputs(40);
    layer0_outputs(10342) <= not(inputs(69)) or (inputs(79));
    layer0_outputs(10343) <= not(inputs(8));
    layer0_outputs(10344) <= (inputs(210)) and not (inputs(239));
    layer0_outputs(10345) <= (inputs(232)) xor (inputs(22));
    layer0_outputs(10346) <= inputs(175);
    layer0_outputs(10347) <= not((inputs(195)) or (inputs(207)));
    layer0_outputs(10348) <= (inputs(195)) and not (inputs(240));
    layer0_outputs(10349) <= not(inputs(58)) or (inputs(114));
    layer0_outputs(10350) <= (inputs(45)) or (inputs(121));
    layer0_outputs(10351) <= (inputs(71)) and not (inputs(166));
    layer0_outputs(10352) <= not((inputs(54)) xor (inputs(212)));
    layer0_outputs(10353) <= inputs(145);
    layer0_outputs(10354) <= not(inputs(68)) or (inputs(143));
    layer0_outputs(10355) <= (inputs(113)) xor (inputs(140));
    layer0_outputs(10356) <= not((inputs(235)) xor (inputs(165)));
    layer0_outputs(10357) <= not(inputs(25));
    layer0_outputs(10358) <= '1';
    layer0_outputs(10359) <= not(inputs(55)) or (inputs(205));
    layer0_outputs(10360) <= not(inputs(122));
    layer0_outputs(10361) <= (inputs(118)) or (inputs(68));
    layer0_outputs(10362) <= (inputs(235)) xor (inputs(9));
    layer0_outputs(10363) <= not((inputs(245)) or (inputs(100)));
    layer0_outputs(10364) <= not(inputs(151));
    layer0_outputs(10365) <= (inputs(80)) xor (inputs(20));
    layer0_outputs(10366) <= not(inputs(74));
    layer0_outputs(10367) <= (inputs(237)) xor (inputs(225));
    layer0_outputs(10368) <= (inputs(18)) and not (inputs(238));
    layer0_outputs(10369) <= (inputs(48)) or (inputs(249));
    layer0_outputs(10370) <= not((inputs(133)) or (inputs(182)));
    layer0_outputs(10371) <= not(inputs(123)) or (inputs(63));
    layer0_outputs(10372) <= inputs(180);
    layer0_outputs(10373) <= (inputs(61)) or (inputs(107));
    layer0_outputs(10374) <= not(inputs(118)) or (inputs(52));
    layer0_outputs(10375) <= not(inputs(4));
    layer0_outputs(10376) <= (inputs(185)) or (inputs(162));
    layer0_outputs(10377) <= not((inputs(164)) xor (inputs(82)));
    layer0_outputs(10378) <= not((inputs(114)) or (inputs(113)));
    layer0_outputs(10379) <= (inputs(27)) and not (inputs(97));
    layer0_outputs(10380) <= not((inputs(157)) xor (inputs(211)));
    layer0_outputs(10381) <= (inputs(224)) and not (inputs(184));
    layer0_outputs(10382) <= not((inputs(120)) or (inputs(45)));
    layer0_outputs(10383) <= inputs(104);
    layer0_outputs(10384) <= (inputs(116)) xor (inputs(139));
    layer0_outputs(10385) <= inputs(217);
    layer0_outputs(10386) <= not(inputs(160)) or (inputs(127));
    layer0_outputs(10387) <= not(inputs(250)) or (inputs(131));
    layer0_outputs(10388) <= not((inputs(208)) or (inputs(214)));
    layer0_outputs(10389) <= not(inputs(91)) or (inputs(175));
    layer0_outputs(10390) <= not((inputs(115)) xor (inputs(84)));
    layer0_outputs(10391) <= not((inputs(17)) or (inputs(125)));
    layer0_outputs(10392) <= (inputs(26)) and not (inputs(205));
    layer0_outputs(10393) <= not(inputs(232)) or (inputs(34));
    layer0_outputs(10394) <= not((inputs(149)) xor (inputs(193)));
    layer0_outputs(10395) <= (inputs(75)) xor (inputs(104));
    layer0_outputs(10396) <= (inputs(162)) xor (inputs(135));
    layer0_outputs(10397) <= (inputs(24)) xor (inputs(138));
    layer0_outputs(10398) <= (inputs(94)) and not (inputs(240));
    layer0_outputs(10399) <= (inputs(211)) xor (inputs(213));
    layer0_outputs(10400) <= (inputs(174)) xor (inputs(117));
    layer0_outputs(10401) <= not(inputs(106)) or (inputs(233));
    layer0_outputs(10402) <= (inputs(26)) xor (inputs(247));
    layer0_outputs(10403) <= not((inputs(242)) or (inputs(248)));
    layer0_outputs(10404) <= not((inputs(62)) or (inputs(13)));
    layer0_outputs(10405) <= inputs(117);
    layer0_outputs(10406) <= (inputs(37)) and not (inputs(166));
    layer0_outputs(10407) <= inputs(15);
    layer0_outputs(10408) <= '0';
    layer0_outputs(10409) <= (inputs(92)) and not (inputs(112));
    layer0_outputs(10410) <= not((inputs(84)) or (inputs(68)));
    layer0_outputs(10411) <= (inputs(147)) and (inputs(116));
    layer0_outputs(10412) <= (inputs(203)) xor (inputs(235));
    layer0_outputs(10413) <= not((inputs(104)) xor (inputs(172)));
    layer0_outputs(10414) <= (inputs(236)) or (inputs(96));
    layer0_outputs(10415) <= not(inputs(58)) or (inputs(103));
    layer0_outputs(10416) <= not((inputs(182)) or (inputs(190)));
    layer0_outputs(10417) <= (inputs(212)) or (inputs(27));
    layer0_outputs(10418) <= not(inputs(196));
    layer0_outputs(10419) <= (inputs(27)) and not (inputs(147));
    layer0_outputs(10420) <= not((inputs(103)) and (inputs(8)));
    layer0_outputs(10421) <= not(inputs(136)) or (inputs(4));
    layer0_outputs(10422) <= not((inputs(216)) xor (inputs(227)));
    layer0_outputs(10423) <= not((inputs(132)) or (inputs(183)));
    layer0_outputs(10424) <= (inputs(25)) xor (inputs(239));
    layer0_outputs(10425) <= not((inputs(90)) xor (inputs(18)));
    layer0_outputs(10426) <= not(inputs(66));
    layer0_outputs(10427) <= (inputs(179)) or (inputs(106));
    layer0_outputs(10428) <= not(inputs(114));
    layer0_outputs(10429) <= (inputs(1)) and not (inputs(170));
    layer0_outputs(10430) <= (inputs(20)) and not (inputs(15));
    layer0_outputs(10431) <= (inputs(211)) and not (inputs(10));
    layer0_outputs(10432) <= not((inputs(161)) xor (inputs(228)));
    layer0_outputs(10433) <= (inputs(10)) or (inputs(20));
    layer0_outputs(10434) <= not(inputs(41));
    layer0_outputs(10435) <= not((inputs(9)) xor (inputs(204)));
    layer0_outputs(10436) <= not(inputs(209));
    layer0_outputs(10437) <= inputs(142);
    layer0_outputs(10438) <= not(inputs(220));
    layer0_outputs(10439) <= inputs(75);
    layer0_outputs(10440) <= inputs(130);
    layer0_outputs(10441) <= not(inputs(176));
    layer0_outputs(10442) <= not(inputs(220)) or (inputs(19));
    layer0_outputs(10443) <= not(inputs(114));
    layer0_outputs(10444) <= not(inputs(124)) or (inputs(220));
    layer0_outputs(10445) <= (inputs(213)) and (inputs(221));
    layer0_outputs(10446) <= (inputs(166)) xor (inputs(167));
    layer0_outputs(10447) <= not((inputs(147)) xor (inputs(158)));
    layer0_outputs(10448) <= (inputs(211)) and not (inputs(25));
    layer0_outputs(10449) <= inputs(181);
    layer0_outputs(10450) <= not((inputs(161)) or (inputs(68)));
    layer0_outputs(10451) <= not(inputs(211)) or (inputs(220));
    layer0_outputs(10452) <= inputs(40);
    layer0_outputs(10453) <= (inputs(194)) or (inputs(198));
    layer0_outputs(10454) <= (inputs(186)) or (inputs(227));
    layer0_outputs(10455) <= not(inputs(232)) or (inputs(189));
    layer0_outputs(10456) <= not(inputs(22));
    layer0_outputs(10457) <= inputs(72);
    layer0_outputs(10458) <= (inputs(164)) or (inputs(171));
    layer0_outputs(10459) <= (inputs(16)) xor (inputs(167));
    layer0_outputs(10460) <= '1';
    layer0_outputs(10461) <= inputs(131);
    layer0_outputs(10462) <= not((inputs(96)) xor (inputs(132)));
    layer0_outputs(10463) <= not((inputs(136)) xor (inputs(117)));
    layer0_outputs(10464) <= not(inputs(221)) or (inputs(212));
    layer0_outputs(10465) <= not((inputs(59)) or (inputs(76)));
    layer0_outputs(10466) <= (inputs(79)) or (inputs(36));
    layer0_outputs(10467) <= (inputs(202)) and not (inputs(103));
    layer0_outputs(10468) <= not((inputs(27)) or (inputs(67)));
    layer0_outputs(10469) <= inputs(230);
    layer0_outputs(10470) <= (inputs(204)) or (inputs(119));
    layer0_outputs(10471) <= inputs(247);
    layer0_outputs(10472) <= not((inputs(16)) or (inputs(154)));
    layer0_outputs(10473) <= inputs(236);
    layer0_outputs(10474) <= not((inputs(54)) xor (inputs(204)));
    layer0_outputs(10475) <= (inputs(164)) and not (inputs(62));
    layer0_outputs(10476) <= not(inputs(6));
    layer0_outputs(10477) <= (inputs(40)) and not (inputs(225));
    layer0_outputs(10478) <= (inputs(140)) or (inputs(34));
    layer0_outputs(10479) <= (inputs(5)) and (inputs(74));
    layer0_outputs(10480) <= (inputs(12)) or (inputs(18));
    layer0_outputs(10481) <= not((inputs(76)) or (inputs(6)));
    layer0_outputs(10482) <= not(inputs(97));
    layer0_outputs(10483) <= (inputs(39)) and not (inputs(80));
    layer0_outputs(10484) <= not((inputs(28)) and (inputs(114)));
    layer0_outputs(10485) <= not(inputs(54)) or (inputs(254));
    layer0_outputs(10486) <= inputs(39);
    layer0_outputs(10487) <= not(inputs(90));
    layer0_outputs(10488) <= (inputs(206)) xor (inputs(85));
    layer0_outputs(10489) <= '0';
    layer0_outputs(10490) <= (inputs(179)) or (inputs(183));
    layer0_outputs(10491) <= (inputs(41)) or (inputs(0));
    layer0_outputs(10492) <= not((inputs(101)) or (inputs(31)));
    layer0_outputs(10493) <= not((inputs(242)) xor (inputs(130)));
    layer0_outputs(10494) <= (inputs(32)) or (inputs(125));
    layer0_outputs(10495) <= not((inputs(212)) or (inputs(160)));
    layer0_outputs(10496) <= (inputs(25)) xor (inputs(240));
    layer0_outputs(10497) <= not((inputs(53)) or (inputs(83)));
    layer0_outputs(10498) <= (inputs(97)) or (inputs(134));
    layer0_outputs(10499) <= not(inputs(136));
    layer0_outputs(10500) <= inputs(237);
    layer0_outputs(10501) <= inputs(63);
    layer0_outputs(10502) <= inputs(130);
    layer0_outputs(10503) <= (inputs(174)) or (inputs(98));
    layer0_outputs(10504) <= (inputs(83)) or (inputs(77));
    layer0_outputs(10505) <= not((inputs(191)) xor (inputs(99)));
    layer0_outputs(10506) <= inputs(66);
    layer0_outputs(10507) <= (inputs(197)) and not (inputs(128));
    layer0_outputs(10508) <= (inputs(122)) and (inputs(107));
    layer0_outputs(10509) <= not(inputs(26));
    layer0_outputs(10510) <= (inputs(56)) xor (inputs(107));
    layer0_outputs(10511) <= not(inputs(98)) or (inputs(124));
    layer0_outputs(10512) <= not(inputs(90)) or (inputs(18));
    layer0_outputs(10513) <= (inputs(171)) or (inputs(79));
    layer0_outputs(10514) <= inputs(213);
    layer0_outputs(10515) <= (inputs(52)) and not (inputs(137));
    layer0_outputs(10516) <= (inputs(206)) or (inputs(174));
    layer0_outputs(10517) <= not((inputs(224)) or (inputs(78)));
    layer0_outputs(10518) <= not((inputs(21)) xor (inputs(73)));
    layer0_outputs(10519) <= '1';
    layer0_outputs(10520) <= not(inputs(57)) or (inputs(41));
    layer0_outputs(10521) <= not(inputs(251));
    layer0_outputs(10522) <= not((inputs(156)) xor (inputs(84)));
    layer0_outputs(10523) <= not(inputs(61));
    layer0_outputs(10524) <= (inputs(212)) or (inputs(240));
    layer0_outputs(10525) <= inputs(149);
    layer0_outputs(10526) <= not((inputs(33)) or (inputs(156)));
    layer0_outputs(10527) <= not((inputs(97)) or (inputs(69)));
    layer0_outputs(10528) <= inputs(166);
    layer0_outputs(10529) <= (inputs(167)) and not (inputs(222));
    layer0_outputs(10530) <= (inputs(194)) or (inputs(110));
    layer0_outputs(10531) <= (inputs(86)) xor (inputs(127));
    layer0_outputs(10532) <= not(inputs(56)) or (inputs(175));
    layer0_outputs(10533) <= (inputs(183)) and not (inputs(94));
    layer0_outputs(10534) <= not(inputs(93)) or (inputs(206));
    layer0_outputs(10535) <= (inputs(142)) or (inputs(128));
    layer0_outputs(10536) <= inputs(135);
    layer0_outputs(10537) <= inputs(35);
    layer0_outputs(10538) <= (inputs(177)) or (inputs(249));
    layer0_outputs(10539) <= not((inputs(61)) xor (inputs(71)));
    layer0_outputs(10540) <= '0';
    layer0_outputs(10541) <= not(inputs(102));
    layer0_outputs(10542) <= not(inputs(66)) or (inputs(209));
    layer0_outputs(10543) <= (inputs(176)) or (inputs(239));
    layer0_outputs(10544) <= not(inputs(136));
    layer0_outputs(10545) <= (inputs(68)) and not (inputs(2));
    layer0_outputs(10546) <= (inputs(247)) xor (inputs(215));
    layer0_outputs(10547) <= (inputs(40)) and (inputs(57));
    layer0_outputs(10548) <= not(inputs(194)) or (inputs(141));
    layer0_outputs(10549) <= not((inputs(2)) or (inputs(230)));
    layer0_outputs(10550) <= (inputs(198)) and not (inputs(100));
    layer0_outputs(10551) <= (inputs(113)) and not (inputs(13));
    layer0_outputs(10552) <= not(inputs(52)) or (inputs(205));
    layer0_outputs(10553) <= inputs(144);
    layer0_outputs(10554) <= (inputs(19)) or (inputs(16));
    layer0_outputs(10555) <= not((inputs(78)) xor (inputs(153)));
    layer0_outputs(10556) <= not(inputs(94)) or (inputs(153));
    layer0_outputs(10557) <= not(inputs(122)) or (inputs(164));
    layer0_outputs(10558) <= (inputs(253)) and not (inputs(155));
    layer0_outputs(10559) <= not(inputs(144)) or (inputs(95));
    layer0_outputs(10560) <= (inputs(32)) xor (inputs(241));
    layer0_outputs(10561) <= inputs(30);
    layer0_outputs(10562) <= not(inputs(192));
    layer0_outputs(10563) <= inputs(218);
    layer0_outputs(10564) <= not(inputs(14));
    layer0_outputs(10565) <= inputs(25);
    layer0_outputs(10566) <= '1';
    layer0_outputs(10567) <= '0';
    layer0_outputs(10568) <= not(inputs(154));
    layer0_outputs(10569) <= not((inputs(116)) xor (inputs(3)));
    layer0_outputs(10570) <= (inputs(115)) and not (inputs(249));
    layer0_outputs(10571) <= (inputs(41)) or (inputs(19));
    layer0_outputs(10572) <= not(inputs(118));
    layer0_outputs(10573) <= (inputs(36)) or (inputs(192));
    layer0_outputs(10574) <= not(inputs(165));
    layer0_outputs(10575) <= (inputs(233)) and not (inputs(4));
    layer0_outputs(10576) <= (inputs(183)) xor (inputs(147));
    layer0_outputs(10577) <= not(inputs(160));
    layer0_outputs(10578) <= inputs(179);
    layer0_outputs(10579) <= (inputs(88)) and not (inputs(88));
    layer0_outputs(10580) <= not(inputs(76)) or (inputs(224));
    layer0_outputs(10581) <= inputs(195);
    layer0_outputs(10582) <= (inputs(235)) or (inputs(161));
    layer0_outputs(10583) <= not(inputs(49));
    layer0_outputs(10584) <= (inputs(102)) and not (inputs(41));
    layer0_outputs(10585) <= not((inputs(113)) or (inputs(248)));
    layer0_outputs(10586) <= (inputs(69)) and not (inputs(179));
    layer0_outputs(10587) <= not(inputs(99));
    layer0_outputs(10588) <= (inputs(45)) or (inputs(206));
    layer0_outputs(10589) <= inputs(104);
    layer0_outputs(10590) <= not((inputs(97)) or (inputs(177)));
    layer0_outputs(10591) <= inputs(100);
    layer0_outputs(10592) <= not((inputs(218)) or (inputs(109)));
    layer0_outputs(10593) <= '1';
    layer0_outputs(10594) <= not(inputs(41));
    layer0_outputs(10595) <= inputs(75);
    layer0_outputs(10596) <= not((inputs(25)) and (inputs(27)));
    layer0_outputs(10597) <= not(inputs(233));
    layer0_outputs(10598) <= inputs(140);
    layer0_outputs(10599) <= not((inputs(51)) or (inputs(22)));
    layer0_outputs(10600) <= not((inputs(23)) or (inputs(37)));
    layer0_outputs(10601) <= inputs(97);
    layer0_outputs(10602) <= (inputs(186)) or (inputs(100));
    layer0_outputs(10603) <= (inputs(140)) xor (inputs(171));
    layer0_outputs(10604) <= (inputs(12)) or (inputs(34));
    layer0_outputs(10605) <= not((inputs(227)) or (inputs(207)));
    layer0_outputs(10606) <= not(inputs(100));
    layer0_outputs(10607) <= (inputs(157)) and not (inputs(7));
    layer0_outputs(10608) <= not(inputs(178));
    layer0_outputs(10609) <= (inputs(23)) or (inputs(145));
    layer0_outputs(10610) <= inputs(90);
    layer0_outputs(10611) <= not(inputs(91)) or (inputs(50));
    layer0_outputs(10612) <= inputs(215);
    layer0_outputs(10613) <= not(inputs(215));
    layer0_outputs(10614) <= not((inputs(196)) or (inputs(107)));
    layer0_outputs(10615) <= not(inputs(204)) or (inputs(31));
    layer0_outputs(10616) <= (inputs(168)) and not (inputs(27));
    layer0_outputs(10617) <= not((inputs(209)) or (inputs(35)));
    layer0_outputs(10618) <= inputs(126);
    layer0_outputs(10619) <= not(inputs(162));
    layer0_outputs(10620) <= not(inputs(228));
    layer0_outputs(10621) <= not((inputs(123)) and (inputs(68)));
    layer0_outputs(10622) <= (inputs(169)) and not (inputs(77));
    layer0_outputs(10623) <= (inputs(254)) or (inputs(113));
    layer0_outputs(10624) <= not(inputs(216));
    layer0_outputs(10625) <= not(inputs(200));
    layer0_outputs(10626) <= (inputs(204)) or (inputs(239));
    layer0_outputs(10627) <= not(inputs(234));
    layer0_outputs(10628) <= not(inputs(99));
    layer0_outputs(10629) <= inputs(4);
    layer0_outputs(10630) <= (inputs(120)) xor (inputs(91));
    layer0_outputs(10631) <= inputs(42);
    layer0_outputs(10632) <= (inputs(190)) and not (inputs(31));
    layer0_outputs(10633) <= (inputs(97)) xor (inputs(34));
    layer0_outputs(10634) <= not(inputs(103)) or (inputs(14));
    layer0_outputs(10635) <= inputs(183);
    layer0_outputs(10636) <= (inputs(82)) or (inputs(220));
    layer0_outputs(10637) <= not(inputs(17));
    layer0_outputs(10638) <= inputs(113);
    layer0_outputs(10639) <= (inputs(225)) or (inputs(212));
    layer0_outputs(10640) <= (inputs(38)) xor (inputs(10));
    layer0_outputs(10641) <= not((inputs(44)) or (inputs(36)));
    layer0_outputs(10642) <= (inputs(70)) xor (inputs(228));
    layer0_outputs(10643) <= (inputs(65)) or (inputs(76));
    layer0_outputs(10644) <= (inputs(255)) or (inputs(222));
    layer0_outputs(10645) <= not((inputs(183)) or (inputs(254)));
    layer0_outputs(10646) <= (inputs(206)) or (inputs(139));
    layer0_outputs(10647) <= (inputs(128)) and not (inputs(136));
    layer0_outputs(10648) <= not(inputs(89));
    layer0_outputs(10649) <= not(inputs(109)) or (inputs(193));
    layer0_outputs(10650) <= '0';
    layer0_outputs(10651) <= not((inputs(85)) or (inputs(217)));
    layer0_outputs(10652) <= inputs(157);
    layer0_outputs(10653) <= not((inputs(115)) xor (inputs(202)));
    layer0_outputs(10654) <= not(inputs(119));
    layer0_outputs(10655) <= not(inputs(186));
    layer0_outputs(10656) <= not(inputs(3)) or (inputs(145));
    layer0_outputs(10657) <= not((inputs(178)) or (inputs(7)));
    layer0_outputs(10658) <= not(inputs(219));
    layer0_outputs(10659) <= (inputs(130)) and not (inputs(49));
    layer0_outputs(10660) <= (inputs(7)) and not (inputs(131));
    layer0_outputs(10661) <= not((inputs(145)) and (inputs(218)));
    layer0_outputs(10662) <= (inputs(46)) xor (inputs(77));
    layer0_outputs(10663) <= inputs(213);
    layer0_outputs(10664) <= not(inputs(149));
    layer0_outputs(10665) <= (inputs(18)) or (inputs(117));
    layer0_outputs(10666) <= inputs(48);
    layer0_outputs(10667) <= (inputs(9)) and not (inputs(190));
    layer0_outputs(10668) <= (inputs(93)) and not (inputs(51));
    layer0_outputs(10669) <= inputs(37);
    layer0_outputs(10670) <= not((inputs(194)) or (inputs(187)));
    layer0_outputs(10671) <= inputs(239);
    layer0_outputs(10672) <= (inputs(184)) and not (inputs(69));
    layer0_outputs(10673) <= '1';
    layer0_outputs(10674) <= inputs(92);
    layer0_outputs(10675) <= (inputs(64)) and not (inputs(208));
    layer0_outputs(10676) <= (inputs(119)) and not (inputs(210));
    layer0_outputs(10677) <= inputs(90);
    layer0_outputs(10678) <= inputs(102);
    layer0_outputs(10679) <= inputs(162);
    layer0_outputs(10680) <= not(inputs(21)) or (inputs(30));
    layer0_outputs(10681) <= not(inputs(0)) or (inputs(127));
    layer0_outputs(10682) <= not(inputs(238)) or (inputs(250));
    layer0_outputs(10683) <= not(inputs(84));
    layer0_outputs(10684) <= (inputs(199)) and not (inputs(66));
    layer0_outputs(10685) <= (inputs(162)) and (inputs(135));
    layer0_outputs(10686) <= (inputs(26)) xor (inputs(42));
    layer0_outputs(10687) <= not((inputs(179)) and (inputs(147)));
    layer0_outputs(10688) <= (inputs(171)) or (inputs(216));
    layer0_outputs(10689) <= (inputs(115)) or (inputs(254));
    layer0_outputs(10690) <= not(inputs(132));
    layer0_outputs(10691) <= (inputs(174)) or (inputs(207));
    layer0_outputs(10692) <= inputs(40);
    layer0_outputs(10693) <= not(inputs(35));
    layer0_outputs(10694) <= not((inputs(210)) or (inputs(102)));
    layer0_outputs(10695) <= (inputs(80)) or (inputs(64));
    layer0_outputs(10696) <= (inputs(75)) or (inputs(43));
    layer0_outputs(10697) <= '0';
    layer0_outputs(10698) <= not(inputs(81));
    layer0_outputs(10699) <= not((inputs(91)) xor (inputs(32)));
    layer0_outputs(10700) <= not((inputs(50)) or (inputs(35)));
    layer0_outputs(10701) <= inputs(180);
    layer0_outputs(10702) <= not((inputs(184)) and (inputs(145)));
    layer0_outputs(10703) <= (inputs(114)) and not (inputs(11));
    layer0_outputs(10704) <= (inputs(119)) and not (inputs(226));
    layer0_outputs(10705) <= not((inputs(95)) xor (inputs(64)));
    layer0_outputs(10706) <= not(inputs(76)) or (inputs(112));
    layer0_outputs(10707) <= not((inputs(157)) and (inputs(1)));
    layer0_outputs(10708) <= '0';
    layer0_outputs(10709) <= inputs(160);
    layer0_outputs(10710) <= (inputs(238)) and not (inputs(141));
    layer0_outputs(10711) <= inputs(114);
    layer0_outputs(10712) <= not(inputs(125));
    layer0_outputs(10713) <= not(inputs(126));
    layer0_outputs(10714) <= not((inputs(253)) xor (inputs(51)));
    layer0_outputs(10715) <= (inputs(238)) and not (inputs(80));
    layer0_outputs(10716) <= not(inputs(195)) or (inputs(27));
    layer0_outputs(10717) <= not(inputs(17)) or (inputs(190));
    layer0_outputs(10718) <= not(inputs(22));
    layer0_outputs(10719) <= (inputs(211)) or (inputs(9));
    layer0_outputs(10720) <= inputs(31);
    layer0_outputs(10721) <= inputs(123);
    layer0_outputs(10722) <= not((inputs(2)) and (inputs(134)));
    layer0_outputs(10723) <= not(inputs(72));
    layer0_outputs(10724) <= not(inputs(197));
    layer0_outputs(10725) <= not(inputs(104));
    layer0_outputs(10726) <= (inputs(17)) or (inputs(25));
    layer0_outputs(10727) <= not(inputs(99)) or (inputs(210));
    layer0_outputs(10728) <= inputs(50);
    layer0_outputs(10729) <= (inputs(166)) and not (inputs(109));
    layer0_outputs(10730) <= (inputs(22)) and not (inputs(198));
    layer0_outputs(10731) <= not((inputs(152)) xor (inputs(149)));
    layer0_outputs(10732) <= inputs(232);
    layer0_outputs(10733) <= inputs(178);
    layer0_outputs(10734) <= not(inputs(101));
    layer0_outputs(10735) <= not((inputs(113)) and (inputs(107)));
    layer0_outputs(10736) <= inputs(184);
    layer0_outputs(10737) <= not(inputs(158));
    layer0_outputs(10738) <= (inputs(6)) xor (inputs(64));
    layer0_outputs(10739) <= inputs(144);
    layer0_outputs(10740) <= (inputs(162)) or (inputs(150));
    layer0_outputs(10741) <= not((inputs(47)) xor (inputs(222)));
    layer0_outputs(10742) <= not((inputs(209)) xor (inputs(246)));
    layer0_outputs(10743) <= (inputs(11)) xor (inputs(111));
    layer0_outputs(10744) <= not((inputs(30)) and (inputs(99)));
    layer0_outputs(10745) <= not((inputs(74)) xor (inputs(1)));
    layer0_outputs(10746) <= not(inputs(74));
    layer0_outputs(10747) <= not(inputs(191));
    layer0_outputs(10748) <= (inputs(104)) and not (inputs(48));
    layer0_outputs(10749) <= not((inputs(48)) xor (inputs(29)));
    layer0_outputs(10750) <= not((inputs(23)) or (inputs(186)));
    layer0_outputs(10751) <= not(inputs(247)) or (inputs(42));
    layer0_outputs(10752) <= not(inputs(200));
    layer0_outputs(10753) <= (inputs(124)) and not (inputs(158));
    layer0_outputs(10754) <= not((inputs(20)) or (inputs(21)));
    layer0_outputs(10755) <= not(inputs(180));
    layer0_outputs(10756) <= not((inputs(123)) or (inputs(66)));
    layer0_outputs(10757) <= not(inputs(72));
    layer0_outputs(10758) <= '0';
    layer0_outputs(10759) <= inputs(201);
    layer0_outputs(10760) <= not((inputs(116)) xor (inputs(226)));
    layer0_outputs(10761) <= not(inputs(165)) or (inputs(80));
    layer0_outputs(10762) <= not(inputs(220));
    layer0_outputs(10763) <= not(inputs(71));
    layer0_outputs(10764) <= not((inputs(72)) and (inputs(191)));
    layer0_outputs(10765) <= not((inputs(238)) or (inputs(34)));
    layer0_outputs(10766) <= not(inputs(137)) or (inputs(26));
    layer0_outputs(10767) <= (inputs(252)) and not (inputs(112));
    layer0_outputs(10768) <= inputs(220);
    layer0_outputs(10769) <= not((inputs(46)) or (inputs(140)));
    layer0_outputs(10770) <= not((inputs(66)) and (inputs(45)));
    layer0_outputs(10771) <= not(inputs(45)) or (inputs(221));
    layer0_outputs(10772) <= (inputs(175)) and not (inputs(254));
    layer0_outputs(10773) <= not(inputs(218));
    layer0_outputs(10774) <= (inputs(73)) or (inputs(225));
    layer0_outputs(10775) <= not(inputs(222));
    layer0_outputs(10776) <= (inputs(208)) or (inputs(224));
    layer0_outputs(10777) <= inputs(101);
    layer0_outputs(10778) <= not((inputs(149)) xor (inputs(231)));
    layer0_outputs(10779) <= (inputs(204)) and not (inputs(142));
    layer0_outputs(10780) <= (inputs(164)) xor (inputs(167));
    layer0_outputs(10781) <= inputs(86);
    layer0_outputs(10782) <= not(inputs(127));
    layer0_outputs(10783) <= not((inputs(228)) or (inputs(84)));
    layer0_outputs(10784) <= inputs(196);
    layer0_outputs(10785) <= '1';
    layer0_outputs(10786) <= (inputs(120)) xor (inputs(28));
    layer0_outputs(10787) <= not(inputs(233)) or (inputs(125));
    layer0_outputs(10788) <= not(inputs(137)) or (inputs(211));
    layer0_outputs(10789) <= inputs(39);
    layer0_outputs(10790) <= not(inputs(25)) or (inputs(200));
    layer0_outputs(10791) <= not(inputs(200));
    layer0_outputs(10792) <= not(inputs(94));
    layer0_outputs(10793) <= inputs(212);
    layer0_outputs(10794) <= not((inputs(59)) xor (inputs(196)));
    layer0_outputs(10795) <= inputs(102);
    layer0_outputs(10796) <= (inputs(63)) or (inputs(214));
    layer0_outputs(10797) <= not((inputs(228)) or (inputs(39)));
    layer0_outputs(10798) <= (inputs(244)) xor (inputs(199));
    layer0_outputs(10799) <= not((inputs(192)) and (inputs(137)));
    layer0_outputs(10800) <= not((inputs(19)) or (inputs(144)));
    layer0_outputs(10801) <= inputs(122);
    layer0_outputs(10802) <= (inputs(226)) or (inputs(87));
    layer0_outputs(10803) <= not(inputs(207));
    layer0_outputs(10804) <= (inputs(170)) and not (inputs(235));
    layer0_outputs(10805) <= not(inputs(148));
    layer0_outputs(10806) <= (inputs(65)) or (inputs(251));
    layer0_outputs(10807) <= (inputs(194)) and not (inputs(93));
    layer0_outputs(10808) <= (inputs(91)) and not (inputs(211));
    layer0_outputs(10809) <= not(inputs(185)) or (inputs(0));
    layer0_outputs(10810) <= not(inputs(65));
    layer0_outputs(10811) <= not((inputs(186)) or (inputs(157)));
    layer0_outputs(10812) <= not(inputs(35)) or (inputs(47));
    layer0_outputs(10813) <= inputs(78);
    layer0_outputs(10814) <= (inputs(255)) or (inputs(113));
    layer0_outputs(10815) <= inputs(12);
    layer0_outputs(10816) <= inputs(59);
    layer0_outputs(10817) <= not((inputs(106)) or (inputs(248)));
    layer0_outputs(10818) <= '0';
    layer0_outputs(10819) <= inputs(54);
    layer0_outputs(10820) <= not((inputs(112)) or (inputs(249)));
    layer0_outputs(10821) <= (inputs(17)) xor (inputs(157));
    layer0_outputs(10822) <= (inputs(103)) xor (inputs(143));
    layer0_outputs(10823) <= inputs(58);
    layer0_outputs(10824) <= not((inputs(220)) or (inputs(81)));
    layer0_outputs(10825) <= (inputs(164)) xor (inputs(68));
    layer0_outputs(10826) <= not((inputs(143)) or (inputs(41)));
    layer0_outputs(10827) <= not((inputs(106)) xor (inputs(141)));
    layer0_outputs(10828) <= '1';
    layer0_outputs(10829) <= (inputs(42)) and (inputs(96));
    layer0_outputs(10830) <= not(inputs(232));
    layer0_outputs(10831) <= not((inputs(105)) xor (inputs(165)));
    layer0_outputs(10832) <= inputs(90);
    layer0_outputs(10833) <= (inputs(14)) or (inputs(107));
    layer0_outputs(10834) <= not((inputs(171)) xor (inputs(119)));
    layer0_outputs(10835) <= inputs(108);
    layer0_outputs(10836) <= not((inputs(251)) or (inputs(104)));
    layer0_outputs(10837) <= inputs(129);
    layer0_outputs(10838) <= (inputs(192)) xor (inputs(179));
    layer0_outputs(10839) <= not(inputs(185)) or (inputs(107));
    layer0_outputs(10840) <= not(inputs(139)) or (inputs(253));
    layer0_outputs(10841) <= not(inputs(11));
    layer0_outputs(10842) <= not(inputs(111));
    layer0_outputs(10843) <= inputs(107);
    layer0_outputs(10844) <= not(inputs(233));
    layer0_outputs(10845) <= not(inputs(236));
    layer0_outputs(10846) <= not(inputs(231));
    layer0_outputs(10847) <= not(inputs(254));
    layer0_outputs(10848) <= not(inputs(228)) or (inputs(40));
    layer0_outputs(10849) <= not(inputs(214));
    layer0_outputs(10850) <= (inputs(205)) and not (inputs(15));
    layer0_outputs(10851) <= (inputs(91)) and not (inputs(158));
    layer0_outputs(10852) <= inputs(90);
    layer0_outputs(10853) <= (inputs(196)) and not (inputs(145));
    layer0_outputs(10854) <= (inputs(52)) and not (inputs(33));
    layer0_outputs(10855) <= not(inputs(154));
    layer0_outputs(10856) <= not((inputs(59)) xor (inputs(17)));
    layer0_outputs(10857) <= (inputs(231)) and not (inputs(128));
    layer0_outputs(10858) <= (inputs(253)) and not (inputs(224));
    layer0_outputs(10859) <= not(inputs(244)) or (inputs(104));
    layer0_outputs(10860) <= not((inputs(133)) or (inputs(133)));
    layer0_outputs(10861) <= not((inputs(244)) or (inputs(156)));
    layer0_outputs(10862) <= not(inputs(69));
    layer0_outputs(10863) <= not(inputs(75));
    layer0_outputs(10864) <= not((inputs(27)) xor (inputs(90)));
    layer0_outputs(10865) <= (inputs(24)) and not (inputs(229));
    layer0_outputs(10866) <= not((inputs(110)) or (inputs(222)));
    layer0_outputs(10867) <= not(inputs(96));
    layer0_outputs(10868) <= '1';
    layer0_outputs(10869) <= (inputs(151)) and not (inputs(245));
    layer0_outputs(10870) <= not(inputs(12));
    layer0_outputs(10871) <= inputs(148);
    layer0_outputs(10872) <= (inputs(109)) or (inputs(52));
    layer0_outputs(10873) <= (inputs(70)) or (inputs(210));
    layer0_outputs(10874) <= not((inputs(232)) xor (inputs(38)));
    layer0_outputs(10875) <= (inputs(66)) xor (inputs(187));
    layer0_outputs(10876) <= not(inputs(25));
    layer0_outputs(10877) <= inputs(212);
    layer0_outputs(10878) <= (inputs(191)) or (inputs(248));
    layer0_outputs(10879) <= not((inputs(230)) xor (inputs(232)));
    layer0_outputs(10880) <= (inputs(137)) xor (inputs(210));
    layer0_outputs(10881) <= not(inputs(125)) or (inputs(136));
    layer0_outputs(10882) <= not((inputs(65)) xor (inputs(115)));
    layer0_outputs(10883) <= inputs(18);
    layer0_outputs(10884) <= not(inputs(22)) or (inputs(206));
    layer0_outputs(10885) <= inputs(201);
    layer0_outputs(10886) <= not((inputs(9)) xor (inputs(117)));
    layer0_outputs(10887) <= not(inputs(62));
    layer0_outputs(10888) <= (inputs(9)) xor (inputs(27));
    layer0_outputs(10889) <= (inputs(10)) and not (inputs(113));
    layer0_outputs(10890) <= not(inputs(233));
    layer0_outputs(10891) <= (inputs(89)) xor (inputs(88));
    layer0_outputs(10892) <= not((inputs(253)) or (inputs(119)));
    layer0_outputs(10893) <= inputs(145);
    layer0_outputs(10894) <= not(inputs(78));
    layer0_outputs(10895) <= (inputs(94)) or (inputs(250));
    layer0_outputs(10896) <= not(inputs(76));
    layer0_outputs(10897) <= not((inputs(223)) or (inputs(173)));
    layer0_outputs(10898) <= (inputs(48)) or (inputs(176));
    layer0_outputs(10899) <= not((inputs(216)) xor (inputs(201)));
    layer0_outputs(10900) <= (inputs(130)) xor (inputs(120));
    layer0_outputs(10901) <= (inputs(213)) or (inputs(105));
    layer0_outputs(10902) <= (inputs(138)) xor (inputs(48));
    layer0_outputs(10903) <= not(inputs(123));
    layer0_outputs(10904) <= not((inputs(50)) or (inputs(122)));
    layer0_outputs(10905) <= inputs(117);
    layer0_outputs(10906) <= not((inputs(236)) or (inputs(84)));
    layer0_outputs(10907) <= not((inputs(226)) xor (inputs(130)));
    layer0_outputs(10908) <= not((inputs(148)) xor (inputs(33)));
    layer0_outputs(10909) <= not((inputs(131)) or (inputs(45)));
    layer0_outputs(10910) <= not((inputs(52)) and (inputs(117)));
    layer0_outputs(10911) <= (inputs(44)) xor (inputs(60));
    layer0_outputs(10912) <= not(inputs(198)) or (inputs(172));
    layer0_outputs(10913) <= inputs(215);
    layer0_outputs(10914) <= inputs(165);
    layer0_outputs(10915) <= (inputs(36)) xor (inputs(75));
    layer0_outputs(10916) <= (inputs(213)) xor (inputs(144));
    layer0_outputs(10917) <= not(inputs(170));
    layer0_outputs(10918) <= not((inputs(138)) xor (inputs(10)));
    layer0_outputs(10919) <= (inputs(85)) and (inputs(52));
    layer0_outputs(10920) <= inputs(59);
    layer0_outputs(10921) <= inputs(149);
    layer0_outputs(10922) <= not(inputs(121)) or (inputs(188));
    layer0_outputs(10923) <= not(inputs(24)) or (inputs(52));
    layer0_outputs(10924) <= inputs(47);
    layer0_outputs(10925) <= (inputs(150)) or (inputs(215));
    layer0_outputs(10926) <= inputs(87);
    layer0_outputs(10927) <= (inputs(32)) xor (inputs(199));
    layer0_outputs(10928) <= (inputs(187)) or (inputs(131));
    layer0_outputs(10929) <= inputs(226);
    layer0_outputs(10930) <= (inputs(249)) and not (inputs(243));
    layer0_outputs(10931) <= not((inputs(222)) or (inputs(80)));
    layer0_outputs(10932) <= (inputs(124)) and not (inputs(29));
    layer0_outputs(10933) <= (inputs(43)) and not (inputs(213));
    layer0_outputs(10934) <= not((inputs(112)) xor (inputs(106)));
    layer0_outputs(10935) <= not((inputs(18)) or (inputs(69)));
    layer0_outputs(10936) <= inputs(83);
    layer0_outputs(10937) <= (inputs(3)) or (inputs(111));
    layer0_outputs(10938) <= (inputs(152)) xor (inputs(1));
    layer0_outputs(10939) <= inputs(85);
    layer0_outputs(10940) <= not(inputs(181));
    layer0_outputs(10941) <= not(inputs(205)) or (inputs(207));
    layer0_outputs(10942) <= '1';
    layer0_outputs(10943) <= not(inputs(42));
    layer0_outputs(10944) <= not(inputs(138));
    layer0_outputs(10945) <= not((inputs(207)) or (inputs(109)));
    layer0_outputs(10946) <= not((inputs(226)) or (inputs(164)));
    layer0_outputs(10947) <= (inputs(112)) or (inputs(87));
    layer0_outputs(10948) <= inputs(241);
    layer0_outputs(10949) <= inputs(10);
    layer0_outputs(10950) <= not(inputs(187)) or (inputs(95));
    layer0_outputs(10951) <= not(inputs(77)) or (inputs(77));
    layer0_outputs(10952) <= not(inputs(164));
    layer0_outputs(10953) <= (inputs(199)) and not (inputs(201));
    layer0_outputs(10954) <= not(inputs(90));
    layer0_outputs(10955) <= inputs(107);
    layer0_outputs(10956) <= not(inputs(233));
    layer0_outputs(10957) <= not((inputs(37)) or (inputs(7)));
    layer0_outputs(10958) <= inputs(86);
    layer0_outputs(10959) <= not((inputs(190)) xor (inputs(19)));
    layer0_outputs(10960) <= inputs(26);
    layer0_outputs(10961) <= not(inputs(9)) or (inputs(240));
    layer0_outputs(10962) <= not((inputs(123)) xor (inputs(103)));
    layer0_outputs(10963) <= not((inputs(3)) xor (inputs(91)));
    layer0_outputs(10964) <= inputs(85);
    layer0_outputs(10965) <= not((inputs(1)) xor (inputs(71)));
    layer0_outputs(10966) <= not((inputs(215)) xor (inputs(231)));
    layer0_outputs(10967) <= inputs(220);
    layer0_outputs(10968) <= (inputs(8)) or (inputs(189));
    layer0_outputs(10969) <= not((inputs(18)) or (inputs(90)));
    layer0_outputs(10970) <= (inputs(231)) and not (inputs(147));
    layer0_outputs(10971) <= (inputs(156)) and not (inputs(4));
    layer0_outputs(10972) <= not(inputs(101));
    layer0_outputs(10973) <= (inputs(5)) and (inputs(26));
    layer0_outputs(10974) <= not((inputs(215)) xor (inputs(202)));
    layer0_outputs(10975) <= (inputs(14)) xor (inputs(239));
    layer0_outputs(10976) <= not((inputs(63)) or (inputs(246)));
    layer0_outputs(10977) <= not(inputs(47)) or (inputs(222));
    layer0_outputs(10978) <= '1';
    layer0_outputs(10979) <= not(inputs(212));
    layer0_outputs(10980) <= inputs(108);
    layer0_outputs(10981) <= inputs(188);
    layer0_outputs(10982) <= (inputs(138)) xor (inputs(21));
    layer0_outputs(10983) <= (inputs(211)) and not (inputs(137));
    layer0_outputs(10984) <= not(inputs(207)) or (inputs(158));
    layer0_outputs(10985) <= (inputs(208)) xor (inputs(206));
    layer0_outputs(10986) <= (inputs(29)) and not (inputs(137));
    layer0_outputs(10987) <= not(inputs(162));
    layer0_outputs(10988) <= not(inputs(214)) or (inputs(73));
    layer0_outputs(10989) <= '0';
    layer0_outputs(10990) <= not((inputs(199)) or (inputs(242)));
    layer0_outputs(10991) <= (inputs(181)) and not (inputs(45));
    layer0_outputs(10992) <= inputs(119);
    layer0_outputs(10993) <= inputs(23);
    layer0_outputs(10994) <= inputs(24);
    layer0_outputs(10995) <= (inputs(247)) and not (inputs(107));
    layer0_outputs(10996) <= not((inputs(9)) xor (inputs(117)));
    layer0_outputs(10997) <= inputs(154);
    layer0_outputs(10998) <= not(inputs(150));
    layer0_outputs(10999) <= not(inputs(179)) or (inputs(43));
    layer0_outputs(11000) <= not((inputs(142)) or (inputs(108)));
    layer0_outputs(11001) <= (inputs(45)) and not (inputs(33));
    layer0_outputs(11002) <= inputs(25);
    layer0_outputs(11003) <= (inputs(54)) xor (inputs(8));
    layer0_outputs(11004) <= (inputs(216)) and not (inputs(130));
    layer0_outputs(11005) <= not(inputs(12));
    layer0_outputs(11006) <= not(inputs(102));
    layer0_outputs(11007) <= not(inputs(248)) or (inputs(57));
    layer0_outputs(11008) <= inputs(187);
    layer0_outputs(11009) <= (inputs(165)) and not (inputs(208));
    layer0_outputs(11010) <= (inputs(6)) and not (inputs(251));
    layer0_outputs(11011) <= not(inputs(244)) or (inputs(97));
    layer0_outputs(11012) <= not((inputs(191)) xor (inputs(163)));
    layer0_outputs(11013) <= inputs(126);
    layer0_outputs(11014) <= (inputs(81)) or (inputs(235));
    layer0_outputs(11015) <= not(inputs(232)) or (inputs(40));
    layer0_outputs(11016) <= (inputs(71)) and not (inputs(112));
    layer0_outputs(11017) <= (inputs(229)) and (inputs(171));
    layer0_outputs(11018) <= inputs(170);
    layer0_outputs(11019) <= not(inputs(196)) or (inputs(97));
    layer0_outputs(11020) <= inputs(108);
    layer0_outputs(11021) <= inputs(214);
    layer0_outputs(11022) <= (inputs(165)) and not (inputs(60));
    layer0_outputs(11023) <= (inputs(161)) xor (inputs(207));
    layer0_outputs(11024) <= not((inputs(43)) and (inputs(25)));
    layer0_outputs(11025) <= (inputs(88)) and not (inputs(235));
    layer0_outputs(11026) <= inputs(94);
    layer0_outputs(11027) <= not(inputs(23)) or (inputs(114));
    layer0_outputs(11028) <= inputs(31);
    layer0_outputs(11029) <= inputs(88);
    layer0_outputs(11030) <= inputs(182);
    layer0_outputs(11031) <= (inputs(17)) or (inputs(181));
    layer0_outputs(11032) <= (inputs(46)) xor (inputs(103));
    layer0_outputs(11033) <= (inputs(7)) or (inputs(243));
    layer0_outputs(11034) <= not(inputs(162));
    layer0_outputs(11035) <= inputs(232);
    layer0_outputs(11036) <= not(inputs(75));
    layer0_outputs(11037) <= (inputs(157)) xor (inputs(123));
    layer0_outputs(11038) <= '1';
    layer0_outputs(11039) <= (inputs(23)) xor (inputs(192));
    layer0_outputs(11040) <= (inputs(142)) xor (inputs(45));
    layer0_outputs(11041) <= inputs(142);
    layer0_outputs(11042) <= not(inputs(227)) or (inputs(74));
    layer0_outputs(11043) <= not(inputs(98));
    layer0_outputs(11044) <= inputs(246);
    layer0_outputs(11045) <= not((inputs(152)) xor (inputs(183)));
    layer0_outputs(11046) <= inputs(149);
    layer0_outputs(11047) <= not(inputs(136));
    layer0_outputs(11048) <= not(inputs(75));
    layer0_outputs(11049) <= inputs(192);
    layer0_outputs(11050) <= (inputs(202)) and not (inputs(241));
    layer0_outputs(11051) <= inputs(59);
    layer0_outputs(11052) <= not((inputs(191)) or (inputs(156)));
    layer0_outputs(11053) <= not((inputs(195)) or (inputs(20)));
    layer0_outputs(11054) <= (inputs(190)) or (inputs(244));
    layer0_outputs(11055) <= not(inputs(114));
    layer0_outputs(11056) <= not(inputs(162));
    layer0_outputs(11057) <= inputs(141);
    layer0_outputs(11058) <= not((inputs(171)) or (inputs(156)));
    layer0_outputs(11059) <= (inputs(138)) or (inputs(235));
    layer0_outputs(11060) <= not(inputs(174));
    layer0_outputs(11061) <= (inputs(239)) and (inputs(13));
    layer0_outputs(11062) <= not(inputs(182));
    layer0_outputs(11063) <= (inputs(6)) and not (inputs(216));
    layer0_outputs(11064) <= (inputs(180)) and not (inputs(175));
    layer0_outputs(11065) <= not(inputs(131));
    layer0_outputs(11066) <= not((inputs(220)) or (inputs(130)));
    layer0_outputs(11067) <= not(inputs(98)) or (inputs(192));
    layer0_outputs(11068) <= inputs(73);
    layer0_outputs(11069) <= (inputs(144)) and (inputs(244));
    layer0_outputs(11070) <= inputs(189);
    layer0_outputs(11071) <= inputs(133);
    layer0_outputs(11072) <= not(inputs(198));
    layer0_outputs(11073) <= not(inputs(180)) or (inputs(45));
    layer0_outputs(11074) <= not(inputs(218)) or (inputs(123));
    layer0_outputs(11075) <= (inputs(232)) and not (inputs(130));
    layer0_outputs(11076) <= not(inputs(133));
    layer0_outputs(11077) <= not((inputs(208)) or (inputs(41)));
    layer0_outputs(11078) <= (inputs(137)) or (inputs(76));
    layer0_outputs(11079) <= (inputs(12)) xor (inputs(134));
    layer0_outputs(11080) <= (inputs(193)) or (inputs(17));
    layer0_outputs(11081) <= not(inputs(11));
    layer0_outputs(11082) <= inputs(197);
    layer0_outputs(11083) <= (inputs(9)) xor (inputs(221));
    layer0_outputs(11084) <= not(inputs(157));
    layer0_outputs(11085) <= (inputs(97)) xor (inputs(84));
    layer0_outputs(11086) <= not(inputs(187)) or (inputs(116));
    layer0_outputs(11087) <= (inputs(167)) xor (inputs(133));
    layer0_outputs(11088) <= (inputs(226)) and (inputs(113));
    layer0_outputs(11089) <= not(inputs(74)) or (inputs(197));
    layer0_outputs(11090) <= not((inputs(244)) or (inputs(108)));
    layer0_outputs(11091) <= (inputs(129)) xor (inputs(54));
    layer0_outputs(11092) <= not((inputs(27)) or (inputs(246)));
    layer0_outputs(11093) <= inputs(131);
    layer0_outputs(11094) <= (inputs(184)) or (inputs(170));
    layer0_outputs(11095) <= not((inputs(49)) xor (inputs(176)));
    layer0_outputs(11096) <= inputs(230);
    layer0_outputs(11097) <= not(inputs(215));
    layer0_outputs(11098) <= (inputs(96)) or (inputs(9));
    layer0_outputs(11099) <= not(inputs(161)) or (inputs(103));
    layer0_outputs(11100) <= inputs(195);
    layer0_outputs(11101) <= not(inputs(222)) or (inputs(125));
    layer0_outputs(11102) <= (inputs(4)) and (inputs(206));
    layer0_outputs(11103) <= inputs(133);
    layer0_outputs(11104) <= (inputs(235)) or (inputs(169));
    layer0_outputs(11105) <= inputs(89);
    layer0_outputs(11106) <= (inputs(239)) or (inputs(196));
    layer0_outputs(11107) <= not((inputs(82)) or (inputs(17)));
    layer0_outputs(11108) <= (inputs(39)) and not (inputs(178));
    layer0_outputs(11109) <= not(inputs(52)) or (inputs(169));
    layer0_outputs(11110) <= (inputs(95)) or (inputs(39));
    layer0_outputs(11111) <= not(inputs(189)) or (inputs(155));
    layer0_outputs(11112) <= inputs(65);
    layer0_outputs(11113) <= (inputs(81)) and not (inputs(198));
    layer0_outputs(11114) <= (inputs(140)) xor (inputs(24));
    layer0_outputs(11115) <= (inputs(18)) and not (inputs(200));
    layer0_outputs(11116) <= not(inputs(141)) or (inputs(14));
    layer0_outputs(11117) <= not(inputs(177));
    layer0_outputs(11118) <= not((inputs(233)) xor (inputs(30)));
    layer0_outputs(11119) <= not((inputs(91)) or (inputs(142)));
    layer0_outputs(11120) <= not(inputs(125)) or (inputs(32));
    layer0_outputs(11121) <= inputs(28);
    layer0_outputs(11122) <= (inputs(49)) and not (inputs(139));
    layer0_outputs(11123) <= (inputs(105)) and not (inputs(34));
    layer0_outputs(11124) <= inputs(98);
    layer0_outputs(11125) <= not(inputs(21));
    layer0_outputs(11126) <= inputs(15);
    layer0_outputs(11127) <= (inputs(50)) or (inputs(236));
    layer0_outputs(11128) <= (inputs(199)) xor (inputs(237));
    layer0_outputs(11129) <= '0';
    layer0_outputs(11130) <= (inputs(116)) xor (inputs(128));
    layer0_outputs(11131) <= not(inputs(228)) or (inputs(14));
    layer0_outputs(11132) <= (inputs(217)) and not (inputs(145));
    layer0_outputs(11133) <= '1';
    layer0_outputs(11134) <= (inputs(71)) or (inputs(109));
    layer0_outputs(11135) <= not(inputs(67));
    layer0_outputs(11136) <= '0';
    layer0_outputs(11137) <= (inputs(88)) or (inputs(159));
    layer0_outputs(11138) <= (inputs(64)) or (inputs(1));
    layer0_outputs(11139) <= not(inputs(41));
    layer0_outputs(11140) <= inputs(213);
    layer0_outputs(11141) <= (inputs(32)) xor (inputs(239));
    layer0_outputs(11142) <= not((inputs(187)) xor (inputs(251)));
    layer0_outputs(11143) <= (inputs(66)) or (inputs(138));
    layer0_outputs(11144) <= not(inputs(63));
    layer0_outputs(11145) <= (inputs(156)) xor (inputs(106));
    layer0_outputs(11146) <= (inputs(122)) and not (inputs(178));
    layer0_outputs(11147) <= (inputs(53)) xor (inputs(45));
    layer0_outputs(11148) <= not((inputs(209)) xor (inputs(174)));
    layer0_outputs(11149) <= not(inputs(29)) or (inputs(102));
    layer0_outputs(11150) <= not(inputs(22)) or (inputs(225));
    layer0_outputs(11151) <= inputs(90);
    layer0_outputs(11152) <= (inputs(127)) or (inputs(82));
    layer0_outputs(11153) <= (inputs(45)) xor (inputs(143));
    layer0_outputs(11154) <= (inputs(1)) xor (inputs(64));
    layer0_outputs(11155) <= not(inputs(94));
    layer0_outputs(11156) <= '0';
    layer0_outputs(11157) <= (inputs(182)) or (inputs(158));
    layer0_outputs(11158) <= inputs(146);
    layer0_outputs(11159) <= inputs(92);
    layer0_outputs(11160) <= inputs(190);
    layer0_outputs(11161) <= not((inputs(171)) xor (inputs(175)));
    layer0_outputs(11162) <= (inputs(14)) xor (inputs(111));
    layer0_outputs(11163) <= not(inputs(118));
    layer0_outputs(11164) <= (inputs(221)) or (inputs(87));
    layer0_outputs(11165) <= (inputs(80)) xor (inputs(191));
    layer0_outputs(11166) <= (inputs(163)) or (inputs(51));
    layer0_outputs(11167) <= inputs(203);
    layer0_outputs(11168) <= (inputs(85)) and not (inputs(92));
    layer0_outputs(11169) <= (inputs(22)) or (inputs(79));
    layer0_outputs(11170) <= not(inputs(90));
    layer0_outputs(11171) <= (inputs(115)) and not (inputs(179));
    layer0_outputs(11172) <= not(inputs(177));
    layer0_outputs(11173) <= inputs(164);
    layer0_outputs(11174) <= '1';
    layer0_outputs(11175) <= not((inputs(55)) xor (inputs(46)));
    layer0_outputs(11176) <= inputs(134);
    layer0_outputs(11177) <= not((inputs(169)) or (inputs(252)));
    layer0_outputs(11178) <= (inputs(198)) and not (inputs(156));
    layer0_outputs(11179) <= (inputs(116)) or (inputs(202));
    layer0_outputs(11180) <= not(inputs(136)) or (inputs(250));
    layer0_outputs(11181) <= not(inputs(25)) or (inputs(176));
    layer0_outputs(11182) <= not((inputs(156)) xor (inputs(103)));
    layer0_outputs(11183) <= not((inputs(126)) or (inputs(85)));
    layer0_outputs(11184) <= (inputs(10)) or (inputs(124));
    layer0_outputs(11185) <= not((inputs(194)) xor (inputs(222)));
    layer0_outputs(11186) <= (inputs(189)) and not (inputs(241));
    layer0_outputs(11187) <= not(inputs(188)) or (inputs(56));
    layer0_outputs(11188) <= not((inputs(175)) xor (inputs(163)));
    layer0_outputs(11189) <= (inputs(24)) and not (inputs(202));
    layer0_outputs(11190) <= (inputs(5)) or (inputs(136));
    layer0_outputs(11191) <= not(inputs(104));
    layer0_outputs(11192) <= not((inputs(234)) or (inputs(35)));
    layer0_outputs(11193) <= not(inputs(221)) or (inputs(205));
    layer0_outputs(11194) <= (inputs(119)) and not (inputs(221));
    layer0_outputs(11195) <= not(inputs(101));
    layer0_outputs(11196) <= not((inputs(62)) xor (inputs(7)));
    layer0_outputs(11197) <= inputs(246);
    layer0_outputs(11198) <= (inputs(51)) xor (inputs(54));
    layer0_outputs(11199) <= not((inputs(37)) xor (inputs(5)));
    layer0_outputs(11200) <= not(inputs(21)) or (inputs(173));
    layer0_outputs(11201) <= (inputs(147)) or (inputs(130));
    layer0_outputs(11202) <= (inputs(65)) and not (inputs(128));
    layer0_outputs(11203) <= not(inputs(244)) or (inputs(105));
    layer0_outputs(11204) <= (inputs(124)) or (inputs(130));
    layer0_outputs(11205) <= not(inputs(88));
    layer0_outputs(11206) <= (inputs(158)) xor (inputs(111));
    layer0_outputs(11207) <= (inputs(204)) and not (inputs(98));
    layer0_outputs(11208) <= not((inputs(139)) and (inputs(1)));
    layer0_outputs(11209) <= not(inputs(95));
    layer0_outputs(11210) <= (inputs(104)) xor (inputs(125));
    layer0_outputs(11211) <= (inputs(149)) or (inputs(8));
    layer0_outputs(11212) <= (inputs(149)) and not (inputs(82));
    layer0_outputs(11213) <= not((inputs(4)) and (inputs(67)));
    layer0_outputs(11214) <= not(inputs(206));
    layer0_outputs(11215) <= inputs(108);
    layer0_outputs(11216) <= not(inputs(81));
    layer0_outputs(11217) <= not((inputs(249)) xor (inputs(250)));
    layer0_outputs(11218) <= inputs(189);
    layer0_outputs(11219) <= not((inputs(133)) or (inputs(209)));
    layer0_outputs(11220) <= (inputs(181)) or (inputs(217));
    layer0_outputs(11221) <= not(inputs(188));
    layer0_outputs(11222) <= '0';
    layer0_outputs(11223) <= (inputs(231)) or (inputs(222));
    layer0_outputs(11224) <= not((inputs(213)) or (inputs(189)));
    layer0_outputs(11225) <= (inputs(147)) or (inputs(251));
    layer0_outputs(11226) <= not((inputs(31)) xor (inputs(229)));
    layer0_outputs(11227) <= (inputs(221)) or (inputs(103));
    layer0_outputs(11228) <= inputs(229);
    layer0_outputs(11229) <= not(inputs(231)) or (inputs(110));
    layer0_outputs(11230) <= (inputs(75)) or (inputs(37));
    layer0_outputs(11231) <= (inputs(63)) or (inputs(77));
    layer0_outputs(11232) <= not((inputs(99)) or (inputs(216)));
    layer0_outputs(11233) <= (inputs(26)) and not (inputs(90));
    layer0_outputs(11234) <= '0';
    layer0_outputs(11235) <= (inputs(165)) and not (inputs(76));
    layer0_outputs(11236) <= (inputs(221)) and not (inputs(93));
    layer0_outputs(11237) <= not((inputs(162)) or (inputs(2)));
    layer0_outputs(11238) <= not(inputs(45));
    layer0_outputs(11239) <= not((inputs(249)) xor (inputs(216)));
    layer0_outputs(11240) <= (inputs(189)) or (inputs(237));
    layer0_outputs(11241) <= not((inputs(64)) xor (inputs(91)));
    layer0_outputs(11242) <= (inputs(195)) or (inputs(129));
    layer0_outputs(11243) <= (inputs(235)) xor (inputs(184));
    layer0_outputs(11244) <= (inputs(173)) and not (inputs(33));
    layer0_outputs(11245) <= not(inputs(86));
    layer0_outputs(11246) <= not((inputs(43)) or (inputs(242)));
    layer0_outputs(11247) <= not((inputs(44)) or (inputs(233)));
    layer0_outputs(11248) <= not((inputs(91)) xor (inputs(211)));
    layer0_outputs(11249) <= (inputs(155)) xor (inputs(70));
    layer0_outputs(11250) <= (inputs(204)) xor (inputs(163));
    layer0_outputs(11251) <= (inputs(159)) xor (inputs(190));
    layer0_outputs(11252) <= (inputs(14)) or (inputs(217));
    layer0_outputs(11253) <= not((inputs(168)) or (inputs(2)));
    layer0_outputs(11254) <= (inputs(68)) or (inputs(66));
    layer0_outputs(11255) <= not(inputs(46));
    layer0_outputs(11256) <= not((inputs(70)) xor (inputs(58)));
    layer0_outputs(11257) <= (inputs(169)) or (inputs(132));
    layer0_outputs(11258) <= not((inputs(156)) xor (inputs(220)));
    layer0_outputs(11259) <= (inputs(65)) or (inputs(28));
    layer0_outputs(11260) <= (inputs(246)) and not (inputs(110));
    layer0_outputs(11261) <= (inputs(65)) and not (inputs(149));
    layer0_outputs(11262) <= not(inputs(233)) or (inputs(161));
    layer0_outputs(11263) <= not((inputs(204)) and (inputs(6)));
    layer0_outputs(11264) <= not(inputs(25));
    layer0_outputs(11265) <= (inputs(19)) xor (inputs(47));
    layer0_outputs(11266) <= not((inputs(38)) xor (inputs(172)));
    layer0_outputs(11267) <= (inputs(197)) and not (inputs(156));
    layer0_outputs(11268) <= not(inputs(149)) or (inputs(137));
    layer0_outputs(11269) <= not(inputs(139));
    layer0_outputs(11270) <= not((inputs(237)) and (inputs(158)));
    layer0_outputs(11271) <= not(inputs(236));
    layer0_outputs(11272) <= (inputs(36)) and not (inputs(56));
    layer0_outputs(11273) <= (inputs(253)) or (inputs(168));
    layer0_outputs(11274) <= not((inputs(11)) xor (inputs(216)));
    layer0_outputs(11275) <= (inputs(67)) and (inputs(235));
    layer0_outputs(11276) <= inputs(209);
    layer0_outputs(11277) <= not((inputs(10)) or (inputs(155)));
    layer0_outputs(11278) <= not(inputs(136));
    layer0_outputs(11279) <= not(inputs(90)) or (inputs(50));
    layer0_outputs(11280) <= (inputs(169)) or (inputs(160));
    layer0_outputs(11281) <= not(inputs(46)) or (inputs(255));
    layer0_outputs(11282) <= not((inputs(138)) xor (inputs(140)));
    layer0_outputs(11283) <= not((inputs(147)) or (inputs(40)));
    layer0_outputs(11284) <= inputs(53);
    layer0_outputs(11285) <= not((inputs(66)) xor (inputs(67)));
    layer0_outputs(11286) <= not(inputs(119)) or (inputs(12));
    layer0_outputs(11287) <= not(inputs(154));
    layer0_outputs(11288) <= inputs(183);
    layer0_outputs(11289) <= not(inputs(45));
    layer0_outputs(11290) <= not(inputs(156)) or (inputs(73));
    layer0_outputs(11291) <= not((inputs(254)) or (inputs(13)));
    layer0_outputs(11292) <= '0';
    layer0_outputs(11293) <= (inputs(216)) or (inputs(161));
    layer0_outputs(11294) <= not((inputs(12)) xor (inputs(55)));
    layer0_outputs(11295) <= not(inputs(181)) or (inputs(241));
    layer0_outputs(11296) <= not((inputs(44)) or (inputs(73)));
    layer0_outputs(11297) <= not((inputs(35)) or (inputs(111)));
    layer0_outputs(11298) <= (inputs(171)) or (inputs(121));
    layer0_outputs(11299) <= not((inputs(133)) or (inputs(155)));
    layer0_outputs(11300) <= '0';
    layer0_outputs(11301) <= not((inputs(218)) or (inputs(174)));
    layer0_outputs(11302) <= inputs(89);
    layer0_outputs(11303) <= inputs(211);
    layer0_outputs(11304) <= not((inputs(204)) and (inputs(167)));
    layer0_outputs(11305) <= (inputs(0)) or (inputs(48));
    layer0_outputs(11306) <= (inputs(241)) or (inputs(191));
    layer0_outputs(11307) <= inputs(72);
    layer0_outputs(11308) <= (inputs(178)) and (inputs(131));
    layer0_outputs(11309) <= not((inputs(103)) or (inputs(61)));
    layer0_outputs(11310) <= (inputs(220)) or (inputs(56));
    layer0_outputs(11311) <= not((inputs(124)) or (inputs(15)));
    layer0_outputs(11312) <= (inputs(20)) or (inputs(223));
    layer0_outputs(11313) <= (inputs(50)) xor (inputs(31));
    layer0_outputs(11314) <= not((inputs(200)) xor (inputs(170)));
    layer0_outputs(11315) <= inputs(216);
    layer0_outputs(11316) <= (inputs(20)) or (inputs(104));
    layer0_outputs(11317) <= not((inputs(61)) xor (inputs(157)));
    layer0_outputs(11318) <= (inputs(74)) and not (inputs(203));
    layer0_outputs(11319) <= not(inputs(148));
    layer0_outputs(11320) <= inputs(250);
    layer0_outputs(11321) <= not(inputs(103));
    layer0_outputs(11322) <= (inputs(156)) and not (inputs(62));
    layer0_outputs(11323) <= (inputs(169)) and not (inputs(30));
    layer0_outputs(11324) <= not(inputs(101));
    layer0_outputs(11325) <= not((inputs(45)) xor (inputs(1)));
    layer0_outputs(11326) <= inputs(10);
    layer0_outputs(11327) <= inputs(202);
    layer0_outputs(11328) <= not((inputs(168)) xor (inputs(121)));
    layer0_outputs(11329) <= not((inputs(91)) and (inputs(75)));
    layer0_outputs(11330) <= not((inputs(159)) or (inputs(112)));
    layer0_outputs(11331) <= not(inputs(44)) or (inputs(102));
    layer0_outputs(11332) <= (inputs(52)) xor (inputs(240));
    layer0_outputs(11333) <= (inputs(173)) xor (inputs(245));
    layer0_outputs(11334) <= not(inputs(74));
    layer0_outputs(11335) <= not((inputs(186)) xor (inputs(205)));
    layer0_outputs(11336) <= inputs(176);
    layer0_outputs(11337) <= not((inputs(22)) or (inputs(141)));
    layer0_outputs(11338) <= inputs(76);
    layer0_outputs(11339) <= '1';
    layer0_outputs(11340) <= (inputs(138)) xor (inputs(248));
    layer0_outputs(11341) <= not(inputs(230));
    layer0_outputs(11342) <= (inputs(215)) xor (inputs(244));
    layer0_outputs(11343) <= inputs(168);
    layer0_outputs(11344) <= (inputs(84)) and not (inputs(153));
    layer0_outputs(11345) <= (inputs(61)) xor (inputs(29));
    layer0_outputs(11346) <= not(inputs(152));
    layer0_outputs(11347) <= (inputs(198)) xor (inputs(226));
    layer0_outputs(11348) <= (inputs(184)) and (inputs(106));
    layer0_outputs(11349) <= (inputs(170)) or (inputs(36));
    layer0_outputs(11350) <= not((inputs(153)) or (inputs(106)));
    layer0_outputs(11351) <= not(inputs(28));
    layer0_outputs(11352) <= (inputs(41)) and not (inputs(243));
    layer0_outputs(11353) <= (inputs(240)) or (inputs(84));
    layer0_outputs(11354) <= not(inputs(67));
    layer0_outputs(11355) <= not(inputs(36));
    layer0_outputs(11356) <= not((inputs(0)) or (inputs(28)));
    layer0_outputs(11357) <= (inputs(142)) xor (inputs(32));
    layer0_outputs(11358) <= not(inputs(23)) or (inputs(31));
    layer0_outputs(11359) <= (inputs(31)) and not (inputs(253));
    layer0_outputs(11360) <= '0';
    layer0_outputs(11361) <= not(inputs(228));
    layer0_outputs(11362) <= (inputs(100)) and not (inputs(26));
    layer0_outputs(11363) <= not((inputs(172)) or (inputs(180)));
    layer0_outputs(11364) <= inputs(179);
    layer0_outputs(11365) <= inputs(231);
    layer0_outputs(11366) <= not(inputs(137)) or (inputs(145));
    layer0_outputs(11367) <= inputs(249);
    layer0_outputs(11368) <= not(inputs(114));
    layer0_outputs(11369) <= (inputs(48)) and not (inputs(26));
    layer0_outputs(11370) <= not((inputs(163)) or (inputs(61)));
    layer0_outputs(11371) <= not(inputs(120));
    layer0_outputs(11372) <= not(inputs(8)) or (inputs(219));
    layer0_outputs(11373) <= not(inputs(161));
    layer0_outputs(11374) <= '0';
    layer0_outputs(11375) <= not(inputs(104)) or (inputs(181));
    layer0_outputs(11376) <= not(inputs(38)) or (inputs(145));
    layer0_outputs(11377) <= (inputs(248)) or (inputs(118));
    layer0_outputs(11378) <= (inputs(49)) and not (inputs(50));
    layer0_outputs(11379) <= (inputs(159)) or (inputs(56));
    layer0_outputs(11380) <= not((inputs(217)) xor (inputs(74)));
    layer0_outputs(11381) <= (inputs(193)) or (inputs(113));
    layer0_outputs(11382) <= not((inputs(7)) xor (inputs(40)));
    layer0_outputs(11383) <= not((inputs(209)) xor (inputs(231)));
    layer0_outputs(11384) <= (inputs(16)) or (inputs(190));
    layer0_outputs(11385) <= inputs(42);
    layer0_outputs(11386) <= not(inputs(187)) or (inputs(31));
    layer0_outputs(11387) <= (inputs(108)) and (inputs(61));
    layer0_outputs(11388) <= (inputs(152)) or (inputs(222));
    layer0_outputs(11389) <= not((inputs(171)) xor (inputs(54)));
    layer0_outputs(11390) <= (inputs(188)) and not (inputs(148));
    layer0_outputs(11391) <= not((inputs(242)) xor (inputs(56)));
    layer0_outputs(11392) <= not(inputs(109)) or (inputs(152));
    layer0_outputs(11393) <= (inputs(37)) and not (inputs(175));
    layer0_outputs(11394) <= inputs(6);
    layer0_outputs(11395) <= inputs(82);
    layer0_outputs(11396) <= inputs(107);
    layer0_outputs(11397) <= not(inputs(114));
    layer0_outputs(11398) <= not((inputs(233)) xor (inputs(216)));
    layer0_outputs(11399) <= not(inputs(77)) or (inputs(244));
    layer0_outputs(11400) <= (inputs(132)) and not (inputs(217));
    layer0_outputs(11401) <= not((inputs(13)) xor (inputs(142)));
    layer0_outputs(11402) <= inputs(228);
    layer0_outputs(11403) <= inputs(62);
    layer0_outputs(11404) <= (inputs(110)) or (inputs(151));
    layer0_outputs(11405) <= not((inputs(18)) or (inputs(19)));
    layer0_outputs(11406) <= not((inputs(192)) or (inputs(63)));
    layer0_outputs(11407) <= not(inputs(148));
    layer0_outputs(11408) <= not(inputs(249));
    layer0_outputs(11409) <= not((inputs(211)) or (inputs(180)));
    layer0_outputs(11410) <= (inputs(109)) xor (inputs(116));
    layer0_outputs(11411) <= not((inputs(58)) and (inputs(172)));
    layer0_outputs(11412) <= (inputs(122)) and (inputs(42));
    layer0_outputs(11413) <= not(inputs(21));
    layer0_outputs(11414) <= not((inputs(248)) xor (inputs(37)));
    layer0_outputs(11415) <= not(inputs(59)) or (inputs(88));
    layer0_outputs(11416) <= inputs(197);
    layer0_outputs(11417) <= not(inputs(210)) or (inputs(30));
    layer0_outputs(11418) <= (inputs(171)) and not (inputs(23));
    layer0_outputs(11419) <= (inputs(198)) and not (inputs(192));
    layer0_outputs(11420) <= (inputs(18)) and not (inputs(214));
    layer0_outputs(11421) <= not(inputs(198)) or (inputs(130));
    layer0_outputs(11422) <= not(inputs(17)) or (inputs(64));
    layer0_outputs(11423) <= (inputs(182)) or (inputs(48));
    layer0_outputs(11424) <= not((inputs(164)) xor (inputs(118)));
    layer0_outputs(11425) <= not((inputs(47)) xor (inputs(18)));
    layer0_outputs(11426) <= (inputs(11)) and not (inputs(203));
    layer0_outputs(11427) <= (inputs(77)) and not (inputs(2));
    layer0_outputs(11428) <= not(inputs(200)) or (inputs(50));
    layer0_outputs(11429) <= not(inputs(105)) or (inputs(159));
    layer0_outputs(11430) <= (inputs(100)) xor (inputs(131));
    layer0_outputs(11431) <= not(inputs(123)) or (inputs(227));
    layer0_outputs(11432) <= (inputs(108)) and not (inputs(250));
    layer0_outputs(11433) <= inputs(165);
    layer0_outputs(11434) <= not((inputs(91)) or (inputs(225)));
    layer0_outputs(11435) <= (inputs(255)) xor (inputs(218));
    layer0_outputs(11436) <= not((inputs(132)) or (inputs(165)));
    layer0_outputs(11437) <= not(inputs(59));
    layer0_outputs(11438) <= (inputs(130)) or (inputs(58));
    layer0_outputs(11439) <= not(inputs(130));
    layer0_outputs(11440) <= (inputs(166)) or (inputs(80));
    layer0_outputs(11441) <= (inputs(116)) and not (inputs(164));
    layer0_outputs(11442) <= not((inputs(63)) xor (inputs(200)));
    layer0_outputs(11443) <= not((inputs(243)) or (inputs(86)));
    layer0_outputs(11444) <= not(inputs(232)) or (inputs(183));
    layer0_outputs(11445) <= (inputs(128)) xor (inputs(116));
    layer0_outputs(11446) <= not(inputs(133));
    layer0_outputs(11447) <= inputs(93);
    layer0_outputs(11448) <= not((inputs(21)) or (inputs(55)));
    layer0_outputs(11449) <= not((inputs(229)) xor (inputs(133)));
    layer0_outputs(11450) <= not(inputs(181));
    layer0_outputs(11451) <= (inputs(41)) and (inputs(149));
    layer0_outputs(11452) <= not(inputs(84));
    layer0_outputs(11453) <= (inputs(76)) and not (inputs(190));
    layer0_outputs(11454) <= not((inputs(33)) xor (inputs(126)));
    layer0_outputs(11455) <= not((inputs(177)) xor (inputs(97)));
    layer0_outputs(11456) <= (inputs(200)) or (inputs(17));
    layer0_outputs(11457) <= (inputs(126)) or (inputs(56));
    layer0_outputs(11458) <= (inputs(221)) xor (inputs(235));
    layer0_outputs(11459) <= not(inputs(170));
    layer0_outputs(11460) <= (inputs(235)) or (inputs(193));
    layer0_outputs(11461) <= inputs(166);
    layer0_outputs(11462) <= not((inputs(130)) or (inputs(198)));
    layer0_outputs(11463) <= not((inputs(118)) xor (inputs(144)));
    layer0_outputs(11464) <= inputs(148);
    layer0_outputs(11465) <= inputs(107);
    layer0_outputs(11466) <= not(inputs(193)) or (inputs(173));
    layer0_outputs(11467) <= not(inputs(152));
    layer0_outputs(11468) <= (inputs(155)) or (inputs(22));
    layer0_outputs(11469) <= not((inputs(214)) and (inputs(213)));
    layer0_outputs(11470) <= not(inputs(22)) or (inputs(128));
    layer0_outputs(11471) <= inputs(234);
    layer0_outputs(11472) <= (inputs(95)) xor (inputs(246));
    layer0_outputs(11473) <= inputs(99);
    layer0_outputs(11474) <= inputs(178);
    layer0_outputs(11475) <= (inputs(229)) xor (inputs(194));
    layer0_outputs(11476) <= not(inputs(6));
    layer0_outputs(11477) <= not(inputs(9)) or (inputs(13));
    layer0_outputs(11478) <= not(inputs(10)) or (inputs(173));
    layer0_outputs(11479) <= (inputs(110)) xor (inputs(56));
    layer0_outputs(11480) <= '0';
    layer0_outputs(11481) <= (inputs(89)) or (inputs(103));
    layer0_outputs(11482) <= not(inputs(145));
    layer0_outputs(11483) <= (inputs(240)) and not (inputs(0));
    layer0_outputs(11484) <= not(inputs(224));
    layer0_outputs(11485) <= not((inputs(14)) xor (inputs(104)));
    layer0_outputs(11486) <= not((inputs(115)) and (inputs(159)));
    layer0_outputs(11487) <= not(inputs(38));
    layer0_outputs(11488) <= not((inputs(183)) xor (inputs(63)));
    layer0_outputs(11489) <= (inputs(110)) xor (inputs(107));
    layer0_outputs(11490) <= (inputs(153)) xor (inputs(103));
    layer0_outputs(11491) <= (inputs(117)) or (inputs(80));
    layer0_outputs(11492) <= not(inputs(27));
    layer0_outputs(11493) <= (inputs(87)) and not (inputs(78));
    layer0_outputs(11494) <= (inputs(91)) xor (inputs(92));
    layer0_outputs(11495) <= not((inputs(176)) xor (inputs(245)));
    layer0_outputs(11496) <= inputs(122);
    layer0_outputs(11497) <= inputs(189);
    layer0_outputs(11498) <= inputs(125);
    layer0_outputs(11499) <= (inputs(192)) and not (inputs(41));
    layer0_outputs(11500) <= not((inputs(233)) xor (inputs(148)));
    layer0_outputs(11501) <= not((inputs(73)) xor (inputs(142)));
    layer0_outputs(11502) <= not((inputs(115)) xor (inputs(219)));
    layer0_outputs(11503) <= not(inputs(211)) or (inputs(111));
    layer0_outputs(11504) <= (inputs(11)) and (inputs(84));
    layer0_outputs(11505) <= not((inputs(237)) xor (inputs(157)));
    layer0_outputs(11506) <= (inputs(100)) and not (inputs(223));
    layer0_outputs(11507) <= (inputs(249)) and not (inputs(109));
    layer0_outputs(11508) <= inputs(138);
    layer0_outputs(11509) <= inputs(106);
    layer0_outputs(11510) <= inputs(131);
    layer0_outputs(11511) <= not((inputs(227)) or (inputs(99)));
    layer0_outputs(11512) <= inputs(203);
    layer0_outputs(11513) <= (inputs(87)) xor (inputs(71));
    layer0_outputs(11514) <= inputs(117);
    layer0_outputs(11515) <= (inputs(248)) and (inputs(182));
    layer0_outputs(11516) <= (inputs(240)) xor (inputs(97));
    layer0_outputs(11517) <= (inputs(244)) or (inputs(1));
    layer0_outputs(11518) <= not(inputs(41));
    layer0_outputs(11519) <= (inputs(106)) and not (inputs(158));
    layer0_outputs(11520) <= (inputs(219)) and (inputs(182));
    layer0_outputs(11521) <= inputs(28);
    layer0_outputs(11522) <= not(inputs(105)) or (inputs(186));
    layer0_outputs(11523) <= (inputs(224)) xor (inputs(121));
    layer0_outputs(11524) <= not((inputs(224)) xor (inputs(6)));
    layer0_outputs(11525) <= (inputs(106)) xor (inputs(244));
    layer0_outputs(11526) <= (inputs(234)) and (inputs(212));
    layer0_outputs(11527) <= (inputs(150)) xor (inputs(106));
    layer0_outputs(11528) <= not((inputs(30)) or (inputs(60)));
    layer0_outputs(11529) <= inputs(111);
    layer0_outputs(11530) <= (inputs(81)) or (inputs(61));
    layer0_outputs(11531) <= (inputs(31)) or (inputs(101));
    layer0_outputs(11532) <= (inputs(178)) and not (inputs(243));
    layer0_outputs(11533) <= not(inputs(178));
    layer0_outputs(11534) <= inputs(76);
    layer0_outputs(11535) <= inputs(238);
    layer0_outputs(11536) <= (inputs(159)) or (inputs(190));
    layer0_outputs(11537) <= (inputs(84)) or (inputs(12));
    layer0_outputs(11538) <= not((inputs(221)) or (inputs(182)));
    layer0_outputs(11539) <= inputs(99);
    layer0_outputs(11540) <= not(inputs(41));
    layer0_outputs(11541) <= not(inputs(163));
    layer0_outputs(11542) <= not(inputs(228)) or (inputs(112));
    layer0_outputs(11543) <= not((inputs(114)) or (inputs(238)));
    layer0_outputs(11544) <= (inputs(124)) and not (inputs(113));
    layer0_outputs(11545) <= not(inputs(89));
    layer0_outputs(11546) <= not(inputs(3));
    layer0_outputs(11547) <= (inputs(163)) xor (inputs(245));
    layer0_outputs(11548) <= not(inputs(94)) or (inputs(35));
    layer0_outputs(11549) <= (inputs(165)) and not (inputs(106));
    layer0_outputs(11550) <= inputs(97);
    layer0_outputs(11551) <= not(inputs(40)) or (inputs(112));
    layer0_outputs(11552) <= (inputs(153)) and not (inputs(143));
    layer0_outputs(11553) <= inputs(98);
    layer0_outputs(11554) <= (inputs(48)) xor (inputs(44));
    layer0_outputs(11555) <= (inputs(76)) or (inputs(23));
    layer0_outputs(11556) <= inputs(135);
    layer0_outputs(11557) <= inputs(146);
    layer0_outputs(11558) <= not(inputs(232));
    layer0_outputs(11559) <= not(inputs(140)) or (inputs(83));
    layer0_outputs(11560) <= inputs(248);
    layer0_outputs(11561) <= inputs(116);
    layer0_outputs(11562) <= inputs(203);
    layer0_outputs(11563) <= (inputs(153)) xor (inputs(107));
    layer0_outputs(11564) <= inputs(209);
    layer0_outputs(11565) <= (inputs(118)) xor (inputs(221));
    layer0_outputs(11566) <= not(inputs(202)) or (inputs(199));
    layer0_outputs(11567) <= not(inputs(143)) or (inputs(38));
    layer0_outputs(11568) <= (inputs(168)) xor (inputs(212));
    layer0_outputs(11569) <= (inputs(201)) or (inputs(182));
    layer0_outputs(11570) <= not((inputs(210)) or (inputs(211)));
    layer0_outputs(11571) <= not(inputs(40));
    layer0_outputs(11572) <= not((inputs(140)) or (inputs(104)));
    layer0_outputs(11573) <= (inputs(111)) xor (inputs(179));
    layer0_outputs(11574) <= not(inputs(184));
    layer0_outputs(11575) <= not(inputs(68)) or (inputs(59));
    layer0_outputs(11576) <= (inputs(128)) or (inputs(205));
    layer0_outputs(11577) <= inputs(179);
    layer0_outputs(11578) <= not(inputs(86)) or (inputs(149));
    layer0_outputs(11579) <= inputs(239);
    layer0_outputs(11580) <= (inputs(143)) xor (inputs(14));
    layer0_outputs(11581) <= not(inputs(163));
    layer0_outputs(11582) <= not(inputs(40)) or (inputs(130));
    layer0_outputs(11583) <= inputs(162);
    layer0_outputs(11584) <= (inputs(99)) xor (inputs(53));
    layer0_outputs(11585) <= (inputs(136)) or (inputs(150));
    layer0_outputs(11586) <= (inputs(115)) and not (inputs(87));
    layer0_outputs(11587) <= not(inputs(118)) or (inputs(2));
    layer0_outputs(11588) <= not((inputs(80)) or (inputs(144)));
    layer0_outputs(11589) <= not(inputs(233));
    layer0_outputs(11590) <= not((inputs(126)) xor (inputs(159)));
    layer0_outputs(11591) <= '1';
    layer0_outputs(11592) <= not(inputs(220)) or (inputs(26));
    layer0_outputs(11593) <= (inputs(250)) or (inputs(174));
    layer0_outputs(11594) <= (inputs(53)) and not (inputs(113));
    layer0_outputs(11595) <= not((inputs(128)) or (inputs(253)));
    layer0_outputs(11596) <= not((inputs(30)) xor (inputs(221)));
    layer0_outputs(11597) <= inputs(23);
    layer0_outputs(11598) <= not((inputs(253)) xor (inputs(179)));
    layer0_outputs(11599) <= not(inputs(105));
    layer0_outputs(11600) <= not((inputs(37)) or (inputs(76)));
    layer0_outputs(11601) <= (inputs(199)) and not (inputs(34));
    layer0_outputs(11602) <= (inputs(40)) and not (inputs(243));
    layer0_outputs(11603) <= not(inputs(218)) or (inputs(79));
    layer0_outputs(11604) <= (inputs(78)) xor (inputs(137));
    layer0_outputs(11605) <= not((inputs(239)) xor (inputs(241)));
    layer0_outputs(11606) <= (inputs(114)) and not (inputs(226));
    layer0_outputs(11607) <= (inputs(195)) xor (inputs(93));
    layer0_outputs(11608) <= inputs(55);
    layer0_outputs(11609) <= not(inputs(98));
    layer0_outputs(11610) <= not(inputs(85));
    layer0_outputs(11611) <= (inputs(132)) xor (inputs(148));
    layer0_outputs(11612) <= not((inputs(176)) or (inputs(183)));
    layer0_outputs(11613) <= (inputs(51)) and (inputs(10));
    layer0_outputs(11614) <= not((inputs(27)) xor (inputs(23)));
    layer0_outputs(11615) <= (inputs(144)) xor (inputs(230));
    layer0_outputs(11616) <= not((inputs(107)) or (inputs(202)));
    layer0_outputs(11617) <= not((inputs(79)) or (inputs(161)));
    layer0_outputs(11618) <= (inputs(2)) and not (inputs(34));
    layer0_outputs(11619) <= (inputs(161)) xor (inputs(234));
    layer0_outputs(11620) <= (inputs(91)) xor (inputs(224));
    layer0_outputs(11621) <= not(inputs(85));
    layer0_outputs(11622) <= not(inputs(110));
    layer0_outputs(11623) <= not((inputs(28)) xor (inputs(192)));
    layer0_outputs(11624) <= inputs(22);
    layer0_outputs(11625) <= not(inputs(92));
    layer0_outputs(11626) <= not(inputs(119));
    layer0_outputs(11627) <= (inputs(112)) xor (inputs(67));
    layer0_outputs(11628) <= inputs(174);
    layer0_outputs(11629) <= not(inputs(38));
    layer0_outputs(11630) <= not(inputs(241)) or (inputs(8));
    layer0_outputs(11631) <= inputs(162);
    layer0_outputs(11632) <= not(inputs(99)) or (inputs(224));
    layer0_outputs(11633) <= (inputs(220)) and not (inputs(51));
    layer0_outputs(11634) <= not((inputs(240)) or (inputs(163)));
    layer0_outputs(11635) <= not((inputs(134)) or (inputs(156)));
    layer0_outputs(11636) <= inputs(67);
    layer0_outputs(11637) <= not(inputs(216));
    layer0_outputs(11638) <= inputs(245);
    layer0_outputs(11639) <= not((inputs(45)) xor (inputs(10)));
    layer0_outputs(11640) <= (inputs(25)) and not (inputs(165));
    layer0_outputs(11641) <= inputs(231);
    layer0_outputs(11642) <= inputs(178);
    layer0_outputs(11643) <= not((inputs(42)) and (inputs(186)));
    layer0_outputs(11644) <= not((inputs(15)) xor (inputs(198)));
    layer0_outputs(11645) <= not(inputs(229));
    layer0_outputs(11646) <= (inputs(157)) and (inputs(129));
    layer0_outputs(11647) <= '1';
    layer0_outputs(11648) <= (inputs(57)) and not (inputs(50));
    layer0_outputs(11649) <= not(inputs(129));
    layer0_outputs(11650) <= not(inputs(42));
    layer0_outputs(11651) <= (inputs(234)) and not (inputs(177));
    layer0_outputs(11652) <= (inputs(83)) xor (inputs(129));
    layer0_outputs(11653) <= not(inputs(120));
    layer0_outputs(11654) <= not(inputs(124));
    layer0_outputs(11655) <= inputs(114);
    layer0_outputs(11656) <= inputs(174);
    layer0_outputs(11657) <= '0';
    layer0_outputs(11658) <= not(inputs(158));
    layer0_outputs(11659) <= not(inputs(198)) or (inputs(221));
    layer0_outputs(11660) <= (inputs(96)) xor (inputs(227));
    layer0_outputs(11661) <= not(inputs(228)) or (inputs(66));
    layer0_outputs(11662) <= not((inputs(165)) or (inputs(103)));
    layer0_outputs(11663) <= inputs(212);
    layer0_outputs(11664) <= (inputs(66)) or (inputs(43));
    layer0_outputs(11665) <= not(inputs(154)) or (inputs(44));
    layer0_outputs(11666) <= (inputs(53)) or (inputs(15));
    layer0_outputs(11667) <= inputs(38);
    layer0_outputs(11668) <= not((inputs(52)) or (inputs(92)));
    layer0_outputs(11669) <= not((inputs(45)) xor (inputs(187)));
    layer0_outputs(11670) <= inputs(227);
    layer0_outputs(11671) <= not((inputs(254)) xor (inputs(179)));
    layer0_outputs(11672) <= not((inputs(231)) or (inputs(16)));
    layer0_outputs(11673) <= (inputs(93)) or (inputs(38));
    layer0_outputs(11674) <= (inputs(176)) xor (inputs(53));
    layer0_outputs(11675) <= inputs(166);
    layer0_outputs(11676) <= not(inputs(94));
    layer0_outputs(11677) <= (inputs(44)) and not (inputs(210));
    layer0_outputs(11678) <= (inputs(230)) xor (inputs(37));
    layer0_outputs(11679) <= (inputs(59)) or (inputs(75));
    layer0_outputs(11680) <= not((inputs(56)) or (inputs(134)));
    layer0_outputs(11681) <= not(inputs(131));
    layer0_outputs(11682) <= not((inputs(158)) xor (inputs(105)));
    layer0_outputs(11683) <= not(inputs(152)) or (inputs(109));
    layer0_outputs(11684) <= (inputs(91)) xor (inputs(16));
    layer0_outputs(11685) <= inputs(119);
    layer0_outputs(11686) <= (inputs(148)) xor (inputs(70));
    layer0_outputs(11687) <= not(inputs(212)) or (inputs(133));
    layer0_outputs(11688) <= not((inputs(79)) or (inputs(176)));
    layer0_outputs(11689) <= not((inputs(72)) xor (inputs(39)));
    layer0_outputs(11690) <= not(inputs(58));
    layer0_outputs(11691) <= (inputs(227)) and (inputs(206));
    layer0_outputs(11692) <= inputs(121);
    layer0_outputs(11693) <= not((inputs(75)) or (inputs(97)));
    layer0_outputs(11694) <= not((inputs(102)) xor (inputs(191)));
    layer0_outputs(11695) <= (inputs(140)) xor (inputs(156));
    layer0_outputs(11696) <= (inputs(7)) xor (inputs(16));
    layer0_outputs(11697) <= inputs(68);
    layer0_outputs(11698) <= (inputs(112)) or (inputs(229));
    layer0_outputs(11699) <= inputs(193);
    layer0_outputs(11700) <= inputs(179);
    layer0_outputs(11701) <= inputs(24);
    layer0_outputs(11702) <= not((inputs(7)) or (inputs(252)));
    layer0_outputs(11703) <= inputs(201);
    layer0_outputs(11704) <= not((inputs(101)) and (inputs(229)));
    layer0_outputs(11705) <= (inputs(85)) or (inputs(31));
    layer0_outputs(11706) <= inputs(60);
    layer0_outputs(11707) <= inputs(93);
    layer0_outputs(11708) <= not(inputs(184)) or (inputs(6));
    layer0_outputs(11709) <= (inputs(102)) and not (inputs(158));
    layer0_outputs(11710) <= not((inputs(81)) and (inputs(112)));
    layer0_outputs(11711) <= not((inputs(241)) or (inputs(88)));
    layer0_outputs(11712) <= (inputs(27)) and (inputs(68));
    layer0_outputs(11713) <= not((inputs(15)) and (inputs(50)));
    layer0_outputs(11714) <= (inputs(76)) xor (inputs(24));
    layer0_outputs(11715) <= not(inputs(194)) or (inputs(59));
    layer0_outputs(11716) <= '0';
    layer0_outputs(11717) <= (inputs(204)) and not (inputs(57));
    layer0_outputs(11718) <= (inputs(7)) and not (inputs(248));
    layer0_outputs(11719) <= (inputs(131)) xor (inputs(207));
    layer0_outputs(11720) <= not(inputs(73)) or (inputs(223));
    layer0_outputs(11721) <= not(inputs(20));
    layer0_outputs(11722) <= not((inputs(79)) or (inputs(241)));
    layer0_outputs(11723) <= not((inputs(52)) or (inputs(133)));
    layer0_outputs(11724) <= inputs(86);
    layer0_outputs(11725) <= (inputs(107)) and not (inputs(189));
    layer0_outputs(11726) <= (inputs(28)) or (inputs(128));
    layer0_outputs(11727) <= not((inputs(238)) xor (inputs(102)));
    layer0_outputs(11728) <= inputs(102);
    layer0_outputs(11729) <= (inputs(138)) or (inputs(166));
    layer0_outputs(11730) <= not((inputs(127)) xor (inputs(139)));
    layer0_outputs(11731) <= not((inputs(43)) and (inputs(34)));
    layer0_outputs(11732) <= inputs(113);
    layer0_outputs(11733) <= not(inputs(62)) or (inputs(126));
    layer0_outputs(11734) <= inputs(124);
    layer0_outputs(11735) <= (inputs(71)) xor (inputs(66));
    layer0_outputs(11736) <= not((inputs(2)) xor (inputs(188)));
    layer0_outputs(11737) <= not(inputs(67));
    layer0_outputs(11738) <= not(inputs(86));
    layer0_outputs(11739) <= not(inputs(219)) or (inputs(46));
    layer0_outputs(11740) <= not(inputs(75)) or (inputs(203));
    layer0_outputs(11741) <= not(inputs(105));
    layer0_outputs(11742) <= (inputs(202)) and not (inputs(46));
    layer0_outputs(11743) <= not(inputs(114));
    layer0_outputs(11744) <= (inputs(168)) or (inputs(225));
    layer0_outputs(11745) <= not((inputs(67)) xor (inputs(177)));
    layer0_outputs(11746) <= (inputs(64)) and not (inputs(30));
    layer0_outputs(11747) <= not((inputs(152)) xor (inputs(48)));
    layer0_outputs(11748) <= inputs(39);
    layer0_outputs(11749) <= not(inputs(166)) or (inputs(143));
    layer0_outputs(11750) <= inputs(20);
    layer0_outputs(11751) <= (inputs(70)) xor (inputs(170));
    layer0_outputs(11752) <= not(inputs(90)) or (inputs(252));
    layer0_outputs(11753) <= (inputs(247)) xor (inputs(239));
    layer0_outputs(11754) <= inputs(171);
    layer0_outputs(11755) <= (inputs(77)) and (inputs(213));
    layer0_outputs(11756) <= inputs(49);
    layer0_outputs(11757) <= (inputs(98)) or (inputs(106));
    layer0_outputs(11758) <= not((inputs(88)) and (inputs(103)));
    layer0_outputs(11759) <= (inputs(218)) or (inputs(145));
    layer0_outputs(11760) <= (inputs(241)) or (inputs(67));
    layer0_outputs(11761) <= (inputs(135)) xor (inputs(34));
    layer0_outputs(11762) <= inputs(169);
    layer0_outputs(11763) <= not(inputs(107));
    layer0_outputs(11764) <= inputs(132);
    layer0_outputs(11765) <= not((inputs(182)) xor (inputs(126)));
    layer0_outputs(11766) <= '1';
    layer0_outputs(11767) <= inputs(40);
    layer0_outputs(11768) <= not(inputs(91)) or (inputs(80));
    layer0_outputs(11769) <= not(inputs(147)) or (inputs(80));
    layer0_outputs(11770) <= not(inputs(51));
    layer0_outputs(11771) <= inputs(227);
    layer0_outputs(11772) <= inputs(232);
    layer0_outputs(11773) <= (inputs(34)) xor (inputs(121));
    layer0_outputs(11774) <= not((inputs(179)) or (inputs(235)));
    layer0_outputs(11775) <= inputs(91);
    layer0_outputs(11776) <= (inputs(200)) and not (inputs(117));
    layer0_outputs(11777) <= (inputs(177)) and not (inputs(70));
    layer0_outputs(11778) <= (inputs(66)) or (inputs(212));
    layer0_outputs(11779) <= not((inputs(114)) or (inputs(147)));
    layer0_outputs(11780) <= (inputs(104)) and not (inputs(214));
    layer0_outputs(11781) <= not(inputs(202));
    layer0_outputs(11782) <= inputs(134);
    layer0_outputs(11783) <= not((inputs(0)) or (inputs(144)));
    layer0_outputs(11784) <= inputs(188);
    layer0_outputs(11785) <= not(inputs(126));
    layer0_outputs(11786) <= inputs(185);
    layer0_outputs(11787) <= not(inputs(176)) or (inputs(95));
    layer0_outputs(11788) <= (inputs(108)) xor (inputs(51));
    layer0_outputs(11789) <= not((inputs(151)) xor (inputs(18)));
    layer0_outputs(11790) <= not((inputs(216)) or (inputs(1)));
    layer0_outputs(11791) <= not((inputs(222)) or (inputs(166)));
    layer0_outputs(11792) <= (inputs(208)) xor (inputs(160));
    layer0_outputs(11793) <= inputs(111);
    layer0_outputs(11794) <= inputs(84);
    layer0_outputs(11795) <= inputs(121);
    layer0_outputs(11796) <= not((inputs(116)) or (inputs(176)));
    layer0_outputs(11797) <= not(inputs(72)) or (inputs(69));
    layer0_outputs(11798) <= (inputs(71)) and (inputs(115));
    layer0_outputs(11799) <= (inputs(57)) xor (inputs(240));
    layer0_outputs(11800) <= (inputs(85)) and not (inputs(17));
    layer0_outputs(11801) <= inputs(146);
    layer0_outputs(11802) <= (inputs(242)) or (inputs(192));
    layer0_outputs(11803) <= (inputs(186)) or (inputs(244));
    layer0_outputs(11804) <= not(inputs(100));
    layer0_outputs(11805) <= '0';
    layer0_outputs(11806) <= (inputs(36)) xor (inputs(149));
    layer0_outputs(11807) <= inputs(25);
    layer0_outputs(11808) <= not(inputs(140)) or (inputs(19));
    layer0_outputs(11809) <= '1';
    layer0_outputs(11810) <= '0';
    layer0_outputs(11811) <= (inputs(58)) and not (inputs(37));
    layer0_outputs(11812) <= '1';
    layer0_outputs(11813) <= not((inputs(59)) xor (inputs(183)));
    layer0_outputs(11814) <= (inputs(118)) xor (inputs(55));
    layer0_outputs(11815) <= not((inputs(133)) or (inputs(229)));
    layer0_outputs(11816) <= '1';
    layer0_outputs(11817) <= (inputs(22)) or (inputs(68));
    layer0_outputs(11818) <= (inputs(236)) and not (inputs(83));
    layer0_outputs(11819) <= (inputs(25)) or (inputs(190));
    layer0_outputs(11820) <= (inputs(154)) or (inputs(88));
    layer0_outputs(11821) <= (inputs(14)) xor (inputs(128));
    layer0_outputs(11822) <= (inputs(119)) and not (inputs(42));
    layer0_outputs(11823) <= not((inputs(187)) or (inputs(208)));
    layer0_outputs(11824) <= not((inputs(22)) and (inputs(51)));
    layer0_outputs(11825) <= not((inputs(64)) or (inputs(19)));
    layer0_outputs(11826) <= not((inputs(55)) or (inputs(141)));
    layer0_outputs(11827) <= (inputs(134)) xor (inputs(42));
    layer0_outputs(11828) <= (inputs(91)) and not (inputs(244));
    layer0_outputs(11829) <= not((inputs(205)) or (inputs(161)));
    layer0_outputs(11830) <= not((inputs(178)) or (inputs(220)));
    layer0_outputs(11831) <= (inputs(17)) xor (inputs(91));
    layer0_outputs(11832) <= (inputs(219)) and not (inputs(148));
    layer0_outputs(11833) <= inputs(193);
    layer0_outputs(11834) <= not(inputs(43));
    layer0_outputs(11835) <= not(inputs(2));
    layer0_outputs(11836) <= inputs(98);
    layer0_outputs(11837) <= '1';
    layer0_outputs(11838) <= (inputs(133)) xor (inputs(86));
    layer0_outputs(11839) <= not(inputs(36));
    layer0_outputs(11840) <= (inputs(202)) and not (inputs(2));
    layer0_outputs(11841) <= not((inputs(46)) xor (inputs(201)));
    layer0_outputs(11842) <= not((inputs(179)) xor (inputs(238)));
    layer0_outputs(11843) <= (inputs(182)) xor (inputs(180));
    layer0_outputs(11844) <= '0';
    layer0_outputs(11845) <= '1';
    layer0_outputs(11846) <= (inputs(173)) or (inputs(171));
    layer0_outputs(11847) <= (inputs(35)) or (inputs(44));
    layer0_outputs(11848) <= not(inputs(58)) or (inputs(15));
    layer0_outputs(11849) <= inputs(178);
    layer0_outputs(11850) <= (inputs(239)) and (inputs(201));
    layer0_outputs(11851) <= (inputs(32)) and (inputs(64));
    layer0_outputs(11852) <= (inputs(22)) and not (inputs(188));
    layer0_outputs(11853) <= not(inputs(28)) or (inputs(149));
    layer0_outputs(11854) <= (inputs(19)) or (inputs(207));
    layer0_outputs(11855) <= not((inputs(85)) or (inputs(62)));
    layer0_outputs(11856) <= inputs(113);
    layer0_outputs(11857) <= (inputs(171)) and (inputs(229));
    layer0_outputs(11858) <= (inputs(161)) xor (inputs(103));
    layer0_outputs(11859) <= (inputs(210)) xor (inputs(189));
    layer0_outputs(11860) <= not((inputs(119)) or (inputs(183)));
    layer0_outputs(11861) <= (inputs(18)) or (inputs(2));
    layer0_outputs(11862) <= (inputs(41)) or (inputs(161));
    layer0_outputs(11863) <= not(inputs(19));
    layer0_outputs(11864) <= not(inputs(200));
    layer0_outputs(11865) <= not(inputs(150)) or (inputs(143));
    layer0_outputs(11866) <= not(inputs(118));
    layer0_outputs(11867) <= not(inputs(150));
    layer0_outputs(11868) <= inputs(108);
    layer0_outputs(11869) <= not((inputs(176)) or (inputs(156)));
    layer0_outputs(11870) <= (inputs(204)) or (inputs(62));
    layer0_outputs(11871) <= (inputs(101)) or (inputs(140));
    layer0_outputs(11872) <= not((inputs(184)) and (inputs(173)));
    layer0_outputs(11873) <= not(inputs(110));
    layer0_outputs(11874) <= not((inputs(106)) xor (inputs(96)));
    layer0_outputs(11875) <= not((inputs(52)) xor (inputs(164)));
    layer0_outputs(11876) <= not(inputs(104));
    layer0_outputs(11877) <= (inputs(27)) and not (inputs(195));
    layer0_outputs(11878) <= (inputs(140)) and not (inputs(227));
    layer0_outputs(11879) <= not((inputs(238)) or (inputs(237)));
    layer0_outputs(11880) <= not((inputs(201)) xor (inputs(233)));
    layer0_outputs(11881) <= not((inputs(148)) or (inputs(247)));
    layer0_outputs(11882) <= not((inputs(155)) or (inputs(183)));
    layer0_outputs(11883) <= not((inputs(48)) xor (inputs(86)));
    layer0_outputs(11884) <= not(inputs(145));
    layer0_outputs(11885) <= not(inputs(106));
    layer0_outputs(11886) <= not((inputs(164)) or (inputs(225)));
    layer0_outputs(11887) <= (inputs(215)) or (inputs(146));
    layer0_outputs(11888) <= (inputs(15)) xor (inputs(195));
    layer0_outputs(11889) <= not((inputs(9)) xor (inputs(57)));
    layer0_outputs(11890) <= inputs(1);
    layer0_outputs(11891) <= (inputs(70)) and not (inputs(126));
    layer0_outputs(11892) <= not(inputs(183));
    layer0_outputs(11893) <= (inputs(21)) or (inputs(19));
    layer0_outputs(11894) <= not((inputs(113)) or (inputs(115)));
    layer0_outputs(11895) <= inputs(116);
    layer0_outputs(11896) <= not((inputs(175)) or (inputs(72)));
    layer0_outputs(11897) <= not((inputs(92)) xor (inputs(2)));
    layer0_outputs(11898) <= '1';
    layer0_outputs(11899) <= not((inputs(177)) or (inputs(157)));
    layer0_outputs(11900) <= (inputs(104)) xor (inputs(5));
    layer0_outputs(11901) <= (inputs(208)) xor (inputs(212));
    layer0_outputs(11902) <= (inputs(212)) xor (inputs(189));
    layer0_outputs(11903) <= (inputs(23)) and not (inputs(224));
    layer0_outputs(11904) <= (inputs(27)) and not (inputs(64));
    layer0_outputs(11905) <= not((inputs(15)) or (inputs(31)));
    layer0_outputs(11906) <= not(inputs(147));
    layer0_outputs(11907) <= not((inputs(43)) xor (inputs(175)));
    layer0_outputs(11908) <= inputs(188);
    layer0_outputs(11909) <= (inputs(19)) or (inputs(35));
    layer0_outputs(11910) <= not(inputs(137));
    layer0_outputs(11911) <= (inputs(24)) and not (inputs(210));
    layer0_outputs(11912) <= (inputs(21)) or (inputs(170));
    layer0_outputs(11913) <= not((inputs(144)) or (inputs(193)));
    layer0_outputs(11914) <= not((inputs(103)) or (inputs(157)));
    layer0_outputs(11915) <= inputs(234);
    layer0_outputs(11916) <= not(inputs(167)) or (inputs(78));
    layer0_outputs(11917) <= inputs(136);
    layer0_outputs(11918) <= (inputs(147)) and not (inputs(45));
    layer0_outputs(11919) <= not((inputs(201)) xor (inputs(191)));
    layer0_outputs(11920) <= (inputs(106)) or (inputs(15));
    layer0_outputs(11921) <= inputs(170);
    layer0_outputs(11922) <= not(inputs(199));
    layer0_outputs(11923) <= '0';
    layer0_outputs(11924) <= not((inputs(116)) or (inputs(7)));
    layer0_outputs(11925) <= (inputs(227)) and (inputs(239));
    layer0_outputs(11926) <= inputs(24);
    layer0_outputs(11927) <= not(inputs(110));
    layer0_outputs(11928) <= not(inputs(235)) or (inputs(66));
    layer0_outputs(11929) <= (inputs(226)) or (inputs(209));
    layer0_outputs(11930) <= not(inputs(30));
    layer0_outputs(11931) <= (inputs(100)) and not (inputs(250));
    layer0_outputs(11932) <= not(inputs(125));
    layer0_outputs(11933) <= (inputs(84)) and not (inputs(145));
    layer0_outputs(11934) <= (inputs(96)) or (inputs(84));
    layer0_outputs(11935) <= inputs(206);
    layer0_outputs(11936) <= not(inputs(243)) or (inputs(73));
    layer0_outputs(11937) <= not(inputs(108)) or (inputs(240));
    layer0_outputs(11938) <= not(inputs(228)) or (inputs(134));
    layer0_outputs(11939) <= not(inputs(98)) or (inputs(47));
    layer0_outputs(11940) <= (inputs(152)) and (inputs(237));
    layer0_outputs(11941) <= not(inputs(53)) or (inputs(242));
    layer0_outputs(11942) <= not(inputs(39)) or (inputs(240));
    layer0_outputs(11943) <= not((inputs(219)) or (inputs(63)));
    layer0_outputs(11944) <= not(inputs(210));
    layer0_outputs(11945) <= not(inputs(214));
    layer0_outputs(11946) <= not((inputs(107)) xor (inputs(125)));
    layer0_outputs(11947) <= not((inputs(165)) xor (inputs(75)));
    layer0_outputs(11948) <= (inputs(77)) and not (inputs(115));
    layer0_outputs(11949) <= (inputs(84)) and not (inputs(234));
    layer0_outputs(11950) <= not(inputs(165));
    layer0_outputs(11951) <= (inputs(171)) or (inputs(191));
    layer0_outputs(11952) <= not(inputs(88));
    layer0_outputs(11953) <= not(inputs(39));
    layer0_outputs(11954) <= (inputs(25)) and (inputs(102));
    layer0_outputs(11955) <= not(inputs(84));
    layer0_outputs(11956) <= not(inputs(228)) or (inputs(64));
    layer0_outputs(11957) <= not(inputs(57));
    layer0_outputs(11958) <= (inputs(209)) xor (inputs(46));
    layer0_outputs(11959) <= not(inputs(54));
    layer0_outputs(11960) <= not(inputs(221));
    layer0_outputs(11961) <= (inputs(169)) or (inputs(251));
    layer0_outputs(11962) <= inputs(205);
    layer0_outputs(11963) <= not((inputs(96)) or (inputs(25)));
    layer0_outputs(11964) <= (inputs(152)) xor (inputs(53));
    layer0_outputs(11965) <= not((inputs(52)) or (inputs(193)));
    layer0_outputs(11966) <= (inputs(157)) xor (inputs(207));
    layer0_outputs(11967) <= inputs(170);
    layer0_outputs(11968) <= (inputs(169)) and not (inputs(71));
    layer0_outputs(11969) <= (inputs(95)) xor (inputs(106));
    layer0_outputs(11970) <= inputs(181);
    layer0_outputs(11971) <= not(inputs(194));
    layer0_outputs(11972) <= not(inputs(89)) or (inputs(153));
    layer0_outputs(11973) <= (inputs(139)) xor (inputs(0));
    layer0_outputs(11974) <= inputs(216);
    layer0_outputs(11975) <= (inputs(91)) and not (inputs(190));
    layer0_outputs(11976) <= (inputs(190)) and not (inputs(42));
    layer0_outputs(11977) <= not(inputs(175)) or (inputs(127));
    layer0_outputs(11978) <= (inputs(213)) and not (inputs(73));
    layer0_outputs(11979) <= (inputs(105)) xor (inputs(141));
    layer0_outputs(11980) <= not(inputs(122));
    layer0_outputs(11981) <= (inputs(135)) xor (inputs(195));
    layer0_outputs(11982) <= not(inputs(37));
    layer0_outputs(11983) <= not(inputs(217));
    layer0_outputs(11984) <= not((inputs(29)) and (inputs(129)));
    layer0_outputs(11985) <= (inputs(236)) and not (inputs(111));
    layer0_outputs(11986) <= '0';
    layer0_outputs(11987) <= not(inputs(216)) or (inputs(162));
    layer0_outputs(11988) <= not((inputs(103)) or (inputs(80)));
    layer0_outputs(11989) <= inputs(14);
    layer0_outputs(11990) <= inputs(24);
    layer0_outputs(11991) <= not(inputs(115));
    layer0_outputs(11992) <= inputs(231);
    layer0_outputs(11993) <= (inputs(201)) and not (inputs(116));
    layer0_outputs(11994) <= (inputs(63)) and not (inputs(190));
    layer0_outputs(11995) <= (inputs(24)) and not (inputs(108));
    layer0_outputs(11996) <= not(inputs(23));
    layer0_outputs(11997) <= (inputs(239)) or (inputs(108));
    layer0_outputs(11998) <= not(inputs(161)) or (inputs(58));
    layer0_outputs(11999) <= '0';
    layer0_outputs(12000) <= not((inputs(187)) xor (inputs(172)));
    layer0_outputs(12001) <= inputs(215);
    layer0_outputs(12002) <= not((inputs(15)) or (inputs(240)));
    layer0_outputs(12003) <= not((inputs(67)) xor (inputs(34)));
    layer0_outputs(12004) <= not(inputs(69));
    layer0_outputs(12005) <= (inputs(115)) xor (inputs(101));
    layer0_outputs(12006) <= (inputs(47)) and not (inputs(111));
    layer0_outputs(12007) <= not(inputs(86));
    layer0_outputs(12008) <= (inputs(28)) or (inputs(241));
    layer0_outputs(12009) <= not(inputs(165));
    layer0_outputs(12010) <= (inputs(91)) and not (inputs(146));
    layer0_outputs(12011) <= not(inputs(84));
    layer0_outputs(12012) <= not((inputs(208)) xor (inputs(40)));
    layer0_outputs(12013) <= not(inputs(40));
    layer0_outputs(12014) <= (inputs(84)) or (inputs(198));
    layer0_outputs(12015) <= not(inputs(107)) or (inputs(119));
    layer0_outputs(12016) <= (inputs(2)) or (inputs(11));
    layer0_outputs(12017) <= not(inputs(69));
    layer0_outputs(12018) <= (inputs(104)) and (inputs(240));
    layer0_outputs(12019) <= not(inputs(196)) or (inputs(206));
    layer0_outputs(12020) <= (inputs(174)) or (inputs(221));
    layer0_outputs(12021) <= inputs(220);
    layer0_outputs(12022) <= (inputs(168)) and not (inputs(173));
    layer0_outputs(12023) <= inputs(221);
    layer0_outputs(12024) <= not((inputs(80)) or (inputs(12)));
    layer0_outputs(12025) <= inputs(7);
    layer0_outputs(12026) <= (inputs(73)) xor (inputs(25));
    layer0_outputs(12027) <= (inputs(92)) or (inputs(138));
    layer0_outputs(12028) <= not((inputs(68)) xor (inputs(222)));
    layer0_outputs(12029) <= inputs(84);
    layer0_outputs(12030) <= inputs(169);
    layer0_outputs(12031) <= not(inputs(183)) or (inputs(131));
    layer0_outputs(12032) <= (inputs(183)) and not (inputs(31));
    layer0_outputs(12033) <= not(inputs(138)) or (inputs(253));
    layer0_outputs(12034) <= not((inputs(61)) or (inputs(20)));
    layer0_outputs(12035) <= not((inputs(163)) or (inputs(92)));
    layer0_outputs(12036) <= (inputs(196)) xor (inputs(211));
    layer0_outputs(12037) <= not(inputs(81));
    layer0_outputs(12038) <= inputs(64);
    layer0_outputs(12039) <= inputs(8);
    layer0_outputs(12040) <= not(inputs(228));
    layer0_outputs(12041) <= '0';
    layer0_outputs(12042) <= not((inputs(127)) or (inputs(81)));
    layer0_outputs(12043) <= not(inputs(73)) or (inputs(127));
    layer0_outputs(12044) <= inputs(135);
    layer0_outputs(12045) <= (inputs(140)) xor (inputs(242));
    layer0_outputs(12046) <= not(inputs(23));
    layer0_outputs(12047) <= (inputs(9)) or (inputs(184));
    layer0_outputs(12048) <= not((inputs(19)) or (inputs(186)));
    layer0_outputs(12049) <= not(inputs(29));
    layer0_outputs(12050) <= '1';
    layer0_outputs(12051) <= not((inputs(199)) xor (inputs(162)));
    layer0_outputs(12052) <= (inputs(187)) or (inputs(255));
    layer0_outputs(12053) <= (inputs(14)) or (inputs(30));
    layer0_outputs(12054) <= not(inputs(230));
    layer0_outputs(12055) <= not((inputs(126)) or (inputs(230)));
    layer0_outputs(12056) <= not(inputs(244));
    layer0_outputs(12057) <= (inputs(254)) or (inputs(251));
    layer0_outputs(12058) <= (inputs(228)) and (inputs(229));
    layer0_outputs(12059) <= '1';
    layer0_outputs(12060) <= not((inputs(218)) xor (inputs(145)));
    layer0_outputs(12061) <= (inputs(137)) and (inputs(219));
    layer0_outputs(12062) <= not(inputs(21)) or (inputs(111));
    layer0_outputs(12063) <= not((inputs(181)) or (inputs(157)));
    layer0_outputs(12064) <= not(inputs(46)) or (inputs(249));
    layer0_outputs(12065) <= not((inputs(100)) or (inputs(48)));
    layer0_outputs(12066) <= (inputs(118)) and not (inputs(217));
    layer0_outputs(12067) <= (inputs(39)) or (inputs(55));
    layer0_outputs(12068) <= not((inputs(196)) or (inputs(174)));
    layer0_outputs(12069) <= inputs(101);
    layer0_outputs(12070) <= (inputs(134)) or (inputs(219));
    layer0_outputs(12071) <= not(inputs(44)) or (inputs(126));
    layer0_outputs(12072) <= (inputs(181)) or (inputs(15));
    layer0_outputs(12073) <= not(inputs(124));
    layer0_outputs(12074) <= not((inputs(187)) xor (inputs(250)));
    layer0_outputs(12075) <= inputs(91);
    layer0_outputs(12076) <= (inputs(59)) xor (inputs(248));
    layer0_outputs(12077) <= (inputs(61)) or (inputs(98));
    layer0_outputs(12078) <= (inputs(5)) xor (inputs(109));
    layer0_outputs(12079) <= not(inputs(130));
    layer0_outputs(12080) <= not((inputs(138)) xor (inputs(34)));
    layer0_outputs(12081) <= inputs(76);
    layer0_outputs(12082) <= not((inputs(218)) or (inputs(191)));
    layer0_outputs(12083) <= inputs(209);
    layer0_outputs(12084) <= not(inputs(37));
    layer0_outputs(12085) <= (inputs(173)) and not (inputs(78));
    layer0_outputs(12086) <= not(inputs(217)) or (inputs(148));
    layer0_outputs(12087) <= not(inputs(37));
    layer0_outputs(12088) <= (inputs(42)) and not (inputs(177));
    layer0_outputs(12089) <= (inputs(68)) or (inputs(66));
    layer0_outputs(12090) <= not((inputs(7)) xor (inputs(225)));
    layer0_outputs(12091) <= not(inputs(228));
    layer0_outputs(12092) <= not(inputs(161)) or (inputs(237));
    layer0_outputs(12093) <= not(inputs(114));
    layer0_outputs(12094) <= (inputs(196)) xor (inputs(62));
    layer0_outputs(12095) <= not((inputs(132)) xor (inputs(86)));
    layer0_outputs(12096) <= (inputs(26)) xor (inputs(11));
    layer0_outputs(12097) <= (inputs(199)) or (inputs(180));
    layer0_outputs(12098) <= not(inputs(11));
    layer0_outputs(12099) <= (inputs(154)) and not (inputs(65));
    layer0_outputs(12100) <= inputs(75);
    layer0_outputs(12101) <= '1';
    layer0_outputs(12102) <= inputs(181);
    layer0_outputs(12103) <= inputs(6);
    layer0_outputs(12104) <= not((inputs(227)) or (inputs(244)));
    layer0_outputs(12105) <= (inputs(130)) or (inputs(119));
    layer0_outputs(12106) <= not((inputs(223)) or (inputs(189)));
    layer0_outputs(12107) <= not((inputs(151)) xor (inputs(231)));
    layer0_outputs(12108) <= not(inputs(101)) or (inputs(162));
    layer0_outputs(12109) <= not(inputs(44)) or (inputs(88));
    layer0_outputs(12110) <= inputs(68);
    layer0_outputs(12111) <= inputs(142);
    layer0_outputs(12112) <= not(inputs(212));
    layer0_outputs(12113) <= not((inputs(85)) xor (inputs(251)));
    layer0_outputs(12114) <= not((inputs(184)) or (inputs(101)));
    layer0_outputs(12115) <= (inputs(103)) xor (inputs(146));
    layer0_outputs(12116) <= not(inputs(42));
    layer0_outputs(12117) <= not(inputs(125));
    layer0_outputs(12118) <= not((inputs(62)) or (inputs(45)));
    layer0_outputs(12119) <= (inputs(167)) or (inputs(60));
    layer0_outputs(12120) <= '1';
    layer0_outputs(12121) <= not(inputs(93)) or (inputs(102));
    layer0_outputs(12122) <= not(inputs(102));
    layer0_outputs(12123) <= inputs(24);
    layer0_outputs(12124) <= not(inputs(10)) or (inputs(31));
    layer0_outputs(12125) <= (inputs(36)) xor (inputs(155));
    layer0_outputs(12126) <= not(inputs(207)) or (inputs(220));
    layer0_outputs(12127) <= not(inputs(158)) or (inputs(152));
    layer0_outputs(12128) <= (inputs(107)) xor (inputs(45));
    layer0_outputs(12129) <= not(inputs(219));
    layer0_outputs(12130) <= not(inputs(57));
    layer0_outputs(12131) <= (inputs(53)) or (inputs(95));
    layer0_outputs(12132) <= inputs(39);
    layer0_outputs(12133) <= not((inputs(155)) xor (inputs(10)));
    layer0_outputs(12134) <= not(inputs(105)) or (inputs(55));
    layer0_outputs(12135) <= not((inputs(195)) xor (inputs(76)));
    layer0_outputs(12136) <= not((inputs(112)) xor (inputs(99)));
    layer0_outputs(12137) <= not(inputs(255));
    layer0_outputs(12138) <= not((inputs(44)) or (inputs(108)));
    layer0_outputs(12139) <= not(inputs(36)) or (inputs(251));
    layer0_outputs(12140) <= not((inputs(120)) or (inputs(191)));
    layer0_outputs(12141) <= inputs(82);
    layer0_outputs(12142) <= (inputs(111)) or (inputs(77));
    layer0_outputs(12143) <= not((inputs(123)) or (inputs(252)));
    layer0_outputs(12144) <= not((inputs(176)) xor (inputs(81)));
    layer0_outputs(12145) <= not((inputs(245)) or (inputs(235)));
    layer0_outputs(12146) <= not((inputs(5)) or (inputs(2)));
    layer0_outputs(12147) <= (inputs(174)) and not (inputs(111));
    layer0_outputs(12148) <= inputs(90);
    layer0_outputs(12149) <= inputs(38);
    layer0_outputs(12150) <= not(inputs(152)) or (inputs(96));
    layer0_outputs(12151) <= (inputs(236)) or (inputs(224));
    layer0_outputs(12152) <= inputs(218);
    layer0_outputs(12153) <= (inputs(33)) and (inputs(152));
    layer0_outputs(12154) <= (inputs(177)) xor (inputs(197));
    layer0_outputs(12155) <= not(inputs(115));
    layer0_outputs(12156) <= (inputs(4)) xor (inputs(192));
    layer0_outputs(12157) <= not(inputs(88));
    layer0_outputs(12158) <= (inputs(222)) and (inputs(97));
    layer0_outputs(12159) <= not(inputs(173)) or (inputs(151));
    layer0_outputs(12160) <= not(inputs(117));
    layer0_outputs(12161) <= not((inputs(17)) or (inputs(32)));
    layer0_outputs(12162) <= not(inputs(216)) or (inputs(113));
    layer0_outputs(12163) <= inputs(194);
    layer0_outputs(12164) <= not((inputs(217)) or (inputs(95)));
    layer0_outputs(12165) <= (inputs(186)) or (inputs(160));
    layer0_outputs(12166) <= not((inputs(94)) and (inputs(18)));
    layer0_outputs(12167) <= not((inputs(184)) or (inputs(254)));
    layer0_outputs(12168) <= not(inputs(20)) or (inputs(207));
    layer0_outputs(12169) <= inputs(222);
    layer0_outputs(12170) <= '1';
    layer0_outputs(12171) <= not(inputs(85));
    layer0_outputs(12172) <= not(inputs(145)) or (inputs(224));
    layer0_outputs(12173) <= (inputs(197)) or (inputs(235));
    layer0_outputs(12174) <= (inputs(198)) xor (inputs(217));
    layer0_outputs(12175) <= not(inputs(219));
    layer0_outputs(12176) <= not(inputs(94));
    layer0_outputs(12177) <= inputs(120);
    layer0_outputs(12178) <= (inputs(194)) or (inputs(178));
    layer0_outputs(12179) <= not((inputs(62)) xor (inputs(219)));
    layer0_outputs(12180) <= (inputs(156)) or (inputs(26));
    layer0_outputs(12181) <= not(inputs(25));
    layer0_outputs(12182) <= not((inputs(177)) xor (inputs(17)));
    layer0_outputs(12183) <= (inputs(232)) and not (inputs(48));
    layer0_outputs(12184) <= not((inputs(60)) or (inputs(217)));
    layer0_outputs(12185) <= not(inputs(169));
    layer0_outputs(12186) <= (inputs(22)) and not (inputs(221));
    layer0_outputs(12187) <= not(inputs(179));
    layer0_outputs(12188) <= not(inputs(10));
    layer0_outputs(12189) <= (inputs(255)) and not (inputs(10));
    layer0_outputs(12190) <= not(inputs(228));
    layer0_outputs(12191) <= (inputs(25)) and not (inputs(69));
    layer0_outputs(12192) <= not((inputs(192)) and (inputs(196)));
    layer0_outputs(12193) <= inputs(65);
    layer0_outputs(12194) <= not((inputs(196)) xor (inputs(54)));
    layer0_outputs(12195) <= (inputs(149)) xor (inputs(190));
    layer0_outputs(12196) <= inputs(101);
    layer0_outputs(12197) <= (inputs(44)) and not (inputs(54));
    layer0_outputs(12198) <= (inputs(112)) or (inputs(51));
    layer0_outputs(12199) <= not((inputs(179)) and (inputs(164)));
    layer0_outputs(12200) <= inputs(195);
    layer0_outputs(12201) <= not((inputs(23)) and (inputs(166)));
    layer0_outputs(12202) <= (inputs(247)) xor (inputs(159));
    layer0_outputs(12203) <= not(inputs(15));
    layer0_outputs(12204) <= inputs(62);
    layer0_outputs(12205) <= not((inputs(18)) or (inputs(4)));
    layer0_outputs(12206) <= inputs(211);
    layer0_outputs(12207) <= (inputs(63)) or (inputs(85));
    layer0_outputs(12208) <= not(inputs(92));
    layer0_outputs(12209) <= not((inputs(88)) xor (inputs(13)));
    layer0_outputs(12210) <= not(inputs(179)) or (inputs(98));
    layer0_outputs(12211) <= not(inputs(21)) or (inputs(115));
    layer0_outputs(12212) <= inputs(167);
    layer0_outputs(12213) <= not((inputs(142)) xor (inputs(107)));
    layer0_outputs(12214) <= inputs(10);
    layer0_outputs(12215) <= not(inputs(114));
    layer0_outputs(12216) <= (inputs(87)) xor (inputs(37));
    layer0_outputs(12217) <= (inputs(98)) and not (inputs(48));
    layer0_outputs(12218) <= (inputs(229)) or (inputs(246));
    layer0_outputs(12219) <= inputs(118);
    layer0_outputs(12220) <= not(inputs(142));
    layer0_outputs(12221) <= not((inputs(33)) or (inputs(37)));
    layer0_outputs(12222) <= inputs(66);
    layer0_outputs(12223) <= (inputs(97)) or (inputs(30));
    layer0_outputs(12224) <= (inputs(112)) or (inputs(85));
    layer0_outputs(12225) <= (inputs(131)) and not (inputs(0));
    layer0_outputs(12226) <= not((inputs(156)) or (inputs(29)));
    layer0_outputs(12227) <= not(inputs(17));
    layer0_outputs(12228) <= not(inputs(84));
    layer0_outputs(12229) <= inputs(25);
    layer0_outputs(12230) <= (inputs(36)) xor (inputs(108));
    layer0_outputs(12231) <= not(inputs(117));
    layer0_outputs(12232) <= not((inputs(213)) and (inputs(165)));
    layer0_outputs(12233) <= not(inputs(199));
    layer0_outputs(12234) <= not((inputs(210)) or (inputs(135)));
    layer0_outputs(12235) <= '0';
    layer0_outputs(12236) <= not(inputs(11)) or (inputs(207));
    layer0_outputs(12237) <= not(inputs(133)) or (inputs(134));
    layer0_outputs(12238) <= (inputs(166)) or (inputs(66));
    layer0_outputs(12239) <= (inputs(60)) and not (inputs(241));
    layer0_outputs(12240) <= inputs(177);
    layer0_outputs(12241) <= not(inputs(198)) or (inputs(2));
    layer0_outputs(12242) <= inputs(248);
    layer0_outputs(12243) <= not(inputs(246));
    layer0_outputs(12244) <= not(inputs(195));
    layer0_outputs(12245) <= not((inputs(149)) xor (inputs(28)));
    layer0_outputs(12246) <= not(inputs(235));
    layer0_outputs(12247) <= not(inputs(214));
    layer0_outputs(12248) <= not(inputs(185));
    layer0_outputs(12249) <= (inputs(10)) or (inputs(206));
    layer0_outputs(12250) <= inputs(164);
    layer0_outputs(12251) <= inputs(246);
    layer0_outputs(12252) <= not((inputs(204)) and (inputs(219)));
    layer0_outputs(12253) <= not(inputs(146)) or (inputs(240));
    layer0_outputs(12254) <= not((inputs(104)) and (inputs(224)));
    layer0_outputs(12255) <= not(inputs(255));
    layer0_outputs(12256) <= (inputs(199)) xor (inputs(0));
    layer0_outputs(12257) <= not((inputs(59)) and (inputs(140)));
    layer0_outputs(12258) <= not((inputs(41)) and (inputs(36)));
    layer0_outputs(12259) <= not(inputs(79));
    layer0_outputs(12260) <= inputs(222);
    layer0_outputs(12261) <= (inputs(160)) or (inputs(221));
    layer0_outputs(12262) <= inputs(36);
    layer0_outputs(12263) <= inputs(249);
    layer0_outputs(12264) <= inputs(144);
    layer0_outputs(12265) <= not(inputs(104)) or (inputs(195));
    layer0_outputs(12266) <= not((inputs(219)) or (inputs(128)));
    layer0_outputs(12267) <= not((inputs(111)) or (inputs(2)));
    layer0_outputs(12268) <= (inputs(77)) and (inputs(243));
    layer0_outputs(12269) <= not((inputs(166)) or (inputs(216)));
    layer0_outputs(12270) <= not(inputs(37)) or (inputs(225));
    layer0_outputs(12271) <= '1';
    layer0_outputs(12272) <= not(inputs(229));
    layer0_outputs(12273) <= not(inputs(234)) or (inputs(126));
    layer0_outputs(12274) <= (inputs(191)) and (inputs(174));
    layer0_outputs(12275) <= not((inputs(246)) or (inputs(221)));
    layer0_outputs(12276) <= not((inputs(183)) xor (inputs(100)));
    layer0_outputs(12277) <= not(inputs(221));
    layer0_outputs(12278) <= (inputs(35)) or (inputs(22));
    layer0_outputs(12279) <= not(inputs(80));
    layer0_outputs(12280) <= not(inputs(125));
    layer0_outputs(12281) <= not(inputs(122)) or (inputs(77));
    layer0_outputs(12282) <= not((inputs(143)) xor (inputs(33)));
    layer0_outputs(12283) <= not(inputs(105));
    layer0_outputs(12284) <= (inputs(15)) and not (inputs(206));
    layer0_outputs(12285) <= not((inputs(51)) xor (inputs(53)));
    layer0_outputs(12286) <= not(inputs(165)) or (inputs(198));
    layer0_outputs(12287) <= (inputs(99)) and not (inputs(127));
    layer0_outputs(12288) <= (inputs(29)) and not (inputs(63));
    layer0_outputs(12289) <= not((inputs(116)) xor (inputs(157)));
    layer0_outputs(12290) <= inputs(104);
    layer0_outputs(12291) <= not(inputs(20)) or (inputs(205));
    layer0_outputs(12292) <= not((inputs(195)) or (inputs(83)));
    layer0_outputs(12293) <= (inputs(201)) and not (inputs(1));
    layer0_outputs(12294) <= inputs(125);
    layer0_outputs(12295) <= not((inputs(43)) or (inputs(140)));
    layer0_outputs(12296) <= (inputs(8)) or (inputs(76));
    layer0_outputs(12297) <= (inputs(21)) or (inputs(136));
    layer0_outputs(12298) <= (inputs(10)) or (inputs(212));
    layer0_outputs(12299) <= not(inputs(236)) or (inputs(1));
    layer0_outputs(12300) <= not((inputs(119)) xor (inputs(178)));
    layer0_outputs(12301) <= not(inputs(114));
    layer0_outputs(12302) <= (inputs(28)) and not (inputs(225));
    layer0_outputs(12303) <= not((inputs(62)) or (inputs(187)));
    layer0_outputs(12304) <= not(inputs(165)) or (inputs(3));
    layer0_outputs(12305) <= inputs(242);
    layer0_outputs(12306) <= inputs(129);
    layer0_outputs(12307) <= not((inputs(205)) xor (inputs(253)));
    layer0_outputs(12308) <= not((inputs(150)) or (inputs(252)));
    layer0_outputs(12309) <= inputs(194);
    layer0_outputs(12310) <= not((inputs(78)) or (inputs(248)));
    layer0_outputs(12311) <= inputs(217);
    layer0_outputs(12312) <= inputs(25);
    layer0_outputs(12313) <= '0';
    layer0_outputs(12314) <= not((inputs(227)) or (inputs(213)));
    layer0_outputs(12315) <= (inputs(189)) xor (inputs(38));
    layer0_outputs(12316) <= inputs(172);
    layer0_outputs(12317) <= not(inputs(164)) or (inputs(127));
    layer0_outputs(12318) <= not((inputs(209)) or (inputs(244)));
    layer0_outputs(12319) <= (inputs(79)) or (inputs(78));
    layer0_outputs(12320) <= not((inputs(208)) xor (inputs(149)));
    layer0_outputs(12321) <= not((inputs(81)) or (inputs(185)));
    layer0_outputs(12322) <= (inputs(93)) or (inputs(215));
    layer0_outputs(12323) <= inputs(125);
    layer0_outputs(12324) <= not((inputs(182)) or (inputs(138)));
    layer0_outputs(12325) <= not(inputs(121));
    layer0_outputs(12326) <= (inputs(77)) and not (inputs(237));
    layer0_outputs(12327) <= (inputs(131)) xor (inputs(19));
    layer0_outputs(12328) <= (inputs(117)) and not (inputs(184));
    layer0_outputs(12329) <= not(inputs(244));
    layer0_outputs(12330) <= (inputs(1)) and (inputs(124));
    layer0_outputs(12331) <= inputs(73);
    layer0_outputs(12332) <= inputs(9);
    layer0_outputs(12333) <= inputs(57);
    layer0_outputs(12334) <= inputs(35);
    layer0_outputs(12335) <= not(inputs(183));
    layer0_outputs(12336) <= not((inputs(109)) and (inputs(18)));
    layer0_outputs(12337) <= (inputs(163)) xor (inputs(165));
    layer0_outputs(12338) <= (inputs(124)) xor (inputs(133));
    layer0_outputs(12339) <= (inputs(142)) and not (inputs(80));
    layer0_outputs(12340) <= not(inputs(96));
    layer0_outputs(12341) <= inputs(114);
    layer0_outputs(12342) <= not(inputs(178)) or (inputs(74));
    layer0_outputs(12343) <= not(inputs(94));
    layer0_outputs(12344) <= inputs(251);
    layer0_outputs(12345) <= (inputs(152)) and (inputs(2));
    layer0_outputs(12346) <= (inputs(72)) xor (inputs(29));
    layer0_outputs(12347) <= not(inputs(110)) or (inputs(229));
    layer0_outputs(12348) <= '0';
    layer0_outputs(12349) <= not((inputs(146)) xor (inputs(187)));
    layer0_outputs(12350) <= (inputs(92)) xor (inputs(119));
    layer0_outputs(12351) <= inputs(130);
    layer0_outputs(12352) <= (inputs(187)) and not (inputs(46));
    layer0_outputs(12353) <= (inputs(30)) xor (inputs(178));
    layer0_outputs(12354) <= inputs(0);
    layer0_outputs(12355) <= not((inputs(93)) or (inputs(251)));
    layer0_outputs(12356) <= not((inputs(164)) or (inputs(197)));
    layer0_outputs(12357) <= (inputs(138)) and not (inputs(159));
    layer0_outputs(12358) <= (inputs(115)) and not (inputs(89));
    layer0_outputs(12359) <= (inputs(165)) and not (inputs(115));
    layer0_outputs(12360) <= inputs(107);
    layer0_outputs(12361) <= (inputs(222)) or (inputs(246));
    layer0_outputs(12362) <= (inputs(105)) and not (inputs(210));
    layer0_outputs(12363) <= inputs(1);
    layer0_outputs(12364) <= (inputs(32)) xor (inputs(187));
    layer0_outputs(12365) <= not(inputs(210));
    layer0_outputs(12366) <= (inputs(10)) and not (inputs(179));
    layer0_outputs(12367) <= (inputs(65)) or (inputs(237));
    layer0_outputs(12368) <= inputs(148);
    layer0_outputs(12369) <= not((inputs(61)) xor (inputs(59)));
    layer0_outputs(12370) <= not(inputs(247));
    layer0_outputs(12371) <= not((inputs(183)) and (inputs(169)));
    layer0_outputs(12372) <= (inputs(252)) or (inputs(218));
    layer0_outputs(12373) <= (inputs(97)) or (inputs(155));
    layer0_outputs(12374) <= not((inputs(179)) or (inputs(219)));
    layer0_outputs(12375) <= inputs(67);
    layer0_outputs(12376) <= (inputs(255)) xor (inputs(53));
    layer0_outputs(12377) <= (inputs(104)) and not (inputs(200));
    layer0_outputs(12378) <= inputs(168);
    layer0_outputs(12379) <= (inputs(70)) xor (inputs(118));
    layer0_outputs(12380) <= (inputs(41)) and not (inputs(186));
    layer0_outputs(12381) <= not(inputs(74)) or (inputs(31));
    layer0_outputs(12382) <= not(inputs(100)) or (inputs(121));
    layer0_outputs(12383) <= (inputs(99)) xor (inputs(31));
    layer0_outputs(12384) <= (inputs(178)) or (inputs(214));
    layer0_outputs(12385) <= inputs(101);
    layer0_outputs(12386) <= (inputs(81)) or (inputs(5));
    layer0_outputs(12387) <= (inputs(1)) xor (inputs(137));
    layer0_outputs(12388) <= not(inputs(225));
    layer0_outputs(12389) <= (inputs(94)) and not (inputs(33));
    layer0_outputs(12390) <= not(inputs(89));
    layer0_outputs(12391) <= inputs(140);
    layer0_outputs(12392) <= not((inputs(81)) and (inputs(20)));
    layer0_outputs(12393) <= not((inputs(231)) xor (inputs(222)));
    layer0_outputs(12394) <= inputs(129);
    layer0_outputs(12395) <= (inputs(62)) xor (inputs(126));
    layer0_outputs(12396) <= inputs(104);
    layer0_outputs(12397) <= not(inputs(47));
    layer0_outputs(12398) <= (inputs(163)) and not (inputs(62));
    layer0_outputs(12399) <= not(inputs(205)) or (inputs(162));
    layer0_outputs(12400) <= inputs(216);
    layer0_outputs(12401) <= not((inputs(183)) and (inputs(179)));
    layer0_outputs(12402) <= not(inputs(130));
    layer0_outputs(12403) <= not(inputs(42)) or (inputs(65));
    layer0_outputs(12404) <= inputs(190);
    layer0_outputs(12405) <= (inputs(238)) xor (inputs(58));
    layer0_outputs(12406) <= not((inputs(39)) or (inputs(27)));
    layer0_outputs(12407) <= not(inputs(94));
    layer0_outputs(12408) <= inputs(41);
    layer0_outputs(12409) <= inputs(157);
    layer0_outputs(12410) <= not(inputs(92));
    layer0_outputs(12411) <= (inputs(155)) and not (inputs(176));
    layer0_outputs(12412) <= not(inputs(172));
    layer0_outputs(12413) <= (inputs(5)) xor (inputs(220));
    layer0_outputs(12414) <= inputs(236);
    layer0_outputs(12415) <= inputs(85);
    layer0_outputs(12416) <= not(inputs(220));
    layer0_outputs(12417) <= not((inputs(99)) or (inputs(78)));
    layer0_outputs(12418) <= '0';
    layer0_outputs(12419) <= not(inputs(135)) or (inputs(28));
    layer0_outputs(12420) <= not((inputs(108)) xor (inputs(120)));
    layer0_outputs(12421) <= not(inputs(45));
    layer0_outputs(12422) <= (inputs(129)) and not (inputs(0));
    layer0_outputs(12423) <= (inputs(236)) or (inputs(62));
    layer0_outputs(12424) <= (inputs(247)) and not (inputs(241));
    layer0_outputs(12425) <= not((inputs(118)) xor (inputs(54)));
    layer0_outputs(12426) <= inputs(162);
    layer0_outputs(12427) <= '0';
    layer0_outputs(12428) <= not((inputs(28)) xor (inputs(142)));
    layer0_outputs(12429) <= not((inputs(47)) or (inputs(90)));
    layer0_outputs(12430) <= inputs(123);
    layer0_outputs(12431) <= (inputs(241)) or (inputs(235));
    layer0_outputs(12432) <= not(inputs(180));
    layer0_outputs(12433) <= not(inputs(4)) or (inputs(114));
    layer0_outputs(12434) <= (inputs(154)) and not (inputs(79));
    layer0_outputs(12435) <= not((inputs(146)) xor (inputs(79)));
    layer0_outputs(12436) <= not(inputs(85)) or (inputs(142));
    layer0_outputs(12437) <= not((inputs(134)) xor (inputs(118)));
    layer0_outputs(12438) <= (inputs(222)) xor (inputs(15));
    layer0_outputs(12439) <= (inputs(241)) or (inputs(223));
    layer0_outputs(12440) <= not(inputs(189));
    layer0_outputs(12441) <= (inputs(103)) xor (inputs(58));
    layer0_outputs(12442) <= inputs(234);
    layer0_outputs(12443) <= not((inputs(227)) or (inputs(239)));
    layer0_outputs(12444) <= not((inputs(156)) xor (inputs(236)));
    layer0_outputs(12445) <= (inputs(90)) and not (inputs(179));
    layer0_outputs(12446) <= not(inputs(107)) or (inputs(226));
    layer0_outputs(12447) <= (inputs(73)) or (inputs(19));
    layer0_outputs(12448) <= not(inputs(169));
    layer0_outputs(12449) <= inputs(77);
    layer0_outputs(12450) <= not((inputs(174)) or (inputs(36)));
    layer0_outputs(12451) <= not(inputs(118)) or (inputs(255));
    layer0_outputs(12452) <= not((inputs(64)) and (inputs(187)));
    layer0_outputs(12453) <= inputs(92);
    layer0_outputs(12454) <= not(inputs(11));
    layer0_outputs(12455) <= not(inputs(114));
    layer0_outputs(12456) <= not(inputs(185)) or (inputs(205));
    layer0_outputs(12457) <= (inputs(42)) and not (inputs(220));
    layer0_outputs(12458) <= not(inputs(24));
    layer0_outputs(12459) <= not(inputs(217)) or (inputs(90));
    layer0_outputs(12460) <= (inputs(137)) xor (inputs(59));
    layer0_outputs(12461) <= (inputs(173)) and not (inputs(46));
    layer0_outputs(12462) <= inputs(57);
    layer0_outputs(12463) <= (inputs(115)) and not (inputs(18));
    layer0_outputs(12464) <= not(inputs(74)) or (inputs(243));
    layer0_outputs(12465) <= (inputs(209)) and not (inputs(249));
    layer0_outputs(12466) <= not((inputs(71)) xor (inputs(190)));
    layer0_outputs(12467) <= (inputs(75)) and not (inputs(235));
    layer0_outputs(12468) <= not(inputs(231));
    layer0_outputs(12469) <= not((inputs(244)) or (inputs(94)));
    layer0_outputs(12470) <= not(inputs(0));
    layer0_outputs(12471) <= not((inputs(213)) or (inputs(191)));
    layer0_outputs(12472) <= not((inputs(128)) or (inputs(52)));
    layer0_outputs(12473) <= not(inputs(178));
    layer0_outputs(12474) <= not(inputs(8));
    layer0_outputs(12475) <= not((inputs(135)) or (inputs(56)));
    layer0_outputs(12476) <= not(inputs(101));
    layer0_outputs(12477) <= inputs(20);
    layer0_outputs(12478) <= not((inputs(172)) or (inputs(186)));
    layer0_outputs(12479) <= not((inputs(109)) xor (inputs(106)));
    layer0_outputs(12480) <= not(inputs(37)) or (inputs(161));
    layer0_outputs(12481) <= not(inputs(98)) or (inputs(252));
    layer0_outputs(12482) <= inputs(0);
    layer0_outputs(12483) <= not(inputs(102)) or (inputs(240));
    layer0_outputs(12484) <= not((inputs(43)) or (inputs(252)));
    layer0_outputs(12485) <= not(inputs(229));
    layer0_outputs(12486) <= not((inputs(68)) or (inputs(12)));
    layer0_outputs(12487) <= not((inputs(23)) xor (inputs(81)));
    layer0_outputs(12488) <= not(inputs(148)) or (inputs(96));
    layer0_outputs(12489) <= inputs(101);
    layer0_outputs(12490) <= not(inputs(228)) or (inputs(29));
    layer0_outputs(12491) <= inputs(107);
    layer0_outputs(12492) <= not(inputs(7));
    layer0_outputs(12493) <= not((inputs(175)) xor (inputs(6)));
    layer0_outputs(12494) <= not(inputs(224)) or (inputs(49));
    layer0_outputs(12495) <= (inputs(168)) xor (inputs(32));
    layer0_outputs(12496) <= not(inputs(85)) or (inputs(199));
    layer0_outputs(12497) <= not(inputs(104)) or (inputs(239));
    layer0_outputs(12498) <= not(inputs(122)) or (inputs(222));
    layer0_outputs(12499) <= '1';
    layer0_outputs(12500) <= not(inputs(116));
    layer0_outputs(12501) <= (inputs(31)) and (inputs(220));
    layer0_outputs(12502) <= (inputs(160)) xor (inputs(14));
    layer0_outputs(12503) <= not((inputs(251)) or (inputs(25)));
    layer0_outputs(12504) <= (inputs(255)) or (inputs(185));
    layer0_outputs(12505) <= inputs(36);
    layer0_outputs(12506) <= (inputs(133)) xor (inputs(68));
    layer0_outputs(12507) <= (inputs(70)) and (inputs(27));
    layer0_outputs(12508) <= not((inputs(18)) or (inputs(43)));
    layer0_outputs(12509) <= not((inputs(231)) xor (inputs(214)));
    layer0_outputs(12510) <= not(inputs(91));
    layer0_outputs(12511) <= not(inputs(80)) or (inputs(212));
    layer0_outputs(12512) <= not((inputs(245)) xor (inputs(4)));
    layer0_outputs(12513) <= not(inputs(18)) or (inputs(207));
    layer0_outputs(12514) <= not((inputs(193)) xor (inputs(67)));
    layer0_outputs(12515) <= (inputs(92)) or (inputs(47));
    layer0_outputs(12516) <= '1';
    layer0_outputs(12517) <= not(inputs(36)) or (inputs(242));
    layer0_outputs(12518) <= not(inputs(29)) or (inputs(48));
    layer0_outputs(12519) <= inputs(35);
    layer0_outputs(12520) <= not((inputs(158)) xor (inputs(124)));
    layer0_outputs(12521) <= (inputs(28)) xor (inputs(61));
    layer0_outputs(12522) <= not((inputs(16)) xor (inputs(249)));
    layer0_outputs(12523) <= not(inputs(199));
    layer0_outputs(12524) <= not((inputs(96)) and (inputs(31)));
    layer0_outputs(12525) <= not((inputs(54)) or (inputs(12)));
    layer0_outputs(12526) <= (inputs(133)) or (inputs(225));
    layer0_outputs(12527) <= (inputs(250)) or (inputs(9));
    layer0_outputs(12528) <= not(inputs(68));
    layer0_outputs(12529) <= (inputs(104)) and not (inputs(91));
    layer0_outputs(12530) <= inputs(247);
    layer0_outputs(12531) <= (inputs(113)) or (inputs(79));
    layer0_outputs(12532) <= (inputs(50)) and not (inputs(56));
    layer0_outputs(12533) <= not((inputs(254)) xor (inputs(74)));
    layer0_outputs(12534) <= not(inputs(248));
    layer0_outputs(12535) <= not((inputs(246)) or (inputs(242)));
    layer0_outputs(12536) <= inputs(1);
    layer0_outputs(12537) <= (inputs(109)) and not (inputs(238));
    layer0_outputs(12538) <= inputs(157);
    layer0_outputs(12539) <= not((inputs(34)) xor (inputs(205)));
    layer0_outputs(12540) <= '1';
    layer0_outputs(12541) <= inputs(230);
    layer0_outputs(12542) <= not(inputs(151));
    layer0_outputs(12543) <= not((inputs(171)) or (inputs(192)));
    layer0_outputs(12544) <= not((inputs(142)) and (inputs(142)));
    layer0_outputs(12545) <= (inputs(74)) xor (inputs(247));
    layer0_outputs(12546) <= not((inputs(102)) xor (inputs(117)));
    layer0_outputs(12547) <= inputs(123);
    layer0_outputs(12548) <= inputs(22);
    layer0_outputs(12549) <= not(inputs(9));
    layer0_outputs(12550) <= inputs(62);
    layer0_outputs(12551) <= not((inputs(240)) or (inputs(65)));
    layer0_outputs(12552) <= not((inputs(201)) and (inputs(242)));
    layer0_outputs(12553) <= not((inputs(47)) xor (inputs(48)));
    layer0_outputs(12554) <= not(inputs(129));
    layer0_outputs(12555) <= inputs(17);
    layer0_outputs(12556) <= inputs(116);
    layer0_outputs(12557) <= not(inputs(173)) or (inputs(23));
    layer0_outputs(12558) <= (inputs(38)) xor (inputs(127));
    layer0_outputs(12559) <= not((inputs(153)) and (inputs(240)));
    layer0_outputs(12560) <= not(inputs(61));
    layer0_outputs(12561) <= not((inputs(4)) xor (inputs(79)));
    layer0_outputs(12562) <= not((inputs(140)) or (inputs(161)));
    layer0_outputs(12563) <= (inputs(151)) xor (inputs(234));
    layer0_outputs(12564) <= not(inputs(190)) or (inputs(200));
    layer0_outputs(12565) <= not((inputs(46)) xor (inputs(49)));
    layer0_outputs(12566) <= not((inputs(190)) xor (inputs(50)));
    layer0_outputs(12567) <= (inputs(3)) or (inputs(39));
    layer0_outputs(12568) <= not((inputs(226)) or (inputs(177)));
    layer0_outputs(12569) <= (inputs(5)) xor (inputs(76));
    layer0_outputs(12570) <= (inputs(123)) or (inputs(28));
    layer0_outputs(12571) <= not((inputs(26)) xor (inputs(88)));
    layer0_outputs(12572) <= inputs(181);
    layer0_outputs(12573) <= '1';
    layer0_outputs(12574) <= (inputs(188)) and not (inputs(114));
    layer0_outputs(12575) <= inputs(188);
    layer0_outputs(12576) <= not((inputs(217)) and (inputs(85)));
    layer0_outputs(12577) <= inputs(67);
    layer0_outputs(12578) <= (inputs(67)) or (inputs(149));
    layer0_outputs(12579) <= (inputs(98)) and not (inputs(57));
    layer0_outputs(12580) <= not((inputs(163)) or (inputs(182)));
    layer0_outputs(12581) <= not((inputs(231)) xor (inputs(48)));
    layer0_outputs(12582) <= (inputs(204)) xor (inputs(110));
    layer0_outputs(12583) <= (inputs(68)) and not (inputs(144));
    layer0_outputs(12584) <= (inputs(69)) or (inputs(189));
    layer0_outputs(12585) <= (inputs(147)) or (inputs(96));
    layer0_outputs(12586) <= not(inputs(164));
    layer0_outputs(12587) <= not((inputs(214)) or (inputs(8)));
    layer0_outputs(12588) <= (inputs(12)) xor (inputs(71));
    layer0_outputs(12589) <= not(inputs(181));
    layer0_outputs(12590) <= (inputs(197)) or (inputs(144));
    layer0_outputs(12591) <= not(inputs(233)) or (inputs(111));
    layer0_outputs(12592) <= inputs(105);
    layer0_outputs(12593) <= (inputs(139)) and not (inputs(229));
    layer0_outputs(12594) <= (inputs(104)) and not (inputs(157));
    layer0_outputs(12595) <= not(inputs(163));
    layer0_outputs(12596) <= not((inputs(187)) xor (inputs(229)));
    layer0_outputs(12597) <= not(inputs(58));
    layer0_outputs(12598) <= (inputs(251)) xor (inputs(73));
    layer0_outputs(12599) <= inputs(180);
    layer0_outputs(12600) <= not((inputs(24)) xor (inputs(156)));
    layer0_outputs(12601) <= (inputs(92)) and not (inputs(223));
    layer0_outputs(12602) <= (inputs(53)) xor (inputs(66));
    layer0_outputs(12603) <= not(inputs(249));
    layer0_outputs(12604) <= (inputs(10)) and (inputs(159));
    layer0_outputs(12605) <= (inputs(95)) xor (inputs(179));
    layer0_outputs(12606) <= inputs(199);
    layer0_outputs(12607) <= inputs(101);
    layer0_outputs(12608) <= '1';
    layer0_outputs(12609) <= (inputs(103)) xor (inputs(133));
    layer0_outputs(12610) <= (inputs(181)) and (inputs(70));
    layer0_outputs(12611) <= not(inputs(144));
    layer0_outputs(12612) <= not(inputs(22));
    layer0_outputs(12613) <= not((inputs(221)) xor (inputs(51)));
    layer0_outputs(12614) <= (inputs(130)) xor (inputs(102));
    layer0_outputs(12615) <= not(inputs(8));
    layer0_outputs(12616) <= '1';
    layer0_outputs(12617) <= inputs(164);
    layer0_outputs(12618) <= (inputs(233)) or (inputs(61));
    layer0_outputs(12619) <= (inputs(251)) xor (inputs(122));
    layer0_outputs(12620) <= (inputs(101)) and not (inputs(80));
    layer0_outputs(12621) <= not(inputs(220)) or (inputs(87));
    layer0_outputs(12622) <= (inputs(218)) xor (inputs(1));
    layer0_outputs(12623) <= not(inputs(247));
    layer0_outputs(12624) <= not(inputs(101)) or (inputs(105));
    layer0_outputs(12625) <= (inputs(133)) and not (inputs(252));
    layer0_outputs(12626) <= not(inputs(69));
    layer0_outputs(12627) <= not((inputs(35)) and (inputs(125)));
    layer0_outputs(12628) <= inputs(22);
    layer0_outputs(12629) <= not(inputs(183));
    layer0_outputs(12630) <= not((inputs(16)) or (inputs(89)));
    layer0_outputs(12631) <= not(inputs(248)) or (inputs(128));
    layer0_outputs(12632) <= not((inputs(246)) xor (inputs(114)));
    layer0_outputs(12633) <= not(inputs(17)) or (inputs(3));
    layer0_outputs(12634) <= not((inputs(168)) or (inputs(247)));
    layer0_outputs(12635) <= not((inputs(129)) xor (inputs(119)));
    layer0_outputs(12636) <= (inputs(69)) or (inputs(70));
    layer0_outputs(12637) <= (inputs(105)) xor (inputs(233));
    layer0_outputs(12638) <= (inputs(251)) or (inputs(143));
    layer0_outputs(12639) <= not((inputs(37)) or (inputs(31)));
    layer0_outputs(12640) <= inputs(93);
    layer0_outputs(12641) <= not(inputs(90));
    layer0_outputs(12642) <= (inputs(15)) or (inputs(100));
    layer0_outputs(12643) <= inputs(116);
    layer0_outputs(12644) <= not(inputs(121)) or (inputs(187));
    layer0_outputs(12645) <= not(inputs(102));
    layer0_outputs(12646) <= inputs(193);
    layer0_outputs(12647) <= (inputs(236)) and not (inputs(208));
    layer0_outputs(12648) <= not((inputs(122)) xor (inputs(1)));
    layer0_outputs(12649) <= not((inputs(177)) xor (inputs(211)));
    layer0_outputs(12650) <= not(inputs(59));
    layer0_outputs(12651) <= inputs(208);
    layer0_outputs(12652) <= not((inputs(61)) and (inputs(137)));
    layer0_outputs(12653) <= not((inputs(93)) or (inputs(179)));
    layer0_outputs(12654) <= not(inputs(169));
    layer0_outputs(12655) <= inputs(247);
    layer0_outputs(12656) <= inputs(181);
    layer0_outputs(12657) <= '1';
    layer0_outputs(12658) <= not(inputs(167));
    layer0_outputs(12659) <= (inputs(98)) or (inputs(63));
    layer0_outputs(12660) <= not(inputs(113));
    layer0_outputs(12661) <= not((inputs(77)) and (inputs(77)));
    layer0_outputs(12662) <= not((inputs(237)) or (inputs(14)));
    layer0_outputs(12663) <= (inputs(68)) xor (inputs(93));
    layer0_outputs(12664) <= (inputs(172)) and not (inputs(145));
    layer0_outputs(12665) <= inputs(114);
    layer0_outputs(12666) <= not((inputs(204)) or (inputs(111)));
    layer0_outputs(12667) <= not((inputs(199)) xor (inputs(88)));
    layer0_outputs(12668) <= not(inputs(166)) or (inputs(37));
    layer0_outputs(12669) <= (inputs(27)) or (inputs(4));
    layer0_outputs(12670) <= not((inputs(93)) xor (inputs(140)));
    layer0_outputs(12671) <= (inputs(51)) and not (inputs(174));
    layer0_outputs(12672) <= not(inputs(60)) or (inputs(241));
    layer0_outputs(12673) <= (inputs(254)) xor (inputs(155));
    layer0_outputs(12674) <= not((inputs(163)) or (inputs(130)));
    layer0_outputs(12675) <= inputs(157);
    layer0_outputs(12676) <= not((inputs(79)) or (inputs(229)));
    layer0_outputs(12677) <= not((inputs(105)) and (inputs(198)));
    layer0_outputs(12678) <= inputs(115);
    layer0_outputs(12679) <= not((inputs(57)) or (inputs(63)));
    layer0_outputs(12680) <= not(inputs(194));
    layer0_outputs(12681) <= (inputs(3)) xor (inputs(239));
    layer0_outputs(12682) <= (inputs(154)) and not (inputs(5));
    layer0_outputs(12683) <= (inputs(215)) and not (inputs(145));
    layer0_outputs(12684) <= inputs(120);
    layer0_outputs(12685) <= not((inputs(106)) xor (inputs(16)));
    layer0_outputs(12686) <= not(inputs(53));
    layer0_outputs(12687) <= not(inputs(247));
    layer0_outputs(12688) <= (inputs(103)) or (inputs(121));
    layer0_outputs(12689) <= inputs(88);
    layer0_outputs(12690) <= not((inputs(218)) xor (inputs(160)));
    layer0_outputs(12691) <= inputs(22);
    layer0_outputs(12692) <= not(inputs(80));
    layer0_outputs(12693) <= (inputs(139)) and not (inputs(79));
    layer0_outputs(12694) <= not(inputs(218));
    layer0_outputs(12695) <= inputs(92);
    layer0_outputs(12696) <= (inputs(156)) or (inputs(69));
    layer0_outputs(12697) <= (inputs(130)) and not (inputs(192));
    layer0_outputs(12698) <= not(inputs(82));
    layer0_outputs(12699) <= (inputs(201)) xor (inputs(83));
    layer0_outputs(12700) <= (inputs(22)) xor (inputs(141));
    layer0_outputs(12701) <= inputs(152);
    layer0_outputs(12702) <= not((inputs(34)) and (inputs(151)));
    layer0_outputs(12703) <= not((inputs(47)) or (inputs(229)));
    layer0_outputs(12704) <= not(inputs(83)) or (inputs(206));
    layer0_outputs(12705) <= not(inputs(99));
    layer0_outputs(12706) <= (inputs(43)) and not (inputs(182));
    layer0_outputs(12707) <= not(inputs(182));
    layer0_outputs(12708) <= not(inputs(25)) or (inputs(117));
    layer0_outputs(12709) <= not((inputs(205)) or (inputs(100)));
    layer0_outputs(12710) <= (inputs(78)) or (inputs(1));
    layer0_outputs(12711) <= not((inputs(24)) or (inputs(192)));
    layer0_outputs(12712) <= not((inputs(85)) or (inputs(207)));
    layer0_outputs(12713) <= not(inputs(59)) or (inputs(64));
    layer0_outputs(12714) <= not(inputs(110));
    layer0_outputs(12715) <= '0';
    layer0_outputs(12716) <= (inputs(192)) or (inputs(98));
    layer0_outputs(12717) <= '1';
    layer0_outputs(12718) <= not(inputs(121)) or (inputs(143));
    layer0_outputs(12719) <= (inputs(83)) and not (inputs(55));
    layer0_outputs(12720) <= (inputs(19)) xor (inputs(49));
    layer0_outputs(12721) <= (inputs(23)) and not (inputs(200));
    layer0_outputs(12722) <= (inputs(251)) or (inputs(38));
    layer0_outputs(12723) <= not((inputs(71)) xor (inputs(138)));
    layer0_outputs(12724) <= inputs(193);
    layer0_outputs(12725) <= inputs(7);
    layer0_outputs(12726) <= (inputs(212)) and not (inputs(103));
    layer0_outputs(12727) <= (inputs(108)) and not (inputs(179));
    layer0_outputs(12728) <= (inputs(39)) or (inputs(49));
    layer0_outputs(12729) <= not(inputs(216));
    layer0_outputs(12730) <= not(inputs(186)) or (inputs(243));
    layer0_outputs(12731) <= (inputs(122)) and not (inputs(93));
    layer0_outputs(12732) <= not(inputs(207));
    layer0_outputs(12733) <= (inputs(191)) or (inputs(65));
    layer0_outputs(12734) <= inputs(52);
    layer0_outputs(12735) <= inputs(194);
    layer0_outputs(12736) <= (inputs(54)) and not (inputs(239));
    layer0_outputs(12737) <= (inputs(203)) and not (inputs(93));
    layer0_outputs(12738) <= not(inputs(157)) or (inputs(167));
    layer0_outputs(12739) <= not(inputs(134));
    layer0_outputs(12740) <= (inputs(203)) or (inputs(37));
    layer0_outputs(12741) <= not((inputs(174)) xor (inputs(117)));
    layer0_outputs(12742) <= inputs(26);
    layer0_outputs(12743) <= (inputs(244)) and not (inputs(68));
    layer0_outputs(12744) <= not(inputs(216));
    layer0_outputs(12745) <= not(inputs(192)) or (inputs(117));
    layer0_outputs(12746) <= (inputs(243)) or (inputs(74));
    layer0_outputs(12747) <= not((inputs(85)) and (inputs(69)));
    layer0_outputs(12748) <= not(inputs(250));
    layer0_outputs(12749) <= not((inputs(137)) and (inputs(71)));
    layer0_outputs(12750) <= not((inputs(78)) xor (inputs(109)));
    layer0_outputs(12751) <= inputs(15);
    layer0_outputs(12752) <= (inputs(86)) xor (inputs(55));
    layer0_outputs(12753) <= '1';
    layer0_outputs(12754) <= inputs(165);
    layer0_outputs(12755) <= (inputs(253)) or (inputs(124));
    layer0_outputs(12756) <= (inputs(218)) and not (inputs(43));
    layer0_outputs(12757) <= (inputs(219)) or (inputs(193));
    layer0_outputs(12758) <= not(inputs(168)) or (inputs(93));
    layer0_outputs(12759) <= not(inputs(205)) or (inputs(170));
    layer0_outputs(12760) <= inputs(164);
    layer0_outputs(12761) <= (inputs(253)) or (inputs(94));
    layer0_outputs(12762) <= not(inputs(24)) or (inputs(158));
    layer0_outputs(12763) <= (inputs(116)) or (inputs(109));
    layer0_outputs(12764) <= (inputs(213)) xor (inputs(194));
    layer0_outputs(12765) <= not((inputs(26)) xor (inputs(127)));
    layer0_outputs(12766) <= (inputs(79)) or (inputs(28));
    layer0_outputs(12767) <= not((inputs(54)) or (inputs(162)));
    layer0_outputs(12768) <= (inputs(245)) or (inputs(175));
    layer0_outputs(12769) <= (inputs(138)) and not (inputs(237));
    layer0_outputs(12770) <= not(inputs(76));
    layer0_outputs(12771) <= (inputs(123)) and not (inputs(189));
    layer0_outputs(12772) <= inputs(247);
    layer0_outputs(12773) <= inputs(181);
    layer0_outputs(12774) <= not(inputs(78)) or (inputs(110));
    layer0_outputs(12775) <= not(inputs(167));
    layer0_outputs(12776) <= not(inputs(151)) or (inputs(111));
    layer0_outputs(12777) <= inputs(231);
    layer0_outputs(12778) <= not(inputs(43));
    layer0_outputs(12779) <= inputs(122);
    layer0_outputs(12780) <= not((inputs(240)) or (inputs(135)));
    layer0_outputs(12781) <= inputs(121);
    layer0_outputs(12782) <= not((inputs(73)) or (inputs(39)));
    layer0_outputs(12783) <= (inputs(172)) and (inputs(111));
    layer0_outputs(12784) <= inputs(245);
    layer0_outputs(12785) <= (inputs(52)) or (inputs(154));
    layer0_outputs(12786) <= not(inputs(122));
    layer0_outputs(12787) <= (inputs(135)) and not (inputs(34));
    layer0_outputs(12788) <= not(inputs(246)) or (inputs(64));
    layer0_outputs(12789) <= not(inputs(37));
    layer0_outputs(12790) <= not(inputs(32));
    layer0_outputs(12791) <= (inputs(83)) and not (inputs(169));
    layer0_outputs(12792) <= (inputs(50)) and not (inputs(188));
    layer0_outputs(12793) <= not(inputs(19));
    layer0_outputs(12794) <= inputs(246);
    layer0_outputs(12795) <= not(inputs(253)) or (inputs(32));
    layer0_outputs(12796) <= (inputs(81)) xor (inputs(212));
    layer0_outputs(12797) <= inputs(102);
    layer0_outputs(12798) <= not(inputs(197));
    layer0_outputs(12799) <= not(inputs(40));
    outputs(0) <= layer0_outputs(5968);
    outputs(1) <= layer0_outputs(5956);
    outputs(2) <= layer0_outputs(8592);
    outputs(3) <= (layer0_outputs(4452)) xor (layer0_outputs(136));
    outputs(4) <= layer0_outputs(4686);
    outputs(5) <= (layer0_outputs(10561)) xor (layer0_outputs(29));
    outputs(6) <= layer0_outputs(6234);
    outputs(7) <= (layer0_outputs(4472)) and not (layer0_outputs(4857));
    outputs(8) <= (layer0_outputs(7624)) xor (layer0_outputs(3888));
    outputs(9) <= not((layer0_outputs(9076)) xor (layer0_outputs(11065)));
    outputs(10) <= not(layer0_outputs(2038));
    outputs(11) <= not((layer0_outputs(5465)) xor (layer0_outputs(168)));
    outputs(12) <= (layer0_outputs(12695)) or (layer0_outputs(10575));
    outputs(13) <= layer0_outputs(1070);
    outputs(14) <= (layer0_outputs(11157)) xor (layer0_outputs(9637));
    outputs(15) <= layer0_outputs(12723);
    outputs(16) <= layer0_outputs(3969);
    outputs(17) <= not(layer0_outputs(11873));
    outputs(18) <= layer0_outputs(8647);
    outputs(19) <= layer0_outputs(7152);
    outputs(20) <= not(layer0_outputs(374)) or (layer0_outputs(7531));
    outputs(21) <= not(layer0_outputs(5982));
    outputs(22) <= not(layer0_outputs(3274));
    outputs(23) <= not((layer0_outputs(1739)) and (layer0_outputs(7455)));
    outputs(24) <= not(layer0_outputs(11099));
    outputs(25) <= not((layer0_outputs(2381)) xor (layer0_outputs(3196)));
    outputs(26) <= not(layer0_outputs(6396)) or (layer0_outputs(7487));
    outputs(27) <= not(layer0_outputs(2142));
    outputs(28) <= layer0_outputs(6511);
    outputs(29) <= not(layer0_outputs(8303));
    outputs(30) <= layer0_outputs(11047);
    outputs(31) <= layer0_outputs(2366);
    outputs(32) <= not((layer0_outputs(6361)) xor (layer0_outputs(4693)));
    outputs(33) <= layer0_outputs(4555);
    outputs(34) <= not((layer0_outputs(7314)) and (layer0_outputs(2523)));
    outputs(35) <= not((layer0_outputs(12545)) and (layer0_outputs(9079)));
    outputs(36) <= not(layer0_outputs(7779)) or (layer0_outputs(9158));
    outputs(37) <= layer0_outputs(8847);
    outputs(38) <= layer0_outputs(11089);
    outputs(39) <= not((layer0_outputs(12466)) and (layer0_outputs(4079)));
    outputs(40) <= not(layer0_outputs(3106));
    outputs(41) <= not(layer0_outputs(6336));
    outputs(42) <= layer0_outputs(5409);
    outputs(43) <= not((layer0_outputs(5591)) and (layer0_outputs(9654)));
    outputs(44) <= layer0_outputs(1002);
    outputs(45) <= not(layer0_outputs(2799));
    outputs(46) <= not(layer0_outputs(4618)) or (layer0_outputs(10147));
    outputs(47) <= not((layer0_outputs(3000)) xor (layer0_outputs(6517)));
    outputs(48) <= layer0_outputs(153);
    outputs(49) <= not((layer0_outputs(8145)) xor (layer0_outputs(1431)));
    outputs(50) <= layer0_outputs(5601);
    outputs(51) <= (layer0_outputs(12589)) xor (layer0_outputs(12402));
    outputs(52) <= layer0_outputs(4285);
    outputs(53) <= not((layer0_outputs(5961)) or (layer0_outputs(6597)));
    outputs(54) <= not((layer0_outputs(2190)) and (layer0_outputs(394)));
    outputs(55) <= (layer0_outputs(1355)) xor (layer0_outputs(805));
    outputs(56) <= layer0_outputs(1934);
    outputs(57) <= not(layer0_outputs(2309));
    outputs(58) <= not(layer0_outputs(9424));
    outputs(59) <= not(layer0_outputs(7719));
    outputs(60) <= not(layer0_outputs(2607));
    outputs(61) <= (layer0_outputs(9082)) xor (layer0_outputs(4209));
    outputs(62) <= layer0_outputs(5341);
    outputs(63) <= (layer0_outputs(12390)) or (layer0_outputs(5836));
    outputs(64) <= not(layer0_outputs(5578));
    outputs(65) <= layer0_outputs(4908);
    outputs(66) <= layer0_outputs(12251);
    outputs(67) <= (layer0_outputs(2378)) and not (layer0_outputs(9976));
    outputs(68) <= not(layer0_outputs(6437));
    outputs(69) <= not(layer0_outputs(9505)) or (layer0_outputs(9373));
    outputs(70) <= layer0_outputs(12685);
    outputs(71) <= layer0_outputs(3573);
    outputs(72) <= not(layer0_outputs(4156));
    outputs(73) <= (layer0_outputs(317)) and not (layer0_outputs(6030));
    outputs(74) <= (layer0_outputs(2520)) xor (layer0_outputs(8855));
    outputs(75) <= layer0_outputs(7514);
    outputs(76) <= (layer0_outputs(7426)) xor (layer0_outputs(10810));
    outputs(77) <= (layer0_outputs(12643)) and (layer0_outputs(10851));
    outputs(78) <= (layer0_outputs(5358)) and not (layer0_outputs(5121));
    outputs(79) <= layer0_outputs(3218);
    outputs(80) <= not(layer0_outputs(11973));
    outputs(81) <= '1';
    outputs(82) <= not((layer0_outputs(2444)) xor (layer0_outputs(12008)));
    outputs(83) <= not(layer0_outputs(1158));
    outputs(84) <= not((layer0_outputs(12241)) xor (layer0_outputs(6549)));
    outputs(85) <= not(layer0_outputs(12432));
    outputs(86) <= not((layer0_outputs(3491)) xor (layer0_outputs(11701)));
    outputs(87) <= not((layer0_outputs(4146)) xor (layer0_outputs(2301)));
    outputs(88) <= not((layer0_outputs(4605)) and (layer0_outputs(4190)));
    outputs(89) <= not(layer0_outputs(7186));
    outputs(90) <= (layer0_outputs(702)) xor (layer0_outputs(1114));
    outputs(91) <= layer0_outputs(11538);
    outputs(92) <= (layer0_outputs(5116)) and (layer0_outputs(2124));
    outputs(93) <= (layer0_outputs(8426)) xor (layer0_outputs(3278));
    outputs(94) <= layer0_outputs(3183);
    outputs(95) <= (layer0_outputs(3352)) and not (layer0_outputs(2832));
    outputs(96) <= (layer0_outputs(5668)) and (layer0_outputs(10904));
    outputs(97) <= not(layer0_outputs(1891)) or (layer0_outputs(3959));
    outputs(98) <= not(layer0_outputs(2993)) or (layer0_outputs(11923));
    outputs(99) <= not(layer0_outputs(12191));
    outputs(100) <= layer0_outputs(12389);
    outputs(101) <= not((layer0_outputs(10902)) or (layer0_outputs(11649)));
    outputs(102) <= (layer0_outputs(10487)) xor (layer0_outputs(216));
    outputs(103) <= not(layer0_outputs(8862));
    outputs(104) <= not((layer0_outputs(773)) xor (layer0_outputs(9855)));
    outputs(105) <= not(layer0_outputs(4043)) or (layer0_outputs(7677));
    outputs(106) <= not((layer0_outputs(6184)) and (layer0_outputs(1330)));
    outputs(107) <= not((layer0_outputs(11774)) and (layer0_outputs(3712)));
    outputs(108) <= layer0_outputs(1345);
    outputs(109) <= (layer0_outputs(5744)) xor (layer0_outputs(1249));
    outputs(110) <= not(layer0_outputs(9554)) or (layer0_outputs(4908));
    outputs(111) <= (layer0_outputs(6268)) or (layer0_outputs(5507));
    outputs(112) <= not(layer0_outputs(9429));
    outputs(113) <= not((layer0_outputs(12484)) xor (layer0_outputs(7002)));
    outputs(114) <= (layer0_outputs(12309)) xor (layer0_outputs(11021));
    outputs(115) <= not((layer0_outputs(12399)) xor (layer0_outputs(10564)));
    outputs(116) <= not(layer0_outputs(9441));
    outputs(117) <= not(layer0_outputs(5867));
    outputs(118) <= not(layer0_outputs(4567));
    outputs(119) <= layer0_outputs(7094);
    outputs(120) <= layer0_outputs(3712);
    outputs(121) <= (layer0_outputs(2865)) xor (layer0_outputs(1946));
    outputs(122) <= not(layer0_outputs(6588));
    outputs(123) <= (layer0_outputs(5881)) xor (layer0_outputs(10970));
    outputs(124) <= layer0_outputs(8262);
    outputs(125) <= not(layer0_outputs(11880)) or (layer0_outputs(1802));
    outputs(126) <= not(layer0_outputs(11724)) or (layer0_outputs(2890));
    outputs(127) <= not((layer0_outputs(12527)) xor (layer0_outputs(9091)));
    outputs(128) <= not(layer0_outputs(3190));
    outputs(129) <= (layer0_outputs(11485)) and not (layer0_outputs(7118));
    outputs(130) <= not(layer0_outputs(5012));
    outputs(131) <= layer0_outputs(3987);
    outputs(132) <= layer0_outputs(3771);
    outputs(133) <= (layer0_outputs(867)) xor (layer0_outputs(8754));
    outputs(134) <= layer0_outputs(11278);
    outputs(135) <= (layer0_outputs(1867)) and not (layer0_outputs(10237));
    outputs(136) <= not(layer0_outputs(1139));
    outputs(137) <= layer0_outputs(9787);
    outputs(138) <= layer0_outputs(2574);
    outputs(139) <= (layer0_outputs(1690)) xor (layer0_outputs(3216));
    outputs(140) <= not(layer0_outputs(4790));
    outputs(141) <= not((layer0_outputs(8045)) xor (layer0_outputs(6921)));
    outputs(142) <= not(layer0_outputs(937));
    outputs(143) <= (layer0_outputs(112)) and (layer0_outputs(12644));
    outputs(144) <= not(layer0_outputs(6061));
    outputs(145) <= layer0_outputs(768);
    outputs(146) <= not(layer0_outputs(11251)) or (layer0_outputs(10767));
    outputs(147) <= layer0_outputs(10044);
    outputs(148) <= layer0_outputs(3642);
    outputs(149) <= (layer0_outputs(1691)) and not (layer0_outputs(9877));
    outputs(150) <= not((layer0_outputs(10057)) xor (layer0_outputs(598)));
    outputs(151) <= (layer0_outputs(10678)) xor (layer0_outputs(7571));
    outputs(152) <= layer0_outputs(1226);
    outputs(153) <= not(layer0_outputs(4267));
    outputs(154) <= not(layer0_outputs(6676));
    outputs(155) <= not(layer0_outputs(7503));
    outputs(156) <= not((layer0_outputs(852)) xor (layer0_outputs(9814)));
    outputs(157) <= not((layer0_outputs(8352)) xor (layer0_outputs(10324)));
    outputs(158) <= (layer0_outputs(12696)) xor (layer0_outputs(7221));
    outputs(159) <= layer0_outputs(9340);
    outputs(160) <= not(layer0_outputs(12374)) or (layer0_outputs(7732));
    outputs(161) <= layer0_outputs(1792);
    outputs(162) <= (layer0_outputs(9895)) and not (layer0_outputs(4784));
    outputs(163) <= not(layer0_outputs(9017));
    outputs(164) <= not((layer0_outputs(6453)) and (layer0_outputs(11927)));
    outputs(165) <= not((layer0_outputs(3822)) xor (layer0_outputs(4292)));
    outputs(166) <= (layer0_outputs(1646)) xor (layer0_outputs(4645));
    outputs(167) <= not(layer0_outputs(6692));
    outputs(168) <= not(layer0_outputs(12469));
    outputs(169) <= layer0_outputs(4368);
    outputs(170) <= not((layer0_outputs(5557)) xor (layer0_outputs(4138)));
    outputs(171) <= layer0_outputs(64);
    outputs(172) <= (layer0_outputs(6791)) xor (layer0_outputs(7281));
    outputs(173) <= (layer0_outputs(11228)) or (layer0_outputs(9045));
    outputs(174) <= not(layer0_outputs(11239)) or (layer0_outputs(10733));
    outputs(175) <= (layer0_outputs(10804)) and not (layer0_outputs(8141));
    outputs(176) <= not((layer0_outputs(110)) xor (layer0_outputs(7868)));
    outputs(177) <= layer0_outputs(8268);
    outputs(178) <= not(layer0_outputs(9155)) or (layer0_outputs(7034));
    outputs(179) <= (layer0_outputs(11529)) xor (layer0_outputs(11406));
    outputs(180) <= not(layer0_outputs(12727)) or (layer0_outputs(3028));
    outputs(181) <= layer0_outputs(48);
    outputs(182) <= not(layer0_outputs(9726)) or (layer0_outputs(12588));
    outputs(183) <= not(layer0_outputs(10190));
    outputs(184) <= not(layer0_outputs(1777));
    outputs(185) <= layer0_outputs(6616);
    outputs(186) <= (layer0_outputs(11678)) or (layer0_outputs(10717));
    outputs(187) <= layer0_outputs(414);
    outputs(188) <= (layer0_outputs(6702)) xor (layer0_outputs(8515));
    outputs(189) <= layer0_outputs(8390);
    outputs(190) <= layer0_outputs(4870);
    outputs(191) <= (layer0_outputs(2149)) and not (layer0_outputs(3586));
    outputs(192) <= layer0_outputs(2513);
    outputs(193) <= not((layer0_outputs(6285)) and (layer0_outputs(1551)));
    outputs(194) <= not(layer0_outputs(4109));
    outputs(195) <= layer0_outputs(424);
    outputs(196) <= layer0_outputs(8508);
    outputs(197) <= layer0_outputs(9672);
    outputs(198) <= not(layer0_outputs(8140));
    outputs(199) <= not((layer0_outputs(4502)) xor (layer0_outputs(5373)));
    outputs(200) <= not(layer0_outputs(8942)) or (layer0_outputs(5802));
    outputs(201) <= not((layer0_outputs(3421)) and (layer0_outputs(4440)));
    outputs(202) <= not(layer0_outputs(9623));
    outputs(203) <= not((layer0_outputs(2563)) xor (layer0_outputs(12416)));
    outputs(204) <= not((layer0_outputs(12670)) and (layer0_outputs(11629)));
    outputs(205) <= not(layer0_outputs(10418));
    outputs(206) <= layer0_outputs(6387);
    outputs(207) <= layer0_outputs(3634);
    outputs(208) <= not(layer0_outputs(784)) or (layer0_outputs(11515));
    outputs(209) <= layer0_outputs(3954);
    outputs(210) <= (layer0_outputs(756)) and not (layer0_outputs(2753));
    outputs(211) <= layer0_outputs(4833);
    outputs(212) <= not(layer0_outputs(10485));
    outputs(213) <= (layer0_outputs(562)) xor (layer0_outputs(7393));
    outputs(214) <= layer0_outputs(5019);
    outputs(215) <= not(layer0_outputs(11968));
    outputs(216) <= not(layer0_outputs(8807));
    outputs(217) <= (layer0_outputs(6739)) xor (layer0_outputs(78));
    outputs(218) <= (layer0_outputs(2319)) and not (layer0_outputs(12720));
    outputs(219) <= (layer0_outputs(1637)) xor (layer0_outputs(12326));
    outputs(220) <= not(layer0_outputs(11548));
    outputs(221) <= not((layer0_outputs(3590)) xor (layer0_outputs(405)));
    outputs(222) <= not(layer0_outputs(1144));
    outputs(223) <= not(layer0_outputs(11388));
    outputs(224) <= not(layer0_outputs(1317)) or (layer0_outputs(10174));
    outputs(225) <= not(layer0_outputs(4741));
    outputs(226) <= layer0_outputs(11314);
    outputs(227) <= layer0_outputs(6559);
    outputs(228) <= not(layer0_outputs(8192)) or (layer0_outputs(6550));
    outputs(229) <= (layer0_outputs(9854)) and not (layer0_outputs(10462));
    outputs(230) <= not(layer0_outputs(6098));
    outputs(231) <= not(layer0_outputs(7534));
    outputs(232) <= layer0_outputs(2187);
    outputs(233) <= not((layer0_outputs(7410)) xor (layer0_outputs(3240)));
    outputs(234) <= layer0_outputs(6293);
    outputs(235) <= not(layer0_outputs(9773)) or (layer0_outputs(3875));
    outputs(236) <= not(layer0_outputs(28));
    outputs(237) <= not(layer0_outputs(1438));
    outputs(238) <= layer0_outputs(12605);
    outputs(239) <= layer0_outputs(5362);
    outputs(240) <= not((layer0_outputs(2817)) and (layer0_outputs(1268)));
    outputs(241) <= (layer0_outputs(5443)) xor (layer0_outputs(6581));
    outputs(242) <= (layer0_outputs(12552)) and not (layer0_outputs(8878));
    outputs(243) <= not((layer0_outputs(9025)) xor (layer0_outputs(11433)));
    outputs(244) <= not((layer0_outputs(6224)) xor (layer0_outputs(11669)));
    outputs(245) <= not(layer0_outputs(10));
    outputs(246) <= not(layer0_outputs(9558));
    outputs(247) <= not((layer0_outputs(6766)) xor (layer0_outputs(8783)));
    outputs(248) <= layer0_outputs(3288);
    outputs(249) <= not(layer0_outputs(2638));
    outputs(250) <= layer0_outputs(2834);
    outputs(251) <= (layer0_outputs(12273)) xor (layer0_outputs(3266));
    outputs(252) <= layer0_outputs(4774);
    outputs(253) <= layer0_outputs(3734);
    outputs(254) <= not((layer0_outputs(9300)) xor (layer0_outputs(11443)));
    outputs(255) <= (layer0_outputs(8070)) xor (layer0_outputs(7490));
    outputs(256) <= layer0_outputs(5672);
    outputs(257) <= (layer0_outputs(3874)) and not (layer0_outputs(7021));
    outputs(258) <= (layer0_outputs(6033)) xor (layer0_outputs(12388));
    outputs(259) <= (layer0_outputs(8725)) xor (layer0_outputs(8394));
    outputs(260) <= (layer0_outputs(10486)) and (layer0_outputs(8512));
    outputs(261) <= not(layer0_outputs(533));
    outputs(262) <= (layer0_outputs(3623)) and not (layer0_outputs(7731));
    outputs(263) <= not(layer0_outputs(4071)) or (layer0_outputs(3480));
    outputs(264) <= layer0_outputs(3884);
    outputs(265) <= not(layer0_outputs(11897));
    outputs(266) <= not(layer0_outputs(11884)) or (layer0_outputs(6071));
    outputs(267) <= layer0_outputs(4630);
    outputs(268) <= not(layer0_outputs(5269));
    outputs(269) <= not((layer0_outputs(6031)) xor (layer0_outputs(9160)));
    outputs(270) <= not(layer0_outputs(8154));
    outputs(271) <= (layer0_outputs(933)) or (layer0_outputs(9939));
    outputs(272) <= not((layer0_outputs(5954)) and (layer0_outputs(2238)));
    outputs(273) <= (layer0_outputs(4404)) xor (layer0_outputs(6529));
    outputs(274) <= not(layer0_outputs(6551));
    outputs(275) <= not(layer0_outputs(10338)) or (layer0_outputs(6727));
    outputs(276) <= not((layer0_outputs(5948)) xor (layer0_outputs(8819)));
    outputs(277) <= layer0_outputs(9716);
    outputs(278) <= not((layer0_outputs(12543)) xor (layer0_outputs(7069)));
    outputs(279) <= layer0_outputs(6560);
    outputs(280) <= not(layer0_outputs(5770));
    outputs(281) <= not(layer0_outputs(4315));
    outputs(282) <= (layer0_outputs(11949)) xor (layer0_outputs(3479));
    outputs(283) <= not(layer0_outputs(9508));
    outputs(284) <= not((layer0_outputs(2054)) xor (layer0_outputs(3500)));
    outputs(285) <= not((layer0_outputs(12476)) or (layer0_outputs(6890)));
    outputs(286) <= not((layer0_outputs(334)) xor (layer0_outputs(7716)));
    outputs(287) <= (layer0_outputs(1309)) and (layer0_outputs(4557));
    outputs(288) <= layer0_outputs(1643);
    outputs(289) <= (layer0_outputs(6496)) and not (layer0_outputs(12244));
    outputs(290) <= layer0_outputs(4294);
    outputs(291) <= (layer0_outputs(11613)) xor (layer0_outputs(5999));
    outputs(292) <= not(layer0_outputs(9882));
    outputs(293) <= (layer0_outputs(10068)) xor (layer0_outputs(4644));
    outputs(294) <= not(layer0_outputs(5711));
    outputs(295) <= (layer0_outputs(6951)) xor (layer0_outputs(10311));
    outputs(296) <= not((layer0_outputs(1381)) xor (layer0_outputs(12606)));
    outputs(297) <= not(layer0_outputs(11094)) or (layer0_outputs(12457));
    outputs(298) <= not((layer0_outputs(11401)) and (layer0_outputs(1650)));
    outputs(299) <= layer0_outputs(7524);
    outputs(300) <= not((layer0_outputs(9572)) and (layer0_outputs(3341)));
    outputs(301) <= not(layer0_outputs(547)) or (layer0_outputs(494));
    outputs(302) <= layer0_outputs(5213);
    outputs(303) <= layer0_outputs(4170);
    outputs(304) <= not(layer0_outputs(3692));
    outputs(305) <= not(layer0_outputs(791));
    outputs(306) <= not(layer0_outputs(3701)) or (layer0_outputs(5710));
    outputs(307) <= (layer0_outputs(9559)) and not (layer0_outputs(3899));
    outputs(308) <= layer0_outputs(8118);
    outputs(309) <= layer0_outputs(1863);
    outputs(310) <= layer0_outputs(9887);
    outputs(311) <= layer0_outputs(5047);
    outputs(312) <= not(layer0_outputs(8335));
    outputs(313) <= not(layer0_outputs(7136));
    outputs(314) <= not(layer0_outputs(5788));
    outputs(315) <= not(layer0_outputs(6991));
    outputs(316) <= layer0_outputs(810);
    outputs(317) <= not(layer0_outputs(5176)) or (layer0_outputs(3153));
    outputs(318) <= (layer0_outputs(12286)) xor (layer0_outputs(8294));
    outputs(319) <= (layer0_outputs(6018)) xor (layer0_outputs(2521));
    outputs(320) <= layer0_outputs(8951);
    outputs(321) <= layer0_outputs(12662);
    outputs(322) <= layer0_outputs(9801);
    outputs(323) <= (layer0_outputs(12274)) or (layer0_outputs(7216));
    outputs(324) <= layer0_outputs(10643);
    outputs(325) <= not((layer0_outputs(5902)) or (layer0_outputs(9661)));
    outputs(326) <= layer0_outputs(6169);
    outputs(327) <= (layer0_outputs(5353)) xor (layer0_outputs(11080));
    outputs(328) <= not((layer0_outputs(12271)) and (layer0_outputs(9634)));
    outputs(329) <= layer0_outputs(12426);
    outputs(330) <= not((layer0_outputs(206)) xor (layer0_outputs(10197)));
    outputs(331) <= not((layer0_outputs(8643)) xor (layer0_outputs(10279)));
    outputs(332) <= not(layer0_outputs(488));
    outputs(333) <= not(layer0_outputs(9083));
    outputs(334) <= not((layer0_outputs(1599)) xor (layer0_outputs(8481)));
    outputs(335) <= not(layer0_outputs(12360)) or (layer0_outputs(6382));
    outputs(336) <= not(layer0_outputs(6160));
    outputs(337) <= not((layer0_outputs(10489)) xor (layer0_outputs(9148)));
    outputs(338) <= layer0_outputs(6188);
    outputs(339) <= layer0_outputs(4789);
    outputs(340) <= not(layer0_outputs(647));
    outputs(341) <= layer0_outputs(7254);
    outputs(342) <= layer0_outputs(10226);
    outputs(343) <= not(layer0_outputs(8426));
    outputs(344) <= layer0_outputs(8519);
    outputs(345) <= not(layer0_outputs(8156));
    outputs(346) <= (layer0_outputs(1819)) xor (layer0_outputs(9058));
    outputs(347) <= layer0_outputs(6730);
    outputs(348) <= not((layer0_outputs(10677)) xor (layer0_outputs(10941)));
    outputs(349) <= '1';
    outputs(350) <= not(layer0_outputs(5945));
    outputs(351) <= not((layer0_outputs(7640)) xor (layer0_outputs(10301)));
    outputs(352) <= layer0_outputs(3241);
    outputs(353) <= layer0_outputs(880);
    outputs(354) <= not(layer0_outputs(8293));
    outputs(355) <= not(layer0_outputs(10716));
    outputs(356) <= not(layer0_outputs(393));
    outputs(357) <= not((layer0_outputs(1469)) xor (layer0_outputs(8360)));
    outputs(358) <= not(layer0_outputs(2479)) or (layer0_outputs(9715));
    outputs(359) <= not(layer0_outputs(8487));
    outputs(360) <= not(layer0_outputs(12346));
    outputs(361) <= (layer0_outputs(8219)) and not (layer0_outputs(932));
    outputs(362) <= (layer0_outputs(9040)) xor (layer0_outputs(3638));
    outputs(363) <= layer0_outputs(6925);
    outputs(364) <= '1';
    outputs(365) <= not(layer0_outputs(1544));
    outputs(366) <= not(layer0_outputs(1743)) or (layer0_outputs(2224));
    outputs(367) <= layer0_outputs(1117);
    outputs(368) <= not((layer0_outputs(3898)) and (layer0_outputs(1623)));
    outputs(369) <= layer0_outputs(5664);
    outputs(370) <= (layer0_outputs(4940)) xor (layer0_outputs(8520));
    outputs(371) <= (layer0_outputs(1303)) xor (layer0_outputs(10784));
    outputs(372) <= not(layer0_outputs(1285));
    outputs(373) <= layer0_outputs(5061);
    outputs(374) <= layer0_outputs(4411);
    outputs(375) <= not(layer0_outputs(4847));
    outputs(376) <= not(layer0_outputs(6736));
    outputs(377) <= layer0_outputs(1888);
    outputs(378) <= not(layer0_outputs(10067));
    outputs(379) <= layer0_outputs(3118);
    outputs(380) <= not(layer0_outputs(7964));
    outputs(381) <= (layer0_outputs(12019)) xor (layer0_outputs(4000));
    outputs(382) <= not(layer0_outputs(9980)) or (layer0_outputs(2919));
    outputs(383) <= not((layer0_outputs(5912)) xor (layer0_outputs(4843)));
    outputs(384) <= not(layer0_outputs(9230));
    outputs(385) <= not(layer0_outputs(5318));
    outputs(386) <= layer0_outputs(9969);
    outputs(387) <= (layer0_outputs(6092)) xor (layer0_outputs(11007));
    outputs(388) <= not(layer0_outputs(12404));
    outputs(389) <= not(layer0_outputs(4220));
    outputs(390) <= layer0_outputs(9791);
    outputs(391) <= not((layer0_outputs(2793)) xor (layer0_outputs(12137)));
    outputs(392) <= not(layer0_outputs(7935));
    outputs(393) <= (layer0_outputs(11574)) and not (layer0_outputs(10022));
    outputs(394) <= not(layer0_outputs(281));
    outputs(395) <= not(layer0_outputs(8713)) or (layer0_outputs(3377));
    outputs(396) <= not(layer0_outputs(7933));
    outputs(397) <= (layer0_outputs(12053)) xor (layer0_outputs(12167));
    outputs(398) <= (layer0_outputs(9039)) and not (layer0_outputs(7231));
    outputs(399) <= not(layer0_outputs(9036)) or (layer0_outputs(9650));
    outputs(400) <= (layer0_outputs(12639)) and not (layer0_outputs(2683));
    outputs(401) <= not(layer0_outputs(5759));
    outputs(402) <= layer0_outputs(5991);
    outputs(403) <= (layer0_outputs(5415)) and not (layer0_outputs(4783));
    outputs(404) <= layer0_outputs(11663);
    outputs(405) <= not(layer0_outputs(10585));
    outputs(406) <= not((layer0_outputs(1834)) or (layer0_outputs(9255)));
    outputs(407) <= not(layer0_outputs(2720));
    outputs(408) <= layer0_outputs(4173);
    outputs(409) <= (layer0_outputs(11290)) and (layer0_outputs(4660));
    outputs(410) <= (layer0_outputs(4107)) and (layer0_outputs(4833));
    outputs(411) <= not(layer0_outputs(11729)) or (layer0_outputs(11623));
    outputs(412) <= not((layer0_outputs(1607)) xor (layer0_outputs(12248)));
    outputs(413) <= not(layer0_outputs(2632));
    outputs(414) <= (layer0_outputs(9821)) xor (layer0_outputs(376));
    outputs(415) <= layer0_outputs(2578);
    outputs(416) <= (layer0_outputs(11350)) or (layer0_outputs(3972));
    outputs(417) <= layer0_outputs(2437);
    outputs(418) <= (layer0_outputs(5402)) and not (layer0_outputs(4483));
    outputs(419) <= layer0_outputs(1550);
    outputs(420) <= (layer0_outputs(12655)) and not (layer0_outputs(8833));
    outputs(421) <= (layer0_outputs(4902)) and (layer0_outputs(3832));
    outputs(422) <= not(layer0_outputs(3723));
    outputs(423) <= not(layer0_outputs(10202));
    outputs(424) <= not((layer0_outputs(700)) xor (layer0_outputs(5283)));
    outputs(425) <= layer0_outputs(9309);
    outputs(426) <= not(layer0_outputs(7897));
    outputs(427) <= layer0_outputs(1714);
    outputs(428) <= not(layer0_outputs(10840)) or (layer0_outputs(666));
    outputs(429) <= not(layer0_outputs(3765));
    outputs(430) <= (layer0_outputs(12135)) and not (layer0_outputs(992));
    outputs(431) <= layer0_outputs(217);
    outputs(432) <= not(layer0_outputs(4414)) or (layer0_outputs(3243));
    outputs(433) <= not(layer0_outputs(9155));
    outputs(434) <= not(layer0_outputs(186));
    outputs(435) <= not(layer0_outputs(9254));
    outputs(436) <= layer0_outputs(5787);
    outputs(437) <= (layer0_outputs(11943)) or (layer0_outputs(3896));
    outputs(438) <= not(layer0_outputs(1489));
    outputs(439) <= not(layer0_outputs(7359)) or (layer0_outputs(6771));
    outputs(440) <= layer0_outputs(8632);
    outputs(441) <= not(layer0_outputs(4977));
    outputs(442) <= not(layer0_outputs(12355)) or (layer0_outputs(11489));
    outputs(443) <= layer0_outputs(7293);
    outputs(444) <= not((layer0_outputs(7641)) and (layer0_outputs(7423)));
    outputs(445) <= not((layer0_outputs(7814)) xor (layer0_outputs(2042)));
    outputs(446) <= not(layer0_outputs(6518));
    outputs(447) <= layer0_outputs(7901);
    outputs(448) <= layer0_outputs(3202);
    outputs(449) <= not(layer0_outputs(2550));
    outputs(450) <= not(layer0_outputs(7741));
    outputs(451) <= not((layer0_outputs(2493)) and (layer0_outputs(8017)));
    outputs(452) <= (layer0_outputs(8199)) and not (layer0_outputs(8771));
    outputs(453) <= not(layer0_outputs(11581));
    outputs(454) <= not((layer0_outputs(2559)) and (layer0_outputs(6777)));
    outputs(455) <= layer0_outputs(1116);
    outputs(456) <= (layer0_outputs(6502)) and not (layer0_outputs(11461));
    outputs(457) <= layer0_outputs(12416);
    outputs(458) <= not((layer0_outputs(11161)) and (layer0_outputs(4344)));
    outputs(459) <= (layer0_outputs(3105)) xor (layer0_outputs(3701));
    outputs(460) <= not((layer0_outputs(6278)) xor (layer0_outputs(12012)));
    outputs(461) <= layer0_outputs(12325);
    outputs(462) <= not((layer0_outputs(9539)) xor (layer0_outputs(8394)));
    outputs(463) <= (layer0_outputs(4494)) and not (layer0_outputs(8317));
    outputs(464) <= layer0_outputs(6456);
    outputs(465) <= not(layer0_outputs(3274));
    outputs(466) <= (layer0_outputs(8052)) xor (layer0_outputs(714));
    outputs(467) <= not(layer0_outputs(7088));
    outputs(468) <= not((layer0_outputs(2877)) xor (layer0_outputs(8924)));
    outputs(469) <= not(layer0_outputs(7947));
    outputs(470) <= not(layer0_outputs(4953));
    outputs(471) <= not((layer0_outputs(11681)) and (layer0_outputs(5314)));
    outputs(472) <= not((layer0_outputs(6996)) and (layer0_outputs(1228)));
    outputs(473) <= (layer0_outputs(520)) xor (layer0_outputs(2766));
    outputs(474) <= (layer0_outputs(3984)) xor (layer0_outputs(3592));
    outputs(475) <= not(layer0_outputs(608)) or (layer0_outputs(10114));
    outputs(476) <= not(layer0_outputs(10481)) or (layer0_outputs(1515));
    outputs(477) <= not(layer0_outputs(10976));
    outputs(478) <= not(layer0_outputs(1039)) or (layer0_outputs(5649));
    outputs(479) <= (layer0_outputs(10404)) and not (layer0_outputs(427));
    outputs(480) <= layer0_outputs(9007);
    outputs(481) <= not(layer0_outputs(7081));
    outputs(482) <= not((layer0_outputs(2790)) xor (layer0_outputs(6926)));
    outputs(483) <= (layer0_outputs(11352)) and (layer0_outputs(2196));
    outputs(484) <= (layer0_outputs(8360)) xor (layer0_outputs(5643));
    outputs(485) <= not(layer0_outputs(7148));
    outputs(486) <= (layer0_outputs(8081)) xor (layer0_outputs(4066));
    outputs(487) <= not(layer0_outputs(5951));
    outputs(488) <= (layer0_outputs(2928)) and not (layer0_outputs(5441));
    outputs(489) <= not(layer0_outputs(10094)) or (layer0_outputs(10171));
    outputs(490) <= layer0_outputs(4370);
    outputs(491) <= (layer0_outputs(45)) xor (layer0_outputs(7493));
    outputs(492) <= layer0_outputs(6448);
    outputs(493) <= not(layer0_outputs(5650)) or (layer0_outputs(12502));
    outputs(494) <= (layer0_outputs(7238)) xor (layer0_outputs(11227));
    outputs(495) <= (layer0_outputs(3509)) xor (layer0_outputs(9784));
    outputs(496) <= (layer0_outputs(4020)) xor (layer0_outputs(10117));
    outputs(497) <= layer0_outputs(120);
    outputs(498) <= not(layer0_outputs(3565));
    outputs(499) <= not((layer0_outputs(6464)) xor (layer0_outputs(12698)));
    outputs(500) <= layer0_outputs(11082);
    outputs(501) <= layer0_outputs(2738);
    outputs(502) <= not(layer0_outputs(9700));
    outputs(503) <= not(layer0_outputs(1857));
    outputs(504) <= layer0_outputs(9306);
    outputs(505) <= layer0_outputs(11438);
    outputs(506) <= not(layer0_outputs(488));
    outputs(507) <= not((layer0_outputs(1266)) and (layer0_outputs(8107)));
    outputs(508) <= layer0_outputs(6263);
    outputs(509) <= not(layer0_outputs(5363));
    outputs(510) <= not((layer0_outputs(12402)) xor (layer0_outputs(2656)));
    outputs(511) <= layer0_outputs(9013);
    outputs(512) <= (layer0_outputs(1429)) and (layer0_outputs(121));
    outputs(513) <= not(layer0_outputs(6999));
    outputs(514) <= (layer0_outputs(12493)) xor (layer0_outputs(7314));
    outputs(515) <= layer0_outputs(7695);
    outputs(516) <= layer0_outputs(8551);
    outputs(517) <= (layer0_outputs(5048)) xor (layer0_outputs(5673));
    outputs(518) <= not(layer0_outputs(5335));
    outputs(519) <= layer0_outputs(11510);
    outputs(520) <= not(layer0_outputs(8036)) or (layer0_outputs(9124));
    outputs(521) <= not((layer0_outputs(11441)) or (layer0_outputs(4935)));
    outputs(522) <= not(layer0_outputs(7197));
    outputs(523) <= layer0_outputs(735);
    outputs(524) <= not((layer0_outputs(8628)) xor (layer0_outputs(1961)));
    outputs(525) <= (layer0_outputs(12335)) or (layer0_outputs(8046));
    outputs(526) <= not(layer0_outputs(7202)) or (layer0_outputs(9383));
    outputs(527) <= layer0_outputs(3814);
    outputs(528) <= not(layer0_outputs(1));
    outputs(529) <= (layer0_outputs(874)) or (layer0_outputs(11037));
    outputs(530) <= (layer0_outputs(2321)) and not (layer0_outputs(3404));
    outputs(531) <= layer0_outputs(4869);
    outputs(532) <= not((layer0_outputs(8822)) xor (layer0_outputs(1153)));
    outputs(533) <= layer0_outputs(5885);
    outputs(534) <= not((layer0_outputs(2062)) and (layer0_outputs(5089)));
    outputs(535) <= not((layer0_outputs(976)) xor (layer0_outputs(1513)));
    outputs(536) <= layer0_outputs(2955);
    outputs(537) <= not(layer0_outputs(11894));
    outputs(538) <= (layer0_outputs(10914)) xor (layer0_outputs(740));
    outputs(539) <= (layer0_outputs(7003)) and not (layer0_outputs(2697));
    outputs(540) <= layer0_outputs(10440);
    outputs(541) <= (layer0_outputs(5104)) xor (layer0_outputs(9470));
    outputs(542) <= not(layer0_outputs(4491));
    outputs(543) <= layer0_outputs(4982);
    outputs(544) <= layer0_outputs(2912);
    outputs(545) <= not(layer0_outputs(10528));
    outputs(546) <= layer0_outputs(2537);
    outputs(547) <= not(layer0_outputs(5411));
    outputs(548) <= layer0_outputs(5572);
    outputs(549) <= not(layer0_outputs(9700));
    outputs(550) <= layer0_outputs(9969);
    outputs(551) <= layer0_outputs(3576);
    outputs(552) <= not(layer0_outputs(11079));
    outputs(553) <= not(layer0_outputs(4114)) or (layer0_outputs(10098));
    outputs(554) <= (layer0_outputs(5753)) xor (layer0_outputs(7977));
    outputs(555) <= layer0_outputs(10039);
    outputs(556) <= not(layer0_outputs(3970));
    outputs(557) <= layer0_outputs(4848);
    outputs(558) <= not(layer0_outputs(9070));
    outputs(559) <= not((layer0_outputs(6103)) xor (layer0_outputs(6197)));
    outputs(560) <= layer0_outputs(10236);
    outputs(561) <= not(layer0_outputs(6157));
    outputs(562) <= layer0_outputs(5118);
    outputs(563) <= (layer0_outputs(1275)) xor (layer0_outputs(11415));
    outputs(564) <= layer0_outputs(3977);
    outputs(565) <= layer0_outputs(961);
    outputs(566) <= not((layer0_outputs(5907)) and (layer0_outputs(12184)));
    outputs(567) <= not(layer0_outputs(4297));
    outputs(568) <= layer0_outputs(1044);
    outputs(569) <= not((layer0_outputs(6566)) and (layer0_outputs(8176)));
    outputs(570) <= (layer0_outputs(487)) and not (layer0_outputs(5897));
    outputs(571) <= not(layer0_outputs(7548));
    outputs(572) <= not(layer0_outputs(836));
    outputs(573) <= not(layer0_outputs(3468)) or (layer0_outputs(10567));
    outputs(574) <= not((layer0_outputs(5885)) xor (layer0_outputs(8871)));
    outputs(575) <= (layer0_outputs(4912)) and not (layer0_outputs(8787));
    outputs(576) <= layer0_outputs(9285);
    outputs(577) <= layer0_outputs(1271);
    outputs(578) <= not(layer0_outputs(1434));
    outputs(579) <= layer0_outputs(8793);
    outputs(580) <= layer0_outputs(12337);
    outputs(581) <= not(layer0_outputs(11946));
    outputs(582) <= not(layer0_outputs(10328)) or (layer0_outputs(7807));
    outputs(583) <= not((layer0_outputs(7400)) and (layer0_outputs(5185)));
    outputs(584) <= not(layer0_outputs(2137));
    outputs(585) <= not(layer0_outputs(5724)) or (layer0_outputs(632));
    outputs(586) <= not((layer0_outputs(3276)) xor (layer0_outputs(7814)));
    outputs(587) <= not((layer0_outputs(9829)) xor (layer0_outputs(6334)));
    outputs(588) <= not(layer0_outputs(7164)) or (layer0_outputs(1713));
    outputs(589) <= not(layer0_outputs(10164));
    outputs(590) <= not(layer0_outputs(6678));
    outputs(591) <= not(layer0_outputs(4145)) or (layer0_outputs(1810));
    outputs(592) <= not(layer0_outputs(2071));
    outputs(593) <= not(layer0_outputs(12701));
    outputs(594) <= layer0_outputs(837);
    outputs(595) <= layer0_outputs(3670);
    outputs(596) <= layer0_outputs(513);
    outputs(597) <= (layer0_outputs(5487)) or (layer0_outputs(5719));
    outputs(598) <= not(layer0_outputs(10444));
    outputs(599) <= layer0_outputs(1445);
    outputs(600) <= layer0_outputs(7529);
    outputs(601) <= not(layer0_outputs(5609));
    outputs(602) <= (layer0_outputs(97)) and not (layer0_outputs(6755));
    outputs(603) <= not(layer0_outputs(8614)) or (layer0_outputs(224));
    outputs(604) <= not(layer0_outputs(10327));
    outputs(605) <= layer0_outputs(9852);
    outputs(606) <= (layer0_outputs(10183)) xor (layer0_outputs(7381));
    outputs(607) <= not(layer0_outputs(12750));
    outputs(608) <= not(layer0_outputs(8468)) or (layer0_outputs(8835));
    outputs(609) <= (layer0_outputs(3206)) or (layer0_outputs(304));
    outputs(610) <= not(layer0_outputs(4480));
    outputs(611) <= (layer0_outputs(3213)) and not (layer0_outputs(11305));
    outputs(612) <= (layer0_outputs(7180)) and (layer0_outputs(5976));
    outputs(613) <= not(layer0_outputs(19));
    outputs(614) <= not((layer0_outputs(2358)) xor (layer0_outputs(1941)));
    outputs(615) <= layer0_outputs(1204);
    outputs(616) <= layer0_outputs(5239);
    outputs(617) <= not((layer0_outputs(10713)) and (layer0_outputs(12020)));
    outputs(618) <= not((layer0_outputs(4145)) or (layer0_outputs(3932)));
    outputs(619) <= (layer0_outputs(3566)) or (layer0_outputs(6774));
    outputs(620) <= layer0_outputs(4650);
    outputs(621) <= not((layer0_outputs(9022)) xor (layer0_outputs(5971)));
    outputs(622) <= not((layer0_outputs(4725)) xor (layer0_outputs(12635)));
    outputs(623) <= not(layer0_outputs(6461)) or (layer0_outputs(3582));
    outputs(624) <= not((layer0_outputs(7428)) and (layer0_outputs(6667)));
    outputs(625) <= layer0_outputs(6012);
    outputs(626) <= (layer0_outputs(10130)) xor (layer0_outputs(3571));
    outputs(627) <= (layer0_outputs(3849)) and (layer0_outputs(5098));
    outputs(628) <= not(layer0_outputs(8732));
    outputs(629) <= not(layer0_outputs(3857));
    outputs(630) <= layer0_outputs(7198);
    outputs(631) <= not(layer0_outputs(6956));
    outputs(632) <= (layer0_outputs(3836)) and not (layer0_outputs(2780));
    outputs(633) <= (layer0_outputs(2459)) xor (layer0_outputs(4928));
    outputs(634) <= not(layer0_outputs(3359)) or (layer0_outputs(5595));
    outputs(635) <= layer0_outputs(3622);
    outputs(636) <= layer0_outputs(1520);
    outputs(637) <= not(layer0_outputs(9324));
    outputs(638) <= not(layer0_outputs(8577));
    outputs(639) <= not(layer0_outputs(11938));
    outputs(640) <= not(layer0_outputs(11854));
    outputs(641) <= not((layer0_outputs(6624)) xor (layer0_outputs(6949)));
    outputs(642) <= (layer0_outputs(3959)) or (layer0_outputs(10333));
    outputs(643) <= not(layer0_outputs(8302)) or (layer0_outputs(4234));
    outputs(644) <= (layer0_outputs(4536)) and not (layer0_outputs(6571));
    outputs(645) <= not((layer0_outputs(9825)) xor (layer0_outputs(7226)));
    outputs(646) <= (layer0_outputs(10855)) xor (layer0_outputs(879));
    outputs(647) <= not(layer0_outputs(2673));
    outputs(648) <= (layer0_outputs(8476)) or (layer0_outputs(10668));
    outputs(649) <= (layer0_outputs(11698)) or (layer0_outputs(7198));
    outputs(650) <= not((layer0_outputs(2023)) and (layer0_outputs(3811)));
    outputs(651) <= not(layer0_outputs(10724)) or (layer0_outputs(2804));
    outputs(652) <= layer0_outputs(1594);
    outputs(653) <= layer0_outputs(10156);
    outputs(654) <= not(layer0_outputs(11219));
    outputs(655) <= layer0_outputs(3619);
    outputs(656) <= (layer0_outputs(2970)) xor (layer0_outputs(11520));
    outputs(657) <= (layer0_outputs(2174)) or (layer0_outputs(5264));
    outputs(658) <= layer0_outputs(2808);
    outputs(659) <= (layer0_outputs(6460)) and not (layer0_outputs(1774));
    outputs(660) <= layer0_outputs(2056);
    outputs(661) <= (layer0_outputs(8521)) xor (layer0_outputs(3525));
    outputs(662) <= not((layer0_outputs(8053)) xor (layer0_outputs(744)));
    outputs(663) <= layer0_outputs(9185);
    outputs(664) <= not((layer0_outputs(12170)) xor (layer0_outputs(3552)));
    outputs(665) <= (layer0_outputs(1179)) or (layer0_outputs(10355));
    outputs(666) <= not(layer0_outputs(1317));
    outputs(667) <= layer0_outputs(6559);
    outputs(668) <= not(layer0_outputs(3027));
    outputs(669) <= layer0_outputs(5886);
    outputs(670) <= not(layer0_outputs(5830));
    outputs(671) <= layer0_outputs(11380);
    outputs(672) <= not((layer0_outputs(5326)) or (layer0_outputs(5302)));
    outputs(673) <= not((layer0_outputs(7098)) or (layer0_outputs(5069)));
    outputs(674) <= not(layer0_outputs(1737)) or (layer0_outputs(593));
    outputs(675) <= not(layer0_outputs(5038)) or (layer0_outputs(5638));
    outputs(676) <= not(layer0_outputs(4143)) or (layer0_outputs(7217));
    outputs(677) <= (layer0_outputs(5528)) xor (layer0_outputs(7265));
    outputs(678) <= (layer0_outputs(5733)) and not (layer0_outputs(1462));
    outputs(679) <= (layer0_outputs(10526)) xor (layer0_outputs(4129));
    outputs(680) <= not(layer0_outputs(11598)) or (layer0_outputs(5803));
    outputs(681) <= not(layer0_outputs(3164));
    outputs(682) <= not(layer0_outputs(10262));
    outputs(683) <= layer0_outputs(11375);
    outputs(684) <= not((layer0_outputs(7100)) or (layer0_outputs(4606)));
    outputs(685) <= layer0_outputs(5173);
    outputs(686) <= layer0_outputs(5755);
    outputs(687) <= not(layer0_outputs(4021));
    outputs(688) <= not((layer0_outputs(1967)) xor (layer0_outputs(3111)));
    outputs(689) <= not((layer0_outputs(10024)) xor (layer0_outputs(9727)));
    outputs(690) <= layer0_outputs(4349);
    outputs(691) <= layer0_outputs(6550);
    outputs(692) <= not((layer0_outputs(10295)) and (layer0_outputs(10989)));
    outputs(693) <= not(layer0_outputs(7244));
    outputs(694) <= not(layer0_outputs(10589));
    outputs(695) <= (layer0_outputs(3310)) and (layer0_outputs(1702));
    outputs(696) <= not(layer0_outputs(8316));
    outputs(697) <= not(layer0_outputs(9923));
    outputs(698) <= not((layer0_outputs(9864)) xor (layer0_outputs(1335)));
    outputs(699) <= layer0_outputs(2791);
    outputs(700) <= not((layer0_outputs(6714)) xor (layer0_outputs(2401)));
    outputs(701) <= not(layer0_outputs(12220)) or (layer0_outputs(6830));
    outputs(702) <= layer0_outputs(5262);
    outputs(703) <= layer0_outputs(3887);
    outputs(704) <= (layer0_outputs(5715)) and (layer0_outputs(7421));
    outputs(705) <= (layer0_outputs(12283)) and (layer0_outputs(2685));
    outputs(706) <= layer0_outputs(9867);
    outputs(707) <= not(layer0_outputs(2562));
    outputs(708) <= (layer0_outputs(9789)) xor (layer0_outputs(8308));
    outputs(709) <= not(layer0_outputs(4003));
    outputs(710) <= layer0_outputs(12209);
    outputs(711) <= layer0_outputs(7480);
    outputs(712) <= layer0_outputs(12319);
    outputs(713) <= (layer0_outputs(5358)) and not (layer0_outputs(12151));
    outputs(714) <= not((layer0_outputs(10655)) and (layer0_outputs(10005)));
    outputs(715) <= layer0_outputs(7523);
    outputs(716) <= layer0_outputs(12780);
    outputs(717) <= not(layer0_outputs(9703)) or (layer0_outputs(9291));
    outputs(718) <= layer0_outputs(2019);
    outputs(719) <= not(layer0_outputs(3922));
    outputs(720) <= not(layer0_outputs(4492));
    outputs(721) <= not(layer0_outputs(10604));
    outputs(722) <= not((layer0_outputs(6779)) xor (layer0_outputs(4095)));
    outputs(723) <= layer0_outputs(12265);
    outputs(724) <= not(layer0_outputs(5030));
    outputs(725) <= not(layer0_outputs(3329));
    outputs(726) <= not((layer0_outputs(759)) or (layer0_outputs(2355)));
    outputs(727) <= layer0_outputs(7892);
    outputs(728) <= not((layer0_outputs(7991)) xor (layer0_outputs(1363)));
    outputs(729) <= (layer0_outputs(9313)) xor (layer0_outputs(6693));
    outputs(730) <= layer0_outputs(262);
    outputs(731) <= layer0_outputs(103);
    outputs(732) <= not((layer0_outputs(9865)) or (layer0_outputs(11273)));
    outputs(733) <= layer0_outputs(5385);
    outputs(734) <= not(layer0_outputs(2464)) or (layer0_outputs(11980));
    outputs(735) <= (layer0_outputs(2648)) or (layer0_outputs(7086));
    outputs(736) <= layer0_outputs(1877);
    outputs(737) <= layer0_outputs(11414);
    outputs(738) <= (layer0_outputs(2161)) and (layer0_outputs(2549));
    outputs(739) <= (layer0_outputs(210)) xor (layer0_outputs(7708));
    outputs(740) <= not(layer0_outputs(6028)) or (layer0_outputs(9746));
    outputs(741) <= not(layer0_outputs(2205));
    outputs(742) <= not(layer0_outputs(7604));
    outputs(743) <= (layer0_outputs(3595)) or (layer0_outputs(12183));
    outputs(744) <= not((layer0_outputs(12023)) or (layer0_outputs(12074)));
    outputs(745) <= (layer0_outputs(1717)) or (layer0_outputs(7445));
    outputs(746) <= layer0_outputs(5301);
    outputs(747) <= (layer0_outputs(7612)) and not (layer0_outputs(5843));
    outputs(748) <= (layer0_outputs(8998)) and not (layer0_outputs(32));
    outputs(749) <= not(layer0_outputs(8385));
    outputs(750) <= layer0_outputs(3435);
    outputs(751) <= layer0_outputs(9531);
    outputs(752) <= (layer0_outputs(6765)) and (layer0_outputs(1995));
    outputs(753) <= layer0_outputs(683);
    outputs(754) <= layer0_outputs(7303);
    outputs(755) <= not(layer0_outputs(8542));
    outputs(756) <= (layer0_outputs(3837)) and not (layer0_outputs(1059));
    outputs(757) <= not((layer0_outputs(11636)) xor (layer0_outputs(3107)));
    outputs(758) <= (layer0_outputs(3713)) xor (layer0_outputs(9750));
    outputs(759) <= not((layer0_outputs(7459)) xor (layer0_outputs(6843)));
    outputs(760) <= (layer0_outputs(5038)) xor (layer0_outputs(3370));
    outputs(761) <= not(layer0_outputs(3397));
    outputs(762) <= not(layer0_outputs(7764)) or (layer0_outputs(7996));
    outputs(763) <= not(layer0_outputs(10717)) or (layer0_outputs(6170));
    outputs(764) <= not((layer0_outputs(8210)) or (layer0_outputs(5075)));
    outputs(765) <= not(layer0_outputs(10842));
    outputs(766) <= (layer0_outputs(5264)) or (layer0_outputs(3706));
    outputs(767) <= not((layer0_outputs(6148)) xor (layer0_outputs(8035)));
    outputs(768) <= (layer0_outputs(8953)) or (layer0_outputs(1503));
    outputs(769) <= not(layer0_outputs(7952));
    outputs(770) <= (layer0_outputs(4984)) and (layer0_outputs(5715));
    outputs(771) <= not(layer0_outputs(1267));
    outputs(772) <= (layer0_outputs(4596)) or (layer0_outputs(10039));
    outputs(773) <= '1';
    outputs(774) <= layer0_outputs(5734);
    outputs(775) <= layer0_outputs(4788);
    outputs(776) <= not((layer0_outputs(3374)) xor (layer0_outputs(5808)));
    outputs(777) <= (layer0_outputs(5183)) and not (layer0_outputs(9114));
    outputs(778) <= layer0_outputs(1570);
    outputs(779) <= layer0_outputs(10314);
    outputs(780) <= not(layer0_outputs(4538));
    outputs(781) <= not(layer0_outputs(1229));
    outputs(782) <= not(layer0_outputs(5285)) or (layer0_outputs(484));
    outputs(783) <= layer0_outputs(9054);
    outputs(784) <= layer0_outputs(11545);
    outputs(785) <= not((layer0_outputs(4360)) and (layer0_outputs(6967)));
    outputs(786) <= layer0_outputs(4856);
    outputs(787) <= not(layer0_outputs(1763));
    outputs(788) <= not(layer0_outputs(5013));
    outputs(789) <= (layer0_outputs(10930)) xor (layer0_outputs(5908));
    outputs(790) <= (layer0_outputs(12183)) and not (layer0_outputs(7884));
    outputs(791) <= not(layer0_outputs(1609));
    outputs(792) <= not((layer0_outputs(6418)) xor (layer0_outputs(5322)));
    outputs(793) <= not((layer0_outputs(9005)) and (layer0_outputs(7425)));
    outputs(794) <= not(layer0_outputs(7857));
    outputs(795) <= not((layer0_outputs(342)) and (layer0_outputs(1556)));
    outputs(796) <= not(layer0_outputs(8068));
    outputs(797) <= not(layer0_outputs(877)) or (layer0_outputs(930));
    outputs(798) <= layer0_outputs(4232);
    outputs(799) <= not(layer0_outputs(9096));
    outputs(800) <= not(layer0_outputs(6340));
    outputs(801) <= (layer0_outputs(2551)) xor (layer0_outputs(4211));
    outputs(802) <= not((layer0_outputs(8188)) xor (layer0_outputs(11059)));
    outputs(803) <= not(layer0_outputs(5304));
    outputs(804) <= not(layer0_outputs(6497));
    outputs(805) <= layer0_outputs(9011);
    outputs(806) <= not((layer0_outputs(12455)) or (layer0_outputs(3505)));
    outputs(807) <= not(layer0_outputs(9713));
    outputs(808) <= not(layer0_outputs(7460));
    outputs(809) <= not(layer0_outputs(6701)) or (layer0_outputs(7199));
    outputs(810) <= not(layer0_outputs(3350));
    outputs(811) <= (layer0_outputs(3494)) and not (layer0_outputs(11266));
    outputs(812) <= (layer0_outputs(12659)) xor (layer0_outputs(11868));
    outputs(813) <= not(layer0_outputs(1587));
    outputs(814) <= (layer0_outputs(8752)) and (layer0_outputs(8008));
    outputs(815) <= layer0_outputs(7248);
    outputs(816) <= layer0_outputs(5295);
    outputs(817) <= not((layer0_outputs(1743)) xor (layer0_outputs(3961)));
    outputs(818) <= layer0_outputs(3129);
    outputs(819) <= layer0_outputs(7261);
    outputs(820) <= layer0_outputs(9490);
    outputs(821) <= (layer0_outputs(7630)) xor (layer0_outputs(11062));
    outputs(822) <= not((layer0_outputs(9636)) xor (layer0_outputs(10756)));
    outputs(823) <= not(layer0_outputs(3852)) or (layer0_outputs(2342));
    outputs(824) <= layer0_outputs(7816);
    outputs(825) <= layer0_outputs(10836);
    outputs(826) <= not((layer0_outputs(1938)) xor (layer0_outputs(1805)));
    outputs(827) <= layer0_outputs(8231);
    outputs(828) <= not(layer0_outputs(7330)) or (layer0_outputs(747));
    outputs(829) <= (layer0_outputs(10823)) or (layer0_outputs(10551));
    outputs(830) <= layer0_outputs(8573);
    outputs(831) <= layer0_outputs(7746);
    outputs(832) <= not(layer0_outputs(4296)) or (layer0_outputs(6629));
    outputs(833) <= layer0_outputs(8870);
    outputs(834) <= not(layer0_outputs(7528)) or (layer0_outputs(11051));
    outputs(835) <= not(layer0_outputs(3281));
    outputs(836) <= not(layer0_outputs(3164));
    outputs(837) <= (layer0_outputs(4944)) xor (layer0_outputs(12164));
    outputs(838) <= layer0_outputs(1939);
    outputs(839) <= layer0_outputs(4641);
    outputs(840) <= not((layer0_outputs(11090)) xor (layer0_outputs(3099)));
    outputs(841) <= not(layer0_outputs(12284));
    outputs(842) <= not(layer0_outputs(9644));
    outputs(843) <= not((layer0_outputs(2823)) and (layer0_outputs(9839)));
    outputs(844) <= (layer0_outputs(5213)) or (layer0_outputs(8775));
    outputs(845) <= (layer0_outputs(4563)) or (layer0_outputs(1026));
    outputs(846) <= not(layer0_outputs(8000));
    outputs(847) <= not(layer0_outputs(3493));
    outputs(848) <= layer0_outputs(7749);
    outputs(849) <= layer0_outputs(5535);
    outputs(850) <= (layer0_outputs(1795)) xor (layer0_outputs(5251));
    outputs(851) <= layer0_outputs(12758);
    outputs(852) <= not(layer0_outputs(12471)) or (layer0_outputs(8270));
    outputs(853) <= not((layer0_outputs(2852)) xor (layer0_outputs(9217)));
    outputs(854) <= not((layer0_outputs(3829)) and (layer0_outputs(4328)));
    outputs(855) <= not((layer0_outputs(10973)) or (layer0_outputs(12587)));
    outputs(856) <= not(layer0_outputs(6311)) or (layer0_outputs(9100));
    outputs(857) <= not((layer0_outputs(8039)) xor (layer0_outputs(6522)));
    outputs(858) <= not(layer0_outputs(6324));
    outputs(859) <= not(layer0_outputs(1902)) or (layer0_outputs(1752));
    outputs(860) <= not((layer0_outputs(9725)) and (layer0_outputs(10563)));
    outputs(861) <= not((layer0_outputs(8198)) and (layer0_outputs(5846)));
    outputs(862) <= not(layer0_outputs(6928)) or (layer0_outputs(737));
    outputs(863) <= (layer0_outputs(9786)) or (layer0_outputs(974));
    outputs(864) <= layer0_outputs(8074);
    outputs(865) <= (layer0_outputs(1678)) and (layer0_outputs(12202));
    outputs(866) <= (layer0_outputs(8168)) and not (layer0_outputs(4690));
    outputs(867) <= (layer0_outputs(12711)) xor (layer0_outputs(12131));
    outputs(868) <= not(layer0_outputs(12092));
    outputs(869) <= (layer0_outputs(1756)) and not (layer0_outputs(8730));
    outputs(870) <= (layer0_outputs(155)) and not (layer0_outputs(5477));
    outputs(871) <= layer0_outputs(2507);
    outputs(872) <= not(layer0_outputs(2262));
    outputs(873) <= not(layer0_outputs(274));
    outputs(874) <= (layer0_outputs(9182)) xor (layer0_outputs(4065));
    outputs(875) <= not(layer0_outputs(3087));
    outputs(876) <= (layer0_outputs(6934)) xor (layer0_outputs(12744));
    outputs(877) <= layer0_outputs(9024);
    outputs(878) <= not(layer0_outputs(1380)) or (layer0_outputs(2139));
    outputs(879) <= layer0_outputs(8093);
    outputs(880) <= (layer0_outputs(10233)) xor (layer0_outputs(9474));
    outputs(881) <= not((layer0_outputs(10132)) xor (layer0_outputs(4478)));
    outputs(882) <= not(layer0_outputs(7358));
    outputs(883) <= layer0_outputs(944);
    outputs(884) <= (layer0_outputs(7879)) xor (layer0_outputs(9702));
    outputs(885) <= not(layer0_outputs(9246));
    outputs(886) <= layer0_outputs(8408);
    outputs(887) <= not((layer0_outputs(5963)) and (layer0_outputs(5807)));
    outputs(888) <= not((layer0_outputs(4546)) and (layer0_outputs(1183)));
    outputs(889) <= layer0_outputs(446);
    outputs(890) <= (layer0_outputs(7136)) xor (layer0_outputs(4346));
    outputs(891) <= layer0_outputs(10353);
    outputs(892) <= (layer0_outputs(8348)) xor (layer0_outputs(10982));
    outputs(893) <= layer0_outputs(4025);
    outputs(894) <= not(layer0_outputs(1655));
    outputs(895) <= (layer0_outputs(999)) xor (layer0_outputs(3338));
    outputs(896) <= (layer0_outputs(7646)) xor (layer0_outputs(5892));
    outputs(897) <= not(layer0_outputs(11509));
    outputs(898) <= not(layer0_outputs(1015)) or (layer0_outputs(1320));
    outputs(899) <= layer0_outputs(7467);
    outputs(900) <= not(layer0_outputs(1494));
    outputs(901) <= (layer0_outputs(9290)) and (layer0_outputs(800));
    outputs(902) <= not(layer0_outputs(9701)) or (layer0_outputs(8464));
    outputs(903) <= not(layer0_outputs(10262));
    outputs(904) <= (layer0_outputs(9273)) xor (layer0_outputs(8720));
    outputs(905) <= '1';
    outputs(906) <= not((layer0_outputs(6657)) or (layer0_outputs(717)));
    outputs(907) <= not(layer0_outputs(766)) or (layer0_outputs(7072));
    outputs(908) <= not(layer0_outputs(3362));
    outputs(909) <= (layer0_outputs(2281)) or (layer0_outputs(6378));
    outputs(910) <= (layer0_outputs(4653)) xor (layer0_outputs(10908));
    outputs(911) <= not(layer0_outputs(5002)) or (layer0_outputs(8870));
    outputs(912) <= (layer0_outputs(11545)) or (layer0_outputs(4327));
    outputs(913) <= (layer0_outputs(10082)) and not (layer0_outputs(2986));
    outputs(914) <= not(layer0_outputs(9094));
    outputs(915) <= not((layer0_outputs(753)) xor (layer0_outputs(6190)));
    outputs(916) <= not(layer0_outputs(4072));
    outputs(917) <= layer0_outputs(175);
    outputs(918) <= not(layer0_outputs(5206));
    outputs(919) <= not((layer0_outputs(3293)) xor (layer0_outputs(4295)));
    outputs(920) <= not(layer0_outputs(8278));
    outputs(921) <= (layer0_outputs(10066)) and not (layer0_outputs(3152));
    outputs(922) <= not(layer0_outputs(554));
    outputs(923) <= (layer0_outputs(5778)) and not (layer0_outputs(2064));
    outputs(924) <= not((layer0_outputs(6589)) xor (layer0_outputs(4936)));
    outputs(925) <= not(layer0_outputs(1031));
    outputs(926) <= (layer0_outputs(2805)) and not (layer0_outputs(11810));
    outputs(927) <= not(layer0_outputs(5120));
    outputs(928) <= layer0_outputs(5002);
    outputs(929) <= (layer0_outputs(5404)) xor (layer0_outputs(2336));
    outputs(930) <= layer0_outputs(6229);
    outputs(931) <= layer0_outputs(10845);
    outputs(932) <= not(layer0_outputs(4493));
    outputs(933) <= layer0_outputs(3776);
    outputs(934) <= (layer0_outputs(1997)) xor (layer0_outputs(667));
    outputs(935) <= layer0_outputs(10739);
    outputs(936) <= not(layer0_outputs(8716));
    outputs(937) <= not((layer0_outputs(11213)) and (layer0_outputs(5113)));
    outputs(938) <= layer0_outputs(11577);
    outputs(939) <= (layer0_outputs(2807)) xor (layer0_outputs(5376));
    outputs(940) <= layer0_outputs(6730);
    outputs(941) <= layer0_outputs(9364);
    outputs(942) <= not((layer0_outputs(1379)) xor (layer0_outputs(1532)));
    outputs(943) <= layer0_outputs(8955);
    outputs(944) <= not((layer0_outputs(1362)) xor (layer0_outputs(5687)));
    outputs(945) <= (layer0_outputs(11319)) xor (layer0_outputs(2409));
    outputs(946) <= layer0_outputs(1674);
    outputs(947) <= (layer0_outputs(11255)) and (layer0_outputs(11835));
    outputs(948) <= layer0_outputs(6797);
    outputs(949) <= not(layer0_outputs(11645));
    outputs(950) <= layer0_outputs(5386);
    outputs(951) <= layer0_outputs(8255);
    outputs(952) <= not((layer0_outputs(2116)) xor (layer0_outputs(8176)));
    outputs(953) <= not(layer0_outputs(6114));
    outputs(954) <= not(layer0_outputs(12112));
    outputs(955) <= (layer0_outputs(10544)) xor (layer0_outputs(722));
    outputs(956) <= not((layer0_outputs(5073)) xor (layer0_outputs(4254)));
    outputs(957) <= layer0_outputs(11972);
    outputs(958) <= not(layer0_outputs(1494));
    outputs(959) <= layer0_outputs(7781);
    outputs(960) <= layer0_outputs(770);
    outputs(961) <= not(layer0_outputs(8284));
    outputs(962) <= not(layer0_outputs(627)) or (layer0_outputs(7036));
    outputs(963) <= not(layer0_outputs(1551));
    outputs(964) <= not(layer0_outputs(12315)) or (layer0_outputs(10235));
    outputs(965) <= not((layer0_outputs(7082)) xor (layer0_outputs(12294)));
    outputs(966) <= layer0_outputs(405);
    outputs(967) <= (layer0_outputs(646)) and not (layer0_outputs(9774));
    outputs(968) <= not(layer0_outputs(12343));
    outputs(969) <= not(layer0_outputs(3265)) or (layer0_outputs(6011));
    outputs(970) <= not(layer0_outputs(8836)) or (layer0_outputs(6343));
    outputs(971) <= not(layer0_outputs(8736));
    outputs(972) <= (layer0_outputs(2148)) xor (layer0_outputs(1468));
    outputs(973) <= layer0_outputs(7008);
    outputs(974) <= layer0_outputs(11583);
    outputs(975) <= layer0_outputs(971);
    outputs(976) <= not((layer0_outputs(5291)) or (layer0_outputs(10302)));
    outputs(977) <= not(layer0_outputs(11056));
    outputs(978) <= (layer0_outputs(3758)) or (layer0_outputs(10911));
    outputs(979) <= not(layer0_outputs(8922));
    outputs(980) <= not(layer0_outputs(6076));
    outputs(981) <= not(layer0_outputs(11099));
    outputs(982) <= not(layer0_outputs(8473));
    outputs(983) <= (layer0_outputs(3437)) or (layer0_outputs(3279));
    outputs(984) <= not((layer0_outputs(10141)) and (layer0_outputs(234)));
    outputs(985) <= (layer0_outputs(921)) xor (layer0_outputs(2502));
    outputs(986) <= (layer0_outputs(8314)) xor (layer0_outputs(651));
    outputs(987) <= not(layer0_outputs(1131));
    outputs(988) <= layer0_outputs(11045);
    outputs(989) <= (layer0_outputs(5288)) xor (layer0_outputs(4201));
    outputs(990) <= layer0_outputs(8438);
    outputs(991) <= layer0_outputs(5646);
    outputs(992) <= layer0_outputs(12142);
    outputs(993) <= layer0_outputs(12739);
    outputs(994) <= (layer0_outputs(264)) xor (layer0_outputs(3013));
    outputs(995) <= not(layer0_outputs(8935));
    outputs(996) <= (layer0_outputs(7748)) and not (layer0_outputs(10318));
    outputs(997) <= not(layer0_outputs(5311));
    outputs(998) <= not(layer0_outputs(5128)) or (layer0_outputs(6851));
    outputs(999) <= not(layer0_outputs(12049)) or (layer0_outputs(6950));
    outputs(1000) <= not((layer0_outputs(8070)) xor (layer0_outputs(7647)));
    outputs(1001) <= (layer0_outputs(9038)) xor (layer0_outputs(7840));
    outputs(1002) <= not(layer0_outputs(11490));
    outputs(1003) <= (layer0_outputs(2994)) xor (layer0_outputs(6663));
    outputs(1004) <= layer0_outputs(9887);
    outputs(1005) <= (layer0_outputs(5920)) xor (layer0_outputs(11687));
    outputs(1006) <= not((layer0_outputs(11353)) xor (layer0_outputs(4602)));
    outputs(1007) <= (layer0_outputs(4759)) and (layer0_outputs(4416));
    outputs(1008) <= layer0_outputs(788);
    outputs(1009) <= layer0_outputs(8431);
    outputs(1010) <= (layer0_outputs(12710)) and (layer0_outputs(251));
    outputs(1011) <= not((layer0_outputs(9588)) xor (layer0_outputs(2273)));
    outputs(1012) <= not(layer0_outputs(5631)) or (layer0_outputs(6552));
    outputs(1013) <= not(layer0_outputs(5343));
    outputs(1014) <= not((layer0_outputs(9516)) xor (layer0_outputs(9656)));
    outputs(1015) <= not(layer0_outputs(9351));
    outputs(1016) <= not((layer0_outputs(6593)) xor (layer0_outputs(4398)));
    outputs(1017) <= (layer0_outputs(8564)) or (layer0_outputs(3167));
    outputs(1018) <= (layer0_outputs(4344)) xor (layer0_outputs(5323));
    outputs(1019) <= not(layer0_outputs(9469));
    outputs(1020) <= not(layer0_outputs(11092));
    outputs(1021) <= not(layer0_outputs(10150));
    outputs(1022) <= not(layer0_outputs(2006));
    outputs(1023) <= not(layer0_outputs(826));
    outputs(1024) <= not(layer0_outputs(2605)) or (layer0_outputs(100));
    outputs(1025) <= (layer0_outputs(6442)) and (layer0_outputs(5139));
    outputs(1026) <= not(layer0_outputs(1914));
    outputs(1027) <= layer0_outputs(5950);
    outputs(1028) <= (layer0_outputs(1936)) or (layer0_outputs(9806));
    outputs(1029) <= not(layer0_outputs(8113)) or (layer0_outputs(4716));
    outputs(1030) <= (layer0_outputs(5938)) and not (layer0_outputs(11935));
    outputs(1031) <= not(layer0_outputs(9228)) or (layer0_outputs(7264));
    outputs(1032) <= layer0_outputs(6636);
    outputs(1033) <= not(layer0_outputs(3341));
    outputs(1034) <= (layer0_outputs(5033)) and not (layer0_outputs(10671));
    outputs(1035) <= not(layer0_outputs(8250)) or (layer0_outputs(4228));
    outputs(1036) <= not(layer0_outputs(8183));
    outputs(1037) <= not((layer0_outputs(2026)) xor (layer0_outputs(5860)));
    outputs(1038) <= not(layer0_outputs(7937));
    outputs(1039) <= layer0_outputs(891);
    outputs(1040) <= (layer0_outputs(9861)) and not (layer0_outputs(5531));
    outputs(1041) <= layer0_outputs(7575);
    outputs(1042) <= not((layer0_outputs(9554)) and (layer0_outputs(11148)));
    outputs(1043) <= layer0_outputs(3220);
    outputs(1044) <= layer0_outputs(7476);
    outputs(1045) <= not((layer0_outputs(6167)) xor (layer0_outputs(11995)));
    outputs(1046) <= not(layer0_outputs(6090));
    outputs(1047) <= not((layer0_outputs(4025)) xor (layer0_outputs(5104)));
    outputs(1048) <= (layer0_outputs(1410)) or (layer0_outputs(10421));
    outputs(1049) <= not(layer0_outputs(4188));
    outputs(1050) <= layer0_outputs(11888);
    outputs(1051) <= (layer0_outputs(168)) or (layer0_outputs(3624));
    outputs(1052) <= layer0_outputs(1345);
    outputs(1053) <= layer0_outputs(2441);
    outputs(1054) <= layer0_outputs(7572);
    outputs(1055) <= layer0_outputs(3022);
    outputs(1056) <= not((layer0_outputs(3229)) xor (layer0_outputs(5289)));
    outputs(1057) <= not(layer0_outputs(5676));
    outputs(1058) <= not(layer0_outputs(4070));
    outputs(1059) <= layer0_outputs(2928);
    outputs(1060) <= not(layer0_outputs(11155));
    outputs(1061) <= layer0_outputs(1154);
    outputs(1062) <= (layer0_outputs(672)) xor (layer0_outputs(6238));
    outputs(1063) <= layer0_outputs(11707);
    outputs(1064) <= not(layer0_outputs(11607));
    outputs(1065) <= layer0_outputs(5099);
    outputs(1066) <= not(layer0_outputs(4424));
    outputs(1067) <= (layer0_outputs(5404)) xor (layer0_outputs(6696));
    outputs(1068) <= not((layer0_outputs(9002)) or (layer0_outputs(8878)));
    outputs(1069) <= (layer0_outputs(6344)) and not (layer0_outputs(10801));
    outputs(1070) <= layer0_outputs(10210);
    outputs(1071) <= not(layer0_outputs(1948));
    outputs(1072) <= (layer0_outputs(8095)) and not (layer0_outputs(11384));
    outputs(1073) <= not(layer0_outputs(12680)) or (layer0_outputs(7162));
    outputs(1074) <= layer0_outputs(6000);
    outputs(1075) <= not(layer0_outputs(815)) or (layer0_outputs(9275));
    outputs(1076) <= (layer0_outputs(12735)) and not (layer0_outputs(184));
    outputs(1077) <= not((layer0_outputs(10965)) xor (layer0_outputs(12185)));
    outputs(1078) <= not(layer0_outputs(1107)) or (layer0_outputs(9949));
    outputs(1079) <= layer0_outputs(3682);
    outputs(1080) <= not(layer0_outputs(2395)) or (layer0_outputs(5729));
    outputs(1081) <= layer0_outputs(10546);
    outputs(1082) <= not((layer0_outputs(6503)) xor (layer0_outputs(5988)));
    outputs(1083) <= layer0_outputs(10499);
    outputs(1084) <= not((layer0_outputs(2606)) xor (layer0_outputs(5753)));
    outputs(1085) <= not((layer0_outputs(2610)) xor (layer0_outputs(9930)));
    outputs(1086) <= not((layer0_outputs(9401)) and (layer0_outputs(3710)));
    outputs(1087) <= (layer0_outputs(708)) and (layer0_outputs(11615));
    outputs(1088) <= not((layer0_outputs(2972)) xor (layer0_outputs(9830)));
    outputs(1089) <= layer0_outputs(9542);
    outputs(1090) <= not((layer0_outputs(5886)) xor (layer0_outputs(12270)));
    outputs(1091) <= not((layer0_outputs(4129)) xor (layer0_outputs(6452)));
    outputs(1092) <= not(layer0_outputs(8285));
    outputs(1093) <= not(layer0_outputs(4538));
    outputs(1094) <= not(layer0_outputs(9515));
    outputs(1095) <= (layer0_outputs(8806)) and not (layer0_outputs(9956));
    outputs(1096) <= (layer0_outputs(4768)) and (layer0_outputs(3309));
    outputs(1097) <= not(layer0_outputs(5013)) or (layer0_outputs(12776));
    outputs(1098) <= not(layer0_outputs(1098));
    outputs(1099) <= layer0_outputs(10077);
    outputs(1100) <= layer0_outputs(3942);
    outputs(1101) <= layer0_outputs(7085);
    outputs(1102) <= (layer0_outputs(2682)) and not (layer0_outputs(5713));
    outputs(1103) <= not(layer0_outputs(3128)) or (layer0_outputs(8750));
    outputs(1104) <= layer0_outputs(11862);
    outputs(1105) <= not(layer0_outputs(8696));
    outputs(1106) <= not(layer0_outputs(4969));
    outputs(1107) <= (layer0_outputs(9544)) and (layer0_outputs(4407));
    outputs(1108) <= not(layer0_outputs(4089));
    outputs(1109) <= not(layer0_outputs(8018));
    outputs(1110) <= not(layer0_outputs(8950));
    outputs(1111) <= (layer0_outputs(4256)) xor (layer0_outputs(239));
    outputs(1112) <= (layer0_outputs(9271)) and not (layer0_outputs(12343));
    outputs(1113) <= not(layer0_outputs(12624)) or (layer0_outputs(8245));
    outputs(1114) <= layer0_outputs(6599);
    outputs(1115) <= (layer0_outputs(11159)) or (layer0_outputs(12531));
    outputs(1116) <= not(layer0_outputs(4222));
    outputs(1117) <= not(layer0_outputs(12731));
    outputs(1118) <= layer0_outputs(12667);
    outputs(1119) <= (layer0_outputs(630)) xor (layer0_outputs(5632));
    outputs(1120) <= layer0_outputs(1632);
    outputs(1121) <= layer0_outputs(7158);
    outputs(1122) <= not((layer0_outputs(10431)) xor (layer0_outputs(8213)));
    outputs(1123) <= not((layer0_outputs(2511)) and (layer0_outputs(6831)));
    outputs(1124) <= not((layer0_outputs(4767)) xor (layer0_outputs(1441)));
    outputs(1125) <= layer0_outputs(5964);
    outputs(1126) <= not(layer0_outputs(6692));
    outputs(1127) <= not(layer0_outputs(12714));
    outputs(1128) <= (layer0_outputs(793)) xor (layer0_outputs(8124));
    outputs(1129) <= layer0_outputs(4322);
    outputs(1130) <= not(layer0_outputs(5133));
    outputs(1131) <= not(layer0_outputs(10556));
    outputs(1132) <= layer0_outputs(9128);
    outputs(1133) <= not(layer0_outputs(7940));
    outputs(1134) <= not((layer0_outputs(449)) or (layer0_outputs(3356)));
    outputs(1135) <= layer0_outputs(5651);
    outputs(1136) <= layer0_outputs(6535);
    outputs(1137) <= not(layer0_outputs(2310));
    outputs(1138) <= not(layer0_outputs(8859)) or (layer0_outputs(7279));
    outputs(1139) <= not((layer0_outputs(1436)) or (layer0_outputs(10246)));
    outputs(1140) <= not((layer0_outputs(4734)) or (layer0_outputs(10467)));
    outputs(1141) <= layer0_outputs(8225);
    outputs(1142) <= layer0_outputs(7971);
    outputs(1143) <= layer0_outputs(5890);
    outputs(1144) <= layer0_outputs(8359);
    outputs(1145) <= not(layer0_outputs(10190));
    outputs(1146) <= not((layer0_outputs(9780)) xor (layer0_outputs(7521)));
    outputs(1147) <= not(layer0_outputs(9911));
    outputs(1148) <= not((layer0_outputs(5816)) or (layer0_outputs(1672)));
    outputs(1149) <= layer0_outputs(6987);
    outputs(1150) <= not((layer0_outputs(11232)) xor (layer0_outputs(9614)));
    outputs(1151) <= not(layer0_outputs(10611)) or (layer0_outputs(9950));
    outputs(1152) <= not(layer0_outputs(6433));
    outputs(1153) <= not(layer0_outputs(8789));
    outputs(1154) <= layer0_outputs(6313);
    outputs(1155) <= not(layer0_outputs(7972));
    outputs(1156) <= layer0_outputs(8112);
    outputs(1157) <= not((layer0_outputs(12011)) xor (layer0_outputs(2129)));
    outputs(1158) <= (layer0_outputs(8861)) and not (layer0_outputs(7096));
    outputs(1159) <= not((layer0_outputs(10670)) xor (layer0_outputs(11765)));
    outputs(1160) <= not(layer0_outputs(11482));
    outputs(1161) <= not(layer0_outputs(6459)) or (layer0_outputs(9071));
    outputs(1162) <= layer0_outputs(1923);
    outputs(1163) <= not((layer0_outputs(785)) xor (layer0_outputs(10230)));
    outputs(1164) <= not(layer0_outputs(3371));
    outputs(1165) <= not(layer0_outputs(10443));
    outputs(1166) <= (layer0_outputs(6547)) and not (layer0_outputs(8311));
    outputs(1167) <= not(layer0_outputs(12237)) or (layer0_outputs(9692));
    outputs(1168) <= not((layer0_outputs(10473)) xor (layer0_outputs(6573)));
    outputs(1169) <= not(layer0_outputs(10116));
    outputs(1170) <= (layer0_outputs(5501)) xor (layer0_outputs(10577));
    outputs(1171) <= layer0_outputs(3348);
    outputs(1172) <= not(layer0_outputs(5880));
    outputs(1173) <= not((layer0_outputs(10259)) xor (layer0_outputs(3805)));
    outputs(1174) <= (layer0_outputs(278)) or (layer0_outputs(6562));
    outputs(1175) <= not(layer0_outputs(3096));
    outputs(1176) <= not(layer0_outputs(8134));
    outputs(1177) <= layer0_outputs(1420);
    outputs(1178) <= layer0_outputs(7818);
    outputs(1179) <= (layer0_outputs(3681)) or (layer0_outputs(6478));
    outputs(1180) <= layer0_outputs(10944);
    outputs(1181) <= not(layer0_outputs(5092));
    outputs(1182) <= not((layer0_outputs(4618)) and (layer0_outputs(4197)));
    outputs(1183) <= not((layer0_outputs(7304)) or (layer0_outputs(8336)));
    outputs(1184) <= not((layer0_outputs(10115)) xor (layer0_outputs(10189)));
    outputs(1185) <= layer0_outputs(2092);
    outputs(1186) <= not(layer0_outputs(9977)) or (layer0_outputs(8115));
    outputs(1187) <= (layer0_outputs(11493)) xor (layer0_outputs(3720));
    outputs(1188) <= not((layer0_outputs(10261)) and (layer0_outputs(3151)));
    outputs(1189) <= layer0_outputs(105);
    outputs(1190) <= not((layer0_outputs(10451)) xor (layer0_outputs(12773)));
    outputs(1191) <= (layer0_outputs(10252)) and not (layer0_outputs(5579));
    outputs(1192) <= not((layer0_outputs(243)) xor (layer0_outputs(2496)));
    outputs(1193) <= (layer0_outputs(12601)) and (layer0_outputs(7949));
    outputs(1194) <= layer0_outputs(9857);
    outputs(1195) <= not(layer0_outputs(4493));
    outputs(1196) <= not(layer0_outputs(3084));
    outputs(1197) <= not(layer0_outputs(7559));
    outputs(1198) <= layer0_outputs(4983);
    outputs(1199) <= not(layer0_outputs(4184));
    outputs(1200) <= not((layer0_outputs(2989)) and (layer0_outputs(4312)));
    outputs(1201) <= (layer0_outputs(11427)) and (layer0_outputs(4972));
    outputs(1202) <= layer0_outputs(5628);
    outputs(1203) <= not(layer0_outputs(2953));
    outputs(1204) <= not((layer0_outputs(1491)) xor (layer0_outputs(3286)));
    outputs(1205) <= not(layer0_outputs(1058)) or (layer0_outputs(4186));
    outputs(1206) <= not((layer0_outputs(11364)) xor (layer0_outputs(3789)));
    outputs(1207) <= (layer0_outputs(12704)) or (layer0_outputs(8111));
    outputs(1208) <= not(layer0_outputs(9647));
    outputs(1209) <= (layer0_outputs(218)) xor (layer0_outputs(10671));
    outputs(1210) <= not(layer0_outputs(11906));
    outputs(1211) <= (layer0_outputs(5573)) xor (layer0_outputs(1134));
    outputs(1212) <= not((layer0_outputs(4765)) xor (layer0_outputs(12134)));
    outputs(1213) <= layer0_outputs(7969);
    outputs(1214) <= (layer0_outputs(3560)) or (layer0_outputs(1481));
    outputs(1215) <= not(layer0_outputs(8223)) or (layer0_outputs(7438));
    outputs(1216) <= (layer0_outputs(6724)) xor (layer0_outputs(5680));
    outputs(1217) <= layer0_outputs(7409);
    outputs(1218) <= layer0_outputs(4223);
    outputs(1219) <= not((layer0_outputs(10072)) or (layer0_outputs(8680)));
    outputs(1220) <= layer0_outputs(9951);
    outputs(1221) <= not(layer0_outputs(3385));
    outputs(1222) <= not((layer0_outputs(12465)) xor (layer0_outputs(941)));
    outputs(1223) <= (layer0_outputs(6978)) xor (layer0_outputs(3187));
    outputs(1224) <= layer0_outputs(3291);
    outputs(1225) <= layer0_outputs(9211);
    outputs(1226) <= not(layer0_outputs(4866)) or (layer0_outputs(11849));
    outputs(1227) <= not(layer0_outputs(6424));
    outputs(1228) <= (layer0_outputs(359)) xor (layer0_outputs(1897));
    outputs(1229) <= not(layer0_outputs(3293)) or (layer0_outputs(10042));
    outputs(1230) <= not((layer0_outputs(3507)) and (layer0_outputs(6317)));
    outputs(1231) <= not((layer0_outputs(8877)) or (layer0_outputs(7378)));
    outputs(1232) <= layer0_outputs(12143);
    outputs(1233) <= (layer0_outputs(1435)) xor (layer0_outputs(1276));
    outputs(1234) <= (layer0_outputs(4544)) xor (layer0_outputs(6217));
    outputs(1235) <= not(layer0_outputs(9807));
    outputs(1236) <= layer0_outputs(4688);
    outputs(1237) <= layer0_outputs(4997);
    outputs(1238) <= not((layer0_outputs(5364)) xor (layer0_outputs(7043)));
    outputs(1239) <= not(layer0_outputs(4364)) or (layer0_outputs(1693));
    outputs(1240) <= not(layer0_outputs(7362)) or (layer0_outputs(907));
    outputs(1241) <= not((layer0_outputs(9041)) xor (layer0_outputs(12055)));
    outputs(1242) <= not(layer0_outputs(6134));
    outputs(1243) <= layer0_outputs(6268);
    outputs(1244) <= (layer0_outputs(9799)) and not (layer0_outputs(12151));
    outputs(1245) <= not(layer0_outputs(5622));
    outputs(1246) <= layer0_outputs(4637);
    outputs(1247) <= not(layer0_outputs(11368));
    outputs(1248) <= layer0_outputs(7398);
    outputs(1249) <= not(layer0_outputs(8273));
    outputs(1250) <= not((layer0_outputs(6367)) or (layer0_outputs(7702)));
    outputs(1251) <= layer0_outputs(11733);
    outputs(1252) <= layer0_outputs(1570);
    outputs(1253) <= layer0_outputs(4809);
    outputs(1254) <= not(layer0_outputs(1563));
    outputs(1255) <= not(layer0_outputs(2780));
    outputs(1256) <= (layer0_outputs(7355)) or (layer0_outputs(9735));
    outputs(1257) <= (layer0_outputs(12283)) or (layer0_outputs(2437));
    outputs(1258) <= (layer0_outputs(9462)) xor (layer0_outputs(5938));
    outputs(1259) <= layer0_outputs(632);
    outputs(1260) <= not((layer0_outputs(3605)) xor (layer0_outputs(12406)));
    outputs(1261) <= (layer0_outputs(5284)) and not (layer0_outputs(8594));
    outputs(1262) <= layer0_outputs(7161);
    outputs(1263) <= (layer0_outputs(3197)) and not (layer0_outputs(11387));
    outputs(1264) <= layer0_outputs(5448);
    outputs(1265) <= (layer0_outputs(6744)) and (layer0_outputs(6681));
    outputs(1266) <= layer0_outputs(9822);
    outputs(1267) <= (layer0_outputs(9617)) and (layer0_outputs(2388));
    outputs(1268) <= layer0_outputs(12216);
    outputs(1269) <= (layer0_outputs(5407)) or (layer0_outputs(10649));
    outputs(1270) <= (layer0_outputs(4389)) xor (layer0_outputs(2992));
    outputs(1271) <= '0';
    outputs(1272) <= layer0_outputs(8639);
    outputs(1273) <= not(layer0_outputs(5103));
    outputs(1274) <= (layer0_outputs(11702)) and (layer0_outputs(8419));
    outputs(1275) <= not(layer0_outputs(10350)) or (layer0_outputs(7257));
    outputs(1276) <= not(layer0_outputs(10284)) or (layer0_outputs(2613));
    outputs(1277) <= layer0_outputs(9603);
    outputs(1278) <= not(layer0_outputs(3420));
    outputs(1279) <= not(layer0_outputs(4260));
    outputs(1280) <= (layer0_outputs(7017)) and not (layer0_outputs(2317));
    outputs(1281) <= not((layer0_outputs(5137)) or (layer0_outputs(70)));
    outputs(1282) <= (layer0_outputs(10524)) and not (layer0_outputs(4785));
    outputs(1283) <= (layer0_outputs(12221)) and (layer0_outputs(10459));
    outputs(1284) <= (layer0_outputs(3796)) xor (layer0_outputs(9872));
    outputs(1285) <= layer0_outputs(3596);
    outputs(1286) <= (layer0_outputs(2121)) xor (layer0_outputs(5806));
    outputs(1287) <= not((layer0_outputs(8060)) or (layer0_outputs(2977)));
    outputs(1288) <= layer0_outputs(2855);
    outputs(1289) <= (layer0_outputs(10159)) xor (layer0_outputs(3409));
    outputs(1290) <= (layer0_outputs(11454)) and (layer0_outputs(14));
    outputs(1291) <= (layer0_outputs(7986)) xor (layer0_outputs(1578));
    outputs(1292) <= (layer0_outputs(1747)) and not (layer0_outputs(98));
    outputs(1293) <= not((layer0_outputs(12261)) or (layer0_outputs(4509)));
    outputs(1294) <= (layer0_outputs(8469)) and (layer0_outputs(7099));
    outputs(1295) <= not((layer0_outputs(5022)) xor (layer0_outputs(10217)));
    outputs(1296) <= (layer0_outputs(8027)) and not (layer0_outputs(2373));
    outputs(1297) <= not((layer0_outputs(10361)) xor (layer0_outputs(11849)));
    outputs(1298) <= not(layer0_outputs(10464));
    outputs(1299) <= (layer0_outputs(7546)) xor (layer0_outputs(10460));
    outputs(1300) <= (layer0_outputs(8177)) and (layer0_outputs(10800));
    outputs(1301) <= not(layer0_outputs(8028));
    outputs(1302) <= layer0_outputs(8423);
    outputs(1303) <= not((layer0_outputs(399)) xor (layer0_outputs(10530)));
    outputs(1304) <= (layer0_outputs(10462)) and not (layer0_outputs(10417));
    outputs(1305) <= not((layer0_outputs(7744)) xor (layer0_outputs(5947)));
    outputs(1306) <= (layer0_outputs(7595)) and not (layer0_outputs(2364));
    outputs(1307) <= (layer0_outputs(11263)) and not (layer0_outputs(12029));
    outputs(1308) <= layer0_outputs(1199);
    outputs(1309) <= layer0_outputs(7735);
    outputs(1310) <= (layer0_outputs(813)) xor (layer0_outputs(2052));
    outputs(1311) <= not((layer0_outputs(7881)) or (layer0_outputs(10626)));
    outputs(1312) <= layer0_outputs(10650);
    outputs(1313) <= (layer0_outputs(1909)) and not (layer0_outputs(11874));
    outputs(1314) <= not(layer0_outputs(7022));
    outputs(1315) <= not(layer0_outputs(6880));
    outputs(1316) <= not((layer0_outputs(478)) xor (layer0_outputs(3340)));
    outputs(1317) <= not(layer0_outputs(6388));
    outputs(1318) <= not((layer0_outputs(11455)) xor (layer0_outputs(7430)));
    outputs(1319) <= not(layer0_outputs(7421));
    outputs(1320) <= not(layer0_outputs(2417));
    outputs(1321) <= not((layer0_outputs(1907)) or (layer0_outputs(12675)));
    outputs(1322) <= not((layer0_outputs(4865)) or (layer0_outputs(10871)));
    outputs(1323) <= not((layer0_outputs(222)) or (layer0_outputs(7795)));
    outputs(1324) <= layer0_outputs(9121);
    outputs(1325) <= not(layer0_outputs(11279));
    outputs(1326) <= not((layer0_outputs(7928)) xor (layer0_outputs(2120)));
    outputs(1327) <= not(layer0_outputs(4636));
    outputs(1328) <= (layer0_outputs(12394)) and not (layer0_outputs(8389));
    outputs(1329) <= layer0_outputs(6852);
    outputs(1330) <= (layer0_outputs(11183)) and not (layer0_outputs(8710));
    outputs(1331) <= not(layer0_outputs(7004));
    outputs(1332) <= (layer0_outputs(7724)) and not (layer0_outputs(69));
    outputs(1333) <= layer0_outputs(176);
    outputs(1334) <= layer0_outputs(5750);
    outputs(1335) <= not((layer0_outputs(400)) xor (layer0_outputs(9316)));
    outputs(1336) <= (layer0_outputs(3375)) and not (layer0_outputs(5157));
    outputs(1337) <= (layer0_outputs(5809)) and (layer0_outputs(3344));
    outputs(1338) <= (layer0_outputs(2867)) xor (layer0_outputs(7945));
    outputs(1339) <= layer0_outputs(9948);
    outputs(1340) <= (layer0_outputs(2010)) and (layer0_outputs(2383));
    outputs(1341) <= not((layer0_outputs(7208)) xor (layer0_outputs(2876)));
    outputs(1342) <= not((layer0_outputs(6794)) xor (layer0_outputs(6019)));
    outputs(1343) <= (layer0_outputs(9709)) and not (layer0_outputs(8201));
    outputs(1344) <= (layer0_outputs(3520)) and (layer0_outputs(4324));
    outputs(1345) <= (layer0_outputs(12489)) xor (layer0_outputs(6886));
    outputs(1346) <= not(layer0_outputs(10141));
    outputs(1347) <= (layer0_outputs(1825)) and not (layer0_outputs(11069));
    outputs(1348) <= '0';
    outputs(1349) <= (layer0_outputs(6154)) xor (layer0_outputs(9101));
    outputs(1350) <= not(layer0_outputs(9116));
    outputs(1351) <= layer0_outputs(3466);
    outputs(1352) <= not((layer0_outputs(1038)) xor (layer0_outputs(9744)));
    outputs(1353) <= not(layer0_outputs(2690));
    outputs(1354) <= (layer0_outputs(9819)) and (layer0_outputs(10680));
    outputs(1355) <= not((layer0_outputs(7516)) xor (layer0_outputs(2836)));
    outputs(1356) <= (layer0_outputs(697)) xor (layer0_outputs(10015));
    outputs(1357) <= layer0_outputs(11287);
    outputs(1358) <= (layer0_outputs(1723)) and not (layer0_outputs(4930));
    outputs(1359) <= layer0_outputs(2853);
    outputs(1360) <= (layer0_outputs(11848)) xor (layer0_outputs(928));
    outputs(1361) <= not((layer0_outputs(8853)) or (layer0_outputs(10409)));
    outputs(1362) <= not(layer0_outputs(1423));
    outputs(1363) <= not((layer0_outputs(9093)) xor (layer0_outputs(1330)));
    outputs(1364) <= not(layer0_outputs(11614));
    outputs(1365) <= (layer0_outputs(948)) xor (layer0_outputs(11893));
    outputs(1366) <= (layer0_outputs(2593)) xor (layer0_outputs(4320));
    outputs(1367) <= not(layer0_outputs(3892)) or (layer0_outputs(6288));
    outputs(1368) <= (layer0_outputs(5974)) xor (layer0_outputs(11579));
    outputs(1369) <= (layer0_outputs(9629)) and not (layer0_outputs(12742));
    outputs(1370) <= (layer0_outputs(3520)) xor (layer0_outputs(9375));
    outputs(1371) <= not((layer0_outputs(7678)) or (layer0_outputs(1260)));
    outputs(1372) <= not((layer0_outputs(372)) or (layer0_outputs(3023)));
    outputs(1373) <= not(layer0_outputs(1581));
    outputs(1374) <= not(layer0_outputs(9225));
    outputs(1375) <= not(layer0_outputs(4037));
    outputs(1376) <= not((layer0_outputs(9575)) xor (layer0_outputs(8282)));
    outputs(1377) <= not((layer0_outputs(4464)) xor (layer0_outputs(7052)));
    outputs(1378) <= (layer0_outputs(10032)) xor (layer0_outputs(11634));
    outputs(1379) <= not(layer0_outputs(6772));
    outputs(1380) <= not(layer0_outputs(6558));
    outputs(1381) <= not((layer0_outputs(2615)) or (layer0_outputs(10076)));
    outputs(1382) <= not(layer0_outputs(9488));
    outputs(1383) <= (layer0_outputs(11947)) xor (layer0_outputs(11747));
    outputs(1384) <= (layer0_outputs(8534)) or (layer0_outputs(4658));
    outputs(1385) <= not(layer0_outputs(9745));
    outputs(1386) <= not((layer0_outputs(1800)) xor (layer0_outputs(2725)));
    outputs(1387) <= layer0_outputs(12181);
    outputs(1388) <= not((layer0_outputs(2268)) or (layer0_outputs(1506)));
    outputs(1389) <= not((layer0_outputs(6123)) xor (layer0_outputs(6951)));
    outputs(1390) <= not((layer0_outputs(8605)) xor (layer0_outputs(941)));
    outputs(1391) <= not((layer0_outputs(4005)) or (layer0_outputs(7143)));
    outputs(1392) <= not((layer0_outputs(8229)) or (layer0_outputs(12734)));
    outputs(1393) <= layer0_outputs(11234);
    outputs(1394) <= not((layer0_outputs(12723)) or (layer0_outputs(11846)));
    outputs(1395) <= not(layer0_outputs(3535));
    outputs(1396) <= not(layer0_outputs(3067));
    outputs(1397) <= (layer0_outputs(2783)) and not (layer0_outputs(361));
    outputs(1398) <= not((layer0_outputs(2957)) xor (layer0_outputs(11066)));
    outputs(1399) <= not((layer0_outputs(10147)) or (layer0_outputs(12307)));
    outputs(1400) <= layer0_outputs(6758);
    outputs(1401) <= (layer0_outputs(7282)) and not (layer0_outputs(12273));
    outputs(1402) <= not(layer0_outputs(1014));
    outputs(1403) <= not((layer0_outputs(5188)) or (layer0_outputs(4387)));
    outputs(1404) <= not((layer0_outputs(10294)) xor (layer0_outputs(10736)));
    outputs(1405) <= not((layer0_outputs(7190)) xor (layer0_outputs(8445)));
    outputs(1406) <= layer0_outputs(2546);
    outputs(1407) <= not((layer0_outputs(9768)) xor (layer0_outputs(77)));
    outputs(1408) <= not((layer0_outputs(12761)) xor (layer0_outputs(10994)));
    outputs(1409) <= layer0_outputs(11448);
    outputs(1410) <= (layer0_outputs(2389)) xor (layer0_outputs(12767));
    outputs(1411) <= (layer0_outputs(1764)) and (layer0_outputs(7717));
    outputs(1412) <= layer0_outputs(5521);
    outputs(1413) <= (layer0_outputs(5492)) and (layer0_outputs(8540));
    outputs(1414) <= layer0_outputs(5494);
    outputs(1415) <= (layer0_outputs(3473)) and (layer0_outputs(3769));
    outputs(1416) <= (layer0_outputs(701)) and not (layer0_outputs(4086));
    outputs(1417) <= not(layer0_outputs(12180));
    outputs(1418) <= (layer0_outputs(8203)) and not (layer0_outputs(4400));
    outputs(1419) <= layer0_outputs(12437);
    outputs(1420) <= (layer0_outputs(1300)) and not (layer0_outputs(6874));
    outputs(1421) <= (layer0_outputs(4984)) and not (layer0_outputs(9260));
    outputs(1422) <= layer0_outputs(9002);
    outputs(1423) <= not((layer0_outputs(7179)) or (layer0_outputs(5278)));
    outputs(1424) <= (layer0_outputs(2329)) and not (layer0_outputs(4210));
    outputs(1425) <= layer0_outputs(1852);
    outputs(1426) <= layer0_outputs(5276);
    outputs(1427) <= (layer0_outputs(8957)) and not (layer0_outputs(11050));
    outputs(1428) <= not((layer0_outputs(7871)) or (layer0_outputs(9523)));
    outputs(1429) <= '0';
    outputs(1430) <= (layer0_outputs(1063)) and (layer0_outputs(11829));
    outputs(1431) <= not((layer0_outputs(12376)) or (layer0_outputs(818)));
    outputs(1432) <= layer0_outputs(2561);
    outputs(1433) <= not(layer0_outputs(2078));
    outputs(1434) <= layer0_outputs(10186);
    outputs(1435) <= (layer0_outputs(1680)) and not (layer0_outputs(423));
    outputs(1436) <= not((layer0_outputs(8560)) or (layer0_outputs(12264)));
    outputs(1437) <= not((layer0_outputs(2051)) or (layer0_outputs(10387)));
    outputs(1438) <= (layer0_outputs(1590)) and (layer0_outputs(6226));
    outputs(1439) <= (layer0_outputs(4661)) and (layer0_outputs(2163));
    outputs(1440) <= (layer0_outputs(3871)) and (layer0_outputs(3786));
    outputs(1441) <= layer0_outputs(4172);
    outputs(1442) <= not((layer0_outputs(8082)) xor (layer0_outputs(5515)));
    outputs(1443) <= (layer0_outputs(8237)) and not (layer0_outputs(10157));
    outputs(1444) <= not((layer0_outputs(1282)) or (layer0_outputs(11291)));
    outputs(1445) <= (layer0_outputs(12397)) and not (layer0_outputs(52));
    outputs(1446) <= layer0_outputs(6728);
    outputs(1447) <= not((layer0_outputs(4218)) or (layer0_outputs(2263)));
    outputs(1448) <= (layer0_outputs(1091)) and not (layer0_outputs(6068));
    outputs(1449) <= (layer0_outputs(11998)) and not (layer0_outputs(6322));
    outputs(1450) <= not((layer0_outputs(1635)) xor (layer0_outputs(2560)));
    outputs(1451) <= not(layer0_outputs(11274)) or (layer0_outputs(11222));
    outputs(1452) <= (layer0_outputs(8651)) and not (layer0_outputs(6654));
    outputs(1453) <= layer0_outputs(10020);
    outputs(1454) <= layer0_outputs(9596);
    outputs(1455) <= (layer0_outputs(6198)) and not (layer0_outputs(3344));
    outputs(1456) <= (layer0_outputs(11588)) and not (layer0_outputs(2441));
    outputs(1457) <= (layer0_outputs(4317)) and not (layer0_outputs(3917));
    outputs(1458) <= (layer0_outputs(8308)) xor (layer0_outputs(6323));
    outputs(1459) <= (layer0_outputs(9571)) and not (layer0_outputs(1122));
    outputs(1460) <= layer0_outputs(8809);
    outputs(1461) <= not(layer0_outputs(6956));
    outputs(1462) <= (layer0_outputs(11014)) xor (layer0_outputs(10869));
    outputs(1463) <= not(layer0_outputs(8586));
    outputs(1464) <= (layer0_outputs(151)) and not (layer0_outputs(8520));
    outputs(1465) <= not((layer0_outputs(10569)) xor (layer0_outputs(2811)));
    outputs(1466) <= layer0_outputs(4220);
    outputs(1467) <= (layer0_outputs(6338)) and not (layer0_outputs(4786));
    outputs(1468) <= not(layer0_outputs(621));
    outputs(1469) <= (layer0_outputs(11102)) and not (layer0_outputs(691));
    outputs(1470) <= not((layer0_outputs(11078)) xor (layer0_outputs(1574)));
    outputs(1471) <= (layer0_outputs(12427)) and (layer0_outputs(470));
    outputs(1472) <= not(layer0_outputs(10156));
    outputs(1473) <= (layer0_outputs(176)) and not (layer0_outputs(11410));
    outputs(1474) <= layer0_outputs(2398);
    outputs(1475) <= (layer0_outputs(1884)) or (layer0_outputs(5901));
    outputs(1476) <= (layer0_outputs(7056)) and not (layer0_outputs(5643));
    outputs(1477) <= not(layer0_outputs(7831));
    outputs(1478) <= (layer0_outputs(8902)) and not (layer0_outputs(9810));
    outputs(1479) <= (layer0_outputs(11372)) and (layer0_outputs(10135));
    outputs(1480) <= layer0_outputs(12787);
    outputs(1481) <= (layer0_outputs(12106)) and not (layer0_outputs(257));
    outputs(1482) <= (layer0_outputs(7530)) xor (layer0_outputs(1659));
    outputs(1483) <= not(layer0_outputs(2225));
    outputs(1484) <= not(layer0_outputs(8143)) or (layer0_outputs(4351));
    outputs(1485) <= layer0_outputs(61);
    outputs(1486) <= layer0_outputs(9341);
    outputs(1487) <= not((layer0_outputs(197)) or (layer0_outputs(2693)));
    outputs(1488) <= not((layer0_outputs(9809)) or (layer0_outputs(9750)));
    outputs(1489) <= layer0_outputs(3351);
    outputs(1490) <= (layer0_outputs(2386)) and not (layer0_outputs(1215));
    outputs(1491) <= not((layer0_outputs(12598)) xor (layer0_outputs(10729)));
    outputs(1492) <= (layer0_outputs(1572)) xor (layer0_outputs(7005));
    outputs(1493) <= not(layer0_outputs(3667));
    outputs(1494) <= (layer0_outputs(5374)) and not (layer0_outputs(11201));
    outputs(1495) <= layer0_outputs(12701);
    outputs(1496) <= (layer0_outputs(8622)) and (layer0_outputs(2768));
    outputs(1497) <= layer0_outputs(7075);
    outputs(1498) <= not((layer0_outputs(12538)) or (layer0_outputs(1636)));
    outputs(1499) <= not(layer0_outputs(6527));
    outputs(1500) <= layer0_outputs(11568);
    outputs(1501) <= layer0_outputs(9475);
    outputs(1502) <= layer0_outputs(2169);
    outputs(1503) <= not((layer0_outputs(94)) xor (layer0_outputs(12017)));
    outputs(1504) <= not((layer0_outputs(9729)) xor (layer0_outputs(3374)));
    outputs(1505) <= layer0_outputs(3061);
    outputs(1506) <= not(layer0_outputs(4443));
    outputs(1507) <= not((layer0_outputs(263)) xor (layer0_outputs(6697)));
    outputs(1508) <= '0';
    outputs(1509) <= (layer0_outputs(1887)) xor (layer0_outputs(3974));
    outputs(1510) <= (layer0_outputs(10794)) and (layer0_outputs(1018));
    outputs(1511) <= not(layer0_outputs(8038));
    outputs(1512) <= (layer0_outputs(3738)) and not (layer0_outputs(7566));
    outputs(1513) <= not((layer0_outputs(5726)) or (layer0_outputs(1267)));
    outputs(1514) <= (layer0_outputs(12224)) and not (layer0_outputs(4772));
    outputs(1515) <= not((layer0_outputs(5879)) xor (layer0_outputs(2890)));
    outputs(1516) <= not((layer0_outputs(1716)) xor (layer0_outputs(3290)));
    outputs(1517) <= layer0_outputs(1974);
    outputs(1518) <= (layer0_outputs(2986)) and (layer0_outputs(8706));
    outputs(1519) <= (layer0_outputs(1010)) and (layer0_outputs(11825));
    outputs(1520) <= layer0_outputs(10351);
    outputs(1521) <= not(layer0_outputs(1042));
    outputs(1522) <= (layer0_outputs(6628)) xor (layer0_outputs(482));
    outputs(1523) <= layer0_outputs(12431);
    outputs(1524) <= not(layer0_outputs(5484));
    outputs(1525) <= layer0_outputs(1622);
    outputs(1526) <= (layer0_outputs(91)) and (layer0_outputs(4844));
    outputs(1527) <= (layer0_outputs(10107)) and not (layer0_outputs(4733));
    outputs(1528) <= (layer0_outputs(4081)) and (layer0_outputs(9305));
    outputs(1529) <= (layer0_outputs(4645)) and not (layer0_outputs(3));
    outputs(1530) <= (layer0_outputs(7739)) and not (layer0_outputs(3621));
    outputs(1531) <= (layer0_outputs(5910)) and not (layer0_outputs(4710));
    outputs(1532) <= (layer0_outputs(12182)) and (layer0_outputs(11283));
    outputs(1533) <= (layer0_outputs(6426)) and not (layer0_outputs(5831));
    outputs(1534) <= not((layer0_outputs(5460)) xor (layer0_outputs(2289)));
    outputs(1535) <= not((layer0_outputs(3149)) or (layer0_outputs(11639)));
    outputs(1536) <= not((layer0_outputs(6909)) xor (layer0_outputs(3251)));
    outputs(1537) <= not(layer0_outputs(4476)) or (layer0_outputs(11495));
    outputs(1538) <= layer0_outputs(11439);
    outputs(1539) <= layer0_outputs(5682);
    outputs(1540) <= (layer0_outputs(1546)) and not (layer0_outputs(12579));
    outputs(1541) <= (layer0_outputs(1872)) and not (layer0_outputs(3056));
    outputs(1542) <= (layer0_outputs(6691)) xor (layer0_outputs(7943));
    outputs(1543) <= layer0_outputs(10599);
    outputs(1544) <= (layer0_outputs(3427)) and not (layer0_outputs(9007));
    outputs(1545) <= (layer0_outputs(7324)) and not (layer0_outputs(11976));
    outputs(1546) <= not((layer0_outputs(5873)) xor (layer0_outputs(6086)));
    outputs(1547) <= (layer0_outputs(7500)) and not (layer0_outputs(12460));
    outputs(1548) <= (layer0_outputs(2142)) and not (layer0_outputs(8218));
    outputs(1549) <= (layer0_outputs(10336)) and (layer0_outputs(1895));
    outputs(1550) <= not((layer0_outputs(11659)) or (layer0_outputs(731)));
    outputs(1551) <= layer0_outputs(4971);
    outputs(1552) <= not((layer0_outputs(6993)) xor (layer0_outputs(11327)));
    outputs(1553) <= not((layer0_outputs(10488)) xor (layer0_outputs(5386)));
    outputs(1554) <= not(layer0_outputs(6694));
    outputs(1555) <= '0';
    outputs(1556) <= (layer0_outputs(9174)) xor (layer0_outputs(7457));
    outputs(1557) <= not(layer0_outputs(4859));
    outputs(1558) <= not((layer0_outputs(3571)) xor (layer0_outputs(2822)));
    outputs(1559) <= (layer0_outputs(7844)) and not (layer0_outputs(6135));
    outputs(1560) <= not((layer0_outputs(3463)) or (layer0_outputs(2272)));
    outputs(1561) <= layer0_outputs(6288);
    outputs(1562) <= (layer0_outputs(1524)) xor (layer0_outputs(11864));
    outputs(1563) <= (layer0_outputs(2182)) and not (layer0_outputs(8857));
    outputs(1564) <= (layer0_outputs(10791)) xor (layer0_outputs(7334));
    outputs(1565) <= not((layer0_outputs(6038)) or (layer0_outputs(1344)));
    outputs(1566) <= not(layer0_outputs(6561)) or (layer0_outputs(3586));
    outputs(1567) <= layer0_outputs(3158);
    outputs(1568) <= not((layer0_outputs(1126)) or (layer0_outputs(4309)));
    outputs(1569) <= not((layer0_outputs(8883)) xor (layer0_outputs(3229)));
    outputs(1570) <= (layer0_outputs(1881)) and not (layer0_outputs(2873));
    outputs(1571) <= (layer0_outputs(3815)) and (layer0_outputs(2231));
    outputs(1572) <= not((layer0_outputs(8648)) xor (layer0_outputs(2035)));
    outputs(1573) <= (layer0_outputs(8048)) xor (layer0_outputs(11511));
    outputs(1574) <= (layer0_outputs(12310)) and not (layer0_outputs(7783));
    outputs(1575) <= layer0_outputs(8907);
    outputs(1576) <= not(layer0_outputs(5045));
    outputs(1577) <= not(layer0_outputs(3610));
    outputs(1578) <= layer0_outputs(6174);
    outputs(1579) <= layer0_outputs(188);
    outputs(1580) <= layer0_outputs(3171);
    outputs(1581) <= not((layer0_outputs(6519)) xor (layer0_outputs(3869)));
    outputs(1582) <= not(layer0_outputs(2433));
    outputs(1583) <= (layer0_outputs(5988)) xor (layer0_outputs(6193));
    outputs(1584) <= (layer0_outputs(605)) and not (layer0_outputs(5005));
    outputs(1585) <= (layer0_outputs(10429)) and not (layer0_outputs(7798));
    outputs(1586) <= (layer0_outputs(9848)) and not (layer0_outputs(9381));
    outputs(1587) <= layer0_outputs(9868);
    outputs(1588) <= not(layer0_outputs(10325));
    outputs(1589) <= not(layer0_outputs(10458)) or (layer0_outputs(3502));
    outputs(1590) <= layer0_outputs(12211);
    outputs(1591) <= (layer0_outputs(3877)) xor (layer0_outputs(6602));
    outputs(1592) <= not(layer0_outputs(6767));
    outputs(1593) <= not((layer0_outputs(4755)) or (layer0_outputs(9646)));
    outputs(1594) <= layer0_outputs(8851);
    outputs(1595) <= (layer0_outputs(7090)) and not (layer0_outputs(5399));
    outputs(1596) <= layer0_outputs(10579);
    outputs(1597) <= (layer0_outputs(7387)) and (layer0_outputs(8291));
    outputs(1598) <= (layer0_outputs(4704)) and (layer0_outputs(9068));
    outputs(1599) <= layer0_outputs(9585);
    outputs(1600) <= (layer0_outputs(11421)) and (layer0_outputs(1419));
    outputs(1601) <= (layer0_outputs(6310)) and not (layer0_outputs(7280));
    outputs(1602) <= not(layer0_outputs(2012));
    outputs(1603) <= (layer0_outputs(6833)) and (layer0_outputs(8730));
    outputs(1604) <= not(layer0_outputs(2143));
    outputs(1605) <= not((layer0_outputs(3414)) or (layer0_outputs(80)));
    outputs(1606) <= not(layer0_outputs(6675));
    outputs(1607) <= not((layer0_outputs(11175)) or (layer0_outputs(10659)));
    outputs(1608) <= layer0_outputs(11691);
    outputs(1609) <= (layer0_outputs(5373)) and not (layer0_outputs(9547));
    outputs(1610) <= layer0_outputs(7298);
    outputs(1611) <= (layer0_outputs(3529)) and (layer0_outputs(9632));
    outputs(1612) <= layer0_outputs(1199);
    outputs(1613) <= not(layer0_outputs(6218));
    outputs(1614) <= (layer0_outputs(1769)) and not (layer0_outputs(11909));
    outputs(1615) <= (layer0_outputs(4922)) and (layer0_outputs(7101));
    outputs(1616) <= not((layer0_outputs(23)) xor (layer0_outputs(5042)));
    outputs(1617) <= (layer0_outputs(4364)) xor (layer0_outputs(7374));
    outputs(1618) <= not(layer0_outputs(12379));
    outputs(1619) <= not((layer0_outputs(5026)) or (layer0_outputs(12312)));
    outputs(1620) <= (layer0_outputs(10754)) xor (layer0_outputs(1304));
    outputs(1621) <= not(layer0_outputs(267));
    outputs(1622) <= layer0_outputs(6751);
    outputs(1623) <= not(layer0_outputs(7440)) or (layer0_outputs(9396));
    outputs(1624) <= not(layer0_outputs(8646));
    outputs(1625) <= not(layer0_outputs(2521));
    outputs(1626) <= not(layer0_outputs(5339));
    outputs(1627) <= not(layer0_outputs(770));
    outputs(1628) <= not(layer0_outputs(11166));
    outputs(1629) <= not((layer0_outputs(8469)) xor (layer0_outputs(2341)));
    outputs(1630) <= not(layer0_outputs(7287));
    outputs(1631) <= not(layer0_outputs(1882));
    outputs(1632) <= not(layer0_outputs(1071));
    outputs(1633) <= '0';
    outputs(1634) <= (layer0_outputs(4891)) and not (layer0_outputs(9605));
    outputs(1635) <= (layer0_outputs(12450)) and (layer0_outputs(10925));
    outputs(1636) <= not(layer0_outputs(2696));
    outputs(1637) <= not((layer0_outputs(7089)) xor (layer0_outputs(12428)));
    outputs(1638) <= not(layer0_outputs(2217));
    outputs(1639) <= not((layer0_outputs(1340)) or (layer0_outputs(9194)));
    outputs(1640) <= '1';
    outputs(1641) <= not((layer0_outputs(8066)) xor (layer0_outputs(853)));
    outputs(1642) <= (layer0_outputs(9026)) and not (layer0_outputs(10709));
    outputs(1643) <= (layer0_outputs(11964)) and not (layer0_outputs(4556));
    outputs(1644) <= not((layer0_outputs(680)) xor (layer0_outputs(2564)));
    outputs(1645) <= layer0_outputs(1034);
    outputs(1646) <= (layer0_outputs(6581)) and (layer0_outputs(9035));
    outputs(1647) <= (layer0_outputs(4909)) and not (layer0_outputs(1118));
    outputs(1648) <= (layer0_outputs(9883)) xor (layer0_outputs(7407));
    outputs(1649) <= layer0_outputs(148);
    outputs(1650) <= (layer0_outputs(6102)) and (layer0_outputs(9977));
    outputs(1651) <= (layer0_outputs(8206)) and not (layer0_outputs(3257));
    outputs(1652) <= layer0_outputs(899);
    outputs(1653) <= '0';
    outputs(1654) <= not(layer0_outputs(9569));
    outputs(1655) <= (layer0_outputs(9988)) and (layer0_outputs(9979));
    outputs(1656) <= (layer0_outputs(4780)) and not (layer0_outputs(5163));
    outputs(1657) <= layer0_outputs(12289);
    outputs(1658) <= not(layer0_outputs(5761));
    outputs(1659) <= (layer0_outputs(5648)) and not (layer0_outputs(9084));
    outputs(1660) <= (layer0_outputs(11125)) and (layer0_outputs(1189));
    outputs(1661) <= (layer0_outputs(90)) and not (layer0_outputs(10565));
    outputs(1662) <= layer0_outputs(6962);
    outputs(1663) <= (layer0_outputs(273)) and not (layer0_outputs(2140));
    outputs(1664) <= '0';
    outputs(1665) <= (layer0_outputs(4275)) xor (layer0_outputs(678));
    outputs(1666) <= (layer0_outputs(7160)) and not (layer0_outputs(10743));
    outputs(1667) <= not((layer0_outputs(9135)) xor (layer0_outputs(11542)));
    outputs(1668) <= '0';
    outputs(1669) <= layer0_outputs(12084);
    outputs(1670) <= (layer0_outputs(1804)) xor (layer0_outputs(11268));
    outputs(1671) <= layer0_outputs(8436);
    outputs(1672) <= (layer0_outputs(4367)) and not (layer0_outputs(5389));
    outputs(1673) <= (layer0_outputs(4868)) xor (layer0_outputs(3678));
    outputs(1674) <= (layer0_outputs(5348)) xor (layer0_outputs(1418));
    outputs(1675) <= not(layer0_outputs(3750));
    outputs(1676) <= not(layer0_outputs(11532));
    outputs(1677) <= not((layer0_outputs(10856)) xor (layer0_outputs(12024)));
    outputs(1678) <= (layer0_outputs(8266)) and not (layer0_outputs(8939));
    outputs(1679) <= not(layer0_outputs(11791));
    outputs(1680) <= layer0_outputs(4322);
    outputs(1681) <= (layer0_outputs(3090)) xor (layer0_outputs(9451));
    outputs(1682) <= not(layer0_outputs(11472));
    outputs(1683) <= (layer0_outputs(4336)) xor (layer0_outputs(3615));
    outputs(1684) <= (layer0_outputs(510)) xor (layer0_outputs(288));
    outputs(1685) <= not(layer0_outputs(924));
    outputs(1686) <= (layer0_outputs(7840)) xor (layer0_outputs(6881));
    outputs(1687) <= (layer0_outputs(5697)) xor (layer0_outputs(8985));
    outputs(1688) <= not((layer0_outputs(6594)) or (layer0_outputs(9046)));
    outputs(1689) <= (layer0_outputs(8433)) and not (layer0_outputs(8400));
    outputs(1690) <= layer0_outputs(1469);
    outputs(1691) <= not((layer0_outputs(8092)) xor (layer0_outputs(5872)));
    outputs(1692) <= not(layer0_outputs(7843));
    outputs(1693) <= not(layer0_outputs(10052));
    outputs(1694) <= not((layer0_outputs(9592)) or (layer0_outputs(5393)));
    outputs(1695) <= (layer0_outputs(3649)) and not (layer0_outputs(5993));
    outputs(1696) <= (layer0_outputs(10230)) and not (layer0_outputs(6937));
    outputs(1697) <= not((layer0_outputs(12607)) xor (layer0_outputs(9761)));
    outputs(1698) <= not((layer0_outputs(6827)) xor (layer0_outputs(1839)));
    outputs(1699) <= (layer0_outputs(8799)) and not (layer0_outputs(12332));
    outputs(1700) <= not((layer0_outputs(2735)) xor (layer0_outputs(858)));
    outputs(1701) <= not((layer0_outputs(10072)) or (layer0_outputs(7031)));
    outputs(1702) <= (layer0_outputs(9035)) and not (layer0_outputs(5945));
    outputs(1703) <= (layer0_outputs(12455)) and not (layer0_outputs(4485));
    outputs(1704) <= not((layer0_outputs(3578)) xor (layer0_outputs(11170)));
    outputs(1705) <= (layer0_outputs(9801)) and (layer0_outputs(1030));
    outputs(1706) <= (layer0_outputs(9476)) and not (layer0_outputs(5489));
    outputs(1707) <= (layer0_outputs(11068)) and not (layer0_outputs(8079));
    outputs(1708) <= (layer0_outputs(12786)) and not (layer0_outputs(5423));
    outputs(1709) <= not((layer0_outputs(5438)) xor (layer0_outputs(10343)));
    outputs(1710) <= (layer0_outputs(7767)) xor (layer0_outputs(2482));
    outputs(1711) <= not(layer0_outputs(9633));
    outputs(1712) <= not((layer0_outputs(3912)) xor (layer0_outputs(6255)));
    outputs(1713) <= not(layer0_outputs(3517));
    outputs(1714) <= '0';
    outputs(1715) <= layer0_outputs(9286);
    outputs(1716) <= not(layer0_outputs(10766));
    outputs(1717) <= (layer0_outputs(918)) and not (layer0_outputs(10605));
    outputs(1718) <= (layer0_outputs(12600)) xor (layer0_outputs(12287));
    outputs(1719) <= '0';
    outputs(1720) <= (layer0_outputs(6056)) and not (layer0_outputs(541));
    outputs(1721) <= layer0_outputs(7014);
    outputs(1722) <= (layer0_outputs(3195)) xor (layer0_outputs(10559));
    outputs(1723) <= (layer0_outputs(8618)) and not (layer0_outputs(9051));
    outputs(1724) <= not((layer0_outputs(9810)) or (layer0_outputs(2718)));
    outputs(1725) <= not((layer0_outputs(7109)) or (layer0_outputs(9152)));
    outputs(1726) <= not(layer0_outputs(7938));
    outputs(1727) <= (layer0_outputs(12282)) xor (layer0_outputs(146));
    outputs(1728) <= not(layer0_outputs(5364));
    outputs(1729) <= not((layer0_outputs(8252)) xor (layer0_outputs(4239)));
    outputs(1730) <= layer0_outputs(499);
    outputs(1731) <= not((layer0_outputs(464)) xor (layer0_outputs(9377)));
    outputs(1732) <= layer0_outputs(4404);
    outputs(1733) <= (layer0_outputs(5709)) and not (layer0_outputs(9276));
    outputs(1734) <= (layer0_outputs(3032)) and not (layer0_outputs(10722));
    outputs(1735) <= not((layer0_outputs(7903)) xor (layer0_outputs(9836)));
    outputs(1736) <= (layer0_outputs(1908)) and not (layer0_outputs(2240));
    outputs(1737) <= layer0_outputs(7981);
    outputs(1738) <= (layer0_outputs(9794)) xor (layer0_outputs(6058));
    outputs(1739) <= layer0_outputs(9929);
    outputs(1740) <= (layer0_outputs(7021)) and not (layer0_outputs(11152));
    outputs(1741) <= (layer0_outputs(6687)) and (layer0_outputs(2365));
    outputs(1742) <= (layer0_outputs(7210)) and not (layer0_outputs(10598));
    outputs(1743) <= (layer0_outputs(741)) xor (layer0_outputs(6312));
    outputs(1744) <= not((layer0_outputs(9139)) xor (layer0_outputs(1682)));
    outputs(1745) <= not(layer0_outputs(4271));
    outputs(1746) <= not((layer0_outputs(591)) xor (layer0_outputs(9107)));
    outputs(1747) <= (layer0_outputs(5293)) and (layer0_outputs(5117));
    outputs(1748) <= not((layer0_outputs(1543)) xor (layer0_outputs(11250)));
    outputs(1749) <= not((layer0_outputs(11693)) xor (layer0_outputs(4572)));
    outputs(1750) <= (layer0_outputs(10309)) xor (layer0_outputs(3910));
    outputs(1751) <= (layer0_outputs(2718)) and (layer0_outputs(396));
    outputs(1752) <= not((layer0_outputs(10207)) xor (layer0_outputs(12065)));
    outputs(1753) <= not(layer0_outputs(3600));
    outputs(1754) <= '0';
    outputs(1755) <= '0';
    outputs(1756) <= (layer0_outputs(11340)) xor (layer0_outputs(4678));
    outputs(1757) <= (layer0_outputs(8186)) xor (layer0_outputs(10146));
    outputs(1758) <= (layer0_outputs(4778)) and not (layer0_outputs(4555));
    outputs(1759) <= not(layer0_outputs(2901));
    outputs(1760) <= not(layer0_outputs(9772));
    outputs(1761) <= (layer0_outputs(519)) and not (layer0_outputs(8403));
    outputs(1762) <= '0';
    outputs(1763) <= (layer0_outputs(6066)) and (layer0_outputs(2866));
    outputs(1764) <= not(layer0_outputs(2685));
    outputs(1765) <= (layer0_outputs(1673)) and not (layer0_outputs(5190));
    outputs(1766) <= layer0_outputs(9213);
    outputs(1767) <= not((layer0_outputs(12121)) xor (layer0_outputs(8189)));
    outputs(1768) <= (layer0_outputs(2176)) xor (layer0_outputs(5860));
    outputs(1769) <= (layer0_outputs(11928)) xor (layer0_outputs(1704));
    outputs(1770) <= (layer0_outputs(8681)) and (layer0_outputs(12714));
    outputs(1771) <= (layer0_outputs(7935)) xor (layer0_outputs(1828));
    outputs(1772) <= not((layer0_outputs(9330)) xor (layer0_outputs(8236)));
    outputs(1773) <= (layer0_outputs(251)) and not (layer0_outputs(11879));
    outputs(1774) <= not((layer0_outputs(6283)) xor (layer0_outputs(8897)));
    outputs(1775) <= (layer0_outputs(6449)) and (layer0_outputs(333));
    outputs(1776) <= (layer0_outputs(9890)) xor (layer0_outputs(1788));
    outputs(1777) <= not(layer0_outputs(9066));
    outputs(1778) <= not((layer0_outputs(7260)) or (layer0_outputs(3253)));
    outputs(1779) <= not((layer0_outputs(688)) xor (layer0_outputs(5518)));
    outputs(1780) <= (layer0_outputs(968)) and not (layer0_outputs(5903));
    outputs(1781) <= (layer0_outputs(10653)) and not (layer0_outputs(6364));
    outputs(1782) <= (layer0_outputs(5619)) xor (layer0_outputs(1554));
    outputs(1783) <= (layer0_outputs(10019)) xor (layer0_outputs(6838));
    outputs(1784) <= layer0_outputs(775);
    outputs(1785) <= layer0_outputs(583);
    outputs(1786) <= layer0_outputs(4929);
    outputs(1787) <= (layer0_outputs(2713)) or (layer0_outputs(4328));
    outputs(1788) <= layer0_outputs(10959);
    outputs(1789) <= not((layer0_outputs(2248)) xor (layer0_outputs(2691)));
    outputs(1790) <= (layer0_outputs(2172)) and not (layer0_outputs(11698));
    outputs(1791) <= not((layer0_outputs(7624)) and (layer0_outputs(10872)));
    outputs(1792) <= not((layer0_outputs(5298)) xor (layer0_outputs(3568)));
    outputs(1793) <= not(layer0_outputs(1639)) or (layer0_outputs(2917));
    outputs(1794) <= (layer0_outputs(1578)) and not (layer0_outputs(5096));
    outputs(1795) <= not(layer0_outputs(8124));
    outputs(1796) <= not(layer0_outputs(8589));
    outputs(1797) <= (layer0_outputs(12191)) xor (layer0_outputs(12638));
    outputs(1798) <= (layer0_outputs(4830)) and not (layer0_outputs(2034));
    outputs(1799) <= not((layer0_outputs(8196)) xor (layer0_outputs(5458)));
    outputs(1800) <= layer0_outputs(3860);
    outputs(1801) <= (layer0_outputs(9733)) and not (layer0_outputs(6627));
    outputs(1802) <= not((layer0_outputs(5612)) xor (layer0_outputs(5138)));
    outputs(1803) <= not((layer0_outputs(5446)) xor (layer0_outputs(7608)));
    outputs(1804) <= (layer0_outputs(1666)) and not (layer0_outputs(946));
    outputs(1805) <= (layer0_outputs(2894)) and not (layer0_outputs(11349));
    outputs(1806) <= (layer0_outputs(2764)) and (layer0_outputs(8838));
    outputs(1807) <= (layer0_outputs(10313)) and not (layer0_outputs(2070));
    outputs(1808) <= not((layer0_outputs(8042)) or (layer0_outputs(10532)));
    outputs(1809) <= (layer0_outputs(3443)) xor (layer0_outputs(11249));
    outputs(1810) <= (layer0_outputs(2016)) and not (layer0_outputs(4409));
    outputs(1811) <= not((layer0_outputs(2375)) or (layer0_outputs(7855)));
    outputs(1812) <= '0';
    outputs(1813) <= not(layer0_outputs(2767));
    outputs(1814) <= not(layer0_outputs(1745));
    outputs(1815) <= not((layer0_outputs(11916)) or (layer0_outputs(2340)));
    outputs(1816) <= (layer0_outputs(9412)) and not (layer0_outputs(3879));
    outputs(1817) <= (layer0_outputs(12251)) xor (layer0_outputs(3797));
    outputs(1818) <= (layer0_outputs(10708)) and not (layer0_outputs(6555));
    outputs(1819) <= (layer0_outputs(9757)) and (layer0_outputs(149));
    outputs(1820) <= (layer0_outputs(10802)) and not (layer0_outputs(2631));
    outputs(1821) <= (layer0_outputs(8374)) and (layer0_outputs(11107));
    outputs(1822) <= (layer0_outputs(2338)) and (layer0_outputs(11813));
    outputs(1823) <= not(layer0_outputs(4712));
    outputs(1824) <= (layer0_outputs(2910)) and not (layer0_outputs(12103));
    outputs(1825) <= not(layer0_outputs(9125));
    outputs(1826) <= (layer0_outputs(7571)) xor (layer0_outputs(1085));
    outputs(1827) <= (layer0_outputs(71)) and (layer0_outputs(6136));
    outputs(1828) <= (layer0_outputs(9272)) xor (layer0_outputs(1782));
    outputs(1829) <= (layer0_outputs(4403)) xor (layer0_outputs(4326));
    outputs(1830) <= layer0_outputs(7904);
    outputs(1831) <= (layer0_outputs(7427)) and (layer0_outputs(1673));
    outputs(1832) <= not(layer0_outputs(225));
    outputs(1833) <= (layer0_outputs(9954)) and (layer0_outputs(11572));
    outputs(1834) <= layer0_outputs(5203);
    outputs(1835) <= (layer0_outputs(3510)) xor (layer0_outputs(4020));
    outputs(1836) <= (layer0_outputs(7992)) and (layer0_outputs(4977));
    outputs(1837) <= not((layer0_outputs(1867)) or (layer0_outputs(4673)));
    outputs(1838) <= (layer0_outputs(1875)) xor (layer0_outputs(5824));
    outputs(1839) <= (layer0_outputs(6584)) xor (layer0_outputs(1487));
    outputs(1840) <= (layer0_outputs(12756)) and not (layer0_outputs(6540));
    outputs(1841) <= not(layer0_outputs(8858)) or (layer0_outputs(5939));
    outputs(1842) <= not(layer0_outputs(11814));
    outputs(1843) <= not(layer0_outputs(7287)) or (layer0_outputs(10457));
    outputs(1844) <= (layer0_outputs(9575)) and not (layer0_outputs(5765));
    outputs(1845) <= (layer0_outputs(687)) xor (layer0_outputs(10956));
    outputs(1846) <= not((layer0_outputs(2419)) or (layer0_outputs(517)));
    outputs(1847) <= (layer0_outputs(1862)) and not (layer0_outputs(10211));
    outputs(1848) <= (layer0_outputs(9088)) and not (layer0_outputs(9992));
    outputs(1849) <= layer0_outputs(8754);
    outputs(1850) <= not((layer0_outputs(8890)) xor (layer0_outputs(2206)));
    outputs(1851) <= (layer0_outputs(12042)) and not (layer0_outputs(1855));
    outputs(1852) <= (layer0_outputs(8381)) and not (layer0_outputs(2360));
    outputs(1853) <= (layer0_outputs(6893)) and not (layer0_outputs(11918));
    outputs(1854) <= not((layer0_outputs(1187)) xor (layer0_outputs(8743)));
    outputs(1855) <= layer0_outputs(10996);
    outputs(1856) <= (layer0_outputs(992)) and (layer0_outputs(5496));
    outputs(1857) <= (layer0_outputs(834)) and not (layer0_outputs(6505));
    outputs(1858) <= not(layer0_outputs(2379));
    outputs(1859) <= not(layer0_outputs(8642));
    outputs(1860) <= '0';
    outputs(1861) <= layer0_outputs(11773);
    outputs(1862) <= not(layer0_outputs(7930));
    outputs(1863) <= not((layer0_outputs(1007)) xor (layer0_outputs(3734)));
    outputs(1864) <= '0';
    outputs(1865) <= not(layer0_outputs(11098));
    outputs(1866) <= not(layer0_outputs(2478));
    outputs(1867) <= layer0_outputs(5637);
    outputs(1868) <= not((layer0_outputs(1960)) or (layer0_outputs(9870)));
    outputs(1869) <= (layer0_outputs(1354)) xor (layer0_outputs(9646));
    outputs(1870) <= (layer0_outputs(8165)) and (layer0_outputs(2518));
    outputs(1871) <= layer0_outputs(2604);
    outputs(1872) <= not(layer0_outputs(9423));
    outputs(1873) <= not((layer0_outputs(3237)) or (layer0_outputs(10483)));
    outputs(1874) <= layer0_outputs(8136);
    outputs(1875) <= (layer0_outputs(2358)) xor (layer0_outputs(3523));
    outputs(1876) <= (layer0_outputs(2964)) and not (layer0_outputs(5375));
    outputs(1877) <= (layer0_outputs(4373)) and not (layer0_outputs(789));
    outputs(1878) <= (layer0_outputs(1473)) and not (layer0_outputs(8333));
    outputs(1879) <= (layer0_outputs(9202)) xor (layer0_outputs(3607));
    outputs(1880) <= not((layer0_outputs(11442)) xor (layer0_outputs(8210)));
    outputs(1881) <= layer0_outputs(10864);
    outputs(1882) <= (layer0_outputs(5324)) and not (layer0_outputs(6982));
    outputs(1883) <= (layer0_outputs(3455)) and (layer0_outputs(4492));
    outputs(1884) <= (layer0_outputs(2978)) xor (layer0_outputs(2408));
    outputs(1885) <= (layer0_outputs(6186)) and not (layer0_outputs(12386));
    outputs(1886) <= (layer0_outputs(4217)) and (layer0_outputs(11964));
    outputs(1887) <= (layer0_outputs(881)) and not (layer0_outputs(4166));
    outputs(1888) <= (layer0_outputs(11248)) xor (layer0_outputs(10017));
    outputs(1889) <= not(layer0_outputs(8614));
    outputs(1890) <= not(layer0_outputs(5891));
    outputs(1891) <= layer0_outputs(8434);
    outputs(1892) <= (layer0_outputs(4732)) xor (layer0_outputs(11540));
    outputs(1893) <= (layer0_outputs(11638)) and not (layer0_outputs(5146));
    outputs(1894) <= (layer0_outputs(3948)) xor (layer0_outputs(7040));
    outputs(1895) <= not((layer0_outputs(10645)) or (layer0_outputs(5294)));
    outputs(1896) <= (layer0_outputs(1787)) and not (layer0_outputs(6027));
    outputs(1897) <= (layer0_outputs(7550)) and not (layer0_outputs(12276));
    outputs(1898) <= (layer0_outputs(7236)) xor (layer0_outputs(10050));
    outputs(1899) <= (layer0_outputs(7908)) and not (layer0_outputs(9322));
    outputs(1900) <= layer0_outputs(3316);
    outputs(1901) <= layer0_outputs(4240);
    outputs(1902) <= layer0_outputs(8286);
    outputs(1903) <= (layer0_outputs(402)) and (layer0_outputs(8537));
    outputs(1904) <= (layer0_outputs(3653)) xor (layer0_outputs(178));
    outputs(1905) <= layer0_outputs(7858);
    outputs(1906) <= not((layer0_outputs(1685)) xor (layer0_outputs(10533)));
    outputs(1907) <= (layer0_outputs(9510)) and not (layer0_outputs(8125));
    outputs(1908) <= layer0_outputs(6740);
    outputs(1909) <= not((layer0_outputs(9696)) xor (layer0_outputs(6998)));
    outputs(1910) <= layer0_outputs(8312);
    outputs(1911) <= layer0_outputs(1107);
    outputs(1912) <= not((layer0_outputs(11718)) or (layer0_outputs(1536)));
    outputs(1913) <= (layer0_outputs(5783)) and not (layer0_outputs(2519));
    outputs(1914) <= layer0_outputs(4571);
    outputs(1915) <= layer0_outputs(1046);
    outputs(1916) <= not((layer0_outputs(10508)) xor (layer0_outputs(6625)));
    outputs(1917) <= not((layer0_outputs(2854)) xor (layer0_outputs(2551)));
    outputs(1918) <= (layer0_outputs(10822)) and (layer0_outputs(8034));
    outputs(1919) <= (layer0_outputs(2623)) and not (layer0_outputs(6350));
    outputs(1920) <= (layer0_outputs(1149)) and (layer0_outputs(5338));
    outputs(1921) <= (layer0_outputs(354)) and (layer0_outputs(9284));
    outputs(1922) <= not((layer0_outputs(2921)) xor (layer0_outputs(1710)));
    outputs(1923) <= not((layer0_outputs(5607)) xor (layer0_outputs(2036)));
    outputs(1924) <= layer0_outputs(1517);
    outputs(1925) <= not((layer0_outputs(11673)) or (layer0_outputs(510)));
    outputs(1926) <= (layer0_outputs(9008)) and not (layer0_outputs(4682));
    outputs(1927) <= (layer0_outputs(7435)) and not (layer0_outputs(8448));
    outputs(1928) <= (layer0_outputs(3389)) and (layer0_outputs(1531));
    outputs(1929) <= layer0_outputs(6995);
    outputs(1930) <= not((layer0_outputs(11846)) or (layer0_outputs(10348)));
    outputs(1931) <= not((layer0_outputs(8981)) or (layer0_outputs(9705)));
    outputs(1932) <= not((layer0_outputs(11631)) or (layer0_outputs(819)));
    outputs(1933) <= layer0_outputs(3946);
    outputs(1934) <= (layer0_outputs(6236)) and (layer0_outputs(9914));
    outputs(1935) <= (layer0_outputs(7915)) and (layer0_outputs(5948));
    outputs(1936) <= not((layer0_outputs(11091)) xor (layer0_outputs(5671)));
    outputs(1937) <= (layer0_outputs(10047)) and (layer0_outputs(5098));
    outputs(1938) <= not((layer0_outputs(4832)) or (layer0_outputs(5160)));
    outputs(1939) <= (layer0_outputs(2861)) and not (layer0_outputs(8417));
    outputs(1940) <= (layer0_outputs(858)) xor (layer0_outputs(3345));
    outputs(1941) <= (layer0_outputs(3015)) and (layer0_outputs(3494));
    outputs(1942) <= (layer0_outputs(7104)) xor (layer0_outputs(6738));
    outputs(1943) <= (layer0_outputs(11320)) and not (layer0_outputs(9254));
    outputs(1944) <= (layer0_outputs(10886)) and not (layer0_outputs(11746));
    outputs(1945) <= (layer0_outputs(9819)) and not (layer0_outputs(1913));
    outputs(1946) <= not((layer0_outputs(8367)) xor (layer0_outputs(7255)));
    outputs(1947) <= (layer0_outputs(716)) and not (layer0_outputs(10911));
    outputs(1948) <= (layer0_outputs(1844)) and not (layer0_outputs(1952));
    outputs(1949) <= layer0_outputs(2430);
    outputs(1950) <= (layer0_outputs(12003)) and not (layer0_outputs(1882));
    outputs(1951) <= (layer0_outputs(12671)) xor (layer0_outputs(1995));
    outputs(1952) <= (layer0_outputs(6955)) and not (layer0_outputs(5508));
    outputs(1953) <= not((layer0_outputs(3508)) xor (layer0_outputs(4823)));
    outputs(1954) <= not(layer0_outputs(468));
    outputs(1955) <= (layer0_outputs(11240)) xor (layer0_outputs(10410));
    outputs(1956) <= not((layer0_outputs(9816)) xor (layer0_outputs(10241)));
    outputs(1957) <= layer0_outputs(3045);
    outputs(1958) <= not((layer0_outputs(778)) or (layer0_outputs(7045)));
    outputs(1959) <= not(layer0_outputs(4999));
    outputs(1960) <= not((layer0_outputs(6362)) or (layer0_outputs(2526)));
    outputs(1961) <= layer0_outputs(6443);
    outputs(1962) <= not((layer0_outputs(1047)) or (layer0_outputs(1078)));
    outputs(1963) <= not((layer0_outputs(7110)) xor (layer0_outputs(6292)));
    outputs(1964) <= not((layer0_outputs(7851)) or (layer0_outputs(3257)));
    outputs(1965) <= not(layer0_outputs(7750));
    outputs(1966) <= (layer0_outputs(10460)) and (layer0_outputs(5628));
    outputs(1967) <= (layer0_outputs(2875)) and not (layer0_outputs(1754));
    outputs(1968) <= not((layer0_outputs(1285)) xor (layer0_outputs(2430)));
    outputs(1969) <= layer0_outputs(9297);
    outputs(1970) <= (layer0_outputs(12060)) and not (layer0_outputs(8826));
    outputs(1971) <= layer0_outputs(10522);
    outputs(1972) <= not((layer0_outputs(12707)) or (layer0_outputs(12031)));
    outputs(1973) <= layer0_outputs(11776);
    outputs(1974) <= not((layer0_outputs(11959)) xor (layer0_outputs(8304)));
    outputs(1975) <= not(layer0_outputs(7728));
    outputs(1976) <= not(layer0_outputs(8378));
    outputs(1977) <= layer0_outputs(9289);
    outputs(1978) <= not(layer0_outputs(10282));
    outputs(1979) <= not(layer0_outputs(6869));
    outputs(1980) <= layer0_outputs(6312);
    outputs(1981) <= not((layer0_outputs(6155)) xor (layer0_outputs(2571)));
    outputs(1982) <= not((layer0_outputs(12224)) xor (layer0_outputs(2158)));
    outputs(1983) <= (layer0_outputs(10335)) and not (layer0_outputs(6237));
    outputs(1984) <= not((layer0_outputs(11449)) or (layer0_outputs(6599)));
    outputs(1985) <= not((layer0_outputs(7229)) xor (layer0_outputs(775)));
    outputs(1986) <= not((layer0_outputs(4208)) or (layer0_outputs(6931)));
    outputs(1987) <= not(layer0_outputs(8912));
    outputs(1988) <= not(layer0_outputs(6865));
    outputs(1989) <= (layer0_outputs(8696)) and not (layer0_outputs(2468));
    outputs(1990) <= not(layer0_outputs(7795));
    outputs(1991) <= not(layer0_outputs(950));
    outputs(1992) <= not(layer0_outputs(11697));
    outputs(1993) <= not((layer0_outputs(11760)) or (layer0_outputs(12677)));
    outputs(1994) <= not(layer0_outputs(7495));
    outputs(1995) <= not(layer0_outputs(6805));
    outputs(1996) <= not((layer0_outputs(3040)) xor (layer0_outputs(3978)));
    outputs(1997) <= layer0_outputs(12155);
    outputs(1998) <= (layer0_outputs(8554)) xor (layer0_outputs(1108));
    outputs(1999) <= not(layer0_outputs(4110));
    outputs(2000) <= '0';
    outputs(2001) <= (layer0_outputs(1870)) and not (layer0_outputs(8593));
    outputs(2002) <= not((layer0_outputs(4422)) or (layer0_outputs(11143)));
    outputs(2003) <= (layer0_outputs(2046)) and not (layer0_outputs(8955));
    outputs(2004) <= (layer0_outputs(574)) and not (layer0_outputs(7289));
    outputs(2005) <= (layer0_outputs(900)) and not (layer0_outputs(9391));
    outputs(2006) <= not((layer0_outputs(9022)) xor (layer0_outputs(564)));
    outputs(2007) <= not(layer0_outputs(6364));
    outputs(2008) <= not((layer0_outputs(4353)) xor (layer0_outputs(2402)));
    outputs(2009) <= (layer0_outputs(83)) and not (layer0_outputs(4226));
    outputs(2010) <= not((layer0_outputs(12373)) or (layer0_outputs(10971)));
    outputs(2011) <= (layer0_outputs(811)) xor (layer0_outputs(6411));
    outputs(2012) <= layer0_outputs(3428);
    outputs(2013) <= (layer0_outputs(4454)) and not (layer0_outputs(4996));
    outputs(2014) <= (layer0_outputs(9932)) and not (layer0_outputs(3157));
    outputs(2015) <= not((layer0_outputs(432)) xor (layer0_outputs(12033)));
    outputs(2016) <= not(layer0_outputs(7988));
    outputs(2017) <= not((layer0_outputs(10213)) or (layer0_outputs(7862)));
    outputs(2018) <= not((layer0_outputs(3705)) xor (layer0_outputs(12619)));
    outputs(2019) <= (layer0_outputs(12158)) and not (layer0_outputs(3850));
    outputs(2020) <= (layer0_outputs(9945)) and not (layer0_outputs(12216));
    outputs(2021) <= '0';
    outputs(2022) <= (layer0_outputs(2911)) xor (layer0_outputs(6182));
    outputs(2023) <= not((layer0_outputs(11622)) xor (layer0_outputs(11239)));
    outputs(2024) <= not(layer0_outputs(3657));
    outputs(2025) <= not((layer0_outputs(2739)) or (layer0_outputs(11536)));
    outputs(2026) <= (layer0_outputs(6041)) and not (layer0_outputs(1747));
    outputs(2027) <= (layer0_outputs(3042)) and not (layer0_outputs(8065));
    outputs(2028) <= not((layer0_outputs(3136)) xor (layer0_outputs(12007)));
    outputs(2029) <= (layer0_outputs(11724)) xor (layer0_outputs(1316));
    outputs(2030) <= (layer0_outputs(2943)) xor (layer0_outputs(4098));
    outputs(2031) <= (layer0_outputs(10456)) and not (layer0_outputs(5420));
    outputs(2032) <= not(layer0_outputs(9127));
    outputs(2033) <= not((layer0_outputs(1720)) xor (layer0_outputs(11702)));
    outputs(2034) <= layer0_outputs(12653);
    outputs(2035) <= (layer0_outputs(8769)) and (layer0_outputs(3303));
    outputs(2036) <= not((layer0_outputs(1351)) xor (layer0_outputs(4432)));
    outputs(2037) <= (layer0_outputs(12444)) and not (layer0_outputs(8279));
    outputs(2038) <= '0';
    outputs(2039) <= (layer0_outputs(5207)) xor (layer0_outputs(1806));
    outputs(2040) <= layer0_outputs(7257);
    outputs(2041) <= not((layer0_outputs(4408)) xor (layer0_outputs(11019)));
    outputs(2042) <= layer0_outputs(672);
    outputs(2043) <= (layer0_outputs(3789)) and (layer0_outputs(5016));
    outputs(2044) <= not((layer0_outputs(6514)) or (layer0_outputs(8493)));
    outputs(2045) <= (layer0_outputs(6181)) and not (layer0_outputs(4810));
    outputs(2046) <= layer0_outputs(10022);
    outputs(2047) <= (layer0_outputs(7195)) and not (layer0_outputs(5794));
    outputs(2048) <= (layer0_outputs(7605)) and not (layer0_outputs(9384));
    outputs(2049) <= not(layer0_outputs(6347));
    outputs(2050) <= layer0_outputs(3562);
    outputs(2051) <= (layer0_outputs(5510)) and not (layer0_outputs(9415));
    outputs(2052) <= layer0_outputs(299);
    outputs(2053) <= not(layer0_outputs(668));
    outputs(2054) <= (layer0_outputs(9614)) and not (layer0_outputs(10551));
    outputs(2055) <= '0';
    outputs(2056) <= (layer0_outputs(3058)) xor (layer0_outputs(12113));
    outputs(2057) <= (layer0_outputs(11221)) xor (layer0_outputs(7510));
    outputs(2058) <= not((layer0_outputs(12409)) or (layer0_outputs(6699)));
    outputs(2059) <= (layer0_outputs(7366)) and not (layer0_outputs(6165));
    outputs(2060) <= not(layer0_outputs(4231));
    outputs(2061) <= (layer0_outputs(4603)) xor (layer0_outputs(11491));
    outputs(2062) <= not(layer0_outputs(4387));
    outputs(2063) <= '0';
    outputs(2064) <= not((layer0_outputs(10217)) or (layer0_outputs(4824)));
    outputs(2065) <= (layer0_outputs(882)) and not (layer0_outputs(11684));
    outputs(2066) <= not(layer0_outputs(4448));
    outputs(2067) <= layer0_outputs(12139);
    outputs(2068) <= not((layer0_outputs(3044)) xor (layer0_outputs(3055)));
    outputs(2069) <= (layer0_outputs(10426)) and (layer0_outputs(1722));
    outputs(2070) <= not((layer0_outputs(1424)) xor (layer0_outputs(12218)));
    outputs(2071) <= (layer0_outputs(8913)) and (layer0_outputs(6350));
    outputs(2072) <= (layer0_outputs(5953)) and (layer0_outputs(6877));
    outputs(2073) <= (layer0_outputs(12618)) and not (layer0_outputs(2250));
    outputs(2074) <= not(layer0_outputs(6393));
    outputs(2075) <= (layer0_outputs(10818)) and (layer0_outputs(11816));
    outputs(2076) <= (layer0_outputs(2276)) and not (layer0_outputs(3876));
    outputs(2077) <= (layer0_outputs(11192)) xor (layer0_outputs(2066));
    outputs(2078) <= (layer0_outputs(11570)) and not (layer0_outputs(4677));
    outputs(2079) <= layer0_outputs(188);
    outputs(2080) <= (layer0_outputs(12387)) and not (layer0_outputs(12535));
    outputs(2081) <= layer0_outputs(7336);
    outputs(2082) <= layer0_outputs(7322);
    outputs(2083) <= (layer0_outputs(8635)) and (layer0_outputs(3758));
    outputs(2084) <= not(layer0_outputs(8073));
    outputs(2085) <= (layer0_outputs(11436)) and not (layer0_outputs(9355));
    outputs(2086) <= (layer0_outputs(580)) and not (layer0_outputs(7496));
    outputs(2087) <= (layer0_outputs(12472)) and not (layer0_outputs(4443));
    outputs(2088) <= not(layer0_outputs(5769));
    outputs(2089) <= not((layer0_outputs(12385)) or (layer0_outputs(9301)));
    outputs(2090) <= (layer0_outputs(1102)) and not (layer0_outputs(6101));
    outputs(2091) <= (layer0_outputs(1558)) xor (layer0_outputs(4149));
    outputs(2092) <= (layer0_outputs(9294)) xor (layer0_outputs(1905));
    outputs(2093) <= not((layer0_outputs(9331)) xor (layer0_outputs(8161)));
    outputs(2094) <= not((layer0_outputs(5313)) xor (layer0_outputs(9432)));
    outputs(2095) <= (layer0_outputs(1103)) and not (layer0_outputs(635));
    outputs(2096) <= not((layer0_outputs(8006)) xor (layer0_outputs(3155)));
    outputs(2097) <= (layer0_outputs(4914)) and not (layer0_outputs(7889));
    outputs(2098) <= (layer0_outputs(6357)) xor (layer0_outputs(12642));
    outputs(2099) <= not(layer0_outputs(988));
    outputs(2100) <= layer0_outputs(8326);
    outputs(2101) <= not((layer0_outputs(10433)) xor (layer0_outputs(1366)));
    outputs(2102) <= not((layer0_outputs(842)) xor (layer0_outputs(8736)));
    outputs(2103) <= (layer0_outputs(2137)) and not (layer0_outputs(5281));
    outputs(2104) <= not((layer0_outputs(570)) or (layer0_outputs(12696)));
    outputs(2105) <= '0';
    outputs(2106) <= (layer0_outputs(4701)) and not (layer0_outputs(4453));
    outputs(2107) <= (layer0_outputs(5557)) xor (layer0_outputs(6544));
    outputs(2108) <= (layer0_outputs(6250)) xor (layer0_outputs(3827));
    outputs(2109) <= '0';
    outputs(2110) <= not((layer0_outputs(3128)) and (layer0_outputs(12157)));
    outputs(2111) <= (layer0_outputs(1001)) and (layer0_outputs(6579));
    outputs(2112) <= (layer0_outputs(4745)) xor (layer0_outputs(1361));
    outputs(2113) <= not((layer0_outputs(8910)) or (layer0_outputs(3400)));
    outputs(2114) <= not(layer0_outputs(12299));
    outputs(2115) <= not((layer0_outputs(4553)) xor (layer0_outputs(3331)));
    outputs(2116) <= layer0_outputs(3567);
    outputs(2117) <= layer0_outputs(10966);
    outputs(2118) <= not((layer0_outputs(4125)) or (layer0_outputs(12131)));
    outputs(2119) <= not((layer0_outputs(9260)) xor (layer0_outputs(3885)));
    outputs(2120) <= not(layer0_outputs(6554));
    outputs(2121) <= not((layer0_outputs(6742)) or (layer0_outputs(215)));
    outputs(2122) <= not(layer0_outputs(3319));
    outputs(2123) <= (layer0_outputs(7394)) and (layer0_outputs(9619));
    outputs(2124) <= (layer0_outputs(4249)) or (layer0_outputs(3258));
    outputs(2125) <= (layer0_outputs(3873)) xor (layer0_outputs(11280));
    outputs(2126) <= (layer0_outputs(2578)) and not (layer0_outputs(2528));
    outputs(2127) <= (layer0_outputs(4676)) and (layer0_outputs(8257));
    outputs(2128) <= (layer0_outputs(1943)) and not (layer0_outputs(3337));
    outputs(2129) <= not((layer0_outputs(3869)) and (layer0_outputs(5429)));
    outputs(2130) <= (layer0_outputs(11382)) and (layer0_outputs(3907));
    outputs(2131) <= not(layer0_outputs(1404));
    outputs(2132) <= (layer0_outputs(6169)) xor (layer0_outputs(12021));
    outputs(2133) <= not((layer0_outputs(12736)) or (layer0_outputs(8850)));
    outputs(2134) <= (layer0_outputs(3804)) and (layer0_outputs(85));
    outputs(2135) <= layer0_outputs(11237);
    outputs(2136) <= (layer0_outputs(10045)) and (layer0_outputs(3355));
    outputs(2137) <= not((layer0_outputs(6719)) xor (layer0_outputs(3521)));
    outputs(2138) <= layer0_outputs(11483);
    outputs(2139) <= not(layer0_outputs(8547));
    outputs(2140) <= not((layer0_outputs(6413)) xor (layer0_outputs(9321)));
    outputs(2141) <= (layer0_outputs(10914)) and not (layer0_outputs(4269));
    outputs(2142) <= layer0_outputs(8011);
    outputs(2143) <= not(layer0_outputs(10366));
    outputs(2144) <= (layer0_outputs(11388)) and not (layer0_outputs(6325));
    outputs(2145) <= not(layer0_outputs(8392));
    outputs(2146) <= (layer0_outputs(11721)) and not (layer0_outputs(6706));
    outputs(2147) <= (layer0_outputs(7601)) and not (layer0_outputs(12128));
    outputs(2148) <= not((layer0_outputs(7824)) and (layer0_outputs(1165)));
    outputs(2149) <= (layer0_outputs(6185)) and (layer0_outputs(3412));
    outputs(2150) <= layer0_outputs(4769);
    outputs(2151) <= not((layer0_outputs(1712)) or (layer0_outputs(5166)));
    outputs(2152) <= layer0_outputs(10694);
    outputs(2153) <= not((layer0_outputs(11652)) xor (layer0_outputs(1505)));
    outputs(2154) <= (layer0_outputs(8650)) and not (layer0_outputs(7566));
    outputs(2155) <= not((layer0_outputs(2850)) xor (layer0_outputs(11549)));
    outputs(2156) <= layer0_outputs(5548);
    outputs(2157) <= layer0_outputs(2431);
    outputs(2158) <= (layer0_outputs(12162)) xor (layer0_outputs(309));
    outputs(2159) <= not((layer0_outputs(12795)) or (layer0_outputs(11758)));
    outputs(2160) <= (layer0_outputs(7620)) and not (layer0_outputs(2746));
    outputs(2161) <= '0';
    outputs(2162) <= layer0_outputs(11493);
    outputs(2163) <= not(layer0_outputs(11256));
    outputs(2164) <= not((layer0_outputs(7617)) xor (layer0_outputs(8424)));
    outputs(2165) <= not(layer0_outputs(6265));
    outputs(2166) <= not(layer0_outputs(3800));
    outputs(2167) <= (layer0_outputs(4780)) and not (layer0_outputs(7237));
    outputs(2168) <= not(layer0_outputs(9473));
    outputs(2169) <= not(layer0_outputs(6292));
    outputs(2170) <= layer0_outputs(10712);
    outputs(2171) <= layer0_outputs(9620);
    outputs(2172) <= (layer0_outputs(2190)) xor (layer0_outputs(5927));
    outputs(2173) <= not((layer0_outputs(1212)) xor (layer0_outputs(3565)));
    outputs(2174) <= (layer0_outputs(5455)) xor (layer0_outputs(10934));
    outputs(2175) <= layer0_outputs(12344);
    outputs(2176) <= (layer0_outputs(5960)) xor (layer0_outputs(11807));
    outputs(2177) <= (layer0_outputs(10065)) and (layer0_outputs(11479));
    outputs(2178) <= layer0_outputs(2959);
    outputs(2179) <= (layer0_outputs(2955)) xor (layer0_outputs(6180));
    outputs(2180) <= '0';
    outputs(2181) <= (layer0_outputs(6647)) and not (layer0_outputs(7151));
    outputs(2182) <= not((layer0_outputs(8117)) xor (layer0_outputs(9173)));
    outputs(2183) <= (layer0_outputs(456)) and not (layer0_outputs(8418));
    outputs(2184) <= layer0_outputs(10935);
    outputs(2185) <= (layer0_outputs(2088)) and not (layer0_outputs(6555));
    outputs(2186) <= not((layer0_outputs(12692)) or (layer0_outputs(5086)));
    outputs(2187) <= layer0_outputs(8836);
    outputs(2188) <= (layer0_outputs(5428)) and (layer0_outputs(1846));
    outputs(2189) <= (layer0_outputs(3281)) and (layer0_outputs(1312));
    outputs(2190) <= (layer0_outputs(4503)) and (layer0_outputs(3867));
    outputs(2191) <= layer0_outputs(10306);
    outputs(2192) <= (layer0_outputs(11907)) and not (layer0_outputs(8071));
    outputs(2193) <= layer0_outputs(8185);
    outputs(2194) <= (layer0_outputs(4713)) and not (layer0_outputs(5890));
    outputs(2195) <= not((layer0_outputs(4024)) or (layer0_outputs(2953)));
    outputs(2196) <= not((layer0_outputs(11137)) xor (layer0_outputs(4365)));
    outputs(2197) <= (layer0_outputs(7165)) and not (layer0_outputs(12386));
    outputs(2198) <= not((layer0_outputs(1293)) xor (layer0_outputs(12541)));
    outputs(2199) <= not(layer0_outputs(5468));
    outputs(2200) <= (layer0_outputs(12370)) and (layer0_outputs(5758));
    outputs(2201) <= (layer0_outputs(6641)) and (layer0_outputs(12470));
    outputs(2202) <= (layer0_outputs(11705)) and not (layer0_outputs(10625));
    outputs(2203) <= not(layer0_outputs(721));
    outputs(2204) <= layer0_outputs(10166);
    outputs(2205) <= (layer0_outputs(6419)) and not (layer0_outputs(6891));
    outputs(2206) <= not((layer0_outputs(5144)) or (layer0_outputs(1927)));
    outputs(2207) <= (layer0_outputs(9583)) and not (layer0_outputs(938));
    outputs(2208) <= not((layer0_outputs(12027)) xor (layer0_outputs(683)));
    outputs(2209) <= layer0_outputs(2449);
    outputs(2210) <= not(layer0_outputs(4421));
    outputs(2211) <= (layer0_outputs(10194)) xor (layer0_outputs(3456));
    outputs(2212) <= (layer0_outputs(12175)) and not (layer0_outputs(3121));
    outputs(2213) <= not((layer0_outputs(12096)) or (layer0_outputs(7877)));
    outputs(2214) <= not((layer0_outputs(6333)) or (layer0_outputs(535)));
    outputs(2215) <= layer0_outputs(7209);
    outputs(2216) <= not(layer0_outputs(3931));
    outputs(2217) <= (layer0_outputs(3145)) and not (layer0_outputs(5936));
    outputs(2218) <= (layer0_outputs(10258)) and not (layer0_outputs(747));
    outputs(2219) <= (layer0_outputs(6051)) and not (layer0_outputs(10813));
    outputs(2220) <= not(layer0_outputs(6139));
    outputs(2221) <= (layer0_outputs(9)) and not (layer0_outputs(12424));
    outputs(2222) <= '0';
    outputs(2223) <= not(layer0_outputs(3198));
    outputs(2224) <= not((layer0_outputs(9373)) xor (layer0_outputs(962)));
    outputs(2225) <= (layer0_outputs(2776)) and (layer0_outputs(3683));
    outputs(2226) <= not((layer0_outputs(4045)) or (layer0_outputs(9399)));
    outputs(2227) <= (layer0_outputs(3445)) and (layer0_outputs(3536));
    outputs(2228) <= not((layer0_outputs(1148)) or (layer0_outputs(10922)));
    outputs(2229) <= not(layer0_outputs(5576));
    outputs(2230) <= (layer0_outputs(10729)) xor (layer0_outputs(3048));
    outputs(2231) <= (layer0_outputs(5762)) and (layer0_outputs(1421));
    outputs(2232) <= (layer0_outputs(3710)) xor (layer0_outputs(6493));
    outputs(2233) <= (layer0_outputs(11217)) and (layer0_outputs(9731));
    outputs(2234) <= (layer0_outputs(4649)) xor (layer0_outputs(3602));
    outputs(2235) <= not((layer0_outputs(270)) xor (layer0_outputs(7458)));
    outputs(2236) <= (layer0_outputs(11161)) and not (layer0_outputs(4955));
    outputs(2237) <= (layer0_outputs(1087)) xor (layer0_outputs(6308));
    outputs(2238) <= not((layer0_outputs(6648)) xor (layer0_outputs(4088)));
    outputs(2239) <= not((layer0_outputs(6228)) xor (layer0_outputs(1568)));
    outputs(2240) <= layer0_outputs(9497);
    outputs(2241) <= (layer0_outputs(10447)) and (layer0_outputs(7804));
    outputs(2242) <= not((layer0_outputs(124)) or (layer0_outputs(4452)));
    outputs(2243) <= not((layer0_outputs(4932)) xor (layer0_outputs(3069)));
    outputs(2244) <= (layer0_outputs(9147)) and not (layer0_outputs(12389));
    outputs(2245) <= layer0_outputs(6954);
    outputs(2246) <= not(layer0_outputs(11699));
    outputs(2247) <= not(layer0_outputs(3395)) or (layer0_outputs(216));
    outputs(2248) <= layer0_outputs(518);
    outputs(2249) <= not((layer0_outputs(7784)) xor (layer0_outputs(7240)));
    outputs(2250) <= (layer0_outputs(3365)) and not (layer0_outputs(7950));
    outputs(2251) <= (layer0_outputs(4137)) and not (layer0_outputs(9342));
    outputs(2252) <= (layer0_outputs(6199)) and not (layer0_outputs(2201));
    outputs(2253) <= (layer0_outputs(10882)) and not (layer0_outputs(3570));
    outputs(2254) <= not(layer0_outputs(5244));
    outputs(2255) <= not((layer0_outputs(7466)) or (layer0_outputs(12395)));
    outputs(2256) <= not(layer0_outputs(6778));
    outputs(2257) <= not(layer0_outputs(3980));
    outputs(2258) <= not((layer0_outputs(6799)) xor (layer0_outputs(2231)));
    outputs(2259) <= not(layer0_outputs(1625));
    outputs(2260) <= not(layer0_outputs(7384));
    outputs(2261) <= layer0_outputs(4427);
    outputs(2262) <= not((layer0_outputs(2544)) or (layer0_outputs(7316)));
    outputs(2263) <= not((layer0_outputs(6097)) xor (layer0_outputs(1683)));
    outputs(2264) <= (layer0_outputs(915)) and not (layer0_outputs(1290));
    outputs(2265) <= (layer0_outputs(8372)) and not (layer0_outputs(4506));
    outputs(2266) <= not(layer0_outputs(1210));
    outputs(2267) <= (layer0_outputs(12559)) and not (layer0_outputs(2254));
    outputs(2268) <= (layer0_outputs(11405)) xor (layer0_outputs(10652));
    outputs(2269) <= (layer0_outputs(5063)) and (layer0_outputs(526));
    outputs(2270) <= not(layer0_outputs(11204));
    outputs(2271) <= (layer0_outputs(3160)) and (layer0_outputs(261));
    outputs(2272) <= not((layer0_outputs(7573)) xor (layer0_outputs(2575)));
    outputs(2273) <= layer0_outputs(1138);
    outputs(2274) <= '0';
    outputs(2275) <= not(layer0_outputs(11862));
    outputs(2276) <= (layer0_outputs(10681)) and not (layer0_outputs(8583));
    outputs(2277) <= (layer0_outputs(12683)) and not (layer0_outputs(165));
    outputs(2278) <= not(layer0_outputs(2991));
    outputs(2279) <= (layer0_outputs(10266)) xor (layer0_outputs(5307));
    outputs(2280) <= not((layer0_outputs(5707)) xor (layer0_outputs(5100)));
    outputs(2281) <= (layer0_outputs(132)) and not (layer0_outputs(3847));
    outputs(2282) <= (layer0_outputs(11048)) and (layer0_outputs(1593));
    outputs(2283) <= (layer0_outputs(1885)) and (layer0_outputs(7876));
    outputs(2284) <= (layer0_outputs(5854)) xor (layer0_outputs(7674));
    outputs(2285) <= (layer0_outputs(2635)) and not (layer0_outputs(4110));
    outputs(2286) <= not(layer0_outputs(6530));
    outputs(2287) <= (layer0_outputs(10970)) xor (layer0_outputs(6483));
    outputs(2288) <= not((layer0_outputs(11520)) xor (layer0_outputs(12519)));
    outputs(2289) <= (layer0_outputs(764)) and (layer0_outputs(10735));
    outputs(2290) <= (layer0_outputs(5752)) xor (layer0_outputs(7980));
    outputs(2291) <= (layer0_outputs(12557)) and not (layer0_outputs(6371));
    outputs(2292) <= (layer0_outputs(8883)) xor (layer0_outputs(9012));
    outputs(2293) <= (layer0_outputs(6721)) xor (layer0_outputs(11351));
    outputs(2294) <= layer0_outputs(2907);
    outputs(2295) <= (layer0_outputs(10999)) and not (layer0_outputs(8701));
    outputs(2296) <= (layer0_outputs(6131)) and not (layer0_outputs(4540));
    outputs(2297) <= (layer0_outputs(3774)) xor (layer0_outputs(5014));
    outputs(2298) <= not(layer0_outputs(1040));
    outputs(2299) <= (layer0_outputs(9808)) and (layer0_outputs(3348));
    outputs(2300) <= not(layer0_outputs(5592));
    outputs(2301) <= not(layer0_outputs(230));
    outputs(2302) <= (layer0_outputs(467)) or (layer0_outputs(8116));
    outputs(2303) <= layer0_outputs(8737);
    outputs(2304) <= not(layer0_outputs(4155));
    outputs(2305) <= (layer0_outputs(11325)) and (layer0_outputs(7435));
    outputs(2306) <= (layer0_outputs(4564)) and not (layer0_outputs(637));
    outputs(2307) <= (layer0_outputs(910)) xor (layer0_outputs(391));
    outputs(2308) <= (layer0_outputs(2072)) xor (layer0_outputs(11363));
    outputs(2309) <= not(layer0_outputs(4191));
    outputs(2310) <= (layer0_outputs(8371)) and (layer0_outputs(10309));
    outputs(2311) <= (layer0_outputs(8258)) and not (layer0_outputs(3367));
    outputs(2312) <= layer0_outputs(5554);
    outputs(2313) <= not(layer0_outputs(576));
    outputs(2314) <= not((layer0_outputs(7729)) or (layer0_outputs(12035)));
    outputs(2315) <= (layer0_outputs(8576)) xor (layer0_outputs(2576));
    outputs(2316) <= (layer0_outputs(7684)) and (layer0_outputs(10300));
    outputs(2317) <= not((layer0_outputs(384)) xor (layer0_outputs(6650)));
    outputs(2318) <= (layer0_outputs(3761)) and not (layer0_outputs(6422));
    outputs(2319) <= (layer0_outputs(4646)) xor (layer0_outputs(12333));
    outputs(2320) <= (layer0_outputs(3943)) and (layer0_outputs(2061));
    outputs(2321) <= (layer0_outputs(3454)) and not (layer0_outputs(1289));
    outputs(2322) <= (layer0_outputs(8522)) and not (layer0_outputs(6672));
    outputs(2323) <= (layer0_outputs(10245)) and not (layer0_outputs(546));
    outputs(2324) <= not((layer0_outputs(11758)) or (layer0_outputs(8099)));
    outputs(2325) <= (layer0_outputs(1925)) or (layer0_outputs(10818));
    outputs(2326) <= (layer0_outputs(486)) and not (layer0_outputs(9166));
    outputs(2327) <= not((layer0_outputs(7010)) xor (layer0_outputs(9818)));
    outputs(2328) <= (layer0_outputs(3396)) xor (layer0_outputs(2762));
    outputs(2329) <= '0';
    outputs(2330) <= not((layer0_outputs(1430)) xor (layer0_outputs(8834)));
    outputs(2331) <= (layer0_outputs(7763)) and not (layer0_outputs(5624));
    outputs(2332) <= (layer0_outputs(11221)) and not (layer0_outputs(5652));
    outputs(2333) <= (layer0_outputs(7239)) and (layer0_outputs(9908));
    outputs(2334) <= (layer0_outputs(8552)) and not (layer0_outputs(8657));
    outputs(2335) <= (layer0_outputs(2980)) and not (layer0_outputs(1736));
    outputs(2336) <= not(layer0_outputs(4247));
    outputs(2337) <= not(layer0_outputs(12753)) or (layer0_outputs(4168));
    outputs(2338) <= not((layer0_outputs(2027)) xor (layer0_outputs(8824)));
    outputs(2339) <= not(layer0_outputs(1083));
    outputs(2340) <= layer0_outputs(4516);
    outputs(2341) <= (layer0_outputs(12387)) xor (layer0_outputs(9832));
    outputs(2342) <= (layer0_outputs(2399)) and (layer0_outputs(7835));
    outputs(2343) <= (layer0_outputs(4738)) and not (layer0_outputs(3114));
    outputs(2344) <= (layer0_outputs(12047)) xor (layer0_outputs(642));
    outputs(2345) <= not((layer0_outputs(10804)) or (layer0_outputs(1371)));
    outputs(2346) <= (layer0_outputs(4053)) or (layer0_outputs(6849));
    outputs(2347) <= (layer0_outputs(11869)) and (layer0_outputs(9284));
    outputs(2348) <= (layer0_outputs(3919)) xor (layer0_outputs(11242));
    outputs(2349) <= (layer0_outputs(9174)) and not (layer0_outputs(9965));
    outputs(2350) <= (layer0_outputs(8304)) and not (layer0_outputs(219));
    outputs(2351) <= layer0_outputs(9333);
    outputs(2352) <= (layer0_outputs(2786)) and (layer0_outputs(7234));
    outputs(2353) <= not((layer0_outputs(9858)) or (layer0_outputs(12)));
    outputs(2354) <= (layer0_outputs(542)) and not (layer0_outputs(1668));
    outputs(2355) <= not((layer0_outputs(1191)) xor (layer0_outputs(8947)));
    outputs(2356) <= not(layer0_outputs(1581));
    outputs(2357) <= (layer0_outputs(743)) xor (layer0_outputs(6083));
    outputs(2358) <= layer0_outputs(5534);
    outputs(2359) <= not(layer0_outputs(3955)) or (layer0_outputs(885));
    outputs(2360) <= layer0_outputs(3633);
    outputs(2361) <= (layer0_outputs(4392)) and (layer0_outputs(10326));
    outputs(2362) <= not((layer0_outputs(2327)) xor (layer0_outputs(3872)));
    outputs(2363) <= (layer0_outputs(8714)) xor (layer0_outputs(5338));
    outputs(2364) <= (layer0_outputs(7248)) xor (layer0_outputs(9358));
    outputs(2365) <= (layer0_outputs(5935)) xor (layer0_outputs(10588));
    outputs(2366) <= not((layer0_outputs(12045)) or (layer0_outputs(3349)));
    outputs(2367) <= not((layer0_outputs(2235)) xor (layer0_outputs(3608)));
    outputs(2368) <= not((layer0_outputs(4794)) or (layer0_outputs(10459)));
    outputs(2369) <= (layer0_outputs(4565)) xor (layer0_outputs(4457));
    outputs(2370) <= (layer0_outputs(7733)) and not (layer0_outputs(4106));
    outputs(2371) <= (layer0_outputs(7364)) and (layer0_outputs(2873));
    outputs(2372) <= (layer0_outputs(7063)) and not (layer0_outputs(12334));
    outputs(2373) <= '0';
    outputs(2374) <= (layer0_outputs(12680)) and not (layer0_outputs(10665));
    outputs(2375) <= not(layer0_outputs(11385));
    outputs(2376) <= (layer0_outputs(7106)) or (layer0_outputs(4278));
    outputs(2377) <= not((layer0_outputs(6809)) or (layer0_outputs(4087)));
    outputs(2378) <= layer0_outputs(7941);
    outputs(2379) <= not(layer0_outputs(9221));
    outputs(2380) <= (layer0_outputs(4482)) and not (layer0_outputs(11912));
    outputs(2381) <= layer0_outputs(8630);
    outputs(2382) <= not((layer0_outputs(7578)) or (layer0_outputs(8491)));
    outputs(2383) <= layer0_outputs(9513);
    outputs(2384) <= (layer0_outputs(10081)) and not (layer0_outputs(4858));
    outputs(2385) <= not(layer0_outputs(10013));
    outputs(2386) <= not((layer0_outputs(1452)) xor (layer0_outputs(8704)));
    outputs(2387) <= not((layer0_outputs(6243)) or (layer0_outputs(1729)));
    outputs(2388) <= not(layer0_outputs(2476));
    outputs(2389) <= (layer0_outputs(692)) and not (layer0_outputs(6377));
    outputs(2390) <= (layer0_outputs(10628)) and (layer0_outputs(5587));
    outputs(2391) <= not(layer0_outputs(10962));
    outputs(2392) <= (layer0_outputs(7625)) xor (layer0_outputs(2061));
    outputs(2393) <= not((layer0_outputs(9350)) xor (layer0_outputs(4019)));
    outputs(2394) <= layer0_outputs(7806);
    outputs(2395) <= (layer0_outputs(3939)) xor (layer0_outputs(4319));
    outputs(2396) <= (layer0_outputs(10715)) xor (layer0_outputs(5091));
    outputs(2397) <= not(layer0_outputs(10778));
    outputs(2398) <= not((layer0_outputs(10951)) xor (layer0_outputs(8596)));
    outputs(2399) <= not(layer0_outputs(447));
    outputs(2400) <= not(layer0_outputs(1760));
    outputs(2401) <= (layer0_outputs(2043)) and not (layer0_outputs(10962));
    outputs(2402) <= (layer0_outputs(6785)) and not (layer0_outputs(4610));
    outputs(2403) <= not(layer0_outputs(495)) or (layer0_outputs(9151));
    outputs(2404) <= not(layer0_outputs(12390));
    outputs(2405) <= not(layer0_outputs(10478));
    outputs(2406) <= not(layer0_outputs(10127));
    outputs(2407) <= not(layer0_outputs(4455));
    outputs(2408) <= not(layer0_outputs(3614)) or (layer0_outputs(6981));
    outputs(2409) <= not((layer0_outputs(9889)) or (layer0_outputs(9282)));
    outputs(2410) <= not(layer0_outputs(8224));
    outputs(2411) <= not((layer0_outputs(3333)) or (layer0_outputs(12609)));
    outputs(2412) <= layer0_outputs(11889);
    outputs(2413) <= not((layer0_outputs(694)) xor (layer0_outputs(8479)));
    outputs(2414) <= not((layer0_outputs(1077)) or (layer0_outputs(12567)));
    outputs(2415) <= (layer0_outputs(10621)) and not (layer0_outputs(492));
    outputs(2416) <= not(layer0_outputs(11262));
    outputs(2417) <= not((layer0_outputs(2175)) or (layer0_outputs(7067)));
    outputs(2418) <= (layer0_outputs(8749)) and (layer0_outputs(2592));
    outputs(2419) <= not((layer0_outputs(9681)) xor (layer0_outputs(2936)));
    outputs(2420) <= (layer0_outputs(2706)) and not (layer0_outputs(10417));
    outputs(2421) <= layer0_outputs(91);
    outputs(2422) <= not((layer0_outputs(4431)) xor (layer0_outputs(2246)));
    outputs(2423) <= (layer0_outputs(9349)) and (layer0_outputs(3992));
    outputs(2424) <= not((layer0_outputs(2677)) or (layer0_outputs(2595)));
    outputs(2425) <= (layer0_outputs(4755)) xor (layer0_outputs(7167));
    outputs(2426) <= (layer0_outputs(8726)) and (layer0_outputs(2334));
    outputs(2427) <= (layer0_outputs(3372)) and not (layer0_outputs(9412));
    outputs(2428) <= (layer0_outputs(3792)) and (layer0_outputs(1565));
    outputs(2429) <= layer0_outputs(11199);
    outputs(2430) <= (layer0_outputs(12226)) and not (layer0_outputs(5095));
    outputs(2431) <= (layer0_outputs(12788)) and not (layer0_outputs(189));
    outputs(2432) <= not(layer0_outputs(5071));
    outputs(2433) <= (layer0_outputs(5479)) xor (layer0_outputs(5082));
    outputs(2434) <= not(layer0_outputs(2682));
    outputs(2435) <= (layer0_outputs(1373)) xor (layer0_outputs(11016));
    outputs(2436) <= layer0_outputs(5758);
    outputs(2437) <= layer0_outputs(6533);
    outputs(2438) <= (layer0_outputs(1838)) and not (layer0_outputs(1795));
    outputs(2439) <= (layer0_outputs(12222)) xor (layer0_outputs(9371));
    outputs(2440) <= (layer0_outputs(10918)) and not (layer0_outputs(10701));
    outputs(2441) <= not((layer0_outputs(3500)) or (layer0_outputs(44)));
    outputs(2442) <= not((layer0_outputs(6847)) or (layer0_outputs(2485)));
    outputs(2443) <= (layer0_outputs(11585)) and (layer0_outputs(8677));
    outputs(2444) <= not(layer0_outputs(11204));
    outputs(2445) <= (layer0_outputs(3490)) and (layer0_outputs(3127));
    outputs(2446) <= not((layer0_outputs(89)) or (layer0_outputs(9947)));
    outputs(2447) <= (layer0_outputs(6473)) and not (layer0_outputs(989));
    outputs(2448) <= (layer0_outputs(8577)) and (layer0_outputs(9945));
    outputs(2449) <= (layer0_outputs(9187)) and (layer0_outputs(4375));
    outputs(2450) <= (layer0_outputs(2591)) xor (layer0_outputs(9690));
    outputs(2451) <= not((layer0_outputs(9413)) xor (layer0_outputs(10385)));
    outputs(2452) <= (layer0_outputs(11689)) and not (layer0_outputs(6891));
    outputs(2453) <= (layer0_outputs(5548)) and (layer0_outputs(3899));
    outputs(2454) <= layer0_outputs(7189);
    outputs(2455) <= not(layer0_outputs(12026));
    outputs(2456) <= layer0_outputs(3001);
    outputs(2457) <= (layer0_outputs(11220)) and not (layer0_outputs(8524));
    outputs(2458) <= not((layer0_outputs(4601)) or (layer0_outputs(10221)));
    outputs(2459) <= (layer0_outputs(8063)) and not (layer0_outputs(11928));
    outputs(2460) <= (layer0_outputs(5832)) and not (layer0_outputs(10256));
    outputs(2461) <= (layer0_outputs(5459)) and not (layer0_outputs(3535));
    outputs(2462) <= not((layer0_outputs(10009)) or (layer0_outputs(3453)));
    outputs(2463) <= not((layer0_outputs(9735)) or (layer0_outputs(1793)));
    outputs(2464) <= not((layer0_outputs(4069)) xor (layer0_outputs(2259)));
    outputs(2465) <= (layer0_outputs(3817)) and (layer0_outputs(5953));
    outputs(2466) <= not((layer0_outputs(6479)) xor (layer0_outputs(6325)));
    outputs(2467) <= layer0_outputs(2181);
    outputs(2468) <= not((layer0_outputs(7061)) xor (layer0_outputs(2646)));
    outputs(2469) <= (layer0_outputs(2787)) and not (layer0_outputs(8321));
    outputs(2470) <= (layer0_outputs(6167)) and not (layer0_outputs(7700));
    outputs(2471) <= (layer0_outputs(2694)) xor (layer0_outputs(11220));
    outputs(2472) <= (layer0_outputs(10843)) and not (layer0_outputs(8152));
    outputs(2473) <= (layer0_outputs(4425)) and (layer0_outputs(9189));
    outputs(2474) <= not(layer0_outputs(8355));
    outputs(2475) <= (layer0_outputs(3024)) and not (layer0_outputs(2674));
    outputs(2476) <= layer0_outputs(9085);
    outputs(2477) <= (layer0_outputs(11024)) and not (layer0_outputs(6099));
    outputs(2478) <= (layer0_outputs(6007)) and not (layer0_outputs(1930));
    outputs(2479) <= not(layer0_outputs(3947));
    outputs(2480) <= not((layer0_outputs(5551)) or (layer0_outputs(7245)));
    outputs(2481) <= not((layer0_outputs(9406)) and (layer0_outputs(4159)));
    outputs(2482) <= (layer0_outputs(2153)) and not (layer0_outputs(4467));
    outputs(2483) <= layer0_outputs(3169);
    outputs(2484) <= (layer0_outputs(175)) and (layer0_outputs(4863));
    outputs(2485) <= layer0_outputs(12396);
    outputs(2486) <= (layer0_outputs(10641)) and not (layer0_outputs(3557));
    outputs(2487) <= layer0_outputs(7125);
    outputs(2488) <= (layer0_outputs(4475)) and not (layer0_outputs(7651));
    outputs(2489) <= (layer0_outputs(4981)) and (layer0_outputs(4694));
    outputs(2490) <= not(layer0_outputs(11418));
    outputs(2491) <= (layer0_outputs(8184)) and (layer0_outputs(2234));
    outputs(2492) <= not(layer0_outputs(5409));
    outputs(2493) <= (layer0_outputs(6842)) and (layer0_outputs(6920));
    outputs(2494) <= '0';
    outputs(2495) <= (layer0_outputs(2535)) and (layer0_outputs(12758));
    outputs(2496) <= layer0_outputs(9349);
    outputs(2497) <= not((layer0_outputs(11471)) xor (layer0_outputs(1953)));
    outputs(2498) <= (layer0_outputs(5012)) and not (layer0_outputs(8934));
    outputs(2499) <= (layer0_outputs(2280)) and (layer0_outputs(9820));
    outputs(2500) <= not(layer0_outputs(8514));
    outputs(2501) <= layer0_outputs(6988);
    outputs(2502) <= (layer0_outputs(7691)) and not (layer0_outputs(18));
    outputs(2503) <= layer0_outputs(12292);
    outputs(2504) <= layer0_outputs(8271);
    outputs(2505) <= (layer0_outputs(5383)) and not (layer0_outputs(3609));
    outputs(2506) <= (layer0_outputs(9781)) xor (layer0_outputs(10341));
    outputs(2507) <= not(layer0_outputs(11262));
    outputs(2508) <= (layer0_outputs(1395)) and (layer0_outputs(5224));
    outputs(2509) <= (layer0_outputs(93)) xor (layer0_outputs(3384));
    outputs(2510) <= (layer0_outputs(9253)) xor (layer0_outputs(9368));
    outputs(2511) <= (layer0_outputs(9356)) and not (layer0_outputs(5838));
    outputs(2512) <= not((layer0_outputs(4496)) or (layer0_outputs(10998)));
    outputs(2513) <= (layer0_outputs(3181)) and (layer0_outputs(6356));
    outputs(2514) <= not((layer0_outputs(9672)) or (layer0_outputs(4956)));
    outputs(2515) <= layer0_outputs(4073);
    outputs(2516) <= not((layer0_outputs(9163)) or (layer0_outputs(3403)));
    outputs(2517) <= (layer0_outputs(10383)) and not (layer0_outputs(7396));
    outputs(2518) <= '0';
    outputs(2519) <= '0';
    outputs(2520) <= (layer0_outputs(3572)) xor (layer0_outputs(4473));
    outputs(2521) <= (layer0_outputs(3082)) and not (layer0_outputs(12196));
    outputs(2522) <= (layer0_outputs(4157)) and (layer0_outputs(806));
    outputs(2523) <= (layer0_outputs(10637)) and (layer0_outputs(383));
    outputs(2524) <= (layer0_outputs(10386)) and not (layer0_outputs(9564));
    outputs(2525) <= (layer0_outputs(8507)) xor (layer0_outputs(4876));
    outputs(2526) <= (layer0_outputs(4266)) and not (layer0_outputs(8228));
    outputs(2527) <= not(layer0_outputs(3865));
    outputs(2528) <= not((layer0_outputs(1969)) xor (layer0_outputs(4270)));
    outputs(2529) <= not(layer0_outputs(9299));
    outputs(2530) <= not((layer0_outputs(10630)) xor (layer0_outputs(2990)));
    outputs(2531) <= not((layer0_outputs(7758)) xor (layer0_outputs(11522)));
    outputs(2532) <= (layer0_outputs(8542)) and (layer0_outputs(12020));
    outputs(2533) <= (layer0_outputs(7285)) xor (layer0_outputs(6957));
    outputs(2534) <= layer0_outputs(5276);
    outputs(2535) <= layer0_outputs(9626);
    outputs(2536) <= not((layer0_outputs(10347)) xor (layer0_outputs(396)));
    outputs(2537) <= layer0_outputs(12508);
    outputs(2538) <= not((layer0_outputs(3168)) xor (layer0_outputs(8288)));
    outputs(2539) <= layer0_outputs(11398);
    outputs(2540) <= (layer0_outputs(283)) and not (layer0_outputs(3297));
    outputs(2541) <= not(layer0_outputs(4540));
    outputs(2542) <= not(layer0_outputs(3668));
    outputs(2543) <= (layer0_outputs(9539)) and not (layer0_outputs(11987));
    outputs(2544) <= not((layer0_outputs(507)) or (layer0_outputs(656)));
    outputs(2545) <= (layer0_outputs(9014)) and not (layer0_outputs(240));
    outputs(2546) <= layer0_outputs(10306);
    outputs(2547) <= not((layer0_outputs(11534)) or (layer0_outputs(7849)));
    outputs(2548) <= not((layer0_outputs(8749)) xor (layer0_outputs(1612)));
    outputs(2549) <= not((layer0_outputs(4745)) xor (layer0_outputs(3731)));
    outputs(2550) <= not((layer0_outputs(5095)) or (layer0_outputs(10662)));
    outputs(2551) <= not(layer0_outputs(7988));
    outputs(2552) <= not(layer0_outputs(6653));
    outputs(2553) <= (layer0_outputs(2471)) and not (layer0_outputs(7133));
    outputs(2554) <= layer0_outputs(1152);
    outputs(2555) <= not(layer0_outputs(5198));
    outputs(2556) <= not(layer0_outputs(3854));
    outputs(2557) <= (layer0_outputs(2597)) and not (layer0_outputs(10932));
    outputs(2558) <= (layer0_outputs(8681)) and not (layer0_outputs(1455));
    outputs(2559) <= layer0_outputs(8015);
    outputs(2560) <= (layer0_outputs(1177)) and (layer0_outputs(2634));
    outputs(2561) <= not(layer0_outputs(2996));
    outputs(2562) <= not(layer0_outputs(8925));
    outputs(2563) <= (layer0_outputs(7955)) or (layer0_outputs(1094));
    outputs(2564) <= not(layer0_outputs(3018));
    outputs(2565) <= (layer0_outputs(8135)) xor (layer0_outputs(4583));
    outputs(2566) <= layer0_outputs(197);
    outputs(2567) <= (layer0_outputs(4318)) or (layer0_outputs(6656));
    outputs(2568) <= not((layer0_outputs(8859)) and (layer0_outputs(6545)));
    outputs(2569) <= not((layer0_outputs(5729)) xor (layer0_outputs(5791)));
    outputs(2570) <= not((layer0_outputs(9183)) xor (layer0_outputs(10124)));
    outputs(2571) <= layer0_outputs(5878);
    outputs(2572) <= not(layer0_outputs(5021)) or (layer0_outputs(4239));
    outputs(2573) <= not(layer0_outputs(10957));
    outputs(2574) <= not((layer0_outputs(10209)) xor (layer0_outputs(8381)));
    outputs(2575) <= not(layer0_outputs(5581));
    outputs(2576) <= not(layer0_outputs(2164));
    outputs(2577) <= not(layer0_outputs(2916)) or (layer0_outputs(12095));
    outputs(2578) <= layer0_outputs(140);
    outputs(2579) <= not(layer0_outputs(12490));
    outputs(2580) <= layer0_outputs(12367);
    outputs(2581) <= layer0_outputs(11324);
    outputs(2582) <= not(layer0_outputs(192));
    outputs(2583) <= not(layer0_outputs(12074)) or (layer0_outputs(1610));
    outputs(2584) <= layer0_outputs(12624);
    outputs(2585) <= layer0_outputs(8965);
    outputs(2586) <= (layer0_outputs(3878)) or (layer0_outputs(3686));
    outputs(2587) <= not(layer0_outputs(12282)) or (layer0_outputs(6652));
    outputs(2588) <= not(layer0_outputs(2497));
    outputs(2589) <= layer0_outputs(12285);
    outputs(2590) <= layer0_outputs(5603);
    outputs(2591) <= not((layer0_outputs(1255)) xor (layer0_outputs(2148)));
    outputs(2592) <= not(layer0_outputs(4671));
    outputs(2593) <= not(layer0_outputs(10845));
    outputs(2594) <= (layer0_outputs(3399)) xor (layer0_outputs(1426));
    outputs(2595) <= layer0_outputs(10065);
    outputs(2596) <= not(layer0_outputs(9560));
    outputs(2597) <= (layer0_outputs(8550)) or (layer0_outputs(12363));
    outputs(2598) <= layer0_outputs(7467);
    outputs(2599) <= (layer0_outputs(915)) xor (layer0_outputs(7397));
    outputs(2600) <= (layer0_outputs(3537)) and (layer0_outputs(6855));
    outputs(2601) <= not((layer0_outputs(6671)) and (layer0_outputs(3089)));
    outputs(2602) <= layer0_outputs(6746);
    outputs(2603) <= layer0_outputs(8435);
    outputs(2604) <= not(layer0_outputs(2113));
    outputs(2605) <= not((layer0_outputs(922)) xor (layer0_outputs(2362)));
    outputs(2606) <= layer0_outputs(1176);
    outputs(2607) <= not(layer0_outputs(9370));
    outputs(2608) <= (layer0_outputs(4510)) xor (layer0_outputs(9957));
    outputs(2609) <= layer0_outputs(11604);
    outputs(2610) <= layer0_outputs(2479);
    outputs(2611) <= not(layer0_outputs(11900));
    outputs(2612) <= layer0_outputs(9612);
    outputs(2613) <= layer0_outputs(2279);
    outputs(2614) <= not(layer0_outputs(10091)) or (layer0_outputs(1188));
    outputs(2615) <= not(layer0_outputs(4547));
    outputs(2616) <= not(layer0_outputs(11878));
    outputs(2617) <= layer0_outputs(10909);
    outputs(2618) <= (layer0_outputs(3925)) xor (layer0_outputs(7405));
    outputs(2619) <= (layer0_outputs(5691)) and (layer0_outputs(9556));
    outputs(2620) <= not((layer0_outputs(1679)) and (layer0_outputs(4037)));
    outputs(2621) <= layer0_outputs(4816);
    outputs(2622) <= layer0_outputs(4282);
    outputs(2623) <= not((layer0_outputs(9623)) or (layer0_outputs(2060)));
    outputs(2624) <= not(layer0_outputs(2515));
    outputs(2625) <= not(layer0_outputs(3652));
    outputs(2626) <= (layer0_outputs(9339)) or (layer0_outputs(358));
    outputs(2627) <= not(layer0_outputs(3033));
    outputs(2628) <= not(layer0_outputs(7543)) or (layer0_outputs(12240));
    outputs(2629) <= not(layer0_outputs(9693));
    outputs(2630) <= not((layer0_outputs(7797)) xor (layer0_outputs(6838)));
    outputs(2631) <= not(layer0_outputs(9085));
    outputs(2632) <= not(layer0_outputs(12358));
    outputs(2633) <= not((layer0_outputs(720)) xor (layer0_outputs(1559)));
    outputs(2634) <= layer0_outputs(8039);
    outputs(2635) <= '1';
    outputs(2636) <= layer0_outputs(9638);
    outputs(2637) <= not(layer0_outputs(7554)) or (layer0_outputs(12102));
    outputs(2638) <= not(layer0_outputs(10161));
    outputs(2639) <= layer0_outputs(981);
    outputs(2640) <= not(layer0_outputs(11455));
    outputs(2641) <= (layer0_outputs(12231)) and (layer0_outputs(7468));
    outputs(2642) <= not(layer0_outputs(6835));
    outputs(2643) <= not((layer0_outputs(9695)) and (layer0_outputs(4019)));
    outputs(2644) <= not((layer0_outputs(7333)) and (layer0_outputs(326)));
    outputs(2645) <= layer0_outputs(6743);
    outputs(2646) <= not(layer0_outputs(9920));
    outputs(2647) <= (layer0_outputs(1136)) xor (layer0_outputs(7549));
    outputs(2648) <= not(layer0_outputs(5483));
    outputs(2649) <= layer0_outputs(10817);
    outputs(2650) <= layer0_outputs(3195);
    outputs(2651) <= (layer0_outputs(523)) xor (layer0_outputs(1256));
    outputs(2652) <= (layer0_outputs(3958)) or (layer0_outputs(2152));
    outputs(2653) <= not(layer0_outputs(4671));
    outputs(2654) <= layer0_outputs(3226);
    outputs(2655) <= not(layer0_outputs(10078));
    outputs(2656) <= not(layer0_outputs(2242));
    outputs(2657) <= layer0_outputs(3900);
    outputs(2658) <= not(layer0_outputs(7622));
    outputs(2659) <= not((layer0_outputs(8796)) and (layer0_outputs(359)));
    outputs(2660) <= not((layer0_outputs(231)) and (layer0_outputs(1531)));
    outputs(2661) <= layer0_outputs(6817);
    outputs(2662) <= layer0_outputs(272);
    outputs(2663) <= not(layer0_outputs(8133));
    outputs(2664) <= not(layer0_outputs(12566)) or (layer0_outputs(3406));
    outputs(2665) <= not((layer0_outputs(11379)) xor (layer0_outputs(4743)));
    outputs(2666) <= not(layer0_outputs(4585));
    outputs(2667) <= not((layer0_outputs(12075)) xor (layer0_outputs(12187)));
    outputs(2668) <= (layer0_outputs(12761)) or (layer0_outputs(3041));
    outputs(2669) <= layer0_outputs(4931);
    outputs(2670) <= not(layer0_outputs(5280));
    outputs(2671) <= layer0_outputs(11401);
    outputs(2672) <= (layer0_outputs(7235)) or (layer0_outputs(849));
    outputs(2673) <= layer0_outputs(5463);
    outputs(2674) <= layer0_outputs(4900);
    outputs(2675) <= layer0_outputs(895);
    outputs(2676) <= not(layer0_outputs(10502));
    outputs(2677) <= layer0_outputs(11632);
    outputs(2678) <= layer0_outputs(1917);
    outputs(2679) <= layer0_outputs(2296);
    outputs(2680) <= layer0_outputs(7606);
    outputs(2681) <= not(layer0_outputs(8250));
    outputs(2682) <= not(layer0_outputs(11454));
    outputs(2683) <= layer0_outputs(5050);
    outputs(2684) <= layer0_outputs(2845);
    outputs(2685) <= not(layer0_outputs(7486));
    outputs(2686) <= not(layer0_outputs(8410)) or (layer0_outputs(12364));
    outputs(2687) <= layer0_outputs(2655);
    outputs(2688) <= not((layer0_outputs(4311)) xor (layer0_outputs(9994)));
    outputs(2689) <= layer0_outputs(8373);
    outputs(2690) <= not(layer0_outputs(6253)) or (layer0_outputs(1337));
    outputs(2691) <= (layer0_outputs(1353)) and (layer0_outputs(6117));
    outputs(2692) <= not((layer0_outputs(11555)) xor (layer0_outputs(7885)));
    outputs(2693) <= layer0_outputs(9262);
    outputs(2694) <= layer0_outputs(8249);
    outputs(2695) <= layer0_outputs(545);
    outputs(2696) <= not(layer0_outputs(2403));
    outputs(2697) <= (layer0_outputs(9986)) xor (layer0_outputs(1744));
    outputs(2698) <= layer0_outputs(4463);
    outputs(2699) <= (layer0_outputs(8579)) and (layer0_outputs(1574));
    outputs(2700) <= (layer0_outputs(4862)) or (layer0_outputs(2232));
    outputs(2701) <= layer0_outputs(4623);
    outputs(2702) <= not((layer0_outputs(9544)) xor (layer0_outputs(12229)));
    outputs(2703) <= not(layer0_outputs(8898)) or (layer0_outputs(11547));
    outputs(2704) <= layer0_outputs(712);
    outputs(2705) <= layer0_outputs(2864);
    outputs(2706) <= (layer0_outputs(1986)) xor (layer0_outputs(10123));
    outputs(2707) <= not(layer0_outputs(12223));
    outputs(2708) <= layer0_outputs(473);
    outputs(2709) <= (layer0_outputs(133)) xor (layer0_outputs(2151));
    outputs(2710) <= layer0_outputs(7746);
    outputs(2711) <= layer0_outputs(1909);
    outputs(2712) <= not(layer0_outputs(4986));
    outputs(2713) <= (layer0_outputs(3347)) and (layer0_outputs(12495));
    outputs(2714) <= not((layer0_outputs(1567)) xor (layer0_outputs(4342)));
    outputs(2715) <= not(layer0_outputs(4575));
    outputs(2716) <= layer0_outputs(8596);
    outputs(2717) <= not((layer0_outputs(7181)) and (layer0_outputs(5962)));
    outputs(2718) <= layer0_outputs(9450);
    outputs(2719) <= layer0_outputs(1161);
    outputs(2720) <= not(layer0_outputs(501));
    outputs(2721) <= not(layer0_outputs(9920));
    outputs(2722) <= (layer0_outputs(5493)) and (layer0_outputs(5941));
    outputs(2723) <= not((layer0_outputs(6815)) xor (layer0_outputs(1308)));
    outputs(2724) <= layer0_outputs(8748);
    outputs(2725) <= not(layer0_outputs(3604));
    outputs(2726) <= layer0_outputs(12108);
    outputs(2727) <= not(layer0_outputs(8868)) or (layer0_outputs(8779));
    outputs(2728) <= not((layer0_outputs(1001)) and (layer0_outputs(8501)));
    outputs(2729) <= not(layer0_outputs(12076));
    outputs(2730) <= layer0_outputs(4385);
    outputs(2731) <= layer0_outputs(7777);
    outputs(2732) <= (layer0_outputs(4606)) and not (layer0_outputs(7635));
    outputs(2733) <= layer0_outputs(10492);
    outputs(2734) <= not((layer0_outputs(2898)) xor (layer0_outputs(6446)));
    outputs(2735) <= not((layer0_outputs(9419)) xor (layer0_outputs(5056)));
    outputs(2736) <= layer0_outputs(8216);
    outputs(2737) <= (layer0_outputs(7469)) xor (layer0_outputs(4120));
    outputs(2738) <= not(layer0_outputs(9809)) or (layer0_outputs(11642));
    outputs(2739) <= not(layer0_outputs(6374));
    outputs(2740) <= not(layer0_outputs(819)) or (layer0_outputs(301));
    outputs(2741) <= not(layer0_outputs(4601));
    outputs(2742) <= (layer0_outputs(5449)) and not (layer0_outputs(12763));
    outputs(2743) <= not((layer0_outputs(1778)) and (layer0_outputs(2032)));
    outputs(2744) <= (layer0_outputs(8779)) and not (layer0_outputs(9715));
    outputs(2745) <= not((layer0_outputs(5145)) xor (layer0_outputs(11801)));
    outputs(2746) <= not(layer0_outputs(11417));
    outputs(2747) <= not((layer0_outputs(12175)) xor (layer0_outputs(3393)));
    outputs(2748) <= layer0_outputs(4243);
    outputs(2749) <= (layer0_outputs(9372)) xor (layer0_outputs(7215));
    outputs(2750) <= layer0_outputs(4463);
    outputs(2751) <= not(layer0_outputs(454));
    outputs(2752) <= layer0_outputs(5342);
    outputs(2753) <= layer0_outputs(1964);
    outputs(2754) <= not(layer0_outputs(4560));
    outputs(2755) <= (layer0_outputs(12403)) xor (layer0_outputs(7850));
    outputs(2756) <= not(layer0_outputs(10718)) or (layer0_outputs(7090));
    outputs(2757) <= not(layer0_outputs(5530));
    outputs(2758) <= layer0_outputs(459);
    outputs(2759) <= (layer0_outputs(6515)) xor (layer0_outputs(3209));
    outputs(2760) <= (layer0_outputs(11276)) or (layer0_outputs(4014));
    outputs(2761) <= (layer0_outputs(9566)) or (layer0_outputs(9233));
    outputs(2762) <= layer0_outputs(6083);
    outputs(2763) <= not(layer0_outputs(10930)) or (layer0_outputs(10948));
    outputs(2764) <= not(layer0_outputs(3979));
    outputs(2765) <= not(layer0_outputs(4547));
    outputs(2766) <= not((layer0_outputs(1414)) xor (layer0_outputs(3922)));
    outputs(2767) <= (layer0_outputs(1541)) xor (layer0_outputs(8398));
    outputs(2768) <= not((layer0_outputs(749)) xor (layer0_outputs(10797)));
    outputs(2769) <= not((layer0_outputs(9524)) and (layer0_outputs(7411)));
    outputs(2770) <= (layer0_outputs(9156)) xor (layer0_outputs(471));
    outputs(2771) <= not((layer0_outputs(1726)) xor (layer0_outputs(6159)));
    outputs(2772) <= not(layer0_outputs(9435));
    outputs(2773) <= layer0_outputs(4112);
    outputs(2774) <= layer0_outputs(1794);
    outputs(2775) <= not(layer0_outputs(9201));
    outputs(2776) <= not(layer0_outputs(11996));
    outputs(2777) <= not(layer0_outputs(11469)) or (layer0_outputs(4341));
    outputs(2778) <= layer0_outputs(4731);
    outputs(2779) <= layer0_outputs(4130);
    outputs(2780) <= not(layer0_outputs(10075));
    outputs(2781) <= (layer0_outputs(777)) and not (layer0_outputs(1390));
    outputs(2782) <= not(layer0_outputs(12659));
    outputs(2783) <= layer0_outputs(11351);
    outputs(2784) <= (layer0_outputs(11961)) and not (layer0_outputs(5111));
    outputs(2785) <= not(layer0_outputs(2584));
    outputs(2786) <= not((layer0_outputs(2415)) and (layer0_outputs(11407)));
    outputs(2787) <= (layer0_outputs(4154)) xor (layer0_outputs(4550));
    outputs(2788) <= layer0_outputs(1527);
    outputs(2789) <= not(layer0_outputs(8480));
    outputs(2790) <= not((layer0_outputs(66)) xor (layer0_outputs(6798)));
    outputs(2791) <= not(layer0_outputs(8790));
    outputs(2792) <= not(layer0_outputs(10854)) or (layer0_outputs(12079));
    outputs(2793) <= (layer0_outputs(9853)) or (layer0_outputs(6989));
    outputs(2794) <= layer0_outputs(9749);
    outputs(2795) <= not(layer0_outputs(4257));
    outputs(2796) <= not((layer0_outputs(3838)) and (layer0_outputs(10008)));
    outputs(2797) <= layer0_outputs(11720);
    outputs(2798) <= (layer0_outputs(2481)) or (layer0_outputs(3776));
    outputs(2799) <= not((layer0_outputs(11017)) xor (layer0_outputs(7031)));
    outputs(2800) <= not(layer0_outputs(7794));
    outputs(2801) <= layer0_outputs(3923);
    outputs(2802) <= (layer0_outputs(8191)) xor (layer0_outputs(8333));
    outputs(2803) <= not((layer0_outputs(1012)) and (layer0_outputs(6789)));
    outputs(2804) <= layer0_outputs(11549);
    outputs(2805) <= layer0_outputs(12788);
    outputs(2806) <= layer0_outputs(5182);
    outputs(2807) <= not(layer0_outputs(875));
    outputs(2808) <= layer0_outputs(5194);
    outputs(2809) <= not(layer0_outputs(10608)) or (layer0_outputs(4206));
    outputs(2810) <= not(layer0_outputs(2891));
    outputs(2811) <= not((layer0_outputs(502)) xor (layer0_outputs(4437)));
    outputs(2812) <= layer0_outputs(6317);
    outputs(2813) <= layer0_outputs(3709);
    outputs(2814) <= not(layer0_outputs(6707));
    outputs(2815) <= not((layer0_outputs(11132)) xor (layer0_outputs(11058)));
    outputs(2816) <= not((layer0_outputs(7747)) or (layer0_outputs(12415)));
    outputs(2817) <= layer0_outputs(3673);
    outputs(2818) <= not(layer0_outputs(10195));
    outputs(2819) <= not((layer0_outputs(1981)) xor (layer0_outputs(3998)));
    outputs(2820) <= not(layer0_outputs(385));
    outputs(2821) <= (layer0_outputs(5)) or (layer0_outputs(3622));
    outputs(2822) <= layer0_outputs(10683);
    outputs(2823) <= layer0_outputs(10160);
    outputs(2824) <= not((layer0_outputs(11655)) or (layer0_outputs(6594)));
    outputs(2825) <= (layer0_outputs(5209)) xor (layer0_outputs(12271));
    outputs(2826) <= not(layer0_outputs(2903));
    outputs(2827) <= (layer0_outputs(9240)) xor (layer0_outputs(1549));
    outputs(2828) <= not(layer0_outputs(4236)) or (layer0_outputs(5259));
    outputs(2829) <= not(layer0_outputs(10400));
    outputs(2830) <= layer0_outputs(10342);
    outputs(2831) <= (layer0_outputs(6710)) or (layer0_outputs(1701));
    outputs(2832) <= not(layer0_outputs(5718));
    outputs(2833) <= not(layer0_outputs(965));
    outputs(2834) <= not(layer0_outputs(4045));
    outputs(2835) <= not((layer0_outputs(9913)) or (layer0_outputs(11811)));
    outputs(2836) <= not(layer0_outputs(11877));
    outputs(2837) <= not((layer0_outputs(588)) and (layer0_outputs(10091)));
    outputs(2838) <= not(layer0_outputs(6992));
    outputs(2839) <= not((layer0_outputs(3497)) xor (layer0_outputs(7447)));
    outputs(2840) <= not(layer0_outputs(6736)) or (layer0_outputs(4195));
    outputs(2841) <= layer0_outputs(10125);
    outputs(2842) <= layer0_outputs(5635);
    outputs(2843) <= not(layer0_outputs(10469));
    outputs(2844) <= layer0_outputs(870);
    outputs(2845) <= (layer0_outputs(5944)) and not (layer0_outputs(3824));
    outputs(2846) <= not(layer0_outputs(217));
    outputs(2847) <= not(layer0_outputs(9990));
    outputs(2848) <= (layer0_outputs(1019)) xor (layer0_outputs(10040));
    outputs(2849) <= not(layer0_outputs(10912));
    outputs(2850) <= layer0_outputs(5505);
    outputs(2851) <= not(layer0_outputs(6457)) or (layer0_outputs(8692));
    outputs(2852) <= not(layer0_outputs(2820));
    outputs(2853) <= (layer0_outputs(8139)) xor (layer0_outputs(7613));
    outputs(2854) <= not(layer0_outputs(7909));
    outputs(2855) <= not(layer0_outputs(5143));
    outputs(2856) <= layer0_outputs(2542);
    outputs(2857) <= not((layer0_outputs(2765)) xor (layer0_outputs(4829)));
    outputs(2858) <= not(layer0_outputs(11634)) or (layer0_outputs(5882));
    outputs(2859) <= layer0_outputs(12169);
    outputs(2860) <= not((layer0_outputs(616)) xor (layer0_outputs(508)));
    outputs(2861) <= not(layer0_outputs(2916));
    outputs(2862) <= not((layer0_outputs(8241)) xor (layer0_outputs(10714)));
    outputs(2863) <= not(layer0_outputs(329));
    outputs(2864) <= layer0_outputs(5070);
    outputs(2865) <= (layer0_outputs(11039)) xor (layer0_outputs(6062));
    outputs(2866) <= not(layer0_outputs(6404));
    outputs(2867) <= (layer0_outputs(9577)) and (layer0_outputs(1837));
    outputs(2868) <= (layer0_outputs(7324)) or (layer0_outputs(11138));
    outputs(2869) <= not(layer0_outputs(6493));
    outputs(2870) <= layer0_outputs(4842);
    outputs(2871) <= not(layer0_outputs(6059));
    outputs(2872) <= layer0_outputs(5683);
    outputs(2873) <= (layer0_outputs(11940)) xor (layer0_outputs(11391));
    outputs(2874) <= not(layer0_outputs(3102));
    outputs(2875) <= not((layer0_outputs(715)) or (layer0_outputs(10481)));
    outputs(2876) <= not((layer0_outputs(6355)) and (layer0_outputs(12299)));
    outputs(2877) <= layer0_outputs(2741);
    outputs(2878) <= layer0_outputs(3844);
    outputs(2879) <= not(layer0_outputs(9665));
    outputs(2880) <= not(layer0_outputs(8484)) or (layer0_outputs(6507));
    outputs(2881) <= not((layer0_outputs(6358)) and (layer0_outputs(12688)));
    outputs(2882) <= layer0_outputs(6498);
    outputs(2883) <= layer0_outputs(10874);
    outputs(2884) <= layer0_outputs(7225);
    outputs(2885) <= not(layer0_outputs(6225));
    outputs(2886) <= not((layer0_outputs(8363)) and (layer0_outputs(11230)));
    outputs(2887) <= not((layer0_outputs(8302)) and (layer0_outputs(11097)));
    outputs(2888) <= layer0_outputs(9520);
    outputs(2889) <= not(layer0_outputs(3212));
    outputs(2890) <= (layer0_outputs(4684)) and not (layer0_outputs(2095));
    outputs(2891) <= not((layer0_outputs(10059)) and (layer0_outputs(12561)));
    outputs(2892) <= (layer0_outputs(11738)) and not (layer0_outputs(6695));
    outputs(2893) <= not((layer0_outputs(2651)) xor (layer0_outputs(4690)));
    outputs(2894) <= (layer0_outputs(10500)) or (layer0_outputs(11202));
    outputs(2895) <= not(layer0_outputs(9148));
    outputs(2896) <= layer0_outputs(9428);
    outputs(2897) <= not(layer0_outputs(5543));
    outputs(2898) <= not((layer0_outputs(3868)) and (layer0_outputs(12649)));
    outputs(2899) <= not(layer0_outputs(3346));
    outputs(2900) <= not(layer0_outputs(6586));
    outputs(2901) <= not(layer0_outputs(7865));
    outputs(2902) <= not((layer0_outputs(1625)) xor (layer0_outputs(12246)));
    outputs(2903) <= not(layer0_outputs(7392));
    outputs(2904) <= (layer0_outputs(1116)) xor (layer0_outputs(8116));
    outputs(2905) <= not(layer0_outputs(12649));
    outputs(2906) <= (layer0_outputs(10166)) xor (layer0_outputs(4740));
    outputs(2907) <= (layer0_outputs(2140)) or (layer0_outputs(5634));
    outputs(2908) <= layer0_outputs(11744);
    outputs(2909) <= layer0_outputs(12125);
    outputs(2910) <= (layer0_outputs(4706)) xor (layer0_outputs(6054));
    outputs(2911) <= (layer0_outputs(6611)) and (layer0_outputs(7209));
    outputs(2912) <= (layer0_outputs(2119)) xor (layer0_outputs(8104));
    outputs(2913) <= (layer0_outputs(3871)) xor (layer0_outputs(9132));
    outputs(2914) <= (layer0_outputs(8127)) and not (layer0_outputs(3287));
    outputs(2915) <= layer0_outputs(5493);
    outputs(2916) <= layer0_outputs(12496);
    outputs(2917) <= not((layer0_outputs(6131)) xor (layer0_outputs(7738)));
    outputs(2918) <= not(layer0_outputs(3343));
    outputs(2919) <= not(layer0_outputs(142)) or (layer0_outputs(9952));
    outputs(2920) <= not(layer0_outputs(2233));
    outputs(2921) <= (layer0_outputs(6616)) xor (layer0_outputs(633));
    outputs(2922) <= layer0_outputs(6817);
    outputs(2923) <= (layer0_outputs(8461)) and (layer0_outputs(8107));
    outputs(2924) <= not(layer0_outputs(11683));
    outputs(2925) <= not((layer0_outputs(3544)) and (layer0_outputs(2460)));
    outputs(2926) <= (layer0_outputs(9010)) and (layer0_outputs(1865));
    outputs(2927) <= not(layer0_outputs(9076));
    outputs(2928) <= layer0_outputs(2255);
    outputs(2929) <= (layer0_outputs(9716)) and (layer0_outputs(119));
    outputs(2930) <= not(layer0_outputs(1466)) or (layer0_outputs(1088));
    outputs(2931) <= not(layer0_outputs(5250));
    outputs(2932) <= layer0_outputs(12554);
    outputs(2933) <= (layer0_outputs(1178)) xor (layer0_outputs(10334));
    outputs(2934) <= (layer0_outputs(8400)) and (layer0_outputs(769));
    outputs(2935) <= layer0_outputs(5580);
    outputs(2936) <= not(layer0_outputs(4845)) or (layer0_outputs(1837));
    outputs(2937) <= not(layer0_outputs(7288)) or (layer0_outputs(3108));
    outputs(2938) <= not(layer0_outputs(4882));
    outputs(2939) <= layer0_outputs(3964);
    outputs(2940) <= layer0_outputs(5996);
    outputs(2941) <= (layer0_outputs(4247)) xor (layer0_outputs(8573));
    outputs(2942) <= not((layer0_outputs(2073)) or (layer0_outputs(5499)));
    outputs(2943) <= (layer0_outputs(4702)) xor (layer0_outputs(6302));
    outputs(2944) <= not(layer0_outputs(12424));
    outputs(2945) <= not(layer0_outputs(2829));
    outputs(2946) <= not((layer0_outputs(5108)) or (layer0_outputs(7383)));
    outputs(2947) <= layer0_outputs(1483);
    outputs(2948) <= not(layer0_outputs(3001)) or (layer0_outputs(1022));
    outputs(2949) <= not(layer0_outputs(2897));
    outputs(2950) <= (layer0_outputs(9722)) and not (layer0_outputs(6873));
    outputs(2951) <= (layer0_outputs(5818)) xor (layer0_outputs(6452));
    outputs(2952) <= not(layer0_outputs(7113));
    outputs(2953) <= (layer0_outputs(1840)) xor (layer0_outputs(11641));
    outputs(2954) <= layer0_outputs(9393);
    outputs(2955) <= (layer0_outputs(12011)) and not (layer0_outputs(4002));
    outputs(2956) <= not(layer0_outputs(1941)) or (layer0_outputs(11100));
    outputs(2957) <= not((layer0_outputs(2025)) and (layer0_outputs(9117)));
    outputs(2958) <= not(layer0_outputs(3012));
    outputs(2959) <= not(layer0_outputs(10375)) or (layer0_outputs(751));
    outputs(2960) <= not(layer0_outputs(2509)) or (layer0_outputs(5674));
    outputs(2961) <= (layer0_outputs(4656)) xor (layer0_outputs(7007));
    outputs(2962) <= not(layer0_outputs(2413));
    outputs(2963) <= not(layer0_outputs(1384));
    outputs(2964) <= not(layer0_outputs(8905));
    outputs(2965) <= not(layer0_outputs(8825));
    outputs(2966) <= not(layer0_outputs(11668)) or (layer0_outputs(4959));
    outputs(2967) <= not(layer0_outputs(7802));
    outputs(2968) <= (layer0_outputs(9502)) and (layer0_outputs(7056));
    outputs(2969) <= not(layer0_outputs(8363)) or (layer0_outputs(5799));
    outputs(2970) <= not((layer0_outputs(10282)) xor (layer0_outputs(2436)));
    outputs(2971) <= not((layer0_outputs(10997)) xor (layer0_outputs(12323)));
    outputs(2972) <= (layer0_outputs(4428)) or (layer0_outputs(5921));
    outputs(2973) <= not(layer0_outputs(5347)) or (layer0_outputs(11558));
    outputs(2974) <= layer0_outputs(9972);
    outputs(2975) <= not((layer0_outputs(11174)) and (layer0_outputs(6535)));
    outputs(2976) <= layer0_outputs(7656);
    outputs(2977) <= (layer0_outputs(10846)) xor (layer0_outputs(8706));
    outputs(2978) <= (layer0_outputs(11914)) or (layer0_outputs(11350));
    outputs(2979) <= layer0_outputs(519);
    outputs(2980) <= (layer0_outputs(6563)) or (layer0_outputs(828));
    outputs(2981) <= layer0_outputs(12574);
    outputs(2982) <= (layer0_outputs(11536)) xor (layer0_outputs(7035));
    outputs(2983) <= layer0_outputs(4050);
    outputs(2984) <= not(layer0_outputs(7618)) or (layer0_outputs(9759));
    outputs(2985) <= (layer0_outputs(4495)) xor (layer0_outputs(10870));
    outputs(2986) <= not(layer0_outputs(6354));
    outputs(2987) <= not(layer0_outputs(377));
    outputs(2988) <= layer0_outputs(3148);
    outputs(2989) <= not(layer0_outputs(2333));
    outputs(2990) <= not(layer0_outputs(2085));
    outputs(2991) <= layer0_outputs(3256);
    outputs(2992) <= (layer0_outputs(5168)) xor (layer0_outputs(5246));
    outputs(2993) <= layer0_outputs(4169);
    outputs(2994) <= (layer0_outputs(10624)) xor (layer0_outputs(8112));
    outputs(2995) <= not(layer0_outputs(4469));
    outputs(2996) <= not(layer0_outputs(4012));
    outputs(2997) <= not(layer0_outputs(3704));
    outputs(2998) <= not((layer0_outputs(7108)) xor (layer0_outputs(140)));
    outputs(2999) <= not(layer0_outputs(1311));
    outputs(3000) <= not(layer0_outputs(5588)) or (layer0_outputs(4959));
    outputs(3001) <= (layer0_outputs(6003)) and (layer0_outputs(5773));
    outputs(3002) <= not(layer0_outputs(6040));
    outputs(3003) <= not(layer0_outputs(8276));
    outputs(3004) <= not(layer0_outputs(6168));
    outputs(3005) <= layer0_outputs(9416);
    outputs(3006) <= layer0_outputs(1403);
    outputs(3007) <= not((layer0_outputs(2628)) xor (layer0_outputs(3679)));
    outputs(3008) <= not(layer0_outputs(12330)) or (layer0_outputs(5190));
    outputs(3009) <= not(layer0_outputs(11438));
    outputs(3010) <= layer0_outputs(2931);
    outputs(3011) <= (layer0_outputs(4718)) xor (layer0_outputs(166));
    outputs(3012) <= (layer0_outputs(9494)) xor (layer0_outputs(11658));
    outputs(3013) <= not(layer0_outputs(11085));
    outputs(3014) <= not(layer0_outputs(9379));
    outputs(3015) <= not(layer0_outputs(8306)) or (layer0_outputs(5889));
    outputs(3016) <= not((layer0_outputs(1214)) and (layer0_outputs(6741)));
    outputs(3017) <= (layer0_outputs(2741)) and not (layer0_outputs(561));
    outputs(3018) <= not(layer0_outputs(1207));
    outputs(3019) <= not((layer0_outputs(475)) xor (layer0_outputs(1595)));
    outputs(3020) <= not(layer0_outputs(10984)) or (layer0_outputs(10467));
    outputs(3021) <= layer0_outputs(3690);
    outputs(3022) <= not(layer0_outputs(2047));
    outputs(3023) <= layer0_outputs(9400);
    outputs(3024) <= (layer0_outputs(980)) or (layer0_outputs(9502));
    outputs(3025) <= not(layer0_outputs(5312)) or (layer0_outputs(3358));
    outputs(3026) <= not((layer0_outputs(7932)) or (layer0_outputs(7129)));
    outputs(3027) <= not((layer0_outputs(2661)) and (layer0_outputs(3309)));
    outputs(3028) <= layer0_outputs(4395);
    outputs(3029) <= not(layer0_outputs(7523)) or (layer0_outputs(10573));
    outputs(3030) <= layer0_outputs(3506);
    outputs(3031) <= (layer0_outputs(5957)) xor (layer0_outputs(7286));
    outputs(3032) <= layer0_outputs(10453);
    outputs(3033) <= layer0_outputs(2517);
    outputs(3034) <= (layer0_outputs(5090)) xor (layer0_outputs(3797));
    outputs(3035) <= not(layer0_outputs(6017));
    outputs(3036) <= not((layer0_outputs(2726)) xor (layer0_outputs(5162)));
    outputs(3037) <= (layer0_outputs(4080)) and (layer0_outputs(9734));
    outputs(3038) <= not((layer0_outputs(5269)) xor (layer0_outputs(649)));
    outputs(3039) <= (layer0_outputs(11958)) or (layer0_outputs(7280));
    outputs(3040) <= (layer0_outputs(4655)) xor (layer0_outputs(3675));
    outputs(3041) <= not((layer0_outputs(8379)) and (layer0_outputs(573)));
    outputs(3042) <= (layer0_outputs(246)) xor (layer0_outputs(12193));
    outputs(3043) <= layer0_outputs(5182);
    outputs(3044) <= (layer0_outputs(382)) or (layer0_outputs(7414));
    outputs(3045) <= not(layer0_outputs(7697));
    outputs(3046) <= not(layer0_outputs(7757));
    outputs(3047) <= (layer0_outputs(6220)) xor (layer0_outputs(3233));
    outputs(3048) <= not((layer0_outputs(1869)) xor (layer0_outputs(2464)));
    outputs(3049) <= (layer0_outputs(8365)) xor (layer0_outputs(6305));
    outputs(3050) <= not(layer0_outputs(10866)) or (layer0_outputs(2666));
    outputs(3051) <= layer0_outputs(5133);
    outputs(3052) <= not(layer0_outputs(957));
    outputs(3053) <= not(layer0_outputs(10161));
    outputs(3054) <= not(layer0_outputs(7710));
    outputs(3055) <= not((layer0_outputs(4008)) and (layer0_outputs(2483)));
    outputs(3056) <= not(layer0_outputs(4592)) or (layer0_outputs(12699));
    outputs(3057) <= not(layer0_outputs(4507));
    outputs(3058) <= not((layer0_outputs(606)) xor (layer0_outputs(8558)));
    outputs(3059) <= (layer0_outputs(7368)) and not (layer0_outputs(6361));
    outputs(3060) <= not(layer0_outputs(11732));
    outputs(3061) <= not(layer0_outputs(7936)) or (layer0_outputs(10434));
    outputs(3062) <= (layer0_outputs(5401)) or (layer0_outputs(1184));
    outputs(3063) <= not(layer0_outputs(2579));
    outputs(3064) <= not(layer0_outputs(5301));
    outputs(3065) <= layer0_outputs(12417);
    outputs(3066) <= layer0_outputs(181);
    outputs(3067) <= layer0_outputs(827);
    outputs(3068) <= not((layer0_outputs(12732)) and (layer0_outputs(12737)));
    outputs(3069) <= not((layer0_outputs(10242)) xor (layer0_outputs(1374)));
    outputs(3070) <= (layer0_outputs(5286)) xor (layer0_outputs(10496));
    outputs(3071) <= (layer0_outputs(10275)) and not (layer0_outputs(10040));
    outputs(3072) <= layer0_outputs(6352);
    outputs(3073) <= layer0_outputs(6944);
    outputs(3074) <= layer0_outputs(137);
    outputs(3075) <= (layer0_outputs(10074)) and (layer0_outputs(5878));
    outputs(3076) <= layer0_outputs(5106);
    outputs(3077) <= not(layer0_outputs(4994)) or (layer0_outputs(11633));
    outputs(3078) <= not(layer0_outputs(2529));
    outputs(3079) <= (layer0_outputs(9577)) and (layer0_outputs(1892));
    outputs(3080) <= (layer0_outputs(11306)) xor (layer0_outputs(3828));
    outputs(3081) <= (layer0_outputs(12064)) xor (layer0_outputs(2101));
    outputs(3082) <= not((layer0_outputs(11886)) and (layer0_outputs(6110)));
    outputs(3083) <= (layer0_outputs(2039)) and not (layer0_outputs(6704));
    outputs(3084) <= not(layer0_outputs(6241)) or (layer0_outputs(4831));
    outputs(3085) <= not(layer0_outputs(1801)) or (layer0_outputs(3777));
    outputs(3086) <= layer0_outputs(12093);
    outputs(3087) <= layer0_outputs(7457);
    outputs(3088) <= not(layer0_outputs(7399));
    outputs(3089) <= layer0_outputs(5618);
    outputs(3090) <= not(layer0_outputs(12620));
    outputs(3091) <= not(layer0_outputs(6784)) or (layer0_outputs(2676));
    outputs(3092) <= layer0_outputs(1450);
    outputs(3093) <= not((layer0_outputs(728)) and (layer0_outputs(12566)));
    outputs(3094) <= layer0_outputs(7374);
    outputs(3095) <= not(layer0_outputs(965));
    outputs(3096) <= not(layer0_outputs(760));
    outputs(3097) <= not((layer0_outputs(431)) and (layer0_outputs(10750)));
    outputs(3098) <= (layer0_outputs(1832)) xor (layer0_outputs(3196));
    outputs(3099) <= not(layer0_outputs(1359));
    outputs(3100) <= layer0_outputs(2762);
    outputs(3101) <= not((layer0_outputs(1286)) or (layer0_outputs(6983)));
    outputs(3102) <= not(layer0_outputs(6967));
    outputs(3103) <= not(layer0_outputs(3368)) or (layer0_outputs(7803));
    outputs(3104) <= layer0_outputs(7092);
    outputs(3105) <= not(layer0_outputs(2830));
    outputs(3106) <= layer0_outputs(462);
    outputs(3107) <= layer0_outputs(7720);
    outputs(3108) <= not(layer0_outputs(12233)) or (layer0_outputs(8851));
    outputs(3109) <= not((layer0_outputs(1301)) or (layer0_outputs(6403)));
    outputs(3110) <= (layer0_outputs(8349)) xor (layer0_outputs(1782));
    outputs(3111) <= not(layer0_outputs(10730));
    outputs(3112) <= layer0_outputs(3940);
    outputs(3113) <= not((layer0_outputs(6045)) xor (layer0_outputs(6638)));
    outputs(3114) <= not(layer0_outputs(338));
    outputs(3115) <= not(layer0_outputs(8202));
    outputs(3116) <= (layer0_outputs(1284)) xor (layer0_outputs(1792));
    outputs(3117) <= layer0_outputs(12635);
    outputs(3118) <= not((layer0_outputs(11995)) xor (layer0_outputs(8849)));
    outputs(3119) <= (layer0_outputs(11967)) or (layer0_outputs(3523));
    outputs(3120) <= not((layer0_outputs(662)) xor (layer0_outputs(4458)));
    outputs(3121) <= layer0_outputs(6331);
    outputs(3122) <= not((layer0_outputs(5861)) and (layer0_outputs(1710)));
    outputs(3123) <= (layer0_outputs(4299)) xor (layer0_outputs(7339));
    outputs(3124) <= not(layer0_outputs(2407)) or (layer0_outputs(7627));
    outputs(3125) <= not((layer0_outputs(10775)) xor (layer0_outputs(1748)));
    outputs(3126) <= not(layer0_outputs(1732));
    outputs(3127) <= layer0_outputs(5636);
    outputs(3128) <= layer0_outputs(5290);
    outputs(3129) <= not(layer0_outputs(11105));
    outputs(3130) <= not(layer0_outputs(10531));
    outputs(3131) <= not(layer0_outputs(7592));
    outputs(3132) <= not(layer0_outputs(7267));
    outputs(3133) <= not(layer0_outputs(3704));
    outputs(3134) <= layer0_outputs(3268);
    outputs(3135) <= (layer0_outputs(7736)) xor (layer0_outputs(3003));
    outputs(3136) <= layer0_outputs(11132);
    outputs(3137) <= (layer0_outputs(11106)) and (layer0_outputs(11004));
    outputs(3138) <= layer0_outputs(2734);
    outputs(3139) <= (layer0_outputs(7268)) xor (layer0_outputs(807));
    outputs(3140) <= (layer0_outputs(12498)) and (layer0_outputs(4412));
    outputs(3141) <= not(layer0_outputs(9208));
    outputs(3142) <= not((layer0_outputs(2950)) and (layer0_outputs(4952)));
    outputs(3143) <= not(layer0_outputs(2796));
    outputs(3144) <= not(layer0_outputs(10297)) or (layer0_outputs(4835));
    outputs(3145) <= not(layer0_outputs(808));
    outputs(3146) <= not(layer0_outputs(12463));
    outputs(3147) <= not((layer0_outputs(8731)) xor (layer0_outputs(12355)));
    outputs(3148) <= not(layer0_outputs(12571));
    outputs(3149) <= layer0_outputs(11080);
    outputs(3150) <= (layer0_outputs(2370)) xor (layer0_outputs(2913));
    outputs(3151) <= not(layer0_outputs(5771)) or (layer0_outputs(12754));
    outputs(3152) <= layer0_outputs(7848);
    outputs(3153) <= (layer0_outputs(9982)) xor (layer0_outputs(3067));
    outputs(3154) <= not(layer0_outputs(11192)) or (layer0_outputs(9280));
    outputs(3155) <= (layer0_outputs(4402)) and not (layer0_outputs(9595));
    outputs(3156) <= (layer0_outputs(6080)) xor (layer0_outputs(8563));
    outputs(3157) <= layer0_outputs(2409);
    outputs(3158) <= (layer0_outputs(1588)) and not (layer0_outputs(66));
    outputs(3159) <= layer0_outputs(6539);
    outputs(3160) <= (layer0_outputs(8209)) xor (layer0_outputs(7960));
    outputs(3161) <= layer0_outputs(2067);
    outputs(3162) <= not(layer0_outputs(4549));
    outputs(3163) <= layer0_outputs(9683);
    outputs(3164) <= not(layer0_outputs(11253));
    outputs(3165) <= not(layer0_outputs(5234));
    outputs(3166) <= (layer0_outputs(171)) xor (layer0_outputs(9866));
    outputs(3167) <= not((layer0_outputs(10619)) and (layer0_outputs(7400)));
    outputs(3168) <= not(layer0_outputs(5478)) or (layer0_outputs(8162));
    outputs(3169) <= not((layer0_outputs(7659)) and (layer0_outputs(1998)));
    outputs(3170) <= layer0_outputs(9567);
    outputs(3171) <= layer0_outputs(1230);
    outputs(3172) <= (layer0_outputs(4062)) and not (layer0_outputs(1977));
    outputs(3173) <= layer0_outputs(228);
    outputs(3174) <= (layer0_outputs(6514)) xor (layer0_outputs(1821));
    outputs(3175) <= not((layer0_outputs(5040)) and (layer0_outputs(4570)));
    outputs(3176) <= not((layer0_outputs(7735)) xor (layer0_outputs(9748)));
    outputs(3177) <= not(layer0_outputs(11506));
    outputs(3178) <= not((layer0_outputs(8483)) xor (layer0_outputs(8703)));
    outputs(3179) <= not(layer0_outputs(7516));
    outputs(3180) <= not((layer0_outputs(4888)) and (layer0_outputs(4113)));
    outputs(3181) <= not((layer0_outputs(12676)) xor (layer0_outputs(48)));
    outputs(3182) <= not(layer0_outputs(1836));
    outputs(3183) <= (layer0_outputs(10103)) xor (layer0_outputs(10759));
    outputs(3184) <= (layer0_outputs(10925)) and not (layer0_outputs(2096));
    outputs(3185) <= not(layer0_outputs(7500));
    outputs(3186) <= (layer0_outputs(1901)) xor (layer0_outputs(11784));
    outputs(3187) <= layer0_outputs(11104);
    outputs(3188) <= layer0_outputs(594);
    outputs(3189) <= layer0_outputs(8737);
    outputs(3190) <= not(layer0_outputs(4466));
    outputs(3191) <= not(layer0_outputs(12051));
    outputs(3192) <= layer0_outputs(11730);
    outputs(3193) <= layer0_outputs(2429);
    outputs(3194) <= not(layer0_outputs(4510));
    outputs(3195) <= (layer0_outputs(4154)) xor (layer0_outputs(5051));
    outputs(3196) <= not(layer0_outputs(10350)) or (layer0_outputs(1016));
    outputs(3197) <= layer0_outputs(7655);
    outputs(3198) <= layer0_outputs(6437);
    outputs(3199) <= not(layer0_outputs(8861));
    outputs(3200) <= layer0_outputs(7759);
    outputs(3201) <= not((layer0_outputs(6486)) xor (layer0_outputs(1794)));
    outputs(3202) <= layer0_outputs(4714);
    outputs(3203) <= not((layer0_outputs(7686)) and (layer0_outputs(9325)));
    outputs(3204) <= layer0_outputs(7306);
    outputs(3205) <= not(layer0_outputs(7422)) or (layer0_outputs(3497));
    outputs(3206) <= not(layer0_outputs(9445)) or (layer0_outputs(5952));
    outputs(3207) <= layer0_outputs(600);
    outputs(3208) <= layer0_outputs(697);
    outputs(3209) <= (layer0_outputs(102)) and not (layer0_outputs(6059));
    outputs(3210) <= not(layer0_outputs(10137)) or (layer0_outputs(2281));
    outputs(3211) <= not(layer0_outputs(4505));
    outputs(3212) <= (layer0_outputs(10830)) xor (layer0_outputs(2221));
    outputs(3213) <= layer0_outputs(9362);
    outputs(3214) <= not(layer0_outputs(12654));
    outputs(3215) <= (layer0_outputs(250)) and not (layer0_outputs(11774));
    outputs(3216) <= not(layer0_outputs(10298));
    outputs(3217) <= (layer0_outputs(4875)) xor (layer0_outputs(9467));
    outputs(3218) <= not((layer0_outputs(8009)) xor (layer0_outputs(7346)));
    outputs(3219) <= not(layer0_outputs(4484));
    outputs(3220) <= not(layer0_outputs(12794));
    outputs(3221) <= not(layer0_outputs(4043));
    outputs(3222) <= not(layer0_outputs(4968));
    outputs(3223) <= not((layer0_outputs(5304)) or (layer0_outputs(11341)));
    outputs(3224) <= not(layer0_outputs(1876));
    outputs(3225) <= not(layer0_outputs(11332)) or (layer0_outputs(8958));
    outputs(3226) <= not((layer0_outputs(3317)) xor (layer0_outputs(1507)));
    outputs(3227) <= layer0_outputs(5385);
    outputs(3228) <= (layer0_outputs(10749)) and not (layer0_outputs(9620));
    outputs(3229) <= layer0_outputs(982);
    outputs(3230) <= layer0_outputs(6623);
    outputs(3231) <= layer0_outputs(2617);
    outputs(3232) <= (layer0_outputs(11141)) or (layer0_outputs(11615));
    outputs(3233) <= layer0_outputs(6117);
    outputs(3234) <= not((layer0_outputs(3932)) xor (layer0_outputs(6525)));
    outputs(3235) <= layer0_outputs(11408);
    outputs(3236) <= not(layer0_outputs(10765));
    outputs(3237) <= not((layer0_outputs(2456)) xor (layer0_outputs(6613)));
    outputs(3238) <= not(layer0_outputs(5046));
    outputs(3239) <= layer0_outputs(4757);
    outputs(3240) <= (layer0_outputs(2870)) xor (layer0_outputs(5035));
    outputs(3241) <= not(layer0_outputs(3147)) or (layer0_outputs(11716));
    outputs(3242) <= (layer0_outputs(11847)) xor (layer0_outputs(11628));
    outputs(3243) <= layer0_outputs(7581);
    outputs(3244) <= not(layer0_outputs(10603));
    outputs(3245) <= not(layer0_outputs(7873));
    outputs(3246) <= (layer0_outputs(11982)) xor (layer0_outputs(4539));
    outputs(3247) <= (layer0_outputs(4465)) and not (layer0_outputs(7526));
    outputs(3248) <= not((layer0_outputs(2451)) and (layer0_outputs(1370)));
    outputs(3249) <= not(layer0_outputs(12076));
    outputs(3250) <= not(layer0_outputs(12290));
    outputs(3251) <= not(layer0_outputs(11412));
    outputs(3252) <= layer0_outputs(7270);
    outputs(3253) <= layer0_outputs(7672);
    outputs(3254) <= layer0_outputs(4964);
    outputs(3255) <= (layer0_outputs(10173)) and not (layer0_outputs(1407));
    outputs(3256) <= not(layer0_outputs(4607));
    outputs(3257) <= layer0_outputs(7815);
    outputs(3258) <= not((layer0_outputs(921)) xor (layer0_outputs(10152)));
    outputs(3259) <= layer0_outputs(3392);
    outputs(3260) <= layer0_outputs(6753);
    outputs(3261) <= (layer0_outputs(1923)) or (layer0_outputs(9243));
    outputs(3262) <= not(layer0_outputs(4012));
    outputs(3263) <= layer0_outputs(8818);
    outputs(3264) <= (layer0_outputs(9404)) xor (layer0_outputs(7948));
    outputs(3265) <= (layer0_outputs(7822)) or (layer0_outputs(5743));
    outputs(3266) <= layer0_outputs(7382);
    outputs(3267) <= not(layer0_outputs(787));
    outputs(3268) <= (layer0_outputs(5388)) and (layer0_outputs(6098));
    outputs(3269) <= layer0_outputs(9357);
    outputs(3270) <= (layer0_outputs(392)) xor (layer0_outputs(1985));
    outputs(3271) <= not(layer0_outputs(10122));
    outputs(3272) <= not((layer0_outputs(7124)) xor (layer0_outputs(5158)));
    outputs(3273) <= layer0_outputs(1860);
    outputs(3274) <= (layer0_outputs(11650)) or (layer0_outputs(3384));
    outputs(3275) <= not(layer0_outputs(22));
    outputs(3276) <= not((layer0_outputs(11523)) or (layer0_outputs(1682)));
    outputs(3277) <= (layer0_outputs(10430)) xor (layer0_outputs(4791));
    outputs(3278) <= layer0_outputs(3784);
    outputs(3279) <= not((layer0_outputs(3173)) xor (layer0_outputs(1361)));
    outputs(3280) <= layer0_outputs(7884);
    outputs(3281) <= not(layer0_outputs(9844));
    outputs(3282) <= not((layer0_outputs(1949)) xor (layer0_outputs(10784)));
    outputs(3283) <= layer0_outputs(9941);
    outputs(3284) <= not(layer0_outputs(1173)) or (layer0_outputs(6378));
    outputs(3285) <= not((layer0_outputs(11023)) xor (layer0_outputs(7208)));
    outputs(3286) <= layer0_outputs(2098);
    outputs(3287) <= not(layer0_outputs(8725));
    outputs(3288) <= not(layer0_outputs(9437));
    outputs(3289) <= not(layer0_outputs(1685));
    outputs(3290) <= layer0_outputs(37);
    outputs(3291) <= not((layer0_outputs(3552)) and (layer0_outputs(3787)));
    outputs(3292) <= not((layer0_outputs(8481)) xor (layer0_outputs(7999)));
    outputs(3293) <= not(layer0_outputs(8925)) or (layer0_outputs(3130));
    outputs(3294) <= not((layer0_outputs(5079)) and (layer0_outputs(11590)));
    outputs(3295) <= layer0_outputs(7979);
    outputs(3296) <= layer0_outputs(4632);
    outputs(3297) <= layer0_outputs(2145);
    outputs(3298) <= not(layer0_outputs(11732));
    outputs(3299) <= not((layer0_outputs(3507)) xor (layer0_outputs(650)));
    outputs(3300) <= layer0_outputs(8001);
    outputs(3301) <= layer0_outputs(11607);
    outputs(3302) <= not(layer0_outputs(7880));
    outputs(3303) <= not((layer0_outputs(9898)) xor (layer0_outputs(9510)));
    outputs(3304) <= not((layer0_outputs(5471)) xor (layer0_outputs(11557)));
    outputs(3305) <= not(layer0_outputs(5717)) or (layer0_outputs(7672));
    outputs(3306) <= not((layer0_outputs(7993)) xor (layer0_outputs(5028)));
    outputs(3307) <= layer0_outputs(4506);
    outputs(3308) <= layer0_outputs(11380);
    outputs(3309) <= not((layer0_outputs(11700)) xor (layer0_outputs(2415)));
    outputs(3310) <= layer0_outputs(7940);
    outputs(3311) <= not(layer0_outputs(12395));
    outputs(3312) <= not(layer0_outputs(1731));
    outputs(3313) <= not(layer0_outputs(5873)) or (layer0_outputs(1073));
    outputs(3314) <= not((layer0_outputs(294)) xor (layer0_outputs(6883)));
    outputs(3315) <= not(layer0_outputs(11506));
    outputs(3316) <= layer0_outputs(9176);
    outputs(3317) <= (layer0_outputs(7297)) and (layer0_outputs(2614));
    outputs(3318) <= layer0_outputs(9209);
    outputs(3319) <= layer0_outputs(8092);
    outputs(3320) <= layer0_outputs(7440);
    outputs(3321) <= (layer0_outputs(2775)) xor (layer0_outputs(1603));
    outputs(3322) <= (layer0_outputs(9511)) and not (layer0_outputs(10074));
    outputs(3323) <= not(layer0_outputs(6077)) or (layer0_outputs(5449));
    outputs(3324) <= not(layer0_outputs(9081));
    outputs(3325) <= layer0_outputs(3921);
    outputs(3326) <= not(layer0_outputs(3791));
    outputs(3327) <= not(layer0_outputs(4365)) or (layer0_outputs(7813));
    outputs(3328) <= (layer0_outputs(10857)) xor (layer0_outputs(12104));
    outputs(3329) <= layer0_outputs(9681);
    outputs(3330) <= not((layer0_outputs(8660)) xor (layer0_outputs(4150)));
    outputs(3331) <= not((layer0_outputs(554)) xor (layer0_outputs(3958)));
    outputs(3332) <= layer0_outputs(7867);
    outputs(3333) <= not(layer0_outputs(3929));
    outputs(3334) <= not((layer0_outputs(9597)) and (layer0_outputs(9964)));
    outputs(3335) <= not(layer0_outputs(10848)) or (layer0_outputs(8908));
    outputs(3336) <= layer0_outputs(2740);
    outputs(3337) <= not((layer0_outputs(1473)) xor (layer0_outputs(5018)));
    outputs(3338) <= not((layer0_outputs(3333)) or (layer0_outputs(566)));
    outputs(3339) <= not(layer0_outputs(6639));
    outputs(3340) <= not(layer0_outputs(5968));
    outputs(3341) <= not(layer0_outputs(12351));
    outputs(3342) <= not(layer0_outputs(5810));
    outputs(3343) <= (layer0_outputs(7144)) and not (layer0_outputs(11757));
    outputs(3344) <= (layer0_outputs(2813)) or (layer0_outputs(12764));
    outputs(3345) <= layer0_outputs(4080);
    outputs(3346) <= not((layer0_outputs(7527)) xor (layer0_outputs(2785)));
    outputs(3347) <= (layer0_outputs(4782)) xor (layer0_outputs(4489));
    outputs(3348) <= not(layer0_outputs(11078));
    outputs(3349) <= not(layer0_outputs(7548));
    outputs(3350) <= not((layer0_outputs(3398)) or (layer0_outputs(2037)));
    outputs(3351) <= layer0_outputs(11675);
    outputs(3352) <= (layer0_outputs(9145)) xor (layer0_outputs(3526));
    outputs(3353) <= (layer0_outputs(4752)) or (layer0_outputs(5876));
    outputs(3354) <= (layer0_outputs(4577)) and (layer0_outputs(3156));
    outputs(3355) <= (layer0_outputs(5909)) and not (layer0_outputs(9782));
    outputs(3356) <= not(layer0_outputs(2352));
    outputs(3357) <= layer0_outputs(10628);
    outputs(3358) <= not((layer0_outputs(2284)) xor (layer0_outputs(10472)));
    outputs(3359) <= layer0_outputs(10786);
    outputs(3360) <= not(layer0_outputs(2286));
    outputs(3361) <= (layer0_outputs(2643)) or (layer0_outputs(7009));
    outputs(3362) <= not(layer0_outputs(3373));
    outputs(3363) <= not((layer0_outputs(2109)) and (layer0_outputs(9281)));
    outputs(3364) <= layer0_outputs(8578);
    outputs(3365) <= layer0_outputs(5949);
    outputs(3366) <= layer0_outputs(10976);
    outputs(3367) <= (layer0_outputs(9622)) xor (layer0_outputs(4787));
    outputs(3368) <= layer0_outputs(12575);
    outputs(3369) <= not((layer0_outputs(9950)) and (layer0_outputs(9140)));
    outputs(3370) <= not(layer0_outputs(955));
    outputs(3371) <= (layer0_outputs(3885)) xor (layer0_outputs(3505));
    outputs(3372) <= not(layer0_outputs(2462));
    outputs(3373) <= not(layer0_outputs(12668)) or (layer0_outputs(10507));
    outputs(3374) <= layer0_outputs(11335);
    outputs(3375) <= not(layer0_outputs(7079));
    outputs(3376) <= not(layer0_outputs(9744));
    outputs(3377) <= not(layer0_outputs(534));
    outputs(3378) <= (layer0_outputs(9238)) and (layer0_outputs(11863));
    outputs(3379) <= not(layer0_outputs(6954));
    outputs(3380) <= not(layer0_outputs(12010));
    outputs(3381) <= not(layer0_outputs(4871));
    outputs(3382) <= (layer0_outputs(8694)) xor (layer0_outputs(6469));
    outputs(3383) <= not((layer0_outputs(3241)) xor (layer0_outputs(2619)));
    outputs(3384) <= not((layer0_outputs(7931)) xor (layer0_outputs(6824)));
    outputs(3385) <= layer0_outputs(11211);
    outputs(3386) <= (layer0_outputs(4325)) or (layer0_outputs(5148));
    outputs(3387) <= not(layer0_outputs(7239));
    outputs(3388) <= not((layer0_outputs(524)) xor (layer0_outputs(7698)));
    outputs(3389) <= not(layer0_outputs(1064));
    outputs(3390) <= (layer0_outputs(9631)) and (layer0_outputs(11741));
    outputs(3391) <= not((layer0_outputs(9370)) and (layer0_outputs(2097)));
    outputs(3392) <= (layer0_outputs(3673)) or (layer0_outputs(3956));
    outputs(3393) <= not(layer0_outputs(10198));
    outputs(3394) <= not(layer0_outputs(12207));
    outputs(3395) <= layer0_outputs(5698);
    outputs(3396) <= (layer0_outputs(11230)) and not (layer0_outputs(3294));
    outputs(3397) <= not(layer0_outputs(12589)) or (layer0_outputs(4028));
    outputs(3398) <= (layer0_outputs(4511)) and not (layer0_outputs(2269));
    outputs(3399) <= layer0_outputs(1984);
    outputs(3400) <= (layer0_outputs(4884)) and (layer0_outputs(4465));
    outputs(3401) <= layer0_outputs(12359);
    outputs(3402) <= layer0_outputs(10240);
    outputs(3403) <= not(layer0_outputs(9242));
    outputs(3404) <= (layer0_outputs(389)) and not (layer0_outputs(7586));
    outputs(3405) <= not(layer0_outputs(1209));
    outputs(3406) <= not((layer0_outputs(7196)) xor (layer0_outputs(4125)));
    outputs(3407) <= not((layer0_outputs(1439)) xor (layer0_outputs(1142)));
    outputs(3408) <= not(layer0_outputs(3202)) or (layer0_outputs(11990));
    outputs(3409) <= not((layer0_outputs(10175)) and (layer0_outputs(7422)));
    outputs(3410) <= (layer0_outputs(598)) or (layer0_outputs(96));
    outputs(3411) <= (layer0_outputs(2077)) and (layer0_outputs(32));
    outputs(3412) <= not(layer0_outputs(3555));
    outputs(3413) <= layer0_outputs(5382);
    outputs(3414) <= (layer0_outputs(12340)) and not (layer0_outputs(6651));
    outputs(3415) <= not((layer0_outputs(5327)) xor (layer0_outputs(9112)));
    outputs(3416) <= not((layer0_outputs(4226)) xor (layer0_outputs(10658)));
    outputs(3417) <= layer0_outputs(12350);
    outputs(3418) <= layer0_outputs(3312);
    outputs(3419) <= layer0_outputs(4943);
    outputs(3420) <= not(layer0_outputs(6842));
    outputs(3421) <= not(layer0_outputs(671)) or (layer0_outputs(2260));
    outputs(3422) <= not(layer0_outputs(8553));
    outputs(3423) <= layer0_outputs(8837);
    outputs(3424) <= not(layer0_outputs(3637));
    outputs(3425) <= not(layer0_outputs(7396));
    outputs(3426) <= layer0_outputs(370);
    outputs(3427) <= not((layer0_outputs(11728)) or (layer0_outputs(4405)));
    outputs(3428) <= not(layer0_outputs(11539));
    outputs(3429) <= not(layer0_outputs(8637));
    outputs(3430) <= not(layer0_outputs(698));
    outputs(3431) <= layer0_outputs(3998);
    outputs(3432) <= not((layer0_outputs(1250)) and (layer0_outputs(5544)));
    outputs(3433) <= layer0_outputs(10449);
    outputs(3434) <= (layer0_outputs(3066)) xor (layer0_outputs(3665));
    outputs(3435) <= not(layer0_outputs(7272)) or (layer0_outputs(4638));
    outputs(3436) <= not(layer0_outputs(2397));
    outputs(3437) <= layer0_outputs(10550);
    outputs(3438) <= not(layer0_outputs(10055));
    outputs(3439) <= (layer0_outputs(5152)) xor (layer0_outputs(11151));
    outputs(3440) <= layer0_outputs(4512);
    outputs(3441) <= (layer0_outputs(7203)) xor (layer0_outputs(10964));
    outputs(3442) <= not(layer0_outputs(9196)) or (layer0_outputs(9142));
    outputs(3443) <= not(layer0_outputs(5205));
    outputs(3444) <= layer0_outputs(6344);
    outputs(3445) <= layer0_outputs(9633);
    outputs(3446) <= not(layer0_outputs(3652));
    outputs(3447) <= not(layer0_outputs(682)) or (layer0_outputs(11010));
    outputs(3448) <= not((layer0_outputs(8061)) and (layer0_outputs(2111)));
    outputs(3449) <= (layer0_outputs(10425)) xor (layer0_outputs(5041));
    outputs(3450) <= not(layer0_outputs(12199));
    outputs(3451) <= (layer0_outputs(5365)) and not (layer0_outputs(8262));
    outputs(3452) <= (layer0_outputs(12660)) and not (layer0_outputs(12642));
    outputs(3453) <= (layer0_outputs(132)) and (layer0_outputs(7652));
    outputs(3454) <= not((layer0_outputs(7343)) xor (layer0_outputs(4893)));
    outputs(3455) <= not(layer0_outputs(5025));
    outputs(3456) <= not((layer0_outputs(6296)) xor (layer0_outputs(8576)));
    outputs(3457) <= (layer0_outputs(7751)) xor (layer0_outputs(3259));
    outputs(3458) <= not(layer0_outputs(11542));
    outputs(3459) <= not(layer0_outputs(5502)) or (layer0_outputs(2864));
    outputs(3460) <= not(layer0_outputs(10777));
    outputs(3461) <= not((layer0_outputs(1571)) xor (layer0_outputs(7576)));
    outputs(3462) <= layer0_outputs(7663);
    outputs(3463) <= (layer0_outputs(4945)) xor (layer0_outputs(8846));
    outputs(3464) <= (layer0_outputs(12787)) xor (layer0_outputs(2942));
    outputs(3465) <= layer0_outputs(39);
    outputs(3466) <= not(layer0_outputs(10067));
    outputs(3467) <= not(layer0_outputs(7710));
    outputs(3468) <= layer0_outputs(7147);
    outputs(3469) <= (layer0_outputs(5142)) and not (layer0_outputs(4779));
    outputs(3470) <= layer0_outputs(12215);
    outputs(3471) <= not(layer0_outputs(423)) or (layer0_outputs(11296));
    outputs(3472) <= (layer0_outputs(8666)) xor (layer0_outputs(9710));
    outputs(3473) <= layer0_outputs(5532);
    outputs(3474) <= (layer0_outputs(8733)) and (layer0_outputs(3606));
    outputs(3475) <= not(layer0_outputs(6232));
    outputs(3476) <= not(layer0_outputs(6225));
    outputs(3477) <= layer0_outputs(5869);
    outputs(3478) <= not(layer0_outputs(6471)) or (layer0_outputs(8961));
    outputs(3479) <= not(layer0_outputs(8697));
    outputs(3480) <= not(layer0_outputs(11362));
    outputs(3481) <= not(layer0_outputs(5412));
    outputs(3482) <= layer0_outputs(9017);
    outputs(3483) <= not(layer0_outputs(164));
    outputs(3484) <= not(layer0_outputs(10959));
    outputs(3485) <= not((layer0_outputs(2033)) xor (layer0_outputs(10883)));
    outputs(3486) <= not(layer0_outputs(12690));
    outputs(3487) <= not(layer0_outputs(1552)) or (layer0_outputs(196));
    outputs(3488) <= not((layer0_outputs(6132)) and (layer0_outputs(1929)));
    outputs(3489) <= not((layer0_outputs(4614)) or (layer0_outputs(2979)));
    outputs(3490) <= not(layer0_outputs(4042)) or (layer0_outputs(11283));
    outputs(3491) <= layer0_outputs(51);
    outputs(3492) <= (layer0_outputs(4599)) and not (layer0_outputs(9540));
    outputs(3493) <= not((layer0_outputs(6642)) and (layer0_outputs(4995)));
    outputs(3494) <= not(layer0_outputs(94)) or (layer0_outputs(4851));
    outputs(3495) <= (layer0_outputs(5094)) xor (layer0_outputs(7798));
    outputs(3496) <= layer0_outputs(10644);
    outputs(3497) <= not(layer0_outputs(9640));
    outputs(3498) <= not((layer0_outputs(9012)) xor (layer0_outputs(6174)));
    outputs(3499) <= layer0_outputs(6352);
    outputs(3500) <= layer0_outputs(2227);
    outputs(3501) <= (layer0_outputs(12008)) xor (layer0_outputs(3643));
    outputs(3502) <= (layer0_outputs(1799)) xor (layer0_outputs(2584));
    outputs(3503) <= not(layer0_outputs(2465));
    outputs(3504) <= not(layer0_outputs(5601));
    outputs(3505) <= not(layer0_outputs(9990)) or (layer0_outputs(1648));
    outputs(3506) <= not((layer0_outputs(2179)) xor (layer0_outputs(11006)));
    outputs(3507) <= layer0_outputs(11191);
    outputs(3508) <= (layer0_outputs(3691)) and not (layer0_outputs(6026));
    outputs(3509) <= not(layer0_outputs(6106)) or (layer0_outputs(10518));
    outputs(3510) <= not(layer0_outputs(4376));
    outputs(3511) <= (layer0_outputs(1734)) and (layer0_outputs(7953));
    outputs(3512) <= not(layer0_outputs(11687));
    outputs(3513) <= not((layer0_outputs(11470)) and (layer0_outputs(2776)));
    outputs(3514) <= not(layer0_outputs(1250));
    outputs(3515) <= (layer0_outputs(2294)) or (layer0_outputs(3513));
    outputs(3516) <= (layer0_outputs(10820)) or (layer0_outputs(6022));
    outputs(3517) <= not(layer0_outputs(6375));
    outputs(3518) <= (layer0_outputs(635)) xor (layer0_outputs(1718));
    outputs(3519) <= (layer0_outputs(5112)) xor (layer0_outputs(6385));
    outputs(3520) <= layer0_outputs(10626);
    outputs(3521) <= not((layer0_outputs(6511)) xor (layer0_outputs(9600)));
    outputs(3522) <= layer0_outputs(8499);
    outputs(3523) <= (layer0_outputs(10263)) and not (layer0_outputs(860));
    outputs(3524) <= (layer0_outputs(6986)) or (layer0_outputs(3123));
    outputs(3525) <= not(layer0_outputs(5559));
    outputs(3526) <= not(layer0_outputs(7994)) or (layer0_outputs(5279));
    outputs(3527) <= layer0_outputs(6207);
    outputs(3528) <= not((layer0_outputs(10269)) xor (layer0_outputs(8711)));
    outputs(3529) <= layer0_outputs(5054);
    outputs(3530) <= not((layer0_outputs(1784)) xor (layer0_outputs(7839)));
    outputs(3531) <= not(layer0_outputs(745)) or (layer0_outputs(7041));
    outputs(3532) <= not(layer0_outputs(9821)) or (layer0_outputs(3501));
    outputs(3533) <= layer0_outputs(11961);
    outputs(3534) <= not((layer0_outputs(5485)) xor (layer0_outputs(5536)));
    outputs(3535) <= not((layer0_outputs(10269)) xor (layer0_outputs(1620)));
    outputs(3536) <= not(layer0_outputs(2166));
    outputs(3537) <= not(layer0_outputs(10743));
    outputs(3538) <= not((layer0_outputs(7815)) xor (layer0_outputs(6153)));
    outputs(3539) <= (layer0_outputs(11134)) xor (layer0_outputs(3595));
    outputs(3540) <= layer0_outputs(4806);
    outputs(3541) <= layer0_outputs(6331);
    outputs(3542) <= not(layer0_outputs(7110));
    outputs(3543) <= not(layer0_outputs(6300)) or (layer0_outputs(1591));
    outputs(3544) <= (layer0_outputs(5728)) xor (layer0_outputs(4381));
    outputs(3545) <= (layer0_outputs(2569)) xor (layer0_outputs(11904));
    outputs(3546) <= not(layer0_outputs(4963));
    outputs(3547) <= (layer0_outputs(8166)) xor (layer0_outputs(11070));
    outputs(3548) <= layer0_outputs(7150);
    outputs(3549) <= (layer0_outputs(9235)) xor (layer0_outputs(5105));
    outputs(3550) <= not((layer0_outputs(9860)) xor (layer0_outputs(12111)));
    outputs(3551) <= not(layer0_outputs(8746));
    outputs(3552) <= not(layer0_outputs(12328)) or (layer0_outputs(11993));
    outputs(3553) <= not((layer0_outputs(10700)) or (layer0_outputs(995)));
    outputs(3554) <= layer0_outputs(3083);
    outputs(3555) <= layer0_outputs(9504);
    outputs(3556) <= layer0_outputs(11317);
    outputs(3557) <= layer0_outputs(3926);
    outputs(3558) <= layer0_outputs(4001);
    outputs(3559) <= (layer0_outputs(6619)) or (layer0_outputs(9204));
    outputs(3560) <= layer0_outputs(11569);
    outputs(3561) <= not(layer0_outputs(12290)) or (layer0_outputs(11474));
    outputs(3562) <= not((layer0_outputs(3417)) xor (layer0_outputs(6668)));
    outputs(3563) <= not(layer0_outputs(8688)) or (layer0_outputs(10409));
    outputs(3564) <= not(layer0_outputs(11533)) or (layer0_outputs(8080));
    outputs(3565) <= not((layer0_outputs(7419)) and (layer0_outputs(6773)));
    outputs(3566) <= not(layer0_outputs(8729));
    outputs(3567) <= not(layer0_outputs(8305));
    outputs(3568) <= not((layer0_outputs(9551)) xor (layer0_outputs(8122)));
    outputs(3569) <= not((layer0_outputs(10781)) and (layer0_outputs(2667)));
    outputs(3570) <= (layer0_outputs(1993)) xor (layer0_outputs(11083));
    outputs(3571) <= not((layer0_outputs(4735)) and (layer0_outputs(4345)));
    outputs(3572) <= (layer0_outputs(5077)) and (layer0_outputs(7957));
    outputs(3573) <= (layer0_outputs(5345)) and not (layer0_outputs(6302));
    outputs(3574) <= layer0_outputs(5154);
    outputs(3575) <= layer0_outputs(5177);
    outputs(3576) <= layer0_outputs(9618);
    outputs(3577) <= layer0_outputs(12754);
    outputs(3578) <= not(layer0_outputs(291)) or (layer0_outputs(12023));
    outputs(3579) <= (layer0_outputs(4811)) or (layer0_outputs(11670));
    outputs(3580) <= layer0_outputs(10557);
    outputs(3581) <= not((layer0_outputs(12532)) xor (layer0_outputs(4965)));
    outputs(3582) <= (layer0_outputs(1196)) xor (layer0_outputs(4938));
    outputs(3583) <= (layer0_outputs(4849)) xor (layer0_outputs(9261));
    outputs(3584) <= not((layer0_outputs(244)) xor (layer0_outputs(9425)));
    outputs(3585) <= not((layer0_outputs(4212)) or (layer0_outputs(10926)));
    outputs(3586) <= layer0_outputs(1767);
    outputs(3587) <= (layer0_outputs(2797)) or (layer0_outputs(2975));
    outputs(3588) <= not(layer0_outputs(1833)) or (layer0_outputs(12746));
    outputs(3589) <= not((layer0_outputs(7621)) xor (layer0_outputs(5910)));
    outputs(3590) <= not((layer0_outputs(11879)) and (layer0_outputs(3779)));
    outputs(3591) <= not((layer0_outputs(6129)) or (layer0_outputs(4159)));
    outputs(3592) <= not(layer0_outputs(3091));
    outputs(3593) <= layer0_outputs(9604);
    outputs(3594) <= not((layer0_outputs(8266)) xor (layer0_outputs(8887)));
    outputs(3595) <= not(layer0_outputs(2909)) or (layer0_outputs(3546));
    outputs(3596) <= (layer0_outputs(4669)) or (layer0_outputs(58));
    outputs(3597) <= not((layer0_outputs(1508)) xor (layer0_outputs(5083)));
    outputs(3598) <= layer0_outputs(4947);
    outputs(3599) <= (layer0_outputs(1443)) xor (layer0_outputs(12162));
    outputs(3600) <= not(layer0_outputs(8132));
    outputs(3601) <= not(layer0_outputs(6041));
    outputs(3602) <= layer0_outputs(2568);
    outputs(3603) <= not((layer0_outputs(11012)) and (layer0_outputs(11581)));
    outputs(3604) <= (layer0_outputs(6684)) xor (layer0_outputs(10491));
    outputs(3605) <= not((layer0_outputs(11602)) xor (layer0_outputs(6621)));
    outputs(3606) <= layer0_outputs(6896);
    outputs(3607) <= layer0_outputs(2641);
    outputs(3608) <= not((layer0_outputs(2412)) and (layer0_outputs(539)));
    outputs(3609) <= layer0_outputs(11288);
    outputs(3610) <= (layer0_outputs(225)) and (layer0_outputs(2851));
    outputs(3611) <= not(layer0_outputs(10193));
    outputs(3612) <= (layer0_outputs(7446)) xor (layer0_outputs(7170));
    outputs(3613) <= not((layer0_outputs(1251)) and (layer0_outputs(10847)));
    outputs(3614) <= not(layer0_outputs(10990));
    outputs(3615) <= layer0_outputs(2548);
    outputs(3616) <= layer0_outputs(7602);
    outputs(3617) <= not(layer0_outputs(4323)) or (layer0_outputs(12041));
    outputs(3618) <= layer0_outputs(9427);
    outputs(3619) <= not((layer0_outputs(10681)) and (layer0_outputs(3484)));
    outputs(3620) <= (layer0_outputs(7057)) and not (layer0_outputs(8814));
    outputs(3621) <= (layer0_outputs(8080)) and (layer0_outputs(9652));
    outputs(3622) <= not(layer0_outputs(6556));
    outputs(3623) <= (layer0_outputs(7337)) or (layer0_outputs(1259));
    outputs(3624) <= (layer0_outputs(932)) or (layer0_outputs(3496));
    outputs(3625) <= not(layer0_outputs(7377));
    outputs(3626) <= not((layer0_outputs(3427)) xor (layer0_outputs(3176)));
    outputs(3627) <= layer0_outputs(11178);
    outputs(3628) <= (layer0_outputs(675)) or (layer0_outputs(5839));
    outputs(3629) <= (layer0_outputs(6540)) xor (layer0_outputs(7886));
    outputs(3630) <= not(layer0_outputs(12619));
    outputs(3631) <= not(layer0_outputs(9146)) or (layer0_outputs(2477));
    outputs(3632) <= (layer0_outputs(7149)) xor (layer0_outputs(9621));
    outputs(3633) <= not(layer0_outputs(7375));
    outputs(3634) <= layer0_outputs(10788);
    outputs(3635) <= not(layer0_outputs(9662));
    outputs(3636) <= not(layer0_outputs(5850));
    outputs(3637) <= not(layer0_outputs(5767)) or (layer0_outputs(7695));
    outputs(3638) <= not(layer0_outputs(7654));
    outputs(3639) <= not(layer0_outputs(4274));
    outputs(3640) <= not((layer0_outputs(5782)) and (layer0_outputs(2587)));
    outputs(3641) <= layer0_outputs(798);
    outputs(3642) <= layer0_outputs(3488);
    outputs(3643) <= not(layer0_outputs(338));
    outputs(3644) <= layer0_outputs(9392);
    outputs(3645) <= not((layer0_outputs(9178)) xor (layer0_outputs(8601)));
    outputs(3646) <= not((layer0_outputs(10865)) or (layer0_outputs(7766)));
    outputs(3647) <= not(layer0_outputs(2107));
    outputs(3648) <= (layer0_outputs(780)) xor (layer0_outputs(8734));
    outputs(3649) <= '1';
    outputs(3650) <= layer0_outputs(4449);
    outputs(3651) <= not((layer0_outputs(7745)) xor (layer0_outputs(5462)));
    outputs(3652) <= not((layer0_outputs(2961)) xor (layer0_outputs(12200)));
    outputs(3653) <= not((layer0_outputs(3747)) xor (layer0_outputs(6788)));
    outputs(3654) <= not(layer0_outputs(12356)) or (layer0_outputs(3801));
    outputs(3655) <= not(layer0_outputs(3660));
    outputs(3656) <= (layer0_outputs(2500)) and not (layer0_outputs(4444));
    outputs(3657) <= not(layer0_outputs(2877)) or (layer0_outputs(3058));
    outputs(3658) <= (layer0_outputs(3152)) and (layer0_outputs(11118));
    outputs(3659) <= not((layer0_outputs(9859)) xor (layer0_outputs(2192)));
    outputs(3660) <= (layer0_outputs(2811)) xor (layer0_outputs(11799));
    outputs(3661) <= layer0_outputs(9058);
    outputs(3662) <= layer0_outputs(8472);
    outputs(3663) <= layer0_outputs(7388);
    outputs(3664) <= not(layer0_outputs(8615)) or (layer0_outputs(2749));
    outputs(3665) <= (layer0_outputs(8224)) xor (layer0_outputs(10181));
    outputs(3666) <= (layer0_outputs(7865)) xor (layer0_outputs(9075));
    outputs(3667) <= not((layer0_outputs(12433)) and (layer0_outputs(9192)));
    outputs(3668) <= (layer0_outputs(842)) and (layer0_outputs(7004));
    outputs(3669) <= layer0_outputs(339);
    outputs(3670) <= not(layer0_outputs(6168));
    outputs(3671) <= (layer0_outputs(9995)) xor (layer0_outputs(6872));
    outputs(3672) <= not(layer0_outputs(9424));
    outputs(3673) <= not(layer0_outputs(11025));
    outputs(3674) <= not(layer0_outputs(11396));
    outputs(3675) <= not(layer0_outputs(2082));
    outputs(3676) <= not(layer0_outputs(5320)) or (layer0_outputs(11055));
    outputs(3677) <= layer0_outputs(12295);
    outputs(3678) <= not(layer0_outputs(6120));
    outputs(3679) <= layer0_outputs(5311);
    outputs(3680) <= (layer0_outputs(9028)) xor (layer0_outputs(3320));
    outputs(3681) <= layer0_outputs(3541);
    outputs(3682) <= layer0_outputs(12138);
    outputs(3683) <= not(layer0_outputs(2665));
    outputs(3684) <= (layer0_outputs(9776)) xor (layer0_outputs(11587));
    outputs(3685) <= (layer0_outputs(2368)) xor (layer0_outputs(7833));
    outputs(3686) <= layer0_outputs(12052);
    outputs(3687) <= layer0_outputs(4879);
    outputs(3688) <= not(layer0_outputs(2841)) or (layer0_outputs(1350));
    outputs(3689) <= layer0_outputs(1861);
    outputs(3690) <= not(layer0_outputs(11027));
    outputs(3691) <= (layer0_outputs(1834)) and not (layer0_outputs(12521));
    outputs(3692) <= not((layer0_outputs(3141)) or (layer0_outputs(558)));
    outputs(3693) <= not(layer0_outputs(8088)) or (layer0_outputs(5642));
    outputs(3694) <= not((layer0_outputs(8888)) xor (layer0_outputs(1050)));
    outputs(3695) <= not((layer0_outputs(1497)) xor (layer0_outputs(189)));
    outputs(3696) <= not((layer0_outputs(5179)) and (layer0_outputs(3306)));
    outputs(3697) <= not(layer0_outputs(11146)) or (layer0_outputs(6811));
    outputs(3698) <= not((layer0_outputs(848)) and (layer0_outputs(3047)));
    outputs(3699) <= not(layer0_outputs(8843));
    outputs(3700) <= not(layer0_outputs(5109));
    outputs(3701) <= (layer0_outputs(6474)) or (layer0_outputs(3948));
    outputs(3702) <= (layer0_outputs(3720)) and (layer0_outputs(2167));
    outputs(3703) <= not(layer0_outputs(4937));
    outputs(3704) <= not(layer0_outputs(9632)) or (layer0_outputs(4568));
    outputs(3705) <= layer0_outputs(4782);
    outputs(3706) <= not(layer0_outputs(7332));
    outputs(3707) <= layer0_outputs(7362);
    outputs(3708) <= not(layer0_outputs(3593)) or (layer0_outputs(6831));
    outputs(3709) <= layer0_outputs(973);
    outputs(3710) <= layer0_outputs(6248);
    outputs(3711) <= not((layer0_outputs(7077)) and (layer0_outputs(6410)));
    outputs(3712) <= layer0_outputs(6213);
    outputs(3713) <= not(layer0_outputs(5748));
    outputs(3714) <= not(layer0_outputs(6579)) or (layer0_outputs(10929));
    outputs(3715) <= (layer0_outputs(2378)) xor (layer0_outputs(5658));
    outputs(3716) <= layer0_outputs(1023);
    outputs(3717) <= (layer0_outputs(1009)) xor (layer0_outputs(1512));
    outputs(3718) <= not(layer0_outputs(1945)) or (layer0_outputs(127));
    outputs(3719) <= not(layer0_outputs(8626));
    outputs(3720) <= (layer0_outputs(1331)) and not (layer0_outputs(6269));
    outputs(3721) <= (layer0_outputs(4730)) or (layer0_outputs(12757));
    outputs(3722) <= not((layer0_outputs(9073)) and (layer0_outputs(12161)));
    outputs(3723) <= not(layer0_outputs(5430));
    outputs(3724) <= not((layer0_outputs(10534)) xor (layer0_outputs(10112)));
    outputs(3725) <= not(layer0_outputs(4636));
    outputs(3726) <= not(layer0_outputs(8686));
    outputs(3727) <= (layer0_outputs(2220)) xor (layer0_outputs(8874));
    outputs(3728) <= layer0_outputs(8094);
    outputs(3729) <= (layer0_outputs(4010)) xor (layer0_outputs(12677));
    outputs(3730) <= (layer0_outputs(3312)) or (layer0_outputs(10710));
    outputs(3731) <= not(layer0_outputs(2939));
    outputs(3732) <= layer0_outputs(12504);
    outputs(3733) <= not(layer0_outputs(11074));
    outputs(3734) <= layer0_outputs(6781);
    outputs(3735) <= (layer0_outputs(8620)) and (layer0_outputs(6533));
    outputs(3736) <= layer0_outputs(6883);
    outputs(3737) <= layer0_outputs(6216);
    outputs(3738) <= (layer0_outputs(2676)) or (layer0_outputs(2470));
    outputs(3739) <= layer0_outputs(6507);
    outputs(3740) <= layer0_outputs(5241);
    outputs(3741) <= layer0_outputs(222);
    outputs(3742) <= not((layer0_outputs(6113)) xor (layer0_outputs(8265)));
    outputs(3743) <= not(layer0_outputs(1654));
    outputs(3744) <= layer0_outputs(2784);
    outputs(3745) <= layer0_outputs(11564);
    outputs(3746) <= (layer0_outputs(7728)) and not (layer0_outputs(11726));
    outputs(3747) <= not((layer0_outputs(435)) xor (layer0_outputs(12260)));
    outputs(3748) <= not(layer0_outputs(6764)) or (layer0_outputs(2995));
    outputs(3749) <= not((layer0_outputs(1537)) xor (layer0_outputs(4293)));
    outputs(3750) <= not(layer0_outputs(2171));
    outputs(3751) <= not(layer0_outputs(11019));
    outputs(3752) <= layer0_outputs(6975);
    outputs(3753) <= not((layer0_outputs(12621)) and (layer0_outputs(12568)));
    outputs(3754) <= layer0_outputs(7508);
    outputs(3755) <= not(layer0_outputs(1166)) or (layer0_outputs(5756));
    outputs(3756) <= layer0_outputs(6722);
    outputs(3757) <= layer0_outputs(4438);
    outputs(3758) <= not(layer0_outputs(3986)) or (layer0_outputs(1202));
    outputs(3759) <= (layer0_outputs(6261)) xor (layer0_outputs(3351));
    outputs(3760) <= not(layer0_outputs(6585));
    outputs(3761) <= not(layer0_outputs(340));
    outputs(3762) <= layer0_outputs(7428);
    outputs(3763) <= layer0_outputs(6010);
    outputs(3764) <= (layer0_outputs(7087)) xor (layer0_outputs(5606));
    outputs(3765) <= not(layer0_outputs(3467));
    outputs(3766) <= not(layer0_outputs(3834));
    outputs(3767) <= not(layer0_outputs(2988));
    outputs(3768) <= layer0_outputs(7250);
    outputs(3769) <= not((layer0_outputs(1092)) xor (layer0_outputs(5040)));
    outputs(3770) <= layer0_outputs(6303);
    outputs(3771) <= not(layer0_outputs(11920));
    outputs(3772) <= not((layer0_outputs(6142)) xor (layer0_outputs(8990)));
    outputs(3773) <= not((layer0_outputs(8280)) xor (layer0_outputs(10928)));
    outputs(3774) <= layer0_outputs(10578);
    outputs(3775) <= layer0_outputs(4383);
    outputs(3776) <= not(layer0_outputs(6373));
    outputs(3777) <= layer0_outputs(2030);
    outputs(3778) <= (layer0_outputs(740)) xor (layer0_outputs(833));
    outputs(3779) <= (layer0_outputs(10044)) and (layer0_outputs(4044));
    outputs(3780) <= layer0_outputs(103);
    outputs(3781) <= layer0_outputs(536);
    outputs(3782) <= not((layer0_outputs(3702)) xor (layer0_outputs(12245)));
    outputs(3783) <= not((layer0_outputs(9760)) xor (layer0_outputs(1210)));
    outputs(3784) <= (layer0_outputs(9660)) xor (layer0_outputs(9847));
    outputs(3785) <= layer0_outputs(85);
    outputs(3786) <= (layer0_outputs(5143)) xor (layer0_outputs(8656));
    outputs(3787) <= not(layer0_outputs(8530));
    outputs(3788) <= not((layer0_outputs(6006)) xor (layer0_outputs(5703)));
    outputs(3789) <= not(layer0_outputs(2901));
    outputs(3790) <= not(layer0_outputs(8930));
    outputs(3791) <= layer0_outputs(9114);
    outputs(3792) <= not(layer0_outputs(3272));
    outputs(3793) <= not(layer0_outputs(401));
    outputs(3794) <= not(layer0_outputs(5920));
    outputs(3795) <= not(layer0_outputs(11266)) or (layer0_outputs(10695));
    outputs(3796) <= not(layer0_outputs(8774)) or (layer0_outputs(2259));
    outputs(3797) <= not((layer0_outputs(12374)) or (layer0_outputs(873)));
    outputs(3798) <= not(layer0_outputs(6953));
    outputs(3799) <= (layer0_outputs(7446)) xor (layer0_outputs(10120));
    outputs(3800) <= layer0_outputs(213);
    outputs(3801) <= not((layer0_outputs(10827)) xor (layer0_outputs(10434)));
    outputs(3802) <= not((layer0_outputs(9184)) xor (layer0_outputs(11060)));
    outputs(3803) <= layer0_outputs(5361);
    outputs(3804) <= not(layer0_outputs(10822));
    outputs(3805) <= not((layer0_outputs(169)) xor (layer0_outputs(5597)));
    outputs(3806) <= layer0_outputs(1118);
    outputs(3807) <= layer0_outputs(6995);
    outputs(3808) <= (layer0_outputs(1483)) xor (layer0_outputs(1599));
    outputs(3809) <= layer0_outputs(9565);
    outputs(3810) <= not((layer0_outputs(7709)) xor (layer0_outputs(9315)));
    outputs(3811) <= (layer0_outputs(936)) or (layer0_outputs(5639));
    outputs(3812) <= not(layer0_outputs(8048));
    outputs(3813) <= not(layer0_outputs(7563));
    outputs(3814) <= not(layer0_outputs(679)) or (layer0_outputs(11792));
    outputs(3815) <= not((layer0_outputs(6773)) or (layer0_outputs(611)));
    outputs(3816) <= not(layer0_outputs(6281));
    outputs(3817) <= not(layer0_outputs(4849));
    outputs(3818) <= layer0_outputs(5343);
    outputs(3819) <= layer0_outputs(7606);
    outputs(3820) <= not(layer0_outputs(9490)) or (layer0_outputs(6405));
    outputs(3821) <= not(layer0_outputs(7636));
    outputs(3822) <= not(layer0_outputs(10833));
    outputs(3823) <= not(layer0_outputs(1614));
    outputs(3824) <= not((layer0_outputs(3225)) xor (layer0_outputs(5850)));
    outputs(3825) <= (layer0_outputs(7682)) or (layer0_outputs(2103));
    outputs(3826) <= not(layer0_outputs(8792));
    outputs(3827) <= layer0_outputs(11397);
    outputs(3828) <= layer0_outputs(557);
    outputs(3829) <= not(layer0_outputs(9857));
    outputs(3830) <= layer0_outputs(9351);
    outputs(3831) <= not(layer0_outputs(10238));
    outputs(3832) <= (layer0_outputs(9446)) xor (layer0_outputs(9302));
    outputs(3833) <= not(layer0_outputs(1128)) or (layer0_outputs(8724));
    outputs(3834) <= layer0_outputs(4410);
    outputs(3835) <= not(layer0_outputs(11612));
    outputs(3836) <= '1';
    outputs(3837) <= not(layer0_outputs(3945));
    outputs(3838) <= layer0_outputs(4189);
    outputs(3839) <= layer0_outputs(25);
    outputs(3840) <= not((layer0_outputs(1481)) or (layer0_outputs(5024)));
    outputs(3841) <= layer0_outputs(6314);
    outputs(3842) <= layer0_outputs(6002);
    outputs(3843) <= not(layer0_outputs(8852));
    outputs(3844) <= (layer0_outputs(12296)) and not (layer0_outputs(12426));
    outputs(3845) <= (layer0_outputs(1496)) and (layer0_outputs(11043));
    outputs(3846) <= not((layer0_outputs(5895)) xor (layer0_outputs(2801)));
    outputs(3847) <= not(layer0_outputs(4819));
    outputs(3848) <= (layer0_outputs(8164)) and (layer0_outputs(4204));
    outputs(3849) <= layer0_outputs(2620);
    outputs(3850) <= not(layer0_outputs(8610));
    outputs(3851) <= layer0_outputs(4616);
    outputs(3852) <= not((layer0_outputs(3939)) or (layer0_outputs(7166)));
    outputs(3853) <= (layer0_outputs(871)) and not (layer0_outputs(4534));
    outputs(3854) <= not(layer0_outputs(5034));
    outputs(3855) <= layer0_outputs(555);
    outputs(3856) <= not(layer0_outputs(235));
    outputs(3857) <= not((layer0_outputs(6991)) xor (layer0_outputs(3803)));
    outputs(3858) <= (layer0_outputs(6194)) and not (layer0_outputs(7172));
    outputs(3859) <= not(layer0_outputs(10120));
    outputs(3860) <= layer0_outputs(10546);
    outputs(3861) <= not(layer0_outputs(11592)) or (layer0_outputs(7319));
    outputs(3862) <= layer0_outputs(203);
    outputs(3863) <= (layer0_outputs(3132)) and not (layer0_outputs(1530));
    outputs(3864) <= not(layer0_outputs(2948)) or (layer0_outputs(735));
    outputs(3865) <= not(layer0_outputs(118));
    outputs(3866) <= not(layer0_outputs(2475));
    outputs(3867) <= (layer0_outputs(3234)) and (layer0_outputs(3927));
    outputs(3868) <= (layer0_outputs(4016)) or (layer0_outputs(11315));
    outputs(3869) <= not(layer0_outputs(8493));
    outputs(3870) <= (layer0_outputs(1785)) xor (layer0_outputs(1456));
    outputs(3871) <= layer0_outputs(1346);
    outputs(3872) <= not(layer0_outputs(7628));
    outputs(3873) <= layer0_outputs(8194);
    outputs(3874) <= not((layer0_outputs(6980)) xor (layer0_outputs(6709)));
    outputs(3875) <= layer0_outputs(3473);
    outputs(3876) <= layer0_outputs(9696);
    outputs(3877) <= (layer0_outputs(2837)) and (layer0_outputs(9345));
    outputs(3878) <= (layer0_outputs(4473)) and (layer0_outputs(9985));
    outputs(3879) <= (layer0_outputs(3736)) xor (layer0_outputs(11752));
    outputs(3880) <= not((layer0_outputs(724)) xor (layer0_outputs(1748)));
    outputs(3881) <= layer0_outputs(1956);
    outputs(3882) <= not(layer0_outputs(10100));
    outputs(3883) <= (layer0_outputs(11434)) xor (layer0_outputs(6723));
    outputs(3884) <= not((layer0_outputs(987)) and (layer0_outputs(12652)));
    outputs(3885) <= not((layer0_outputs(2020)) xor (layer0_outputs(1852)));
    outputs(3886) <= not((layer0_outputs(12189)) xor (layer0_outputs(922)));
    outputs(3887) <= (layer0_outputs(11614)) xor (layer0_outputs(4423));
    outputs(3888) <= not(layer0_outputs(8441));
    outputs(3889) <= (layer0_outputs(8277)) or (layer0_outputs(8465));
    outputs(3890) <= not(layer0_outputs(11087));
    outputs(3891) <= (layer0_outputs(4399)) and (layer0_outputs(11894));
    outputs(3892) <= layer0_outputs(10232);
    outputs(3893) <= (layer0_outputs(2502)) and not (layer0_outputs(3879));
    outputs(3894) <= (layer0_outputs(3641)) or (layer0_outputs(8330));
    outputs(3895) <= (layer0_outputs(6233)) and not (layer0_outputs(7633));
    outputs(3896) <= not(layer0_outputs(3073)) or (layer0_outputs(1730));
    outputs(3897) <= layer0_outputs(11628);
    outputs(3898) <= layer0_outputs(12292);
    outputs(3899) <= not(layer0_outputs(4202)) or (layer0_outputs(6521));
    outputs(3900) <= (layer0_outputs(10796)) and (layer0_outputs(9171));
    outputs(3901) <= layer0_outputs(5883);
    outputs(3902) <= (layer0_outputs(4339)) and not (layer0_outputs(472));
    outputs(3903) <= (layer0_outputs(466)) xor (layer0_outputs(10706));
    outputs(3904) <= (layer0_outputs(2648)) xor (layer0_outputs(11667));
    outputs(3905) <= layer0_outputs(6688);
    outputs(3906) <= (layer0_outputs(1590)) and not (layer0_outputs(3364));
    outputs(3907) <= not((layer0_outputs(6251)) and (layer0_outputs(3953)));
    outputs(3908) <= (layer0_outputs(4478)) and not (layer0_outputs(4467));
    outputs(3909) <= layer0_outputs(8175);
    outputs(3910) <= not(layer0_outputs(9101));
    outputs(3911) <= (layer0_outputs(10270)) and (layer0_outputs(6255));
    outputs(3912) <= (layer0_outputs(7979)) and (layer0_outputs(11177));
    outputs(3913) <= not(layer0_outputs(8998)) or (layer0_outputs(2017));
    outputs(3914) <= not((layer0_outputs(5820)) xor (layer0_outputs(3674)));
    outputs(3915) <= layer0_outputs(5177);
    outputs(3916) <= (layer0_outputs(11598)) and not (layer0_outputs(12005));
    outputs(3917) <= (layer0_outputs(3188)) xor (layer0_outputs(10800));
    outputs(3918) <= not(layer0_outputs(9159)) or (layer0_outputs(900));
    outputs(3919) <= (layer0_outputs(9149)) and not (layer0_outputs(1694));
    outputs(3920) <= layer0_outputs(8692);
    outputs(3921) <= layer0_outputs(4089);
    outputs(3922) <= (layer0_outputs(8037)) and not (layer0_outputs(7771));
    outputs(3923) <= (layer0_outputs(4409)) and not (layer0_outputs(7896));
    outputs(3924) <= layer0_outputs(8237);
    outputs(3925) <= not(layer0_outputs(3184));
    outputs(3926) <= layer0_outputs(4955);
    outputs(3927) <= layer0_outputs(12541);
    outputs(3928) <= (layer0_outputs(10850)) and (layer0_outputs(1521));
    outputs(3929) <= not((layer0_outputs(6972)) or (layer0_outputs(4419)));
    outputs(3930) <= (layer0_outputs(1618)) xor (layer0_outputs(8534));
    outputs(3931) <= layer0_outputs(11043);
    outputs(3932) <= layer0_outputs(8345);
    outputs(3933) <= layer0_outputs(9511);
    outputs(3934) <= layer0_outputs(11749);
    outputs(3935) <= not(layer0_outputs(1958)) or (layer0_outputs(5078));
    outputs(3936) <= not(layer0_outputs(11972)) or (layer0_outputs(4682));
    outputs(3937) <= not((layer0_outputs(8150)) xor (layer0_outputs(9157)));
    outputs(3938) <= layer0_outputs(7211);
    outputs(3939) <= (layer0_outputs(5440)) and not (layer0_outputs(4998));
    outputs(3940) <= layer0_outputs(206);
    outputs(3941) <= not((layer0_outputs(3088)) xor (layer0_outputs(4542)));
    outputs(3942) <= (layer0_outputs(10610)) and (layer0_outputs(4326));
    outputs(3943) <= (layer0_outputs(2313)) xor (layer0_outputs(4347));
    outputs(3944) <= not(layer0_outputs(2878));
    outputs(3945) <= (layer0_outputs(650)) and (layer0_outputs(12576));
    outputs(3946) <= (layer0_outputs(2168)) xor (layer0_outputs(9528));
    outputs(3947) <= not(layer0_outputs(9295));
    outputs(3948) <= (layer0_outputs(10501)) or (layer0_outputs(6909));
    outputs(3949) <= not(layer0_outputs(1409));
    outputs(3950) <= (layer0_outputs(11624)) or (layer0_outputs(6256));
    outputs(3951) <= not(layer0_outputs(12223));
    outputs(3952) <= not(layer0_outputs(10024));
    outputs(3953) <= not((layer0_outputs(4461)) or (layer0_outputs(5978)));
    outputs(3954) <= (layer0_outputs(7320)) xor (layer0_outputs(1841));
    outputs(3955) <= (layer0_outputs(9665)) and not (layer0_outputs(3222));
    outputs(3956) <= layer0_outputs(11870);
    outputs(3957) <= (layer0_outputs(5536)) and not (layer0_outputs(6905));
    outputs(3958) <= not((layer0_outputs(2756)) or (layer0_outputs(955)));
    outputs(3959) <= not(layer0_outputs(1529));
    outputs(3960) <= layer0_outputs(5381);
    outputs(3961) <= layer0_outputs(7339);
    outputs(3962) <= (layer0_outputs(31)) or (layer0_outputs(2737));
    outputs(3963) <= not(layer0_outputs(4838));
    outputs(3964) <= not((layer0_outputs(2784)) or (layer0_outputs(3175)));
    outputs(3965) <= not(layer0_outputs(11321)) or (layer0_outputs(10061));
    outputs(3966) <= not(layer0_outputs(10475));
    outputs(3967) <= not((layer0_outputs(8582)) xor (layer0_outputs(2850)));
    outputs(3968) <= not(layer0_outputs(10214)) or (layer0_outputs(2639));
    outputs(3969) <= not(layer0_outputs(4368));
    outputs(3970) <= (layer0_outputs(3121)) xor (layer0_outputs(4396));
    outputs(3971) <= (layer0_outputs(1897)) or (layer0_outputs(6711));
    outputs(3972) <= not((layer0_outputs(8526)) and (layer0_outputs(10438)));
    outputs(3973) <= layer0_outputs(1959);
    outputs(3974) <= (layer0_outputs(1983)) xor (layer0_outputs(840));
    outputs(3975) <= not(layer0_outputs(7223));
    outputs(3976) <= not(layer0_outputs(1413)) or (layer0_outputs(11941));
    outputs(3977) <= not(layer0_outputs(9126));
    outputs(3978) <= not(layer0_outputs(1969));
    outputs(3979) <= not((layer0_outputs(5775)) xor (layer0_outputs(12699)));
    outputs(3980) <= not(layer0_outputs(1910));
    outputs(3981) <= layer0_outputs(12078);
    outputs(3982) <= not((layer0_outputs(6220)) and (layer0_outputs(2806)));
    outputs(3983) <= (layer0_outputs(8723)) and (layer0_outputs(3249));
    outputs(3984) <= (layer0_outputs(2731)) and not (layer0_outputs(5822));
    outputs(3985) <= (layer0_outputs(364)) or (layer0_outputs(1427));
    outputs(3986) <= (layer0_outputs(3746)) xor (layer0_outputs(9335));
    outputs(3987) <= not(layer0_outputs(3038));
    outputs(3988) <= layer0_outputs(4749);
    outputs(3989) <= (layer0_outputs(737)) or (layer0_outputs(12339));
    outputs(3990) <= (layer0_outputs(10251)) and not (layer0_outputs(5692));
    outputs(3991) <= layer0_outputs(12037);
    outputs(3992) <= not((layer0_outputs(6289)) xor (layer0_outputs(8943)));
    outputs(3993) <= not(layer0_outputs(11347)) or (layer0_outputs(6737));
    outputs(3994) <= (layer0_outputs(6119)) and not (layer0_outputs(1092));
    outputs(3995) <= layer0_outputs(8473);
    outputs(3996) <= (layer0_outputs(5623)) and not (layer0_outputs(8443));
    outputs(3997) <= not((layer0_outputs(6050)) or (layer0_outputs(1758)));
    outputs(3998) <= not(layer0_outputs(9648)) or (layer0_outputs(6939));
    outputs(3999) <= not((layer0_outputs(2996)) xor (layer0_outputs(5144)));
    outputs(4000) <= not(layer0_outputs(11794));
    outputs(4001) <= layer0_outputs(9244);
    outputs(4002) <= (layer0_outputs(12626)) and not (layer0_outputs(2740));
    outputs(4003) <= not(layer0_outputs(3813));
    outputs(4004) <= (layer0_outputs(10239)) and (layer0_outputs(9742));
    outputs(4005) <= not((layer0_outputs(2759)) or (layer0_outputs(2636)));
    outputs(4006) <= (layer0_outputs(10642)) and not (layer0_outputs(9224));
    outputs(4007) <= not(layer0_outputs(12578));
    outputs(4008) <= (layer0_outputs(8938)) and not (layer0_outputs(2755));
    outputs(4009) <= not(layer0_outputs(5179));
    outputs(4010) <= not(layer0_outputs(307));
    outputs(4011) <= not((layer0_outputs(4267)) xor (layer0_outputs(4881)));
    outputs(4012) <= not((layer0_outputs(6874)) or (layer0_outputs(5060)));
    outputs(4013) <= not((layer0_outputs(6647)) and (layer0_outputs(410)));
    outputs(4014) <= (layer0_outputs(2663)) or (layer0_outputs(3381));
    outputs(4015) <= not((layer0_outputs(3855)) or (layer0_outputs(2939)));
    outputs(4016) <= not((layer0_outputs(8506)) and (layer0_outputs(7449)));
    outputs(4017) <= layer0_outputs(10288);
    outputs(4018) <= not(layer0_outputs(7583));
    outputs(4019) <= layer0_outputs(11108);
    outputs(4020) <= layer0_outputs(10424);
    outputs(4021) <= not((layer0_outputs(8521)) and (layer0_outputs(11411)));
    outputs(4022) <= layer0_outputs(7574);
    outputs(4023) <= not(layer0_outputs(5153));
    outputs(4024) <= (layer0_outputs(408)) and not (layer0_outputs(12159));
    outputs(4025) <= not((layer0_outputs(6791)) xor (layer0_outputs(4010)));
    outputs(4026) <= layer0_outputs(529);
    outputs(4027) <= (layer0_outputs(1222)) and not (layer0_outputs(2637));
    outputs(4028) <= not((layer0_outputs(4796)) or (layer0_outputs(2163)));
    outputs(4029) <= layer0_outputs(12629);
    outputs(4030) <= not((layer0_outputs(2093)) xor (layer0_outputs(550)));
    outputs(4031) <= not((layer0_outputs(11152)) or (layer0_outputs(120)));
    outputs(4032) <= not((layer0_outputs(1760)) xor (layer0_outputs(2312)));
    outputs(4033) <= not((layer0_outputs(12062)) xor (layer0_outputs(6544)));
    outputs(4034) <= not((layer0_outputs(6140)) xor (layer0_outputs(10393)));
    outputs(4035) <= (layer0_outputs(10790)) or (layer0_outputs(11252));
    outputs(4036) <= (layer0_outputs(6520)) and not (layer0_outputs(5120));
    outputs(4037) <= not(layer0_outputs(11968));
    outputs(4038) <= not((layer0_outputs(5711)) or (layer0_outputs(5898)));
    outputs(4039) <= layer0_outputs(7611);
    outputs(4040) <= (layer0_outputs(9181)) and (layer0_outputs(11260));
    outputs(4041) <= not(layer0_outputs(4880));
    outputs(4042) <= not(layer0_outputs(1826));
    outputs(4043) <= layer0_outputs(7991);
    outputs(4044) <= not(layer0_outputs(8676)) or (layer0_outputs(10676));
    outputs(4045) <= layer0_outputs(12554);
    outputs(4046) <= layer0_outputs(8611);
    outputs(4047) <= not(layer0_outputs(1262));
    outputs(4048) <= not(layer0_outputs(4823));
    outputs(4049) <= layer0_outputs(3308);
    outputs(4050) <= not(layer0_outputs(5853)) or (layer0_outputs(10461));
    outputs(4051) <= not((layer0_outputs(7685)) xor (layer0_outputs(7501)));
    outputs(4052) <= not(layer0_outputs(10654));
    outputs(4053) <= (layer0_outputs(10471)) xor (layer0_outputs(10148));
    outputs(4054) <= (layer0_outputs(1085)) xor (layer0_outputs(6275));
    outputs(4055) <= not(layer0_outputs(2822));
    outputs(4056) <= not(layer0_outputs(10837));
    outputs(4057) <= (layer0_outputs(9264)) and not (layer0_outputs(10003));
    outputs(4058) <= layer0_outputs(12147);
    outputs(4059) <= '0';
    outputs(4060) <= layer0_outputs(5325);
    outputs(4061) <= not((layer0_outputs(10087)) xor (layer0_outputs(1135)));
    outputs(4062) <= not((layer0_outputs(12577)) and (layer0_outputs(11077)));
    outputs(4063) <= not(layer0_outputs(474)) or (layer0_outputs(6813));
    outputs(4064) <= not(layer0_outputs(12127));
    outputs(4065) <= (layer0_outputs(11740)) and not (layer0_outputs(1151));
    outputs(4066) <= (layer0_outputs(11589)) and not (layer0_outputs(7456));
    outputs(4067) <= not((layer0_outputs(4148)) and (layer0_outputs(3100)));
    outputs(4068) <= layer0_outputs(1622);
    outputs(4069) <= (layer0_outputs(1266)) and not (layer0_outputs(11222));
    outputs(4070) <= not(layer0_outputs(6564));
    outputs(4071) <= not((layer0_outputs(5030)) xor (layer0_outputs(10359)));
    outputs(4072) <= not((layer0_outputs(8678)) and (layer0_outputs(1226)));
    outputs(4073) <= (layer0_outputs(3640)) and (layer0_outputs(5445));
    outputs(4074) <= (layer0_outputs(5093)) and (layer0_outputs(227));
    outputs(4075) <= not(layer0_outputs(12738)) or (layer0_outputs(2792));
    outputs(4076) <= layer0_outputs(7787);
    outputs(4077) <= (layer0_outputs(5036)) and not (layer0_outputs(8336));
    outputs(4078) <= (layer0_outputs(10981)) and (layer0_outputs(7584));
    outputs(4079) <= layer0_outputs(5290);
    outputs(4080) <= not(layer0_outputs(2856));
    outputs(4081) <= not(layer0_outputs(2004));
    outputs(4082) <= (layer0_outputs(3379)) xor (layer0_outputs(9477));
    outputs(4083) <= (layer0_outputs(3478)) xor (layer0_outputs(3168));
    outputs(4084) <= (layer0_outputs(3583)) and (layer0_outputs(7850));
    outputs(4085) <= not(layer0_outputs(6713));
    outputs(4086) <= not(layer0_outputs(4788)) or (layer0_outputs(6918));
    outputs(4087) <= not(layer0_outputs(302)) or (layer0_outputs(397));
    outputs(4088) <= not((layer0_outputs(6720)) xor (layer0_outputs(12152)));
    outputs(4089) <= layer0_outputs(2240);
    outputs(4090) <= not((layer0_outputs(12022)) or (layer0_outputs(3171)));
    outputs(4091) <= not(layer0_outputs(861));
    outputs(4092) <= not((layer0_outputs(5951)) or (layer0_outputs(10159)));
    outputs(4093) <= not((layer0_outputs(6181)) xor (layer0_outputs(10185)));
    outputs(4094) <= (layer0_outputs(1472)) or (layer0_outputs(1688));
    outputs(4095) <= (layer0_outputs(11248)) and not (layer0_outputs(6154));
    outputs(4096) <= not(layer0_outputs(8718));
    outputs(4097) <= (layer0_outputs(8857)) and (layer0_outputs(5286));
    outputs(4098) <= not(layer0_outputs(6660));
    outputs(4099) <= layer0_outputs(11595);
    outputs(4100) <= layer0_outputs(8641);
    outputs(4101) <= layer0_outputs(6321);
    outputs(4102) <= layer0_outputs(466);
    outputs(4103) <= not(layer0_outputs(472));
    outputs(4104) <= not((layer0_outputs(10544)) or (layer0_outputs(846)));
    outputs(4105) <= not((layer0_outputs(4036)) xor (layer0_outputs(8939)));
    outputs(4106) <= (layer0_outputs(8551)) and not (layer0_outputs(4250));
    outputs(4107) <= not((layer0_outputs(6469)) xor (layer0_outputs(2016)));
    outputs(4108) <= not(layer0_outputs(2110));
    outputs(4109) <= layer0_outputs(493);
    outputs(4110) <= layer0_outputs(5874);
    outputs(4111) <= (layer0_outputs(2120)) and not (layer0_outputs(8301));
    outputs(4112) <= not((layer0_outputs(4477)) or (layer0_outputs(8297)));
    outputs(4113) <= (layer0_outputs(3915)) or (layer0_outputs(10651));
    outputs(4114) <= layer0_outputs(5649);
    outputs(4115) <= (layer0_outputs(6133)) xor (layer0_outputs(7896));
    outputs(4116) <= not(layer0_outputs(8682));
    outputs(4117) <= not((layer0_outputs(3886)) xor (layer0_outputs(9324)));
    outputs(4118) <= (layer0_outputs(11073)) and not (layer0_outputs(10741));
    outputs(4119) <= not((layer0_outputs(3279)) and (layer0_outputs(412)));
    outputs(4120) <= not(layer0_outputs(2050));
    outputs(4121) <= not(layer0_outputs(12029));
    outputs(4122) <= layer0_outputs(5119);
    outputs(4123) <= (layer0_outputs(3259)) and not (layer0_outputs(963));
    outputs(4124) <= (layer0_outputs(311)) and not (layer0_outputs(4462));
    outputs(4125) <= not(layer0_outputs(11559));
    outputs(4126) <= not((layer0_outputs(7556)) and (layer0_outputs(10003)));
    outputs(4127) <= (layer0_outputs(156)) or (layer0_outputs(3616));
    outputs(4128) <= not((layer0_outputs(9414)) xor (layer0_outputs(9842)));
    outputs(4129) <= not(layer0_outputs(1841));
    outputs(4130) <= layer0_outputs(6615);
    outputs(4131) <= layer0_outputs(6588);
    outputs(4132) <= (layer0_outputs(11759)) and not (layer0_outputs(4307));
    outputs(4133) <= not(layer0_outputs(7186));
    outputs(4134) <= not(layer0_outputs(6477));
    outputs(4135) <= not((layer0_outputs(5305)) or (layer0_outputs(4140)));
    outputs(4136) <= layer0_outputs(9560);
    outputs(4137) <= not((layer0_outputs(10228)) and (layer0_outputs(12471)));
    outputs(4138) <= not((layer0_outputs(630)) and (layer0_outputs(2335)));
    outputs(4139) <= (layer0_outputs(1602)) and (layer0_outputs(10450));
    outputs(4140) <= (layer0_outputs(5452)) and (layer0_outputs(6078));
    outputs(4141) <= not((layer0_outputs(1762)) or (layer0_outputs(4589)));
    outputs(4142) <= layer0_outputs(5694);
    outputs(4143) <= not(layer0_outputs(11425));
    outputs(4144) <= (layer0_outputs(4329)) and (layer0_outputs(1302));
    outputs(4145) <= not((layer0_outputs(10530)) or (layer0_outputs(4793)));
    outputs(4146) <= (layer0_outputs(10809)) xor (layer0_outputs(7027));
    outputs(4147) <= not(layer0_outputs(3514));
    outputs(4148) <= not((layer0_outputs(1518)) and (layer0_outputs(3418)));
    outputs(4149) <= not(layer0_outputs(4594)) or (layer0_outputs(11755));
    outputs(4150) <= (layer0_outputs(7144)) and not (layer0_outputs(8386));
    outputs(4151) <= not((layer0_outputs(4696)) xor (layer0_outputs(5630)));
    outputs(4152) <= layer0_outputs(11861);
    outputs(4153) <= not((layer0_outputs(9305)) and (layer0_outputs(5360)));
    outputs(4154) <= not(layer0_outputs(5024)) or (layer0_outputs(5707));
    outputs(4155) <= not(layer0_outputs(6231)) or (layer0_outputs(9198));
    outputs(4156) <= not((layer0_outputs(9655)) xor (layer0_outputs(1564)));
    outputs(4157) <= not(layer0_outputs(6009)) or (layer0_outputs(2176));
    outputs(4158) <= not((layer0_outputs(6235)) or (layer0_outputs(11284)));
    outputs(4159) <= not((layer0_outputs(6970)) xor (layer0_outputs(8969)));
    outputs(4160) <= (layer0_outputs(9770)) and not (layer0_outputs(12330));
    outputs(4161) <= not(layer0_outputs(515));
    outputs(4162) <= layer0_outputs(12010);
    outputs(4163) <= (layer0_outputs(3311)) or (layer0_outputs(6377));
    outputs(4164) <= not(layer0_outputs(7544));
    outputs(4165) <= not((layer0_outputs(12410)) and (layer0_outputs(4746)));
    outputs(4166) <= layer0_outputs(10452);
    outputs(4167) <= not((layer0_outputs(9802)) or (layer0_outputs(8817)));
    outputs(4168) <= layer0_outputs(9268);
    outputs(4169) <= not(layer0_outputs(7782)) or (layer0_outputs(12293));
    outputs(4170) <= layer0_outputs(8954);
    outputs(4171) <= not((layer0_outputs(3999)) xor (layer0_outputs(6415)));
    outputs(4172) <= not((layer0_outputs(5309)) xor (layer0_outputs(8961)));
    outputs(4173) <= (layer0_outputs(2243)) or (layer0_outputs(8242));
    outputs(4174) <= not(layer0_outputs(9069));
    outputs(4175) <= (layer0_outputs(7175)) and (layer0_outputs(7306));
    outputs(4176) <= not(layer0_outputs(6531));
    outputs(4177) <= not((layer0_outputs(5922)) xor (layer0_outputs(6051)));
    outputs(4178) <= layer0_outputs(399);
    outputs(4179) <= (layer0_outputs(3052)) and not (layer0_outputs(1010));
    outputs(4180) <= not(layer0_outputs(12252));
    outputs(4181) <= not((layer0_outputs(12732)) and (layer0_outputs(9803)));
    outputs(4182) <= (layer0_outputs(10727)) and not (layer0_outputs(6193));
    outputs(4183) <= not(layer0_outputs(8133));
    outputs(4184) <= layer0_outputs(5849);
    outputs(4185) <= not(layer0_outputs(10545));
    outputs(4186) <= not(layer0_outputs(757)) or (layer0_outputs(8405));
    outputs(4187) <= not((layer0_outputs(332)) or (layer0_outputs(8556)));
    outputs(4188) <= not((layer0_outputs(12279)) xor (layer0_outputs(6634)));
    outputs(4189) <= (layer0_outputs(6264)) xor (layer0_outputs(2320));
    outputs(4190) <= layer0_outputs(3808);
    outputs(4191) <= not(layer0_outputs(882));
    outputs(4192) <= layer0_outputs(9858);
    outputs(4193) <= layer0_outputs(2480);
    outputs(4194) <= not(layer0_outputs(3725)) or (layer0_outputs(1060));
    outputs(4195) <= not(layer0_outputs(9138));
    outputs(4196) <= layer0_outputs(6439);
    outputs(4197) <= not(layer0_outputs(8609));
    outputs(4198) <= layer0_outputs(11390);
    outputs(4199) <= layer0_outputs(8037);
    outputs(4200) <= (layer0_outputs(5520)) or (layer0_outputs(9756));
    outputs(4201) <= (layer0_outputs(6013)) xor (layer0_outputs(2348));
    outputs(4202) <= not(layer0_outputs(5027));
    outputs(4203) <= not(layer0_outputs(10241));
    outputs(4204) <= layer0_outputs(4281);
    outputs(4205) <= not(layer0_outputs(195));
    outputs(4206) <= not(layer0_outputs(5178));
    outputs(4207) <= (layer0_outputs(6427)) xor (layer0_outputs(685));
    outputs(4208) <= (layer0_outputs(11446)) xor (layer0_outputs(2514));
    outputs(4209) <= layer0_outputs(9720);
    outputs(4210) <= layer0_outputs(8190);
    outputs(4211) <= not((layer0_outputs(5704)) xor (layer0_outputs(12208)));
    outputs(4212) <= (layer0_outputs(4453)) xor (layer0_outputs(12658));
    outputs(4213) <= layer0_outputs(11232);
    outputs(4214) <= not((layer0_outputs(8162)) or (layer0_outputs(10303)));
    outputs(4215) <= (layer0_outputs(11731)) and not (layer0_outputs(6135));
    outputs(4216) <= layer0_outputs(2292);
    outputs(4217) <= not(layer0_outputs(8745));
    outputs(4218) <= layer0_outputs(9297);
    outputs(4219) <= not(layer0_outputs(6892));
    outputs(4220) <= (layer0_outputs(6355)) and not (layer0_outputs(1298));
    outputs(4221) <= layer0_outputs(4631);
    outputs(4222) <= not(layer0_outputs(463));
    outputs(4223) <= not(layer0_outputs(8081));
    outputs(4224) <= (layer0_outputs(2494)) xor (layer0_outputs(1814));
    outputs(4225) <= (layer0_outputs(3446)) xor (layer0_outputs(12142));
    outputs(4226) <= layer0_outputs(7891);
    outputs(4227) <= layer0_outputs(8282);
    outputs(4228) <= (layer0_outputs(4884)) and not (layer0_outputs(9347));
    outputs(4229) <= not((layer0_outputs(2998)) xor (layer0_outputs(11280)));
    outputs(4230) <= (layer0_outputs(5703)) xor (layer0_outputs(3362));
    outputs(4231) <= layer0_outputs(3647);
    outputs(4232) <= not(layer0_outputs(4897)) or (layer0_outputs(7433));
    outputs(4233) <= (layer0_outputs(4151)) and not (layer0_outputs(9233));
    outputs(4234) <= '1';
    outputs(4235) <= (layer0_outputs(6548)) xor (layer0_outputs(11569));
    outputs(4236) <= (layer0_outputs(6660)) xor (layer0_outputs(6760));
    outputs(4237) <= not((layer0_outputs(10596)) or (layer0_outputs(3826)));
    outputs(4238) <= (layer0_outputs(11463)) xor (layer0_outputs(9496));
    outputs(4239) <= not(layer0_outputs(11064)) or (layer0_outputs(3676));
    outputs(4240) <= (layer0_outputs(12253)) and not (layer0_outputs(5252));
    outputs(4241) <= layer0_outputs(1823);
    outputs(4242) <= (layer0_outputs(3438)) and not (layer0_outputs(6440));
    outputs(4243) <= not(layer0_outputs(12110));
    outputs(4244) <= layer0_outputs(10862);
    outputs(4245) <= layer0_outputs(8619);
    outputs(4246) <= layer0_outputs(2667);
    outputs(4247) <= (layer0_outputs(7773)) and (layer0_outputs(12249));
    outputs(4248) <= layer0_outputs(2155);
    outputs(4249) <= not((layer0_outputs(948)) and (layer0_outputs(2325)));
    outputs(4250) <= not(layer0_outputs(9079));
    outputs(4251) <= layer0_outputs(3979);
    outputs(4252) <= (layer0_outputs(5901)) xor (layer0_outputs(11135));
    outputs(4253) <= layer0_outputs(33);
    outputs(4254) <= (layer0_outputs(11070)) or (layer0_outputs(3839));
    outputs(4255) <= layer0_outputs(5455);
    outputs(4256) <= not((layer0_outputs(10499)) xor (layer0_outputs(9451)));
    outputs(4257) <= not(layer0_outputs(1121)) or (layer0_outputs(10832));
    outputs(4258) <= not((layer0_outputs(11790)) and (layer0_outputs(8647)));
    outputs(4259) <= not((layer0_outputs(3866)) xor (layer0_outputs(10088)));
    outputs(4260) <= not(layer0_outputs(7058));
    outputs(4261) <= not(layer0_outputs(4620));
    outputs(4262) <= (layer0_outputs(5652)) xor (layer0_outputs(12430));
    outputs(4263) <= layer0_outputs(12700);
    outputs(4264) <= not(layer0_outputs(3675));
    outputs(4265) <= (layer0_outputs(11231)) and not (layer0_outputs(9899));
    outputs(4266) <= not((layer0_outputs(2983)) or (layer0_outputs(1545)));
    outputs(4267) <= (layer0_outputs(1279)) and not (layer0_outputs(2082));
    outputs(4268) <= layer0_outputs(2598);
    outputs(4269) <= not(layer0_outputs(10520));
    outputs(4270) <= (layer0_outputs(5714)) and (layer0_outputs(3221));
    outputs(4271) <= not(layer0_outputs(11553));
    outputs(4272) <= not(layer0_outputs(5691));
    outputs(4273) <= (layer0_outputs(4275)) and (layer0_outputs(4167));
    outputs(4274) <= not(layer0_outputs(7157));
    outputs(4275) <= not(layer0_outputs(10345));
    outputs(4276) <= layer0_outputs(10310);
    outputs(4277) <= layer0_outputs(9967);
    outputs(4278) <= not(layer0_outputs(9361));
    outputs(4279) <= not((layer0_outputs(12073)) or (layer0_outputs(7742)));
    outputs(4280) <= not((layer0_outputs(9599)) or (layer0_outputs(4817)));
    outputs(4281) <= layer0_outputs(12004);
    outputs(4282) <= (layer0_outputs(363)) and (layer0_outputs(7873));
    outputs(4283) <= layer0_outputs(1181);
    outputs(4284) <= not(layer0_outputs(9903));
    outputs(4285) <= not(layer0_outputs(11286));
    outputs(4286) <= not((layer0_outputs(2442)) xor (layer0_outputs(913)));
    outputs(4287) <= not((layer0_outputs(7969)) and (layer0_outputs(2542)));
    outputs(4288) <= (layer0_outputs(9563)) xor (layer0_outputs(887));
    outputs(4289) <= layer0_outputs(3821);
    outputs(4290) <= (layer0_outputs(4058)) or (layer0_outputs(11305));
    outputs(4291) <= not((layer0_outputs(9955)) xor (layer0_outputs(9911)));
    outputs(4292) <= not((layer0_outputs(381)) or (layer0_outputs(11557)));
    outputs(4293) <= not((layer0_outputs(6776)) xor (layer0_outputs(11983)));
    outputs(4294) <= (layer0_outputs(11284)) or (layer0_outputs(4885));
    outputs(4295) <= not((layer0_outputs(12745)) and (layer0_outputs(4672)));
    outputs(4296) <= not((layer0_outputs(9210)) and (layer0_outputs(4176)));
    outputs(4297) <= not(layer0_outputs(4970));
    outputs(4298) <= not((layer0_outputs(11309)) or (layer0_outputs(2232)));
    outputs(4299) <= (layer0_outputs(8221)) xor (layer0_outputs(4479));
    outputs(4300) <= not(layer0_outputs(6650)) or (layer0_outputs(9392));
    outputs(4301) <= (layer0_outputs(3350)) and not (layer0_outputs(1244));
    outputs(4302) <= (layer0_outputs(7888)) and not (layer0_outputs(11933));
    outputs(4303) <= (layer0_outputs(12524)) xor (layer0_outputs(2978));
    outputs(4304) <= (layer0_outputs(3711)) xor (layer0_outputs(3025));
    outputs(4305) <= (layer0_outputs(10062)) and not (layer0_outputs(8800));
    outputs(4306) <= not(layer0_outputs(9021));
    outputs(4307) <= (layer0_outputs(12321)) and not (layer0_outputs(10526));
    outputs(4308) <= layer0_outputs(1565);
    outputs(4309) <= (layer0_outputs(3296)) and (layer0_outputs(7692));
    outputs(4310) <= not(layer0_outputs(2803));
    outputs(4311) <= layer0_outputs(3245);
    outputs(4312) <= (layer0_outputs(11644)) and (layer0_outputs(2219));
    outputs(4313) <= not(layer0_outputs(6258));
    outputs(4314) <= (layer0_outputs(10423)) and not (layer0_outputs(5937));
    outputs(4315) <= '0';
    outputs(4316) <= not(layer0_outputs(10679));
    outputs(4317) <= layer0_outputs(2144);
    outputs(4318) <= layer0_outputs(8633);
    outputs(4319) <= layer0_outputs(12194);
    outputs(4320) <= not((layer0_outputs(5963)) xor (layer0_outputs(4951)));
    outputs(4321) <= (layer0_outputs(1283)) and not (layer0_outputs(10675));
    outputs(4322) <= layer0_outputs(4978);
    outputs(4323) <= (layer0_outputs(2900)) and not (layer0_outputs(1122));
    outputs(4324) <= (layer0_outputs(5295)) xor (layer0_outputs(6284));
    outputs(4325) <= not(layer0_outputs(3864));
    outputs(4326) <= not(layer0_outputs(2619)) or (layer0_outputs(10912));
    outputs(4327) <= (layer0_outputs(832)) and not (layer0_outputs(8936));
    outputs(4328) <= not(layer0_outputs(5716));
    outputs(4329) <= layer0_outputs(1474);
    outputs(4330) <= not((layer0_outputs(7904)) or (layer0_outputs(5993)));
    outputs(4331) <= not(layer0_outputs(1393)) or (layer0_outputs(9658));
    outputs(4332) <= layer0_outputs(12405);
    outputs(4333) <= layer0_outputs(5188);
    outputs(4334) <= not(layer0_outputs(2575));
    outputs(4335) <= not(layer0_outputs(7294));
    outputs(4336) <= layer0_outputs(2045);
    outputs(4337) <= layer0_outputs(7413);
    outputs(4338) <= not((layer0_outputs(8428)) or (layer0_outputs(9779)));
    outputs(4339) <= not(layer0_outputs(6928));
    outputs(4340) <= layer0_outputs(6613);
    outputs(4341) <= not(layer0_outputs(2423));
    outputs(4342) <= layer0_outputs(6612);
    outputs(4343) <= not(layer0_outputs(1587));
    outputs(4344) <= not(layer0_outputs(1220));
    outputs(4345) <= not(layer0_outputs(11313));
    outputs(4346) <= not(layer0_outputs(5983));
    outputs(4347) <= (layer0_outputs(10455)) or (layer0_outputs(9595));
    outputs(4348) <= not(layer0_outputs(6508)) or (layer0_outputs(2080));
    outputs(4349) <= not(layer0_outputs(2297));
    outputs(4350) <= not((layer0_outputs(5277)) xor (layer0_outputs(7453)));
    outputs(4351) <= not(layer0_outputs(4699));
    outputs(4352) <= not((layer0_outputs(7758)) or (layer0_outputs(6089)));
    outputs(4353) <= layer0_outputs(6796);
    outputs(4354) <= not(layer0_outputs(5681));
    outputs(4355) <= not(layer0_outputs(4863));
    outputs(4356) <= layer0_outputs(1349);
    outputs(4357) <= (layer0_outputs(10881)) xor (layer0_outputs(5274));
    outputs(4358) <= layer0_outputs(11902);
    outputs(4359) <= layer0_outputs(1430);
    outputs(4360) <= layer0_outputs(2333);
    outputs(4361) <= not(layer0_outputs(241));
    outputs(4362) <= not((layer0_outputs(1828)) xor (layer0_outputs(4773)));
    outputs(4363) <= (layer0_outputs(1846)) xor (layer0_outputs(5249));
    outputs(4364) <= layer0_outputs(4561);
    outputs(4365) <= not((layer0_outputs(4913)) or (layer0_outputs(6244)));
    outputs(4366) <= (layer0_outputs(876)) xor (layer0_outputs(444));
    outputs(4367) <= not((layer0_outputs(6910)) xor (layer0_outputs(3947)));
    outputs(4368) <= not(layer0_outputs(6313));
    outputs(4369) <= layer0_outputs(11206);
    outputs(4370) <= (layer0_outputs(699)) and not (layer0_outputs(4139));
    outputs(4371) <= layer0_outputs(2159);
    outputs(4372) <= layer0_outputs(8956);
    outputs(4373) <= not(layer0_outputs(10525));
    outputs(4374) <= (layer0_outputs(459)) and not (layer0_outputs(12068));
    outputs(4375) <= (layer0_outputs(2275)) and (layer0_outputs(3313));
    outputs(4376) <= (layer0_outputs(2758)) xor (layer0_outputs(5341));
    outputs(4377) <= layer0_outputs(11639);
    outputs(4378) <= not((layer0_outputs(5050)) xor (layer0_outputs(7078)));
    outputs(4379) <= not((layer0_outputs(10997)) xor (layer0_outputs(4304)));
    outputs(4380) <= (layer0_outputs(1109)) and not (layer0_outputs(4979));
    outputs(4381) <= layer0_outputs(12338);
    outputs(4382) <= (layer0_outputs(4147)) xor (layer0_outputs(1389));
    outputs(4383) <= not(layer0_outputs(5257));
    outputs(4384) <= not(layer0_outputs(3581));
    outputs(4385) <= (layer0_outputs(4103)) xor (layer0_outputs(12249));
    outputs(4386) <= not(layer0_outputs(9631));
    outputs(4387) <= layer0_outputs(11883);
    outputs(4388) <= not(layer0_outputs(9385));
    outputs(4389) <= (layer0_outputs(8079)) or (layer0_outputs(6816));
    outputs(4390) <= layer0_outputs(11621);
    outputs(4391) <= not(layer0_outputs(1409));
    outputs(4392) <= not(layer0_outputs(10420));
    outputs(4393) <= not(layer0_outputs(8758));
    outputs(4394) <= layer0_outputs(1602);
    outputs(4395) <= not(layer0_outputs(177)) or (layer0_outputs(12051));
    outputs(4396) <= layer0_outputs(4255);
    outputs(4397) <= layer0_outputs(3613);
    outputs(4398) <= not(layer0_outputs(12303));
    outputs(4399) <= not(layer0_outputs(1632));
    outputs(4400) <= not(layer0_outputs(4305));
    outputs(4401) <= not(layer0_outputs(8729));
    outputs(4402) <= (layer0_outputs(6984)) xor (layer0_outputs(9418));
    outputs(4403) <= layer0_outputs(4407);
    outputs(4404) <= (layer0_outputs(5391)) or (layer0_outputs(2503));
    outputs(4405) <= not(layer0_outputs(11957));
    outputs(4406) <= not((layer0_outputs(6768)) or (layer0_outputs(9542)));
    outputs(4407) <= not(layer0_outputs(7389)) or (layer0_outputs(1859));
    outputs(4408) <= not((layer0_outputs(1230)) xor (layer0_outputs(9426)));
    outputs(4409) <= not((layer0_outputs(11150)) or (layer0_outputs(10136)));
    outputs(4410) <= (layer0_outputs(3448)) xor (layer0_outputs(698));
    outputs(4411) <= layer0_outputs(6481);
    outputs(4412) <= layer0_outputs(9701);
    outputs(4413) <= layer0_outputs(9080);
    outputs(4414) <= not((layer0_outputs(11596)) or (layer0_outputs(2749)));
    outputs(4415) <= not((layer0_outputs(1847)) xor (layer0_outputs(3413)));
    outputs(4416) <= not(layer0_outputs(1851));
    outputs(4417) <= layer0_outputs(11482);
    outputs(4418) <= (layer0_outputs(12342)) and not (layer0_outputs(5773));
    outputs(4419) <= not(layer0_outputs(7478)) or (layer0_outputs(3283));
    outputs(4420) <= (layer0_outputs(7994)) and not (layer0_outputs(10752));
    outputs(4421) <= not((layer0_outputs(4143)) and (layer0_outputs(7829)));
    outputs(4422) <= not(layer0_outputs(10339));
    outputs(4423) <= (layer0_outputs(6669)) xor (layer0_outputs(2064));
    outputs(4424) <= (layer0_outputs(5374)) and not (layer0_outputs(6968));
    outputs(4425) <= not((layer0_outputs(9219)) or (layer0_outputs(9906)));
    outputs(4426) <= not(layer0_outputs(7901)) or (layer0_outputs(12449));
    outputs(4427) <= not(layer0_outputs(10395));
    outputs(4428) <= (layer0_outputs(12058)) xor (layer0_outputs(844));
    outputs(4429) <= not((layer0_outputs(214)) xor (layer0_outputs(7328)));
    outputs(4430) <= not(layer0_outputs(4807)) or (layer0_outputs(12346));
    outputs(4431) <= not(layer0_outputs(1559)) or (layer0_outputs(7005));
    outputs(4432) <= (layer0_outputs(10640)) and not (layer0_outputs(4007));
    outputs(4433) <= layer0_outputs(8454);
    outputs(4434) <= layer0_outputs(3450);
    outputs(4435) <= not((layer0_outputs(418)) or (layer0_outputs(5319)));
    outputs(4436) <= (layer0_outputs(8765)) and not (layer0_outputs(8869));
    outputs(4437) <= (layer0_outputs(9475)) and not (layer0_outputs(9765));
    outputs(4438) <= (layer0_outputs(4231)) xor (layer0_outputs(6757));
    outputs(4439) <= not((layer0_outputs(7967)) or (layer0_outputs(1904)));
    outputs(4440) <= not(layer0_outputs(769));
    outputs(4441) <= (layer0_outputs(2526)) and (layer0_outputs(11567));
    outputs(4442) <= (layer0_outputs(1447)) or (layer0_outputs(9322));
    outputs(4443) <= layer0_outputs(3560);
    outputs(4444) <= (layer0_outputs(1658)) xor (layer0_outputs(8416));
    outputs(4445) <= (layer0_outputs(3007)) xor (layer0_outputs(12747));
    outputs(4446) <= not(layer0_outputs(4193));
    outputs(4447) <= (layer0_outputs(8664)) and not (layer0_outputs(3554));
    outputs(4448) <= layer0_outputs(4814);
    outputs(4449) <= not(layer0_outputs(8863));
    outputs(4450) <= (layer0_outputs(1739)) and not (layer0_outputs(2262));
    outputs(4451) <= not(layer0_outputs(669));
    outputs(4452) <= not(layer0_outputs(5174));
    outputs(4453) <= (layer0_outputs(8783)) xor (layer0_outputs(8260));
    outputs(4454) <= (layer0_outputs(12272)) xor (layer0_outputs(2236));
    outputs(4455) <= layer0_outputs(5792);
    outputs(4456) <= not((layer0_outputs(8123)) xor (layer0_outputs(10999)));
    outputs(4457) <= not(layer0_outputs(1803));
    outputs(4458) <= layer0_outputs(5566);
    outputs(4459) <= layer0_outputs(10565);
    outputs(4460) <= (layer0_outputs(1825)) xor (layer0_outputs(3372));
    outputs(4461) <= not((layer0_outputs(9876)) xor (layer0_outputs(7176)));
    outputs(4462) <= (layer0_outputs(10320)) xor (layer0_outputs(6441));
    outputs(4463) <= layer0_outputs(3207);
    outputs(4464) <= not(layer0_outputs(2516)) or (layer0_outputs(4872));
    outputs(4465) <= not(layer0_outputs(4818));
    outputs(4466) <= layer0_outputs(10906);
    outputs(4467) <= layer0_outputs(6646);
    outputs(4468) <= not((layer0_outputs(11895)) or (layer0_outputs(7187)));
    outputs(4469) <= layer0_outputs(11367);
    outputs(4470) <= not(layer0_outputs(859)) or (layer0_outputs(1661));
    outputs(4471) <= not(layer0_outputs(12159));
    outputs(4472) <= not(layer0_outputs(648)) or (layer0_outputs(845));
    outputs(4473) <= (layer0_outputs(5169)) xor (layer0_outputs(12277));
    outputs(4474) <= layer0_outputs(7684);
    outputs(4475) <= not((layer0_outputs(11086)) and (layer0_outputs(10799)));
    outputs(4476) <= not(layer0_outputs(4668));
    outputs(4477) <= not((layer0_outputs(814)) xor (layer0_outputs(6542)));
    outputs(4478) <= layer0_outputs(10968);
    outputs(4479) <= not(layer0_outputs(10680));
    outputs(4480) <= not(layer0_outputs(4793));
    outputs(4481) <= not((layer0_outputs(10117)) or (layer0_outputs(9192)));
    outputs(4482) <= not(layer0_outputs(776));
    outputs(4483) <= (layer0_outputs(9110)) xor (layer0_outputs(5064));
    outputs(4484) <= (layer0_outputs(11820)) and not (layer0_outputs(9645));
    outputs(4485) <= not(layer0_outputs(2363)) or (layer0_outputs(9786));
    outputs(4486) <= (layer0_outputs(7809)) and (layer0_outputs(7115));
    outputs(4487) <= (layer0_outputs(7551)) or (layer0_outputs(3503));
    outputs(4488) <= (layer0_outputs(4713)) xor (layer0_outputs(768));
    outputs(4489) <= layer0_outputs(430);
    outputs(4490) <= not(layer0_outputs(11635)) or (layer0_outputs(9785));
    outputs(4491) <= not(layer0_outputs(1940));
    outputs(4492) <= not((layer0_outputs(6525)) or (layer0_outputs(3295)));
    outputs(4493) <= not(layer0_outputs(11335));
    outputs(4494) <= layer0_outputs(8109);
    outputs(4495) <= (layer0_outputs(3201)) xor (layer0_outputs(172));
    outputs(4496) <= not(layer0_outputs(5728)) or (layer0_outputs(8598));
    outputs(4497) <= layer0_outputs(3663);
    outputs(4498) <= layer0_outputs(10805);
    outputs(4499) <= (layer0_outputs(3611)) or (layer0_outputs(1864));
    outputs(4500) <= not((layer0_outputs(626)) or (layer0_outputs(2392)));
    outputs(4501) <= not(layer0_outputs(1815));
    outputs(4502) <= not(layer0_outputs(9782));
    outputs(4503) <= layer0_outputs(4737);
    outputs(4504) <= (layer0_outputs(6472)) xor (layer0_outputs(5709));
    outputs(4505) <= not(layer0_outputs(8453));
    outputs(4506) <= layer0_outputs(5403);
    outputs(4507) <= not(layer0_outputs(4891)) or (layer0_outputs(7697));
    outputs(4508) <= (layer0_outputs(8243)) and not (layer0_outputs(12751));
    outputs(4509) <= not(layer0_outputs(6619)) or (layer0_outputs(9471));
    outputs(4510) <= layer0_outputs(6096);
    outputs(4511) <= (layer0_outputs(5471)) and not (layer0_outputs(6713));
    outputs(4512) <= layer0_outputs(3217);
    outputs(4513) <= layer0_outputs(1898);
    outputs(4514) <= not(layer0_outputs(2265)) or (layer0_outputs(7211));
    outputs(4515) <= layer0_outputs(1065);
    outputs(4516) <= not(layer0_outputs(12300));
    outputs(4517) <= layer0_outputs(10664);
    outputs(4518) <= not(layer0_outputs(10144));
    outputs(4519) <= not(layer0_outputs(10219));
    outputs(4520) <= layer0_outputs(2807);
    outputs(4521) <= not(layer0_outputs(1300));
    outputs(4522) <= not(layer0_outputs(839));
    outputs(4523) <= (layer0_outputs(3601)) xor (layer0_outputs(7570));
    outputs(4524) <= not((layer0_outputs(1649)) xor (layer0_outputs(9074)));
    outputs(4525) <= not((layer0_outputs(7887)) xor (layer0_outputs(4812)));
    outputs(4526) <= layer0_outputs(4582);
    outputs(4527) <= (layer0_outputs(1889)) xor (layer0_outputs(1776));
    outputs(4528) <= (layer0_outputs(8500)) xor (layer0_outputs(9407));
    outputs(4529) <= layer0_outputs(8287);
    outputs(4530) <= not((layer0_outputs(4855)) xor (layer0_outputs(8032)));
    outputs(4531) <= not(layer0_outputs(2909));
    outputs(4532) <= not(layer0_outputs(3124));
    outputs(4533) <= (layer0_outputs(7152)) and not (layer0_outputs(7982));
    outputs(4534) <= (layer0_outputs(6162)) xor (layer0_outputs(5258));
    outputs(4535) <= layer0_outputs(2576);
    outputs(4536) <= not(layer0_outputs(11224));
    outputs(4537) <= not(layer0_outputs(6273));
    outputs(4538) <= (layer0_outputs(620)) xor (layer0_outputs(3165));
    outputs(4539) <= (layer0_outputs(7391)) and not (layer0_outputs(1758));
    outputs(4540) <= not((layer0_outputs(3034)) or (layer0_outputs(1994)));
    outputs(4541) <= not(layer0_outputs(2662));
    outputs(4542) <= layer0_outputs(8052);
    outputs(4543) <= layer0_outputs(6363);
    outputs(4544) <= (layer0_outputs(3313)) xor (layer0_outputs(2383));
    outputs(4545) <= layer0_outputs(6404);
    outputs(4546) <= layer0_outputs(1564);
    outputs(4547) <= not((layer0_outputs(12278)) xor (layer0_outputs(5627)));
    outputs(4548) <= not((layer0_outputs(1253)) xor (layer0_outputs(5723)));
    outputs(4549) <= layer0_outputs(2835);
    outputs(4550) <= layer0_outputs(6918);
    outputs(4551) <= (layer0_outputs(1666)) and (layer0_outputs(12347));
    outputs(4552) <= not(layer0_outputs(1492));
    outputs(4553) <= layer0_outputs(2580);
    outputs(4554) <= layer0_outputs(5020);
    outputs(4555) <= not(layer0_outputs(2734));
    outputs(4556) <= layer0_outputs(8475);
    outputs(4557) <= (layer0_outputs(9982)) and not (layer0_outputs(5503));
    outputs(4558) <= not((layer0_outputs(6587)) xor (layer0_outputs(11112)));
    outputs(4559) <= layer0_outputs(6031);
    outputs(4560) <= (layer0_outputs(12144)) and not (layer0_outputs(10798));
    outputs(4561) <= (layer0_outputs(2649)) xor (layer0_outputs(7443));
    outputs(4562) <= (layer0_outputs(5835)) and (layer0_outputs(7799));
    outputs(4563) <= layer0_outputs(7503);
    outputs(4564) <= (layer0_outputs(11555)) and not (layer0_outputs(5208));
    outputs(4565) <= (layer0_outputs(1619)) and not (layer0_outputs(12625));
    outputs(4566) <= not((layer0_outputs(6202)) or (layer0_outputs(11503)));
    outputs(4567) <= (layer0_outputs(6257)) and not (layer0_outputs(1492));
    outputs(4568) <= not(layer0_outputs(3065)) or (layer0_outputs(6421));
    outputs(4569) <= not(layer0_outputs(5815));
    outputs(4570) <= (layer0_outputs(11034)) and not (layer0_outputs(9306));
    outputs(4571) <= not((layer0_outputs(7550)) xor (layer0_outputs(11183)));
    outputs(4572) <= not(layer0_outputs(8431));
    outputs(4573) <= (layer0_outputs(1606)) and not (layer0_outputs(8364));
    outputs(4574) <= not(layer0_outputs(9409));
    outputs(4575) <= not((layer0_outputs(10705)) xor (layer0_outputs(12449)));
    outputs(4576) <= not(layer0_outputs(469));
    outputs(4577) <= (layer0_outputs(3723)) xor (layer0_outputs(7460));
    outputs(4578) <= not(layer0_outputs(11500));
    outputs(4579) <= not(layer0_outputs(9329)) or (layer0_outputs(8618));
    outputs(4580) <= layer0_outputs(9160);
    outputs(4581) <= not(layer0_outputs(8911)) or (layer0_outputs(9150));
    outputs(4582) <= not(layer0_outputs(8244));
    outputs(4583) <= layer0_outputs(6064);
    outputs(4584) <= (layer0_outputs(9242)) and (layer0_outputs(1504));
    outputs(4585) <= (layer0_outputs(5206)) xor (layer0_outputs(1063));
    outputs(4586) <= not((layer0_outputs(4171)) xor (layer0_outputs(7246)));
    outputs(4587) <= not(layer0_outputs(6414));
    outputs(4588) <= not((layer0_outputs(8759)) xor (layer0_outputs(7390)));
    outputs(4589) <= layer0_outputs(11436);
    outputs(4590) <= not(layer0_outputs(8322));
    outputs(4591) <= (layer0_outputs(3276)) xor (layer0_outputs(9987));
    outputs(4592) <= not((layer0_outputs(9481)) and (layer0_outputs(11945)));
    outputs(4593) <= (layer0_outputs(4068)) and not (layer0_outputs(5217));
    outputs(4594) <= layer0_outputs(5654);
    outputs(4595) <= not(layer0_outputs(6782));
    outputs(4596) <= (layer0_outputs(9032)) and not (layer0_outputs(12412));
    outputs(4597) <= (layer0_outputs(6298)) xor (layer0_outputs(2471));
    outputs(4598) <= layer0_outputs(8170);
    outputs(4599) <= not(layer0_outputs(10859));
    outputs(4600) <= layer0_outputs(10587);
    outputs(4601) <= not(layer0_outputs(5857));
    outputs(4602) <= (layer0_outputs(10312)) xor (layer0_outputs(7134));
    outputs(4603) <= not((layer0_outputs(4321)) xor (layer0_outputs(7089)));
    outputs(4604) <= not(layer0_outputs(193)) or (layer0_outputs(11771));
    outputs(4605) <= (layer0_outputs(9651)) xor (layer0_outputs(11361));
    outputs(4606) <= not(layer0_outputs(4052)) or (layer0_outputs(9212));
    outputs(4607) <= not(layer0_outputs(469));
    outputs(4608) <= (layer0_outputs(9123)) xor (layer0_outputs(8171));
    outputs(4609) <= layer0_outputs(8376);
    outputs(4610) <= not(layer0_outputs(7247));
    outputs(4611) <= (layer0_outputs(1053)) and not (layer0_outputs(4086));
    outputs(4612) <= layer0_outputs(8546);
    outputs(4613) <= (layer0_outputs(6926)) and (layer0_outputs(9107));
    outputs(4614) <= (layer0_outputs(6046)) xor (layer0_outputs(1725));
    outputs(4615) <= not(layer0_outputs(11116)) or (layer0_outputs(9259));
    outputs(4616) <= layer0_outputs(7197);
    outputs(4617) <= not((layer0_outputs(12625)) xor (layer0_outputs(2336)));
    outputs(4618) <= (layer0_outputs(1349)) and not (layer0_outputs(5813));
    outputs(4619) <= not(layer0_outputs(489));
    outputs(4620) <= not((layer0_outputs(11656)) xor (layer0_outputs(6204)));
    outputs(4621) <= not((layer0_outputs(4362)) and (layer0_outputs(12553)));
    outputs(4622) <= not((layer0_outputs(8490)) xor (layer0_outputs(12378)));
    outputs(4623) <= not(layer0_outputs(3261)) or (layer0_outputs(7836));
    outputs(4624) <= not(layer0_outputs(10375)) or (layer0_outputs(7302));
    outputs(4625) <= layer0_outputs(10731);
    outputs(4626) <= layer0_outputs(2357);
    outputs(4627) <= not(layer0_outputs(9504));
    outputs(4628) <= not((layer0_outputs(3543)) or (layer0_outputs(11627)));
    outputs(4629) <= (layer0_outputs(12750)) and not (layer0_outputs(11474));
    outputs(4630) <= (layer0_outputs(10005)) and not (layer0_outputs(10115));
    outputs(4631) <= not((layer0_outputs(10307)) xor (layer0_outputs(2152)));
    outputs(4632) <= not((layer0_outputs(12429)) xor (layer0_outputs(125)));
    outputs(4633) <= not((layer0_outputs(3483)) or (layer0_outputs(10778)));
    outputs(4634) <= not((layer0_outputs(4762)) and (layer0_outputs(5942)));
    outputs(4635) <= layer0_outputs(2461);
    outputs(4636) <= layer0_outputs(7825);
    outputs(4637) <= layer0_outputs(2597);
    outputs(4638) <= layer0_outputs(5861);
    outputs(4639) <= not(layer0_outputs(249));
    outputs(4640) <= not(layer0_outputs(9090)) or (layer0_outputs(10695));
    outputs(4641) <= (layer0_outputs(10099)) xor (layer0_outputs(1633));
    outputs(4642) <= layer0_outputs(9070);
    outputs(4643) <= not(layer0_outputs(12522));
    outputs(4644) <= not(layer0_outputs(9962)) or (layer0_outputs(8169));
    outputs(4645) <= not((layer0_outputs(6543)) xor (layer0_outputs(7754)));
    outputs(4646) <= layer0_outputs(2863);
    outputs(4647) <= layer0_outputs(11298);
    outputs(4648) <= not(layer0_outputs(5479));
    outputs(4649) <= not(layer0_outputs(822)) or (layer0_outputs(3430));
    outputs(4650) <= not(layer0_outputs(4393));
    outputs(4651) <= (layer0_outputs(8016)) and not (layer0_outputs(11241));
    outputs(4652) <= not((layer0_outputs(10144)) and (layer0_outputs(11484)));
    outputs(4653) <= (layer0_outputs(5419)) xor (layer0_outputs(6444));
    outputs(4654) <= (layer0_outputs(7386)) xor (layer0_outputs(4517));
    outputs(4655) <= layer0_outputs(2663);
    outputs(4656) <= not(layer0_outputs(7599));
    outputs(4657) <= not(layer0_outputs(4800));
    outputs(4658) <= (layer0_outputs(8031)) and not (layer0_outputs(10101));
    outputs(4659) <= (layer0_outputs(393)) and not (layer0_outputs(271));
    outputs(4660) <= not(layer0_outputs(1934));
    outputs(4661) <= not(layer0_outputs(4378));
    outputs(4662) <= (layer0_outputs(10103)) and not (layer0_outputs(3037));
    outputs(4663) <= not(layer0_outputs(1671));
    outputs(4664) <= not((layer0_outputs(1788)) xor (layer0_outputs(5797)));
    outputs(4665) <= not((layer0_outputs(336)) or (layer0_outputs(6236)));
    outputs(4666) <= not((layer0_outputs(9299)) xor (layer0_outputs(11610)));
    outputs(4667) <= (layer0_outputs(10231)) and not (layer0_outputs(817));
    outputs(4668) <= layer0_outputs(5735);
    outputs(4669) <= not((layer0_outputs(1325)) xor (layer0_outputs(9653)));
    outputs(4670) <= (layer0_outputs(11477)) xor (layer0_outputs(3733));
    outputs(4671) <= (layer0_outputs(453)) and (layer0_outputs(3244));
    outputs(4672) <= layer0_outputs(6662);
    outputs(4673) <= not(layer0_outputs(9330));
    outputs(4674) <= not((layer0_outputs(60)) xor (layer0_outputs(9812)));
    outputs(4675) <= (layer0_outputs(3579)) and not (layer0_outputs(8294));
    outputs(4676) <= not((layer0_outputs(12425)) xor (layer0_outputs(9691)));
    outputs(4677) <= not(layer0_outputs(465));
    outputs(4678) <= (layer0_outputs(10454)) and (layer0_outputs(6053));
    outputs(4679) <= not(layer0_outputs(10510));
    outputs(4680) <= not(layer0_outputs(11386));
    outputs(4681) <= not((layer0_outputs(5742)) xor (layer0_outputs(3191)));
    outputs(4682) <= (layer0_outputs(3951)) and not (layer0_outputs(1475));
    outputs(4683) <= not(layer0_outputs(2012));
    outputs(4684) <= not(layer0_outputs(4520));
    outputs(4685) <= layer0_outputs(6406);
    outputs(4686) <= not((layer0_outputs(3385)) xor (layer0_outputs(4272)));
    outputs(4687) <= layer0_outputs(7504);
    outputs(4688) <= layer0_outputs(3098);
    outputs(4689) <= (layer0_outputs(1962)) and (layer0_outputs(7673));
    outputs(4690) <= not(layer0_outputs(978));
    outputs(4691) <= not(layer0_outputs(12521));
    outputs(4692) <= (layer0_outputs(11753)) or (layer0_outputs(8147));
    outputs(4693) <= not((layer0_outputs(3243)) or (layer0_outputs(1136)));
    outputs(4694) <= not((layer0_outputs(2446)) xor (layer0_outputs(6635)));
    outputs(4695) <= not((layer0_outputs(5722)) xor (layer0_outputs(9642)));
    outputs(4696) <= (layer0_outputs(3796)) xor (layer0_outputs(7905));
    outputs(4697) <= not((layer0_outputs(11926)) xor (layer0_outputs(30)));
    outputs(4698) <= (layer0_outputs(380)) xor (layer0_outputs(8465));
    outputs(4699) <= not(layer0_outputs(3453));
    outputs(4700) <= (layer0_outputs(12436)) and not (layer0_outputs(10432));
    outputs(4701) <= not(layer0_outputs(9099));
    outputs(4702) <= (layer0_outputs(8517)) and not (layer0_outputs(9573));
    outputs(4703) <= (layer0_outputs(10795)) xor (layer0_outputs(143));
    outputs(4704) <= not((layer0_outputs(8271)) or (layer0_outputs(10372)));
    outputs(4705) <= (layer0_outputs(12689)) and (layer0_outputs(4553));
    outputs(4706) <= layer0_outputs(2599);
    outputs(4707) <= layer0_outputs(10265);
    outputs(4708) <= (layer0_outputs(12628)) and not (layer0_outputs(1990));
    outputs(4709) <= not((layer0_outputs(5147)) or (layer0_outputs(1762)));
    outputs(4710) <= not((layer0_outputs(4163)) xor (layer0_outputs(5426)));
    outputs(4711) <= layer0_outputs(4584);
    outputs(4712) <= (layer0_outputs(190)) or (layer0_outputs(7700));
    outputs(4713) <= layer0_outputs(5998);
    outputs(4714) <= not((layer0_outputs(6556)) xor (layer0_outputs(7357)));
    outputs(4715) <= not((layer0_outputs(1479)) xor (layer0_outputs(7289)));
    outputs(4716) <= layer0_outputs(6596);
    outputs(4717) <= not((layer0_outputs(8982)) or (layer0_outputs(420)));
    outputs(4718) <= (layer0_outputs(3205)) and not (layer0_outputs(12090));
    outputs(4719) <= not((layer0_outputs(11047)) xor (layer0_outputs(6324)));
    outputs(4720) <= not((layer0_outputs(12544)) and (layer0_outputs(4228)));
    outputs(4721) <= layer0_outputs(3060);
    outputs(4722) <= layer0_outputs(7621);
    outputs(4723) <= not(layer0_outputs(6271)) or (layer0_outputs(10095));
    outputs(4724) <= not((layer0_outputs(7268)) or (layer0_outputs(122)));
    outputs(4725) <= not((layer0_outputs(10873)) or (layer0_outputs(12563)));
    outputs(4726) <= layer0_outputs(5410);
    outputs(4727) <= not((layer0_outputs(2041)) or (layer0_outputs(3760)));
    outputs(4728) <= '1';
    outputs(4729) <= layer0_outputs(4890);
    outputs(4730) <= (layer0_outputs(7626)) xor (layer0_outputs(11703));
    outputs(4731) <= layer0_outputs(10286);
    outputs(4732) <= (layer0_outputs(11977)) xor (layer0_outputs(732));
    outputs(4733) <= (layer0_outputs(10588)) or (layer0_outputs(7913));
    outputs(4734) <= (layer0_outputs(3708)) and not (layer0_outputs(10010));
    outputs(4735) <= layer0_outputs(3305);
    outputs(4736) <= not(layer0_outputs(10136));
    outputs(4737) <= layer0_outputs(5686);
    outputs(4738) <= not(layer0_outputs(8539));
    outputs(4739) <= (layer0_outputs(7910)) xor (layer0_outputs(6271));
    outputs(4740) <= not(layer0_outputs(2323));
    outputs(4741) <= (layer0_outputs(11812)) xor (layer0_outputs(8817));
    outputs(4742) <= layer0_outputs(4985);
    outputs(4743) <= layer0_outputs(4760);
    outputs(4744) <= not((layer0_outputs(1778)) and (layer0_outputs(10321)));
    outputs(4745) <= (layer0_outputs(9213)) and not (layer0_outputs(11374));
    outputs(4746) <= (layer0_outputs(7379)) or (layer0_outputs(9477));
    outputs(4747) <= not(layer0_outputs(836));
    outputs(4748) <= not((layer0_outputs(2751)) xor (layer0_outputs(2845)));
    outputs(4749) <= (layer0_outputs(8668)) and not (layer0_outputs(5464));
    outputs(4750) <= not((layer0_outputs(6147)) xor (layer0_outputs(1241)));
    outputs(4751) <= not(layer0_outputs(11375)) or (layer0_outputs(3722));
    outputs(4752) <= not(layer0_outputs(11308));
    outputs(4753) <= (layer0_outputs(5975)) xor (layer0_outputs(12601));
    outputs(4754) <= not((layer0_outputs(2594)) and (layer0_outputs(11484)));
    outputs(4755) <= layer0_outputs(8284);
    outputs(4756) <= (layer0_outputs(8607)) and not (layer0_outputs(10919));
    outputs(4757) <= not(layer0_outputs(1775));
    outputs(4758) <= not((layer0_outputs(10923)) or (layer0_outputs(10858)));
    outputs(4759) <= not(layer0_outputs(5621));
    outputs(4760) <= not((layer0_outputs(9758)) or (layer0_outputs(2625)));
    outputs(4761) <= not(layer0_outputs(4599));
    outputs(4762) <= layer0_outputs(1482);
    outputs(4763) <= layer0_outputs(274);
    outputs(4764) <= not(layer0_outputs(6502));
    outputs(4765) <= (layer0_outputs(12115)) and not (layer0_outputs(9431));
    outputs(4766) <= not((layer0_outputs(11038)) xor (layer0_outputs(8862)));
    outputs(4767) <= not(layer0_outputs(10725));
    outputs(4768) <= not((layer0_outputs(10496)) and (layer0_outputs(12208)));
    outputs(4769) <= layer0_outputs(10669);
    outputs(4770) <= not((layer0_outputs(433)) xor (layer0_outputs(8856)));
    outputs(4771) <= layer0_outputs(5225);
    outputs(4772) <= layer0_outputs(11265);
    outputs(4773) <= (layer0_outputs(4300)) or (layer0_outputs(5109));
    outputs(4774) <= not((layer0_outputs(12532)) and (layer0_outputs(12518)));
    outputs(4775) <= layer0_outputs(654);
    outputs(4776) <= not(layer0_outputs(644));
    outputs(4777) <= not(layer0_outputs(3411)) or (layer0_outputs(155));
    outputs(4778) <= layer0_outputs(12460);
    outputs(4779) <= layer0_outputs(1016);
    outputs(4780) <= not(layer0_outputs(3433));
    outputs(4781) <= (layer0_outputs(12048)) xor (layer0_outputs(9675));
    outputs(4782) <= (layer0_outputs(4992)) or (layer0_outputs(9503));
    outputs(4783) <= (layer0_outputs(10450)) and not (layer0_outputs(9398));
    outputs(4784) <= not((layer0_outputs(5393)) xor (layer0_outputs(5751)));
    outputs(4785) <= not(layer0_outputs(3433));
    outputs(4786) <= not(layer0_outputs(6762));
    outputs(4787) <= layer0_outputs(11462);
    outputs(4788) <= not((layer0_outputs(11469)) and (layer0_outputs(4471)));
    outputs(4789) <= (layer0_outputs(5831)) and not (layer0_outputs(11093));
    outputs(4790) <= (layer0_outputs(2531)) xor (layer0_outputs(7614));
    outputs(4791) <= (layer0_outputs(553)) xor (layer0_outputs(8246));
    outputs(4792) <= not((layer0_outputs(12071)) xor (layer0_outputs(208)));
    outputs(4793) <= layer0_outputs(10106);
    outputs(4794) <= not(layer0_outputs(1541));
    outputs(4795) <= (layer0_outputs(10368)) and not (layer0_outputs(4537));
    outputs(4796) <= layer0_outputs(6303);
    outputs(4797) <= not(layer0_outputs(3130)) or (layer0_outputs(2940));
    outputs(4798) <= not(layer0_outputs(2728)) or (layer0_outputs(7084));
    outputs(4799) <= (layer0_outputs(1665)) xor (layer0_outputs(1607));
    outputs(4800) <= (layer0_outputs(7968)) and not (layer0_outputs(1814));
    outputs(4801) <= (layer0_outputs(1687)) xor (layer0_outputs(9688));
    outputs(4802) <= (layer0_outputs(11354)) and not (layer0_outputs(4183));
    outputs(4803) <= (layer0_outputs(133)) xor (layer0_outputs(2920));
    outputs(4804) <= not(layer0_outputs(3465));
    outputs(4805) <= not((layer0_outputs(12392)) xor (layer0_outputs(12674)));
    outputs(4806) <= layer0_outputs(8125);
    outputs(4807) <= not(layer0_outputs(783));
    outputs(4808) <= not((layer0_outputs(7579)) xor (layer0_outputs(2011)));
    outputs(4809) <= not(layer0_outputs(11845)) or (layer0_outputs(5119));
    outputs(4810) <= not(layer0_outputs(8340));
    outputs(4811) <= (layer0_outputs(10955)) and not (layer0_outputs(11625));
    outputs(4812) <= (layer0_outputs(5135)) and not (layer0_outputs(10618));
    outputs(4813) <= (layer0_outputs(12789)) xor (layer0_outputs(12230));
    outputs(4814) <= (layer0_outputs(3616)) or (layer0_outputs(2959));
    outputs(4815) <= not(layer0_outputs(8021)) or (layer0_outputs(11010));
    outputs(4816) <= not(layer0_outputs(11599));
    outputs(4817) <= not(layer0_outputs(3557));
    outputs(4818) <= not(layer0_outputs(12678));
    outputs(4819) <= layer0_outputs(3965);
    outputs(4820) <= not(layer0_outputs(11103));
    outputs(4821) <= not((layer0_outputs(6803)) and (layer0_outputs(1989)));
    outputs(4822) <= layer0_outputs(1824);
    outputs(4823) <= not(layer0_outputs(6532));
    outputs(4824) <= not((layer0_outputs(4206)) or (layer0_outputs(10165)));
    outputs(4825) <= (layer0_outputs(42)) and not (layer0_outputs(12507));
    outputs(4826) <= not((layer0_outputs(12306)) or (layer0_outputs(11444)));
    outputs(4827) <= not(layer0_outputs(9133));
    outputs(4828) <= (layer0_outputs(659)) xor (layer0_outputs(10867));
    outputs(4829) <= layer0_outputs(3859);
    outputs(4830) <= (layer0_outputs(6128)) or (layer0_outputs(2678));
    outputs(4831) <= layer0_outputs(6706);
    outputs(4832) <= layer0_outputs(314);
    outputs(4833) <= layer0_outputs(2318);
    outputs(4834) <= (layer0_outputs(3095)) xor (layer0_outputs(10299));
    outputs(4835) <= layer0_outputs(4864);
    outputs(4836) <= layer0_outputs(8686);
    outputs(4837) <= not((layer0_outputs(8958)) xor (layer0_outputs(9745)));
    outputs(4838) <= layer0_outputs(1256);
    outputs(4839) <= not((layer0_outputs(11725)) xor (layer0_outputs(6101)));
    outputs(4840) <= not((layer0_outputs(6733)) and (layer0_outputs(2992)));
    outputs(4841) <= (layer0_outputs(7412)) and (layer0_outputs(10329));
    outputs(4842) <= not(layer0_outputs(11225));
    outputs(4843) <= layer0_outputs(6130);
    outputs(4844) <= not(layer0_outputs(9737));
    outputs(4845) <= layer0_outputs(5747);
    outputs(4846) <= (layer0_outputs(3037)) xor (layer0_outputs(8184));
    outputs(4847) <= not((layer0_outputs(1097)) xor (layer0_outputs(2984)));
    outputs(4848) <= not((layer0_outputs(7718)) or (layer0_outputs(6663)));
    outputs(4849) <= layer0_outputs(4763);
    outputs(4850) <= not((layer0_outputs(1654)) xor (layer0_outputs(7407)));
    outputs(4851) <= not(layer0_outputs(3661)) or (layer0_outputs(4674));
    outputs(4852) <= layer0_outputs(4056);
    outputs(4853) <= layer0_outputs(3741);
    outputs(4854) <= not(layer0_outputs(5434));
    outputs(4855) <= (layer0_outputs(998)) xor (layer0_outputs(11923));
    outputs(4856) <= not(layer0_outputs(8631));
    outputs(4857) <= not(layer0_outputs(1719));
    outputs(4858) <= not((layer0_outputs(8993)) xor (layer0_outputs(11714)));
    outputs(4859) <= not(layer0_outputs(8999));
    outputs(4860) <= layer0_outputs(4112);
    outputs(4861) <= (layer0_outputs(3614)) xor (layer0_outputs(2629));
    outputs(4862) <= layer0_outputs(6002);
    outputs(4863) <= not(layer0_outputs(1522)) or (layer0_outputs(9359));
    outputs(4864) <= (layer0_outputs(162)) xor (layer0_outputs(2660));
    outputs(4865) <= (layer0_outputs(7670)) xor (layer0_outputs(3410));
    outputs(4866) <= not((layer0_outputs(6927)) xor (layer0_outputs(2032)));
    outputs(4867) <= layer0_outputs(11743);
    outputs(4868) <= not(layer0_outputs(12469));
    outputs(4869) <= layer0_outputs(3593);
    outputs(4870) <= not(layer0_outputs(4843)) or (layer0_outputs(9535));
    outputs(4871) <= not(layer0_outputs(389)) or (layer0_outputs(11723));
    outputs(4872) <= layer0_outputs(4335);
    outputs(4873) <= (layer0_outputs(5780)) and (layer0_outputs(4386));
    outputs(4874) <= not((layer0_outputs(2969)) xor (layer0_outputs(1817)));
    outputs(4875) <= layer0_outputs(296);
    outputs(4876) <= not((layer0_outputs(6420)) or (layer0_outputs(774)));
    outputs(4877) <= not(layer0_outputs(4373));
    outputs(4878) <= (layer0_outputs(3793)) xor (layer0_outputs(596));
    outputs(4879) <= not((layer0_outputs(11674)) xor (layer0_outputs(9797)));
    outputs(4880) <= layer0_outputs(5593);
    outputs(4881) <= not((layer0_outputs(3837)) and (layer0_outputs(3791)));
    outputs(4882) <= (layer0_outputs(8764)) xor (layer0_outputs(11164));
    outputs(4883) <= layer0_outputs(8153);
    outputs(4884) <= (layer0_outputs(7077)) and not (layer0_outputs(7307));
    outputs(4885) <= not(layer0_outputs(8441));
    outputs(4886) <= not(layer0_outputs(7546));
    outputs(4887) <= (layer0_outputs(4983)) xor (layer0_outputs(8471));
    outputs(4888) <= layer0_outputs(9259);
    outputs(4889) <= layer0_outputs(11917);
    outputs(4890) <= layer0_outputs(11946);
    outputs(4891) <= (layer0_outputs(334)) xor (layer0_outputs(434));
    outputs(4892) <= not((layer0_outputs(9006)) and (layer0_outputs(4807)));
    outputs(4893) <= not(layer0_outputs(4952));
    outputs(4894) <= not((layer0_outputs(2825)) and (layer0_outputs(12140)));
    outputs(4895) <= layer0_outputs(9998);
    outputs(4896) <= layer0_outputs(3396);
    outputs(4897) <= layer0_outputs(6521);
    outputs(4898) <= not((layer0_outputs(8722)) xor (layer0_outputs(5889)));
    outputs(4899) <= (layer0_outputs(5854)) and not (layer0_outputs(5413));
    outputs(4900) <= not((layer0_outputs(8673)) and (layer0_outputs(1699)));
    outputs(4901) <= (layer0_outputs(3901)) and not (layer0_outputs(2511));
    outputs(4902) <= not((layer0_outputs(11458)) and (layer0_outputs(1534)));
    outputs(4903) <= not(layer0_outputs(5003)) or (layer0_outputs(8560));
    outputs(4904) <= (layer0_outputs(10883)) xor (layer0_outputs(11396));
    outputs(4905) <= not(layer0_outputs(12773));
    outputs(4906) <= layer0_outputs(1992);
    outputs(4907) <= (layer0_outputs(1539)) xor (layer0_outputs(354));
    outputs(4908) <= layer0_outputs(8579);
    outputs(4909) <= not(layer0_outputs(9390));
    outputs(4910) <= layer0_outputs(9063);
    outputs(4911) <= not(layer0_outputs(2183));
    outputs(4912) <= not(layer0_outputs(9619));
    outputs(4913) <= (layer0_outputs(2690)) and not (layer0_outputs(11655));
    outputs(4914) <= not(layer0_outputs(5859));
    outputs(4915) <= not(layer0_outputs(3984));
    outputs(4916) <= layer0_outputs(8679);
    outputs(4917) <= not((layer0_outputs(3985)) or (layer0_outputs(10661)));
    outputs(4918) <= (layer0_outputs(12180)) and (layer0_outputs(4569));
    outputs(4919) <= (layer0_outputs(9379)) or (layer0_outputs(5214));
    outputs(4920) <= (layer0_outputs(6752)) and not (layer0_outputs(9009));
    outputs(4921) <= not(layer0_outputs(2345)) or (layer0_outputs(618));
    outputs(4922) <= (layer0_outputs(1273)) xor (layer0_outputs(1079));
    outputs(4923) <= (layer0_outputs(6614)) and (layer0_outputs(1955));
    outputs(4924) <= not((layer0_outputs(2917)) xor (layer0_outputs(8537)));
    outputs(4925) <= layer0_outputs(973);
    outputs(4926) <= layer0_outputs(1786);
    outputs(4927) <= layer0_outputs(9723);
    outputs(4928) <= (layer0_outputs(2508)) and not (layer0_outputs(3409));
    outputs(4929) <= not(layer0_outputs(104));
    outputs(4930) <= (layer0_outputs(1101)) xor (layer0_outputs(10803));
    outputs(4931) <= (layer0_outputs(1307)) and not (layer0_outputs(2608));
    outputs(4932) <= not((layer0_outputs(4079)) xor (layer0_outputs(10038)));
    outputs(4933) <= not(layer0_outputs(7464));
    outputs(4934) <= (layer0_outputs(5954)) and not (layer0_outputs(9435));
    outputs(4935) <= (layer0_outputs(6885)) or (layer0_outputs(7699));
    outputs(4936) <= layer0_outputs(924);
    outputs(4937) <= not((layer0_outputs(8460)) xor (layer0_outputs(9843)));
    outputs(4938) <= not((layer0_outputs(7650)) and (layer0_outputs(10760)));
    outputs(4939) <= layer0_outputs(2128);
    outputs(4940) <= not(layer0_outputs(10047));
    outputs(4941) <= (layer0_outputs(276)) xor (layer0_outputs(10399));
    outputs(4942) <= not(layer0_outputs(2049)) or (layer0_outputs(3217));
    outputs(4943) <= not(layer0_outputs(1728)) or (layer0_outputs(5914));
    outputs(4944) <= not(layer0_outputs(3820));
    outputs(4945) <= not(layer0_outputs(8893)) or (layer0_outputs(3415));
    outputs(4946) <= not(layer0_outputs(3896));
    outputs(4947) <= not((layer0_outputs(6270)) xor (layer0_outputs(4219)));
    outputs(4948) <= layer0_outputs(10028);
    outputs(4949) <= not(layer0_outputs(2135));
    outputs(4950) <= not(layer0_outputs(4715));
    outputs(4951) <= layer0_outputs(437);
    outputs(4952) <= not(layer0_outputs(5561));
    outputs(4953) <= not(layer0_outputs(12656));
    outputs(4954) <= not(layer0_outputs(4545));
    outputs(4955) <= not(layer0_outputs(4689));
    outputs(4956) <= not((layer0_outputs(4413)) and (layer0_outputs(10154)));
    outputs(4957) <= layer0_outputs(1288);
    outputs(4958) <= not((layer0_outputs(9783)) xor (layer0_outputs(9056)));
    outputs(4959) <= (layer0_outputs(8138)) xor (layer0_outputs(4279));
    outputs(4960) <= not(layer0_outputs(10545));
    outputs(4961) <= not((layer0_outputs(9344)) xor (layer0_outputs(3301)));
    outputs(4962) <= not(layer0_outputs(2711)) or (layer0_outputs(7036));
    outputs(4963) <= not((layer0_outputs(9313)) xor (layer0_outputs(11672)));
    outputs(4964) <= layer0_outputs(3437);
    outputs(4965) <= layer0_outputs(12592);
    outputs(4966) <= '0';
    outputs(4967) <= not(layer0_outputs(10285)) or (layer0_outputs(10351));
    outputs(4968) <= not((layer0_outputs(2109)) and (layer0_outputs(7623)));
    outputs(4969) <= (layer0_outputs(3894)) and not (layer0_outputs(4966));
    outputs(4970) <= (layer0_outputs(6712)) and not (layer0_outputs(1442));
    outputs(4971) <= not(layer0_outputs(3124));
    outputs(4972) <= layer0_outputs(2210);
    outputs(4973) <= not(layer0_outputs(9307)) or (layer0_outputs(3447));
    outputs(4974) <= not((layer0_outputs(9562)) and (layer0_outputs(6655)));
    outputs(4975) <= layer0_outputs(4978);
    outputs(4976) <= layer0_outputs(10687);
    outputs(4977) <= layer0_outputs(11779);
    outputs(4978) <= (layer0_outputs(11785)) and not (layer0_outputs(7806));
    outputs(4979) <= not((layer0_outputs(9220)) xor (layer0_outputs(6356)));
    outputs(4980) <= (layer0_outputs(7106)) and (layer0_outputs(6029));
    outputs(4981) <= not(layer0_outputs(4678));
    outputs(4982) <= (layer0_outputs(10261)) and not (layer0_outputs(8249));
    outputs(4983) <= (layer0_outputs(7091)) or (layer0_outputs(11193));
    outputs(4984) <= not(layer0_outputs(2994));
    outputs(4985) <= (layer0_outputs(10034)) xor (layer0_outputs(3086));
    outputs(4986) <= layer0_outputs(11450);
    outputs(4987) <= (layer0_outputs(1437)) or (layer0_outputs(1772));
    outputs(4988) <= not((layer0_outputs(4430)) xor (layer0_outputs(12616)));
    outputs(4989) <= (layer0_outputs(10810)) and not (layer0_outputs(12174));
    outputs(4990) <= (layer0_outputs(8511)) or (layer0_outputs(8947));
    outputs(4991) <= layer0_outputs(3191);
    outputs(4992) <= (layer0_outputs(9673)) and not (layer0_outputs(1812));
    outputs(4993) <= not(layer0_outputs(8383));
    outputs(4994) <= not(layer0_outputs(885));
    outputs(4995) <= (layer0_outputs(8873)) and (layer0_outputs(12099));
    outputs(4996) <= layer0_outputs(11312);
    outputs(4997) <= (layer0_outputs(10782)) and (layer0_outputs(1820));
    outputs(4998) <= (layer0_outputs(11824)) and not (layer0_outputs(2456));
    outputs(4999) <= layer0_outputs(12177);
    outputs(5000) <= not((layer0_outputs(11925)) xor (layer0_outputs(12676)));
    outputs(5001) <= (layer0_outputs(10952)) and not (layer0_outputs(7648));
    outputs(5002) <= not(layer0_outputs(10211));
    outputs(5003) <= layer0_outputs(10776);
    outputs(5004) <= not(layer0_outputs(8697));
    outputs(5005) <= not((layer0_outputs(10610)) xor (layer0_outputs(4995)));
    outputs(5006) <= not(layer0_outputs(2793));
    outputs(5007) <= (layer0_outputs(11950)) and (layer0_outputs(5625));
    outputs(5008) <= (layer0_outputs(12620)) xor (layer0_outputs(9300));
    outputs(5009) <= (layer0_outputs(11407)) and (layer0_outputs(1428));
    outputs(5010) <= (layer0_outputs(8096)) and not (layer0_outputs(9099));
    outputs(5011) <= not((layer0_outputs(9162)) xor (layer0_outputs(5321)));
    outputs(5012) <= not(layer0_outputs(10100));
    outputs(5013) <= not(layer0_outputs(1529));
    outputs(5014) <= not((layer0_outputs(1402)) or (layer0_outputs(4398)));
    outputs(5015) <= not(layer0_outputs(439));
    outputs(5016) <= layer0_outputs(7271);
    outputs(5017) <= not((layer0_outputs(2057)) xor (layer0_outputs(3768)));
    outputs(5018) <= layer0_outputs(9915);
    outputs(5019) <= (layer0_outputs(5379)) and not (layer0_outputs(111));
    outputs(5020) <= not(layer0_outputs(6298)) or (layer0_outputs(3983));
    outputs(5021) <= not(layer0_outputs(10247));
    outputs(5022) <= not(layer0_outputs(4182));
    outputs(5023) <= (layer0_outputs(7545)) or (layer0_outputs(991));
    outputs(5024) <= layer0_outputs(6643);
    outputs(5025) <= not(layer0_outputs(12154));
    outputs(5026) <= not(layer0_outputs(12072));
    outputs(5027) <= layer0_outputs(4474);
    outputs(5028) <= not(layer0_outputs(6583));
    outputs(5029) <= not((layer0_outputs(6399)) xor (layer0_outputs(5020)));
    outputs(5030) <= not(layer0_outputs(4612));
    outputs(5031) <= (layer0_outputs(11854)) and not (layer0_outputs(7848));
    outputs(5032) <= layer0_outputs(1416);
    outputs(5033) <= not(layer0_outputs(8654));
    outputs(5034) <= layer0_outputs(2460);
    outputs(5035) <= (layer0_outputs(4720)) and not (layer0_outputs(1806));
    outputs(5036) <= not((layer0_outputs(3471)) xor (layer0_outputs(2034)));
    outputs(5037) <= layer0_outputs(12228);
    outputs(5038) <= layer0_outputs(3450);
    outputs(5039) <= not((layer0_outputs(2444)) xor (layer0_outputs(1501)));
    outputs(5040) <= not(layer0_outputs(9814)) or (layer0_outputs(310));
    outputs(5041) <= not(layer0_outputs(3038));
    outputs(5042) <= not((layer0_outputs(8921)) xor (layer0_outputs(4829)));
    outputs(5043) <= (layer0_outputs(9097)) xor (layer0_outputs(923));
    outputs(5044) <= not(layer0_outputs(2529)) or (layer0_outputs(4252));
    outputs(5045) <= layer0_outputs(6871);
    outputs(5046) <= not((layer0_outputs(6065)) xor (layer0_outputs(2958)));
    outputs(5047) <= layer0_outputs(2264);
    outputs(5048) <= not(layer0_outputs(8299));
    outputs(5049) <= not((layer0_outputs(8331)) or (layer0_outputs(11052)));
    outputs(5050) <= not(layer0_outputs(1876));
    outputs(5051) <= not(layer0_outputs(10529));
    outputs(5052) <= not(layer0_outputs(2249));
    outputs(5053) <= not(layer0_outputs(5706));
    outputs(5054) <= (layer0_outputs(3490)) xor (layer0_outputs(8556));
    outputs(5055) <= layer0_outputs(1657);
    outputs(5056) <= not(layer0_outputs(9923)) or (layer0_outputs(6965));
    outputs(5057) <= not(layer0_outputs(11433));
    outputs(5058) <= layer0_outputs(4251);
    outputs(5059) <= layer0_outputs(634);
    outputs(5060) <= not((layer0_outputs(4375)) and (layer0_outputs(10042)));
    outputs(5061) <= layer0_outputs(328);
    outputs(5062) <= not(layer0_outputs(5540));
    outputs(5063) <= (layer0_outputs(3732)) and not (layer0_outputs(5273));
    outputs(5064) <= (layer0_outputs(6184)) and (layer0_outputs(8876));
    outputs(5065) <= layer0_outputs(8263);
    outputs(5066) <= (layer0_outputs(10547)) and not (layer0_outputs(8355));
    outputs(5067) <= not((layer0_outputs(4162)) xor (layer0_outputs(6057)));
    outputs(5068) <= not(layer0_outputs(4077));
    outputs(5069) <= (layer0_outputs(6119)) xor (layer0_outputs(8246));
    outputs(5070) <= layer0_outputs(10265);
    outputs(5071) <= not(layer0_outputs(3106));
    outputs(5072) <= (layer0_outputs(8090)) or (layer0_outputs(9676));
    outputs(5073) <= not(layer0_outputs(2913));
    outputs(5074) <= not(layer0_outputs(407));
    outputs(5075) <= not(layer0_outputs(8996));
    outputs(5076) <= not(layer0_outputs(3955));
    outputs(5077) <= not(layer0_outputs(12141));
    outputs(5078) <= not(layer0_outputs(6578));
    outputs(5079) <= (layer0_outputs(2860)) and not (layer0_outputs(9528));
    outputs(5080) <= layer0_outputs(6213);
    outputs(5081) <= not((layer0_outputs(6770)) xor (layer0_outputs(2732)));
    outputs(5082) <= (layer0_outputs(4912)) xor (layer0_outputs(1247));
    outputs(5083) <= not(layer0_outputs(2872));
    outputs(5084) <= not(layer0_outputs(10222));
    outputs(5085) <= (layer0_outputs(8100)) xor (layer0_outputs(9873));
    outputs(5086) <= not(layer0_outputs(9824)) or (layer0_outputs(6813));
    outputs(5087) <= layer0_outputs(7323);
    outputs(5088) <= (layer0_outputs(860)) and (layer0_outputs(11680));
    outputs(5089) <= (layer0_outputs(7066)) and not (layer0_outputs(3945));
    outputs(5090) <= not(layer0_outputs(158)) or (layer0_outputs(7978));
    outputs(5091) <= layer0_outputs(367);
    outputs(5092) <= (layer0_outputs(12101)) and (layer0_outputs(5268));
    outputs(5093) <= layer0_outputs(8208);
    outputs(5094) <= not(layer0_outputs(7163));
    outputs(5095) <= (layer0_outputs(11848)) xor (layer0_outputs(791));
    outputs(5096) <= not(layer0_outputs(1200)) or (layer0_outputs(3857));
    outputs(5097) <= layer0_outputs(12462);
    outputs(5098) <= not((layer0_outputs(9963)) xor (layer0_outputs(5733)));
    outputs(5099) <= (layer0_outputs(2895)) and not (layer0_outputs(12434));
    outputs(5100) <= not(layer0_outputs(925)) or (layer0_outputs(9157));
    outputs(5101) <= not((layer0_outputs(5933)) or (layer0_outputs(4181)));
    outputs(5102) <= not(layer0_outputs(685)) or (layer0_outputs(11333));
    outputs(5103) <= (layer0_outputs(4102)) and not (layer0_outputs(7473));
    outputs(5104) <= (layer0_outputs(9740)) xor (layer0_outputs(11089));
    outputs(5105) <= (layer0_outputs(1689)) and (layer0_outputs(5141));
    outputs(5106) <= (layer0_outputs(1120)) and not (layer0_outputs(10934));
    outputs(5107) <= layer0_outputs(12301);
    outputs(5108) <= (layer0_outputs(8269)) and (layer0_outputs(3254));
    outputs(5109) <= not(layer0_outputs(5759)) or (layer0_outputs(7903));
    outputs(5110) <= not(layer0_outputs(10771));
    outputs(5111) <= not(layer0_outputs(9712));
    outputs(5112) <= layer0_outputs(805);
    outputs(5113) <= not((layer0_outputs(6004)) or (layer0_outputs(4539)));
    outputs(5114) <= not(layer0_outputs(1073));
    outputs(5115) <= (layer0_outputs(5414)) or (layer0_outputs(12664));
    outputs(5116) <= not(layer0_outputs(5490));
    outputs(5117) <= not(layer0_outputs(2025));
    outputs(5118) <= (layer0_outputs(2888)) and not (layer0_outputs(5895));
    outputs(5119) <= not((layer0_outputs(10382)) xor (layer0_outputs(5431)));
    outputs(5120) <= layer0_outputs(6249);
    outputs(5121) <= layer0_outputs(2272);
    outputs(5122) <= (layer0_outputs(11620)) and not (layer0_outputs(4414));
    outputs(5123) <= not((layer0_outputs(5865)) or (layer0_outputs(6474)));
    outputs(5124) <= not(layer0_outputs(2983));
    outputs(5125) <= not(layer0_outputs(12026));
    outputs(5126) <= not((layer0_outputs(10218)) xor (layer0_outputs(324)));
    outputs(5127) <= not(layer0_outputs(12298)) or (layer0_outputs(3938));
    outputs(5128) <= (layer0_outputs(3049)) and not (layer0_outputs(7961));
    outputs(5129) <= layer0_outputs(7326);
    outputs(5130) <= not(layer0_outputs(12436));
    outputs(5131) <= layer0_outputs(152);
    outputs(5132) <= not(layer0_outputs(3261));
    outputs(5133) <= not((layer0_outputs(9380)) xor (layer0_outputs(10654)));
    outputs(5134) <= not((layer0_outputs(3043)) and (layer0_outputs(2492)));
    outputs(5135) <= (layer0_outputs(8617)) and not (layer0_outputs(16));
    outputs(5136) <= not((layer0_outputs(8603)) xor (layer0_outputs(391)));
    outputs(5137) <= not(layer0_outputs(4007));
    outputs(5138) <= not(layer0_outputs(11543));
    outputs(5139) <= not((layer0_outputs(3070)) xor (layer0_outputs(11406)));
    outputs(5140) <= layer0_outputs(3031);
    outputs(5141) <= not((layer0_outputs(1218)) and (layer0_outputs(4429)));
    outputs(5142) <= not(layer0_outputs(6877)) or (layer0_outputs(11734));
    outputs(5143) <= layer0_outputs(5558);
    outputs(5144) <= not(layer0_outputs(5181));
    outputs(5145) <= not((layer0_outputs(111)) xor (layer0_outputs(5917)));
    outputs(5146) <= (layer0_outputs(2215)) xor (layer0_outputs(8148));
    outputs(5147) <= not(layer0_outputs(11670)) or (layer0_outputs(7690));
    outputs(5148) <= (layer0_outputs(6020)) xor (layer0_outputs(3156));
    outputs(5149) <= (layer0_outputs(12013)) and not (layer0_outputs(3026));
    outputs(5150) <= layer0_outputs(11942);
    outputs(5151) <= layer0_outputs(4893);
    outputs(5152) <= not(layer0_outputs(4646));
    outputs(5153) <= layer0_outputs(3326);
    outputs(5154) <= not(layer0_outputs(12796));
    outputs(5155) <= not((layer0_outputs(10789)) or (layer0_outputs(7463)));
    outputs(5156) <= not((layer0_outputs(7529)) or (layer0_outputs(6856)));
    outputs(5157) <= layer0_outputs(4046);
    outputs(5158) <= (layer0_outputs(8402)) and (layer0_outputs(4672));
    outputs(5159) <= layer0_outputs(5842);
    outputs(5160) <= (layer0_outputs(8672)) and not (layer0_outputs(1877));
    outputs(5161) <= (layer0_outputs(4392)) and not (layer0_outputs(10732));
    outputs(5162) <= layer0_outputs(9835);
    outputs(5163) <= not(layer0_outputs(1099)) or (layer0_outputs(1597));
    outputs(5164) <= not(layer0_outputs(658));
    outputs(5165) <= not((layer0_outputs(8320)) or (layer0_outputs(9480)));
    outputs(5166) <= not((layer0_outputs(11790)) xor (layer0_outputs(7995)));
    outputs(5167) <= (layer0_outputs(12030)) and (layer0_outputs(8532));
    outputs(5168) <= not(layer0_outputs(1394));
    outputs(5169) <= layer0_outputs(6111);
    outputs(5170) <= not((layer0_outputs(8474)) xor (layer0_outputs(2242)));
    outputs(5171) <= layer0_outputs(8974);
    outputs(5172) <= layer0_outputs(7769);
    outputs(5173) <= layer0_outputs(5347);
    outputs(5174) <= not((layer0_outputs(8700)) xor (layer0_outputs(5523)));
    outputs(5175) <= not(layer0_outputs(966));
    outputs(5176) <= layer0_outputs(3767);
    outputs(5177) <= (layer0_outputs(2291)) and not (layer0_outputs(6495));
    outputs(5178) <= (layer0_outputs(2806)) xor (layer0_outputs(6095));
    outputs(5179) <= layer0_outputs(2165);
    outputs(5180) <= not((layer0_outputs(9908)) xor (layer0_outputs(8186)));
    outputs(5181) <= layer0_outputs(7019);
    outputs(5182) <= (layer0_outputs(12614)) and (layer0_outputs(2675));
    outputs(5183) <= not(layer0_outputs(3625));
    outputs(5184) <= (layer0_outputs(5719)) xor (layer0_outputs(1276));
    outputs(5185) <= not((layer0_outputs(1875)) xor (layer0_outputs(5843)));
    outputs(5186) <= (layer0_outputs(6149)) and not (layer0_outputs(1724));
    outputs(5187) <= layer0_outputs(6853);
    outputs(5188) <= not(layer0_outputs(8197)) or (layer0_outputs(1465));
    outputs(5189) <= not((layer0_outputs(1636)) or (layer0_outputs(4483)));
    outputs(5190) <= not(layer0_outputs(11056));
    outputs(5191) <= layer0_outputs(3219);
    outputs(5192) <= not(layer0_outputs(9960));
    outputs(5193) <= not(layer0_outputs(10944));
    outputs(5194) <= (layer0_outputs(344)) and not (layer0_outputs(1401));
    outputs(5195) <= not(layer0_outputs(3242));
    outputs(5196) <= layer0_outputs(8084);
    outputs(5197) <= not(layer0_outputs(3742));
    outputs(5198) <= not(layer0_outputs(1446)) or (layer0_outputs(4415));
    outputs(5199) <= not((layer0_outputs(1697)) xor (layer0_outputs(4708)));
    outputs(5200) <= not(layer0_outputs(5990));
    outputs(5201) <= (layer0_outputs(5387)) and (layer0_outputs(10562));
    outputs(5202) <= layer0_outputs(11836);
    outputs(5203) <= (layer0_outputs(996)) xor (layer0_outputs(4084));
    outputs(5204) <= layer0_outputs(3135);
    outputs(5205) <= layer0_outputs(8254);
    outputs(5206) <= not(layer0_outputs(9936));
    outputs(5207) <= '0';
    outputs(5208) <= layer0_outputs(8117);
    outputs(5209) <= (layer0_outputs(6013)) xor (layer0_outputs(1708));
    outputs(5210) <= layer0_outputs(6376);
    outputs(5211) <= not(layer0_outputs(8496));
    outputs(5212) <= not((layer0_outputs(3632)) xor (layer0_outputs(3589)));
    outputs(5213) <= not((layer0_outputs(10907)) or (layer0_outputs(8361)));
    outputs(5214) <= not(layer0_outputs(12749)) or (layer0_outputs(10797));
    outputs(5215) <= layer0_outputs(7591);
    outputs(5216) <= not((layer0_outputs(6129)) xor (layer0_outputs(4484)));
    outputs(5217) <= layer0_outputs(11856);
    outputs(5218) <= layer0_outputs(6827);
    outputs(5219) <= layer0_outputs(5519);
    outputs(5220) <= not(layer0_outputs(12781)) or (layer0_outputs(1948));
    outputs(5221) <= not(layer0_outputs(10987));
    outputs(5222) <= (layer0_outputs(3963)) xor (layer0_outputs(7100));
    outputs(5223) <= not(layer0_outputs(4303));
    outputs(5224) <= layer0_outputs(2172);
    outputs(5225) <= (layer0_outputs(7857)) and not (layer0_outputs(7070));
    outputs(5226) <= (layer0_outputs(12511)) xor (layer0_outputs(10568));
    outputs(5227) <= (layer0_outputs(10273)) xor (layer0_outputs(4186));
    outputs(5228) <= not((layer0_outputs(7805)) and (layer0_outputs(5221)));
    outputs(5229) <= not((layer0_outputs(4961)) xor (layer0_outputs(1730)));
    outputs(5230) <= layer0_outputs(124);
    outputs(5231) <= (layer0_outputs(9784)) and not (layer0_outputs(3805));
    outputs(5232) <= layer0_outputs(7061);
    outputs(5233) <= (layer0_outputs(7251)) xor (layer0_outputs(10248));
    outputs(5234) <= '1';
    outputs(5235) <= (layer0_outputs(1497)) xor (layer0_outputs(1534));
    outputs(5236) <= layer0_outputs(6844);
    outputs(5237) <= not(layer0_outputs(5600));
    outputs(5238) <= not(layer0_outputs(9722));
    outputs(5239) <= (layer0_outputs(4036)) and not (layer0_outputs(4638));
    outputs(5240) <= (layer0_outputs(4808)) xor (layer0_outputs(9842));
    outputs(5241) <= not((layer0_outputs(11329)) or (layer0_outputs(6664)));
    outputs(5242) <= layer0_outputs(3514);
    outputs(5243) <= (layer0_outputs(458)) or (layer0_outputs(11580));
    outputs(5244) <= (layer0_outputs(2132)) xor (layer0_outputs(1885));
    outputs(5245) <= layer0_outputs(1074);
    outputs(5246) <= not(layer0_outputs(3412)) or (layer0_outputs(12284));
    outputs(5247) <= not(layer0_outputs(8877));
    outputs(5248) <= not(layer0_outputs(10138));
    outputs(5249) <= not(layer0_outputs(12158));
    outputs(5250) <= (layer0_outputs(2354)) xor (layer0_outputs(8848));
    outputs(5251) <= layer0_outputs(7168);
    outputs(5252) <= not(layer0_outputs(3399)) or (layer0_outputs(7537));
    outputs(5253) <= not(layer0_outputs(7466)) or (layer0_outputs(12439));
    outputs(5254) <= (layer0_outputs(1546)) or (layer0_outputs(6835));
    outputs(5255) <= (layer0_outputs(5062)) and (layer0_outputs(6691));
    outputs(5256) <= not((layer0_outputs(6391)) xor (layer0_outputs(6504)));
    outputs(5257) <= (layer0_outputs(12306)) xor (layer0_outputs(11891));
    outputs(5258) <= not(layer0_outputs(5432));
    outputs(5259) <= not(layer0_outputs(3880));
    outputs(5260) <= layer0_outputs(7524);
    outputs(5261) <= layer0_outputs(5486);
    outputs(5262) <= layer0_outputs(9125);
    outputs(5263) <= not(layer0_outputs(4785));
    outputs(5264) <= not((layer0_outputs(7931)) xor (layer0_outputs(4820)));
    outputs(5265) <= (layer0_outputs(11112)) xor (layer0_outputs(5822));
    outputs(5266) <= (layer0_outputs(1158)) xor (layer0_outputs(1145));
    outputs(5267) <= (layer0_outputs(2918)) and (layer0_outputs(4736));
    outputs(5268) <= not((layer0_outputs(718)) or (layer0_outputs(9641)));
    outputs(5269) <= (layer0_outputs(9097)) and not (layer0_outputs(5089));
    outputs(5270) <= (layer0_outputs(5001)) and not (layer0_outputs(6966));
    outputs(5271) <= not(layer0_outputs(8189));
    outputs(5272) <= not(layer0_outputs(9292));
    outputs(5273) <= layer0_outputs(12415);
    outputs(5274) <= layer0_outputs(2625);
    outputs(5275) <= not(layer0_outputs(2420)) or (layer0_outputs(5999));
    outputs(5276) <= layer0_outputs(1110);
    outputs(5277) <= not(layer0_outputs(10325));
    outputs(5278) <= not((layer0_outputs(465)) xor (layer0_outputs(1978)));
    outputs(5279) <= (layer0_outputs(12577)) xor (layer0_outputs(2340));
    outputs(5280) <= (layer0_outputs(7321)) and (layer0_outputs(10745));
    outputs(5281) <= not(layer0_outputs(1863));
    outputs(5282) <= (layer0_outputs(4508)) xor (layer0_outputs(12513));
    outputs(5283) <= not((layer0_outputs(3703)) xor (layer0_outputs(7003)));
    outputs(5284) <= not(layer0_outputs(2743));
    outputs(5285) <= layer0_outputs(11527);
    outputs(5286) <= not((layer0_outputs(8260)) or (layer0_outputs(9775)));
    outputs(5287) <= not(layer0_outputs(6020));
    outputs(5288) <= not(layer0_outputs(11075));
    outputs(5289) <= not(layer0_outputs(1343)) or (layer0_outputs(9294));
    outputs(5290) <= layer0_outputs(9423);
    outputs(5291) <= (layer0_outputs(4874)) and not (layer0_outputs(864));
    outputs(5292) <= layer0_outputs(4004);
    outputs(5293) <= (layer0_outputs(1458)) and not (layer0_outputs(12743));
    outputs(5294) <= layer0_outputs(80);
    outputs(5295) <= layer0_outputs(11053);
    outputs(5296) <= (layer0_outputs(2973)) xor (layer0_outputs(2556));
    outputs(5297) <= not(layer0_outputs(367));
    outputs(5298) <= not((layer0_outputs(3227)) xor (layer0_outputs(9040)));
    outputs(5299) <= not(layer0_outputs(10342));
    outputs(5300) <= (layer0_outputs(12090)) and (layer0_outputs(36));
    outputs(5301) <= (layer0_outputs(8325)) xor (layer0_outputs(928));
    outputs(5302) <= (layer0_outputs(6624)) xor (layer0_outputs(4081));
    outputs(5303) <= not(layer0_outputs(311));
    outputs(5304) <= (layer0_outputs(3318)) and not (layer0_outputs(7667));
    outputs(5305) <= (layer0_outputs(12044)) xor (layer0_outputs(2048));
    outputs(5306) <= (layer0_outputs(9902)) or (layer0_outputs(7229));
    outputs(5307) <= not((layer0_outputs(9608)) or (layer0_outputs(1562)));
    outputs(5308) <= layer0_outputs(6637);
    outputs(5309) <= not(layer0_outputs(5473));
    outputs(5310) <= (layer0_outputs(912)) and not (layer0_outputs(138));
    outputs(5311) <= not(layer0_outputs(3408));
    outputs(5312) <= layer0_outputs(8488);
    outputs(5313) <= layer0_outputs(8126);
    outputs(5314) <= layer0_outputs(4184);
    outputs(5315) <= layer0_outputs(4541);
    outputs(5316) <= layer0_outputs(9695);
    outputs(5317) <= (layer0_outputs(6306)) and (layer0_outputs(11037));
    outputs(5318) <= (layer0_outputs(3306)) and (layer0_outputs(7661));
    outputs(5319) <= not(layer0_outputs(2555));
    outputs(5320) <= not(layer0_outputs(2848));
    outputs(5321) <= not(layer0_outputs(7488));
    outputs(5322) <= (layer0_outputs(12556)) and not (layer0_outputs(2677));
    outputs(5323) <= layer0_outputs(9553);
    outputs(5324) <= not(layer0_outputs(6971));
    outputs(5325) <= (layer0_outputs(1)) and not (layer0_outputs(6932));
    outputs(5326) <= not(layer0_outputs(5806));
    outputs(5327) <= layer0_outputs(3999);
    outputs(5328) <= (layer0_outputs(757)) and not (layer0_outputs(9538));
    outputs(5329) <= layer0_outputs(10128);
    outputs(5330) <= not((layer0_outputs(6694)) xor (layer0_outputs(2754)));
    outputs(5331) <= (layer0_outputs(9312)) and not (layer0_outputs(1154));
    outputs(5332) <= not(layer0_outputs(2277));
    outputs(5333) <= layer0_outputs(10212);
    outputs(5334) <= not(layer0_outputs(6480));
    outputs(5335) <= not((layer0_outputs(11954)) xor (layer0_outputs(3146)));
    outputs(5336) <= not(layer0_outputs(2440));
    outputs(5337) <= not(layer0_outputs(1014));
    outputs(5338) <= not(layer0_outputs(388));
    outputs(5339) <= layer0_outputs(2042);
    outputs(5340) <= layer0_outputs(5307);
    outputs(5341) <= not(layer0_outputs(12479));
    outputs(5342) <= not((layer0_outputs(4337)) xor (layer0_outputs(6252)));
    outputs(5343) <= not(layer0_outputs(754));
    outputs(5344) <= (layer0_outputs(1919)) or (layer0_outputs(4937));
    outputs(5345) <= not(layer0_outputs(4962));
    outputs(5346) <= layer0_outputs(11780);
    outputs(5347) <= not((layer0_outputs(2463)) or (layer0_outputs(899)));
    outputs(5348) <= (layer0_outputs(8767)) and not (layer0_outputs(7667));
    outputs(5349) <= layer0_outputs(4574);
    outputs(5350) <= not(layer0_outputs(1056)) or (layer0_outputs(11836));
    outputs(5351) <= not(layer0_outputs(583));
    outputs(5352) <= not(layer0_outputs(4252));
    outputs(5353) <= not((layer0_outputs(10428)) and (layer0_outputs(12160)));
    outputs(5354) <= layer0_outputs(5514);
    outputs(5355) <= (layer0_outputs(4631)) or (layer0_outputs(2699));
    outputs(5356) <= not((layer0_outputs(7444)) or (layer0_outputs(10889)));
    outputs(5357) <= not((layer0_outputs(154)) xor (layer0_outputs(2701)));
    outputs(5358) <= layer0_outputs(11378);
    outputs(5359) <= (layer0_outputs(8286)) or (layer0_outputs(3635));
    outputs(5360) <= not(layer0_outputs(11067));
    outputs(5361) <= not(layer0_outputs(5245));
    outputs(5362) <= layer0_outputs(1991);
    outputs(5363) <= not((layer0_outputs(2843)) xor (layer0_outputs(2980)));
    outputs(5364) <= (layer0_outputs(12463)) and not (layer0_outputs(356));
    outputs(5365) <= not(layer0_outputs(10595));
    outputs(5366) <= (layer0_outputs(8270)) or (layer0_outputs(9440));
    outputs(5367) <= not((layer0_outputs(4687)) xor (layer0_outputs(3863)));
    outputs(5368) <= not((layer0_outputs(12214)) or (layer0_outputs(2702)));
    outputs(5369) <= layer0_outputs(4248);
    outputs(5370) <= (layer0_outputs(12441)) xor (layer0_outputs(4822));
    outputs(5371) <= layer0_outputs(622);
    outputs(5372) <= not(layer0_outputs(981)) or (layer0_outputs(8003));
    outputs(5373) <= not(layer0_outputs(9364));
    outputs(5374) <= not(layer0_outputs(1474));
    outputs(5375) <= (layer0_outputs(10936)) and (layer0_outputs(2093));
    outputs(5376) <= layer0_outputs(4844);
    outputs(5377) <= (layer0_outputs(7541)) and not (layer0_outputs(2931));
    outputs(5378) <= not((layer0_outputs(10332)) and (layer0_outputs(4909)));
    outputs(5379) <= not(layer0_outputs(1391));
    outputs(5380) <= (layer0_outputs(12003)) and not (layer0_outputs(8287));
    outputs(5381) <= not((layer0_outputs(3448)) and (layer0_outputs(11287)));
    outputs(5382) <= not(layer0_outputs(11160));
    outputs(5383) <= not((layer0_outputs(8256)) xor (layer0_outputs(947)));
    outputs(5384) <= not((layer0_outputs(10887)) xor (layer0_outputs(11996)));
    outputs(5385) <= (layer0_outputs(9478)) and not (layer0_outputs(4525));
    outputs(5386) <= (layer0_outputs(3458)) xor (layer0_outputs(4276));
    outputs(5387) <= not((layer0_outputs(7295)) and (layer0_outputs(12254)));
    outputs(5388) <= not((layer0_outputs(1475)) xor (layer0_outputs(12316)));
    outputs(5389) <= (layer0_outputs(11531)) or (layer0_outputs(12681));
    outputs(5390) <= layer0_outputs(7954);
    outputs(5391) <= '1';
    outputs(5392) <= (layer0_outputs(10509)) and (layer0_outputs(8022));
    outputs(5393) <= layer0_outputs(10638);
    outputs(5394) <= (layer0_outputs(9840)) xor (layer0_outputs(4459));
    outputs(5395) <= (layer0_outputs(2297)) and not (layer0_outputs(496));
    outputs(5396) <= (layer0_outputs(9521)) and (layer0_outputs(1029));
    outputs(5397) <= not(layer0_outputs(10621));
    outputs(5398) <= layer0_outputs(5820);
    outputs(5399) <= (layer0_outputs(8901)) and not (layer0_outputs(4417));
    outputs(5400) <= layer0_outputs(11565);
    outputs(5401) <= not(layer0_outputs(8131)) or (layer0_outputs(9922));
    outputs(5402) <= (layer0_outputs(3228)) or (layer0_outputs(4302));
    outputs(5403) <= not(layer0_outputs(10466));
    outputs(5404) <= layer0_outputs(2757);
    outputs(5405) <= layer0_outputs(3549);
    outputs(5406) <= not(layer0_outputs(7564));
    outputs(5407) <= not(layer0_outputs(7406)) or (layer0_outputs(8685));
    outputs(5408) <= not(layer0_outputs(2835));
    outputs(5409) <= layer0_outputs(5702);
    outputs(5410) <= not(layer0_outputs(10889));
    outputs(5411) <= layer0_outputs(5762);
    outputs(5412) <= layer0_outputs(2657);
    outputs(5413) <= (layer0_outputs(3009)) and not (layer0_outputs(4213));
    outputs(5414) <= layer0_outputs(8091);
    outputs(5415) <= (layer0_outputs(6176)) and not (layer0_outputs(3580));
    outputs(5416) <= (layer0_outputs(7956)) or (layer0_outputs(5595));
    outputs(5417) <= layer0_outputs(5529);
    outputs(5418) <= not(layer0_outputs(4416));
    outputs(5419) <= layer0_outputs(6311);
    outputs(5420) <= not(layer0_outputs(5406));
    outputs(5421) <= layer0_outputs(11540);
    outputs(5422) <= layer0_outputs(1125);
    outputs(5423) <= (layer0_outputs(1194)) and not (layer0_outputs(11593));
    outputs(5424) <= layer0_outputs(11553);
    outputs(5425) <= not(layer0_outputs(8763));
    outputs(5426) <= layer0_outputs(7020);
    outputs(5427) <= layer0_outputs(2396);
    outputs(5428) <= layer0_outputs(4846);
    outputs(5429) <= (layer0_outputs(10317)) or (layer0_outputs(5069));
    outputs(5430) <= layer0_outputs(5238);
    outputs(5431) <= (layer0_outputs(4799)) and not (layer0_outputs(3726));
    outputs(5432) <= (layer0_outputs(463)) or (layer0_outputs(5664));
    outputs(5433) <= not(layer0_outputs(3623));
    outputs(5434) <= (layer0_outputs(12212)) and not (layer0_outputs(10629));
    outputs(5435) <= (layer0_outputs(7201)) and not (layer0_outputs(11276));
    outputs(5436) <= layer0_outputs(3853);
    outputs(5437) <= (layer0_outputs(357)) and not (layer0_outputs(6580));
    outputs(5438) <= not((layer0_outputs(5271)) or (layer0_outputs(2316)));
    outputs(5439) <= (layer0_outputs(939)) and not (layer0_outputs(10772));
    outputs(5440) <= not(layer0_outputs(2688));
    outputs(5441) <= (layer0_outputs(10108)) xor (layer0_outputs(10430));
    outputs(5442) <= not(layer0_outputs(10985));
    outputs(5443) <= not(layer0_outputs(4237));
    outputs(5444) <= not(layer0_outputs(1808));
    outputs(5445) <= (layer0_outputs(8973)) xor (layer0_outputs(1453));
    outputs(5446) <= not((layer0_outputs(12156)) xor (layer0_outputs(9136)));
    outputs(5447) <= not(layer0_outputs(6959));
    outputs(5448) <= not((layer0_outputs(8710)) and (layer0_outputs(1184)));
    outputs(5449) <= (layer0_outputs(10646)) xor (layer0_outputs(200));
    outputs(5450) <= (layer0_outputs(1638)) xor (layer0_outputs(11122));
    outputs(5451) <= not((layer0_outputs(8084)) xor (layer0_outputs(1592)));
    outputs(5452) <= not(layer0_outputs(1123));
    outputs(5453) <= (layer0_outputs(2122)) or (layer0_outputs(11537));
    outputs(5454) <= not((layer0_outputs(1061)) or (layer0_outputs(10356)));
    outputs(5455) <= layer0_outputs(5162);
    outputs(5456) <= layer0_outputs(11931);
    outputs(5457) <= not(layer0_outputs(9262)) or (layer0_outputs(5102));
    outputs(5458) <= layer0_outputs(11494);
    outputs(5459) <= not((layer0_outputs(7966)) xor (layer0_outputs(3181)));
    outputs(5460) <= not((layer0_outputs(7189)) or (layer0_outputs(5641)));
    outputs(5461) <= not(layer0_outputs(2966)) or (layer0_outputs(8799));
    outputs(5462) <= not((layer0_outputs(6007)) or (layer0_outputs(12204)));
    outputs(5463) <= (layer0_outputs(1912)) xor (layer0_outputs(10411));
    outputs(5464) <= (layer0_outputs(764)) and (layer0_outputs(6345));
    outputs(5465) <= layer0_outputs(2452);
    outputs(5466) <= not((layer0_outputs(4459)) xor (layer0_outputs(590)));
    outputs(5467) <= (layer0_outputs(6144)) or (layer0_outputs(1555));
    outputs(5468) <= not((layer0_outputs(11218)) xor (layer0_outputs(689)));
    outputs(5469) <= layer0_outputs(2188);
    outputs(5470) <= layer0_outputs(11196);
    outputs(5471) <= (layer0_outputs(3669)) and not (layer0_outputs(10898));
    outputs(5472) <= (layer0_outputs(11024)) and (layer0_outputs(1051));
    outputs(5473) <= not((layer0_outputs(10812)) xor (layer0_outputs(4284)));
    outputs(5474) <= '1';
    outputs(5475) <= layer0_outputs(4779);
    outputs(5476) <= not(layer0_outputs(4520));
    outputs(5477) <= not((layer0_outputs(3967)) xor (layer0_outputs(5761)));
    outputs(5478) <= layer0_outputs(7285);
    outputs(5479) <= (layer0_outputs(5027)) and not (layer0_outputs(1246));
    outputs(5480) <= not(layer0_outputs(749));
    outputs(5481) <= layer0_outputs(5740);
    outputs(5482) <= not((layer0_outputs(12134)) and (layer0_outputs(2941)));
    outputs(5483) <= layer0_outputs(8327);
    outputs(5484) <= layer0_outputs(2247);
    outputs(5485) <= (layer0_outputs(7658)) or (layer0_outputs(10109));
    outputs(5486) <= (layer0_outputs(332)) xor (layer0_outputs(2384));
    outputs(5487) <= layer0_outputs(5436);
    outputs(5488) <= not(layer0_outputs(1097)) or (layer0_outputs(10979));
    outputs(5489) <= (layer0_outputs(7908)) xor (layer0_outputs(1975));
    outputs(5490) <= not((layer0_outputs(6450)) xor (layer0_outputs(12675)));
    outputs(5491) <= not(layer0_outputs(9682));
    outputs(5492) <= not((layer0_outputs(9576)) xor (layer0_outputs(3534)));
    outputs(5493) <= (layer0_outputs(7788)) xor (layer0_outputs(1383));
    outputs(5494) <= (layer0_outputs(9065)) and not (layer0_outputs(8338));
    outputs(5495) <= (layer0_outputs(6449)) and (layer0_outputs(352));
    outputs(5496) <= not(layer0_outputs(12447)) or (layer0_outputs(3402));
    outputs(5497) <= not(layer0_outputs(7734));
    outputs(5498) <= (layer0_outputs(5379)) xor (layer0_outputs(5267));
    outputs(5499) <= layer0_outputs(6764);
    outputs(5500) <= not(layer0_outputs(6478));
    outputs(5501) <= not((layer0_outputs(5110)) xor (layer0_outputs(12025)));
    outputs(5502) <= not(layer0_outputs(5615));
    outputs(5503) <= (layer0_outputs(6429)) and (layer0_outputs(8377));
    outputs(5504) <= not(layer0_outputs(4911));
    outputs(5505) <= (layer0_outputs(1550)) xor (layer0_outputs(2515));
    outputs(5506) <= not(layer0_outputs(11763));
    outputs(5507) <= (layer0_outputs(11257)) and (layer0_outputs(5103));
    outputs(5508) <= not((layer0_outputs(1848)) or (layer0_outputs(2129)));
    outputs(5509) <= (layer0_outputs(6655)) xor (layer0_outputs(3802));
    outputs(5510) <= (layer0_outputs(4127)) xor (layer0_outputs(9675));
    outputs(5511) <= (layer0_outputs(11049)) xor (layer0_outputs(7135));
    outputs(5512) <= (layer0_outputs(4024)) and (layer0_outputs(10613));
    outputs(5513) <= not((layer0_outputs(9461)) xor (layer0_outputs(12535)));
    outputs(5514) <= (layer0_outputs(8251)) and not (layer0_outputs(1526));
    outputs(5515) <= not(layer0_outputs(9439));
    outputs(5516) <= layer0_outputs(6484);
    outputs(5517) <= layer0_outputs(6251);
    outputs(5518) <= (layer0_outputs(11237)) and (layer0_outputs(8588));
    outputs(5519) <= not((layer0_outputs(9135)) or (layer0_outputs(10472)));
    outputs(5520) <= (layer0_outputs(9987)) and (layer0_outputs(2414));
    outputs(5521) <= layer0_outputs(8972);
    outputs(5522) <= not((layer0_outputs(2427)) and (layer0_outputs(11245)));
    outputs(5523) <= not((layer0_outputs(1323)) xor (layer0_outputs(9647)));
    outputs(5524) <= not(layer0_outputs(10972));
    outputs(5525) <= (layer0_outputs(9524)) xor (layer0_outputs(7284));
    outputs(5526) <= not(layer0_outputs(2519));
    outputs(5527) <= layer0_outputs(2684);
    outputs(5528) <= (layer0_outputs(7635)) and not (layer0_outputs(2079));
    outputs(5529) <= not(layer0_outputs(8096));
    outputs(5530) <= not((layer0_outputs(788)) or (layer0_outputs(5896)));
    outputs(5531) <= not((layer0_outputs(2818)) xor (layer0_outputs(12034)));
    outputs(5532) <= not((layer0_outputs(3820)) xor (layer0_outputs(11590)));
    outputs(5533) <= (layer0_outputs(10698)) xor (layer0_outputs(10229));
    outputs(5534) <= (layer0_outputs(7649)) xor (layer0_outputs(11626));
    outputs(5535) <= not((layer0_outputs(8547)) xor (layer0_outputs(853)));
    outputs(5536) <= layer0_outputs(2227);
    outputs(5537) <= not(layer0_outputs(2533));
    outputs(5538) <= (layer0_outputs(10655)) xor (layer0_outputs(1356));
    outputs(5539) <= not(layer0_outputs(10143));
    outputs(5540) <= layer0_outputs(6309);
    outputs(5541) <= not(layer0_outputs(1052));
    outputs(5542) <= not(layer0_outputs(11621));
    outputs(5543) <= layer0_outputs(9537);
    outputs(5544) <= layer0_outputs(5256);
    outputs(5545) <= layer0_outputs(12679);
    outputs(5546) <= layer0_outputs(2107);
    outputs(5547) <= layer0_outputs(3302);
    outputs(5548) <= not((layer0_outputs(7251)) xor (layer0_outputs(5131)));
    outputs(5549) <= not(layer0_outputs(8461));
    outputs(5550) <= not(layer0_outputs(1616));
    outputs(5551) <= not(layer0_outputs(5255));
    outputs(5552) <= (layer0_outputs(9851)) xor (layer0_outputs(11197));
    outputs(5553) <= not(layer0_outputs(6043));
    outputs(5554) <= (layer0_outputs(8721)) and (layer0_outputs(5124));
    outputs(5555) <= (layer0_outputs(7883)) xor (layer0_outputs(11029));
    outputs(5556) <= layer0_outputs(8031);
    outputs(5557) <= layer0_outputs(1132);
    outputs(5558) <= not(layer0_outputs(624));
    outputs(5559) <= not(layer0_outputs(3138));
    outputs(5560) <= (layer0_outputs(7225)) xor (layer0_outputs(1111));
    outputs(5561) <= (layer0_outputs(3271)) and (layer0_outputs(4477));
    outputs(5562) <= not(layer0_outputs(12333)) or (layer0_outputs(11556));
    outputs(5563) <= layer0_outputs(619);
    outputs(5564) <= not(layer0_outputs(11769));
    outputs(5565) <= (layer0_outputs(1134)) xor (layer0_outputs(5685));
    outputs(5566) <= layer0_outputs(6376);
    outputs(5567) <= (layer0_outputs(695)) xor (layer0_outputs(8164));
    outputs(5568) <= (layer0_outputs(2838)) xor (layer0_outputs(7561));
    outputs(5569) <= not(layer0_outputs(807));
    outputs(5570) <= not(layer0_outputs(7970));
    outputs(5571) <= not(layer0_outputs(12726));
    outputs(5572) <= not((layer0_outputs(3417)) xor (layer0_outputs(345)));
    outputs(5573) <= not(layer0_outputs(6937));
    outputs(5574) <= not(layer0_outputs(11990));
    outputs(5575) <= (layer0_outputs(6091)) and not (layer0_outputs(5921));
    outputs(5576) <= layer0_outputs(7309);
    outputs(5577) <= not(layer0_outputs(6919));
    outputs(5578) <= not(layer0_outputs(8307));
    outputs(5579) <= not((layer0_outputs(4752)) or (layer0_outputs(12281)));
    outputs(5580) <= (layer0_outputs(2763)) and (layer0_outputs(11018));
    outputs(5581) <= layer0_outputs(136);
    outputs(5582) <= (layer0_outputs(1249)) xor (layer0_outputs(12689));
    outputs(5583) <= not(layer0_outputs(8751));
    outputs(5584) <= not(layer0_outputs(8397));
    outputs(5585) <= not(layer0_outputs(6887));
    outputs(5586) <= not(layer0_outputs(2736));
    outputs(5587) <= not(layer0_outputs(3717)) or (layer0_outputs(6541));
    outputs(5588) <= layer0_outputs(2403);
    outputs(5589) <= layer0_outputs(705);
    outputs(5590) <= (layer0_outputs(343)) and (layer0_outputs(3547));
    outputs(5591) <= not((layer0_outputs(11518)) xor (layer0_outputs(3320)));
    outputs(5592) <= not(layer0_outputs(2136)) or (layer0_outputs(1519));
    outputs(5593) <= not(layer0_outputs(5647));
    outputs(5594) <= not((layer0_outputs(6301)) or (layer0_outputs(6387)));
    outputs(5595) <= not((layer0_outputs(796)) and (layer0_outputs(11065)));
    outputs(5596) <= not(layer0_outputs(8846)) or (layer0_outputs(2841));
    outputs(5597) <= (layer0_outputs(1121)) xor (layer0_outputs(11528));
    outputs(5598) <= not((layer0_outputs(4628)) or (layer0_outputs(9415)));
    outputs(5599) <= not((layer0_outputs(7898)) xor (layer0_outputs(11934)));
    outputs(5600) <= layer0_outputs(2649);
    outputs(5601) <= (layer0_outputs(10400)) xor (layer0_outputs(1390));
    outputs(5602) <= (layer0_outputs(1292)) and not (layer0_outputs(9833));
    outputs(5603) <= not(layer0_outputs(1669));
    outputs(5604) <= (layer0_outputs(9121)) xor (layer0_outputs(6885));
    outputs(5605) <= layer0_outputs(9875);
    outputs(5606) <= (layer0_outputs(3011)) xor (layer0_outputs(8988));
    outputs(5607) <= layer0_outputs(5842);
    outputs(5608) <= (layer0_outputs(2388)) xor (layer0_outputs(8367));
    outputs(5609) <= not(layer0_outputs(2369));
    outputs(5610) <= not((layer0_outputs(3361)) or (layer0_outputs(5041)));
    outputs(5611) <= layer0_outputs(6682);
    outputs(5612) <= not(layer0_outputs(1688));
    outputs(5613) <= layer0_outputs(238);
    outputs(5614) <= (layer0_outputs(10961)) and not (layer0_outputs(7000));
    outputs(5615) <= layer0_outputs(386);
    outputs(5616) <= not(layer0_outputs(3386));
    outputs(5617) <= not(layer0_outputs(7298));
    outputs(5618) <= (layer0_outputs(9851)) and not (layer0_outputs(9282));
    outputs(5619) <= not(layer0_outputs(2833));
    outputs(5620) <= not(layer0_outputs(6892));
    outputs(5621) <= layer0_outputs(12779);
    outputs(5622) <= (layer0_outputs(3210)) and not (layer0_outputs(9341));
    outputs(5623) <= (layer0_outputs(2222)) xor (layer0_outputs(1090));
    outputs(5624) <= not(layer0_outputs(5255));
    outputs(5625) <= layer0_outputs(8625);
    outputs(5626) <= (layer0_outputs(10096)) xor (layer0_outputs(8216));
    outputs(5627) <= (layer0_outputs(11562)) xor (layer0_outputs(3785));
    outputs(5628) <= (layer0_outputs(795)) and not (layer0_outputs(11572));
    outputs(5629) <= layer0_outputs(147);
    outputs(5630) <= (layer0_outputs(959)) and (layer0_outputs(11074));
    outputs(5631) <= not((layer0_outputs(5815)) xor (layer0_outputs(6787)));
    outputs(5632) <= not((layer0_outputs(4245)) xor (layer0_outputs(12697)));
    outputs(5633) <= layer0_outputs(7044);
    outputs(5634) <= not((layer0_outputs(2320)) or (layer0_outputs(8930)));
    outputs(5635) <= not(layer0_outputs(3332));
    outputs(5636) <= layer0_outputs(5305);
    outputs(5637) <= not(layer0_outputs(3690));
    outputs(5638) <= layer0_outputs(10405);
    outputs(5639) <= not(layer0_outputs(1057)) or (layer0_outputs(7182));
    outputs(5640) <= layer0_outputs(7368);
    outputs(5641) <= not(layer0_outputs(10341));
    outputs(5642) <= not(layer0_outputs(5966));
    outputs(5643) <= layer0_outputs(3253);
    outputs(5644) <= not(layer0_outputs(6008));
    outputs(5645) <= layer0_outputs(2723);
    outputs(5646) <= layer0_outputs(9328);
    outputs(5647) <= (layer0_outputs(7805)) and not (layer0_outputs(1048));
    outputs(5648) <= layer0_outputs(28);
    outputs(5649) <= layer0_outputs(5135);
    outputs(5650) <= layer0_outputs(8944);
    outputs(5651) <= not((layer0_outputs(645)) xor (layer0_outputs(4840)));
    outputs(5652) <= not((layer0_outputs(5864)) or (layer0_outputs(10452)));
    outputs(5653) <= not(layer0_outputs(7981));
    outputs(5654) <= layer0_outputs(10825);
    outputs(5655) <= (layer0_outputs(9501)) and not (layer0_outputs(6374));
    outputs(5656) <= not(layer0_outputs(4918));
    outputs(5657) <= layer0_outputs(11552);
    outputs(5658) <= (layer0_outputs(10856)) xor (layer0_outputs(64));
    outputs(5659) <= layer0_outputs(10704);
    outputs(5660) <= not(layer0_outputs(1687));
    outputs(5661) <= (layer0_outputs(3020)) xor (layer0_outputs(8330));
    outputs(5662) <= (layer0_outputs(2897)) and (layer0_outputs(903));
    outputs(5663) <= layer0_outputs(409);
    outputs(5664) <= (layer0_outputs(9769)) xor (layer0_outputs(1371));
    outputs(5665) <= '1';
    outputs(5666) <= (layer0_outputs(3516)) and (layer0_outputs(7898));
    outputs(5667) <= '0';
    outputs(5668) <= (layer0_outputs(6509)) xor (layer0_outputs(3744));
    outputs(5669) <= (layer0_outputs(4981)) and not (layer0_outputs(4119));
    outputs(5670) <= not((layer0_outputs(3556)) xor (layer0_outputs(1887)));
    outputs(5671) <= not((layer0_outputs(11057)) and (layer0_outputs(11865)));
    outputs(5672) <= not(layer0_outputs(342));
    outputs(5673) <= not((layer0_outputs(10369)) or (layer0_outputs(10733)));
    outputs(5674) <= not(layer0_outputs(5186));
    outputs(5675) <= not(layer0_outputs(823));
    outputs(5676) <= layer0_outputs(9250);
    outputs(5677) <= not((layer0_outputs(10647)) or (layer0_outputs(12772)));
    outputs(5678) <= not((layer0_outputs(1797)) or (layer0_outputs(6062)));
    outputs(5679) <= not((layer0_outputs(3375)) or (layer0_outputs(6077)));
    outputs(5680) <= not((layer0_outputs(7902)) xor (layer0_outputs(5781)));
    outputs(5681) <= not(layer0_outputs(10899)) or (layer0_outputs(11685));
    outputs(5682) <= not(layer0_outputs(8199));
    outputs(5683) <= not((layer0_outputs(7283)) xor (layer0_outputs(8490)));
    outputs(5684) <= layer0_outputs(6240);
    outputs(5685) <= not(layer0_outputs(9005));
    outputs(5686) <= not((layer0_outputs(711)) xor (layer0_outputs(5421)));
    outputs(5687) <= not((layer0_outputs(8198)) or (layer0_outputs(6136)));
    outputs(5688) <= layer0_outputs(910);
    outputs(5689) <= not(layer0_outputs(10034));
    outputs(5690) <= not(layer0_outputs(4644));
    outputs(5691) <= (layer0_outputs(12509)) and (layer0_outputs(440));
    outputs(5692) <= layer0_outputs(11042);
    outputs(5693) <= (layer0_outputs(11224)) and not (layer0_outputs(2541));
    outputs(5694) <= (layer0_outputs(11334)) and not (layer0_outputs(11654));
    outputs(5695) <= (layer0_outputs(5474)) and (layer0_outputs(12388));
    outputs(5696) <= not(layer0_outputs(11682));
    outputs(5697) <= not(layer0_outputs(8094));
    outputs(5698) <= (layer0_outputs(2284)) and not (layer0_outputs(7342));
    outputs(5699) <= layer0_outputs(6808);
    outputs(5700) <= not((layer0_outputs(12347)) and (layer0_outputs(2081)));
    outputs(5701) <= not((layer0_outputs(12650)) and (layer0_outputs(11332)));
    outputs(5702) <= not((layer0_outputs(4399)) xor (layer0_outputs(4380)));
    outputs(5703) <= (layer0_outputs(7580)) and (layer0_outputs(11423));
    outputs(5704) <= not(layer0_outputs(4332));
    outputs(5705) <= not(layer0_outputs(1339));
    outputs(5706) <= not((layer0_outputs(9495)) xor (layer0_outputs(9533)));
    outputs(5707) <= not((layer0_outputs(2422)) or (layer0_outputs(12427)));
    outputs(5708) <= not((layer0_outputs(3035)) or (layer0_outputs(12311)));
    outputs(5709) <= layer0_outputs(3186);
    outputs(5710) <= (layer0_outputs(6266)) and not (layer0_outputs(7923));
    outputs(5711) <= not(layer0_outputs(1496)) or (layer0_outputs(11786));
    outputs(5712) <= (layer0_outputs(4958)) xor (layer0_outputs(8518));
    outputs(5713) <= layer0_outputs(11225);
    outputs(5714) <= (layer0_outputs(12104)) and not (layer0_outputs(11206));
    outputs(5715) <= layer0_outputs(7721);
    outputs(5716) <= layer0_outputs(9223);
    outputs(5717) <= not(layer0_outputs(4280));
    outputs(5718) <= layer0_outputs(8823);
    outputs(5719) <= not(layer0_outputs(3873));
    outputs(5720) <= not(layer0_outputs(901));
    outputs(5721) <= not((layer0_outputs(7820)) xor (layer0_outputs(830)));
    outputs(5722) <= not((layer0_outputs(10571)) xor (layer0_outputs(1164)));
    outputs(5723) <= not((layer0_outputs(5085)) or (layer0_outputs(10609)));
    outputs(5724) <= not(layer0_outputs(7843));
    outputs(5725) <= not(layer0_outputs(11660));
    outputs(5726) <= layer0_outputs(360);
    outputs(5727) <= layer0_outputs(10009);
    outputs(5728) <= not(layer0_outputs(280));
    outputs(5729) <= not((layer0_outputs(1643)) xor (layer0_outputs(2535)));
    outputs(5730) <= not((layer0_outputs(9198)) xor (layer0_outputs(10664)));
    outputs(5731) <= not(layer0_outputs(5461));
    outputs(5732) <= not(layer0_outputs(10474));
    outputs(5733) <= not((layer0_outputs(5571)) xor (layer0_outputs(6120)));
    outputs(5734) <= layer0_outputs(1034);
    outputs(5735) <= layer0_outputs(9570);
    outputs(5736) <= not(layer0_outputs(12149));
    outputs(5737) <= (layer0_outputs(4588)) xor (layer0_outputs(1656));
    outputs(5738) <= not(layer0_outputs(2054)) or (layer0_outputs(4797));
    outputs(5739) <= layer0_outputs(8373);
    outputs(5740) <= layer0_outputs(8901);
    outputs(5741) <= not(layer0_outputs(3905));
    outputs(5742) <= layer0_outputs(6834);
    outputs(5743) <= not(layer0_outputs(9264));
    outputs(5744) <= not(layer0_outputs(11290));
    outputs(5745) <= layer0_outputs(561);
    outputs(5746) <= not(layer0_outputs(2183));
    outputs(5747) <= (layer0_outputs(8952)) and not (layer0_outputs(8023));
    outputs(5748) <= not((layer0_outputs(5592)) xor (layer0_outputs(1495)));
    outputs(5749) <= layer0_outputs(3816);
    outputs(5750) <= (layer0_outputs(2583)) and not (layer0_outputs(1769));
    outputs(5751) <= (layer0_outputs(3759)) xor (layer0_outputs(4308));
    outputs(5752) <= (layer0_outputs(12719)) and (layer0_outputs(7570));
    outputs(5753) <= layer0_outputs(1426);
    outputs(5754) <= layer0_outputs(7051);
    outputs(5755) <= layer0_outputs(266);
    outputs(5756) <= layer0_outputs(11362);
    outputs(5757) <= not(layer0_outputs(11991));
    outputs(5758) <= not((layer0_outputs(11263)) xor (layer0_outputs(11005)));
    outputs(5759) <= not(layer0_outputs(1924));
    outputs(5760) <= not(layer0_outputs(4774)) or (layer0_outputs(10529));
    outputs(5761) <= layer0_outputs(6863);
    outputs(5762) <= not(layer0_outputs(6492));
    outputs(5763) <= (layer0_outputs(1111)) xor (layer0_outputs(5494));
    outputs(5764) <= layer0_outputs(10966);
    outputs(5765) <= not(layer0_outputs(7824));
    outputs(5766) <= not(layer0_outputs(11039));
    outputs(5767) <= not(layer0_outputs(4291));
    outputs(5768) <= not((layer0_outputs(5847)) xor (layer0_outputs(8273)));
    outputs(5769) <= not((layer0_outputs(5371)) xor (layer0_outputs(12785)));
    outputs(5770) <= layer0_outputs(10246);
    outputs(5771) <= (layer0_outputs(8707)) xor (layer0_outputs(7649));
    outputs(5772) <= layer0_outputs(8144);
    outputs(5773) <= layer0_outputs(10801);
    outputs(5774) <= not(layer0_outputs(10011));
    outputs(5775) <= not((layer0_outputs(2857)) or (layer0_outputs(7525)));
    outputs(5776) <= not(layer0_outputs(578));
    outputs(5777) <= not(layer0_outputs(10330));
    outputs(5778) <= not(layer0_outputs(9482));
    outputs(5779) <= not((layer0_outputs(11452)) xor (layer0_outputs(11891)));
    outputs(5780) <= layer0_outputs(647);
    outputs(5781) <= not(layer0_outputs(709)) or (layer0_outputs(11215));
    outputs(5782) <= layer0_outputs(12428);
    outputs(5783) <= layer0_outputs(6780);
    outputs(5784) <= not((layer0_outputs(2478)) xor (layer0_outputs(1859)));
    outputs(5785) <= (layer0_outputs(12399)) and not (layer0_outputs(7823));
    outputs(5786) <= (layer0_outputs(6523)) and not (layer0_outputs(4947));
    outputs(5787) <= (layer0_outputs(5481)) and not (layer0_outputs(7536));
    outputs(5788) <= not((layer0_outputs(8621)) and (layer0_outputs(4744)));
    outputs(5789) <= layer0_outputs(12631);
    outputs(5790) <= layer0_outputs(126);
    outputs(5791) <= (layer0_outputs(2721)) xor (layer0_outputs(1402));
    outputs(5792) <= layer0_outputs(12098);
    outputs(5793) <= not(layer0_outputs(9462));
    outputs(5794) <= (layer0_outputs(7199)) or (layer0_outputs(7140));
    outputs(5795) <= (layer0_outputs(1271)) xor (layer0_outputs(3759));
    outputs(5796) <= not(layer0_outputs(10378));
    outputs(5797) <= layer0_outputs(6900);
    outputs(5798) <= layer0_outputs(7256);
    outputs(5799) <= not((layer0_outputs(8825)) xor (layer0_outputs(8420)));
    outputs(5800) <= not(layer0_outputs(1463));
    outputs(5801) <= not(layer0_outputs(5028));
    outputs(5802) <= not(layer0_outputs(8277));
    outputs(5803) <= not(layer0_outputs(7630));
    outputs(5804) <= layer0_outputs(353);
    outputs(5805) <= not(layer0_outputs(9845));
    outputs(5806) <= not((layer0_outputs(5406)) or (layer0_outputs(5242)));
    outputs(5807) <= (layer0_outputs(4058)) xor (layer0_outputs(4359));
    outputs(5808) <= (layer0_outputs(4600)) xor (layer0_outputs(3831));
    outputs(5809) <= not((layer0_outputs(4550)) xor (layer0_outputs(6779)));
    outputs(5810) <= (layer0_outputs(10387)) and not (layer0_outputs(10142));
    outputs(5811) <= not(layer0_outputs(12698)) or (layer0_outputs(1592));
    outputs(5812) <= not(layer0_outputs(8384));
    outputs(5813) <= (layer0_outputs(1987)) and not (layer0_outputs(12300));
    outputs(5814) <= not((layer0_outputs(6603)) or (layer0_outputs(8089)));
    outputs(5815) <= not(layer0_outputs(228));
    outputs(5816) <= not(layer0_outputs(12627)) or (layer0_outputs(12647));
    outputs(5817) <= (layer0_outputs(7632)) xor (layer0_outputs(10933));
    outputs(5818) <= not(layer0_outputs(3936)) or (layer0_outputs(920));
    outputs(5819) <= (layer0_outputs(5101)) and not (layer0_outputs(2402));
    outputs(5820) <= layer0_outputs(8254);
    outputs(5821) <= not(layer0_outputs(7968));
    outputs(5822) <= (layer0_outputs(11450)) and not (layer0_outputs(9247));
    outputs(5823) <= (layer0_outputs(4886)) and not (layer0_outputs(4556));
    outputs(5824) <= not(layer0_outputs(10998));
    outputs(5825) <= not((layer0_outputs(2298)) xor (layer0_outputs(3240)));
    outputs(5826) <= not((layer0_outputs(11307)) xor (layer0_outputs(6659)));
    outputs(5827) <= (layer0_outputs(11864)) xor (layer0_outputs(11243));
    outputs(5828) <= not(layer0_outputs(68));
    outputs(5829) <= layer0_outputs(63);
    outputs(5830) <= not(layer0_outputs(9443));
    outputs(5831) <= layer0_outputs(9725);
    outputs(5832) <= (layer0_outputs(6895)) and not (layer0_outputs(10539));
    outputs(5833) <= not(layer0_outputs(9783));
    outputs(5834) <= not(layer0_outputs(8662)) or (layer0_outputs(8319));
    outputs(5835) <= not(layer0_outputs(4119));
    outputs(5836) <= not(layer0_outputs(11875));
    outputs(5837) <= not(layer0_outputs(5262));
    outputs(5838) <= not(layer0_outputs(41));
    outputs(5839) <= (layer0_outputs(10582)) xor (layer0_outputs(2454));
    outputs(5840) <= layer0_outputs(11144);
    outputs(5841) <= (layer0_outputs(8819)) and (layer0_outputs(1341));
    outputs(5842) <= not(layer0_outputs(694));
    outputs(5843) <= (layer0_outputs(3008)) xor (layer0_outputs(8349));
    outputs(5844) <= not(layer0_outputs(2729)) or (layer0_outputs(4161));
    outputs(5845) <= layer0_outputs(9710);
    outputs(5846) <= not(layer0_outputs(11416));
    outputs(5847) <= not((layer0_outputs(774)) xor (layer0_outputs(863)));
    outputs(5848) <= not((layer0_outputs(4494)) xor (layer0_outputs(3936)));
    outputs(5849) <= (layer0_outputs(11871)) and (layer0_outputs(6506));
    outputs(5850) <= not(layer0_outputs(3630));
    outputs(5851) <= (layer0_outputs(6362)) xor (layer0_outputs(7360));
    outputs(5852) <= not(layer0_outputs(1663)) or (layer0_outputs(10858));
    outputs(5853) <= layer0_outputs(7262);
    outputs(5854) <= not(layer0_outputs(8078)) or (layer0_outputs(3455));
    outputs(5855) <= layer0_outputs(7989);
    outputs(5856) <= (layer0_outputs(8258)) and not (layer0_outputs(12319));
    outputs(5857) <= (layer0_outputs(4933)) and not (layer0_outputs(7026));
    outputs(5858) <= not((layer0_outputs(7522)) and (layer0_outputs(5097)));
    outputs(5859) <= layer0_outputs(8963);
    outputs(5860) <= (layer0_outputs(11213)) and not (layer0_outputs(12550));
    outputs(5861) <= not((layer0_outputs(12058)) or (layer0_outputs(6854)));
    outputs(5862) <= not((layer0_outputs(6388)) xor (layer0_outputs(8513)));
    outputs(5863) <= (layer0_outputs(12702)) xor (layer0_outputs(2816));
    outputs(5864) <= layer0_outputs(1913);
    outputs(5865) <= (layer0_outputs(5302)) xor (layer0_outputs(8612));
    outputs(5866) <= layer0_outputs(577);
    outputs(5867) <= layer0_outputs(348);
    outputs(5868) <= not(layer0_outputs(4578)) or (layer0_outputs(7505));
    outputs(5869) <= not(layer0_outputs(9861));
    outputs(5870) <= layer0_outputs(1899);
    outputs(5871) <= (layer0_outputs(8467)) and (layer0_outputs(10012));
    outputs(5872) <= not(layer0_outputs(2795));
    outputs(5873) <= layer0_outputs(12129);
    outputs(5874) <= (layer0_outputs(9196)) xor (layer0_outputs(11915));
    outputs(5875) <= not(layer0_outputs(12743)) or (layer0_outputs(357));
    outputs(5876) <= not((layer0_outputs(9273)) xor (layer0_outputs(2361)));
    outputs(5877) <= (layer0_outputs(4641)) xor (layer0_outputs(9907));
    outputs(5878) <= (layer0_outputs(956)) xor (layer0_outputs(215));
    outputs(5879) <= layer0_outputs(6522);
    outputs(5880) <= (layer0_outputs(7214)) xor (layer0_outputs(2077));
    outputs(5881) <= layer0_outputs(11825);
    outputs(5882) <= layer0_outputs(6375);
    outputs(5883) <= layer0_outputs(8674);
    outputs(5884) <= layer0_outputs(8969);
    outputs(5885) <= (layer0_outputs(6864)) or (layer0_outputs(1281));
    outputs(5886) <= not((layer0_outputs(6705)) xor (layer0_outputs(8590)));
    outputs(5887) <= not(layer0_outputs(12484)) or (layer0_outputs(11158));
    outputs(5888) <= not(layer0_outputs(6297));
    outputs(5889) <= (layer0_outputs(2432)) and not (layer0_outputs(8283));
    outputs(5890) <= (layer0_outputs(9916)) xor (layer0_outputs(4034));
    outputs(5891) <= layer0_outputs(12181);
    outputs(5892) <= not(layer0_outputs(3201));
    outputs(5893) <= layer0_outputs(5261);
    outputs(5894) <= not(layer0_outputs(12401)) or (layer0_outputs(8329));
    outputs(5895) <= not(layer0_outputs(5277)) or (layer0_outputs(3161));
    outputs(5896) <= layer0_outputs(4356);
    outputs(5897) <= not(layer0_outputs(1675)) or (layer0_outputs(9639));
    outputs(5898) <= layer0_outputs(929);
    outputs(5899) <= not((layer0_outputs(5802)) xor (layer0_outputs(3247)));
    outputs(5900) <= not((layer0_outputs(7990)) and (layer0_outputs(8323)));
    outputs(5901) <= (layer0_outputs(4612)) and not (layer0_outputs(1326));
    outputs(5902) <= not(layer0_outputs(8683));
    outputs(5903) <= layer0_outputs(9721);
    outputs(5904) <= layer0_outputs(4821);
    outputs(5905) <= not(layer0_outputs(11866)) or (layer0_outputs(5724));
    outputs(5906) <= layer0_outputs(5590);
    outputs(5907) <= not(layer0_outputs(6881));
    outputs(5908) <= (layer0_outputs(6899)) and not (layer0_outputs(2127));
    outputs(5909) <= not(layer0_outputs(3065));
    outputs(5910) <= not(layer0_outputs(9741));
    outputs(5911) <= not(layer0_outputs(8139));
    outputs(5912) <= layer0_outputs(474);
    outputs(5913) <= layer0_outputs(6391);
    outputs(5914) <= (layer0_outputs(12272)) and (layer0_outputs(3429));
    outputs(5915) <= layer0_outputs(953);
    outputs(5916) <= layer0_outputs(12765);
    outputs(5917) <= layer0_outputs(4666);
    outputs(5918) <= (layer0_outputs(7774)) and (layer0_outputs(12314));
    outputs(5919) <= layer0_outputs(12636);
    outputs(5920) <= layer0_outputs(5663);
    outputs(5921) <= not(layer0_outputs(7093)) or (layer0_outputs(1538));
    outputs(5922) <= not(layer0_outputs(11326));
    outputs(5923) <= (layer0_outputs(8004)) or (layer0_outputs(8501));
    outputs(5924) <= layer0_outputs(3828);
    outputs(5925) <= layer0_outputs(6229);
    outputs(5926) <= layer0_outputs(11896);
    outputs(5927) <= not(layer0_outputs(12215));
    outputs(5928) <= not(layer0_outputs(4924));
    outputs(5929) <= not(layer0_outputs(2868));
    outputs(5930) <= layer0_outputs(12474);
    outputs(5931) <= (layer0_outputs(7708)) or (layer0_outputs(10776));
    outputs(5932) <= not(layer0_outputs(7458));
    outputs(5933) <= layer0_outputs(3597);
    outputs(5934) <= (layer0_outputs(8791)) and (layer0_outputs(3533));
    outputs(5935) <= not((layer0_outputs(2926)) xor (layer0_outputs(6034)));
    outputs(5936) <= not(layer0_outputs(1079));
    outputs(5937) <= layer0_outputs(7097);
    outputs(5938) <= not(layer0_outputs(3524)) or (layer0_outputs(6673));
    outputs(5939) <= not((layer0_outputs(12202)) or (layer0_outputs(11635)));
    outputs(5940) <= layer0_outputs(6475);
    outputs(5941) <= not((layer0_outputs(205)) xor (layer0_outputs(9430)));
    outputs(5942) <= not((layer0_outputs(10077)) xor (layer0_outputs(8380)));
    outputs(5943) <= (layer0_outputs(7351)) and not (layer0_outputs(10079));
    outputs(5944) <= layer0_outputs(8459);
    outputs(5945) <= (layer0_outputs(4367)) xor (layer0_outputs(9203));
    outputs(5946) <= layer0_outputs(5017);
    outputs(5947) <= not((layer0_outputs(1000)) xor (layer0_outputs(11049)));
    outputs(5948) <= (layer0_outputs(619)) and not (layer0_outputs(2191));
    outputs(5949) <= not(layer0_outputs(695));
    outputs(5950) <= not(layer0_outputs(2750)) or (layer0_outputs(6739));
    outputs(5951) <= not(layer0_outputs(9256));
    outputs(5952) <= layer0_outputs(10605);
    outputs(5953) <= not((layer0_outputs(983)) or (layer0_outputs(4101)));
    outputs(5954) <= not(layer0_outputs(6114)) or (layer0_outputs(8310));
    outputs(5955) <= (layer0_outputs(8146)) and not (layer0_outputs(11597));
    outputs(5956) <= (layer0_outputs(7540)) xor (layer0_outputs(8339));
    outputs(5957) <= not(layer0_outputs(5845)) or (layer0_outputs(322));
    outputs(5958) <= not(layer0_outputs(5995));
    outputs(5959) <= layer0_outputs(10085);
    outputs(5960) <= (layer0_outputs(6335)) and not (layer0_outputs(4728));
    outputs(5961) <= not(layer0_outputs(10853)) or (layer0_outputs(6001));
    outputs(5962) <= layer0_outputs(3112);
    outputs(5963) <= not(layer0_outputs(8606));
    outputs(5964) <= not((layer0_outputs(4391)) or (layer0_outputs(9981)));
    outputs(5965) <= not((layer0_outputs(8088)) xor (layer0_outputs(293)));
    outputs(5966) <= not((layer0_outputs(5756)) xor (layer0_outputs(7545)));
    outputs(5967) <= not(layer0_outputs(10001));
    outputs(5968) <= not(layer0_outputs(1631)) or (layer0_outputs(5049));
    outputs(5969) <= not((layer0_outputs(1977)) xor (layer0_outputs(1234)));
    outputs(5970) <= (layer0_outputs(590)) and not (layer0_outputs(11040));
    outputs(5971) <= layer0_outputs(4753);
    outputs(5972) <= not(layer0_outputs(7442));
    outputs(5973) <= not(layer0_outputs(7484));
    outputs(5974) <= (layer0_outputs(11736)) xor (layer0_outputs(2285));
    outputs(5975) <= not(layer0_outputs(771));
    outputs(5976) <= layer0_outputs(11524);
    outputs(5977) <= (layer0_outputs(3377)) or (layer0_outputs(8605));
    outputs(5978) <= not(layer0_outputs(803));
    outputs(5979) <= not((layer0_outputs(1611)) xor (layer0_outputs(3930)));
    outputs(5980) <= layer0_outputs(962);
    outputs(5981) <= not(layer0_outputs(10274));
    outputs(5982) <= not(layer0_outputs(2536));
    outputs(5983) <= (layer0_outputs(625)) and (layer0_outputs(9637));
    outputs(5984) <= not((layer0_outputs(7962)) or (layer0_outputs(3036)));
    outputs(5985) <= (layer0_outputs(4209)) and not (layer0_outputs(7965));
    outputs(5986) <= not(layer0_outputs(9788));
    outputs(5987) <= not((layer0_outputs(12768)) or (layer0_outputs(2810)));
    outputs(5988) <= not(layer0_outputs(4647)) or (layer0_outputs(2827));
    outputs(5989) <= not(layer0_outputs(4795)) or (layer0_outputs(572));
    outputs(5990) <= not(layer0_outputs(960)) or (layer0_outputs(10703));
    outputs(5991) <= not((layer0_outputs(12709)) or (layer0_outputs(7837)));
    outputs(5992) <= layer0_outputs(8392);
    outputs(5993) <= not(layer0_outputs(841));
    outputs(5994) <= (layer0_outputs(10905)) and not (layer0_outputs(1903));
    outputs(5995) <= not((layer0_outputs(4841)) or (layer0_outputs(4549)));
    outputs(5996) <= (layer0_outputs(5184)) xor (layer0_outputs(5284));
    outputs(5997) <= (layer0_outputs(5320)) or (layer0_outputs(5924));
    outputs(5998) <= not(layer0_outputs(3852));
    outputs(5999) <= layer0_outputs(11298);
    outputs(6000) <= not((layer0_outputs(138)) or (layer0_outputs(7706)));
    outputs(6001) <= layer0_outputs(7767);
    outputs(6002) <= layer0_outputs(5661);
    outputs(6003) <= not((layer0_outputs(1238)) or (layer0_outputs(9558)));
    outputs(6004) <= layer0_outputs(2962);
    outputs(6005) <= layer0_outputs(2652);
    outputs(6006) <= layer0_outputs(663);
    outputs(6007) <= (layer0_outputs(587)) xor (layer0_outputs(10330));
    outputs(6008) <= (layer0_outputs(12414)) or (layer0_outputs(11057));
    outputs(6009) <= not((layer0_outputs(4613)) or (layer0_outputs(7874)));
    outputs(6010) <= not((layer0_outputs(9013)) or (layer0_outputs(11378)));
    outputs(6011) <= (layer0_outputs(5309)) and not (layer0_outputs(12044));
    outputs(6012) <= (layer0_outputs(5185)) and not (layer0_outputs(7006));
    outputs(6013) <= (layer0_outputs(8801)) xor (layer0_outputs(7932));
    outputs(6014) <= not(layer0_outputs(3208));
    outputs(6015) <= not(layer0_outputs(951)) or (layer0_outputs(1768));
    outputs(6016) <= not(layer0_outputs(1507)) or (layer0_outputs(1471));
    outputs(6017) <= not((layer0_outputs(2997)) xor (layer0_outputs(2763)));
    outputs(6018) <= layer0_outputs(10043);
    outputs(6019) <= (layer0_outputs(5840)) and not (layer0_outputs(977));
    outputs(6020) <= layer0_outputs(6272);
    outputs(6021) <= not((layer0_outputs(9270)) or (layer0_outputs(6438)));
    outputs(6022) <= (layer0_outputs(7275)) xor (layer0_outputs(2368));
    outputs(6023) <= not(layer0_outputs(6945));
    outputs(6024) <= layer0_outputs(11977);
    outputs(6025) <= (layer0_outputs(533)) and not (layer0_outputs(3125));
    outputs(6026) <= not(layer0_outputs(10140));
    outputs(6027) <= (layer0_outputs(6816)) xor (layer0_outputs(7722));
    outputs(6028) <= not((layer0_outputs(299)) xor (layer0_outputs(134)));
    outputs(6029) <= not(layer0_outputs(8301));
    outputs(6030) <= not(layer0_outputs(4142));
    outputs(6031) <= (layer0_outputs(10548)) xor (layer0_outputs(9800));
    outputs(6032) <= (layer0_outputs(4412)) xor (layer0_outputs(6821));
    outputs(6033) <= not((layer0_outputs(7207)) or (layer0_outputs(5048)));
    outputs(6034) <= not((layer0_outputs(2056)) xor (layer0_outputs(1261)));
    outputs(6035) <= (layer0_outputs(6032)) or (layer0_outputs(7174));
    outputs(6036) <= layer0_outputs(2486);
    outputs(6037) <= not(layer0_outputs(11992));
    outputs(6038) <= layer0_outputs(11123);
    outputs(6039) <= (layer0_outputs(859)) and not (layer0_outputs(5527));
    outputs(6040) <= (layer0_outputs(7785)) and (layer0_outputs(5653));
    outputs(6041) <= not(layer0_outputs(1605)) or (layer0_outputs(10711));
    outputs(6042) <= not((layer0_outputs(6683)) xor (layer0_outputs(11302)));
    outputs(6043) <= (layer0_outputs(3147)) or (layer0_outputs(4349));
    outputs(6044) <= layer0_outputs(3329);
    outputs(6045) <= not(layer0_outputs(3966));
    outputs(6046) <= (layer0_outputs(9711)) or (layer0_outputs(4135));
    outputs(6047) <= (layer0_outputs(3349)) and not (layer0_outputs(8777));
    outputs(6048) <= layer0_outputs(4389);
    outputs(6049) <= not(layer0_outputs(9320));
    outputs(6050) <= layer0_outputs(560);
    outputs(6051) <= (layer0_outputs(12146)) xor (layer0_outputs(7263));
    outputs(6052) <= (layer0_outputs(1425)) and not (layer0_outputs(10635));
    outputs(6053) <= not(layer0_outputs(4303));
    outputs(6054) <= (layer0_outputs(10014)) xor (layer0_outputs(7780));
    outputs(6055) <= not(layer0_outputs(157));
    outputs(6056) <= not(layer0_outputs(7032));
    outputs(6057) <= (layer0_outputs(3002)) and (layer0_outputs(11617));
    outputs(6058) <= not((layer0_outputs(3836)) xor (layer0_outputs(6402)));
    outputs(6059) <= (layer0_outputs(11408)) and (layer0_outputs(8393));
    outputs(6060) <= layer0_outputs(9751);
    outputs(6061) <= (layer0_outputs(112)) xor (layer0_outputs(5283));
    outputs(6062) <= (layer0_outputs(3988)) xor (layer0_outputs(5956));
    outputs(6063) <= (layer0_outputs(5695)) and not (layer0_outputs(2557));
    outputs(6064) <= not((layer0_outputs(12548)) xor (layer0_outputs(5018)));
    outputs(6065) <= layer0_outputs(7681);
    outputs(6066) <= not(layer0_outputs(6027)) or (layer0_outputs(9670));
    outputs(6067) <= not(layer0_outputs(7890));
    outputs(6068) <= not(layer0_outputs(12775)) or (layer0_outputs(3554));
    outputs(6069) <= (layer0_outputs(10811)) xor (layer0_outputs(6744));
    outputs(6070) <= layer0_outputs(3264);
    outputs(6071) <= (layer0_outputs(10321)) xor (layer0_outputs(9223));
    outputs(6072) <= (layer0_outputs(9664)) or (layer0_outputs(3902));
    outputs(6073) <= not(layer0_outputs(8562));
    outputs(6074) <= layer0_outputs(5234);
    outputs(6075) <= not(layer0_outputs(4776)) or (layer0_outputs(10971));
    outputs(6076) <= layer0_outputs(4310);
    outputs(6077) <= not(layer0_outputs(10719));
    outputs(6078) <= not(layer0_outputs(11365));
    outputs(6079) <= not(layer0_outputs(9225));
    outputs(6080) <= (layer0_outputs(343)) and (layer0_outputs(1931));
    outputs(6081) <= not((layer0_outputs(5488)) or (layer0_outputs(5884)));
    outputs(6082) <= layer0_outputs(5209);
    outputs(6083) <= layer0_outputs(9156);
    outputs(6084) <= not(layer0_outputs(7235));
    outputs(6085) <= not(layer0_outputs(951));
    outputs(6086) <= not(layer0_outputs(413));
    outputs(6087) <= (layer0_outputs(889)) or (layer0_outputs(10982));
    outputs(6088) <= not((layer0_outputs(6482)) xor (layer0_outputs(3111)));
    outputs(6089) <= (layer0_outputs(11551)) and not (layer0_outputs(4633));
    outputs(6090) <= (layer0_outputs(10128)) and (layer0_outputs(8312));
    outputs(6091) <= not((layer0_outputs(1660)) xor (layer0_outputs(10685)));
    outputs(6092) <= layer0_outputs(5900);
    outputs(6093) <= (layer0_outputs(3960)) and not (layer0_outputs(1600));
    outputs(6094) <= not(layer0_outputs(7540));
    outputs(6095) <= (layer0_outputs(6369)) xor (layer0_outputs(4288));
    outputs(6096) <= not((layer0_outputs(4085)) xor (layer0_outputs(9507)));
    outputs(6097) <= not((layer0_outputs(5194)) or (layer0_outputs(5961)));
    outputs(6098) <= (layer0_outputs(5258)) and not (layer0_outputs(10296));
    outputs(6099) <= not(layer0_outputs(7475));
    outputs(6100) <= layer0_outputs(2757);
    outputs(6101) <= layer0_outputs(6162);
    outputs(6102) <= (layer0_outputs(3677)) xor (layer0_outputs(12799));
    outputs(6103) <= not(layer0_outputs(6093));
    outputs(6104) <= not(layer0_outputs(11293));
    outputs(6105) <= not(layer0_outputs(11233));
    outputs(6106) <= not(layer0_outputs(6865));
    outputs(6107) <= not((layer0_outputs(8607)) xor (layer0_outputs(1388)));
    outputs(6108) <= not((layer0_outputs(4950)) xor (layer0_outputs(1108)));
    outputs(6109) <= not((layer0_outputs(11662)) or (layer0_outputs(356)));
    outputs(6110) <= layer0_outputs(8256);
    outputs(6111) <= not((layer0_outputs(4619)) and (layer0_outputs(6152)));
    outputs(6112) <= not((layer0_outputs(7252)) and (layer0_outputs(10682)));
    outputs(6113) <= not(layer0_outputs(7866));
    outputs(6114) <= not(layer0_outputs(10744)) or (layer0_outputs(7861));
    outputs(6115) <= not(layer0_outputs(3104));
    outputs(6116) <= not((layer0_outputs(10981)) xor (layer0_outputs(3521)));
    outputs(6117) <= not((layer0_outputs(9293)) xor (layer0_outputs(2730)));
    outputs(6118) <= not(layer0_outputs(170)) or (layer0_outputs(4998));
    outputs(6119) <= layer0_outputs(5782);
    outputs(6120) <= layer0_outputs(3634);
    outputs(6121) <= not((layer0_outputs(1594)) xor (layer0_outputs(8479)));
    outputs(6122) <= (layer0_outputs(823)) xor (layer0_outputs(8212));
    outputs(6123) <= not((layer0_outputs(8362)) xor (layer0_outputs(2474)));
    outputs(6124) <= not(layer0_outputs(7558));
    outputs(6125) <= layer0_outputs(3493);
    outputs(6126) <= not(layer0_outputs(8204)) or (layer0_outputs(3827));
    outputs(6127) <= not(layer0_outputs(4898));
    outputs(6128) <= layer0_outputs(3671);
    outputs(6129) <= (layer0_outputs(6466)) and (layer0_outputs(1098));
    outputs(6130) <= not(layer0_outputs(6804));
    outputs(6131) <= not(layer0_outputs(12080));
    outputs(6132) <= (layer0_outputs(9061)) xor (layer0_outputs(4354));
    outputs(6133) <= (layer0_outputs(1357)) and not (layer0_outputs(1935));
    outputs(6134) <= not((layer0_outputs(6137)) xor (layer0_outputs(5552)));
    outputs(6135) <= (layer0_outputs(7380)) xor (layer0_outputs(1096));
    outputs(6136) <= not((layer0_outputs(9204)) and (layer0_outputs(8167)));
    outputs(6137) <= (layer0_outputs(9439)) xor (layer0_outputs(10279));
    outputs(6138) <= layer0_outputs(12512);
    outputs(6139) <= not(layer0_outputs(5949));
    outputs(6140) <= layer0_outputs(12238);
    outputs(6141) <= (layer0_outputs(3585)) and (layer0_outputs(12468));
    outputs(6142) <= layer0_outputs(3799);
    outputs(6143) <= layer0_outputs(588);
    outputs(6144) <= (layer0_outputs(8045)) xor (layer0_outputs(11186));
    outputs(6145) <= layer0_outputs(919);
    outputs(6146) <= (layer0_outputs(7071)) xor (layer0_outputs(7647));
    outputs(6147) <= not(layer0_outputs(1724));
    outputs(6148) <= not(layer0_outputs(5829)) or (layer0_outputs(10748));
    outputs(6149) <= layer0_outputs(2647);
    outputs(6150) <= layer0_outputs(12322);
    outputs(6151) <= (layer0_outputs(682)) and not (layer0_outputs(8356));
    outputs(6152) <= (layer0_outputs(5129)) and not (layer0_outputs(9206));
    outputs(6153) <= not(layer0_outputs(1790));
    outputs(6154) <= not((layer0_outputs(7556)) or (layer0_outputs(6037)));
    outputs(6155) <= not(layer0_outputs(3646));
    outputs(6156) <= not(layer0_outputs(2221));
    outputs(6157) <= layer0_outputs(7385);
    outputs(6158) <= not((layer0_outputs(10579)) or (layer0_outputs(3221)));
    outputs(6159) <= not((layer0_outputs(4042)) or (layer0_outputs(1420)));
    outputs(6160) <= not(layer0_outputs(1364));
    outputs(6161) <= not(layer0_outputs(4358));
    outputs(6162) <= not(layer0_outputs(260));
    outputs(6163) <= not(layer0_outputs(9487));
    outputs(6164) <= not((layer0_outputs(7616)) xor (layer0_outputs(4345)));
    outputs(6165) <= not(layer0_outputs(11002));
    outputs(6166) <= not(layer0_outputs(8412));
    outputs(6167) <= layer0_outputs(1840);
    outputs(6168) <= layer0_outputs(5483);
    outputs(6169) <= not(layer0_outputs(10563));
    outputs(6170) <= layer0_outputs(1584);
    outputs(6171) <= layer0_outputs(1471);
    outputs(6172) <= not(layer0_outputs(9124));
    outputs(6173) <= not(layer0_outputs(11749)) or (layer0_outputs(5344));
    outputs(6174) <= (layer0_outputs(6491)) xor (layer0_outputs(11978));
    outputs(6175) <= not(layer0_outputs(1451));
    outputs(6176) <= not(layer0_outputs(10685));
    outputs(6177) <= not(layer0_outputs(2425)) or (layer0_outputs(11563));
    outputs(6178) <= not(layer0_outputs(7055)) or (layer0_outputs(11800));
    outputs(6179) <= not(layer0_outputs(2005));
    outputs(6180) <= layer0_outputs(8484);
    outputs(6181) <= (layer0_outputs(11767)) xor (layer0_outputs(2075));
    outputs(6182) <= not((layer0_outputs(2076)) and (layer0_outputs(9060)));
    outputs(6183) <= not(layer0_outputs(7535)) or (layer0_outputs(3457));
    outputs(6184) <= not(layer0_outputs(3711));
    outputs(6185) <= layer0_outputs(6927);
    outputs(6186) <= layer0_outputs(9893);
    outputs(6187) <= not(layer0_outputs(2857));
    outputs(6188) <= (layer0_outputs(11117)) and (layer0_outputs(5754));
    outputs(6189) <= not(layer0_outputs(2207));
    outputs(6190) <= (layer0_outputs(11425)) xor (layer0_outputs(3123));
    outputs(6191) <= (layer0_outputs(10133)) xor (layer0_outputs(8941));
    outputs(6192) <= not((layer0_outputs(1412)) xor (layer0_outputs(4200)));
    outputs(6193) <= (layer0_outputs(2130)) or (layer0_outputs(9369));
    outputs(6194) <= not(layer0_outputs(8622));
    outputs(6195) <= not(layer0_outputs(8151));
    outputs(6196) <= (layer0_outputs(59)) xor (layer0_outputs(7748));
    outputs(6197) <= (layer0_outputs(9527)) and not (layer0_outputs(8233));
    outputs(6198) <= (layer0_outputs(2173)) xor (layer0_outputs(6476));
    outputs(6199) <= not(layer0_outputs(6400));
    outputs(6200) <= not((layer0_outputs(3584)) and (layer0_outputs(7791)));
    outputs(6201) <= not(layer0_outputs(12408)) or (layer0_outputs(12529));
    outputs(6202) <= not(layer0_outputs(11163));
    outputs(6203) <= not(layer0_outputs(8370));
    outputs(6204) <= not((layer0_outputs(9931)) and (layer0_outputs(8805)));
    outputs(6205) <= not(layer0_outputs(7577));
    outputs(6206) <= layer0_outputs(7489);
    outputs(6207) <= layer0_outputs(6814);
    outputs(6208) <= (layer0_outputs(506)) and (layer0_outputs(12385));
    outputs(6209) <= layer0_outputs(3889);
    outputs(6210) <= (layer0_outputs(8232)) and not (layer0_outputs(7057));
    outputs(6211) <= layer0_outputs(10179);
    outputs(6212) <= (layer0_outputs(3376)) and not (layer0_outputs(892));
    outputs(6213) <= layer0_outputs(10310);
    outputs(6214) <= not(layer0_outputs(8152));
    outputs(6215) <= not(layer0_outputs(12622));
    outputs(6216) <= (layer0_outputs(7925)) and not (layer0_outputs(9548));
    outputs(6217) <= (layer0_outputs(241)) xor (layer0_outputs(414));
    outputs(6218) <= not(layer0_outputs(4710));
    outputs(6219) <= (layer0_outputs(5196)) xor (layer0_outputs(3068));
    outputs(6220) <= layer0_outputs(10591);
    outputs(6221) <= not((layer0_outputs(16)) xor (layer0_outputs(493)));
    outputs(6222) <= layer0_outputs(993);
    outputs(6223) <= not((layer0_outputs(5263)) xor (layer0_outputs(9555)));
    outputs(6224) <= (layer0_outputs(10145)) and not (layer0_outputs(12305));
    outputs(6225) <= not(layer0_outputs(5570));
    outputs(6226) <= (layer0_outputs(1452)) and (layer0_outputs(3688));
    outputs(6227) <= not(layer0_outputs(6801));
    outputs(6228) <= (layer0_outputs(3053)) and not (layer0_outputs(8442));
    outputs(6229) <= layer0_outputs(10689);
    outputs(6230) <= not((layer0_outputs(9787)) xor (layer0_outputs(10256)));
    outputs(6231) <= (layer0_outputs(10961)) xor (layer0_outputs(6520));
    outputs(6232) <= layer0_outputs(3765);
    outputs(6233) <= (layer0_outputs(1820)) and (layer0_outputs(12119));
    outputs(6234) <= (layer0_outputs(3137)) xor (layer0_outputs(5391));
    outputs(6235) <= not(layer0_outputs(10428));
    outputs(6236) <= layer0_outputs(10859);
    outputs(6237) <= layer0_outputs(5436);
    outputs(6238) <= layer0_outputs(5776);
    outputs(6239) <= layer0_outputs(3419);
    outputs(6240) <= not((layer0_outputs(7597)) and (layer0_outputs(8727)));
    outputs(6241) <= layer0_outputs(9927);
    outputs(6242) <= not(layer0_outputs(7156));
    outputs(6243) <= (layer0_outputs(4751)) xor (layer0_outputs(8880));
    outputs(6244) <= not(layer0_outputs(1321)) or (layer0_outputs(5809));
    outputs(6245) <= (layer0_outputs(5929)) and not (layer0_outputs(6939));
    outputs(6246) <= not((layer0_outputs(9465)) xor (layer0_outputs(370)));
    outputs(6247) <= (layer0_outputs(11026)) xor (layer0_outputs(8343));
    outputs(6248) <= not(layer0_outputs(8727));
    outputs(6249) <= not((layer0_outputs(8160)) xor (layer0_outputs(1612)));
    outputs(6250) <= not((layer0_outputs(6138)) and (layer0_outputs(2941)));
    outputs(6251) <= layer0_outputs(8631);
    outputs(6252) <= layer0_outputs(10852);
    outputs(6253) <= (layer0_outputs(8179)) xor (layer0_outputs(4971));
    outputs(6254) <= not(layer0_outputs(9479)) or (layer0_outputs(4936));
    outputs(6255) <= layer0_outputs(8382);
    outputs(6256) <= not(layer0_outputs(5475));
    outputs(6257) <= not(layer0_outputs(3230));
    outputs(6258) <= not(layer0_outputs(5354)) or (layer0_outputs(9237));
    outputs(6259) <= layer0_outputs(3328);
    outputs(6260) <= (layer0_outputs(12188)) and (layer0_outputs(12782));
    outputs(6261) <= (layer0_outputs(832)) xor (layer0_outputs(5219));
    outputs(6262) <= layer0_outputs(4804);
    outputs(6263) <= layer0_outputs(1157);
    outputs(6264) <= (layer0_outputs(11738)) xor (layer0_outputs(850));
    outputs(6265) <= not(layer0_outputs(4751));
    outputs(6266) <= (layer0_outputs(10753)) and (layer0_outputs(8807));
    outputs(6267) <= not((layer0_outputs(5522)) and (layer0_outputs(5382)));
    outputs(6268) <= not(layer0_outputs(9686));
    outputs(6269) <= (layer0_outputs(12637)) xor (layer0_outputs(7126));
    outputs(6270) <= layer0_outputs(4772);
    outputs(6271) <= (layer0_outputs(2118)) and not (layer0_outputs(6465));
    outputs(6272) <= (layer0_outputs(6568)) and not (layer0_outputs(3471));
    outputs(6273) <= (layer0_outputs(9369)) and not (layer0_outputs(2192));
    outputs(6274) <= not(layer0_outputs(1444));
    outputs(6275) <= not(layer0_outputs(8321)) or (layer0_outputs(9995));
    outputs(6276) <= not((layer0_outputs(3564)) xor (layer0_outputs(3638)));
    outputs(6277) <= not((layer0_outputs(7657)) xor (layer0_outputs(627)));
    outputs(6278) <= (layer0_outputs(10849)) and (layer0_outputs(5767));
    outputs(6279) <= not(layer0_outputs(1032)) or (layer0_outputs(10657));
    outputs(6280) <= (layer0_outputs(12112)) and (layer0_outputs(2896));
    outputs(6281) <= not((layer0_outputs(11076)) and (layer0_outputs(11439)));
    outputs(6282) <= (layer0_outputs(2659)) and (layer0_outputs(12711));
    outputs(6283) <= not(layer0_outputs(1759));
    outputs(6284) <= (layer0_outputs(4450)) xor (layer0_outputs(255));
    outputs(6285) <= not(layer0_outputs(11673));
    outputs(6286) <= (layer0_outputs(5600)) xor (layer0_outputs(2884));
    outputs(6287) <= not(layer0_outputs(8514)) or (layer0_outputs(1467));
    outputs(6288) <= (layer0_outputs(10119)) and (layer0_outputs(9134));
    outputs(6289) <= not((layer0_outputs(12148)) xor (layer0_outputs(6994)));
    outputs(6290) <= layer0_outputs(4397);
    outputs(6291) <= '1';
    outputs(6292) <= not(layer0_outputs(2467));
    outputs(6293) <= not(layer0_outputs(9049));
    outputs(6294) <= (layer0_outputs(9405)) and (layer0_outputs(11198));
    outputs(6295) <= (layer0_outputs(2094)) xor (layer0_outputs(7111));
    outputs(6296) <= not((layer0_outputs(7095)) or (layer0_outputs(4016)));
    outputs(6297) <= (layer0_outputs(7165)) and not (layer0_outputs(9366));
    outputs(6298) <= layer0_outputs(12040);
    outputs(6299) <= (layer0_outputs(12442)) xor (layer0_outputs(6762));
    outputs(6300) <= layer0_outputs(2607);
    outputs(6301) <= not((layer0_outputs(79)) xor (layer0_outputs(4558)));
    outputs(6302) <= (layer0_outputs(1074)) and not (layer0_outputs(1373));
    outputs(6303) <= not(layer0_outputs(7249)) or (layer0_outputs(2101));
    outputs(6304) <= layer0_outputs(2150);
    outputs(6305) <= not(layer0_outputs(1790));
    outputs(6306) <= not(layer0_outputs(10507));
    outputs(6307) <= not(layer0_outputs(4904));
    outputs(6308) <= layer0_outputs(7653);
    outputs(6309) <= (layer0_outputs(1055)) or (layer0_outputs(7801));
    outputs(6310) <= not(layer0_outputs(2018)) or (layer0_outputs(6153));
    outputs(6311) <= not(layer0_outputs(6353)) or (layer0_outputs(4436));
    outputs(6312) <= not(layer0_outputs(2492));
    outputs(6313) <= not((layer0_outputs(11467)) xor (layer0_outputs(7153)));
    outputs(6314) <= layer0_outputs(11959);
    outputs(6315) <= (layer0_outputs(11701)) xor (layer0_outputs(7074));
    outputs(6316) <= layer0_outputs(11194);
    outputs(6317) <= not(layer0_outputs(10527));
    outputs(6318) <= (layer0_outputs(4614)) xor (layer0_outputs(10376));
    outputs(6319) <= layer0_outputs(6349);
    outputs(6320) <= layer0_outputs(10502);
    outputs(6321) <= layer0_outputs(10172);
    outputs(6322) <= (layer0_outputs(1916)) xor (layer0_outputs(7921));
    outputs(6323) <= layer0_outputs(8100);
    outputs(6324) <= not(layer0_outputs(6423)) or (layer0_outputs(9265));
    outputs(6325) <= not((layer0_outputs(11899)) xor (layer0_outputs(2453)));
    outputs(6326) <= not((layer0_outputs(8797)) xor (layer0_outputs(10597)));
    outputs(6327) <= (layer0_outputs(8875)) xor (layer0_outputs(2072));
    outputs(6328) <= (layer0_outputs(4923)) xor (layer0_outputs(11587));
    outputs(6329) <= not(layer0_outputs(692));
    outputs(6330) <= (layer0_outputs(11032)) xor (layer0_outputs(9628));
    outputs(6331) <= (layer0_outputs(3558)) xor (layer0_outputs(10032));
    outputs(6332) <= (layer0_outputs(10693)) and not (layer0_outputs(1362));
    outputs(6333) <= layer0_outputs(4188);
    outputs(6334) <= layer0_outputs(8072);
    outputs(6335) <= not((layer0_outputs(6790)) xor (layer0_outputs(6454)));
    outputs(6336) <= layer0_outputs(11358);
    outputs(6337) <= not((layer0_outputs(10770)) xor (layer0_outputs(2882)));
    outputs(6338) <= (layer0_outputs(6589)) and not (layer0_outputs(11512));
    outputs(6339) <= (layer0_outputs(9374)) and (layer0_outputs(8458));
    outputs(6340) <= layer0_outputs(3153);
    outputs(6341) <= (layer0_outputs(10763)) xor (layer0_outputs(3339));
    outputs(6342) <= not(layer0_outputs(2548));
    outputs(6343) <= not(layer0_outputs(2289));
    outputs(6344) <= not(layer0_outputs(10188));
    outputs(6345) <= not(layer0_outputs(3345));
    outputs(6346) <= not((layer0_outputs(2695)) xor (layer0_outputs(11876)));
    outputs(6347) <= layer0_outputs(395);
    outputs(6348) <= layer0_outputs(9585);
    outputs(6349) <= not(layer0_outputs(2792));
    outputs(6350) <= not((layer0_outputs(12115)) xor (layer0_outputs(2086)));
    outputs(6351) <= (layer0_outputs(726)) and not (layer0_outputs(1937));
    outputs(6352) <= layer0_outputs(1486);
    outputs(6353) <= (layer0_outputs(2790)) xor (layer0_outputs(4063));
    outputs(6354) <= (layer0_outputs(9877)) xor (layer0_outputs(2812));
    outputs(6355) <= not((layer0_outputs(3021)) xor (layer0_outputs(1949)));
    outputs(6356) <= layer0_outputs(9922);
    outputs(6357) <= (layer0_outputs(10979)) and not (layer0_outputs(2216));
    outputs(6358) <= layer0_outputs(4655);
    outputs(6359) <= not(layer0_outputs(1383)) or (layer0_outputs(9447));
    outputs(6360) <= (layer0_outputs(5807)) and (layer0_outputs(10328));
    outputs(6361) <= (layer0_outputs(4097)) and (layer0_outputs(365));
    outputs(6362) <= (layer0_outputs(12039)) or (layer0_outputs(7951));
    outputs(6363) <= layer0_outputs(9318);
    outputs(6364) <= not(layer0_outputs(4157));
    outputs(6365) <= layer0_outputs(4111);
    outputs(6366) <= not((layer0_outputs(3300)) xor (layer0_outputs(9063)));
    outputs(6367) <= not(layer0_outputs(74));
    outputs(6368) <= not((layer0_outputs(2966)) and (layer0_outputs(7372)));
    outputs(6369) <= layer0_outputs(2539);
    outputs(6370) <= not(layer0_outputs(6675));
    outputs(6371) <= (layer0_outputs(9894)) and (layer0_outputs(1906));
    outputs(6372) <= layer0_outputs(1376);
    outputs(6373) <= not((layer0_outputs(6496)) or (layer0_outputs(8049)));
    outputs(6374) <= layer0_outputs(8884);
    outputs(6375) <= (layer0_outputs(10253)) xor (layer0_outputs(4899));
    outputs(6376) <= (layer0_outputs(5533)) and not (layer0_outputs(9999));
    outputs(6377) <= (layer0_outputs(11071)) or (layer0_outputs(4818));
    outputs(6378) <= layer0_outputs(8760);
    outputs(6379) <= (layer0_outputs(8532)) and not (layer0_outputs(708));
    outputs(6380) <= not(layer0_outputs(10486));
    outputs(6381) <= not(layer0_outputs(6037));
    outputs(6382) <= not(layer0_outputs(496));
    outputs(6383) <= not(layer0_outputs(8430));
    outputs(6384) <= not(layer0_outputs(12654));
    outputs(6385) <= not(layer0_outputs(3777));
    outputs(6386) <= layer0_outputs(11009);
    outputs(6387) <= (layer0_outputs(11444)) and not (layer0_outputs(3854));
    outputs(6388) <= not(layer0_outputs(655)) or (layer0_outputs(12351));
    outputs(6389) <= layer0_outputs(7262);
    outputs(6390) <= layer0_outputs(10181);
    outputs(6391) <= layer0_outputs(6806);
    outputs(6392) <= not(layer0_outputs(6878));
    outputs(6393) <= (layer0_outputs(9466)) xor (layer0_outputs(6034));
    outputs(6394) <= (layer0_outputs(12596)) xor (layer0_outputs(8563));
    outputs(6395) <= (layer0_outputs(8247)) and (layer0_outputs(1518));
    outputs(6396) <= not(layer0_outputs(10917));
    outputs(6397) <= (layer0_outputs(659)) and (layer0_outputs(8154));
    outputs(6398) <= (layer0_outputs(11737)) xor (layer0_outputs(11453));
    outputs(6399) <= layer0_outputs(9088);
    outputs(6400) <= not(layer0_outputs(3110));
    outputs(6401) <= not(layer0_outputs(12771));
    outputs(6402) <= not(layer0_outputs(5448));
    outputs(6403) <= layer0_outputs(289);
    outputs(6404) <= not(layer0_outputs(3778));
    outputs(6405) <= not(layer0_outputs(10345));
    outputs(6406) <= layer0_outputs(12542);
    outputs(6407) <= not(layer0_outputs(3674)) or (layer0_outputs(3696));
    outputs(6408) <= not(layer0_outputs(9381));
    outputs(6409) <= not((layer0_outputs(824)) and (layer0_outputs(6526)));
    outputs(6410) <= not(layer0_outputs(11013));
    outputs(6411) <= not((layer0_outputs(10104)) xor (layer0_outputs(10746)));
    outputs(6412) <= layer0_outputs(6822);
    outputs(6413) <= (layer0_outputs(7836)) xor (layer0_outputs(3741));
    outputs(6414) <= layer0_outputs(8067);
    outputs(6415) <= not(layer0_outputs(1478)) or (layer0_outputs(7532));
    outputs(6416) <= not((layer0_outputs(392)) xor (layer0_outputs(11992)));
    outputs(6417) <= not((layer0_outputs(7637)) and (layer0_outputs(3532)));
    outputs(6418) <= not(layer0_outputs(1589)) or (layer0_outputs(7615));
    outputs(6419) <= layer0_outputs(3246);
    outputs(6420) <= (layer0_outputs(7939)) xor (layer0_outputs(1236));
    outputs(6421) <= not(layer0_outputs(4116));
    outputs(6422) <= (layer0_outputs(11281)) xor (layer0_outputs(5577));
    outputs(6423) <= not((layer0_outputs(10660)) or (layer0_outputs(5362)));
    outputs(6424) <= not(layer0_outputs(464));
    outputs(6425) <= (layer0_outputs(10349)) and not (layer0_outputs(10697));
    outputs(6426) <= layer0_outputs(10940);
    outputs(6427) <= (layer0_outputs(12551)) xor (layer0_outputs(7246));
    outputs(6428) <= (layer0_outputs(5175)) xor (layer0_outputs(5605));
    outputs(6429) <= layer0_outputs(10805);
    outputs(6430) <= not(layer0_outputs(4027));
    outputs(6431) <= layer0_outputs(10337);
    outputs(6432) <= (layer0_outputs(563)) xor (layer0_outputs(756));
    outputs(6433) <= layer0_outputs(12641);
    outputs(6434) <= not(layer0_outputs(4834));
    outputs(6435) <= (layer0_outputs(7138)) or (layer0_outputs(1417));
    outputs(6436) <= not((layer0_outputs(2398)) or (layer0_outputs(3715)));
    outputs(6437) <= (layer0_outputs(8617)) and (layer0_outputs(6305));
    outputs(6438) <= (layer0_outputs(9394)) xor (layer0_outputs(11194));
    outputs(6439) <= (layer0_outputs(10521)) and not (layer0_outputs(2692));
    outputs(6440) <= not(layer0_outputs(1101)) or (layer0_outputs(1547));
    outputs(6441) <= not((layer0_outputs(6428)) and (layer0_outputs(8615)));
    outputs(6442) <= layer0_outputs(9551);
    outputs(6443) <= not((layer0_outputs(6439)) xor (layer0_outputs(5164)));
    outputs(6444) <= not((layer0_outputs(3893)) xor (layer0_outputs(3660)));
    outputs(6445) <= layer0_outputs(9336);
    outputs(6446) <= (layer0_outputs(508)) xor (layer0_outputs(5521));
    outputs(6447) <= layer0_outputs(2217);
    outputs(6448) <= (layer0_outputs(12102)) xor (layer0_outputs(5547));
    outputs(6449) <= not(layer0_outputs(4386));
    outputs(6450) <= not(layer0_outputs(7645));
    outputs(6451) <= layer0_outputs(3718);
    outputs(6452) <= (layer0_outputs(9880)) xor (layer0_outputs(3982));
    outputs(6453) <= not((layer0_outputs(7668)) xor (layer0_outputs(5971)));
    outputs(6454) <= not(layer0_outputs(12228));
    outputs(6455) <= not(layer0_outputs(1766));
    outputs(6456) <= not(layer0_outputs(3991));
    outputs(6457) <= (layer0_outputs(11768)) and (layer0_outputs(1476));
    outputs(6458) <= not((layer0_outputs(1972)) and (layer0_outputs(2733)));
    outputs(6459) <= (layer0_outputs(7177)) xor (layer0_outputs(5348));
    outputs(6460) <= not(layer0_outputs(8211));
    outputs(6461) <= not(layer0_outputs(7509));
    outputs(6462) <= (layer0_outputs(2866)) and (layer0_outputs(2076));
    outputs(6463) <= (layer0_outputs(4499)) and (layer0_outputs(4015));
    outputs(6464) <= layer0_outputs(8492);
    outputs(6465) <= not(layer0_outputs(11195));
    outputs(6466) <= not(layer0_outputs(7028));
    outputs(6467) <= (layer0_outputs(9653)) and not (layer0_outputs(12564));
    outputs(6468) <= not(layer0_outputs(6738));
    outputs(6469) <= not(layer0_outputs(3252)) or (layer0_outputs(5731));
    outputs(6470) <= not(layer0_outputs(2278));
    outputs(6471) <= not((layer0_outputs(1321)) xor (layer0_outputs(10118)));
    outputs(6472) <= not(layer0_outputs(5498));
    outputs(6473) <= not(layer0_outputs(2162));
    outputs(6474) <= not((layer0_outputs(1080)) xor (layer0_outputs(11011)));
    outputs(6475) <= (layer0_outputs(9936)) xor (layer0_outputs(8628));
    outputs(6476) <= not(layer0_outputs(3177)) or (layer0_outputs(11028));
    outputs(6477) <= not((layer0_outputs(876)) or (layer0_outputs(1558)));
    outputs(6478) <= (layer0_outputs(3913)) xor (layer0_outputs(9738));
    outputs(6479) <= (layer0_outputs(5037)) and not (layer0_outputs(4255));
    outputs(6480) <= not(layer0_outputs(3308));
    outputs(6481) <= layer0_outputs(6941);
    outputs(6482) <= layer0_outputs(8620);
    outputs(6483) <= layer0_outputs(5868);
    outputs(6484) <= layer0_outputs(7963);
    outputs(6485) <= (layer0_outputs(4796)) or (layer0_outputs(5155));
    outputs(6486) <= not(layer0_outputs(12437));
    outputs(6487) <= not(layer0_outputs(12774));
    outputs(6488) <= layer0_outputs(6629);
    outputs(6489) <= (layer0_outputs(5240)) xor (layer0_outputs(8531));
    outputs(6490) <= not(layer0_outputs(10085)) or (layer0_outputs(12141));
    outputs(6491) <= not(layer0_outputs(10891));
    outputs(6492) <= (layer0_outputs(6775)) xor (layer0_outputs(9974));
    outputs(6493) <= (layer0_outputs(6837)) xor (layer0_outputs(10870));
    outputs(6494) <= (layer0_outputs(7841)) xor (layer0_outputs(3819));
    outputs(6495) <= (layer0_outputs(573)) and (layer0_outputs(11226));
    outputs(6496) <= not((layer0_outputs(2874)) xor (layer0_outputs(9740)));
    outputs(6497) <= (layer0_outputs(10205)) or (layer0_outputs(11115));
    outputs(6498) <= not(layer0_outputs(11905));
    outputs(6499) <= (layer0_outputs(10226)) xor (layer0_outputs(9403));
    outputs(6500) <= layer0_outputs(3077);
    outputs(6501) <= layer0_outputs(4864);
    outputs(6502) <= (layer0_outputs(6057)) xor (layer0_outputs(8841));
    outputs(6503) <= not((layer0_outputs(444)) xor (layer0_outputs(4201)));
    outputs(6504) <= (layer0_outputs(607)) xor (layer0_outputs(3764));
    outputs(6505) <= not(layer0_outputs(1488));
    outputs(6506) <= layer0_outputs(3192);
    outputs(6507) <= not((layer0_outputs(7721)) xor (layer0_outputs(2934)));
    outputs(6508) <= layer0_outputs(337);
    outputs(6509) <= (layer0_outputs(4217)) and not (layer0_outputs(7490));
    outputs(6510) <= layer0_outputs(8975);
    outputs(6511) <= layer0_outputs(263);
    outputs(6512) <= not((layer0_outputs(2605)) and (layer0_outputs(7785)));
    outputs(6513) <= (layer0_outputs(9266)) xor (layer0_outputs(9450));
    outputs(6514) <= not(layer0_outputs(7970));
    outputs(6515) <= not((layer0_outputs(4067)) xor (layer0_outputs(6500)));
    outputs(6516) <= not((layer0_outputs(11357)) or (layer0_outputs(325)));
    outputs(6517) <= not((layer0_outputs(2211)) xor (layer0_outputs(8475)));
    outputs(6518) <= (layer0_outputs(9975)) xor (layer0_outputs(4011));
    outputs(6519) <= (layer0_outputs(1479)) xor (layer0_outputs(1501));
    outputs(6520) <= layer0_outputs(2556);
    outputs(6521) <= (layer0_outputs(10170)) and not (layer0_outputs(10674));
    outputs(6522) <= (layer0_outputs(8448)) xor (layer0_outputs(1604));
    outputs(6523) <= layer0_outputs(2887);
    outputs(6524) <= not(layer0_outputs(2237));
    outputs(6525) <= not(layer0_outputs(128));
    outputs(6526) <= (layer0_outputs(7195)) xor (layer0_outputs(11246));
    outputs(6527) <= (layer0_outputs(11035)) xor (layer0_outputs(2138));
    outputs(6528) <= not(layer0_outputs(939));
    outputs(6529) <= not(layer0_outputs(7204)) or (layer0_outputs(12190));
    outputs(6530) <= (layer0_outputs(4113)) and (layer0_outputs(2450));
    outputs(6531) <= not((layer0_outputs(328)) xor (layer0_outputs(5489)));
    outputs(6532) <= not(layer0_outputs(10707)) or (layer0_outputs(4501));
    outputs(6533) <= not((layer0_outputs(3874)) xor (layer0_outputs(8497)));
    outputs(6534) <= layer0_outputs(6532);
    outputs(6535) <= (layer0_outputs(1523)) xor (layer0_outputs(8656));
    outputs(6536) <= layer0_outputs(3753);
    outputs(6537) <= (layer0_outputs(10939)) or (layer0_outputs(6737));
    outputs(6538) <= not(layer0_outputs(3424));
    outputs(6539) <= not(layer0_outputs(8003));
    outputs(6540) <= (layer0_outputs(8695)) xor (layer0_outputs(5893));
    outputs(6541) <= (layer0_outputs(3489)) and (layer0_outputs(11769));
    outputs(6542) <= layer0_outputs(5252);
    outputs(6543) <= layer0_outputs(11906);
    outputs(6544) <= not((layer0_outputs(3185)) and (layer0_outputs(9482)));
    outputs(6545) <= not((layer0_outputs(1051)) xor (layer0_outputs(5168)));
    outputs(6546) <= (layer0_outputs(11762)) xor (layer0_outputs(34));
    outputs(6547) <= (layer0_outputs(12006)) or (layer0_outputs(11911));
    outputs(6548) <= not(layer0_outputs(9496));
    outputs(6549) <= layer0_outputs(10487);
    outputs(6550) <= not(layer0_outputs(9195));
    outputs(6551) <= (layer0_outputs(11144)) xor (layer0_outputs(11722));
    outputs(6552) <= layer0_outputs(7862);
    outputs(6553) <= not(layer0_outputs(6875));
    outputs(6554) <= layer0_outputs(8888);
    outputs(6555) <= not(layer0_outputs(4974));
    outputs(6556) <= not(layer0_outputs(8421));
    outputs(6557) <= not(layer0_outputs(7730));
    outputs(6558) <= not(layer0_outputs(9226));
    outputs(6559) <= not(layer0_outputs(7821)) or (layer0_outputs(9177));
    outputs(6560) <= (layer0_outputs(5066)) xor (layer0_outputs(12329));
    outputs(6561) <= not((layer0_outputs(7706)) xor (layer0_outputs(2911)));
    outputs(6562) <= not((layer0_outputs(8066)) xor (layer0_outputs(1324)));
    outputs(6563) <= not(layer0_outputs(9170));
    outputs(6564) <= not((layer0_outputs(12765)) xor (layer0_outputs(11453)));
    outputs(6565) <= not(layer0_outputs(6118));
    outputs(6566) <= (layer0_outputs(4697)) and not (layer0_outputs(6151));
    outputs(6567) <= (layer0_outputs(12140)) xor (layer0_outputs(1540));
    outputs(6568) <= layer0_outputs(6668);
    outputs(6569) <= not(layer0_outputs(4464)) or (layer0_outputs(11091));
    outputs(6570) <= layer0_outputs(11344);
    outputs(6571) <= (layer0_outputs(6420)) xor (layer0_outputs(10688));
    outputs(6572) <= (layer0_outputs(11921)) xor (layer0_outputs(1004));
    outputs(6573) <= (layer0_outputs(3211)) xor (layer0_outputs(4689));
    outputs(6574) <= not((layer0_outputs(3093)) xor (layer0_outputs(5763)));
    outputs(6575) <= not(layer0_outputs(5481)) or (layer0_outputs(4312));
    outputs(6576) <= (layer0_outputs(12237)) or (layer0_outputs(1767));
    outputs(6577) <= layer0_outputs(4957);
    outputs(6578) <= not(layer0_outputs(9256)) or (layer0_outputs(4661));
    outputs(6579) <= not((layer0_outputs(11033)) xor (layer0_outputs(150)));
    outputs(6580) <= layer0_outputs(3611);
    outputs(6581) <= (layer0_outputs(4712)) and not (layer0_outputs(5851));
    outputs(6582) <= not((layer0_outputs(6716)) xor (layer0_outputs(3757)));
    outputs(6583) <= (layer0_outputs(2139)) or (layer0_outputs(4214));
    outputs(6584) <= not(layer0_outputs(1072));
    outputs(6585) <= (layer0_outputs(2307)) xor (layer0_outputs(2153));
    outputs(6586) <= (layer0_outputs(8364)) xor (layer0_outputs(12672));
    outputs(6587) <= layer0_outputs(4548);
    outputs(6588) <= not((layer0_outputs(9303)) xor (layer0_outputs(10110)));
    outputs(6589) <= not(layer0_outputs(12578));
    outputs(6590) <= layer0_outputs(10766);
    outputs(6591) <= not(layer0_outputs(110));
    outputs(6592) <= not(layer0_outputs(6950));
    outputs(6593) <= not((layer0_outputs(242)) xor (layer0_outputs(10570)));
    outputs(6594) <= not(layer0_outputs(4290));
    outputs(6595) <= (layer0_outputs(504)) xor (layer0_outputs(150));
    outputs(6596) <= layer0_outputs(98);
    outputs(6597) <= (layer0_outputs(1714)) xor (layer0_outputs(8989));
    outputs(6598) <= not(layer0_outputs(2099)) or (layer0_outputs(4608));
    outputs(6599) <= (layer0_outputs(3159)) xor (layer0_outputs(1699));
    outputs(6600) <= not((layer0_outputs(7686)) xor (layer0_outputs(4658)));
    outputs(6601) <= (layer0_outputs(106)) and not (layer0_outputs(9453));
    outputs(6602) <= (layer0_outputs(11582)) xor (layer0_outputs(1231));
    outputs(6603) <= not(layer0_outputs(10396));
    outputs(6604) <= layer0_outputs(2715);
    outputs(6605) <= not(layer0_outputs(9957)) or (layer0_outputs(535));
    outputs(6606) <= (layer0_outputs(9556)) xor (layer0_outputs(2552));
    outputs(6607) <= (layer0_outputs(9818)) and not (layer0_outputs(9717));
    outputs(6608) <= layer0_outputs(7750);
    outputs(6609) <= not(layer0_outputs(12094)) or (layer0_outputs(10614));
    outputs(6610) <= not((layer0_outputs(5539)) xor (layer0_outputs(8990)));
    outputs(6611) <= not(layer0_outputs(9311)) or (layer0_outputs(1189));
    outputs(6612) <= not(layer0_outputs(11843));
    outputs(6613) <= not(layer0_outputs(6257));
    outputs(6614) <= (layer0_outputs(8580)) xor (layer0_outputs(8738));
    outputs(6615) <= not(layer0_outputs(5982));
    outputs(6616) <= not((layer0_outputs(4722)) and (layer0_outputs(10642)));
    outputs(6617) <= layer0_outputs(10101);
    outputs(6618) <= not(layer0_outputs(10225)) or (layer0_outputs(7143));
    outputs(6619) <= (layer0_outputs(7867)) xor (layer0_outputs(12186));
    outputs(6620) <= (layer0_outputs(3511)) or (layer0_outputs(6661));
    outputs(6621) <= layer0_outputs(6134);
    outputs(6622) <= (layer0_outputs(11550)) or (layer0_outputs(5940));
    outputs(6623) <= (layer0_outputs(11377)) and not (layer0_outputs(8784));
    outputs(6624) <= not(layer0_outputs(8351));
    outputs(6625) <= (layer0_outputs(3465)) xor (layer0_outputs(3725));
    outputs(6626) <= (layer0_outputs(3237)) and (layer0_outputs(3323));
    outputs(6627) <= (layer0_outputs(8170)) xor (layer0_outputs(9493));
    outputs(6628) <= (layer0_outputs(1950)) and (layer0_outputs(6902));
    outputs(6629) <= (layer0_outputs(6072)) xor (layer0_outputs(2769));
    outputs(6630) <= not((layer0_outputs(12079)) xor (layer0_outputs(4281)));
    outputs(6631) <= not(layer0_outputs(26));
    outputs(6632) <= (layer0_outputs(5858)) or (layer0_outputs(718));
    outputs(6633) <= (layer0_outputs(6997)) xor (layer0_outputs(2530));
    outputs(6634) <= not(layer0_outputs(2130));
    outputs(6635) <= (layer0_outputs(9456)) xor (layer0_outputs(12035));
    outputs(6636) <= (layer0_outputs(9666)) xor (layer0_outputs(567));
    outputs(6637) <= not(layer0_outputs(4831));
    outputs(6638) <= not(layer0_outputs(4627));
    outputs(6639) <= not(layer0_outputs(11966));
    outputs(6640) <= layer0_outputs(6962);
    outputs(6641) <= (layer0_outputs(7530)) and (layer0_outputs(5140));
    outputs(6642) <= (layer0_outputs(9212)) and not (layer0_outputs(4023));
    outputs(6643) <= not((layer0_outputs(7493)) xor (layer0_outputs(253)));
    outputs(6644) <= (layer0_outputs(7154)) xor (layer0_outputs(3343));
    outputs(6645) <= not(layer0_outputs(1821));
    outputs(6646) <= not((layer0_outputs(12293)) xor (layer0_outputs(8463)));
    outputs(6647) <= layer0_outputs(1750);
    outputs(6648) <= not((layer0_outputs(869)) xor (layer0_outputs(9538)));
    outputs(6649) <= not(layer0_outputs(1780));
    outputs(6650) <= not((layer0_outputs(12412)) xor (layer0_outputs(2750)));
    outputs(6651) <= layer0_outputs(1423);
    outputs(6652) <= (layer0_outputs(9452)) xor (layer0_outputs(4044));
    outputs(6653) <= (layer0_outputs(7665)) and not (layer0_outputs(9411));
    outputs(6654) <= layer0_outputs(12085);
    outputs(6655) <= not((layer0_outputs(6904)) xor (layer0_outputs(12024)));
    outputs(6656) <= not(layer0_outputs(7783));
    outputs(6657) <= not(layer0_outputs(171));
    outputs(6658) <= not(layer0_outputs(7725)) or (layer0_outputs(6879));
    outputs(6659) <= (layer0_outputs(6227)) and not (layer0_outputs(11165));
    outputs(6660) <= not(layer0_outputs(2119));
    outputs(6661) <= not((layer0_outputs(1873)) xor (layer0_outputs(5630)));
    outputs(6662) <= not((layer0_outputs(3843)) or (layer0_outputs(2525)));
    outputs(6663) <= not(layer0_outputs(3773));
    outputs(6664) <= (layer0_outputs(8806)) xor (layer0_outputs(4651));
    outputs(6665) <= not((layer0_outputs(9752)) xor (layer0_outputs(5765)));
    outputs(6666) <= not(layer0_outputs(40));
    outputs(6667) <= not(layer0_outputs(2009));
    outputs(6668) <= not((layer0_outputs(2141)) xor (layer0_outputs(12144)));
    outputs(6669) <= (layer0_outputs(11381)) xor (layer0_outputs(2485));
    outputs(6670) <= not(layer0_outputs(754));
    outputs(6671) <= layer0_outputs(6731);
    outputs(6672) <= (layer0_outputs(8038)) xor (layer0_outputs(10540));
    outputs(6673) <= not(layer0_outputs(233));
    outputs(6674) <= (layer0_outputs(2295)) xor (layer0_outputs(4102));
    outputs(6675) <= layer0_outputs(5565);
    outputs(6676) <= (layer0_outputs(2382)) xor (layer0_outputs(2266));
    outputs(6677) <= layer0_outputs(2208);
    outputs(6678) <= not((layer0_outputs(995)) xor (layer0_outputs(1615)));
    outputs(6679) <= (layer0_outputs(8920)) xor (layer0_outputs(902));
    outputs(6680) <= (layer0_outputs(7579)) and not (layer0_outputs(6307));
    outputs(6681) <= (layer0_outputs(4932)) xor (layer0_outputs(10894));
    outputs(6682) <= not(layer0_outputs(7456));
    outputs(6683) <= (layer0_outputs(7353)) xor (layer0_outputs(11611));
    outputs(6684) <= layer0_outputs(2539);
    outputs(6685) <= layer0_outputs(3182);
    outputs(6686) <= (layer0_outputs(1856)) xor (layer0_outputs(4323));
    outputs(6687) <= layer0_outputs(8743);
    outputs(6688) <= not(layer0_outputs(11364));
    outputs(6689) <= (layer0_outputs(3090)) or (layer0_outputs(12502));
    outputs(6690) <= (layer0_outputs(1314)) and (layer0_outputs(4229));
    outputs(6691) <= not(layer0_outputs(9757));
    outputs(6692) <= not(layer0_outputs(4920));
    outputs(6693) <= not(layer0_outputs(8326));
    outputs(6694) <= (layer0_outputs(4287)) or (layer0_outputs(6680));
    outputs(6695) <= layer0_outputs(3684);
    outputs(6696) <= not((layer0_outputs(10102)) xor (layer0_outputs(4265)));
    outputs(6697) <= layer0_outputs(5803);
    outputs(6698) <= (layer0_outputs(11177)) or (layer0_outputs(6966));
    outputs(6699) <= not(layer0_outputs(5578));
    outputs(6700) <= layer0_outputs(7654);
    outputs(6701) <= layer0_outputs(4320);
    outputs(6702) <= (layer0_outputs(4656)) and not (layer0_outputs(3256));
    outputs(6703) <= not(layer0_outputs(7424));
    outputs(6704) <= layer0_outputs(9180);
    outputs(6705) <= not(layer0_outputs(9327));
    outputs(6706) <= not((layer0_outputs(7014)) xor (layer0_outputs(9209)));
    outputs(6707) <= not(layer0_outputs(969));
    outputs(6708) <= (layer0_outputs(83)) xor (layer0_outputs(4633));
    outputs(6709) <= not(layer0_outputs(3487));
    outputs(6710) <= layer0_outputs(11259);
    outputs(6711) <= not((layer0_outputs(864)) or (layer0_outputs(7473)));
    outputs(6712) <= not(layer0_outputs(7441));
    outputs(6713) <= layer0_outputs(5940);
    outputs(6714) <= layer0_outputs(9326);
    outputs(6715) <= not(layer0_outputs(7863)) or (layer0_outputs(8144));
    outputs(6716) <= not((layer0_outputs(10162)) or (layer0_outputs(2209)));
    outputs(6717) <= layer0_outputs(8404);
    outputs(6718) <= not(layer0_outputs(978));
    outputs(6719) <= not(layer0_outputs(5855)) or (layer0_outputs(4182));
    outputs(6720) <= (layer0_outputs(5659)) xor (layer0_outputs(398));
    outputs(6721) <= not(layer0_outputs(12565));
    outputs(6722) <= (layer0_outputs(11111)) xor (layer0_outputs(11755));
    outputs(6723) <= (layer0_outputs(6608)) xor (layer0_outputs(10420));
    outputs(6724) <= layer0_outputs(8181);
    outputs(6725) <= (layer0_outputs(10543)) xor (layer0_outputs(11666));
    outputs(6726) <= not(layer0_outputs(3199));
    outputs(6727) <= (layer0_outputs(2014)) xor (layer0_outputs(3817));
    outputs(6728) <= (layer0_outputs(11339)) and not (layer0_outputs(443));
    outputs(6729) <= not((layer0_outputs(3844)) xor (layer0_outputs(17)));
    outputs(6730) <= layer0_outputs(2719);
    outputs(6731) <= not(layer0_outputs(10069));
    outputs(6732) <= not(layer0_outputs(8865));
    outputs(6733) <= (layer0_outputs(8425)) xor (layer0_outputs(8527));
    outputs(6734) <= not(layer0_outputs(3110));
    outputs(6735) <= (layer0_outputs(1448)) xor (layer0_outputs(2382));
    outputs(6736) <= (layer0_outputs(6389)) xor (layer0_outputs(10126));
    outputs(6737) <= not(layer0_outputs(8420));
    outputs(6738) <= not((layer0_outputs(6345)) xor (layer0_outputs(2572)));
    outputs(6739) <= not(layer0_outputs(12760));
    outputs(6740) <= not(layer0_outputs(9679));
    outputs(6741) <= (layer0_outputs(8259)) or (layer0_outputs(9281));
    outputs(6742) <= layer0_outputs(10792);
    outputs(6743) <= not((layer0_outputs(5722)) or (layer0_outputs(449)));
    outputs(6744) <= not(layer0_outputs(4446)) or (layer0_outputs(9763));
    outputs(6745) <= layer0_outputs(10413);
    outputs(6746) <= not(layer0_outputs(11404));
    outputs(6747) <= (layer0_outputs(8315)) or (layer0_outputs(4509));
    outputs(6748) <= (layer0_outputs(10090)) xor (layer0_outputs(1907));
    outputs(6749) <= layer0_outputs(10054);
    outputs(6750) <= (layer0_outputs(12607)) or (layer0_outputs(8801));
    outputs(6751) <= layer0_outputs(6528);
    outputs(6752) <= not((layer0_outputs(9812)) xor (layer0_outputs(8384)));
    outputs(6753) <= (layer0_outputs(479)) and (layer0_outputs(11422));
    outputs(6754) <= layer0_outputs(8196);
    outputs(6755) <= layer0_outputs(904);
    outputs(6756) <= (layer0_outputs(9953)) or (layer0_outputs(3310));
    outputs(6757) <= (layer0_outputs(10082)) or (layer0_outputs(4342));
    outputs(6758) <= layer0_outputs(3019);
    outputs(6759) <= (layer0_outputs(6860)) xor (layer0_outputs(10192));
    outputs(6760) <= not(layer0_outputs(4773));
    outputs(6761) <= layer0_outputs(3003);
    outputs(6762) <= not(layer0_outputs(1596));
    outputs(6763) <= (layer0_outputs(12647)) or (layer0_outputs(1721));
    outputs(6764) <= not(layer0_outputs(5513));
    outputs(6765) <= layer0_outputs(1783);
    outputs(6766) <= (layer0_outputs(653)) xor (layer0_outputs(5839));
    outputs(6767) <= not(layer0_outputs(7161));
    outputs(6768) <= not((layer0_outputs(9347)) xor (layer0_outputs(5146)));
    outputs(6769) <= not((layer0_outputs(11671)) xor (layer0_outputs(351)));
    outputs(6770) <= (layer0_outputs(207)) xor (layer0_outputs(12353));
    outputs(6771) <= not(layer0_outputs(10564)) or (layer0_outputs(7507));
    outputs(6772) <= (layer0_outputs(795)) xor (layer0_outputs(3641));
    outputs(6773) <= layer0_outputs(10165);
    outputs(6774) <= not(layer0_outputs(2350)) or (layer0_outputs(11277));
    outputs(6775) <= not((layer0_outputs(12264)) xor (layer0_outputs(7917)));
    outputs(6776) <= (layer0_outputs(6934)) xor (layer0_outputs(5793));
    outputs(6777) <= not(layer0_outputs(7627));
    outputs(6778) <= layer0_outputs(9513);
    outputs(6779) <= not((layer0_outputs(11114)) xor (layer0_outputs(11756)));
    outputs(6780) <= (layer0_outputs(9168)) and not (layer0_outputs(2487));
    outputs(6781) <= (layer0_outputs(5785)) and not (layer0_outputs(913));
    outputs(6782) <= not(layer0_outputs(3973));
    outputs(6783) <= not(layer0_outputs(6515));
    outputs(6784) <= layer0_outputs(11625);
    outputs(6785) <= (layer0_outputs(11765)) and not (layer0_outputs(9834));
    outputs(6786) <= not(layer0_outputs(11827)) or (layer0_outputs(10249));
    outputs(6787) <= not(layer0_outputs(5790)) or (layer0_outputs(1555));
    outputs(6788) <= (layer0_outputs(862)) xor (layer0_outputs(7137));
    outputs(6789) <= layer0_outputs(2925);
    outputs(6790) <= (layer0_outputs(4350)) xor (layer0_outputs(468));
    outputs(6791) <= not(layer0_outputs(3143));
    outputs(6792) <= not(layer0_outputs(7826)) or (layer0_outputs(8891));
    outputs(6793) <= not(layer0_outputs(2878));
    outputs(6794) <= layer0_outputs(3423);
    outputs(6795) <= not((layer0_outputs(6233)) xor (layer0_outputs(4861)));
    outputs(6796) <= (layer0_outputs(11416)) xor (layer0_outputs(11971));
    outputs(6797) <= layer0_outputs(6907);
    outputs(6798) <= not(layer0_outputs(6840));
    outputs(6799) <= (layer0_outputs(5087)) or (layer0_outputs(4987));
    outputs(6800) <= layer0_outputs(1824);
    outputs(6801) <= not((layer0_outputs(801)) and (layer0_outputs(11291)));
    outputs(6802) <= not(layer0_outputs(7290)) or (layer0_outputs(2503));
    outputs(6803) <= (layer0_outputs(8522)) xor (layer0_outputs(1152));
    outputs(6804) <= (layer0_outputs(818)) xor (layer0_outputs(1025));
    outputs(6805) <= not(layer0_outputs(11960)) or (layer0_outputs(10018));
    outputs(6806) <= (layer0_outputs(2363)) xor (layer0_outputs(6290));
    outputs(6807) <= layer0_outputs(11182);
    outputs(6808) <= layer0_outputs(481);
    outputs(6809) <= not((layer0_outputs(10992)) xor (layer0_outputs(9584)));
    outputs(6810) <= not(layer0_outputs(4953));
    outputs(6811) <= (layer0_outputs(12612)) xor (layer0_outputs(11711));
    outputs(6812) <= (layer0_outputs(6024)) xor (layer0_outputs(4034));
    outputs(6813) <= (layer0_outputs(7455)) and not (layer0_outputs(9983));
    outputs(6814) <= (layer0_outputs(5204)) and not (layer0_outputs(11535));
    outputs(6815) <= (layer0_outputs(5882)) xor (layer0_outputs(1515));
    outputs(6816) <= layer0_outputs(12586);
    outputs(6817) <= (layer0_outputs(4382)) xor (layer0_outputs(6987));
    outputs(6818) <= not(layer0_outputs(7715)) or (layer0_outputs(6797));
    outputs(6819) <= not(layer0_outputs(9339));
    outputs(6820) <= not(layer0_outputs(7371));
    outputs(6821) <= (layer0_outputs(6090)) xor (layer0_outputs(2702));
    outputs(6822) <= not(layer0_outputs(12093));
    outputs(6823) <= not(layer0_outputs(54));
    outputs(6824) <= (layer0_outputs(2450)) and (layer0_outputs(2558));
    outputs(6825) <= not((layer0_outputs(9361)) xor (layer0_outputs(5700)));
    outputs(6826) <= (layer0_outputs(289)) and (layer0_outputs(8362));
    outputs(6827) <= not(layer0_outputs(5110));
    outputs(6828) <= (layer0_outputs(8023)) xor (layer0_outputs(1766));
    outputs(6829) <= not(layer0_outputs(12268));
    outputs(6830) <= (layer0_outputs(8451)) and not (layer0_outputs(3098));
    outputs(6831) <= layer0_outputs(11622);
    outputs(6832) <= not(layer0_outputs(8753));
    outputs(6833) <= (layer0_outputs(1335)) xor (layer0_outputs(6326));
    outputs(6834) <= not((layer0_outputs(12630)) xor (layer0_outputs(5627)));
    outputs(6835) <= (layer0_outputs(1548)) and not (layer0_outputs(3921));
    outputs(6836) <= (layer0_outputs(10958)) and not (layer0_outputs(1738));
    outputs(6837) <= not((layer0_outputs(1826)) xor (layer0_outputs(6205)));
    outputs(6838) <= layer0_outputs(10401);
    outputs(6839) <= (layer0_outputs(3255)) xor (layer0_outputs(6319));
    outputs(6840) <= not(layer0_outputs(12111));
    outputs(6841) <= not((layer0_outputs(8875)) xor (layer0_outputs(7371)));
    outputs(6842) <= layer0_outputs(909);
    outputs(6843) <= layer0_outputs(1962);
    outputs(6844) <= not((layer0_outputs(2108)) xor (layer0_outputs(8166)));
    outputs(6845) <= not(layer0_outputs(8041)) or (layer0_outputs(4227));
    outputs(6846) <= not(layer0_outputs(10187));
    outputs(6847) <= (layer0_outputs(8253)) xor (layer0_outputs(477));
    outputs(6848) <= not(layer0_outputs(10932));
    outputs(6849) <= not(layer0_outputs(4307));
    outputs(6850) <= layer0_outputs(12176);
    outputs(6851) <= (layer0_outputs(9607)) xor (layer0_outputs(10707));
    outputs(6852) <= layer0_outputs(6028);
    outputs(6853) <= (layer0_outputs(12297)) xor (layer0_outputs(6947));
    outputs(6854) <= layer0_outputs(5261);
    outputs(6855) <= not(layer0_outputs(5503));
    outputs(6856) <= not(layer0_outputs(8886));
    outputs(6857) <= layer0_outputs(3452);
    outputs(6858) <= layer0_outputs(5684);
    outputs(6859) <= layer0_outputs(3050);
    outputs(6860) <= not((layer0_outputs(12760)) xor (layer0_outputs(4598)));
    outputs(6861) <= layer0_outputs(7778);
    outputs(6862) <= (layer0_outputs(11172)) xor (layer0_outputs(7961));
    outputs(6863) <= not((layer0_outputs(8523)) xor (layer0_outputs(1439)));
    outputs(6864) <= not((layer0_outputs(11783)) xor (layer0_outputs(10292)));
    outputs(6865) <= layer0_outputs(4165);
    outputs(6866) <= not(layer0_outputs(9935));
    outputs(6867) <= (layer0_outputs(742)) or (layer0_outputs(3447));
    outputs(6868) <= not((layer0_outputs(9188)) xor (layer0_outputs(8670)));
    outputs(6869) <= (layer0_outputs(5735)) xor (layer0_outputs(10071));
    outputs(6870) <= not(layer0_outputs(10495));
    outputs(6871) <= not(layer0_outputs(10048));
    outputs(6872) <= not((layer0_outputs(10438)) xor (layer0_outputs(537)));
    outputs(6873) <= not((layer0_outputs(12327)) xor (layer0_outputs(3224)));
    outputs(6874) <= layer0_outputs(2736);
    outputs(6875) <= layer0_outputs(6035);
    outputs(6876) <= not(layer0_outputs(8510)) or (layer0_outputs(4160));
    outputs(6877) <= not(layer0_outputs(5260));
    outputs(6878) <= not(layer0_outputs(11725));
    outputs(6879) <= (layer0_outputs(10689)) and not (layer0_outputs(2668));
    outputs(6880) <= not(layer0_outputs(9292)) or (layer0_outputs(9694));
    outputs(6881) <= layer0_outputs(10940);
    outputs(6882) <= (layer0_outputs(6014)) xor (layer0_outputs(1606));
    outputs(6883) <= not(layer0_outputs(10134));
    outputs(6884) <= not(layer0_outputs(7641));
    outputs(6885) <= (layer0_outputs(8005)) xor (layer0_outputs(1858));
    outputs(6886) <= not(layer0_outputs(12593));
    outputs(6887) <= not((layer0_outputs(5970)) xor (layer0_outputs(1336)));
    outputs(6888) <= not(layer0_outputs(5164)) or (layer0_outputs(11346));
    outputs(6889) <= layer0_outputs(2814);
    outputs(6890) <= not(layer0_outputs(161));
    outputs(6891) <= layer0_outputs(437);
    outputs(6892) <= not(layer0_outputs(3663));
    outputs(6893) <= (layer0_outputs(10086)) xor (layer0_outputs(9249));
    outputs(6894) <= (layer0_outputs(229)) xor (layer0_outputs(599));
    outputs(6895) <= not(layer0_outputs(660));
    outputs(6896) <= layer0_outputs(9396);
    outputs(6897) <= not(layer0_outputs(10295)) or (layer0_outputs(4350));
    outputs(6898) <= not(layer0_outputs(6990));
    outputs(6899) <= not((layer0_outputs(11129)) xor (layer0_outputs(8831)));
    outputs(6900) <= (layer0_outputs(6297)) xor (layer0_outputs(8215));
    outputs(6901) <= not((layer0_outputs(6126)) xor (layer0_outputs(7236)));
    outputs(6902) <= not(layer0_outputs(10439)) or (layer0_outputs(9485));
    outputs(6903) <= (layer0_outputs(2214)) xor (layer0_outputs(5976));
    outputs(6904) <= not(layer0_outputs(10880));
    outputs(6905) <= (layer0_outputs(3134)) xor (layer0_outputs(12764));
    outputs(6906) <= not((layer0_outputs(2710)) xor (layer0_outputs(6084)));
    outputs(6907) <= not((layer0_outputs(5587)) or (layer0_outputs(12605)));
    outputs(6908) <= layer0_outputs(3508);
    outputs(6909) <= not(layer0_outputs(8214)) or (layer0_outputs(6578));
    outputs(6910) <= not((layer0_outputs(11492)) xor (layer0_outputs(559)));
    outputs(6911) <= layer0_outputs(11859);
    outputs(6912) <= not(layer0_outputs(12250));
    outputs(6913) <= not(layer0_outputs(2461));
    outputs(6914) <= not(layer0_outputs(1537));
    outputs(6915) <= not(layer0_outputs(8332));
    outputs(6916) <= not((layer0_outputs(12544)) xor (layer0_outputs(6368)));
    outputs(6917) <= (layer0_outputs(7558)) xor (layer0_outputs(5516));
    outputs(6918) <= not(layer0_outputs(12148)) or (layer0_outputs(7977));
    outputs(6919) <= not((layer0_outputs(2566)) or (layer0_outputs(11804)));
    outputs(6920) <= not(layer0_outputs(12491));
    outputs(6921) <= not(layer0_outputs(5563));
    outputs(6922) <= not((layer0_outputs(10294)) xor (layer0_outputs(4073)));
    outputs(6923) <= not(layer0_outputs(12615));
    outputs(6924) <= not(layer0_outputs(300));
    outputs(6925) <= not((layer0_outputs(11869)) or (layer0_outputs(1007)));
    outputs(6926) <= not(layer0_outputs(5625)) or (layer0_outputs(1269));
    outputs(6927) <= not((layer0_outputs(11338)) xor (layer0_outputs(1033)));
    outputs(6928) <= (layer0_outputs(6267)) xor (layer0_outputs(6957));
    outputs(6929) <= not(layer0_outputs(5208));
    outputs(6930) <= (layer0_outputs(11368)) xor (layer0_outputs(7542));
    outputs(6931) <= layer0_outputs(10834);
    outputs(6932) <= (layer0_outputs(1364)) and not (layer0_outputs(5091));
    outputs(6933) <= layer0_outputs(1405);
    outputs(6934) <= (layer0_outputs(10555)) and not (layer0_outputs(7120));
    outputs(6935) <= not((layer0_outputs(10370)) xor (layer0_outputs(1384)));
    outputs(6936) <= not(layer0_outputs(1319));
    outputs(6937) <= (layer0_outputs(7974)) or (layer0_outputs(5278));
    outputs(6938) <= (layer0_outputs(701)) xor (layer0_outputs(5855));
    outputs(6939) <= not(layer0_outputs(3431));
    outputs(6940) <= not(layer0_outputs(10362));
    outputs(6941) <= (layer0_outputs(9177)) or (layer0_outputs(6725));
    outputs(6942) <= not(layer0_outputs(4767));
    outputs(6943) <= (layer0_outputs(11820)) xor (layer0_outputs(10823));
    outputs(6944) <= (layer0_outputs(10158)) and not (layer0_outputs(11707));
    outputs(6945) <= not((layer0_outputs(2138)) or (layer0_outputs(5498)));
    outputs(6946) <= layer0_outputs(2772);
    outputs(6947) <= layer0_outputs(5026);
    outputs(6948) <= (layer0_outputs(11124)) xor (layer0_outputs(8109));
    outputs(6949) <= (layer0_outputs(9941)) xor (layer0_outputs(10031));
    outputs(6950) <= (layer0_outputs(1429)) or (layer0_outputs(2631));
    outputs(6951) <= (layer0_outputs(11561)) or (layer0_outputs(5052));
    outputs(6952) <= layer0_outputs(4028);
    outputs(6953) <= not((layer0_outputs(3393)) and (layer0_outputs(10566)));
    outputs(6954) <= not(layer0_outputs(11148));
    outputs(6955) <= not((layer0_outputs(2553)) xor (layer0_outputs(2984)));
    outputs(6956) <= (layer0_outputs(7811)) xor (layer0_outputs(11312));
    outputs(6957) <= not(layer0_outputs(5360)) or (layer0_outputs(9367));
    outputs(6958) <= layer0_outputs(10264);
    outputs(6959) <= (layer0_outputs(6055)) xor (layer0_outputs(501));
    outputs(6960) <= not(layer0_outputs(9165));
    outputs(6961) <= layer0_outputs(4657);
    outputs(6962) <= not((layer0_outputs(9863)) or (layer0_outputs(4558)));
    outputs(6963) <= not((layer0_outputs(5115)) xor (layer0_outputs(5076)));
    outputs(6964) <= not((layer0_outputs(3298)) xor (layer0_outputs(677)));
    outputs(6965) <= not((layer0_outputs(5167)) xor (layer0_outputs(12434)));
    outputs(6966) <= (layer0_outputs(3985)) xor (layer0_outputs(11223));
    outputs(6967) <= layer0_outputs(1435);
    outputs(6968) <= not(layer0_outputs(1387));
    outputs(6969) <= not((layer0_outputs(4316)) xor (layer0_outputs(6857)));
    outputs(6970) <= layer0_outputs(8072);
    outputs(6971) <= (layer0_outputs(8020)) xor (layer0_outputs(254));
    outputs(6972) <= not(layer0_outputs(808));
    outputs(6973) <= layer0_outputs(2880);
    outputs(6974) <= (layer0_outputs(4976)) and not (layer0_outputs(224));
    outputs(6975) <= not(layer0_outputs(3107));
    outputs(6976) <= layer0_outputs(5967);
    outputs(6977) <= not((layer0_outputs(11855)) or (layer0_outputs(4903)));
    outputs(6978) <= not((layer0_outputs(3078)) xor (layer0_outputs(4931)));
    outputs(6979) <= (layer0_outputs(9466)) and not (layer0_outputs(664));
    outputs(6980) <= (layer0_outputs(8798)) xor (layer0_outputs(7253));
    outputs(6981) <= layer0_outputs(1535);
    outputs(6982) <= layer0_outputs(5058);
    outputs(6983) <= layer0_outputs(11430);
    outputs(6984) <= not(layer0_outputs(2612));
    outputs(6985) <= (layer0_outputs(3902)) and (layer0_outputs(8292));
    outputs(6986) <= (layer0_outputs(5821)) and not (layer0_outputs(8833));
    outputs(6987) <= (layer0_outputs(4164)) xor (layer0_outputs(12367));
    outputs(6988) <= layer0_outputs(5422);
    outputs(6989) <= layer0_outputs(509);
    outputs(6990) <= layer0_outputs(11170);
    outputs(6991) <= not(layer0_outputs(8026));
    outputs(6992) <= not(layer0_outputs(1874));
    outputs(6993) <= not(layer0_outputs(10173));
    outputs(6994) <= (layer0_outputs(3025)) xor (layer0_outputs(7723));
    outputs(6995) <= not(layer0_outputs(2821));
    outputs(6996) <= not(layer0_outputs(6442));
    outputs(6997) <= not(layer0_outputs(12281)) or (layer0_outputs(10004));
    outputs(6998) <= (layer0_outputs(2538)) xor (layer0_outputs(5470));
    outputs(6999) <= not((layer0_outputs(10703)) xor (layer0_outputs(1947)));
    outputs(7000) <= (layer0_outputs(12378)) xor (layer0_outputs(4324));
    outputs(7001) <= not((layer0_outputs(4122)) or (layer0_outputs(12095)));
    outputs(7002) <= not((layer0_outputs(12443)) xor (layer0_outputs(3422)));
    outputs(7003) <= not((layer0_outputs(1325)) xor (layer0_outputs(11624)));
    outputs(7004) <= not(layer0_outputs(867));
    outputs(7005) <= not(layer0_outputs(5443)) or (layer0_outputs(11253));
    outputs(7006) <= not(layer0_outputs(10674));
    outputs(7007) <= (layer0_outputs(9241)) xor (layer0_outputs(2601));
    outputs(7008) <= not(layer0_outputs(4719));
    outputs(7009) <= (layer0_outputs(3481)) xor (layer0_outputs(2193));
    outputs(7010) <= not(layer0_outputs(575));
    outputs(7011) <= (layer0_outputs(12753)) and (layer0_outputs(9921));
    outputs(7012) <= (layer0_outputs(5084)) and (layer0_outputs(3272));
    outputs(7013) <= not(layer0_outputs(7381)) or (layer0_outputs(1932));
    outputs(7014) <= not((layer0_outputs(7796)) xor (layer0_outputs(12565)));
    outputs(7015) <= (layer0_outputs(1076)) xor (layer0_outputs(11139));
    outputs(7016) <= not((layer0_outputs(7376)) or (layer0_outputs(10640)));
    outputs(7017) <= (layer0_outputs(11841)) xor (layer0_outputs(3811));
    outputs(7018) <= not(layer0_outputs(5034));
    outputs(7019) <= not(layer0_outputs(1658));
    outputs(7020) <= layer0_outputs(3530);
    outputs(7021) <= not(layer0_outputs(6673));
    outputs(7022) <= not((layer0_outputs(5751)) xor (layer0_outputs(7369)));
    outputs(7023) <= layer0_outputs(10090);
    outputs(7024) <= (layer0_outputs(2761)) and not (layer0_outputs(11273));
    outputs(7025) <= not(layer0_outputs(9872));
    outputs(7026) <= (layer0_outputs(3031)) xor (layer0_outputs(322));
    outputs(7027) <= (layer0_outputs(5076)) xor (layer0_outputs(1445));
    outputs(7028) <= layer0_outputs(10035);
    outputs(7029) <= not((layer0_outputs(6296)) xor (layer0_outputs(10339)));
    outputs(7030) <= not((layer0_outputs(11681)) xor (layer0_outputs(8025)));
    outputs(7031) <= not((layer0_outputs(10523)) xor (layer0_outputs(9569)));
    outputs(7032) <= (layer0_outputs(4552)) and not (layer0_outputs(11706));
    outputs(7033) <= not(layer0_outputs(9250));
    outputs(7034) <= not((layer0_outputs(3853)) xor (layer0_outputs(506)));
    outputs(7035) <= (layer0_outputs(10623)) and not (layer0_outputs(5171));
    outputs(7036) <= (layer0_outputs(2785)) xor (layer0_outputs(2533));
    outputs(7037) <= (layer0_outputs(3286)) xor (layer0_outputs(9417));
    outputs(7038) <= (layer0_outputs(9994)) and not (layer0_outputs(248));
    outputs(7039) <= (layer0_outputs(8464)) xor (layer0_outputs(5067));
    outputs(7040) <= layer0_outputs(8927);
    outputs(7041) <= '1';
    outputs(7042) <= not((layer0_outputs(1735)) xor (layer0_outputs(2914)));
    outputs(7043) <= (layer0_outputs(9888)) or (layer0_outputs(7292));
    outputs(7044) <= (layer0_outputs(8272)) and not (layer0_outputs(10525));
    outputs(7045) <= not(layer0_outputs(4822));
    outputs(7046) <= not((layer0_outputs(4566)) xor (layer0_outputs(8489)));
    outputs(7047) <= layer0_outputs(6676);
    outputs(7048) <= not((layer0_outputs(1180)) xor (layer0_outputs(4480)));
    outputs(7049) <= (layer0_outputs(145)) or (layer0_outputs(12556));
    outputs(7050) <= (layer0_outputs(10713)) and not (layer0_outputs(167));
    outputs(7051) <= not(layer0_outputs(934));
    outputs(7052) <= not((layer0_outputs(11806)) or (layer0_outputs(10763)));
    outputs(7053) <= layer0_outputs(2621);
    outputs(7054) <= not((layer0_outputs(7818)) and (layer0_outputs(5322)));
    outputs(7055) <= not(layer0_outputs(6793));
    outputs(7056) <= not((layer0_outputs(186)) xor (layer0_outputs(8168)));
    outputs(7057) <= not((layer0_outputs(2018)) xor (layer0_outputs(6231)));
    outputs(7058) <= not((layer0_outputs(9231)) xor (layer0_outputs(11121)));
    outputs(7059) <= not(layer0_outputs(11930));
    outputs(7060) <= not(layer0_outputs(2435));
    outputs(7061) <= not((layer0_outputs(7109)) xor (layer0_outputs(6036)));
    outputs(7062) <= (layer0_outputs(7459)) and (layer0_outputs(7488));
    outputs(7063) <= layer0_outputs(12117);
    outputs(7064) <= layer0_outputs(9071);
    outputs(7065) <= not((layer0_outputs(8244)) xor (layer0_outputs(4581)));
    outputs(7066) <= not(layer0_outputs(3847));
    outputs(7067) <= not(layer0_outputs(4094));
    outputs(7068) <= layer0_outputs(2748);
    outputs(7069) <= layer0_outputs(1305);
    outputs(7070) <= not(layer0_outputs(9320));
    outputs(7071) <= not((layer0_outputs(7768)) and (layer0_outputs(11713)));
    outputs(7072) <= not(layer0_outputs(7551));
    outputs(7073) <= not(layer0_outputs(643));
    outputs(7074) <= not(layer0_outputs(12514));
    outputs(7075) <= not((layer0_outputs(5383)) xor (layer0_outputs(3004)));
    outputs(7076) <= layer0_outputs(9594);
    outputs(7077) <= not((layer0_outputs(10905)) xor (layer0_outputs(6732)));
    outputs(7078) <= layer0_outputs(7259);
    outputs(7079) <= not((layer0_outputs(9912)) xor (layer0_outputs(8455)));
    outputs(7080) <= not(layer0_outputs(5704));
    outputs(7081) <= not(layer0_outputs(2815)) or (layer0_outputs(3678));
    outputs(7082) <= not(layer0_outputs(9383));
    outputs(7083) <= layer0_outputs(12410);
    outputs(7084) <= layer0_outputs(9747);
    outputs(7085) <= layer0_outputs(279);
    outputs(7086) <= (layer0_outputs(8661)) xor (layer0_outputs(3125));
    outputs(7087) <= (layer0_outputs(6192)) xor (layer0_outputs(933));
    outputs(7088) <= not((layer0_outputs(1706)) xor (layer0_outputs(4934)));
    outputs(7089) <= layer0_outputs(10916);
    outputs(7090) <= layer0_outputs(12493);
    outputs(7091) <= (layer0_outputs(4264)) xor (layer0_outputs(5189));
    outputs(7092) <= not((layer0_outputs(4053)) xor (layer0_outputs(12396)));
    outputs(7093) <= layer0_outputs(8380);
    outputs(7094) <= (layer0_outputs(6146)) xor (layer0_outputs(12190));
    outputs(7095) <= not((layer0_outputs(8307)) xor (layer0_outputs(5629)));
    outputs(7096) <= not(layer0_outputs(1853));
    outputs(7097) <= not((layer0_outputs(2302)) xor (layer0_outputs(7105)));
    outputs(7098) <= (layer0_outputs(10331)) and not (layer0_outputs(7681));
    outputs(7099) <= (layer0_outputs(1695)) and not (layer0_outputs(12007));
    outputs(7100) <= not((layer0_outputs(9032)) xor (layer0_outputs(12740)));
    outputs(7101) <= not(layer0_outputs(7975)) or (layer0_outputs(9019));
    outputs(7102) <= layer0_outputs(11867);
    outputs(7103) <= (layer0_outputs(1770)) xor (layer0_outputs(8549));
    outputs(7104) <= layer0_outputs(6889);
    outputs(7105) <= layer0_outputs(246);
    outputs(7106) <= (layer0_outputs(211)) and not (layer0_outputs(10494));
    outputs(7107) <= not(layer0_outputs(6917));
    outputs(7108) <= layer0_outputs(5372);
    outputs(7109) <= not(layer0_outputs(480)) or (layer0_outputs(5297));
    outputs(7110) <= not((layer0_outputs(2113)) xor (layer0_outputs(4726)));
    outputs(7111) <= not(layer0_outputs(2964));
    outputs(7112) <= not(layer0_outputs(9098));
    outputs(7113) <= not((layer0_outputs(12467)) xor (layer0_outputs(7301)));
    outputs(7114) <= not((layer0_outputs(5163)) and (layer0_outputs(8672)));
    outputs(7115) <= (layer0_outputs(10084)) xor (layer0_outputs(10250));
    outputs(7116) <= not((layer0_outputs(6385)) and (layer0_outputs(2679)));
    outputs(7117) <= (layer0_outputs(7346)) and not (layer0_outputs(11083));
    outputs(7118) <= not(layer0_outputs(10149));
    outputs(7119) <= not((layer0_outputs(3054)) xor (layer0_outputs(9942)));
    outputs(7120) <= not((layer0_outputs(7033)) xor (layer0_outputs(1046)));
    outputs(7121) <= (layer0_outputs(3602)) or (layer0_outputs(11395));
    outputs(7122) <= not(layer0_outputs(4039)) or (layer0_outputs(4761));
    outputs(7123) <= not((layer0_outputs(3689)) xor (layer0_outputs(7860)));
    outputs(7124) <= layer0_outputs(11441);
    outputs(7125) <= not((layer0_outputs(1593)) xor (layer0_outputs(5556)));
    outputs(7126) <= (layer0_outputs(5108)) and not (layer0_outputs(3636));
    outputs(7127) <= (layer0_outputs(3459)) xor (layer0_outputs(4169));
    outputs(7128) <= (layer0_outputs(5665)) xor (layer0_outputs(8516));
    outputs(7129) <= layer0_outputs(11381);
    outputs(7130) <= (layer0_outputs(4904)) xor (layer0_outputs(11700));
    outputs(7131) <= (layer0_outputs(4363)) xor (layer0_outputs(11302));
    outputs(7132) <= layer0_outputs(6063);
    outputs(7133) <= layer0_outputs(778);
    outputs(7134) <= not(layer0_outputs(6219));
    outputs(7135) <= not((layer0_outputs(10157)) or (layer0_outputs(4396)));
    outputs(7136) <= (layer0_outputs(11125)) xor (layer0_outputs(949));
    outputs(7137) <= not((layer0_outputs(7517)) xor (layer0_outputs(1440)));
    outputs(7138) <= not(layer0_outputs(8907));
    outputs(7139) <= layer0_outputs(9318);
    outputs(7140) <= (layer0_outputs(1697)) and (layer0_outputs(11370));
    outputs(7141) <= (layer0_outputs(11185)) xor (layer0_outputs(8351));
    outputs(7142) <= not(layer0_outputs(10236));
    outputs(7143) <= not((layer0_outputs(10196)) or (layer0_outputs(10617)));
    outputs(7144) <= not(layer0_outputs(9352));
    outputs(7145) <= layer0_outputs(9028);
    outputs(7146) <= (layer0_outputs(5047)) or (layer0_outputs(11851));
    outputs(7147) <= layer0_outputs(4882);
    outputs(7148) <= layer0_outputs(6241);
    outputs(7149) <= not((layer0_outputs(1664)) xor (layer0_outputs(11754)));
    outputs(7150) <= not(layer0_outputs(705));
    outputs(7151) <= layer0_outputs(7356);
    outputs(7152) <= (layer0_outputs(893)) xor (layer0_outputs(6543));
    outputs(7153) <= layer0_outputs(5402);
    outputs(7154) <= not(layer0_outputs(7589));
    outputs(7155) <= not(layer0_outputs(2223));
    outputs(7156) <= layer0_outputs(6126);
    outputs(7157) <= not((layer0_outputs(9188)) or (layer0_outputs(11853)));
    outputs(7158) <= layer0_outputs(5068);
    outputs(7159) <= (layer0_outputs(3057)) and not (layer0_outputs(2318));
    outputs(7160) <= not((layer0_outputs(9016)) and (layer0_outputs(4964)));
    outputs(7161) <= not((layer0_outputs(3562)) xor (layer0_outputs(5739)));
    outputs(7162) <= (layer0_outputs(6071)) or (layer0_outputs(12391));
    outputs(7163) <= (layer0_outputs(2727)) and not (layer0_outputs(8231));
    outputs(7164) <= not((layer0_outputs(2920)) xor (layer0_outputs(92)));
    outputs(7165) <= layer0_outputs(11258);
    outputs(7166) <= (layer0_outputs(4603)) xor (layer0_outputs(4230));
    outputs(7167) <= layer0_outputs(10422);
    outputs(7168) <= (layer0_outputs(3677)) or (layer0_outputs(4896));
    outputs(7169) <= not((layer0_outputs(4439)) and (layer0_outputs(9691)));
    outputs(7170) <= not((layer0_outputs(3751)) xor (layer0_outputs(3756)));
    outputs(7171) <= not(layer0_outputs(1984));
    outputs(7172) <= (layer0_outputs(6208)) xor (layer0_outputs(3012));
    outputs(7173) <= layer0_outputs(9108);
    outputs(7174) <= not((layer0_outputs(12562)) xor (layer0_outputs(12710)));
    outputs(7175) <= not(layer0_outputs(7070)) or (layer0_outputs(1763));
    outputs(7176) <= not(layer0_outputs(11404));
    outputs(7177) <= not((layer0_outputs(1142)) and (layer0_outputs(9687)));
    outputs(7178) <= not((layer0_outputs(7736)) and (layer0_outputs(10129)));
    outputs(7179) <= not(layer0_outputs(3225));
    outputs(7180) <= not(layer0_outputs(8145));
    outputs(7181) <= (layer0_outputs(8209)) xor (layer0_outputs(2391));
    outputs(7182) <= layer0_outputs(10556);
    outputs(7183) <= layer0_outputs(10601);
    outputs(7184) <= (layer0_outputs(10611)) and not (layer0_outputs(829));
    outputs(7185) <= not(layer0_outputs(3446));
    outputs(7186) <= (layer0_outputs(1571)) or (layer0_outputs(8205));
    outputs(7187) <= layer0_outputs(6565);
    outputs(7188) <= not(layer0_outputs(9205));
    outputs(7189) <= layer0_outputs(10874);
    outputs(7190) <= not((layer0_outputs(4530)) xor (layer0_outputs(108)));
    outputs(7191) <= (layer0_outputs(8051)) xor (layer0_outputs(2396));
    outputs(7192) <= (layer0_outputs(9815)) xor (layer0_outputs(4358));
    outputs(7193) <= (layer0_outputs(7401)) xor (layer0_outputs(2879));
    outputs(7194) <= not((layer0_outputs(1807)) xor (layer0_outputs(10017)));
    outputs(7195) <= not(layer0_outputs(10255));
    outputs(7196) <= not(layer0_outputs(5754));
    outputs(7197) <= layer0_outputs(10041);
    outputs(7198) <= layer0_outputs(1829);
    outputs(7199) <= not((layer0_outputs(4514)) xor (layer0_outputs(182)));
    outputs(7200) <= layer0_outputs(12121);
    outputs(7201) <= not((layer0_outputs(6998)) and (layer0_outputs(163)));
    outputs(7202) <= layer0_outputs(595);
    outputs(7203) <= layer0_outputs(11233);
    outputs(7204) <= layer0_outputs(10539);
    outputs(7205) <= not(layer0_outputs(1148));
    outputs(7206) <= not(layer0_outputs(3832)) or (layer0_outputs(8701));
    outputs(7207) <= '1';
    outputs(7208) <= not(layer0_outputs(6103));
    outputs(7209) <= (layer0_outputs(1149)) xor (layer0_outputs(7010));
    outputs(7210) <= (layer0_outputs(5567)) or (layer0_outputs(9087));
    outputs(7211) <= not(layer0_outputs(8505)) or (layer0_outputs(8548));
    outputs(7212) <= (layer0_outputs(3468)) xor (layer0_outputs(5025));
    outputs(7213) <= layer0_outputs(4142);
    outputs(7214) <= not(layer0_outputs(2477)) or (layer0_outputs(9670));
    outputs(7215) <= not((layer0_outputs(4916)) xor (layer0_outputs(4924)));
    outputs(7216) <= not(layer0_outputs(9214));
    outputs(7217) <= not(layer0_outputs(7023)) or (layer0_outputs(702));
    outputs(7218) <= (layer0_outputs(595)) and not (layer0_outputs(5485));
    outputs(7219) <= layer0_outputs(9868);
    outputs(7220) <= layer0_outputs(10686);
    outputs(7221) <= layer0_outputs(9127);
    outputs(7222) <= (layer0_outputs(10490)) xor (layer0_outputs(548));
    outputs(7223) <= (layer0_outputs(6498)) xor (layer0_outputs(2514));
    outputs(7224) <= not((layer0_outputs(6595)) xor (layer0_outputs(3030)));
    outputs(7225) <= not(layer0_outputs(3109));
    outputs(7226) <= (layer0_outputs(11116)) and not (layer0_outputs(11357));
    outputs(7227) <= layer0_outputs(1638);
    outputs(7228) <= not(layer0_outputs(2334));
    outputs(7229) <= (layer0_outputs(3707)) xor (layer0_outputs(371));
    outputs(7230) <= not(layer0_outputs(20));
    outputs(7231) <= not(layer0_outputs(9376)) or (layer0_outputs(12533));
    outputs(7232) <= (layer0_outputs(2615)) and not (layer0_outputs(6244));
    outputs(7233) <= not(layer0_outputs(6783));
    outputs(7234) <= layer0_outputs(12009);
    outputs(7235) <= not(layer0_outputs(2946));
    outputs(7236) <= (layer0_outputs(5375)) xor (layer0_outputs(7639));
    outputs(7237) <= not(layer0_outputs(8054));
    outputs(7238) <= not((layer0_outputs(4190)) xor (layer0_outputs(3416)));
    outputs(7239) <= (layer0_outputs(9874)) and not (layer0_outputs(12017));
    outputs(7240) <= not((layer0_outputs(10497)) and (layer0_outputs(2326)));
    outputs(7241) <= not(layer0_outputs(3042));
    outputs(7242) <= not(layer0_outputs(287));
    outputs(7243) <= layer0_outputs(1432);
    outputs(7244) <= not(layer0_outputs(9891)) or (layer0_outputs(3556));
    outputs(7245) <= (layer0_outputs(7905)) and not (layer0_outputs(665));
    outputs(7246) <= not(layer0_outputs(12362));
    outputs(7247) <= not(layer0_outputs(10808));
    outputs(7248) <= (layer0_outputs(154)) and not (layer0_outputs(7589));
    outputs(7249) <= not((layer0_outputs(6164)) xor (layer0_outputs(943)));
    outputs(7250) <= layer0_outputs(2720);
    outputs(7251) <= (layer0_outputs(9031)) xor (layer0_outputs(657));
    outputs(7252) <= not((layer0_outputs(6622)) or (layer0_outputs(9457)));
    outputs(7253) <= (layer0_outputs(5123)) and not (layer0_outputs(11348));
    outputs(7254) <= layer0_outputs(9314);
    outputs(7255) <= (layer0_outputs(10636)) xor (layer0_outputs(3146));
    outputs(7256) <= layer0_outputs(5100);
    outputs(7257) <= not(layer0_outputs(8057));
    outputs(7258) <= (layer0_outputs(12280)) and (layer0_outputs(8204));
    outputs(7259) <= not(layer0_outputs(2343)) or (layer0_outputs(513));
    outputs(7260) <= layer0_outputs(23);
    outputs(7261) <= layer0_outputs(11538);
    outputs(7262) <= (layer0_outputs(8940)) xor (layer0_outputs(4803));
    outputs(7263) <= layer0_outputs(10945);
    outputs(7264) <= (layer0_outputs(6164)) or (layer0_outputs(7786));
    outputs(7265) <= not(layer0_outputs(9218));
    outputs(7266) <= not(layer0_outputs(11502));
    outputs(7267) <= (layer0_outputs(8625)) xor (layer0_outputs(3432));
    outputs(7268) <= not((layer0_outputs(10597)) xor (layer0_outputs(11822)));
    outputs(7269) <= not((layer0_outputs(642)) xor (layer0_outputs(8887)));
    outputs(7270) <= not((layer0_outputs(6841)) xor (layer0_outputs(6769)));
    outputs(7271) <= (layer0_outputs(6973)) and (layer0_outputs(11686));
    outputs(7272) <= (layer0_outputs(6823)) and not (layer0_outputs(10549));
    outputs(7273) <= not(layer0_outputs(3724));
    outputs(7274) <= not((layer0_outputs(9802)) and (layer0_outputs(115)));
    outputs(7275) <= (layer0_outputs(6045)) xor (layer0_outputs(4943));
    outputs(7276) <= not(layer0_outputs(11341));
    outputs(7277) <= (layer0_outputs(11919)) xor (layer0_outputs(11339));
    outputs(7278) <= not(layer0_outputs(10760));
    outputs(7279) <= not((layer0_outputs(499)) xor (layer0_outputs(36)));
    outputs(7280) <= layer0_outputs(5087);
    outputs(7281) <= not((layer0_outputs(5998)) or (layer0_outputs(10893)));
    outputs(7282) <= not(layer0_outputs(6471)) or (layer0_outputs(4064));
    outputs(7283) <= not((layer0_outputs(5655)) or (layer0_outputs(6563)));
    outputs(7284) <= not((layer0_outputs(7129)) xor (layer0_outputs(3983)));
    outputs(7285) <= layer0_outputs(4670);
    outputs(7286) <= (layer0_outputs(3782)) and (layer0_outputs(7791));
    outputs(7287) <= layer0_outputs(4244);
    outputs(7288) <= layer0_outputs(7108);
    outputs(7289) <= not(layer0_outputs(11815));
    outputs(7290) <= (layer0_outputs(448)) xor (layer0_outputs(6036));
    outputs(7291) <= not(layer0_outputs(4341));
    outputs(7292) <= not(layer0_outputs(5351)) or (layer0_outputs(2998));
    outputs(7293) <= layer0_outputs(3319);
    outputs(7294) <= not(layer0_outputs(10000));
    outputs(7295) <= not(layer0_outputs(6961));
    outputs(7296) <= (layer0_outputs(2752)) and not (layer0_outputs(3908));
    outputs(7297) <= (layer0_outputs(2687)) xor (layer0_outputs(11872));
    outputs(7298) <= not(layer0_outputs(11632));
    outputs(7299) <= layer0_outputs(10802);
    outputs(7300) <= not((layer0_outputs(8029)) xor (layer0_outputs(293)));
    outputs(7301) <= '1';
    outputs(7302) <= (layer0_outputs(12409)) or (layer0_outputs(8682));
    outputs(7303) <= not((layer0_outputs(9515)) xor (layer0_outputs(940)));
    outputs(7304) <= (layer0_outputs(5594)) xor (layer0_outputs(3075));
    outputs(7305) <= (layer0_outputs(8341)) or (layer0_outputs(8135));
    outputs(7306) <= not((layer0_outputs(2834)) xor (layer0_outputs(5279)));
    outputs(7307) <= (layer0_outputs(3097)) or (layer0_outputs(11429));
    outputs(7308) <= not((layer0_outputs(12325)) xor (layer0_outputs(7565)));
    outputs(7309) <= (layer0_outputs(9050)) xor (layer0_outputs(11420));
    outputs(7310) <= not(layer0_outputs(7034));
    outputs(7311) <= layer0_outputs(7149);
    outputs(7312) <= not(layer0_outputs(84));
    outputs(7313) <= not(layer0_outputs(12746)) or (layer0_outputs(8399));
    outputs(7314) <= not(layer0_outputs(11419));
    outputs(7315) <= not((layer0_outputs(10058)) xor (layer0_outputs(9760)));
    outputs(7316) <= (layer0_outputs(12089)) xor (layer0_outputs(10553));
    outputs(7317) <= not((layer0_outputs(3925)) and (layer0_outputs(7592)));
    outputs(7318) <= (layer0_outputs(7420)) and not (layer0_outputs(10453));
    outputs(7319) <= layer0_outputs(3193);
    outputs(7320) <= not((layer0_outputs(8056)) xor (layer0_outputs(5915)));
    outputs(7321) <= not(layer0_outputs(1043)) or (layer0_outputs(9667));
    outputs(7322) <= not((layer0_outputs(8926)) and (layer0_outputs(7066)));
    outputs(7323) <= (layer0_outputs(8458)) xor (layer0_outputs(10457));
    outputs(7324) <= layer0_outputs(9610);
    outputs(7325) <= not(layer0_outputs(390));
    outputs(7326) <= not(layer0_outputs(12382));
    outputs(7327) <= not(layer0_outputs(6093));
    outputs(7328) <= (layer0_outputs(2429)) xor (layer0_outputs(10691));
    outputs(7329) <= layer0_outputs(4957);
    outputs(7330) <= not((layer0_outputs(7305)) or (layer0_outputs(6873)));
    outputs(7331) <= (layer0_outputs(4768)) and (layer0_outputs(5531));
    outputs(7332) <= not(layer0_outputs(9109)) or (layer0_outputs(6735));
    outputs(7333) <= layer0_outputs(211);
    outputs(7334) <= (layer0_outputs(6876)) xor (layer0_outputs(6924));
    outputs(7335) <= not((layer0_outputs(11589)) xor (layer0_outputs(4739)));
    outputs(7336) <= not(layer0_outputs(2516));
    outputs(7337) <= not((layer0_outputs(1509)) xor (layer0_outputs(12560)));
    outputs(7338) <= layer0_outputs(9761);
    outputs(7339) <= layer0_outputs(11813);
    outputs(7340) <= layer0_outputs(10463);
    outputs(7341) <= layer0_outputs(2248);
    outputs(7342) <= not(layer0_outputs(187)) or (layer0_outputs(3131));
    outputs(7343) <= not(layer0_outputs(6600));
    outputs(7344) <= (layer0_outputs(4001)) and not (layer0_outputs(10378));
    outputs(7345) <= (layer0_outputs(9382)) xor (layer0_outputs(2802));
    outputs(7346) <= not(layer0_outputs(4537));
    outputs(7347) <= (layer0_outputs(5937)) xor (layer0_outputs(3315));
    outputs(7348) <= layer0_outputs(4198);
    outputs(7349) <= (layer0_outputs(6137)) xor (layer0_outputs(2883));
    outputs(7350) <= layer0_outputs(1243);
    outputs(7351) <= not((layer0_outputs(11847)) xor (layer0_outputs(3126)));
    outputs(7352) <= (layer0_outputs(2104)) xor (layer0_outputs(9850));
    outputs(7353) <= not((layer0_outputs(10878)) xor (layer0_outputs(9227)));
    outputs(7354) <= not((layer0_outputs(5748)) xor (layer0_outputs(6397)));
    outputs(7355) <= layer0_outputs(10574);
    outputs(7356) <= (layer0_outputs(2200)) xor (layer0_outputs(8679));
    outputs(7357) <= (layer0_outputs(1734)) and not (layer0_outputs(8954));
    outputs(7358) <= layer0_outputs(4970);
    outputs(7359) <= (layer0_outputs(11278)) and not (layer0_outputs(8207));
    outputs(7360) <= not(layer0_outputs(3989));
    outputs(7361) <= not(layer0_outputs(5736));
    outputs(7362) <= (layer0_outputs(10584)) or (layer0_outputs(11359));
    outputs(7363) <= (layer0_outputs(3524)) xor (layer0_outputs(1130));
    outputs(7364) <= not((layer0_outputs(4816)) xor (layer0_outputs(3597)));
    outputs(7365) <= (layer0_outputs(12383)) or (layer0_outputs(804));
    outputs(7366) <= (layer0_outputs(9762)) and not (layer0_outputs(6531));
    outputs(7367) <= layer0_outputs(6868);
    outputs(7368) <= (layer0_outputs(12182)) xor (layer0_outputs(8591));
    outputs(7369) <= layer0_outputs(11034);
    outputs(7370) <= not((layer0_outputs(2144)) xor (layer0_outputs(1751)));
    outputs(7371) <= (layer0_outputs(1651)) xor (layer0_outputs(11094));
    outputs(7372) <= not((layer0_outputs(7157)) xor (layer0_outputs(10592)));
    outputs(7373) <= not((layer0_outputs(4333)) xor (layer0_outputs(4561)));
    outputs(7374) <= not((layer0_outputs(7018)) xor (layer0_outputs(9158)));
    outputs(7375) <= not(layer0_outputs(5253));
    outputs(7376) <= not((layer0_outputs(7124)) xor (layer0_outputs(6545)));
    outputs(7377) <= layer0_outputs(12492);
    outputs(7378) <= not(layer0_outputs(12075));
    outputs(7379) <= not((layer0_outputs(11122)) xor (layer0_outputs(12103)));
    outputs(7380) <= not((layer0_outputs(3470)) or (layer0_outputs(1207)));
    outputs(7381) <= layer0_outputs(11513);
    outputs(7382) <= not(layer0_outputs(6633));
    outputs(7383) <= layer0_outputs(1561);
    outputs(7384) <= (layer0_outputs(1709)) and not (layer0_outputs(11944));
    outputs(7385) <= not((layer0_outputs(2999)) xor (layer0_outputs(11798)));
    outputs(7386) <= not((layer0_outputs(10484)) xor (layer0_outputs(8353)));
    outputs(7387) <= (layer0_outputs(8253)) and (layer0_outputs(7928));
    outputs(7388) <= not(layer0_outputs(7809));
    outputs(7389) <= not((layer0_outputs(5472)) xor (layer0_outputs(12496)));
    outputs(7390) <= not(layer0_outputs(4836));
    outputs(7391) <= not(layer0_outputs(6986));
    outputs(7392) <= layer0_outputs(5718);
    outputs(7393) <= not((layer0_outputs(1192)) xor (layer0_outputs(7567)));
    outputs(7394) <= (layer0_outputs(786)) and not (layer0_outputs(7998));
    outputs(7395) <= layer0_outputs(9980);
    outputs(7396) <= (layer0_outputs(11445)) and (layer0_outputs(8936));
    outputs(7397) <= not(layer0_outputs(5435));
    outputs(7398) <= layer0_outputs(2976);
    outputs(7399) <= not((layer0_outputs(1115)) xor (layer0_outputs(5090)));
    outputs(7400) <= not(layer0_outputs(5216));
    outputs(7401) <= (layer0_outputs(7584)) and (layer0_outputs(259));
    outputs(7402) <= not((layer0_outputs(613)) and (layer0_outputs(2195)));
    outputs(7403) <= not(layer0_outputs(1830));
    outputs(7404) <= not(layer0_outputs(6195));
    outputs(7405) <= (layer0_outputs(4371)) xor (layer0_outputs(3518));
    outputs(7406) <= not((layer0_outputs(2112)) xor (layer0_outputs(9483)));
    outputs(7407) <= not(layer0_outputs(11917)) or (layer0_outputs(492));
    outputs(7408) <= not((layer0_outputs(1375)) xor (layer0_outputs(6977)));
    outputs(7409) <= (layer0_outputs(4698)) and (layer0_outputs(10781));
    outputs(7410) <= not(layer0_outputs(12637));
    outputs(7411) <= (layer0_outputs(4061)) xor (layer0_outputs(12433));
    outputs(7412) <= not(layer0_outputs(9053));
    outputs(7413) <= layer0_outputs(4283);
    outputs(7414) <= (layer0_outputs(8873)) and not (layer0_outputs(1454));
    outputs(7415) <= (layer0_outputs(5461)) xor (layer0_outputs(301));
    outputs(7416) <= layer0_outputs(10915);
    outputs(7417) <= not(layer0_outputs(9043));
    outputs(7418) <= not(layer0_outputs(3011));
    outputs(7419) <= layer0_outputs(11155);
    outputs(7420) <= not((layer0_outputs(7317)) xor (layer0_outputs(12196)));
    outputs(7421) <= not(layer0_outputs(5702)) or (layer0_outputs(2394));
    outputs(7422) <= layer0_outputs(585);
    outputs(7423) <= layer0_outputs(888);
    outputs(7424) <= not(layer0_outputs(7683));
    outputs(7425) <= (layer0_outputs(1890)) xor (layer0_outputs(6107));
    outputs(7426) <= not((layer0_outputs(11041)) xor (layer0_outputs(10178)));
    outputs(7427) <= not(layer0_outputs(2771)) or (layer0_outputs(8726));
    outputs(7428) <= (layer0_outputs(11247)) xor (layer0_outputs(1623));
    outputs(7429) <= (layer0_outputs(11819)) xor (layer0_outputs(9304));
    outputs(7430) <= '0';
    outputs(7431) <= (layer0_outputs(4898)) xor (layer0_outputs(7790));
    outputs(7432) <= layer0_outputs(10915);
    outputs(7433) <= (layer0_outputs(4518)) xor (layer0_outputs(1633));
    outputs(7434) <= not(layer0_outputs(2956));
    outputs(7435) <= layer0_outputs(2304);
    outputs(7436) <= not(layer0_outputs(7062));
    outputs(7437) <= not((layer0_outputs(9046)) xor (layer0_outputs(1704)));
    outputs(7438) <= not((layer0_outputs(11989)) xor (layer0_outputs(7625)));
    outputs(7439) <= not((layer0_outputs(9495)) xor (layer0_outputs(10392)));
    outputs(7440) <= not(layer0_outputs(7347));
    outputs(7441) <= layer0_outputs(11714);
    outputs(7442) <= not((layer0_outputs(12155)) xor (layer0_outputs(10821)));
    outputs(7443) <= not(layer0_outputs(5181));
    outputs(7444) <= layer0_outputs(6110);
    outputs(7445) <= not((layer0_outputs(7167)) xor (layer0_outputs(7220)));
    outputs(7446) <= not((layer0_outputs(6903)) xor (layer0_outputs(6287)));
    outputs(7447) <= not((layer0_outputs(2108)) or (layer0_outputs(113)));
    outputs(7448) <= not(layer0_outputs(12382)) or (layer0_outputs(117));
    outputs(7449) <= layer0_outputs(10095);
    outputs(7450) <= not((layer0_outputs(12312)) xor (layer0_outputs(12570)));
    outputs(7451) <= (layer0_outputs(2469)) xor (layer0_outputs(1166));
    outputs(7452) <= not((layer0_outputs(12516)) and (layer0_outputs(6862)));
    outputs(7453) <= (layer0_outputs(6534)) xor (layer0_outputs(75));
    outputs(7454) <= layer0_outputs(7296);
    outputs(7455) <= layer0_outputs(11697);
    outputs(7456) <= not((layer0_outputs(2168)) xor (layer0_outputs(7552)));
    outputs(7457) <= not((layer0_outputs(2210)) and (layer0_outputs(3749)));
    outputs(7458) <= layer0_outputs(7356);
    outputs(7459) <= layer0_outputs(12053);
    outputs(7460) <= layer0_outputs(7053);
    outputs(7461) <= not(layer0_outputs(10511));
    outputs(7462) <= (layer0_outputs(5617)) xor (layer0_outputs(9869));
    outputs(7463) <= not(layer0_outputs(3786));
    outputs(7464) <= (layer0_outputs(5490)) and not (layer0_outputs(10239));
    outputs(7465) <= (layer0_outputs(9843)) and not (layer0_outputs(4512));
    outputs(7466) <= (layer0_outputs(8856)) or (layer0_outputs(7677));
    outputs(7467) <= (layer0_outputs(6156)) and not (layer0_outputs(9232));
    outputs(7468) <= layer0_outputs(11947);
    outputs(7469) <= (layer0_outputs(6346)) xor (layer0_outputs(11727));
    outputs(7470) <= not((layer0_outputs(5245)) xor (layer0_outputs(2522)));
    outputs(7471) <= not(layer0_outputs(10414));
    outputs(7472) <= layer0_outputs(10289);
    outputs(7473) <= layer0_outputs(6513);
    outputs(7474) <= not(layer0_outputs(8328));
    outputs(7475) <= layer0_outputs(4576);
    outputs(7476) <= layer0_outputs(9850);
    outputs(7477) <= (layer0_outputs(10842)) and not (layer0_outputs(10458));
    outputs(7478) <= layer0_outputs(8042);
    outputs(7479) <= not((layer0_outputs(170)) or (layer0_outputs(3239)));
    outputs(7480) <= layer0_outputs(9921);
    outputs(7481) <= layer0_outputs(8557);
    outputs(7482) <= (layer0_outputs(11927)) and not (layer0_outputs(1892));
    outputs(7483) <= not(layer0_outputs(6858));
    outputs(7484) <= not((layer0_outputs(12705)) xor (layer0_outputs(1741)));
    outputs(7485) <= (layer0_outputs(7918)) xor (layer0_outputs(2256));
    outputs(7486) <= not(layer0_outputs(1270)) or (layer0_outputs(6606));
    outputs(7487) <= (layer0_outputs(174)) xor (layer0_outputs(1779));
    outputs(7488) <= layer0_outputs(12116);
    outputs(7489) <= not((layer0_outputs(9457)) or (layer0_outputs(7555)));
    outputs(7490) <= not((layer0_outputs(1255)) xor (layer0_outputs(11694)));
    outputs(7491) <= not(layer0_outputs(2512));
    outputs(7492) <= layer0_outputs(10360);
    outputs(7493) <= not((layer0_outputs(4617)) or (layer0_outputs(198)));
    outputs(7494) <= not((layer0_outputs(11178)) xor (layer0_outputs(9296)));
    outputs(7495) <= not((layer0_outputs(6819)) xor (layer0_outputs(1201)));
    outputs(7496) <= not(layer0_outputs(7737));
    outputs(7497) <= not(layer0_outputs(12576));
    outputs(7498) <= not(layer0_outputs(1836));
    outputs(7499) <= layer0_outputs(8976);
    outputs(7500) <= layer0_outputs(11663);
    outputs(7501) <= not(layer0_outputs(11713)) or (layer0_outputs(4131));
    outputs(7502) <= layer0_outputs(12542);
    outputs(7503) <= not(layer0_outputs(6607));
    outputs(7504) <= (layer0_outputs(9129)) and not (layer0_outputs(6698));
    outputs(7505) <= not((layer0_outputs(9064)) or (layer0_outputs(2364)));
    outputs(7506) <= not(layer0_outputs(11979));
    outputs(7507) <= not(layer0_outputs(6921));
    outputs(7508) <= not((layer0_outputs(6484)) xor (layer0_outputs(5904)));
    outputs(7509) <= not(layer0_outputs(9308));
    outputs(7510) <= (layer0_outputs(3223)) xor (layer0_outputs(1953));
    outputs(7511) <= not(layer0_outputs(10769)) or (layer0_outputs(3298));
    outputs(7512) <= layer0_outputs(3398);
    outputs(7513) <= not(layer0_outputs(6789));
    outputs(7514) <= (layer0_outputs(11575)) xor (layer0_outputs(5114));
    outputs(7515) <= layer0_outputs(9483);
    outputs(7516) <= not(layer0_outputs(6958)) or (layer0_outputs(873));
    outputs(7517) <= not(layer0_outputs(8303)) or (layer0_outputs(7318));
    outputs(7518) <= not(layer0_outputs(5273));
    outputs(7519) <= layer0_outputs(4927);
    outputs(7520) <= not((layer0_outputs(9178)) xor (layer0_outputs(3183)));
    outputs(7521) <= not((layer0_outputs(4055)) or (layer0_outputs(10477)));
    outputs(7522) <= (layer0_outputs(8517)) and not (layer0_outputs(8953));
    outputs(7523) <= not((layer0_outputs(2426)) xor (layer0_outputs(11446)));
    outputs(7524) <= (layer0_outputs(1813)) xor (layer0_outputs(1884));
    outputs(7525) <= (layer0_outputs(4256)) xor (layer0_outputs(5620));
    outputs(7526) <= not(layer0_outputs(10402));
    outputs(7527) <= (layer0_outputs(2381)) and not (layer0_outputs(6348));
    outputs(7528) <= not(layer0_outputs(6984)) or (layer0_outputs(8049));
    outputs(7529) <= not(layer0_outputs(8545));
    outputs(7530) <= layer0_outputs(9418);
    outputs(7531) <= (layer0_outputs(4458)) xor (layer0_outputs(10403));
    outputs(7532) <= not(layer0_outputs(11427));
    outputs(7533) <= not((layer0_outputs(57)) and (layer0_outputs(6648)));
    outputs(7534) <= (layer0_outputs(12234)) or (layer0_outputs(10344));
    outputs(7535) <= not(layer0_outputs(2627));
    outputs(7536) <= not((layer0_outputs(7499)) xor (layer0_outputs(6044)));
    outputs(7537) <= layer0_outputs(9159);
    outputs(7538) <= layer0_outputs(3590);
    outputs(7539) <= (layer0_outputs(9082)) xor (layer0_outputs(10528));
    outputs(7540) <= not(layer0_outputs(11114)) or (layer0_outputs(2062));
    outputs(7541) <= not(layer0_outputs(8395));
    outputs(7542) <= not((layer0_outputs(2862)) xor (layer0_outputs(388)));
    outputs(7543) <= layer0_outputs(12488);
    outputs(7544) <= layer0_outputs(4246);
    outputs(7545) <= (layer0_outputs(9280)) xor (layer0_outputs(9500));
    outputs(7546) <= (layer0_outputs(7739)) and not (layer0_outputs(8427));
    outputs(7547) <= (layer0_outputs(9290)) or (layer0_outputs(8525));
    outputs(7548) <= layer0_outputs(4474);
    outputs(7549) <= not(layer0_outputs(118));
    outputs(7550) <= (layer0_outputs(11945)) xor (layer0_outputs(2395));
    outputs(7551) <= not((layer0_outputs(12037)) and (layer0_outputs(7577)));
    outputs(7552) <= (layer0_outputs(10435)) or (layer0_outputs(8747));
    outputs(7553) <= layer0_outputs(12353);
    outputs(7554) <= not((layer0_outputs(8502)) xor (layer0_outputs(10901)));
    outputs(7555) <= (layer0_outputs(4308)) and not (layer0_outputs(8831));
    outputs(7556) <= not(layer0_outputs(8293));
    outputs(7557) <= not(layer0_outputs(12192)) or (layer0_outputs(4910));
    outputs(7558) <= layer0_outputs(2858);
    outputs(7559) <= not(layer0_outputs(8007));
    outputs(7560) <= not((layer0_outputs(7941)) and (layer0_outputs(7574)));
    outputs(7561) <= not(layer0_outputs(8923));
    outputs(7562) <= layer0_outputs(8705);
    outputs(7563) <= not(layer0_outputs(12028));
    outputs(7564) <= not((layer0_outputs(11804)) and (layer0_outputs(4203)));
    outputs(7565) <= not((layer0_outputs(10953)) or (layer0_outputs(10055)));
    outputs(7566) <= (layer0_outputs(7705)) xor (layer0_outputs(12277));
    outputs(7567) <= not((layer0_outputs(3915)) xor (layer0_outputs(10011)));
    outputs(7568) <= not((layer0_outputs(1720)) xor (layer0_outputs(7361)));
    outputs(7569) <= layer0_outputs(883);
    outputs(7570) <= (layer0_outputs(3719)) xor (layer0_outputs(7920));
    outputs(7571) <= (layer0_outputs(6625)) xor (layer0_outputs(3159));
    outputs(7572) <= (layer0_outputs(1272)) xor (layer0_outputs(8766));
    outputs(7573) <= not((layer0_outputs(6017)) xor (layer0_outputs(5907)));
    outputs(7574) <= (layer0_outputs(9492)) or (layer0_outputs(11459));
    outputs(7575) <= not(layer0_outputs(5624));
    outputs(7576) <= layer0_outputs(3755);
    outputs(7577) <= (layer0_outputs(5310)) or (layer0_outputs(10608));
    outputs(7578) <= layer0_outputs(7838);
    outputs(7579) <= not((layer0_outputs(12684)) or (layer0_outputs(5613)));
    outputs(7580) <= layer0_outputs(2599);
    outputs(7581) <= not((layer0_outputs(12734)) xor (layer0_outputs(4013)));
    outputs(7582) <= (layer0_outputs(7155)) and not (layer0_outputs(8056));
    outputs(7583) <= not(layer0_outputs(982));
    outputs(7584) <= (layer0_outputs(2098)) xor (layer0_outputs(686));
    outputs(7585) <= (layer0_outputs(5667)) and not (layer0_outputs(5742));
    outputs(7586) <= layer0_outputs(10503);
    outputs(7587) <= not(layer0_outputs(2314)) or (layer0_outputs(10616));
    outputs(7588) <= (layer0_outputs(9613)) xor (layer0_outputs(2538));
    outputs(7589) <= '0';
    outputs(7590) <= layer0_outputs(12257);
    outputs(7591) <= (layer0_outputs(10244)) xor (layer0_outputs(7340));
    outputs(7592) <= not((layer0_outputs(2838)) xor (layer0_outputs(11190)));
    outputs(7593) <= (layer0_outputs(6158)) xor (layer0_outputs(4586));
    outputs(7594) <= layer0_outputs(3303);
    outputs(7595) <= not((layer0_outputs(2738)) xor (layer0_outputs(11834)));
    outputs(7596) <= not((layer0_outputs(5421)) or (layer0_outputs(2753)));
    outputs(7597) <= layer0_outputs(4878);
    outputs(7598) <= layer0_outputs(10316);
    outputs(7599) <= not(layer0_outputs(11788)) or (layer0_outputs(3176));
    outputs(7600) <= (layer0_outputs(9141)) xor (layer0_outputs(12177));
    outputs(7601) <= not(layer0_outputs(908));
    outputs(7602) <= not((layer0_outputs(4544)) and (layer0_outputs(8694)));
    outputs(7603) <= not(layer0_outputs(10721));
    outputs(7604) <= not((layer0_outputs(9537)) and (layer0_outputs(6554)));
    outputs(7605) <= not(layer0_outputs(3118));
    outputs(7606) <= layer0_outputs(5337);
    outputs(7607) <= (layer0_outputs(11721)) xor (layer0_outputs(11466));
    outputs(7608) <= not((layer0_outputs(8044)) xor (layer0_outputs(12133)));
    outputs(7609) <= not(layer0_outputs(1369));
    outputs(7610) <= (layer0_outputs(11924)) xor (layer0_outputs(2704));
    outputs(7611) <= (layer0_outputs(1104)) and not (layer0_outputs(3170));
    outputs(7612) <= (layer0_outputs(9417)) xor (layer0_outputs(6996));
    outputs(7613) <= layer0_outputs(1324);
    outputs(7614) <= not((layer0_outputs(5454)) xor (layer0_outputs(8121)));
    outputs(7615) <= (layer0_outputs(7982)) and not (layer0_outputs(3051));
    outputs(7616) <= (layer0_outputs(12633)) and (layer0_outputs(256));
    outputs(7617) <= not(layer0_outputs(8948));
    outputs(7618) <= layer0_outputs(11477);
    outputs(7619) <= (layer0_outputs(11069)) xor (layer0_outputs(4665));
    outputs(7620) <= (layer0_outputs(4630)) xor (layer0_outputs(10006));
    outputs(7621) <= not(layer0_outputs(3585)) or (layer0_outputs(6527));
    outputs(7622) <= (layer0_outputs(10398)) xor (layer0_outputs(8626));
    outputs(7623) <= not((layer0_outputs(9640)) xor (layer0_outputs(10337)));
    outputs(7624) <= (layer0_outputs(9899)) xor (layer0_outputs(3215));
    outputs(7625) <= not(layer0_outputs(9789));
    outputs(7626) <= (layer0_outputs(810)) xor (layer0_outputs(10114));
    outputs(7627) <= (layer0_outputs(9582)) xor (layer0_outputs(2295));
    outputs(7628) <= layer0_outputs(3335);
    outputs(7629) <= not(layer0_outputs(1927));
    outputs(7630) <= (layer0_outputs(12089)) xor (layer0_outputs(9375));
    outputs(7631) <= not((layer0_outputs(641)) xor (layer0_outputs(4808)));
    outputs(7632) <= layer0_outputs(1677);
    outputs(7633) <= layer0_outputs(9081);
    outputs(7634) <= (layer0_outputs(2735)) or (layer0_outputs(5547));
    outputs(7635) <= not((layer0_outputs(2162)) and (layer0_outputs(2277)));
    outputs(7636) <= not(layer0_outputs(11503));
    outputs(7637) <= not(layer0_outputs(1385));
    outputs(7638) <= layer0_outputs(9400);
    outputs(7639) <= layer0_outputs(8470);
    outputs(7640) <= not((layer0_outputs(3032)) xor (layer0_outputs(9926)));
    outputs(7641) <= layer0_outputs(3457);
    outputs(7642) <= not(layer0_outputs(1843));
    outputs(7643) <= (layer0_outputs(7787)) xor (layer0_outputs(11832));
    outputs(7644) <= (layer0_outputs(10866)) and (layer0_outputs(4902));
    outputs(7645) <= not(layer0_outputs(5265));
    outputs(7646) <= layer0_outputs(1377);
    outputs(7647) <= not(layer0_outputs(3954)) or (layer0_outputs(298));
    outputs(7648) <= layer0_outputs(344);
    outputs(7649) <= (layer0_outputs(7184)) xor (layer0_outputs(7373));
    outputs(7650) <= not(layer0_outputs(3589)) or (layer0_outputs(6687));
    outputs(7651) <= layer0_outputs(10794);
    outputs(7652) <= layer0_outputs(3480);
    outputs(7653) <= (layer0_outputs(9487)) and not (layer0_outputs(3543));
    outputs(7654) <= layer0_outputs(821);
    outputs(7655) <= layer0_outputs(1314);
    outputs(7656) <= (layer0_outputs(3178)) xor (layer0_outputs(7586));
    outputs(7657) <= layer0_outputs(7882);
    outputs(7658) <= (layer0_outputs(9741)) and not (layer0_outputs(6743));
    outputs(7659) <= (layer0_outputs(7933)) xor (layer0_outputs(3667));
    outputs(7660) <= (layer0_outputs(5384)) xor (layer0_outputs(8816));
    outputs(7661) <= (layer0_outputs(9442)) xor (layer0_outputs(7664));
    outputs(7662) <= not(layer0_outputs(8675));
    outputs(7663) <= not((layer0_outputs(11138)) xor (layer0_outputs(4446)));
    outputs(7664) <= (layer0_outputs(6820)) xor (layer0_outputs(8252));
    outputs(7665) <= (layer0_outputs(1156)) xor (layer0_outputs(11514));
    outputs(7666) <= not((layer0_outputs(2745)) xor (layer0_outputs(11342)));
    outputs(7667) <= layer0_outputs(9191);
    outputs(7668) <= (layer0_outputs(1845)) xor (layer0_outputs(11048));
    outputs(7669) <= layer0_outputs(8533);
    outputs(7670) <= layer0_outputs(12792);
    outputs(7671) <= not(layer0_outputs(9697));
    outputs(7672) <= not((layer0_outputs(6197)) xor (layer0_outputs(5505)));
    outputs(7673) <= not(layer0_outputs(6806));
    outputs(7674) <= layer0_outputs(8569);
    outputs(7675) <= layer0_outputs(10515);
    outputs(7676) <= not(layer0_outputs(4462));
    outputs(7677) <= (layer0_outputs(11465)) xor (layer0_outputs(7290));
    outputs(7678) <= not(layer0_outputs(2199));
    outputs(7679) <= not(layer0_outputs(12327)) or (layer0_outputs(6460));
    outputs(7680) <= not(layer0_outputs(7859)) or (layer0_outputs(2021));
    outputs(7681) <= not(layer0_outputs(3775));
    outputs(7682) <= not(layer0_outputs(8940));
    outputs(7683) <= not((layer0_outputs(2945)) and (layer0_outputs(11226)));
    outputs(7684) <= not(layer0_outputs(1815));
    outputs(7685) <= layer0_outputs(7644);
    outputs(7686) <= layer0_outputs(7638);
    outputs(7687) <= (layer0_outputs(9308)) and not (layer0_outputs(10728));
    outputs(7688) <= layer0_outputs(7154);
    outputs(7689) <= layer0_outputs(5064);
    outputs(7690) <= not(layer0_outputs(10244));
    outputs(7691) <= not(layer0_outputs(12314));
    outputs(7692) <= (layer0_outputs(10092)) xor (layer0_outputs(3863));
    outputs(7693) <= layer0_outputs(448);
    outputs(7694) <= not(layer0_outputs(10118));
    outputs(7695) <= (layer0_outputs(8157)) xor (layer0_outputs(12227));
    outputs(7696) <= layer0_outputs(6422);
    outputs(7697) <= not((layer0_outputs(5776)) xor (layer0_outputs(11531)));
    outputs(7698) <= not(layer0_outputs(6747));
    outputs(7699) <= (layer0_outputs(4903)) xor (layer0_outputs(1567));
    outputs(7700) <= not(layer0_outputs(4049));
    outputs(7701) <= layer0_outputs(9612);
    outputs(7702) <= layer0_outputs(2881);
    outputs(7703) <= (layer0_outputs(6906)) xor (layer0_outputs(11011));
    outputs(7704) <= not((layer0_outputs(11534)) or (layer0_outputs(12326)));
    outputs(7705) <= layer0_outputs(212);
    outputs(7706) <= (layer0_outputs(6179)) and not (layer0_outputs(8687));
    outputs(7707) <= (layer0_outputs(2376)) xor (layer0_outputs(12278));
    outputs(7708) <= (layer0_outputs(11472)) and (layer0_outputs(11022));
    outputs(7709) <= layer0_outputs(10431);
    outputs(7710) <= not(layer0_outputs(9278));
    outputs(7711) <= (layer0_outputs(2726)) and not (layer0_outputs(9682));
    outputs(7712) <= (layer0_outputs(5442)) xor (layer0_outputs(7261));
    outputs(7713) <= (layer0_outputs(5955)) xor (layer0_outputs(6504));
    outputs(7714) <= not((layer0_outputs(2374)) xor (layer0_outputs(2160)));
    outputs(7715) <= not(layer0_outputs(7662));
    outputs(7716) <= layer0_outputs(6004);
    outputs(7717) <= not(layer0_outputs(10312));
    outputs(7718) <= not(layer0_outputs(5553));
    outputs(7719) <= not((layer0_outputs(6287)) xor (layer0_outputs(11870)));
    outputs(7720) <= not(layer0_outputs(7502));
    outputs(7721) <= not(layer0_outputs(4634));
    outputs(7722) <= not((layer0_outputs(3425)) or (layer0_outputs(1442)));
    outputs(7723) <= (layer0_outputs(4850)) and not (layer0_outputs(2713));
    outputs(7724) <= (layer0_outputs(8267)) and not (layer0_outputs(11828));
    outputs(7725) <= not(layer0_outputs(643));
    outputs(7726) <= layer0_outputs(345);
    outputs(7727) <= (layer0_outputs(10861)) xor (layer0_outputs(8585));
    outputs(7728) <= not(layer0_outputs(1306));
    outputs(7729) <= not(layer0_outputs(935));
    outputs(7730) <= not((layer0_outputs(5904)) xor (layer0_outputs(9023)));
    outputs(7731) <= not((layer0_outputs(4639)) or (layer0_outputs(1645)));
    outputs(7732) <= layer0_outputs(8892);
    outputs(7733) <= (layer0_outputs(3080)) xor (layer0_outputs(3727));
    outputs(7734) <= layer0_outputs(9678);
    outputs(7735) <= layer0_outputs(1242);
    outputs(7736) <= layer0_outputs(9115);
    outputs(7737) <= layer0_outputs(9518);
    outputs(7738) <= not((layer0_outputs(5418)) xor (layer0_outputs(181)));
    outputs(7739) <= not(layer0_outputs(10751)) or (layer0_outputs(11046));
    outputs(7740) <= layer0_outputs(8739);
    outputs(7741) <= layer0_outputs(3186);
    outputs(7742) <= layer0_outputs(6016);
    outputs(7743) <= not((layer0_outputs(2589)) or (layer0_outputs(10929)));
    outputs(7744) <= not(layer0_outputs(12063));
    outputs(7745) <= not(layer0_outputs(3933));
    outputs(7746) <= layer0_outputs(11573);
    outputs(7747) <= not(layer0_outputs(11783)) or (layer0_outputs(4352));
    outputs(7748) <= not(layer0_outputs(8347));
    outputs(7749) <= layer0_outputs(7277);
    outputs(7750) <= layer0_outputs(4498);
    outputs(7751) <= not((layer0_outputs(5699)) and (layer0_outputs(4942)));
    outputs(7752) <= layer0_outputs(597);
    outputs(7753) <= not(layer0_outputs(7663)) or (layer0_outputs(281));
    outputs(7754) <= (layer0_outputs(7638)) xor (layer0_outputs(347));
    outputs(7755) <= (layer0_outputs(12401)) xor (layer0_outputs(989));
    outputs(7756) <= (layer0_outputs(911)) xor (layer0_outputs(10841));
    outputs(7757) <= not(layer0_outputs(2547)) or (layer0_outputs(2821));
    outputs(7758) <= (layer0_outputs(2595)) xor (layer0_outputs(7132));
    outputs(7759) <= layer0_outputs(5789);
    outputs(7760) <= not((layer0_outputs(6804)) xor (layer0_outputs(551)));
    outputs(7761) <= (layer0_outputs(10242)) xor (layer0_outputs(7064));
    outputs(7762) <= not(layer0_outputs(7569));
    outputs(7763) <= layer0_outputs(62);
    outputs(7764) <= (layer0_outputs(9769)) and not (layer0_outputs(3099));
    outputs(7765) <= not(layer0_outputs(5039));
    outputs(7766) <= not((layer0_outputs(8900)) and (layer0_outputs(6912)));
    outputs(7767) <= layer0_outputs(10635);
    outputs(7768) <= (layer0_outputs(2255)) xor (layer0_outputs(8007));
    outputs(7769) <= not(layer0_outputs(2678));
    outputs(7770) <= not(layer0_outputs(4925));
    outputs(7771) <= layer0_outputs(7907);
    outputs(7772) <= not(layer0_outputs(8357));
    outputs(7773) <= not(layer0_outputs(4196));
    outputs(7774) <= not(layer0_outputs(4792));
    outputs(7775) <= layer0_outputs(11578);
    outputs(7776) <= not(layer0_outputs(9949));
    outputs(7777) <= (layer0_outputs(3481)) xor (layer0_outputs(6406));
    outputs(7778) <= (layer0_outputs(7048)) xor (layer0_outputs(3262));
    outputs(7779) <= not(layer0_outputs(411));
    outputs(7780) <= layer0_outputs(7331);
    outputs(7781) <= layer0_outputs(7122);
    outputs(7782) <= not(layer0_outputs(10848));
    outputs(7783) <= (layer0_outputs(12751)) or (layer0_outputs(587));
    outputs(7784) <= layer0_outputs(2694);
    outputs(7785) <= not((layer0_outputs(5887)) and (layer0_outputs(2086)));
    outputs(7786) <= layer0_outputs(7642);
    outputs(7787) <= not(layer0_outputs(4919));
    outputs(7788) <= not(layer0_outputs(7922));
    outputs(7789) <= not(layer0_outputs(3545));
    outputs(7790) <= (layer0_outputs(8905)) xor (layer0_outputs(3572));
    outputs(7791) <= not((layer0_outputs(8992)) or (layer0_outputs(2186)));
    outputs(7792) <= not((layer0_outputs(10377)) or (layer0_outputs(11677)));
    outputs(7793) <= not(layer0_outputs(6953));
    outputs(7794) <= not(layer0_outputs(8097));
    outputs(7795) <= (layer0_outputs(4175)) and not (layer0_outputs(12377));
    outputs(7796) <= not(layer0_outputs(6408)) or (layer0_outputs(5009));
    outputs(7797) <= not(layer0_outputs(834));
    outputs(7798) <= layer0_outputs(12503);
    outputs(7799) <= not(layer0_outputs(5867));
    outputs(7800) <= not(layer0_outputs(4134));
    outputs(7801) <= not(layer0_outputs(12529)) or (layer0_outputs(7942));
    outputs(7802) <= layer0_outputs(9010);
    outputs(7803) <= layer0_outputs(11485);
    outputs(7804) <= not((layer0_outputs(4980)) or (layer0_outputs(2962)));
    outputs(7805) <= (layer0_outputs(2293)) xor (layer0_outputs(9183));
    outputs(7806) <= not((layer0_outputs(69)) or (layer0_outputs(10195)));
    outputs(7807) <= layer0_outputs(89);
    outputs(7808) <= (layer0_outputs(177)) and (layer0_outputs(8412));
    outputs(7809) <= layer0_outputs(5930);
    outputs(7810) <= (layer0_outputs(7897)) and not (layer0_outputs(12056));
    outputs(7811) <= not((layer0_outputs(1866)) and (layer0_outputs(2935)));
    outputs(7812) <= not(layer0_outputs(6604));
    outputs(7813) <= not(layer0_outputs(1050)) or (layer0_outputs(3109));
    outputs(7814) <= not(layer0_outputs(230));
    outputs(7815) <= not(layer0_outputs(3576));
    outputs(7816) <= layer0_outputs(11577);
    outputs(7817) <= (layer0_outputs(4990)) and (layer0_outputs(10390));
    outputs(7818) <= '0';
    outputs(7819) <= not(layer0_outputs(2369));
    outputs(7820) <= layer0_outputs(11650);
    outputs(7821) <= layer0_outputs(10888);
    outputs(7822) <= layer0_outputs(8230);
    outputs(7823) <= layer0_outputs(12138);
    outputs(7824) <= (layer0_outputs(4287)) and (layer0_outputs(12168));
    outputs(7825) <= layer0_outputs(8413);
    outputs(7826) <= not(layer0_outputs(12187)) or (layer0_outputs(9959));
    outputs(7827) <= not(layer0_outputs(10254));
    outputs(7828) <= not((layer0_outputs(71)) or (layer0_outputs(608)));
    outputs(7829) <= (layer0_outputs(7531)) and not (layer0_outputs(11073));
    outputs(7830) <= (layer0_outputs(10742)) xor (layer0_outputs(1522));
    outputs(7831) <= (layer0_outputs(11461)) and not (layer0_outputs(9956));
    outputs(7832) <= not(layer0_outputs(266));
    outputs(7833) <= (layer0_outputs(5616)) and not (layer0_outputs(2268));
    outputs(7834) <= (layer0_outputs(2855)) xor (layer0_outputs(1981));
    outputs(7835) <= (layer0_outputs(4195)) and (layer0_outputs(10240));
    outputs(7836) <= layer0_outputs(12639);
    outputs(7837) <= layer0_outputs(7429);
    outputs(7838) <= (layer0_outputs(3981)) xor (layer0_outputs(467));
    outputs(7839) <= (layer0_outputs(6280)) and (layer0_outputs(10492));
    outputs(7840) <= not(layer0_outputs(6272));
    outputs(7841) <= (layer0_outputs(1761)) and not (layer0_outputs(11933));
    outputs(7842) <= layer0_outputs(3781);
    outputs(7843) <= (layer0_outputs(8798)) and not (layer0_outputs(7151));
    outputs(7844) <= not((layer0_outputs(1273)) xor (layer0_outputs(8849)));
    outputs(7845) <= (layer0_outputs(5852)) and not (layer0_outputs(7247));
    outputs(7846) <= layer0_outputs(9645);
    outputs(7847) <= not(layer0_outputs(10363));
    outputs(7848) <= not(layer0_outputs(5697));
    outputs(7849) <= not(layer0_outputs(10595));
    outputs(7850) <= (layer0_outputs(10026)) and not (layer0_outputs(5752));
    outputs(7851) <= layer0_outputs(376);
    outputs(7852) <= (layer0_outputs(10877)) and not (layer0_outputs(4286));
    outputs(7853) <= layer0_outputs(7494);
    outputs(7854) <= not(layer0_outputs(4070));
    outputs(7855) <= not(layer0_outputs(3027));
    outputs(7856) <= layer0_outputs(8776);
    outputs(7857) <= not(layer0_outputs(8934));
    outputs(7858) <= not((layer0_outputs(12258)) xor (layer0_outputs(577)));
    outputs(7859) <= (layer0_outputs(2665)) xor (layer0_outputs(2847));
    outputs(7860) <= not(layer0_outputs(10537));
    outputs(7861) <= not(layer0_outputs(1147));
    outputs(7862) <= layer0_outputs(1727);
    outputs(7863) <= not(layer0_outputs(6202));
    outputs(7864) <= (layer0_outputs(5768)) and not (layer0_outputs(3238));
    outputs(7865) <= (layer0_outputs(6771)) xor (layer0_outputs(9151));
    outputs(7866) <= layer0_outputs(838);
    outputs(7867) <= (layer0_outputs(4813)) and not (layer0_outputs(10561));
    outputs(7868) <= not(layer0_outputs(4724));
    outputs(7869) <= (layer0_outputs(9446)) xor (layer0_outputs(9060));
    outputs(7870) <= not((layer0_outputs(5229)) xor (layer0_outputs(1726)));
    outputs(7871) <= layer0_outputs(712);
    outputs(7872) <= not(layer0_outputs(8997));
    outputs(7873) <= layer0_outputs(6029);
    outputs(7874) <= layer0_outputs(10963);
    outputs(7875) <= (layer0_outputs(4438)) and not (layer0_outputs(7687));
    outputs(7876) <= not(layer0_outputs(2501));
    outputs(7877) <= not(layer0_outputs(4177)) or (layer0_outputs(2194));
    outputs(7878) <= layer0_outputs(7299);
    outputs(7879) <= layer0_outputs(1211);
    outputs(7880) <= (layer0_outputs(2860)) xor (layer0_outputs(10862));
    outputs(7881) <= layer0_outputs(7064);
    outputs(7882) <= layer0_outputs(7804);
    outputs(7883) <= not(layer0_outputs(5469));
    outputs(7884) <= (layer0_outputs(5333)) and not (layer0_outputs(3285));
    outputs(7885) <= layer0_outputs(11560);
    outputs(7886) <= (layer0_outputs(1069)) and (layer0_outputs(11096));
    outputs(7887) <= not(layer0_outputs(4680));
    outputs(7888) <= (layer0_outputs(6603)) and not (layer0_outputs(7278));
    outputs(7889) <= (layer0_outputs(8658)) and not (layer0_outputs(1627));
    outputs(7890) <= not(layer0_outputs(10140));
    outputs(7891) <= not(layer0_outputs(758));
    outputs(7892) <= not(layer0_outputs(9214));
    outputs(7893) <= not(layer0_outputs(2684));
    outputs(7894) <= not(layer0_outputs(549)) or (layer0_outputs(7276));
    outputs(7895) <= (layer0_outputs(7889)) or (layer0_outputs(382));
    outputs(7896) <= not(layer0_outputs(8575));
    outputs(7897) <= layer0_outputs(3904);
    outputs(7898) <= (layer0_outputs(5732)) and not (layer0_outputs(4315));
    outputs(7899) <= not(layer0_outputs(5495));
    outputs(7900) <= layer0_outputs(11806);
    outputs(7901) <= not((layer0_outputs(4136)) xor (layer0_outputs(8406)));
    outputs(7902) <= (layer0_outputs(4383)) xor (layer0_outputs(8767));
    outputs(7903) <= (layer0_outputs(5568)) xor (layer0_outputs(7652));
    outputs(7904) <= not(layer0_outputs(11956)) or (layer0_outputs(5083));
    outputs(7905) <= layer0_outputs(7185);
    outputs(7906) <= layer0_outputs(5451);
    outputs(7907) <= not(layer0_outputs(7594));
    outputs(7908) <= layer0_outputs(5856);
    outputs(7909) <= (layer0_outputs(579)) xor (layer0_outputs(7058));
    outputs(7910) <= not(layer0_outputs(8575));
    outputs(7911) <= not(layer0_outputs(12478));
    outputs(7912) <= (layer0_outputs(7301)) xor (layer0_outputs(10327));
    outputs(7913) <= layer0_outputs(6005);
    outputs(7914) <= (layer0_outputs(11932)) xor (layer0_outputs(10977));
    outputs(7915) <= not(layer0_outputs(4847));
    outputs(7916) <= not((layer0_outputs(1894)) xor (layer0_outputs(10002)));
    outputs(7917) <= not(layer0_outputs(12594));
    outputs(7918) <= (layer0_outputs(6640)) and not (layer0_outputs(12129));
    outputs(7919) <= not((layer0_outputs(5675)) and (layer0_outputs(2974)));
    outputs(7920) <= not(layer0_outputs(5296));
    outputs(7921) <= layer0_outputs(4781);
    outputs(7922) <= (layer0_outputs(10334)) and not (layer0_outputs(8908));
    outputs(7923) <= not(layer0_outputs(194));
    outputs(7924) <= layer0_outputs(471);
    outputs(7925) <= not(layer0_outputs(11468)) or (layer0_outputs(7310));
    outputs(7926) <= not((layer0_outputs(8183)) or (layer0_outputs(1862)));
    outputs(7927) <= layer0_outputs(3729);
    outputs(7928) <= (layer0_outputs(9516)) or (layer0_outputs(7582));
    outputs(7929) <= (layer0_outputs(9830)) and (layer0_outputs(440));
    outputs(7930) <= (layer0_outputs(6923)) and (layer0_outputs(10113));
    outputs(7931) <= not((layer0_outputs(1533)) or (layer0_outputs(8599)));
    outputs(7932) <= not(layer0_outputs(5848));
    outputs(7933) <= not(layer0_outputs(3534)) or (layer0_outputs(8810));
    outputs(7934) <= layer0_outputs(2337);
    outputs(7935) <= (layer0_outputs(11897)) and (layer0_outputs(12211));
    outputs(7936) <= (layer0_outputs(4725)) and (layer0_outputs(6626));
    outputs(7937) <= layer0_outputs(12036);
    outputs(7938) <= not(layer0_outputs(7115));
    outputs(7939) <= layer0_outputs(5604);
    outputs(7940) <= not(layer0_outputs(1228));
    outputs(7941) <= layer0_outputs(1694);
    outputs(7942) <= layer0_outputs(5863);
    outputs(7943) <= not(layer0_outputs(11328));
    outputs(7944) <= not(layer0_outputs(1411)) or (layer0_outputs(10382));
    outputs(7945) <= (layer0_outputs(7871)) and not (layer0_outputs(7202));
    outputs(7946) <= not(layer0_outputs(11231));
    outputs(7947) <= not(layer0_outputs(8848));
    outputs(7948) <= not(layer0_outputs(7888)) or (layer0_outputs(878));
    outputs(7949) <= (layer0_outputs(11576)) or (layer0_outputs(8328));
    outputs(7950) <= not(layer0_outputs(9651));
    outputs(7951) <= layer0_outputs(4574);
    outputs(7952) <= not((layer0_outputs(4861)) or (layer0_outputs(12262)));
    outputs(7953) <= (layer0_outputs(11840)) or (layer0_outputs(997));
    outputs(7954) <= not(layer0_outputs(4491));
    outputs(7955) <= not(layer0_outputs(11748));
    outputs(7956) <= not((layer0_outputs(10142)) xor (layer0_outputs(11373)));
    outputs(7957) <= layer0_outputs(5300);
    outputs(7958) <= not(layer0_outputs(4293));
    outputs(7959) <= (layer0_outputs(6485)) xor (layer0_outputs(9053));
    outputs(7960) <= not((layer0_outputs(9605)) xor (layer0_outputs(3270)));
    outputs(7961) <= layer0_outputs(3172);
    outputs(7962) <= not((layer0_outputs(3294)) or (layer0_outputs(2573)));
    outputs(7963) <= layer0_outputs(3200);
    outputs(7964) <= (layer0_outputs(5661)) and (layer0_outputs(10048));
    outputs(7965) <= layer0_outputs(2606);
    outputs(7966) <= not(layer0_outputs(7611));
    outputs(7967) <= (layer0_outputs(12118)) and (layer0_outputs(3989));
    outputs(7968) <= (layer0_outputs(850)) and not (layer0_outputs(6768));
    outputs(7969) <= layer0_outputs(4401);
    outputs(7970) <= not(layer0_outputs(2157)) or (layer0_outputs(9122));
    outputs(7971) <= (layer0_outputs(1242)) and not (layer0_outputs(7749));
    outputs(7972) <= layer0_outputs(5088);
    outputs(7973) <= (layer0_outputs(5170)) and (layer0_outputs(4011));
    outputs(7974) <= (layer0_outputs(2681)) xor (layer0_outputs(1180));
    outputs(7975) <= not(layer0_outputs(4697));
    outputs(7976) <= (layer0_outputs(2889)) and (layer0_outputs(3382));
    outputs(7977) <= not((layer0_outputs(9532)) xor (layer0_outputs(1227)));
    outputs(7978) <= layer0_outputs(6546);
    outputs(7979) <= (layer0_outputs(11200)) and not (layer0_outputs(2391));
    outputs(7980) <= not(layer0_outputs(8193)) or (layer0_outputs(9925));
    outputs(7981) <= not(layer0_outputs(10078));
    outputs(7982) <= not(layer0_outputs(8299));
    outputs(7983) <= not(layer0_outputs(1757));
    outputs(7984) <= (layer0_outputs(10456)) or (layer0_outputs(6552));
    outputs(7985) <= not(layer0_outputs(3743));
    outputs(7986) <= not(layer0_outputs(1147)) or (layer0_outputs(9805));
    outputs(7987) <= not(layer0_outputs(3813));
    outputs(7988) <= layer0_outputs(11642);
    outputs(7989) <= layer0_outputs(6332);
    outputs(7990) <= layer0_outputs(3856);
    outputs(7991) <= layer0_outputs(898);
    outputs(7992) <= (layer0_outputs(12213)) and not (layer0_outputs(994));
    outputs(7993) <= not((layer0_outputs(2487)) or (layer0_outputs(2302)));
    outputs(7994) <= not(layer0_outputs(8663));
    outputs(7995) <= (layer0_outputs(10019)) and (layer0_outputs(9931));
    outputs(7996) <= not(layer0_outputs(11072));
    outputs(7997) <= layer0_outputs(4253);
    outputs(7998) <= layer0_outputs(7465);
    outputs(7999) <= layer0_outputs(3583);
    outputs(8000) <= (layer0_outputs(502)) and not (layer0_outputs(2452));
    outputs(8001) <= (layer0_outputs(6189)) and not (layer0_outputs(12724));
    outputs(8002) <= not((layer0_outputs(6799)) and (layer0_outputs(3930)));
    outputs(8003) <= not((layer0_outputs(3299)) xor (layer0_outputs(1516)));
    outputs(8004) <= not(layer0_outputs(7770));
    outputs(8005) <= layer0_outputs(9314);
    outputs(8006) <= (layer0_outputs(2261)) and not (layer0_outputs(7470));
    outputs(8007) <= (layer0_outputs(9692)) xor (layer0_outputs(2732));
    outputs(8008) <= not(layer0_outputs(540)) or (layer0_outputs(4996));
    outputs(8009) <= layer0_outputs(8374);
    outputs(8010) <= (layer0_outputs(12331)) xor (layer0_outputs(11238));
    outputs(8011) <= not(layer0_outputs(9897));
    outputs(8012) <= not(layer0_outputs(5303));
    outputs(8013) <= not(layer0_outputs(8309));
    outputs(8014) <= layer0_outputs(6078);
    outputs(8015) <= not(layer0_outputs(6853));
    outputs(8016) <= (layer0_outputs(9251)) xor (layer0_outputs(7533));
    outputs(8017) <= (layer0_outputs(10137)) and not (layer0_outputs(10416));
    outputs(8018) <= (layer0_outputs(3158)) and not (layer0_outputs(10687));
    outputs(8019) <= layer0_outputs(4579);
    outputs(8020) <= not(layer0_outputs(6104));
    outputs(8021) <= layer0_outputs(4309);
    outputs(8022) <= layer0_outputs(284);
    outputs(8023) <= layer0_outputs(8864);
    outputs(8024) <= not(layer0_outputs(3691));
    outputs(8025) <= '0';
    outputs(8026) <= layer0_outputs(10446);
    outputs(8027) <= layer0_outputs(5308);
    outputs(8028) <= not(layer0_outputs(5224));
    outputs(8029) <= (layer0_outputs(12656)) or (layer0_outputs(2209));
    outputs(8030) <= not((layer0_outputs(5563)) or (layer0_outputs(4680)));
    outputs(8031) <= not(layer0_outputs(6326));
    outputs(8032) <= (layer0_outputs(5887)) and (layer0_outputs(9884));
    outputs(8033) <= not(layer0_outputs(3082)) or (layer0_outputs(6591));
    outputs(8034) <= not(layer0_outputs(2710));
    outputs(8035) <= (layer0_outputs(11742)) or (layer0_outputs(8787));
    outputs(8036) <= not(layer0_outputs(11831));
    outputs(8037) <= not(layer0_outputs(6433));
    outputs(8038) <= layer0_outputs(12648);
    outputs(8039) <= not(layer0_outputs(4391));
    outputs(8040) <= not((layer0_outputs(7506)) and (layer0_outputs(4093)));
    outputs(8041) <= layer0_outputs(9207);
    outputs(8042) <= layer0_outputs(3788);
    outputs(8043) <= not((layer0_outputs(11792)) xor (layer0_outputs(8069)));
    outputs(8044) <= (layer0_outputs(1086)) and (layer0_outputs(8014));
    outputs(8045) <= layer0_outputs(4269);
    outputs(8046) <= (layer0_outputs(7245)) xor (layer0_outputs(11418));
    outputs(8047) <= not(layer0_outputs(1156));
    outputs(8048) <= (layer0_outputs(3956)) or (layer0_outputs(5426));
    outputs(8049) <= (layer0_outputs(10251)) xor (layer0_outputs(6963));
    outputs(8050) <= (layer0_outputs(5674)) and (layer0_outputs(1297));
    outputs(8051) <= not(layer0_outputs(687));
    outputs(8052) <= layer0_outputs(2567);
    outputs(8053) <= layer0_outputs(2571);
    outputs(8054) <= layer0_outputs(8159);
    outputs(8055) <= not(layer0_outputs(8110)) or (layer0_outputs(5468));
    outputs(8056) <= (layer0_outputs(2937)) and not (layer0_outputs(7544));
    outputs(8057) <= (layer0_outputs(8680)) xor (layer0_outputs(6448));
    outputs(8058) <= not(layer0_outputs(1129));
    outputs(8059) <= layer0_outputs(4837);
    outputs(8060) <= (layer0_outputs(9754)) or (layer0_outputs(8352));
    outputs(8061) <= not(layer0_outputs(6393));
    outputs(8062) <= layer0_outputs(3087);
    outputs(8063) <= layer0_outputs(5714);
    outputs(8064) <= not(layer0_outputs(9073));
    outputs(8065) <= not(layer0_outputs(12741));
    outputs(8066) <= not((layer0_outputs(9336)) xor (layer0_outputs(9119)));
    outputs(8067) <= (layer0_outputs(9615)) or (layer0_outputs(931));
    outputs(8068) <= not((layer0_outputs(10371)) xor (layer0_outputs(374)));
    outputs(8069) <= (layer0_outputs(6666)) and not (layer0_outputs(8818));
    outputs(8070) <= (layer0_outputs(6373)) xor (layer0_outputs(801));
    outputs(8071) <= not((layer0_outputs(1260)) xor (layer0_outputs(8941)));
    outputs(8072) <= not(layer0_outputs(7406));
    outputs(8073) <= (layer0_outputs(7223)) and not (layer0_outputs(8872));
    outputs(8074) <= (layer0_outputs(1880)) xor (layer0_outputs(10996));
    outputs(8075) <= not((layer0_outputs(11837)) xor (layer0_outputs(8438)));
    outputs(8076) <= not(layer0_outputs(7900));
    outputs(8077) <= layer0_outputs(10793);
    outputs(8078) <= not((layer0_outputs(7461)) xor (layer0_outputs(6049)));
    outputs(8079) <= not(layer0_outputs(6795));
    outputs(8080) <= not(layer0_outputs(11316));
    outputs(8081) <= not(layer0_outputs(9111));
    outputs(8082) <= not(layer0_outputs(2328));
    outputs(8083) <= (layer0_outputs(3197)) and not (layer0_outputs(869));
    outputs(8084) <= layer0_outputs(8613);
    outputs(8085) <= layer0_outputs(3901);
    outputs(8086) <= not(layer0_outputs(5325));
    outputs(8087) <= not(layer0_outputs(8012));
    outputs(8088) <= (layer0_outputs(553)) and not (layer0_outputs(7416));
    outputs(8089) <= not((layer0_outputs(2499)) or (layer0_outputs(5292)));
    outputs(8090) <= (layer0_outputs(10928)) and not (layer0_outputs(2555));
    outputs(8091) <= layer0_outputs(4199);
    outputs(8092) <= not(layer0_outputs(12580));
    outputs(8093) <= layer0_outputs(1890);
    outputs(8094) <= layer0_outputs(8975);
    outputs(8095) <= not(layer0_outputs(2640));
    outputs(8096) <= not(layer0_outputs(1973));
    outputs(8097) <= not(layer0_outputs(4754));
    outputs(8098) <= not(layer0_outputs(607));
    outputs(8099) <= not(layer0_outputs(4622)) or (layer0_outputs(9048));
    outputs(8100) <= not(layer0_outputs(6291));
    outputs(8101) <= layer0_outputs(8447);
    outputs(8102) <= layer0_outputs(1545);
    outputs(8103) <= layer0_outputs(4777);
    outputs(8104) <= layer0_outputs(470);
    outputs(8105) <= (layer0_outputs(4262)) and not (layer0_outputs(1566));
    outputs(8106) <= layer0_outputs(12195);
    outputs(8107) <= layer0_outputs(3014);
    outputs(8108) <= (layer0_outputs(7563)) xor (layer0_outputs(6915));
    outputs(8109) <= (layer0_outputs(8222)) and (layer0_outputs(5875));
    outputs(8110) <= (layer0_outputs(9378)) and not (layer0_outputs(4041));
    outputs(8111) <= not(layer0_outputs(6708));
    outputs(8112) <= layer0_outputs(6304);
    outputs(8113) <= not(layer0_outputs(8796));
    outputs(8114) <= not((layer0_outputs(2089)) xor (layer0_outputs(3133)));
    outputs(8115) <= layer0_outputs(7614);
    outputs(8116) <= not(layer0_outputs(10224));
    outputs(8117) <= layer0_outputs(1451);
    outputs(8118) <= layer0_outputs(9772);
    outputs(8119) <= layer0_outputs(11487);
    outputs(8120) <= not(layer0_outputs(6844));
    outputs(8121) <= not(layer0_outputs(456));
    outputs(8122) <= layer0_outputs(11633);
    outputs(8123) <= layer0_outputs(7286);
    outputs(8124) <= (layer0_outputs(5721)) and not (layer0_outputs(8599));
    outputs(8125) <= layer0_outputs(1163);
    outputs(8126) <= (layer0_outputs(7719)) xor (layer0_outputs(2748));
    outputs(8127) <= layer0_outputs(6240);
    outputs(8128) <= not((layer0_outputs(5189)) xor (layer0_outputs(2469)));
    outputs(8129) <= layer0_outputs(169);
    outputs(8130) <= not((layer0_outputs(7963)) and (layer0_outputs(5151)));
    outputs(8131) <= not(layer0_outputs(2510)) or (layer0_outputs(3807));
    outputs(8132) <= not(layer0_outputs(10988));
    outputs(8133) <= layer0_outputs(2567);
    outputs(8134) <= not(layer0_outputs(5541));
    outputs(8135) <= (layer0_outputs(10287)) and not (layer0_outputs(1951));
    outputs(8136) <= (layer0_outputs(8159)) and not (layer0_outputs(2459));
    outputs(8137) <= layer0_outputs(5838);
    outputs(8138) <= not(layer0_outputs(7752));
    outputs(8139) <= not(layer0_outputs(6282));
    outputs(8140) <= not(layer0_outputs(745));
    outputs(8141) <= not(layer0_outputs(12534)) or (layer0_outputs(8093));
    outputs(8142) <= not(layer0_outputs(9939));
    outputs(8143) <= not(layer0_outputs(9234));
    outputs(8144) <= (layer0_outputs(2356)) and not (layer0_outputs(1146));
    outputs(8145) <= not(layer0_outputs(6109)) or (layer0_outputs(4153));
    outputs(8146) <= layer0_outputs(3971);
    outputs(8147) <= not((layer0_outputs(1077)) or (layer0_outputs(5416)));
    outputs(8148) <= layer0_outputs(6916);
    outputs(8149) <= not((layer0_outputs(3278)) xor (layer0_outputs(10690)));
    outputs(8150) <= not(layer0_outputs(6614));
    outputs(8151) <= layer0_outputs(7385);
    outputs(8152) <= (layer0_outputs(213)) or (layer0_outputs(2267));
    outputs(8153) <= layer0_outputs(10415);
    outputs(8154) <= not(layer0_outputs(7383));
    outputs(8155) <= not(layer0_outputs(8175));
    outputs(8156) <= not((layer0_outputs(115)) or (layer0_outputs(5126)));
    outputs(8157) <= not(layer0_outputs(419));
    outputs(8158) <= layer0_outputs(4988);
    outputs(8159) <= not(layer0_outputs(3911));
    outputs(8160) <= (layer0_outputs(10984)) and (layer0_outputs(3906));
    outputs(8161) <= not(layer0_outputs(6335));
    outputs(8162) <= layer0_outputs(4356);
    outputs(8163) <= layer0_outputs(9576);
    outputs(8164) <= not((layer0_outputs(7325)) xor (layer0_outputs(9648)));
    outputs(8165) <= not((layer0_outputs(9465)) xor (layer0_outputs(10975)));
    outputs(8166) <= layer0_outputs(11157);
    outputs(8167) <= (layer0_outputs(584)) and not (layer0_outputs(8896));
    outputs(8168) <= not(layer0_outputs(11015));
    outputs(8169) <= layer0_outputs(2808);
    outputs(8170) <= not(layer0_outputs(4051));
    outputs(8171) <= not(layer0_outputs(1208));
    outputs(8172) <= layer0_outputs(10838);
    outputs(8173) <= (layer0_outputs(1432)) and not (layer0_outputs(11620));
    outputs(8174) <= not((layer0_outputs(7819)) xor (layer0_outputs(5259)));
    outputs(8175) <= not(layer0_outputs(792));
    outputs(8176) <= layer0_outputs(7685);
    outputs(8177) <= (layer0_outputs(12358)) or (layer0_outputs(9751));
    outputs(8178) <= not(layer0_outputs(12100));
    outputs(8179) <= layer0_outputs(10233);
    outputs(8180) <= layer0_outputs(4726);
    outputs(8181) <= not((layer0_outputs(5567)) xor (layer0_outputs(411)));
    outputs(8182) <= (layer0_outputs(9546)) and (layer0_outputs(5706));
    outputs(8183) <= not((layer0_outputs(9011)) and (layer0_outputs(151)));
    outputs(8184) <= not(layer0_outputs(8016));
    outputs(8185) <= not(layer0_outputs(2385));
    outputs(8186) <= not(layer0_outputs(3692));
    outputs(8187) <= not(layer0_outputs(10813));
    outputs(8188) <= (layer0_outputs(10601)) and not (layer0_outputs(8828));
    outputs(8189) <= not(layer0_outputs(1904));
    outputs(8190) <= layer0_outputs(10807);
    outputs(8191) <= not(layer0_outputs(11481));
    outputs(8192) <= layer0_outputs(3048);
    outputs(8193) <= (layer0_outputs(12420)) and not (layer0_outputs(2544));
    outputs(8194) <= (layer0_outputs(348)) xor (layer0_outputs(7217));
    outputs(8195) <= not(layer0_outputs(5830));
    outputs(8196) <= not(layer0_outputs(9380));
    outputs(8197) <= not(layer0_outputs(11533));
    outputs(8198) <= not(layer0_outputs(4278));
    outputs(8199) <= (layer0_outputs(3752)) and not (layer0_outputs(1403));
    outputs(8200) <= layer0_outputs(8929);
    outputs(8201) <= layer0_outputs(4347);
    outputs(8202) <= (layer0_outputs(1485)) and not (layer0_outputs(10315));
    outputs(8203) <= layer0_outputs(2802);
    outputs(8204) <= not(layer0_outputs(5869));
    outputs(8205) <= (layer0_outputs(3512)) or (layer0_outputs(6727));
    outputs(8206) <= not(layer0_outputs(9791));
    outputs(8207) <= layer0_outputs(3428);
    outputs(8208) <= (layer0_outputs(865)) and not (layer0_outputs(1675));
    outputs(8209) <= layer0_outputs(10639);
    outputs(8210) <= layer0_outputs(5031);
    outputs(8211) <= layer0_outputs(6091);
    outputs(8212) <= layer0_outputs(8414);
    outputs(8213) <= layer0_outputs(10691);
    outputs(8214) <= (layer0_outputs(4296)) xor (layer0_outputs(1580));
    outputs(8215) <= (layer0_outputs(7263)) or (layer0_outputs(5308));
    outputs(8216) <= not((layer0_outputs(3898)) xor (layer0_outputs(143)));
    outputs(8217) <= not(layer0_outputs(4429));
    outputs(8218) <= not(layer0_outputs(4207));
    outputs(8219) <= layer0_outputs(10672);
    outputs(8220) <= layer0_outputs(7604);
    outputs(8221) <= not(layer0_outputs(67));
    outputs(8222) <= not(layer0_outputs(6299));
    outputs(8223) <= not(layer0_outputs(706));
    outputs(8224) <= not(layer0_outputs(6833));
    outputs(8225) <= not(layer0_outputs(9901));
    outputs(8226) <= (layer0_outputs(1787)) and not (layer0_outputs(11574));
    outputs(8227) <= layer0_outputs(1653);
    outputs(8228) <= not(layer0_outputs(1693));
    outputs(8229) <= layer0_outputs(12517);
    outputs(8230) <= not((layer0_outputs(8057)) xor (layer0_outputs(6859)));
    outputs(8231) <= not(layer0_outputs(7179));
    outputs(8232) <= not((layer0_outputs(7886)) xor (layer0_outputs(2427)));
    outputs(8233) <= (layer0_outputs(1086)) and (layer0_outputs(8629));
    outputs(8234) <= not(layer0_outputs(1102)) or (layer0_outputs(4271));
    outputs(8235) <= (layer0_outputs(10191)) or (layer0_outputs(12379));
    outputs(8236) <= layer0_outputs(5504);
    outputs(8237) <= not((layer0_outputs(1296)) xor (layer0_outputs(2831)));
    outputs(8238) <= layer0_outputs(10954);
    outputs(8239) <= not(layer0_outputs(9407));
    outputs(8240) <= layer0_outputs(7037);
    outputs(8241) <= (layer0_outputs(1671)) and not (layer0_outputs(6930));
    outputs(8242) <= layer0_outputs(12139);
    outputs(8243) <= (layer0_outputs(9093)) xor (layer0_outputs(10252));
    outputs(8244) <= (layer0_outputs(2078)) and not (layer0_outputs(606));
    outputs(8245) <= not(layer0_outputs(10393));
    outputs(8246) <= (layer0_outputs(8824)) and not (layer0_outputs(11997));
    outputs(8247) <= layer0_outputs(576);
    outputs(8248) <= not((layer0_outputs(9606)) and (layer0_outputs(8906)));
    outputs(8249) <= layer0_outputs(179);
    outputs(8250) <= (layer0_outputs(11727)) xor (layer0_outputs(1956));
    outputs(8251) <= not((layer0_outputs(3909)) xor (layer0_outputs(3258)));
    outputs(8252) <= (layer0_outputs(6223)) and not (layer0_outputs(8422));
    outputs(8253) <= (layer0_outputs(11630)) and not (layer0_outputs(5370));
    outputs(8254) <= (layer0_outputs(7039)) and not (layer0_outputs(494));
    outputs(8255) <= not(layer0_outputs(10491));
    outputs(8256) <= not(layer0_outputs(2300));
    outputs(8257) <= not(layer0_outputs(2982));
    outputs(8258) <= not(layer0_outputs(10249));
    outputs(8259) <= not((layer0_outputs(240)) xor (layer0_outputs(8889)));
    outputs(8260) <= not((layer0_outputs(9486)) or (layer0_outputs(6060)));
    outputs(8261) <= not((layer0_outputs(562)) or (layer0_outputs(1185)));
    outputs(8262) <= not((layer0_outputs(1190)) xor (layer0_outputs(12719)));
    outputs(8263) <= layer0_outputs(11293);
    outputs(8264) <= not(layer0_outputs(7723));
    outputs(8265) <= (layer0_outputs(8147)) and not (layer0_outputs(2345));
    outputs(8266) <= (layer0_outputs(8120)) xor (layer0_outputs(5534));
    outputs(8267) <= not(layer0_outputs(3848));
    outputs(8268) <= layer0_outputs(8435);
    outputs(8269) <= not(layer0_outputs(7377));
    outputs(8270) <= layer0_outputs(5380);
    outputs(8271) <= not(layer0_outputs(7939));
    outputs(8272) <= not(layer0_outputs(12252)) or (layer0_outputs(9059));
    outputs(8273) <= layer0_outputs(11623);
    outputs(8274) <= not((layer0_outputs(4146)) xor (layer0_outputs(1336)));
    outputs(8275) <= (layer0_outputs(1864)) xor (layer0_outputs(1353));
    outputs(8276) <= not(layer0_outputs(10547));
    outputs(8277) <= layer0_outputs(12446);
    outputs(8278) <= (layer0_outputs(9420)) xor (layer0_outputs(8503));
    outputs(8279) <= layer0_outputs(8255);
    outputs(8280) <= not(layer0_outputs(12798));
    outputs(8281) <= not(layer0_outputs(2704));
    outputs(8282) <= not((layer0_outputs(2074)) xor (layer0_outputs(12669)));
    outputs(8283) <= layer0_outputs(8466);
    outputs(8284) <= (layer0_outputs(10872)) xor (layer0_outputs(626));
    outputs(8285) <= (layer0_outputs(3314)) xor (layer0_outputs(6646));
    outputs(8286) <= (layer0_outputs(11373)) xor (layer0_outputs(4557));
    outputs(8287) <= not(layer0_outputs(4564));
    outputs(8288) <= layer0_outputs(5893);
    outputs(8289) <= layer0_outputs(1038);
    outputs(8290) <= layer0_outputs(3559);
    outputs(8291) <= not((layer0_outputs(1171)) or (layer0_outputs(9150)));
    outputs(8292) <= not(layer0_outputs(7190));
    outputs(8293) <= (layer0_outputs(1983)) xor (layer0_outputs(11588));
    outputs(8294) <= layer0_outputs(2798);
    outputs(8295) <= layer0_outputs(8146);
    outputs(8296) <= layer0_outputs(9855);
    outputs(8297) <= not((layer0_outputs(10222)) xor (layer0_outputs(7825)));
    outputs(8298) <= (layer0_outputs(10427)) xor (layer0_outputs(1514));
    outputs(8299) <= (layer0_outputs(7983)) xor (layer0_outputs(1879));
    outputs(8300) <= not((layer0_outputs(7132)) xor (layer0_outputs(2071)));
    outputs(8301) <= not(layer0_outputs(6122)) or (layer0_outputs(7731));
    outputs(8302) <= not(layer0_outputs(10439));
    outputs(8303) <= not(layer0_outputs(2695));
    outputs(8304) <= not((layer0_outputs(6626)) xor (layer0_outputs(6889)));
    outputs(8305) <= (layer0_outputs(4235)) xor (layer0_outputs(3059));
    outputs(8306) <= not(layer0_outputs(1676));
    outputs(8307) <= not((layer0_outputs(9310)) xor (layer0_outputs(11402)));
    outputs(8308) <= (layer0_outputs(2517)) xor (layer0_outputs(2106));
    outputs(8309) <= layer0_outputs(8902);
    outputs(8310) <= not((layer0_outputs(12569)) xor (layer0_outputs(868)));
    outputs(8311) <= not(layer0_outputs(9312));
    outputs(8312) <= not(layer0_outputs(9360));
    outputs(8313) <= (layer0_outputs(3887)) and not (layer0_outputs(6254));
    outputs(8314) <= (layer0_outputs(5250)) xor (layer0_outputs(2125));
    outputs(8315) <= layer0_outputs(6214);
    outputs(8316) <= (layer0_outputs(1462)) xor (layer0_outputs(11120));
    outputs(8317) <= (layer0_outputs(4163)) xor (layer0_outputs(2253));
    outputs(8318) <= not(layer0_outputs(9967));
    outputs(8319) <= layer0_outputs(4224);
    outputs(8320) <= (layer0_outputs(35)) xor (layer0_outputs(3976));
    outputs(8321) <= (layer0_outputs(11050)) and (layer0_outputs(5229));
    outputs(8322) <= not(layer0_outputs(2084));
    outputs(8323) <= layer0_outputs(7054);
    outputs(8324) <= not(layer0_outputs(4854));
    outputs(8325) <= layer0_outputs(8654);
    outputs(8326) <= layer0_outputs(12530);
    outputs(8327) <= not((layer0_outputs(5519)) xor (layer0_outputs(1334)));
    outputs(8328) <= (layer0_outputs(11539)) and not (layer0_outputs(3972));
    outputs(8329) <= not(layer0_outputs(4801));
    outputs(8330) <= not((layer0_outputs(6022)) xor (layer0_outputs(4442)));
    outputs(8331) <= not(layer0_outputs(5808));
    outputs(8332) <= not(layer0_outputs(12586));
    outputs(8333) <= layer0_outputs(9345);
    outputs(8334) <= not((layer0_outputs(9755)) and (layer0_outputs(3550)));
    outputs(8335) <= layer0_outputs(12597);
    outputs(8336) <= not(layer0_outputs(1035)) or (layer0_outputs(5584));
    outputs(8337) <= not(layer0_outputs(2253));
    outputs(8338) <= not((layer0_outputs(4003)) and (layer0_outputs(11919)));
    outputs(8339) <= layer0_outputs(10622);
    outputs(8340) <= layer0_outputs(8702);
    outputs(8341) <= layer0_outputs(3835);
    outputs(8342) <= layer0_outputs(9489);
    outputs(8343) <= layer0_outputs(9231);
    outputs(8344) <= (layer0_outputs(3203)) and (layer0_outputs(11311));
    outputs(8345) <= layer0_outputs(254);
    outputs(8346) <= '1';
    outputs(8347) <= layer0_outputs(5817);
    outputs(8348) <= layer0_outputs(9367);
    outputs(8349) <= not(layer0_outputs(2769));
    outputs(8350) <= (layer0_outputs(890)) xor (layer0_outputs(3405));
    outputs(8351) <= not(layer0_outputs(3392));
    outputs(8352) <= not(layer0_outputs(6708)) or (layer0_outputs(2574));
    outputs(8353) <= layer0_outputs(6196);
    outputs(8354) <= not(layer0_outputs(8550));
    outputs(8355) <= not(layer0_outputs(6977));
    outputs(8356) <= (layer0_outputs(10896)) and (layer0_outputs(137));
    outputs(8357) <= layer0_outputs(6475);
    outputs(8358) <= (layer0_outputs(4527)) xor (layer0_outputs(5942));
    outputs(8359) <= layer0_outputs(10884);
    outputs(8360) <= (layer0_outputs(12682)) and not (layer0_outputs(10419));
    outputs(8361) <= layer0_outputs(11096);
    outputs(8362) <= not(layer0_outputs(4109)) or (layer0_outputs(6366));
    outputs(8363) <= not((layer0_outputs(202)) xor (layer0_outputs(2390)));
    outputs(8364) <= layer0_outputs(1753);
    outputs(8365) <= not(layer0_outputs(10993)) or (layer0_outputs(6416));
    outputs(8366) <= not((layer0_outputs(3788)) xor (layer0_outputs(6992)));
    outputs(8367) <= not(layer0_outputs(4248));
    outputs(8368) <= (layer0_outputs(9752)) and (layer0_outputs(7451));
    outputs(8369) <= layer0_outputs(10575);
    outputs(8370) <= not(layer0_outputs(3942)) or (layer0_outputs(1041));
    outputs(8371) <= not((layer0_outputs(649)) or (layer0_outputs(5896)));
    outputs(8372) <= not(layer0_outputs(4198));
    outputs(8373) <= not(layer0_outputs(1521));
    outputs(8374) <= (layer0_outputs(10109)) and not (layer0_outputs(9817));
    outputs(8375) <= layer0_outputs(11030);
    outputs(8376) <= layer0_outputs(12242);
    outputs(8377) <= not(layer0_outputs(12523));
    outputs(8378) <= not((layer0_outputs(843)) or (layer0_outputs(3575)));
    outputs(8379) <= not(layer0_outputs(1183));
    outputs(8380) <= layer0_outputs(5930);
    outputs(8381) <= not((layer0_outputs(2400)) or (layer0_outputs(3122)));
    outputs(8382) <= not(layer0_outputs(9235));
    outputs(8383) <= (layer0_outputs(4856)) and not (layer0_outputs(451));
    outputs(8384) <= not((layer0_outputs(9094)) xor (layer0_outputs(3962)));
    outputs(8385) <= not(layer0_outputs(11295));
    outputs(8386) <= (layer0_outputs(72)) and (layer0_outputs(2149));
    outputs(8387) <= not(layer0_outputs(2828));
    outputs(8388) <= not(layer0_outputs(6315));
    outputs(8389) <= layer0_outputs(8703);
    outputs(8390) <= (layer0_outputs(10903)) and not (layer0_outputs(786));
    outputs(8391) <= not(layer0_outputs(1745));
    outputs(8392) <= (layer0_outputs(6867)) and not (layer0_outputs(10924));
    outputs(8393) <= layer0_outputs(7083);
    outputs(8394) <= layer0_outputs(8739);
    outputs(8395) <= not((layer0_outputs(7323)) xor (layer0_outputs(11369)));
    outputs(8396) <= not(layer0_outputs(2387));
    outputs(8397) <= layer0_outputs(7220);
    outputs(8398) <= (layer0_outputs(6365)) or (layer0_outputs(2881));
    outputs(8399) <= not(layer0_outputs(2030));
    outputs(8400) <= not(layer0_outputs(5518));
    outputs(8401) <= not(layer0_outputs(76));
    outputs(8402) <= not(layer0_outputs(3928));
    outputs(8403) <= not(layer0_outputs(8174));
    outputs(8404) <= layer0_outputs(3134);
    outputs(8405) <= layer0_outputs(8974);
    outputs(8406) <= layer0_outputs(5596);
    outputs(8407) <= not(layer0_outputs(2512)) or (layer0_outputs(794));
    outputs(8408) <= layer0_outputs(3231);
    outputs(8409) <= layer0_outputs(5059);
    outputs(8410) <= not(layer0_outputs(11922)) or (layer0_outputs(10709));
    outputs(8411) <= not((layer0_outputs(4659)) xor (layer0_outputs(7921)));
    outputs(8412) <= not(layer0_outputs(9095));
    outputs(8413) <= layer0_outputs(5444);
    outputs(8414) <= not(layer0_outputs(10946));
    outputs(8415) <= layer0_outputs(3120);
    outputs(8416) <= not((layer0_outputs(5827)) xor (layer0_outputs(5314)));
    outputs(8417) <= layer0_outputs(8485);
    outputs(8418) <= (layer0_outputs(5738)) xor (layer0_outputs(11254));
    outputs(8419) <= layer0_outputs(6039);
    outputs(8420) <= not(layer0_outputs(6930));
    outputs(8421) <= not(layer0_outputs(10773));
    outputs(8422) <= not(layer0_outputs(384));
    outputs(8423) <= not(layer0_outputs(10645)) or (layer0_outputs(4848));
    outputs(8424) <= not(layer0_outputs(7096));
    outputs(8425) <= (layer0_outputs(4640)) and not (layer0_outputs(851));
    outputs(8426) <= not(layer0_outputs(8499));
    outputs(8427) <= layer0_outputs(4253);
    outputs(8428) <= layer0_outputs(5813);
    outputs(8429) <= (layer0_outputs(6938)) or (layer0_outputs(12206));
    outputs(8430) <= layer0_outputs(9781);
    outputs(8431) <= layer0_outputs(4013);
    outputs(8432) <= not(layer0_outputs(12320));
    outputs(8433) <= not(layer0_outputs(4418));
    outputs(8434) <= not(layer0_outputs(6684)) or (layer0_outputs(1576));
    outputs(8435) <= not(layer0_outputs(10163));
    outputs(8436) <= layer0_outputs(2134);
    outputs(8437) <= not(layer0_outputs(9764));
    outputs(8438) <= not(layer0_outputs(12537));
    outputs(8439) <= (layer0_outputs(5408)) and not (layer0_outputs(6707));
    outputs(8440) <= (layer0_outputs(10405)) or (layer0_outputs(7364));
    outputs(8441) <= not(layer0_outputs(8541));
    outputs(8442) <= (layer0_outputs(9191)) and not (layer0_outputs(9348));
    outputs(8443) <= not(layer0_outputs(1650)) or (layer0_outputs(2228));
    outputs(8444) <= not((layer0_outputs(8695)) xor (layer0_outputs(2287)));
    outputs(8445) <= not((layer0_outputs(12514)) and (layer0_outputs(3918)));
    outputs(8446) <= layer0_outputs(7243);
    outputs(8447) <= not(layer0_outputs(2863));
    outputs(8448) <= not(layer0_outputs(4066));
    outputs(8449) <= layer0_outputs(3340);
    outputs(8450) <= (layer0_outputs(10827)) and (layer0_outputs(9571));
    outputs(8451) <= layer0_outputs(2719);
    outputs(8452) <= not(layer0_outputs(6235));
    outputs(8453) <= layer0_outputs(4258);
    outputs(8454) <= not(layer0_outputs(6620));
    outputs(8455) <= (layer0_outputs(484)) or (layer0_outputs(11322));
    outputs(8456) <= (layer0_outputs(9889)) or (layer0_outputs(4541));
    outputs(8457) <= layer0_outputs(8130);
    outputs(8458) <= not(layer0_outputs(428));
    outputs(8459) <= (layer0_outputs(4090)) or (layer0_outputs(11009));
    outputs(8460) <= not(layer0_outputs(2658));
    outputs(8461) <= layer0_outputs(11514);
    outputs(8462) <= not(layer0_outputs(4691));
    outputs(8463) <= layer0_outputs(10517);
    outputs(8464) <= not(layer0_outputs(5476));
    outputs(8465) <= (layer0_outputs(9884)) and (layer0_outputs(4705));
    outputs(8466) <= not(layer0_outputs(9708));
    outputs(8467) <= not(layer0_outputs(11570));
    outputs(8468) <= layer0_outputs(1698);
    outputs(8469) <= (layer0_outputs(8212)) and not (layer0_outputs(8440));
    outputs(8470) <= (layer0_outputs(7349)) or (layer0_outputs(5397));
    outputs(8471) <= not(layer0_outputs(1771));
    outputs(8472) <= (layer0_outputs(10876)) or (layer0_outputs(3816));
    outputs(8473) <= not(layer0_outputs(12342));
    outputs(8474) <= not(layer0_outputs(12204));
    outputs(8475) <= (layer0_outputs(8604)) xor (layer0_outputs(3071));
    outputs(8476) <= not((layer0_outputs(12435)) xor (layer0_outputs(455)));
    outputs(8477) <= not(layer0_outputs(10511)) or (layer0_outputs(10362));
    outputs(8478) <= layer0_outputs(2833);
    outputs(8479) <= not(layer0_outputs(6177));
    outputs(8480) <= not(layer0_outputs(11145));
    outputs(8481) <= layer0_outputs(10001);
    outputs(8482) <= layer0_outputs(8587);
    outputs(8483) <= layer0_outputs(6239);
    outputs(8484) <= (layer0_outputs(10184)) and not (layer0_outputs(8918));
    outputs(8485) <= layer0_outputs(1401);
    outputs(8486) <= not(layer0_outputs(8446));
    outputs(8487) <= (layer0_outputs(283)) and (layer0_outputs(12712));
    outputs(8488) <= not((layer0_outputs(11898)) xor (layer0_outputs(1310)));
    outputs(8489) <= not(layer0_outputs(1586));
    outputs(8490) <= layer0_outputs(11777);
    outputs(8491) <= layer0_outputs(10214);
    outputs(8492) <= not((layer0_outputs(6876)) and (layer0_outputs(1655)));
    outputs(8493) <= not(layer0_outputs(4338));
    outputs(8494) <= (layer0_outputs(2473)) and not (layer0_outputs(11543));
    outputs(8495) <= not(layer0_outputs(11881)) or (layer0_outputs(5775));
    outputs(8496) <= (layer0_outputs(4078)) xor (layer0_outputs(1741));
    outputs(8497) <= layer0_outputs(11876);
    outputs(8498) <= not(layer0_outputs(12380));
    outputs(8499) <= not(layer0_outputs(3607));
    outputs(8500) <= not((layer0_outputs(126)) or (layer0_outputs(7754)));
    outputs(8501) <= (layer0_outputs(2160)) xor (layer0_outputs(5212));
    outputs(8502) <= not(layer0_outputs(6729));
    outputs(8503) <= not((layer0_outputs(5517)) and (layer0_outputs(536)));
    outputs(8504) <= layer0_outputs(3254);
    outputs(8505) <= not((layer0_outputs(12547)) xor (layer0_outputs(11013)));
    outputs(8506) <= (layer0_outputs(2234)) and not (layer0_outputs(1506));
    outputs(8507) <= (layer0_outputs(6178)) or (layer0_outputs(894));
    outputs(8508) <= layer0_outputs(404);
    outputs(8509) <= (layer0_outputs(2730)) xor (layer0_outputs(12481));
    outputs(8510) <= layer0_outputs(8413);
    outputs(8511) <= not(layer0_outputs(6669));
    outputs(8512) <= not(layer0_outputs(3192));
    outputs(8513) <= layer0_outputs(2739);
    outputs(8514) <= (layer0_outputs(11892)) xor (layer0_outputs(2788));
    outputs(8515) <= layer0_outputs(7707);
    outputs(8516) <= layer0_outputs(3747);
    outputs(8517) <= (layer0_outputs(8949)) and not (layer0_outputs(9248));
    outputs(8518) <= not(layer0_outputs(8106));
    outputs(8519) <= (layer0_outputs(8529)) or (layer0_outputs(3655));
    outputs(8520) <= layer0_outputs(5345);
    outputs(8521) <= not(layer0_outputs(295));
    outputs(8522) <= not(layer0_outputs(4828));
    outputs(8523) <= layer0_outputs(2117);
    outputs(8524) <= not(layer0_outputs(2068));
    outputs(8525) <= layer0_outputs(1133);
    outputs(8526) <= layer0_outputs(11241);
    outputs(8527) <= not(layer0_outputs(10221));
    outputs(8528) <= not(layer0_outputs(1306));
    outputs(8529) <= layer0_outputs(10706);
    outputs(8530) <= not(layer0_outputs(2404));
    outputs(8531) <= layer0_outputs(12034);
    outputs(8532) <= not(layer0_outputs(10394));
    outputs(8533) <= not(layer0_outputs(12068));
    outputs(8534) <= (layer0_outputs(166)) xor (layer0_outputs(8994));
    outputs(8535) <= not((layer0_outputs(11708)) and (layer0_outputs(2421)));
    outputs(8536) <= not(layer0_outputs(9663));
    outputs(8537) <= not(layer0_outputs(11110));
    outputs(8538) <= (layer0_outputs(4687)) and not (layer0_outputs(1008));
    outputs(8539) <= not((layer0_outputs(3812)) and (layer0_outputs(1579)));
    outputs(8540) <= layer0_outputs(10369);
    outputs(8541) <= (layer0_outputs(8564)) or (layer0_outputs(2638));
    outputs(8542) <= not(layer0_outputs(3860));
    outputs(8543) <= not(layer0_outputs(11998)) or (layer0_outputs(5906));
    outputs(8544) <= not((layer0_outputs(5912)) xor (layer0_outputs(7679)));
    outputs(8545) <= layer0_outputs(4775);
    outputs(8546) <= layer0_outputs(12777);
    outputs(8547) <= layer0_outputs(7552);
    outputs(8548) <= not(layer0_outputs(6516));
    outputs(8549) <= not(layer0_outputs(9055)) or (layer0_outputs(6630));
    outputs(8550) <= layer0_outputs(6778);
    outputs(8551) <= not(layer0_outputs(7080));
    outputs(8552) <= layer0_outputs(4798);
    outputs(8553) <= not(layer0_outputs(6398));
    outputs(8554) <= not(layer0_outputs(8128));
    outputs(8555) <= not(layer0_outputs(12567));
    outputs(8556) <= layer0_outputs(102);
    outputs(8557) <= not(layer0_outputs(6709));
    outputs(8558) <= not(layer0_outputs(8022));
    outputs(8559) <= not(layer0_outputs(6702));
    outputs(8560) <= '0';
    outputs(8561) <= not(layer0_outputs(12459));
    outputs(8562) <= not(layer0_outputs(7536));
    outputs(8563) <= not(layer0_outputs(10254));
    outputs(8564) <= not(layer0_outputs(12370));
    outputs(8565) <= (layer0_outputs(917)) and not (layer0_outputs(7692));
    outputs(8566) <= layer0_outputs(8892);
    outputs(8567) <= not((layer0_outputs(5656)) or (layer0_outputs(1915)));
    outputs(8568) <= not(layer0_outputs(8318));
    outputs(8569) <= layer0_outputs(9378);
    outputs(8570) <= not(layer0_outputs(11346)) or (layer0_outputs(3506));
    outputs(8571) <= layer0_outputs(5681);
    outputs(8572) <= not((layer0_outputs(12786)) xor (layer0_outputs(9105)));
    outputs(8573) <= not(layer0_outputs(5369));
    outputs(8574) <= layer0_outputs(7883);
    outputs(8575) <= layer0_outputs(4873);
    outputs(8576) <= layer0_outputs(4166);
    outputs(8577) <= layer0_outputs(7357);
    outputs(8578) <= layer0_outputs(639);
    outputs(8579) <= layer0_outputs(11382);
    outputs(8580) <= not(layer0_outputs(6882));
    outputs(8581) <= layer0_outputs(7711);
    outputs(8582) <= not(layer0_outputs(3531));
    outputs(8583) <= not(layer0_outputs(9881));
    outputs(8584) <= layer0_outputs(12411);
    outputs(8585) <= (layer0_outputs(9432)) and not (layer0_outputs(12441));
    outputs(8586) <= layer0_outputs(9878);
    outputs(8587) <= (layer0_outputs(9694)) xor (layer0_outputs(6242));
    outputs(8588) <= layer0_outputs(4888);
    outputs(8589) <= not(layer0_outputs(9616));
    outputs(8590) <= not(layer0_outputs(8821));
    outputs(8591) <= not(layer0_outputs(2630));
    outputs(8592) <= (layer0_outputs(5725)) xor (layer0_outputs(2956));
    outputs(8593) <= (layer0_outputs(3266)) and not (layer0_outputs(6372));
    outputs(8594) <= layer0_outputs(4390);
    outputs(8595) <= layer0_outputs(2681);
    outputs(8596) <= not(layer0_outputs(2229));
    outputs(8597) <= (layer0_outputs(6759)) and not (layer0_outputs(10830));
    outputs(8598) <= layer0_outputs(9618);
    outputs(8599) <= not(layer0_outputs(11696));
    outputs(8600) <= not(layer0_outputs(3046));
    outputs(8601) <= not(layer0_outputs(1705)) or (layer0_outputs(3325));
    outputs(8602) <= (layer0_outputs(3647)) and not (layer0_outputs(5456));
    outputs(8603) <= not((layer0_outputs(5268)) or (layer0_outputs(4956)));
    outputs(8604) <= (layer0_outputs(11953)) and (layer0_outputs(10028));
    outputs(8605) <= layer0_outputs(7705);
    outputs(8606) <= not((layer0_outputs(9988)) xor (layer0_outputs(10922)));
    outputs(8607) <= not((layer0_outputs(8891)) or (layer0_outputs(11092)));
    outputs(8608) <= not(layer0_outputs(9811)) or (layer0_outputs(4748));
    outputs(8609) <= layer0_outputs(12495);
    outputs(8610) <= layer0_outputs(3596);
    outputs(8611) <= not((layer0_outputs(4652)) xor (layer0_outputs(7329)));
    outputs(8612) <= (layer0_outputs(1395)) and (layer0_outputs(3291));
    outputs(8613) <= layer0_outputs(8234);
    outputs(8614) <= (layer0_outputs(12070)) and (layer0_outputs(2443));
    outputs(8615) <= (layer0_outputs(4300)) xor (layer0_outputs(3029));
    outputs(8616) <= not((layer0_outputs(490)) xor (layer0_outputs(8242)));
    outputs(8617) <= (layer0_outputs(6485)) or (layer0_outputs(5877));
    outputs(8618) <= not((layer0_outputs(9018)) xor (layer0_outputs(9434)));
    outputs(8619) <= not(layer0_outputs(5331));
    outputs(8620) <= not(layer0_outputs(9611));
    outputs(8621) <= not((layer0_outputs(4610)) and (layer0_outputs(3063)));
    outputs(8622) <= not(layer0_outputs(4948));
    outputs(8623) <= not((layer0_outputs(9536)) or (layer0_outputs(11113)));
    outputs(8624) <= layer0_outputs(10884);
    outputs(8625) <= not(layer0_outputs(7206));
    outputs(8626) <= not(layer0_outputs(12468));
    outputs(8627) <= layer0_outputs(11199);
    outputs(8628) <= layer0_outputs(7243);
    outputs(8629) <= not(layer0_outputs(10627));
    outputs(8630) <= (layer0_outputs(8401)) and not (layer0_outputs(8741));
    outputs(8631) <= not((layer0_outputs(10772)) xor (layer0_outputs(10619)));
    outputs(8632) <= layer0_outputs(4855);
    outputs(8633) <= (layer0_outputs(12483)) or (layer0_outputs(9711));
    outputs(8634) <= not((layer0_outputs(3809)) xor (layer0_outputs(10738)));
    outputs(8635) <= not(layer0_outputs(8217));
    outputs(8636) <= (layer0_outputs(11719)) xor (layer0_outputs(10014));
    outputs(8637) <= not((layer0_outputs(6814)) or (layer0_outputs(12041)));
    outputs(8638) <= layer0_outputs(7105);
    outputs(8639) <= layer0_outputs(7797);
    outputs(8640) <= layer0_outputs(5947);
    outputs(8641) <= not((layer0_outputs(5480)) and (layer0_outputs(8820)));
    outputs(8642) <= layer0_outputs(6570);
    outputs(8643) <= layer0_outputs(6100);
    outputs(8644) <= layer0_outputs(3103);
    outputs(8645) <= layer0_outputs(839);
    outputs(8646) <= not(layer0_outputs(10329)) or (layer0_outputs(38));
    outputs(8647) <= (layer0_outputs(980)) xor (layer0_outputs(5841));
    outputs(8648) <= not(layer0_outputs(7079)) or (layer0_outputs(2495));
    outputs(8649) <= not(layer0_outputs(10506));
    outputs(8650) <= layer0_outputs(3218);
    outputs(8651) <= (layer0_outputs(8149)) or (layer0_outputs(10317));
    outputs(8652) <= not((layer0_outputs(5639)) or (layer0_outputs(6116)));
    outputs(8653) <= not(layer0_outputs(4261));
    outputs(8654) <= (layer0_outputs(1634)) and not (layer0_outputs(8106));
    outputs(8655) <= not((layer0_outputs(7629)) xor (layer0_outputs(10669)));
    outputs(8656) <= layer0_outputs(10366);
    outputs(8657) <= layer0_outputs(820);
    outputs(8658) <= not(layer0_outputs(9866)) or (layer0_outputs(8334));
    outputs(8659) <= (layer0_outputs(139)) and not (layer0_outputs(2633));
    outputs(8660) <= (layer0_outputs(11271)) xor (layer0_outputs(2040));
    outputs(8661) <= not(layer0_outputs(11409));
    outputs(8662) <= not(layer0_outputs(7906));
    outputs(8663) <= not(layer0_outputs(10286));
    outputs(8664) <= not((layer0_outputs(12133)) xor (layer0_outputs(5946)));
    outputs(8665) <= layer0_outputs(3236);
    outputs(8666) <= not(layer0_outputs(6142)) or (layer0_outputs(6761));
    outputs(8667) <= (layer0_outputs(3198)) xor (layer0_outputs(10060));
    outputs(8668) <= not(layer0_outputs(12425));
    outputs(8669) <= not(layer0_outputs(5419));
    outputs(8670) <= layer0_outputs(6509);
    outputs(8671) <= (layer0_outputs(1422)) and not (layer0_outputs(8261));
    outputs(8672) <= not(layer0_outputs(1238));
    outputs(8673) <= not(layer0_outputs(6506));
    outputs(8674) <= not(layer0_outputs(8641));
    outputs(8675) <= layer0_outputs(323);
    outputs(8676) <= layer0_outputs(1742);
    outputs(8677) <= not((layer0_outputs(12690)) and (layer0_outputs(4435)));
    outputs(8678) <= layer0_outputs(545);
    outputs(8679) <= layer0_outputs(9026);
    outputs(8680) <= not(layer0_outputs(2488));
    outputs(8681) <= not(layer0_outputs(7916));
    outputs(8682) <= (layer0_outputs(10904)) xor (layer0_outputs(7909));
    outputs(8683) <= (layer0_outputs(10666)) xor (layer0_outputs(2813));
    outputs(8684) <= not(layer0_outputs(6065));
    outputs(8685) <= not(layer0_outputs(5501));
    outputs(8686) <= not(layer0_outputs(3117));
    outputs(8687) <= (layer0_outputs(6205)) xor (layer0_outputs(11151));
    outputs(8688) <= not(layer0_outputs(3962));
    outputs(8689) <= layer0_outputs(1878);
    outputs(8690) <= layer0_outputs(1400);
    outputs(8691) <= layer0_outputs(12661);
    outputs(8692) <= not(layer0_outputs(12232));
    outputs(8693) <= layer0_outputs(1036);
    outputs(8694) <= layer0_outputs(5497);
    outputs(8695) <= (layer0_outputs(7855)) and not (layer0_outputs(4639));
    outputs(8696) <= not(layer0_outputs(9319));
    outputs(8697) <= (layer0_outputs(12613)) xor (layer0_outputs(314));
    outputs(8698) <= not(layer0_outputs(3072));
    outputs(8699) <= layer0_outputs(7760);
    outputs(8700) <= layer0_outputs(2344);
    outputs(8701) <= not((layer0_outputs(12452)) xor (layer0_outputs(3519)));
    outputs(8702) <= (layer0_outputs(3115)) xor (layer0_outputs(11));
    outputs(8703) <= layer0_outputs(11334);
    outputs(8704) <= not(layer0_outputs(8823)) or (layer0_outputs(4225));
    outputs(8705) <= layer0_outputs(2439);
    outputs(8706) <= (layer0_outputs(5023)) xor (layer0_outputs(3499));
    outputs(8707) <= layer0_outputs(11563);
    outputs(8708) <= layer0_outputs(11915);
    outputs(8709) <= not(layer0_outputs(11304));
    outputs(8710) <= not(layer0_outputs(5771));
    outputs(8711) <= layer0_outputs(4289);
    outputs(8712) <= layer0_outputs(5072);
    outputs(8713) <= not(layer0_outputs(3541));
    outputs(8714) <= not(layer0_outputs(1773));
    outputs(8715) <= not(layer0_outputs(346));
    outputs(8716) <= (layer0_outputs(12065)) xor (layer0_outputs(3598));
    outputs(8717) <= layer0_outputs(8671);
    outputs(8718) <= not(layer0_outputs(5812));
    outputs(8719) <= layer0_outputs(11953);
    outputs(8720) <= not((layer0_outputs(2177)) or (layer0_outputs(1845)));
    outputs(8721) <= not(layer0_outputs(10394));
    outputs(8722) <= not(layer0_outputs(1456));
    outputs(8723) <= not(layer0_outputs(8206));
    outputs(8724) <= not((layer0_outputs(6085)) or (layer0_outputs(6092)));
    outputs(8725) <= not((layer0_outputs(3004)) xor (layer0_outputs(10)));
    outputs(8726) <= (layer0_outputs(11980)) and not (layer0_outputs(11612));
    outputs(8727) <= not((layer0_outputs(3693)) xor (layer0_outputs(4611)));
    outputs(8728) <= (layer0_outputs(10710)) xor (layer0_outputs(4960));
    outputs(8729) <= not(layer0_outputs(4681));
    outputs(8730) <= not(layer0_outputs(3163)) or (layer0_outputs(4035));
    outputs(8731) <= not(layer0_outputs(8375));
    outputs(8732) <= not(layer0_outputs(1258));
    outputs(8733) <= layer0_outputs(8395);
    outputs(8734) <= not((layer0_outputs(5811)) xor (layer0_outputs(8691)));
    outputs(8735) <= (layer0_outputs(2218)) xor (layer0_outputs(7130));
    outputs(8736) <= layer0_outputs(1020);
    outputs(8737) <= not(layer0_outputs(12040)) or (layer0_outputs(11978));
    outputs(8738) <= (layer0_outputs(1237)) xor (layer0_outputs(926));
    outputs(8739) <= not(layer0_outputs(2701));
    outputs(8740) <= layer0_outputs(6075);
    outputs(8741) <= layer0_outputs(1847);
    outputs(8742) <= (layer0_outputs(2467)) xor (layer0_outputs(8860));
    outputs(8743) <= layer0_outputs(742);
    outputs(8744) <= layer0_outputs(8699);
    outputs(8745) <= layer0_outputs(3952);
    outputs(8746) <= not(layer0_outputs(11467));
    outputs(8747) <= not(layer0_outputs(12581));
    outputs(8748) <= layer0_outputs(4490);
    outputs(8749) <= not((layer0_outputs(145)) or (layer0_outputs(11172)));
    outputs(8750) <= layer0_outputs(2250);
    outputs(8751) <= not(layer0_outputs(2009));
    outputs(8752) <= (layer0_outputs(2577)) and not (layer0_outputs(1975));
    outputs(8753) <= not(layer0_outputs(2291));
    outputs(8754) <= not(layer0_outputs(5377));
    outputs(8755) <= not(layer0_outputs(6054));
    outputs(8756) <= layer0_outputs(8979);
    outputs(8757) <= not(layer0_outputs(9419));
    outputs(8758) <= layer0_outputs(4580);
    outputs(8759) <= (layer0_outputs(1563)) and not (layer0_outputs(657));
    outputs(8760) <= layer0_outputs(12464);
    outputs(8761) <= layer0_outputs(4573);
    outputs(8762) <= layer0_outputs(9328);
    outputs(8763) <= (layer0_outputs(8324)) xor (layer0_outputs(5132));
    outputs(8764) <= (layer0_outputs(9608)) xor (layer0_outputs(7093));
    outputs(8765) <= not(layer0_outputs(7598)) or (layer0_outputs(2373));
    outputs(8766) <= layer0_outputs(11593);
    outputs(8767) <= not(layer0_outputs(4560)) or (layer0_outputs(9886));
    outputs(8768) <= not((layer0_outputs(3861)) xor (layer0_outputs(1681)));
    outputs(8769) <= (layer0_outputs(7830)) xor (layer0_outputs(11997));
    outputs(8770) <= (layer0_outputs(5994)) or (layer0_outputs(6183));
    outputs(8771) <= (layer0_outputs(8938)) and not (layer0_outputs(3766));
    outputs(8772) <= layer0_outputs(6790);
    outputs(8773) <= not((layer0_outputs(5456)) or (layer0_outputs(9794)));
    outputs(8774) <= not(layer0_outputs(11430));
    outputs(8775) <= not(layer0_outputs(10207)) or (layer0_outputs(11235));
    outputs(8776) <= layer0_outputs(3706);
    outputs(8777) <= layer0_outputs(7102);
    outputs(8778) <= layer0_outputs(1823);
    outputs(8779) <= not((layer0_outputs(11775)) or (layer0_outputs(7945)));
    outputs(8780) <= layer0_outputs(10197);
    outputs(8781) <= (layer0_outputs(7329)) xor (layer0_outputs(11041));
    outputs(8782) <= (layer0_outputs(4988)) xor (layer0_outputs(11359));
    outputs(8783) <= layer0_outputs(3116);
    outputs(8784) <= not(layer0_outputs(227));
    outputs(8785) <= not(layer0_outputs(4074)) or (layer0_outputs(284));
    outputs(8786) <= (layer0_outputs(5408)) and not (layer0_outputs(2203));
    outputs(8787) <= not((layer0_outputs(1338)) xor (layer0_outputs(2799)));
    outputs(8788) <= layer0_outputs(11201);
    outputs(8789) <= (layer0_outputs(3204)) xor (layer0_outputs(6748));
    outputs(8790) <= layer0_outputs(11260);
    outputs(8791) <= (layer0_outputs(8239)) and not (layer0_outputs(11994));
    outputs(8792) <= layer0_outputs(5253);
    outputs(8793) <= layer0_outputs(8472);
    outputs(8794) <= (layer0_outputs(7810)) and (layer0_outputs(5450));
    outputs(8795) <= layer0_outputs(10603);
    outputs(8796) <= not(layer0_outputs(6072));
    outputs(8797) <= (layer0_outputs(8111)) xor (layer0_outputs(1205));
    outputs(8798) <= layer0_outputs(2999);
    outputs(8799) <= not(layer0_outputs(12054));
    outputs(8800) <= (layer0_outputs(11437)) and not (layer0_outputs(5853));
    outputs(8801) <= not((layer0_outputs(8552)) or (layer0_outputs(10882)));
    outputs(8802) <= layer0_outputs(12209);
    outputs(8803) <= not(layer0_outputs(7538));
    outputs(8804) <= not(layer0_outputs(7094));
    outputs(8805) <= (layer0_outputs(10839)) xor (layer0_outputs(7178));
    outputs(8806) <= not(layer0_outputs(6602));
    outputs(8807) <= not(layer0_outputs(6175));
    outputs(8808) <= layer0_outputs(4876);
    outputs(8809) <= layer0_outputs(3846);
    outputs(8810) <= not(layer0_outputs(11521));
    outputs(8811) <= (layer0_outputs(11601)) and not (layer0_outputs(11760));
    outputs(8812) <= not(layer0_outputs(8103)) or (layer0_outputs(6463));
    outputs(8813) <= layer0_outputs(10523);
    outputs(8814) <= (layer0_outputs(11824)) and (layer0_outputs(2689));
    outputs(8815) <= (layer0_outputs(2408)) xor (layer0_outputs(5506));
    outputs(8816) <= not(layer0_outputs(9411));
    outputs(8817) <= (layer0_outputs(6066)) and (layer0_outputs(7989));
    outputs(8818) <= not((layer0_outputs(3408)) xor (layer0_outputs(9976)));
    outputs(8819) <= layer0_outputs(12400);
    outputs(8820) <= layer0_outputs(12062);
    outputs(8821) <= (layer0_outputs(4091)) and not (layer0_outputs(4026));
    outputs(8822) <= not((layer0_outputs(2069)) or (layer0_outputs(10374)));
    outputs(8823) <= layer0_outputs(10354);
    outputs(8824) <= not((layer0_outputs(6632)) xor (layer0_outputs(12002)));
    outputs(8825) <= not(layer0_outputs(568));
    outputs(8826) <= layer0_outputs(3137);
    outputs(8827) <= not(layer0_outputs(10786));
    outputs(8828) <= layer0_outputs(2285);
    outputs(8829) <= layer0_outputs(11772);
    outputs(8830) <= layer0_outputs(270);
    outputs(8831) <= not(layer0_outputs(767));
    outputs(8832) <= not(layer0_outputs(4919));
    outputs(8833) <= not(layer0_outputs(1502)) or (layer0_outputs(7441));
    outputs(8834) <= layer0_outputs(4257);
    outputs(8835) <= not(layer0_outputs(11739));
    outputs(8836) <= not((layer0_outputs(6234)) xor (layer0_outputs(3342)));
    outputs(8837) <= layer0_outputs(6734);
    outputs(8838) <= layer0_outputs(11744);
    outputs(8839) <= not(layer0_outputs(10043));
    outputs(8840) <= layer0_outputs(10875);
    outputs(8841) <= layer0_outputs(10469);
    outputs(8842) <= not(layer0_outputs(2782));
    outputs(8843) <= not(layer0_outputs(10050));
    outputs(8844) <= layer0_outputs(7402);
    outputs(8845) <= layer0_outputs(1796);
    outputs(8846) <= not((layer0_outputs(6628)) xor (layer0_outputs(11356)));
    outputs(8847) <= (layer0_outputs(9664)) and not (layer0_outputs(9713));
    outputs(8848) <= not(layer0_outputs(6405));
    outputs(8849) <= not(layer0_outputs(10447));
    outputs(8850) <= layer0_outputs(3041);
    outputs(8851) <= not((layer0_outputs(7828)) or (layer0_outputs(10277)));
    outputs(8852) <= (layer0_outputs(11212)) and not (layer0_outputs(1613));
    outputs(8853) <= not(layer0_outputs(11705));
    outputs(8854) <= not((layer0_outputs(1780)) and (layer0_outputs(4980)));
    outputs(8855) <= layer0_outputs(11957);
    outputs(8856) <= (layer0_outputs(3702)) xor (layer0_outputs(12064));
    outputs(8857) <= layer0_outputs(2491);
    outputs(8858) <= not((layer0_outputs(11338)) or (layer0_outputs(4629)));
    outputs(8859) <= (layer0_outputs(4357)) xor (layer0_outputs(1302));
    outputs(8860) <= not(layer0_outputs(6747));
    outputs(8861) <= not(layer0_outputs(1549));
    outputs(8862) <= not((layer0_outputs(10102)) or (layer0_outputs(10433)));
    outputs(8863) <= not(layer0_outputs(581));
    outputs(8864) <= not((layer0_outputs(3645)) or (layer0_outputs(11105)));
    outputs(8865) <= (layer0_outputs(12038)) xor (layer0_outputs(8700));
    outputs(8866) <= not(layer0_outputs(7366));
    outputs(8867) <= not(layer0_outputs(358));
    outputs(8868) <= not(layer0_outputs(4834));
    outputs(8869) <= not(layer0_outputs(8903)) or (layer0_outputs(1293));
    outputs(8870) <= (layer0_outputs(10031)) xor (layer0_outputs(190));
    outputs(8871) <= (layer0_outputs(3429)) and not (layer0_outputs(11584));
    outputs(8872) <= not(layer0_outputs(4586));
    outputs(8873) <= layer0_outputs(4242);
    outputs(8874) <= layer0_outputs(9184);
    outputs(8875) <= (layer0_outputs(3346)) and not (layer0_outputs(8898));
    outputs(8876) <= not(layer0_outputs(7341));
    outputs(8877) <= layer0_outputs(5056);
    outputs(8878) <= not(layer0_outputs(11462));
    outputs(8879) <= not(layer0_outputs(9807)) or (layer0_outputs(5053));
    outputs(8880) <= (layer0_outputs(3323)) xor (layer0_outputs(8635));
    outputs(8881) <= (layer0_outputs(10918)) xor (layer0_outputs(9997));
    outputs(8882) <= not((layer0_outputs(3709)) xor (layer0_outputs(8396)));
    outputs(8883) <= layer0_outputs(10995);
    outputs(8884) <= not(layer0_outputs(8805));
    outputs(8885) <= (layer0_outputs(6156)) and not (layer0_outputs(11877));
    outputs(8886) <= layer0_outputs(1582);
    outputs(8887) <= not(layer0_outputs(11664)) or (layer0_outputs(12431));
    outputs(8888) <= layer0_outputs(10740);
    outputs(8889) <= (layer0_outputs(7025)) and (layer0_outputs(4078));
    outputs(8890) <= not(layer0_outputs(5550));
    outputs(8891) <= (layer0_outputs(618)) xor (layer0_outputs(12769));
    outputs(8892) <= not((layer0_outputs(11781)) xor (layer0_outputs(3685)));
    outputs(8893) <= (layer0_outputs(12608)) and (layer0_outputs(12644));
    outputs(8894) <= not((layer0_outputs(11475)) or (layer0_outputs(10443)));
    outputs(8895) <= not((layer0_outputs(8837)) xor (layer0_outputs(5545)));
    outputs(8896) <= not(layer0_outputs(7891));
    outputs(8897) <= (layer0_outputs(6815)) and (layer0_outputs(8815));
    outputs(8898) <= not(layer0_outputs(9892));
    outputs(8899) <= layer0_outputs(7394);
    outputs(8900) <= (layer0_outputs(3851)) and not (layer0_outputs(2532));
    outputs(8901) <= not(layer0_outputs(12640));
    outputs(8902) <= not((layer0_outputs(6800)) xor (layer0_outputs(7210)));
    outputs(8903) <= (layer0_outputs(1583)) xor (layer0_outputs(2534));
    outputs(8904) <= (layer0_outputs(5466)) and (layer0_outputs(402));
    outputs(8905) <= layer0_outputs(3317);
    outputs(8906) <= (layer0_outputs(2428)) and not (layer0_outputs(1809));
    outputs(8907) <= layer0_outputs(11742);
    outputs(8908) <= (layer0_outputs(6330)) and not (layer0_outputs(248));
    outputs(8909) <= not((layer0_outputs(55)) or (layer0_outputs(6913)));
    outputs(8910) <= not(layer0_outputs(6795));
    outputs(8911) <= not(layer0_outputs(9106)) or (layer0_outputs(4340));
    outputs(8912) <= not((layer0_outputs(9200)) or (layer0_outputs(3513)));
    outputs(8913) <= (layer0_outputs(9329)) xor (layer0_outputs(10949));
    outputs(8914) <= layer0_outputs(3975);
    outputs(8915) <= (layer0_outputs(9220)) and not (layer0_outputs(2116));
    outputs(8916) <= (layer0_outputs(11839)) and not (layer0_outputs(12716));
    outputs(8917) <= not(layer0_outputs(6489));
    outputs(8918) <= not((layer0_outputs(10536)) xor (layer0_outputs(4353)));
    outputs(8919) <= layer0_outputs(12528);
    outputs(8920) <= not((layer0_outputs(5172)) xor (layer0_outputs(1689)));
    outputs(8921) <= layer0_outputs(2178);
    outputs(8922) <= not(layer0_outputs(6151));
    outputs(8923) <= not(layer0_outputs(1344));
    outputs(8924) <= (layer0_outputs(10131)) and not (layer0_outputs(5825));
    outputs(8925) <= not(layer0_outputs(4049));
    outputs(8926) <= (layer0_outputs(5170)) and not (layer0_outputs(7639));
    outputs(8927) <= (layer0_outputs(3451)) and not (layer0_outputs(3967));
    outputs(8928) <= layer0_outputs(3511);
    outputs(8929) <= (layer0_outputs(12499)) and not (layer0_outputs(8408));
    outputs(8930) <= layer0_outputs(4739);
    outputs(8931) <= (layer0_outputs(4298)) and not (layer0_outputs(4723));
    outputs(8932) <= not((layer0_outputs(9841)) or (layer0_outputs(8567)));
    outputs(8933) <= layer0_outputs(8230);
    outputs(8934) <= not(layer0_outputs(8580));
    outputs(8935) <= not(layer0_outputs(114));
    outputs(8936) <= (layer0_outputs(9591)) and not (layer0_outputs(4664));
    outputs(8937) <= layer0_outputs(10718);
    outputs(8938) <= (layer0_outputs(12780)) xor (layer0_outputs(12684));
    outputs(8939) <= (layer0_outputs(12097)) and not (layer0_outputs(4865));
    outputs(8940) <= layer0_outputs(3088);
    outputs(8941) <= layer0_outputs(4023);
    outputs(8942) <= not(layer0_outputs(8015));
    outputs(8943) <= layer0_outputs(2136);
    outputs(8944) <= not(layer0_outputs(9564));
    outputs(8945) <= layer0_outputs(8028);
    outputs(8946) <= layer0_outputs(375);
    outputs(8947) <= layer0_outputs(12650);
    outputs(8948) <= not(layer0_outputs(9985)) or (layer0_outputs(6445));
    outputs(8949) <= layer0_outputs(897);
    outputs(8950) <= layer0_outputs(2770);
    outputs(8951) <= not((layer0_outputs(7436)) or (layer0_outputs(7680)));
    outputs(8952) <= (layer0_outputs(2482)) and (layer0_outputs(6425));
    outputs(8953) <= not((layer0_outputs(9526)) and (layer0_outputs(8541)));
    outputs(8954) <= layer0_outputs(6605);
    outputs(8955) <= (layer0_outputs(8316)) and not (layer0_outputs(9486));
    outputs(8956) <= not((layer0_outputs(7894)) or (layer0_outputs(443)));
    outputs(8957) <= not(layer0_outputs(3194));
    outputs(8958) <= not((layer0_outputs(8059)) xor (layer0_outputs(8895)));
    outputs(8959) <= not((layer0_outputs(3639)) and (layer0_outputs(3275)));
    outputs(8960) <= not(layer0_outputs(6653));
    outputs(8961) <= not(layer0_outputs(9332));
    outputs(8962) <= layer0_outputs(3883);
    outputs(8963) <= not((layer0_outputs(12161)) and (layer0_outputs(1861)));
    outputs(8964) <= not((layer0_outputs(7526)) or (layer0_outputs(5033)));
    outputs(8965) <= layer0_outputs(8557);
    outputs(8966) <= not(layer0_outputs(4758));
    outputs(8967) <= layer0_outputs(1290);
    outputs(8968) <= not(layer0_outputs(9468));
    outputs(8969) <= not((layer0_outputs(11431)) and (layer0_outputs(3907)));
    outputs(8970) <= (layer0_outputs(9274)) and not (layer0_outputs(10768));
    outputs(8971) <= (layer0_outputs(5816)) and (layer0_outputs(1917));
    outputs(8972) <= not(layer0_outputs(7484));
    outputs(8973) <= (layer0_outputs(6417)) and not (layer0_outputs(12673));
    outputs(8974) <= layer0_outputs(12720);
    outputs(8975) <= (layer0_outputs(5051)) and not (layer0_outputs(1178));
    outputs(8976) <= not(layer0_outputs(11887));
    outputs(8977) <= (layer0_outputs(8684)) or (layer0_outputs(11828));
    outputs(8978) <= not(layer0_outputs(7676));
    outputs(8979) <= (layer0_outputs(3631)) and not (layer0_outputs(10728));
    outputs(8980) <= layer0_outputs(6875);
    outputs(8981) <= not(layer0_outputs(6055));
    outputs(8982) <= (layer0_outputs(11417)) and not (layer0_outputs(790));
    outputs(8983) <= not(layer0_outputs(5798));
    outputs(8984) <= not(layer0_outputs(5003));
    outputs(8985) <= layer0_outputs(1707);
    outputs(8986) <= layer0_outputs(12132);
    outputs(8987) <= (layer0_outputs(4394)) xor (layer0_outputs(1816));
    outputs(8988) <= not(layer0_outputs(7065));
    outputs(8989) <= layer0_outputs(10751);
    outputs(8990) <= (layer0_outputs(11187)) and not (layer0_outputs(2453));
    outputs(8991) <= '1';
    outputs(8992) <= not(layer0_outputs(10391));
    outputs(8993) <= layer0_outputs(11203);
    outputs(8994) <= not((layer0_outputs(12267)) and (layer0_outputs(12259)));
    outputs(8995) <= not(layer0_outputs(8839));
    outputs(8996) <= not((layer0_outputs(4771)) or (layer0_outputs(2332)));
    outputs(8997) <= (layer0_outputs(5248)) and (layer0_outputs(5662));
    outputs(8998) <= (layer0_outputs(3736)) xor (layer0_outputs(6840));
    outputs(8999) <= not(layer0_outputs(7418));
    outputs(9000) <= not((layer0_outputs(6014)) xor (layer0_outputs(6492)));
    outputs(9001) <= not(layer0_outputs(6888));
    outputs(9002) <= layer0_outputs(3466);
    outputs(9003) <= (layer0_outputs(1627)) and (layer0_outputs(5657));
    outputs(9004) <= not(layer0_outputs(11619));
    outputs(9005) <= layer0_outputs(7334);
    outputs(9006) <= not((layer0_outputs(4472)) xor (layer0_outputs(9930)));
    outputs(9007) <= layer0_outputs(7717);
    outputs(9008) <= (layer0_outputs(10618)) or (layer0_outputs(6495));
    outputs(9009) <= not((layer0_outputs(2303)) or (layer0_outputs(854)));
    outputs(9010) <= (layer0_outputs(11184)) and not (layer0_outputs(10070));
    outputs(9011) <= not(layer0_outputs(2389));
    outputs(9012) <= not((layer0_outputs(7720)) or (layer0_outputs(8119)));
    outputs(9013) <= not(layer0_outputs(724));
    outputs(9014) <= layer0_outputs(2029);
    outputs(9015) <= not(layer0_outputs(10700));
    outputs(9016) <= layer0_outputs(2593);
    outputs(9017) <= (layer0_outputs(5004)) xor (layer0_outputs(8989));
    outputs(9018) <= layer0_outputs(7030);
    outputs(9019) <= layer0_outputs(4805);
    outputs(9020) <= not(layer0_outputs(6152));
    outputs(9021) <= (layer0_outputs(9937)) and not (layer0_outputs(12486));
    outputs(9022) <= layer0_outputs(11142);
    outputs(9023) <= layer0_outputs(485);
    outputs(9024) <= layer0_outputs(5010);
    outputs(9025) <= (layer0_outputs(9458)) and not (layer0_outputs(11764));
    outputs(9026) <= layer0_outputs(1258);
    outputs(9027) <= not(layer0_outputs(1028));
    outputs(9028) <= not((layer0_outputs(9499)) xor (layer0_outputs(528)));
    outputs(9029) <= (layer0_outputs(1234)) xor (layer0_outputs(10527));
    outputs(9030) <= (layer0_outputs(12546)) and not (layer0_outputs(4600));
    outputs(9031) <= not(layer0_outputs(5150)) or (layer0_outputs(10533));
    outputs(9032) <= not((layer0_outputs(4122)) xor (layer0_outputs(7312)));
    outputs(9033) <= not((layer0_outputs(9601)) xor (layer0_outputs(204)));
    outputs(9034) <= not(layer0_outputs(9885));
    outputs(9035) <= (layer0_outputs(7562)) and (layer0_outputs(8058));
    outputs(9036) <= (layer0_outputs(7173)) xor (layer0_outputs(2023));
    outputs(9037) <= not(layer0_outputs(3016));
    outputs(9038) <= not((layer0_outputs(6230)) or (layer0_outputs(12438)));
    outputs(9039) <= (layer0_outputs(2411)) and (layer0_outputs(2742));
    outputs(9040) <= layer0_outputs(400);
    outputs(9041) <= (layer0_outputs(589)) xor (layer0_outputs(12091));
    outputs(9042) <= (layer0_outputs(5983)) or (layer0_outputs(6576));
    outputs(9043) <= '1';
    outputs(9044) <= (layer0_outputs(5350)) and not (layer0_outputs(2827));
    outputs(9045) <= not(layer0_outputs(2585));
    outputs(9046) <= not(layer0_outputs(11551));
    outputs(9047) <= (layer0_outputs(9455)) xor (layer0_outputs(4047));
    outputs(9048) <= not(layer0_outputs(10169));
    outputs(9049) <= layer0_outputs(6627);
    outputs(9050) <= not((layer0_outputs(9669)) xor (layer0_outputs(3928)));
    outputs(9051) <= not((layer0_outputs(9951)) or (layer0_outputs(11384)));
    outputs(9052) <= not(layer0_outputs(865));
    outputs(9053) <= not(layer0_outputs(12487));
    outputs(9054) <= layer0_outputs(5247);
    outputs(9055) <= not(layer0_outputs(7389));
    outputs(9056) <= (layer0_outputs(4123)) and not (layer0_outputs(11857));
    outputs(9057) <= not(layer0_outputs(3246));
    outputs(9058) <= not((layer0_outputs(9823)) and (layer0_outputs(5236)));
    outputs(9059) <= layer0_outputs(2523);
    outputs(9060) <= layer0_outputs(3184);
    outputs(9061) <= (layer0_outputs(10988)) and not (layer0_outputs(6094));
    outputs(9062) <= (layer0_outputs(7133)) and not (layer0_outputs(1958));
    outputs(9063) <= not(layer0_outputs(7733));
    outputs(9064) <= not(layer0_outputs(8689));
    outputs(9065) <= layer0_outputs(5131);
    outputs(9066) <= not((layer0_outputs(9164)) or (layer0_outputs(9126)));
    outputs(9067) <= layer0_outputs(11301);
    outputs(9068) <= not(layer0_outputs(11559));
    outputs(9069) <= (layer0_outputs(13)) and not (layer0_outputs(10594));
    outputs(9070) <= not((layer0_outputs(681)) xor (layer0_outputs(7192)));
    outputs(9071) <= not((layer0_outputs(1236)) xor (layer0_outputs(7520)));
    outputs(9072) <= not(layer0_outputs(4259));
    outputs(9073) <= (layer0_outputs(5941)) and (layer0_outputs(2905));
    outputs(9074) <= not(layer0_outputs(5243));
    outputs(9075) <= not(layer0_outputs(8652));
    outputs(9076) <= layer0_outputs(852);
    outputs(9077) <= not((layer0_outputs(1354)) xor (layer0_outputs(5507)));
    outputs(9078) <= (layer0_outputs(6322)) or (layer0_outputs(532));
    outputs(9079) <= not(layer0_outputs(11576));
    outputs(9080) <= (layer0_outputs(6018)) and not (layer0_outputs(9604));
    outputs(9081) <= not(layer0_outputs(2610));
    outputs(9082) <= layer0_outputs(10824);
    outputs(9083) <= not((layer0_outputs(11435)) or (layer0_outputs(4720)));
    outputs(9084) <= layer0_outputs(929);
    outputs(9085) <= not(layer0_outputs(6946));
    outputs(9086) <= (layer0_outputs(11863)) xor (layer0_outputs(4523));
    outputs(9087) <= layer0_outputs(7293);
    outputs(9088) <= layer0_outputs(9579);
    outputs(9089) <= not(layer0_outputs(7131));
    outputs(9090) <= layer0_outputs(12016);
    outputs(9091) <= (layer0_outputs(5848)) and not (layer0_outputs(8489));
    outputs(9092) <= not((layer0_outputs(603)) or (layer0_outputs(11942)));
    outputs(9093) <= (layer0_outputs(8653)) xor (layer0_outputs(3228));
    outputs(9094) <= layer0_outputs(623);
    outputs(9095) <= layer0_outputs(906);
    outputs(9096) <= (layer0_outputs(974)) and not (layer0_outputs(6025));
    outputs(9097) <= not(layer0_outputs(3668));
    outputs(9098) <= not(layer0_outputs(9395));
    outputs(9099) <= (layer0_outputs(1150)) and not (layer0_outputs(11564));
    outputs(9100) <= not((layer0_outputs(4117)) or (layer0_outputs(10205)));
    outputs(9101) <= (layer0_outputs(11983)) xor (layer0_outputs(8982));
    outputs(9102) <= not(layer0_outputs(8765));
    outputs(9103) <= layer0_outputs(6538);
    outputs(9104) <= not(layer0_outputs(7462));
    outputs(9105) <= (layer0_outputs(3378)) and (layer0_outputs(1755));
    outputs(9106) <= (layer0_outputs(9333)) and (layer0_outputs(1900));
    outputs(9107) <= (layer0_outputs(5619)) and not (layer0_outputs(11127));
    outputs(9108) <= layer0_outputs(11914);
    outputs(9109) <= layer0_outputs(4069);
    outputs(9110) <= layer0_outputs(4187);
    outputs(9111) <= not((layer0_outputs(6281)) or (layer0_outputs(12260)));
    outputs(9112) <= not(layer0_outputs(10749));
    outputs(9113) <= not((layer0_outputs(2015)) and (layer0_outputs(5054)));
    outputs(9114) <= layer0_outputs(8757);
    outputs(9115) <= not(layer0_outputs(1318));
    outputs(9116) <= (layer0_outputs(8029)) xor (layer0_outputs(4993));
    outputs(9117) <= (layer0_outputs(4099)) and not (layer0_outputs(2184));
    outputs(9118) <= layer0_outputs(12462);
    outputs(9119) <= not((layer0_outputs(2794)) and (layer0_outputs(7387)));
    outputs(9120) <= layer0_outputs(8325);
    outputs(9121) <= (layer0_outputs(7580)) and not (layer0_outputs(10644));
    outputs(9122) <= (layer0_outputs(1105)) and not (layer0_outputs(5433));
    outputs(9123) <= not(layer0_outputs(6341));
    outputs(9124) <= not((layer0_outputs(368)) and (layer0_outputs(11740)));
    outputs(9125) <= layer0_outputs(1221);
    outputs(9126) <= layer0_outputs(7043);
    outputs(9127) <= not(layer0_outputs(10007));
    outputs(9128) <= (layer0_outputs(11842)) and not (layer0_outputs(2031));
    outputs(9129) <= not((layer0_outputs(4065)) or (layer0_outputs(4038)));
    outputs(9130) <= not(layer0_outputs(10412));
    outputs(9131) <= (layer0_outputs(12546)) and (layer0_outputs(8546));
    outputs(9132) <= layer0_outputs(11169);
    outputs(9133) <= layer0_outputs(5787);
    outputs(9134) <= not((layer0_outputs(6836)) xor (layer0_outputs(10947)));
    outputs(9135) <= not(layer0_outputs(857));
    outputs(9136) <= layer0_outputs(10163);
    outputs(9137) <= layer0_outputs(5543);
    outputs(9138) <= not(layer0_outputs(6410)) or (layer0_outputs(54));
    outputs(9139) <= layer0_outputs(9708);
    outputs(9140) <= (layer0_outputs(6454)) and (layer0_outputs(8758));
    outputs(9141) <= not(layer0_outputs(2375));
    outputs(9142) <= (layer0_outputs(1301)) and (layer0_outputs(8669));
    outputs(9143) <= not((layer0_outputs(7083)) xor (layer0_outputs(4800)));
    outputs(9144) <= not(layer0_outputs(3821));
    outputs(9145) <= layer0_outputs(5068);
    outputs(9146) <= not(layer0_outputs(253));
    outputs(9147) <= not((layer0_outputs(4283)) xor (layer0_outputs(2670)));
    outputs(9148) <= (layer0_outputs(7866)) xor (layer0_outputs(8723));
    outputs(9149) <= not((layer0_outputs(10602)) or (layer0_outputs(4532)));
    outputs(9150) <= not(layer0_outputs(12291));
    outputs(9151) <= not((layer0_outputs(3626)) xor (layer0_outputs(7497)));
    outputs(9152) <= not((layer0_outputs(2161)) or (layer0_outputs(10885)));
    outputs(9153) <= not(layer0_outputs(4087));
    outputs(9154) <= layer0_outputs(2151);
    outputs(9155) <= not(layer0_outputs(4426));
    outputs(9156) <= layer0_outputs(12380);
    outputs(9157) <= not((layer0_outputs(7434)) xor (layer0_outputs(8006)));
    outputs(9158) <= not(layer0_outputs(3155));
    outputs(9159) <= not(layer0_outputs(855)) or (layer0_outputs(8909));
    outputs(9160) <= not(layer0_outputs(56));
    outputs(9161) <= not(layer0_outputs(12291));
    outputs(9162) <= layer0_outputs(3553);
    outputs(9163) <= (layer0_outputs(7452)) xor (layer0_outputs(11355));
    outputs(9164) <= not((layer0_outputs(3744)) or (layer0_outputs(3269)));
    outputs(9165) <= not(layer0_outputs(4524)) or (layer0_outputs(11973));
    outputs(9166) <= not((layer0_outputs(5462)) or (layer0_outputs(11139)));
    outputs(9167) <= (layer0_outputs(8429)) and not (layer0_outputs(2781));
    outputs(9168) <= not(layer0_outputs(4266));
    outputs(9169) <= (layer0_outputs(8036)) and (layer0_outputs(10223));
    outputs(9170) <= layer0_outputs(4165);
    outputs(9171) <= layer0_outputs(848);
    outputs(9172) <= layer0_outputs(7583);
    outputs(9173) <= (layer0_outputs(6172)) and not (layer0_outputs(10167));
    outputs(9174) <= layer0_outputs(5657);
    outputs(9175) <= not(layer0_outputs(4608));
    outputs(9176) <= (layer0_outputs(7603)) xor (layer0_outputs(8074));
    outputs(9177) <= layer0_outputs(8220);
    outputs(9178) <= (layer0_outputs(5377)) and not (layer0_outputs(1257));
    outputs(9179) <= layer0_outputs(8977);
    outputs(9180) <= (layer0_outputs(5008)) and (layer0_outputs(11969));
    outputs(9181) <= (layer0_outputs(8642)) xor (layer0_outputs(3212));
    outputs(9182) <= layer0_outputs(7616);
    outputs(9183) <= (layer0_outputs(8446)) xor (layer0_outputs(1511));
    outputs(9184) <= not(layer0_outputs(2193)) or (layer0_outputs(10955));
    outputs(9185) <= (layer0_outputs(1807)) and (layer0_outputs(1212));
    outputs(9186) <= layer0_outputs(4092);
    outputs(9187) <= not(layer0_outputs(12480)) or (layer0_outputs(7342));
    outputs(9188) <= not(layer0_outputs(9331));
    outputs(9189) <= layer0_outputs(10692);
    outputs(9190) <= not(layer0_outputs(11399));
    outputs(9191) <= (layer0_outputs(11975)) xor (layer0_outputs(44));
    outputs(9192) <= (layer0_outputs(7352)) and (layer0_outputs(5650));
    outputs(9193) <= (layer0_outputs(5220)) and not (layer0_outputs(10172));
    outputs(9194) <= (layer0_outputs(1457)) and not (layer0_outputs(824));
    outputs(9195) <= not((layer0_outputs(11180)) xor (layer0_outputs(11473)));
    outputs(9196) <= layer0_outputs(9208);
    outputs(9197) <= not((layer0_outputs(3763)) or (layer0_outputs(11200)));
    outputs(9198) <= (layer0_outputs(723)) and not (layer0_outputs(10748));
    outputs(9199) <= (layer0_outputs(3205)) xor (layer0_outputs(7875));
    outputs(9200) <= layer0_outputs(3867);
    outputs(9201) <= not(layer0_outputs(3527)) or (layer0_outputs(2451));
    outputs(9202) <= not(layer0_outputs(11160));
    outputs(9203) <= layer0_outputs(306);
    outputs(9204) <= not((layer0_outputs(6922)) and (layer0_outputs(10557)));
    outputs(9205) <= layer0_outputs(2836);
    outputs(9206) <= not(layer0_outputs(7226));
    outputs(9207) <= layer0_outputs(7424);
    outputs(9208) <= not(layer0_outputs(10935)) or (layer0_outputs(9643));
    outputs(9209) <= not(layer0_outputs(610));
    outputs(9210) <= not(layer0_outputs(6111));
    outputs(9211) <= not((layer0_outputs(242)) xor (layer0_outputs(1176)));
    outputs(9212) <= layer0_outputs(6195);
    outputs(9213) <= not((layer0_outputs(1598)) and (layer0_outputs(8689)));
    outputs(9214) <= layer0_outputs(12467);
    outputs(9215) <= not(layer0_outputs(5487));
    outputs(9216) <= not(layer0_outputs(9123));
    outputs(9217) <= (layer0_outputs(3469)) and not (layer0_outputs(3330));
    outputs(9218) <= not(layer0_outputs(2706));
    outputs(9219) <= (layer0_outputs(1244)) and not (layer0_outputs(9409));
    outputs(9220) <= (layer0_outputs(12067)) and (layer0_outputs(9075));
    outputs(9221) <= layer0_outputs(5804);
    outputs(9222) <= not((layer0_outputs(11218)) or (layer0_outputs(10600)));
    outputs(9223) <= (layer0_outputs(2229)) and not (layer0_outputs(3781));
    outputs(9224) <= not(layer0_outputs(12516)) or (layer0_outputs(3645));
    outputs(9225) <= not(layer0_outputs(3650));
    outputs(9226) <= not((layer0_outputs(4899)) or (layer0_outputs(11818)));
    outputs(9227) <= layer0_outputs(12231);
    outputs(9228) <= (layer0_outputs(8897)) or (layer0_outputs(7738));
    outputs(9229) <= (layer0_outputs(10243)) and (layer0_outputs(7410));
    outputs(9230) <= not((layer0_outputs(8418)) xor (layer0_outputs(3539)));
    outputs(9231) <= layer0_outputs(5233);
    outputs(9232) <= layer0_outputs(1094);
    outputs(9233) <= (layer0_outputs(10505)) and not (layer0_outputs(12268));
    outputs(9234) <= not(layer0_outputs(3802));
    outputs(9235) <= not(layer0_outputs(2849));
    outputs(9236) <= (layer0_outputs(5296)) xor (layer0_outputs(3157));
    outputs(9237) <= layer0_outputs(10423);
    outputs(9238) <= (layer0_outputs(2680)) and not (layer0_outputs(3283));
    outputs(9239) <= (layer0_outputs(3076)) and (layer0_outputs(11909));
    outputs(9240) <= not((layer0_outputs(11583)) or (layer0_outputs(8609)));
    outputs(9241) <= not(layer0_outputs(11719));
    outputs(9242) <= (layer0_outputs(9689)) and not (layer0_outputs(9047));
    outputs(9243) <= not((layer0_outputs(497)) and (layer0_outputs(6717)));
    outputs(9244) <= not(layer0_outputs(4242));
    outputs(9245) <= not(layer0_outputs(5191)) or (layer0_outputs(2085));
    outputs(9246) <= not(layer0_outputs(7575));
    outputs(9247) <= layer0_outputs(11602);
    outputs(9248) <= (layer0_outputs(6053)) and not (layer0_outputs(12582));
    outputs(9249) <= not((layer0_outputs(12704)) xor (layer0_outputs(12479)));
    outputs(9250) <= not((layer0_outputs(2021)) or (layer0_outputs(9796)));
    outputs(9251) <= not((layer0_outputs(9291)) or (layer0_outputs(11223)));
    outputs(9252) <= layer0_outputs(723);
    outputs(9253) <= not((layer0_outputs(7437)) or (layer0_outputs(11999)));
    outputs(9254) <= (layer0_outputs(6538)) and not (layer0_outputs(12716));
    outputs(9255) <= layer0_outputs(6812);
    outputs(9256) <= not((layer0_outputs(6528)) xor (layer0_outputs(12357)));
    outputs(9257) <= not(layer0_outputs(4379));
    outputs(9258) <= (layer0_outputs(4068)) xor (layer0_outputs(914));
    outputs(9259) <= not(layer0_outputs(8528));
    outputs(9260) <= (layer0_outputs(8131)) and not (layer0_outputs(6631));
    outputs(9261) <= layer0_outputs(10590);
    outputs(9262) <= (layer0_outputs(1287)) and (layer0_outputs(6866));
    outputs(9263) <= (layer0_outputs(11032)) xor (layer0_outputs(10228));
    outputs(9264) <= not(layer0_outputs(2143));
    outputs(9265) <= not((layer0_outputs(10379)) xor (layer0_outputs(5355)));
    outputs(9266) <= (layer0_outputs(7985)) and not (layer0_outputs(11735));
    outputs(9267) <= not(layer0_outputs(4929));
    outputs(9268) <= not(layer0_outputs(4273)) or (layer0_outputs(397));
    outputs(9269) <= layer0_outputs(12628);
    outputs(9270) <= (layer0_outputs(6861)) and not (layer0_outputs(10672));
    outputs(9271) <= not((layer0_outputs(5357)) or (layer0_outputs(9385)));
    outputs(9272) <= (layer0_outputs(4958)) and not (layer0_outputs(6597));
    outputs(9273) <= (layer0_outputs(11857)) xor (layer0_outputs(12712));
    outputs(9274) <= (layer0_outputs(10324)) and (layer0_outputs(9283));
    outputs(9275) <= layer0_outputs(6609);
    outputs(9276) <= not(layer0_outputs(1525));
    outputs(9277) <= not((layer0_outputs(3892)) xor (layer0_outputs(1968)));
    outputs(9278) <= not(layer0_outputs(6115));
    outputs(9279) <= layer0_outputs(11185);
    outputs(9280) <= not((layer0_outputs(2951)) or (layer0_outputs(2105)));
    outputs(9281) <= (layer0_outputs(3421)) xor (layer0_outputs(10701));
    outputs(9282) <= not(layer0_outputs(3793));
    outputs(9283) <= layer0_outputs(1573);
    outputs(9284) <= not((layer0_outputs(5905)) or (layer0_outputs(1082)));
    outputs(9285) <= not((layer0_outputs(7279)) or (layer0_outputs(1583)));
    outputs(9286) <= layer0_outputs(5689);
    outputs(9287) <= (layer0_outputs(11267)) xor (layer0_outputs(12063));
    outputs(9288) <= not(layer0_outputs(5102));
    outputs(9289) <= not(layer0_outputs(7826));
    outputs(9290) <= layer0_outputs(1188);
    outputs(9291) <= layer0_outputs(10865);
    outputs(9292) <= layer0_outputs(7740);
    outputs(9293) <= layer0_outputs(7709);
    outputs(9294) <= not(layer0_outputs(4802));
    outputs(9295) <= (layer0_outputs(480)) and (layer0_outputs(8978));
    outputs(9296) <= not((layer0_outputs(6121)) or (layer0_outputs(1509)));
    outputs(9297) <= not(layer0_outputs(8919)) or (layer0_outputs(6913));
    outputs(9298) <= not((layer0_outputs(11488)) and (layer0_outputs(6690)));
    outputs(9299) <= not(layer0_outputs(1341));
    outputs(9300) <= not(layer0_outputs(1530));
    outputs(9301) <= (layer0_outputs(6611)) xor (layer0_outputs(6477));
    outputs(9302) <= (layer0_outputs(11789)) xor (layer0_outputs(11796));
    outputs(9303) <= not(layer0_outputs(11123));
    outputs(9304) <= (layer0_outputs(6025)) xor (layer0_outputs(2923));
    outputs(9305) <= not((layer0_outputs(1709)) and (layer0_outputs(8201)));
    outputs(9306) <= layer0_outputs(4027);
    outputs(9307) <= (layer0_outputs(7912)) and not (layer0_outputs(7380));
    outputs(9308) <= layer0_outputs(8835);
    outputs(9309) <= (layer0_outputs(8690)) xor (layer0_outputs(11219));
    outputs(9310) <= not(layer0_outputs(8932));
    outputs(9311) <= (layer0_outputs(5574)) xor (layer0_outputs(6642));
    outputs(9312) <= (layer0_outputs(8422)) xor (layer0_outputs(9764));
    outputs(9313) <= layer0_outputs(2058);
    outputs(9314) <= layer0_outputs(5390);
    outputs(9315) <= not(layer0_outputs(1785));
    outputs(9316) <= (layer0_outputs(10864)) xor (layer0_outputs(9944));
    outputs(9317) <= not(layer0_outputs(3951));
    outputs(9318) <= (layer0_outputs(1417)) xor (layer0_outputs(3488));
    outputs(9319) <= layer0_outputs(6398);
    outputs(9320) <= layer0_outputs(8638);
    outputs(9321) <= layer0_outputs(265);
    outputs(9322) <= not(layer0_outputs(1315));
    outputs(9323) <= (layer0_outputs(6113)) and not (layer0_outputs(12250));
    outputs(9324) <= layer0_outputs(2458);
    outputs(9325) <= not(layer0_outputs(2294));
    outputs(9326) <= not((layer0_outputs(2103)) and (layer0_outputs(2306)));
    outputs(9327) <= (layer0_outputs(9944)) and not (layer0_outputs(7633));
    outputs(9328) <= not(layer0_outputs(7993)) or (layer0_outputs(7486));
    outputs(9329) <= not(layer0_outputs(12530));
    outputs(9330) <= (layer0_outputs(9566)) and not (layer0_outputs(4210));
    outputs(9331) <= not(layer0_outputs(2585));
    outputs(9332) <= layer0_outputs(4940);
    outputs(9333) <= not(layer0_outputs(6429)) or (layer0_outputs(2580));
    outputs(9334) <= layer0_outputs(8802);
    outputs(9335) <= not(layer0_outputs(6248));
    outputs(9336) <= not(layer0_outputs(1835));
    outputs(9337) <= (layer0_outputs(6337)) and (layer0_outputs(5851));
    outputs(9338) <= not(layer0_outputs(11075));
    outputs(9339) <= not(layer0_outputs(8809));
    outputs(9340) <= (layer0_outputs(10755)) and not (layer0_outputs(11113));
    outputs(9341) <= layer0_outputs(2972);
    outputs(9342) <= layer0_outputs(3780);
    outputs(9343) <= layer0_outputs(8077);
    outputs(9344) <= not(layer0_outputs(11008));
    outputs(9345) <= layer0_outputs(9357);
    outputs(9346) <= (layer0_outputs(11216)) and (layer0_outputs(3387));
    outputs(9347) <= not(layer0_outputs(4749));
    outputs(9348) <= (layer0_outputs(2926)) and not (layer0_outputs(4695));
    outputs(9349) <= not(layer0_outputs(5929));
    outputs(9350) <= (layer0_outputs(673)) and not (layer0_outputs(12245));
    outputs(9351) <= layer0_outputs(1502);
    outputs(9352) <= not(layer0_outputs(5359));
    outputs(9353) <= (layer0_outputs(6146)) and not (layer0_outputs(552));
    outputs(9354) <= not(layer0_outputs(316));
    outputs(9355) <= not(layer0_outputs(2534));
    outputs(9356) <= layer0_outputs(4609);
    outputs(9357) <= (layer0_outputs(5067)) and not (layer0_outputs(4758));
    outputs(9358) <= layer0_outputs(9592);
    outputs(9359) <= (layer0_outputs(10521)) and (layer0_outputs(12591));
    outputs(9360) <= not(layer0_outputs(1547));
    outputs(9361) <= not((layer0_outputs(3292)) or (layer0_outputs(11985)));
    outputs(9362) <= (layer0_outputs(580)) and (layer0_outputs(4250));
    outputs(9363) <= (layer0_outputs(12645)) xor (layer0_outputs(2531));
    outputs(9364) <= not(layer0_outputs(734));
    outputs(9365) <= layer0_outputs(4194);
    outputs(9366) <= layer0_outputs(3482);
    outputs(9367) <= not(layer0_outputs(7588));
    outputs(9368) <= (layer0_outputs(3818)) or (layer0_outputs(10437));
    outputs(9369) <= (layer0_outputs(5475)) or (layer0_outputs(7253));
    outputs(9370) <= not(layer0_outputs(2872));
    outputs(9371) <= layer0_outputs(78);
    outputs(9372) <= (layer0_outputs(773)) xor (layer0_outputs(8353));
    outputs(9373) <= not((layer0_outputs(9480)) xor (layer0_outputs(750)));
    outputs(9374) <= not(layer0_outputs(2530)) or (layer0_outputs(5969));
    outputs(9375) <= layer0_outputs(10177);
    outputs(9376) <= (layer0_outputs(2007)) xor (layer0_outputs(7495));
    outputs(9377) <= (layer0_outputs(7661)) and (layer0_outputs(12302));
    outputs(9378) <= layer0_outputs(1197);
    outputs(9379) <= not(layer0_outputs(12205));
    outputs(9380) <= not(layer0_outputs(11445)) or (layer0_outputs(6729));
    outputs(9381) <= (layer0_outputs(5063)) or (layer0_outputs(11154));
    outputs(9382) <= layer0_outputs(11637);
    outputs(9383) <= layer0_outputs(12447);
    outputs(9384) <= not((layer0_outputs(12458)) or (layer0_outputs(9460)));
    outputs(9385) <= (layer0_outputs(3719)) and (layer0_outputs(6487));
    outputs(9386) <= layer0_outputs(7443);
    outputs(9387) <= not(layer0_outputs(11168));
    outputs(9388) <= (layer0_outputs(2347)) and not (layer0_outputs(11753));
    outputs(9389) <= layer0_outputs(9912);
    outputs(9390) <= layer0_outputs(9574);
    outputs(9391) <= not((layer0_outputs(7713)) or (layer0_outputs(5799)));
    outputs(9392) <= not(layer0_outputs(9705));
    outputs(9393) <= not((layer0_outputs(7875)) and (layer0_outputs(6426)));
    outputs(9394) <= layer0_outputs(5812);
    outputs(9395) <= not((layer0_outputs(3575)) xor (layer0_outputs(7947)));
    outputs(9396) <= layer0_outputs(1064);
    outputs(9397) <= not(layer0_outputs(9543));
    outputs(9398) <= not(layer0_outputs(11179));
    outputs(9399) <= not((layer0_outputs(3542)) xor (layer0_outputs(2321)));
    outputs(9400) <= not((layer0_outputs(11982)) or (layer0_outputs(12400)));
    outputs(9401) <= not((layer0_outputs(11571)) or (layer0_outputs(4809)));
    outputs(9402) <= not(layer0_outputs(761));
    outputs(9403) <= layer0_outputs(4015);
    outputs(9404) <= not((layer0_outputs(2924)) or (layer0_outputs(5016)));
    outputs(9405) <= (layer0_outputs(10051)) and not (layer0_outputs(2024));
    outputs(9406) <= layer0_outputs(6459);
    outputs(9407) <= layer0_outputs(2904);
    outputs(9408) <= (layer0_outputs(12748)) and (layer0_outputs(11205));
    outputs(9409) <= (layer0_outputs(5226)) and (layer0_outputs(10631));
    outputs(9410) <= not(layer0_outputs(8882));
    outputs(9411) <= (layer0_outputs(11823)) and not (layer0_outputs(2778));
    outputs(9412) <= layer0_outputs(2703);
    outputs(9413) <= layer0_outputs(6038);
    outputs(9414) <= not(layer0_outputs(3975));
    outputs(9415) <= (layer0_outputs(6239)) xor (layer0_outputs(2399));
    outputs(9416) <= (layer0_outputs(4099)) and not (layer0_outputs(7525));
    outputs(9417) <= not(layer0_outputs(5772));
    outputs(9418) <= (layer0_outputs(8491)) and not (layer0_outputs(505));
    outputs(9419) <= not(layer0_outputs(339));
    outputs(9420) <= (layer0_outputs(4866)) and (layer0_outputs(6453));
    outputs(9421) <= layer0_outputs(6019);
    outputs(9422) <= not((layer0_outputs(6445)) xor (layer0_outputs(1333)));
    outputs(9423) <= (layer0_outputs(2360)) or (layer0_outputs(9078));
    outputs(9424) <= layer0_outputs(3114);
    outputs(9425) <= not(layer0_outputs(2699));
    outputs(9426) <= (layer0_outputs(5862)) and (layer0_outputs(1500));
    outputs(9427) <= not((layer0_outputs(11908)) xor (layer0_outputs(9491)));
    outputs(9428) <= not((layer0_outputs(5235)) xor (layer0_outputs(4756)));
    outputs(9429) <= (layer0_outputs(2319)) and (layer0_outputs(8693));
    outputs(9430) <= (layer0_outputs(11994)) xor (layer0_outputs(256));
    outputs(9431) <= not(layer0_outputs(4573));
    outputs(9432) <= (layer0_outputs(617)) or (layer0_outputs(8065));
    outputs(9433) <= not(layer0_outputs(11405));
    outputs(9434) <= not(layer0_outputs(1945)) or (layer0_outputs(8226));
    outputs(9435) <= layer0_outputs(6095);
    outputs(9436) <= layer0_outputs(9837);
    outputs(9437) <= layer0_outputs(2819);
    outputs(9438) <= (layer0_outputs(7463)) and not (layer0_outputs(1513));
    outputs(9439) <= layer0_outputs(6333);
    outputs(9440) <= layer0_outputs(9650);
    outputs(9441) <= not((layer0_outputs(2824)) xor (layer0_outputs(286)));
    outputs(9442) <= not((layer0_outputs(2724)) or (layer0_outputs(7128)));
    outputs(9443) <= not(layer0_outputs(5236));
    outputs(9444) <= not(layer0_outputs(2662));
    outputs(9445) <= (layer0_outputs(7022)) and not (layer0_outputs(8151));
    outputs(9446) <= layer0_outputs(1227);
    outputs(9447) <= layer0_outputs(9529);
    outputs(9448) <= layer0_outputs(8375);
    outputs(9449) <= not((layer0_outputs(9968)) or (layer0_outputs(2600)));
    outputs(9450) <= (layer0_outputs(10958)) xor (layer0_outputs(4778));
    outputs(9451) <= layer0_outputs(1246);
    outputs(9452) <= layer0_outputs(3740);
    outputs(9453) <= not(layer0_outputs(395));
    outputs(9454) <= not(layer0_outputs(4660));
    outputs(9455) <= not(layer0_outputs(4663));
    outputs(9456) <= not(layer0_outputs(1163));
    outputs(9457) <= not((layer0_outputs(8790)) xor (layer0_outputs(6464)));
    outputs(9458) <= layer0_outputs(167);
    outputs(9459) <= not((layer0_outputs(4434)) or (layer0_outputs(2410)));
    outputs(9460) <= not(layer0_outputs(1935));
    outputs(9461) <= not(layer0_outputs(5800));
    outputs(9462) <= not(layer0_outputs(6263));
    outputs(9463) <= layer0_outputs(5232);
    outputs(9464) <= (layer0_outputs(3249)) and (layer0_outputs(365));
    outputs(9465) <= layer0_outputs(5554);
    outputs(9466) <= layer0_outputs(6116);
    outputs(9467) <= (layer0_outputs(8669)) xor (layer0_outputs(11164));
    outputs(9468) <= (layer0_outputs(7670)) xor (layer0_outputs(1006));
    outputs(9469) <= not((layer0_outputs(489)) and (layer0_outputs(10273)));
    outputs(9470) <= not(layer0_outputs(1151));
    outputs(9471) <= (layer0_outputs(5500)) and not (layer0_outputs(1294));
    outputs(9472) <= not(layer0_outputs(3383));
    outputs(9473) <= (layer0_outputs(10336)) and (layer0_outputs(12568));
    outputs(9474) <= layer0_outputs(2102);
    outputs(9475) <= not(layer0_outputs(11518));
    outputs(9476) <= layer0_outputs(2537);
    outputs(9477) <= not(layer0_outputs(10444));
    outputs(9478) <= not((layer0_outputs(10308)) xor (layer0_outputs(7507)));
    outputs(9479) <= not(layer0_outputs(8747));
    outputs(9480) <= not((layer0_outputs(4927)) or (layer0_outputs(2691)));
    outputs(9481) <= layer0_outputs(355);
    outputs(9482) <= layer0_outputs(11189);
    outputs(9483) <= not(layer0_outputs(7569));
    outputs(9484) <= not(layer0_outputs(11929));
    outputs(9485) <= not((layer0_outputs(3900)) xor (layer0_outputs(4005)));
    outputs(9486) <= (layer0_outputs(8494)) xor (layer0_outputs(8983));
    outputs(9487) <= not((layer0_outputs(11044)) or (layer0_outputs(9410)));
    outputs(9488) <= (layer0_outputs(10066)) and not (layer0_outputs(5395));
    outputs(9489) <= not((layer0_outputs(7398)) xor (layer0_outputs(12721)));
    outputs(9490) <= layer0_outputs(6958);
    outputs(9491) <= (layer0_outputs(10480)) or (layer0_outputs(2570));
    outputs(9492) <= (layer0_outputs(12477)) and (layer0_outputs(8535));
    outputs(9493) <= not((layer0_outputs(7084)) or (layer0_outputs(11981)));
    outputs(9494) <= (layer0_outputs(1365)) xor (layer0_outputs(7228));
    outputs(9495) <= not(layer0_outputs(2312));
    outputs(9496) <= not(layer0_outputs(2310));
    outputs(9497) <= (layer0_outputs(4108)) xor (layer0_outputs(5589));
    outputs(9498) <= layer0_outputs(9459);
    outputs(9499) <= (layer0_outputs(11886)) and not (layer0_outputs(11550));
    outputs(9500) <= not(layer0_outputs(8327));
    outputs(9501) <= layer0_outputs(9894);
    outputs(9502) <= layer0_outputs(12534);
    outputs(9503) <= not(layer0_outputs(3949));
    outputs(9504) <= layer0_outputs(8444);
    outputs(9505) <= not(layer0_outputs(9770));
    outputs(9506) <= not((layer0_outputs(9431)) or (layer0_outputs(11437)));
    outputs(9507) <= (layer0_outputs(160)) and not (layer0_outputs(3548));
    outputs(9508) <= (layer0_outputs(229)) and not (layer0_outputs(9049));
    outputs(9509) <= not((layer0_outputs(7360)) or (layer0_outputs(11415)));
    outputs(9510) <= not(layer0_outputs(337));
    outputs(9511) <= not((layer0_outputs(8803)) or (layer0_outputs(12793)));
    outputs(9512) <= not(layer0_outputs(8714));
    outputs(9513) <= (layer0_outputs(2777)) or (layer0_outputs(11420));
    outputs(9514) <= (layer0_outputs(3178)) and not (layer0_outputs(6829));
    outputs(9515) <= not(layer0_outputs(3739));
    outputs(9516) <= not(layer0_outputs(11778));
    outputs(9517) <= not((layer0_outputs(12073)) xor (layer0_outputs(2220)));
    outputs(9518) <= layer0_outputs(3239);
    outputs(9519) <= layer0_outputs(2274);
    outputs(9520) <= not((layer0_outputs(8895)) or (layer0_outputs(886)));
    outputs(9521) <= (layer0_outputs(3077)) and not (layer0_outputs(1686));
    outputs(9522) <= not(layer0_outputs(10257));
    outputs(9523) <= not((layer0_outputs(6418)) or (layer0_outputs(4415)));
    outputs(9524) <= (layer0_outputs(11609)) and not (layer0_outputs(9048));
    outputs(9525) <= not(layer0_outputs(2935)) or (layer0_outputs(9523));
    outputs(9526) <= (layer0_outputs(5447)) xor (layer0_outputs(3770));
    outputs(9527) <= layer0_outputs(1973);
    outputs(9528) <= layer0_outputs(7547);
    outputs(9529) <= not((layer0_outputs(8598)) or (layer0_outputs(6618)));
    outputs(9530) <= (layer0_outputs(9658)) or (layer0_outputs(9077));
    outputs(9531) <= (layer0_outputs(8407)) and not (layer0_outputs(8724));
    outputs(9532) <= not(layer0_outputs(8324));
    outputs(9533) <= (layer0_outputs(12276)) and (layer0_outputs(10280));
    outputs(9534) <= not((layer0_outputs(2417)) or (layer0_outputs(1634)));
    outputs(9535) <= (layer0_outputs(7156)) and not (layer0_outputs(8813));
    outputs(9536) <= (layer0_outputs(902)) and (layer0_outputs(12674));
    outputs(9537) <= layer0_outputs(12766);
    outputs(9538) <= layer0_outputs(1722);
    outputs(9539) <= (layer0_outputs(9095)) and not (layer0_outputs(11491));
    outputs(9540) <= not((layer0_outputs(7233)) or (layer0_outputs(8879)));
    outputs(9541) <= (layer0_outputs(2899)) and not (layer0_outputs(12609));
    outputs(9542) <= not(layer0_outputs(2447)) or (layer0_outputs(7755));
    outputs(9543) <= not(layer0_outputs(5559));
    outputs(9544) <= layer0_outputs(4836);
    outputs(9545) <= (layer0_outputs(11797)) and (layer0_outputs(11892));
    outputs(9546) <= layer0_outputs(8698);
    outputs(9547) <= not((layer0_outputs(9541)) xor (layer0_outputs(11794)));
    outputs(9548) <= not(layer0_outputs(1392));
    outputs(9549) <= not(layer0_outputs(11460));
    outputs(9550) <= layer0_outputs(4299);
    outputs(9551) <= not((layer0_outputs(2703)) xor (layer0_outputs(9228)));
    outputs(9552) <= not(layer0_outputs(9627));
    outputs(9553) <= layer0_outputs(8800);
    outputs(9554) <= (layer0_outputs(3680)) and not (layer0_outputs(5868));
    outputs(9555) <= not(layer0_outputs(9039));
    outputs(9556) <= not((layer0_outputs(3819)) and (layer0_outputs(2623)));
    outputs(9557) <= (layer0_outputs(3533)) and not (layer0_outputs(10807));
    outputs(9558) <= not(layer0_outputs(3215));
    outputs(9559) <= not((layer0_outputs(416)) xor (layer0_outputs(12275)));
    outputs(9560) <= not(layer0_outputs(4732));
    outputs(9561) <= not(layer0_outputs(7026));
    outputs(9562) <= not((layer0_outputs(11261)) xor (layer0_outputs(6215)));
    outputs(9563) <= (layer0_outputs(648)) and not (layer0_outputs(9776));
    outputs(9564) <= (layer0_outputs(2196)) and not (layer0_outputs(1716));
    outputs(9565) <= layer0_outputs(1299);
    outputs(9566) <= (layer0_outputs(3850)) xor (layer0_outputs(333));
    outputs(9567) <= (layer0_outputs(9876)) and not (layer0_outputs(7213));
    outputs(9568) <= not(layer0_outputs(10188));
    outputs(9569) <= (layer0_outputs(7348)) and not (layer0_outputs(3484));
    outputs(9570) <= not(layer0_outputs(11249));
    outputs(9571) <= (layer0_outputs(4282)) and (layer0_outputs(4530));
    outputs(9572) <= not(layer0_outputs(9428));
    outputs(9573) <= layer0_outputs(7171);
    outputs(9574) <= not((layer0_outputs(9834)) or (layer0_outputs(12421)));
    outputs(9575) <= (layer0_outputs(895)) and not (layer0_outputs(4029));
    outputs(9576) <= not(layer0_outputs(9115));
    outputs(9577) <= (layer0_outputs(3305)) xor (layer0_outputs(6483));
    outputs(9578) <= not((layer0_outputs(12240)) or (layer0_outputs(4662)));
    outputs(9579) <= (layer0_outputs(5525)) and (layer0_outputs(655));
    outputs(9580) <= not((layer0_outputs(10868)) xor (layer0_outputs(2700)));
    outputs(9581) <= not(layer0_outputs(4370));
    outputs(9582) <= not((layer0_outputs(7344)) xor (layer0_outputs(2380)));
    outputs(9583) <= not(layer0_outputs(8980));
    outputs(9584) <= not(layer0_outputs(5792));
    outputs(9585) <= not((layer0_outputs(11133)) xor (layer0_outputs(2954)));
    outputs(9586) <= layer0_outputs(3629);
    outputs(9587) <= not((layer0_outputs(10994)) xor (layer0_outputs(6399)));
    outputs(9588) <= not(layer0_outputs(990)) or (layer0_outputs(7653));
    outputs(9589) <= not(layer0_outputs(7899));
    outputs(9590) <= layer0_outputs(1012);
    outputs(9591) <= layer0_outputs(8844);
    outputs(9592) <= (layer0_outputs(9942)) and not (layer0_outputs(2839));
    outputs(9593) <= not(layer0_outputs(49));
    outputs(9594) <= (layer0_outputs(10358)) and not (layer0_outputs(4554));
    outputs(9595) <= (layer0_outputs(11796)) and (layer0_outputs(11890));
    outputs(9596) <= not(layer0_outputs(8797));
    outputs(9597) <= not(layer0_outputs(11448));
    outputs(9598) <= not(layer0_outputs(3920));
    outputs(9599) <= layer0_outputs(3463);
    outputs(9600) <= layer0_outputs(1251);
    outputs(9601) <= (layer0_outputs(8568)) xor (layer0_outputs(8593));
    outputs(9602) <= not((layer0_outputs(35)) xor (layer0_outputs(4765)));
    outputs(9603) <= not((layer0_outputs(7607)) or (layer0_outputs(1037)));
    outputs(9604) <= not(layer0_outputs(5760));
    outputs(9605) <= not(layer0_outputs(1860));
    outputs(9606) <= layer0_outputs(2425);
    outputs(9607) <= (layer0_outputs(968)) and (layer0_outputs(1087));
    outputs(9608) <= layer0_outputs(9929);
    outputs(9609) <= not((layer0_outputs(6755)) xor (layer0_outputs(2861)));
    outputs(9610) <= layer0_outputs(7479);
    outputs(9611) <= layer0_outputs(3498);
    outputs(9612) <= layer0_outputs(2744);
    outputs(9613) <= (layer0_outputs(70)) xor (layer0_outputs(4703));
    outputs(9614) <= layer0_outputs(10906);
    outputs(9615) <= layer0_outputs(2819);
    outputs(9616) <= not(layer0_outputs(12614));
    outputs(9617) <= (layer0_outputs(528)) and not (layer0_outputs(2849));
    outputs(9618) <= layer0_outputs(12473);
    outputs(9619) <= not(layer0_outputs(5737));
    outputs(9620) <= not(layer0_outputs(4406));
    outputs(9621) <= not(layer0_outputs(5881)) or (layer0_outputs(4945));
    outputs(9622) <= layer0_outputs(4366);
    outputs(9623) <= layer0_outputs(3469);
    outputs(9624) <= not(layer0_outputs(12600));
    outputs(9625) <= not(layer0_outputs(1982));
    outputs(9626) <= not((layer0_outputs(12025)) xor (layer0_outputs(7442)));
    outputs(9627) <= layer0_outputs(5679);
    outputs(9628) <= (layer0_outputs(7423)) and not (layer0_outputs(12604));
    outputs(9629) <= (layer0_outputs(4074)) and not (layer0_outputs(7779));
    outputs(9630) <= (layer0_outputs(8372)) and (layer0_outputs(1544));
    outputs(9631) <= (layer0_outputs(5969)) and not (layer0_outputs(6085));
    outputs(9632) <= (layer0_outputs(3189)) xor (layer0_outputs(620));
    outputs(9633) <= (layer0_outputs(6204)) and not (layer0_outputs(10500));
    outputs(9634) <= layer0_outputs(10572);
    outputs(9635) <= not(layer0_outputs(1967));
    outputs(9636) <= layer0_outputs(10212);
    outputs(9637) <= layer0_outputs(5006);
    outputs(9638) <= not(layer0_outputs(8678));
    outputs(9639) <= (layer0_outputs(9429)) and not (layer0_outputs(11292));
    outputs(9640) <= (layer0_outputs(7726)) or (layer0_outputs(7476));
    outputs(9641) <= not((layer0_outputs(12109)) and (layer0_outputs(12336)));
    outputs(9642) <= not((layer0_outputs(7640)) or (layer0_outputs(11470)));
    outputs(9643) <= (layer0_outputs(12762)) xor (layer0_outputs(9319));
    outputs(9644) <= layer0_outputs(2716);
    outputs(9645) <= not(layer0_outputs(1912));
    outputs(9646) <= (layer0_outputs(7761)) and not (layer0_outputs(1525));
    outputs(9647) <= (layer0_outputs(3287)) xor (layer0_outputs(1631));
    outputs(9648) <= layer0_outputs(11020);
    outputs(9649) <= layer0_outputs(8318);
    outputs(9650) <= not(layer0_outputs(11954));
    outputs(9651) <= layer0_outputs(5492);
    outputs(9652) <= not(layer0_outputs(2723));
    outputs(9653) <= (layer0_outputs(1239)) and not (layer0_outputs(11140));
    outputs(9654) <= not((layer0_outputs(10675)) or (layer0_outputs(2269)));
    outputs(9655) <= (layer0_outputs(11423)) and (layer0_outputs(9003));
    outputs(9656) <= (layer0_outputs(7777)) and (layer0_outputs(10199));
    outputs(9657) <= not(layer0_outputs(6689)) or (layer0_outputs(12506));
    outputs(9658) <= layer0_outputs(2154);
    outputs(9659) <= not(layer0_outputs(7273));
    outputs(9660) <= not(layer0_outputs(10840));
    outputs(9661) <= (layer0_outputs(5365)) xor (layer0_outputs(9205));
    outputs(9662) <= not((layer0_outputs(8354)) xor (layer0_outputs(12375)));
    outputs(9663) <= not(layer0_outputs(179));
    outputs(9664) <= layer0_outputs(3051);
    outputs(9665) <= layer0_outputs(5583);
    outputs(9666) <= (layer0_outputs(1061)) and not (layer0_outputs(10465));
    outputs(9667) <= layer0_outputs(4346);
    outputs(9668) <= not(layer0_outputs(4627));
    outputs(9669) <= not((layer0_outputs(10838)) or (layer0_outputs(1431)));
    outputs(9670) <= (layer0_outputs(8085)) xor (layer0_outputs(5226));
    outputs(9671) <= (layer0_outputs(10890)) and not (layer0_outputs(1996));
    outputs(9672) <= layer0_outputs(6097);
    outputs(9673) <= not((layer0_outputs(4642)) or (layer0_outputs(9224)));
    outputs(9674) <= (layer0_outputs(8257)) or (layer0_outputs(2932));
    outputs(9675) <= not(layer0_outputs(11331));
    outputs(9676) <= not(layer0_outputs(7121));
    outputs(9677) <= (layer0_outputs(6291)) xor (layer0_outputs(976));
    outputs(9678) <= (layer0_outputs(11468)) and not (layer0_outputs(2804));
    outputs(9679) <= layer0_outputs(3418);
    outputs(9680) <= (layer0_outputs(366)) xor (layer0_outputs(1810));
    outputs(9681) <= not(layer0_outputs(11289));
    outputs(9682) <= (layer0_outputs(6432)) and (layer0_outputs(11715));
    outputs(9683) <= layer0_outputs(3687);
    outputs(9684) <= (layer0_outputs(8713)) and not (layer0_outputs(7727));
    outputs(9685) <= (layer0_outputs(9376)) xor (layer0_outputs(582));
    outputs(9686) <= (layer0_outputs(3840)) and (layer0_outputs(4319));
    outputs(9687) <= not((layer0_outputs(10702)) xor (layer0_outputs(3877)));
    outputs(9688) <= (layer0_outputs(5833)) or (layer0_outputs(8828));
    outputs(9689) <= not(layer0_outputs(3756));
    outputs(9690) <= layer0_outputs(6123);
    outputs(9691) <= not((layer0_outputs(8838)) and (layer0_outputs(11171)));
    outputs(9692) <= not((layer0_outputs(4590)) xor (layer0_outputs(2805)));
    outputs(9693) <= (layer0_outputs(10677)) and not (layer0_outputs(6787));
    outputs(9694) <= (layer0_outputs(11631)) xor (layer0_outputs(9257));
    outputs(9695) <= not((layer0_outputs(6714)) and (layer0_outputs(8137)));
    outputs(9696) <= layer0_outputs(12795);
    outputs(9697) <= layer0_outputs(409);
    outputs(9698) <= (layer0_outputs(5370)) and (layer0_outputs(1979));
    outputs(9699) <= layer0_outputs(1177);
    outputs(9700) <= not(layer0_outputs(10538));
    outputs(9701) <= layer0_outputs(11855);
    outputs(9702) <= not((layer0_outputs(8311)) or (layer0_outputs(4623)));
    outputs(9703) <= not(layer0_outputs(12178));
    outputs(9704) <= (layer0_outputs(1577)) or (layer0_outputs(3502));
    outputs(9705) <= not(layer0_outputs(10174));
    outputs(9706) <= not(layer0_outputs(1976)) or (layer0_outputs(10986));
    outputs(9707) <= not(layer0_outputs(4437));
    outputs(9708) <= not((layer0_outputs(2967)) xor (layer0_outputs(5201)));
    outputs(9709) <= not((layer0_outputs(958)) or (layer0_outputs(10461)));
    outputs(9710) <= not(layer0_outputs(8414));
    outputs(9711) <= (layer0_outputs(11352)) and (layer0_outputs(5973));
    outputs(9712) <= not((layer0_outputs(11736)) and (layer0_outputs(4371)));
    outputs(9713) <= layer0_outputs(5496);
    outputs(9714) <= not(layer0_outputs(11840));
    outputs(9715) <= not(layer0_outputs(10131));
    outputs(9716) <= (layer0_outputs(6076)) and (layer0_outputs(5960));
    outputs(9717) <= layer0_outputs(3635);
    outputs(9718) <= not((layer0_outputs(2705)) xor (layer0_outputs(2636)));
    outputs(9719) <= (layer0_outputs(3231)) xor (layer0_outputs(257));
    outputs(9720) <= (layer0_outputs(113)) xor (layer0_outputs(8915));
    outputs(9721) <= not(layer0_outputs(8882));
    outputs(9722) <= (layer0_outputs(9325)) and (layer0_outputs(12668));
    outputs(9723) <= layer0_outputs(2356);
    outputs(9724) <= (layer0_outputs(9118)) xor (layer0_outputs(11501));
    outputs(9725) <= not(layer0_outputs(9018));
    outputs(9726) <= (layer0_outputs(1652)) xor (layer0_outputs(2712));
    outputs(9727) <= not(layer0_outputs(7910));
    outputs(9728) <= layer0_outputs(1235);
    outputs(9729) <= not((layer0_outputs(8010)) xor (layer0_outputs(4552)));
    outputs(9730) <= not(layer0_outputs(9933));
    outputs(9731) <= layer0_outputs(8863);
    outputs(9732) <= not(layer0_outputs(1028));
    outputs(9733) <= not(layer0_outputs(6758));
    outputs(9734) <= (layer0_outputs(6940)) and (layer0_outputs(3897));
    outputs(9735) <= not((layer0_outputs(8634)) xor (layer0_outputs(4837)));
    outputs(9736) <= not((layer0_outputs(11464)) xor (layer0_outputs(8512)));
    outputs(9737) <= not((layer0_outputs(7169)) or (layer0_outputs(5257)));
    outputs(9738) <= (layer0_outputs(5928)) and not (layer0_outputs(10771));
    outputs(9739) <= (layer0_outputs(6206)) xor (layer0_outputs(5140));
    outputs(9740) <= not((layer0_outputs(4077)) xor (layer0_outputs(10059)));
    outputs(9741) <= not((layer0_outputs(4507)) or (layer0_outputs(8442)));
    outputs(9742) <= layer0_outputs(12709);
    outputs(9743) <= not(layer0_outputs(308));
    outputs(9744) <= not((layer0_outputs(8554)) and (layer0_outputs(8274)));
    outputs(9745) <= not(layer0_outputs(12105));
    outputs(9746) <= not(layer0_outputs(7762));
    outputs(9747) <= (layer0_outputs(6672)) and (layer0_outputs(2654));
    outputs(9748) <= not((layer0_outputs(8766)) or (layer0_outputs(8735)));
    outputs(9749) <= (layer0_outputs(4635)) and not (layer0_outputs(2843));
    outputs(9750) <= not(layer0_outputs(2189));
    outputs(9751) <= layer0_outputs(4335);
    outputs(9752) <= not(layer0_outputs(10476));
    outputs(9753) <= not(layer0_outputs(12590));
    outputs(9754) <= (layer0_outputs(8623)) xor (layer0_outputs(11451));
    outputs(9755) <= (layer0_outputs(11147)) xor (layer0_outputs(5801));
    outputs(9756) <= not(layer0_outputs(8451)) or (layer0_outputs(2258));
    outputs(9757) <= (layer0_outputs(5011)) and not (layer0_outputs(1848));
    outputs(9758) <= not(layer0_outputs(6907));
    outputs(9759) <= (layer0_outputs(5648)) and (layer0_outputs(10392));
    outputs(9760) <= not(layer0_outputs(9004));
    outputs(9761) <= not((layer0_outputs(5805)) or (layer0_outputs(6490)));
    outputs(9762) <= not(layer0_outputs(7688));
    outputs(9763) <= layer0_outputs(1387);
    outputs(9764) <= not(layer0_outputs(6100));
    outputs(9765) <= not(layer0_outputs(12446));
    outputs(9766) <= (layer0_outputs(8570)) and not (layer0_outputs(4284));
    outputs(9767) <= not((layer0_outputs(8597)) or (layer0_outputs(62)));
    outputs(9768) <= (layer0_outputs(7949)) and not (layer0_outputs(9185));
    outputs(9769) <= not(layer0_outputs(11027));
    outputs(9770) <= not(layer0_outputs(9561)) or (layer0_outputs(12430));
    outputs(9771) <= (layer0_outputs(2083)) and not (layer0_outputs(517));
    outputs(9772) <= not(layer0_outputs(9792));
    outputs(9773) <= not(layer0_outputs(6933));
    outputs(9774) <= not(layer0_outputs(6872));
    outputs(9775) <= (layer0_outputs(3242)) and not (layer0_outputs(7803));
    outputs(9776) <= (layer0_outputs(2954)) xor (layer0_outputs(8653));
    outputs(9777) <= layer0_outputs(457);
    outputs(9778) <= (layer0_outputs(6329)) xor (layer0_outputs(4675));
    outputs(9779) <= (layer0_outputs(65)) xor (layer0_outputs(10390));
    outputs(9780) <= not((layer0_outputs(2238)) or (layer0_outputs(1480)));
    outputs(9781) <= not((layer0_outputs(2906)) xor (layer0_outputs(4054)));
    outputs(9782) <= layer0_outputs(10479);
    outputs(9783) <= not(layer0_outputs(11244));
    outputs(9784) <= not(layer0_outputs(11228));
    outputs(9785) <= not(layer0_outputs(10454));
    outputs(9786) <= (layer0_outputs(9833)) or (layer0_outputs(12785));
    outputs(9787) <= not(layer0_outputs(11053));
    outputs(9788) <= layer0_outputs(12728);
    outputs(9789) <= (layer0_outputs(9660)) and (layer0_outputs(1360));
    outputs(9790) <= (layer0_outputs(4420)) and not (layer0_outputs(6569));
    outputs(9791) <= not(layer0_outputs(3068));
    outputs(9792) <= not((layer0_outputs(3783)) or (layer0_outputs(9846)));
    outputs(9793) <= not((layer0_outputs(863)) or (layer0_outputs(6200)));
    outputs(9794) <= (layer0_outputs(2716)) or (layer0_outputs(10721));
    outputs(9795) <= not(layer0_outputs(10723)) or (layer0_outputs(10920));
    outputs(9796) <= layer0_outputs(7147);
    outputs(9797) <= not(layer0_outputs(739));
    outputs(9798) <= not((layer0_outputs(108)) xor (layer0_outputs(10897)));
    outputs(9799) <= (layer0_outputs(9557)) and not (layer0_outputs(10632));
    outputs(9800) <= layer0_outputs(4698);
    outputs(9801) <= (layer0_outputs(843)) xor (layer0_outputs(6243));
    outputs(9802) <= not(layer0_outputs(2862));
    outputs(9803) <= not(layer0_outputs(7307));
    outputs(9804) <= (layer0_outputs(4141)) and (layer0_outputs(12199));
    outputs(9805) <= not((layer0_outputs(2031)) or (layer0_outputs(4992)));
    outputs(9806) <= layer0_outputs(9803);
    outputs(9807) <= (layer0_outputs(3000)) and not (layer0_outputs(7141));
    outputs(9808) <= (layer0_outputs(7532)) xor (layer0_outputs(4596));
    outputs(9809) <= layer0_outputs(9992);
    outputs(9810) <= not((layer0_outputs(11413)) xor (layer0_outputs(7842)));
    outputs(9811) <= (layer0_outputs(5673)) xor (layer0_outputs(10812));
    outputs(9812) <= not(layer0_outputs(12685)) or (layer0_outputs(10494));
    outputs(9813) <= not((layer0_outputs(4535)) and (layer0_outputs(5716)));
    outputs(9814) <= not(layer0_outputs(56));
    outputs(9815) <= not(layer0_outputs(11686)) or (layer0_outputs(889));
    outputs(9816) <= layer0_outputs(10860);
    outputs(9817) <= not((layer0_outputs(12169)) or (layer0_outputs(10213)));
    outputs(9818) <= not(layer0_outputs(7926)) or (layer0_outputs(714));
    outputs(9819) <= (layer0_outputs(12149)) or (layer0_outputs(4634));
    outputs(9820) <= not((layer0_outputs(4916)) or (layer0_outputs(6221)));
    outputs(9821) <= (layer0_outputs(2664)) and (layer0_outputs(2552));
    outputs(9822) <= not(layer0_outputs(8884));
    outputs(9823) <= layer0_outputs(8097);
    outputs(9824) <= not((layer0_outputs(2600)) or (layer0_outputs(4362)));
    outputs(9825) <= layer0_outputs(7150);
    outputs(9826) <= not(layer0_outputs(763));
    outputs(9827) <= (layer0_outputs(8832)) and not (layer0_outputs(4285));
    outputs(9828) <= (layer0_outputs(4352)) xor (layer0_outputs(3757));
    outputs(9829) <= layer0_outputs(4245);
    outputs(9830) <= not((layer0_outputs(7256)) or (layer0_outputs(1274)));
    outputs(9831) <= not((layer0_outputs(34)) xor (layer0_outputs(88)));
    outputs(9832) <= not(layer0_outputs(12489));
    outputs(9833) <= (layer0_outputs(11591)) and not (layer0_outputs(4348));
    outputs(9834) <= layer0_outputs(6127);
    outputs(9835) <= layer0_outputs(6320);
    outputs(9836) <= (layer0_outputs(5846)) and (layer0_outputs(4654));
    outputs(9837) <= not((layer0_outputs(12485)) xor (layer0_outputs(6351)));
    outputs(9838) <= not((layer0_outputs(8410)) or (layer0_outputs(12404)));
    outputs(9839) <= not((layer0_outputs(3338)) xor (layer0_outputs(1252)));
    outputs(9840) <= (layer0_outputs(6145)) and (layer0_outputs(4585));
    outputs(9841) <= not(layer0_outputs(3190));
    outputs(9842) <= layer0_outputs(6961);
    outputs(9843) <= (layer0_outputs(5355)) and not (layer0_outputs(11728));
    outputs(9844) <= not((layer0_outputs(8013)) xor (layer0_outputs(8191)));
    outputs(9845) <= layer0_outputs(8290);
    outputs(9846) <= (layer0_outputs(10111)) and not (layer0_outputs(10514));
    outputs(9847) <= layer0_outputs(970);
    outputs(9848) <= (layer0_outputs(9863)) xor (layer0_outputs(6718));
    outputs(9849) <= (layer0_outputs(275)) and not (layer0_outputs(12225));
    outputs(9850) <= not((layer0_outputs(11852)) xor (layer0_outputs(7511)));
    outputs(9851) <= (layer0_outputs(5057)) and (layer0_outputs(10606));
    outputs(9852) <= layer0_outputs(11893);
    outputs(9853) <= not((layer0_outputs(12336)) and (layer0_outputs(6536)));
    outputs(9854) <= not(layer0_outputs(8960)) or (layer0_outputs(1575));
    outputs(9855) <= (layer0_outputs(5248)) and (layer0_outputs(7454));
    outputs(9856) <= not((layer0_outputs(7320)) xor (layer0_outputs(3754)));
    outputs(9857) <= not(layer0_outputs(3882)) or (layer0_outputs(2923));
    outputs(9858) <= (layer0_outputs(11173)) xor (layer0_outputs(8047));
    outputs(9859) <= not(layer0_outputs(11951));
    outputs(9860) <= (layer0_outputs(1936)) and (layer0_outputs(5272));
    outputs(9861) <= layer0_outputs(2825);
    outputs(9862) <= not(layer0_outputs(2351));
    outputs(9863) <= (layer0_outputs(4648)) xor (layer0_outputs(7656));
    outputs(9864) <= (layer0_outputs(7477)) and not (layer0_outputs(1366));
    outputs(9865) <= not(layer0_outputs(8793));
    outputs(9866) <= not(layer0_outputs(5400));
    outputs(9867) <= (layer0_outputs(4022)) and not (layer0_outputs(5394));
    outputs(9868) <= not(layer0_outputs(5228));
    outputs(9869) <= not((layer0_outputs(8899)) xor (layer0_outputs(5491)));
    outputs(9870) <= not((layer0_outputs(4301)) and (layer0_outputs(6716)));
    outputs(9871) <= not(layer0_outputs(7830));
    outputs(9872) <= layer0_outputs(3434);
    outputs(9873) <= (layer0_outputs(6541)) xor (layer0_outputs(10094));
    outputs(9874) <= not((layer0_outputs(5902)) xor (layer0_outputs(4376)));
    outputs(9875) <= layer0_outputs(205);
    outputs(9876) <= not(layer0_outputs(961));
    outputs(9877) <= not(layer0_outputs(8445));
    outputs(9878) <= layer0_outputs(2679);
    outputs(9879) <= (layer0_outputs(8486)) and not (layer0_outputs(9128));
    outputs(9880) <= layer0_outputs(2985);
    outputs(9881) <= not(layer0_outputs(8652));
    outputs(9882) <= layer0_outputs(3414);
    outputs(9883) <= not(layer0_outputs(12178));
    outputs(9884) <= not(layer0_outputs(7174));
    outputs(9885) <= layer0_outputs(9800);
    outputs(9886) <= (layer0_outputs(1062)) and not (layer0_outputs(403));
    outputs(9887) <= not(layer0_outputs(11044));
    outputs(9888) <= layer0_outputs(2830);
    outputs(9889) <= (layer0_outputs(8918)) xor (layer0_outputs(3763));
    outputs(9890) <= (layer0_outputs(4085)) or (layer0_outputs(10346));
    outputs(9891) <= not(layer0_outputs(7404)) or (layer0_outputs(6896));
    outputs(9892) <= not(layer0_outputs(12087));
    outputs(9893) <= not(layer0_outputs(4218));
    outputs(9894) <= layer0_outputs(4236);
    outputs(9895) <= not(layer0_outputs(2060));
    outputs(9896) <= (layer0_outputs(8452)) and (layer0_outputs(949));
    outputs(9897) <= (layer0_outputs(8396)) and not (layer0_outputs(11337));
    outputs(9898) <= layer0_outputs(10267);
    outputs(9899) <= (layer0_outputs(6783)) and not (layer0_outputs(2184));
    outputs(9900) <= layer0_outputs(8844);
    outputs(9901) <= not(layer0_outputs(4576));
    outputs(9902) <= not(layer0_outputs(2801));
    outputs(9903) <= not(layer0_outputs(586));
    outputs(9904) <= (layer0_outputs(9491)) xor (layer0_outputs(6911));
    outputs(9905) <= (layer0_outputs(7734)) and not (layer0_outputs(12646));
    outputs(9906) <= not((layer0_outputs(7784)) or (layer0_outputs(11211)));
    outputs(9907) <= layer0_outputs(10323);
    outputs(9908) <= (layer0_outputs(2296)) and not (layer0_outputs(3381));
    outputs(9909) <= not(layer0_outputs(1842)) or (layer0_outputs(10666));
    outputs(9910) <= (layer0_outputs(5330)) and (layer0_outputs(39));
    outputs(9911) <= layer0_outputs(5330);
    outputs(9912) <= layer0_outputs(3749);
    outputs(9913) <= not((layer0_outputs(1015)) xor (layer0_outputs(3113)));
    outputs(9914) <= (layer0_outputs(9179)) xor (layer0_outputs(1006));
    outputs(9915) <= layer0_outputs(3960);
    outputs(9916) <= layer0_outputs(4764);
    outputs(9917) <= not(layer0_outputs(904)) or (layer0_outputs(9323));
    outputs(9918) <= not((layer0_outputs(8439)) xor (layer0_outputs(8120)));
    outputs(9919) <= not(layer0_outputs(1026));
    outputs(9920) <= (layer0_outputs(47)) or (layer0_outputs(192));
    outputs(9921) <= not((layer0_outputs(9334)) xor (layer0_outputs(2737)));
    outputs(9922) <= not((layer0_outputs(12442)) xor (layer0_outputs(772)));
    outputs(9923) <= not((layer0_outputs(8227)) xor (layer0_outputs(8401)));
    outputs(9924) <= not(layer0_outputs(4910));
    outputs(9925) <= (layer0_outputs(6419)) and not (layer0_outputs(12708));
    outputs(9926) <= not(layer0_outputs(5580));
    outputs(9927) <= (layer0_outputs(1414)) xor (layer0_outputs(10495));
    outputs(9928) <= layer0_outputs(7294);
    outputs(9929) <= layer0_outputs(5931);
    outputs(9930) <= layer0_outputs(10571);
    outputs(9931) <= (layer0_outputs(10993)) and not (layer0_outputs(7264));
    outputs(9932) <= layer0_outputs(9179);
    outputs(9933) <= not((layer0_outputs(3113)) xor (layer0_outputs(5723)));
    outputs(9934) <= not((layer0_outputs(2729)) xor (layer0_outputs(6955)));
    outputs(9935) <= not(layer0_outputs(884));
    outputs(9936) <= not(layer0_outputs(8533));
    outputs(9937) <= (layer0_outputs(12136)) and (layer0_outputs(8047));
    outputs(9938) <= not((layer0_outputs(4298)) xor (layer0_outputs(3476)));
    outputs(9939) <= layer0_outputs(9831);
    outputs(9940) <= (layer0_outputs(12033)) xor (layer0_outputs(5916));
    outputs(9941) <= not((layer0_outputs(3682)) xor (layer0_outputs(5871)));
    outputs(9942) <= (layer0_outputs(8903)) and not (layer0_outputs(6069));
    outputs(9943) <= (layer0_outputs(7359)) and not (layer0_outputs(9045));
    outputs(9944) <= (layer0_outputs(4797)) or (layer0_outputs(210));
    outputs(9945) <= (layer0_outputs(7269)) or (layer0_outputs(9785));
    outputs(9946) <= layer0_outputs(3695);
    outputs(9947) <= not(layer0_outputs(4180));
    outputs(9948) <= (layer0_outputs(3101)) xor (layer0_outputs(1100));
    outputs(9949) <= layer0_outputs(8627);
    outputs(9950) <= not((layer0_outputs(5265)) xor (layer0_outputs(1732)));
    outputs(9951) <= (layer0_outputs(8063)) and (layer0_outputs(2260));
    outputs(9952) <= layer0_outputs(10615);
    outputs(9953) <= layer0_outputs(12060);
    outputs(9954) <= not(layer0_outputs(5399));
    outputs(9955) <= not(layer0_outputs(1572));
    outputs(9956) <= not(layer0_outputs(5460));
    outputs(9957) <= not(layer0_outputs(308));
    outputs(9958) <= (layer0_outputs(11830)) and not (layer0_outputs(1591));
    outputs(9959) <= not(layer0_outputs(5701));
    outputs(9960) <= not(layer0_outputs(6763));
    outputs(9961) <= layer0_outputs(5291);
    outputs(9962) <= (layer0_outputs(12537)) and not (layer0_outputs(10913));
    outputs(9963) <= layer0_outputs(5035);
    outputs(9964) <= layer0_outputs(12473);
    outputs(9965) <= not(layer0_outputs(3977));
    outputs(9966) <= not(layer0_outputs(11296));
    outputs(9967) <= not(layer0_outputs(7743));
    outputs(9968) <= not(layer0_outputs(2435));
    outputs(9969) <= (layer0_outputs(1040)) and (layer0_outputs(3815));
    outputs(9970) <= not(layer0_outputs(2455));
    outputs(9971) <= layer0_outputs(6035);
    outputs(9972) <= layer0_outputs(164);
    outputs(9973) <= (layer0_outputs(7042)) xor (layer0_outputs(87));
    outputs(9974) <= not((layer0_outputs(794)) or (layer0_outputs(6546)));
    outputs(9975) <= (layer0_outputs(6825)) xor (layer0_outputs(8812));
    outputs(9976) <= not(layer0_outputs(1598));
    outputs(9977) <= not(layer0_outputs(1348));
    outputs(9978) <= (layer0_outputs(4193)) and (layer0_outputs(9391));
    outputs(9979) <= not(layer0_outputs(387)) or (layer0_outputs(4551));
    outputs(9980) <= not((layer0_outputs(4314)) or (layer0_outputs(1203)));
    outputs(9981) <= (layer0_outputs(2258)) and (layer0_outputs(2683));
    outputs(9982) <= not((layer0_outputs(11498)) xor (layer0_outputs(11295)));
    outputs(9983) <= not((layer0_outputs(6946)) or (layer0_outputs(1796)));
    outputs(9984) <= not(layer0_outputs(7041));
    outputs(9985) <= layer0_outputs(6260);
    outputs(9986) <= not((layer0_outputs(4579)) xor (layer0_outputs(3644)));
    outputs(9987) <= layer0_outputs(638);
    outputs(9988) <= layer0_outputs(12393);
    outputs(9989) <= not((layer0_outputs(11861)) xor (layer0_outputs(9134)));
    outputs(9990) <= (layer0_outputs(9963)) and (layer0_outputs(1827));
    outputs(9991) <= layer0_outputs(8513);
    outputs(9992) <= (layer0_outputs(2380)) and (layer0_outputs(7690));
    outputs(9993) <= (layer0_outputs(12476)) and (layer0_outputs(5246));
    outputs(9994) <= not(layer0_outputs(4258));
    outputs(9995) <= (layer0_outputs(8933)) and not (layer0_outputs(3538));
    outputs(9996) <= layer0_outputs(11412);
    outputs(9997) <= layer0_outputs(7258);
    outputs(9998) <= not(layer0_outputs(2211));
    outputs(9999) <= not((layer0_outputs(897)) or (layer0_outputs(12406)));
    outputs(10000) <= not(layer0_outputs(12508));
    outputs(10001) <= not(layer0_outputs(4424));
    outputs(10002) <= (layer0_outputs(8636)) and (layer0_outputs(11647));
    outputs(10003) <= not((layer0_outputs(7596)) or (layer0_outputs(4905)));
    outputs(10004) <= (layer0_outputs(3104)) or (layer0_outputs(7756));
    outputs(10005) <= layer0_outputs(6609);
    outputs(10006) <= not(layer0_outputs(2035));
    outputs(10007) <= (layer0_outputs(8643)) and (layer0_outputs(1270));
    outputs(10008) <= not(layer0_outputs(12116));
    outputs(10009) <= (layer0_outputs(11060)) and not (layer0_outputs(6775));
    outputs(10010) <= layer0_outputs(5167);
    outputs(10011) <= (layer0_outputs(2722)) and not (layer0_outputs(12361));
    outputs(10012) <= not(layer0_outputs(6155));
    outputs(10013) <= not(layer0_outputs(1485));
    outputs(10014) <= not(layer0_outputs(12001));
    outputs(10015) <= layer0_outputs(12145);
    outputs(10016) <= layer0_outputs(2832);
    outputs(10017) <= not(layer0_outputs(8937));
    outputs(10018) <= not(layer0_outputs(9933));
    outputs(10019) <= not(layer0_outputs(1751));
    outputs(10020) <= (layer0_outputs(10155)) and (layer0_outputs(12266));
    outputs(10021) <= layer0_outputs(2501);
    outputs(10022) <= (layer0_outputs(2440)) and not (layer0_outputs(7793));
    outputs(10023) <= layer0_outputs(7499);
    outputs(10024) <= (layer0_outputs(12485)) xor (layer0_outputs(3267));
    outputs(10025) <= not(layer0_outputs(3260));
    outputs(10026) <= layer0_outputs(7308);
    outputs(10027) <= (layer0_outputs(11428)) and (layer0_outputs(9442));
    outputs(10028) <= not(layer0_outputs(2490)) or (layer0_outputs(9514));
    outputs(10029) <= layer0_outputs(4097);
    outputs(10030) <= (layer0_outputs(11476)) xor (layer0_outputs(9061));
    outputs(10031) <= not(layer0_outputs(2200));
    outputs(10032) <= (layer0_outputs(1648)) and (layer0_outputs(524));
    outputs(10033) <= not(layer0_outputs(292));
    outputs(10034) <= layer0_outputs(8245);
    outputs(10035) <= layer0_outputs(10931);
    outputs(10036) <= not(layer0_outputs(12520));
    outputs(10037) <= (layer0_outputs(10408)) xor (layer0_outputs(9753));
    outputs(10038) <= (layer0_outputs(12694)) xor (layer0_outputs(3666));
    outputs(10039) <= (layer0_outputs(7335)) xor (layer0_outputs(7391));
    outputs(10040) <= not(layer0_outputs(6518));
    outputs(10041) <= (layer0_outputs(4677)) and not (layer0_outputs(8983));
    outputs(10042) <= (layer0_outputs(7831)) and (layer0_outputs(1621));
    outputs(10043) <= not((layer0_outputs(4148)) xor (layer0_outputs(5612)));
    outputs(10044) <= (layer0_outputs(8717)) and not (layer0_outputs(8476));
    outputs(10045) <= not(layer0_outputs(3708)) or (layer0_outputs(2370));
    outputs(10046) <= layer0_outputs(12078);
    outputs(10047) <= (layer0_outputs(8416)) and not (layer0_outputs(4699));
    outputs(10048) <= not(layer0_outputs(9143)) or (layer0_outputs(352));
    outputs(10049) <= (layer0_outputs(733)) and (layer0_outputs(6329));
    outputs(10050) <= (layer0_outputs(1214)) and not (layer0_outputs(6796));
    outputs(10051) <= layer0_outputs(1376);
    outputs(10052) <= (layer0_outputs(2851)) or (layer0_outputs(3275));
    outputs(10053) <= (layer0_outputs(8058)) and not (layer0_outputs(3659));
    outputs(10054) <= layer0_outputs(1239);
    outputs(10055) <= (layer0_outputs(9170)) and (layer0_outputs(12171));
    outputs(10056) <= (layer0_outputs(3699)) and not (layer0_outputs(9853));
    outputs(10057) <= (layer0_outputs(9674)) and not (layer0_outputs(1466));
    outputs(10058) <= (layer0_outputs(12632)) and (layer0_outputs(461));
    outputs(10059) <= not((layer0_outputs(5331)) xor (layer0_outputs(952)));
    outputs(10060) <= not((layer0_outputs(4905)) or (layer0_outputs(12461)));
    outputs(10061) <= layer0_outputs(10657);
    outputs(10062) <= not(layer0_outputs(7772));
    outputs(10063) <= not((layer0_outputs(10623)) or (layer0_outputs(12316)));
    outputs(10064) <= layer0_outputs(6446);
    outputs(10065) <= (layer0_outputs(7183)) and not (layer0_outputs(1248));
    outputs(10066) <= not((layer0_outputs(10943)) xor (layer0_outputs(483)));
    outputs(10067) <= layer0_outputs(6431);
    outputs(10068) <= (layer0_outputs(10270)) and not (layer0_outputs(11932));
    outputs(10069) <= layer0_outputs(9243);
    outputs(10070) <= not(layer0_outputs(8137));
    outputs(10071) <= layer0_outputs(3431);
    outputs(10072) <= layer0_outputs(9384);
    outputs(10073) <= (layer0_outputs(9498)) and not (layer0_outputs(5898));
    outputs(10074) <= (layer0_outputs(8099)) xor (layer0_outputs(4173));
    outputs(10075) <= not(layer0_outputs(11171));
    outputs(10076) <= layer0_outputs(4489);
    outputs(10077) <= not(layer0_outputs(9037));
    outputs(10078) <= not(layer0_outputs(11507));
    outputs(10079) <= not(layer0_outputs(8966));
    outputs(10080) <= not(layer0_outputs(8342));
    outputs(10081) <= not((layer0_outputs(1127)) or (layer0_outputs(9778)));
    outputs(10082) <= (layer0_outputs(5712)) and not (layer0_outputs(5678));
    outputs(10083) <= not(layer0_outputs(2147));
    outputs(10084) <= layer0_outputs(11767);
    outputs(10085) <= (layer0_outputs(1434)) xor (layer0_outputs(6163));
    outputs(10086) <= layer0_outputs(9245);
    outputs(10087) <= not(layer0_outputs(4667)) or (layer0_outputs(9084));
    outputs(10088) <= not(layer0_outputs(4795));
    outputs(10089) <= (layer0_outputs(1562)) or (layer0_outputs(6264));
    outputs(10090) <= (layer0_outputs(8265)) and not (layer0_outputs(4815));
    outputs(10091) <= (layer0_outputs(3326)) and not (layer0_outputs(11288));
    outputs(10092) <= not(layer0_outputs(7013));
    outputs(10093) <= not((layer0_outputs(4775)) xor (layer0_outputs(6370)));
    outputs(10094) <= layer0_outputs(9133);
    outputs(10095) <= layer0_outputs(10200);
    outputs(10096) <= not(layer0_outputs(4969));
    outputs(10097) <= not(layer0_outputs(6295)) or (layer0_outputs(7895));
    outputs(10098) <= layer0_outputs(3075);
    outputs(10099) <= layer0_outputs(11398);
    outputs(10100) <= layer0_outputs(6384);
    outputs(10101) <= not(layer0_outputs(8322));
    outputs(10102) <= not(layer0_outputs(7962));
    outputs(10103) <= not(layer0_outputs(11826));
    outputs(10104) <= layer0_outputs(3698);
    outputs(10105) <= not(layer0_outputs(2891));
    outputs(10106) <= (layer0_outputs(8335)) or (layer0_outputs(1789));
    outputs(10107) <= layer0_outputs(7073);
    outputs(10108) <= layer0_outputs(7135);
    outputs(10109) <= layer0_outputs(6585);
    outputs(10110) <= (layer0_outputs(574)) xor (layer0_outputs(10852));
    outputs(10111) <= (layer0_outputs(2454)) and not (layer0_outputs(9788));
    outputs(10112) <= not((layer0_outputs(11277)) or (layer0_outputs(3538)));
    outputs(10113) <= layer0_outputs(3628);
    outputs(10114) <= not(layer0_outputs(9736));
    outputs(10115) <= (layer0_outputs(8971)) and not (layer0_outputs(2371));
    outputs(10116) <= not((layer0_outputs(8439)) xor (layer0_outputs(3449)));
    outputs(10117) <= layer0_outputs(2982);
    outputs(10118) <= not(layer0_outputs(4717));
    outputs(10119) <= layer0_outputs(10130);
    outputs(10120) <= (layer0_outputs(362)) and not (layer0_outputs(11071));
    outputs(10121) <= not(layer0_outputs(4174));
    outputs(10122) <= layer0_outputs(8666);
    outputs(10123) <= not(layer0_outputs(4568));
    outputs(10124) <= not(layer0_outputs(12015)) or (layer0_outputs(8155));
    outputs(10125) <= not(layer0_outputs(11832));
    outputs(10126) <= not((layer0_outputs(279)) and (layer0_outputs(7420)));
    outputs(10127) <= (layer0_outputs(1296)) and not (layer0_outputs(2325));
    outputs(10128) <= (layer0_outputs(1350)) and (layer0_outputs(12611));
    outputs(10129) <= not(layer0_outputs(11158));
    outputs(10130) <= not(layer0_outputs(9217));
    outputs(10131) <= (layer0_outputs(2105)) xor (layer0_outputs(3081));
    outputs(10132) <= layer0_outputs(2774);
    outputs(10133) <= not((layer0_outputs(10299)) xor (layer0_outputs(2504)));
    outputs(10134) <= (layer0_outputs(5880)) xor (layer0_outputs(1680));
    outputs(10135) <= not(layer0_outputs(3407)) or (layer0_outputs(4760));
    outputs(10136) <= (layer0_outputs(1991)) and (layer0_outputs(11913));
    outputs(10137) <= not(layer0_outputs(4852));
    outputs(10138) <= not(layer0_outputs(4263));
    outputs(10139) <= not(layer0_outputs(9525));
    outputs(10140) <= not((layer0_outputs(12653)) or (layer0_outputs(10271)));
    outputs(10141) <= not(layer0_outputs(5835));
    outputs(10142) <= layer0_outputs(3277);
    outputs(10143) <= layer0_outputs(4889);
    outputs(10144) <= not(layer0_outputs(4040));
    outputs(10145) <= layer0_outputs(10787);
    outputs(10146) <= not(layer0_outputs(12117));
    outputs(10147) <= layer0_outputs(3180);
    outputs(10148) <= not((layer0_outputs(476)) or (layer0_outputs(3371)));
    outputs(10149) <= not(layer0_outputs(8142)) or (layer0_outputs(6390));
    outputs(10150) <= not(layer0_outputs(1618));
    outputs(10151) <= layer0_outputs(3890);
    outputs(10152) <= not((layer0_outputs(8565)) xor (layer0_outputs(6030)));
    outputs(10153) <= not((layer0_outputs(5777)) xor (layer0_outputs(7269)));
    outputs(10154) <= not(layer0_outputs(11778));
    outputs(10155) <= layer0_outputs(369);
    outputs(10156) <= not(layer0_outputs(320));
    outputs(10157) <= not((layer0_outputs(6416)) or (layer0_outputs(1822)));
    outputs(10158) <= not(layer0_outputs(11035));
    outputs(10159) <= layer0_outputs(5832);
    outputs(10160) <= (layer0_outputs(9606)) and not (layer0_outputs(1838));
    outputs(10161) <= not((layer0_outputs(2771)) or (layer0_outputs(4592)));
    outputs(10162) <= not((layer0_outputs(4139)) or (layer0_outputs(9978)));
    outputs(10163) <= (layer0_outputs(4062)) and (layer0_outputs(2157));
    outputs(10164) <= not(layer0_outputs(8398));
    outputs(10165) <= not(layer0_outputs(7643));
    outputs(10166) <= not((layer0_outputs(2592)) or (layer0_outputs(3991)));
    outputs(10167) <= (layer0_outputs(8931)) and not (layer0_outputs(10806));
    outputs(10168) <= not(layer0_outputs(38));
    outputs(10169) <= layer0_outputs(10368);
    outputs(10170) <= layer0_outputs(8240);
    outputs(10171) <= not((layer0_outputs(6700)) xor (layer0_outputs(9171)));
    outputs(10172) <= (layer0_outputs(3553)) and not (layer0_outputs(6372));
    outputs(10173) <= not(layer0_outputs(3354));
    outputs(10174) <= (layer0_outputs(6295)) xor (layer0_outputs(1338));
    outputs(10175) <= not((layer0_outputs(12269)) xor (layer0_outputs(12372)));
    outputs(10176) <= not(layer0_outputs(2940));
    outputs(10177) <= (layer0_outputs(9856)) and not (layer0_outputs(9136));
    outputs(10178) <= layer0_outputs(1683);
    outputs(10179) <= layer0_outputs(8432);
    outputs(10180) <= not((layer0_outputs(12313)) xor (layer0_outputs(12708)));
    outputs(10181) <= not(layer0_outputs(5149));
    outputs(10182) <= not(layer0_outputs(12384));
    outputs(10183) <= layer0_outputs(8712);
    outputs(10184) <= layer0_outputs(452);
    outputs(10185) <= (layer0_outputs(4584)) and not (layer0_outputs(8114));
    outputs(10186) <= not((layer0_outputs(12626)) xor (layer0_outputs(10410)));
    outputs(10187) <= not(layer0_outputs(9684));
    outputs(10188) <= not((layer0_outputs(3835)) or (layer0_outputs(2745)));
    outputs(10189) <= layer0_outputs(4504);
    outputs(10190) <= not(layer0_outputs(2449)) or (layer0_outputs(5932));
    outputs(10191) <= not(layer0_outputs(12152));
    outputs(10192) <= layer0_outputs(7559);
    outputs(10193) <= not(layer0_outputs(4707));
    outputs(10194) <= not(layer0_outputs(3336));
    outputs(10195) <= layer0_outputs(5270);
    outputs(10196) <= (layer0_outputs(3862)) xor (layer0_outputs(2865));
    outputs(10197) <= (layer0_outputs(1291)) and not (layer0_outputs(7713));
    outputs(10198) <= (layer0_outputs(2438)) xor (layer0_outputs(4219));
    outputs(10199) <= layer0_outputs(11958);
    outputs(10200) <= not((layer0_outputs(12421)) and (layer0_outputs(6273)));
    outputs(10201) <= layer0_outputs(8357);
    outputs(10202) <= not((layer0_outputs(3454)) xor (layer0_outputs(452)));
    outputs(10203) <= not(layer0_outputs(5906));
    outputs(10204) <= not(layer0_outputs(10404));
    outputs(10205) <= (layer0_outputs(3179)) and not (layer0_outputs(5772));
    outputs(10206) <= (layer0_outputs(4033)) and not (layer0_outputs(3405));
    outputs(10207) <= not(layer0_outputs(11803));
    outputs(10208) <= layer0_outputs(194);
    outputs(10209) <= (layer0_outputs(6982)) xor (layer0_outputs(5425));
    outputs(10210) <= not((layer0_outputs(6382)) xor (layer0_outputs(4624)));
    outputs(10211) <= layer0_outputs(3486);
    outputs(10212) <= not(layer0_outputs(5235)) or (layer0_outputs(4393));
    outputs(10213) <= not((layer0_outputs(3439)) or (layer0_outputs(9805)));
    outputs(10214) <= layer0_outputs(5318);
    outputs(10215) <= not(layer0_outputs(689));
    outputs(10216) <= not(layer0_outputs(1484));
    outputs(10217) <= (layer0_outputs(10799)) and not (layer0_outputs(11119));
    outputs(10218) <= layer0_outputs(2742);
    outputs(10219) <= not((layer0_outputs(725)) or (layer0_outputs(1868)));
    outputs(10220) <= layer0_outputs(906);
    outputs(10221) <= not(layer0_outputs(9590));
    outputs(10222) <= (layer0_outputs(10441)) and not (layer0_outputs(1083));
    outputs(10223) <= (layer0_outputs(11191)) and not (layer0_outputs(5607));
    outputs(10224) <= not(layer0_outputs(12263));
    outputs(10225) <= not(layer0_outputs(12287));
    outputs(10226) <= layer0_outputs(9444);
    outputs(10227) <= not(layer0_outputs(9362));
    outputs(10228) <= layer0_outputs(2095);
    outputs(10229) <= not(layer0_outputs(10779));
    outputs(10230) <= not((layer0_outputs(8914)) or (layer0_outputs(827)));
    outputs(10231) <= not(layer0_outputs(7505));
    outputs(10232) <= not((layer0_outputs(9878)) xor (layer0_outputs(6575)));
    outputs(10233) <= not(layer0_outputs(8108)) or (layer0_outputs(12550));
    outputs(10234) <= layer0_outputs(4868);
    outputs(10235) <= not((layer0_outputs(11255)) and (layer0_outputs(7702)));
    outputs(10236) <= (layer0_outputs(7327)) and not (layer0_outputs(1930));
    outputs(10237) <= not(layer0_outputs(8108));
    outputs(10238) <= layer0_outputs(3079);
    outputs(10239) <= layer0_outputs(5943);
    outputs(10240) <= layer0_outputs(5178);
    outputs(10241) <= not(layer0_outputs(6395));
    outputs(10242) <= not(layer0_outputs(7008));
    outputs(10243) <= (layer0_outputs(9365)) xor (layer0_outputs(3268));
    outputs(10244) <= layer0_outputs(5326);
    outputs(10245) <= not(layer0_outputs(3064)) or (layer0_outputs(1921));
    outputs(10246) <= (layer0_outputs(4306)) xor (layer0_outputs(3288));
    outputs(10247) <= (layer0_outputs(11497)) xor (layer0_outputs(8141));
    outputs(10248) <= not((layer0_outputs(10815)) xor (layer0_outputs(12046)));
    outputs(10249) <= layer0_outputs(5677);
    outputs(10250) <= not((layer0_outputs(12114)) xor (layer0_outputs(677)));
    outputs(10251) <= not(layer0_outputs(3540));
    outputs(10252) <= (layer0_outputs(2566)) xor (layer0_outputs(1756));
    outputs(10253) <= not((layer0_outputs(6400)) and (layer0_outputs(3740)));
    outputs(10254) <= layer0_outputs(8923);
    outputs(10255) <= (layer0_outputs(10740)) and not (layer0_outputs(9078));
    outputs(10256) <= (layer0_outputs(6224)) xor (layer0_outputs(2645));
    outputs(10257) <= (layer0_outputs(8077)) xor (layer0_outputs(4171));
    outputs(10258) <= not((layer0_outputs(5243)) xor (layer0_outputs(5060)));
    outputs(10259) <= layer0_outputs(11440);
    outputs(10260) <= layer0_outputs(5570);
    outputs(10261) <= not(layer0_outputs(6542));
    outputs(10262) <= layer0_outputs(7959);
    outputs(10263) <= not((layer0_outputs(9421)) xor (layer0_outputs(9934)));
    outputs(10264) <= (layer0_outputs(3580)) xor (layer0_outputs(2249));
    outputs(10265) <= not((layer0_outputs(4115)) xor (layer0_outputs(6622)));
    outputs(10266) <= not(layer0_outputs(10151)) or (layer0_outputs(6871));
    outputs(10267) <= not(layer0_outputs(2654)) or (layer0_outputs(3670));
    outputs(10268) <= not(layer0_outputs(27));
    outputs(10269) <= (layer0_outputs(7081)) and not (layer0_outputs(3097));
    outputs(10270) <= not((layer0_outputs(6949)) and (layer0_outputs(9932)));
    outputs(10271) <= layer0_outputs(6917);
    outputs(10272) <= not(layer0_outputs(4374));
    outputs(10273) <= layer0_outputs(2416);
    outputs(10274) <= (layer0_outputs(10271)) or (layer0_outputs(12592));
    outputs(10275) <= (layer0_outputs(3839)) xor (layer0_outputs(6430));
    outputs(10276) <= not(layer0_outputs(11163)) or (layer0_outputs(10612));
    outputs(10277) <= not(layer0_outputs(9570));
    outputs(10278) <= not(layer0_outputs(4132));
    outputs(10279) <= not(layer0_outputs(1499)) or (layer0_outputs(12725));
    outputs(10280) <= layer0_outputs(87);
    outputs(10281) <= not(layer0_outputs(1081));
    outputs(10282) <= (layer0_outputs(12482)) xor (layer0_outputs(3716));
    outputs(10283) <= not(layer0_outputs(10073));
    outputs(10284) <= layer0_outputs(5222);
    outputs(10285) <= not(layer0_outputs(3630));
    outputs(10286) <= not(layer0_outputs(7471));
    outputs(10287) <= (layer0_outputs(12188)) xor (layer0_outputs(8528));
    outputs(10288) <= layer0_outputs(9638);
    outputs(10289) <= not(layer0_outputs(2257));
    outputs(10290) <= not((layer0_outputs(6801)) xor (layer0_outputs(11715)));
    outputs(10291) <= layer0_outputs(6353);
    outputs(10292) <= not(layer0_outputs(7845));
    outputs(10293) <= not((layer0_outputs(375)) xor (layer0_outputs(8055)));
    outputs(10294) <= not(layer0_outputs(7628));
    outputs(10295) <= not(layer0_outputs(5962));
    outputs(10296) <= not(layer0_outputs(12176));
    outputs(10297) <= not(layer0_outputs(622)) or (layer0_outputs(6882));
    outputs(10298) <= layer0_outputs(12752);
    outputs(10299) <= not((layer0_outputs(7191)) and (layer0_outputs(11789)));
    outputs(10300) <= (layer0_outputs(6408)) xor (layer0_outputs(1033));
    outputs(10301) <= not(layer0_outputs(2777));
    outputs(10302) <= layer0_outputs(2438);
    outputs(10303) <= not((layer0_outputs(9953)) xor (layer0_outputs(10863)));
    outputs(10304) <= layer0_outputs(12027);
    outputs(10305) <= '1';
    outputs(10306) <= not(layer0_outputs(3604));
    outputs(10307) <= not(layer0_outputs(2)) or (layer0_outputs(3978));
    outputs(10308) <= layer0_outputs(12583);
    outputs(10309) <= (layer0_outputs(11948)) xor (layer0_outputs(975));
    outputs(10310) <= (layer0_outputs(5407)) xor (layer0_outputs(12352));
    outputs(10311) <= (layer0_outputs(6819)) xor (layer0_outputs(161));
    outputs(10312) <= not((layer0_outputs(4915)) and (layer0_outputs(1895)));
    outputs(10313) <= layer0_outputs(2114);
    outputs(10314) <= not((layer0_outputs(6901)) xor (layer0_outputs(12481)));
    outputs(10315) <= not(layer0_outputs(3996)) or (layer0_outputs(8050));
    outputs(10316) <= not((layer0_outputs(1386)) and (layer0_outputs(9893)));
    outputs(10317) <= not(layer0_outputs(5451));
    outputs(10318) <= layer0_outputs(9246);
    outputs(10319) <= not((layer0_outputs(12663)) xor (layer0_outputs(8952)));
    outputs(10320) <= not(layer0_outputs(8200)) or (layer0_outputs(1662));
    outputs(10321) <= (layer0_outputs(9427)) xor (layer0_outputs(6973));
    outputs(10322) <= layer0_outputs(3173);
    outputs(10323) <= (layer0_outputs(11979)) and not (layer0_outputs(660));
    outputs(10324) <= (layer0_outputs(5884)) xor (layer0_outputs(1833));
    outputs(10325) <= not(layer0_outputs(12031)) or (layer0_outputs(9222));
    outputs(10326) <= not(layer0_outputs(372));
    outputs(10327) <= (layer0_outputs(11002)) or (layer0_outputs(7689));
    outputs(10328) <= (layer0_outputs(201)) and not (layer0_outputs(12315));
    outputs(10329) <= layer0_outputs(10148);
    outputs(10330) <= layer0_outputs(2271);
    outputs(10331) <= layer0_outputs(2497);
    outputs(10332) <= layer0_outputs(3940);
    outputs(10333) <= not((layer0_outputs(1600)) or (layer0_outputs(1286)));
    outputs(10334) <= not(layer0_outputs(9408));
    outputs(10335) <= layer0_outputs(7050);
    outputs(10336) <= (layer0_outputs(3220)) xor (layer0_outputs(1484));
    outputs(10337) <= not((layer0_outputs(1029)) and (layer0_outputs(8948)));
    outputs(10338) <= not(layer0_outputs(10356));
    outputs(10339) <= (layer0_outputs(11392)) xor (layer0_outputs(11492));
    outputs(10340) <= not((layer0_outputs(9266)) xor (layer0_outputs(9916)));
    outputs(10341) <= layer0_outputs(1071);
    outputs(10342) <= layer0_outputs(8740);
    outputs(10343) <= not((layer0_outputs(12164)) xor (layer0_outputs(9395)));
    outputs(10344) <= not(layer0_outputs(994)) or (layer0_outputs(4221));
    outputs(10345) <= (layer0_outputs(10576)) or (layer0_outputs(11063));
    outputs(10346) <= not((layer0_outputs(10182)) xor (layer0_outputs(8060)));
    outputs(10347) <= not(layer0_outputs(5847)) or (layer0_outputs(12383));
    outputs(10348) <= (layer0_outputs(3890)) xor (layer0_outputs(7337));
    outputs(10349) <= not((layer0_outputs(12381)) xor (layer0_outputs(5538)));
    outputs(10350) <= not((layer0_outputs(9910)) xor (layer0_outputs(7730)));
    outputs(10351) <= not(layer0_outputs(8771)) or (layer0_outputs(7913));
    outputs(10352) <= (layer0_outputs(7511)) xor (layer0_outputs(7900));
    outputs(10353) <= not(layer0_outputs(255)) or (layer0_outputs(3214));
    outputs(10354) <= layer0_outputs(6246);
    outputs(10355) <= layer0_outputs(6592);
    outputs(10356) <= not((layer0_outputs(8571)) and (layer0_outputs(3752)));
    outputs(10357) <= not((layer0_outputs(10814)) and (layer0_outputs(1871)));
    outputs(10358) <= not(layer0_outputs(3085)) or (layer0_outputs(8995));
    outputs(10359) <= (layer0_outputs(6908)) xor (layer0_outputs(8980));
    outputs(10360) <= (layer0_outputs(7023)) and not (layer0_outputs(1109));
    outputs(10361) <= not(layer0_outputs(1398));
    outputs(10362) <= layer0_outputs(1110);
    outputs(10363) <= layer0_outputs(321);
    outputs(10364) <= not(layer0_outputs(2133)) or (layer0_outputs(3658));
    outputs(10365) <= (layer0_outputs(9707)) xor (layer0_outputs(11342));
    outputs(10366) <= (layer0_outputs(11402)) xor (layer0_outputs(3944));
    outputs(10367) <= not((layer0_outputs(4466)) xor (layer0_outputs(1039)));
    outputs(10368) <= not(layer0_outputs(9350));
    outputs(10369) <= not(layer0_outputs(5398));
    outputs(10370) <= not(layer0_outputs(5865));
    outputs(10371) <= not((layer0_outputs(6636)) xor (layer0_outputs(9860)));
    outputs(10372) <= (layer0_outputs(2199)) and not (layer0_outputs(2590));
    outputs(10373) <= layer0_outputs(11843);
    outputs(10374) <= not((layer0_outputs(11031)) xor (layer0_outputs(2313)));
    outputs(10375) <= layer0_outputs(1580);
    outputs(10376) <= not(layer0_outputs(12418));
    outputs(10377) <= not(layer0_outputs(5043)) or (layer0_outputs(6677));
    outputs(10378) <= not(layer0_outputs(4681)) or (layer0_outputs(8160));
    outputs(10379) <= not((layer0_outputs(8637)) xor (layer0_outputs(5486)));
    outputs(10380) <= layer0_outputs(9666);
    outputs(10381) <= not(layer0_outputs(12770)) or (layer0_outputs(2392));
    outputs(10382) <= (layer0_outputs(4351)) and not (layer0_outputs(3603));
    outputs(10383) <= not(layer0_outputs(11429));
    outputs(10384) <= (layer0_outputs(457)) or (layer0_outputs(9874));
    outputs(10385) <= (layer0_outputs(6748)) or (layer0_outputs(7557));
    outputs(10386) <= not(layer0_outputs(4380));
    outputs(10387) <= not((layer0_outputs(410)) xor (layer0_outputs(4516)));
    outputs(10388) <= layer0_outputs(6893);
    outputs(10389) <= not(layer0_outputs(2494)) or (layer0_outputs(11449));
    outputs(10390) <= not((layer0_outputs(6147)) xor (layer0_outputs(2252)));
    outputs(10391) <= not(layer0_outputs(6952));
    outputs(10392) <= (layer0_outputs(75)) xor (layer0_outputs(7666));
    outputs(10393) <= not((layer0_outputs(9731)) and (layer0_outputs(9896)));
    outputs(10394) <= layer0_outputs(12663);
    outputs(10395) <= (layer0_outputs(8238)) or (layer0_outputs(1932));
    outputs(10396) <= not((layer0_outputs(3222)) and (layer0_outputs(8405)));
    outputs(10397) <= not((layer0_outputs(12000)) and (layer0_outputs(1126)));
    outputs(10398) <= not(layer0_outputs(4294));
    outputs(10399) <= not((layer0_outputs(1569)) xor (layer0_outputs(11904)));
    outputs(10400) <= layer0_outputs(12423);
    outputs(10401) <= layer0_outputs(7743);
    outputs(10402) <= layer0_outputs(12510);
    outputs(10403) <= not((layer0_outputs(21)) xor (layer0_outputs(10216)));
    outputs(10404) <= (layer0_outputs(5006)) xor (layer0_outputs(6259));
    outputs(10405) <= not(layer0_outputs(3151)) or (layer0_outputs(4668));
    outputs(10406) <= not((layer0_outputs(4629)) xor (layer0_outputs(2988)));
    outputs(10407) <= not((layer0_outputs(11921)) xor (layer0_outputs(12365)));
    outputs(10408) <= layer0_outputs(11594);
    outputs(10409) <= (layer0_outputs(0)) xor (layer0_outputs(3926));
    outputs(10410) <= (layer0_outputs(4942)) or (layer0_outputs(8134));
    outputs(10411) <= layer0_outputs(3142);
    outputs(10412) <= (layer0_outputs(9869)) xor (layer0_outputs(232));
    outputs(10413) <= not(layer0_outputs(1460));
    outputs(10414) <= layer0_outputs(12255);
    outputs(10415) <= not((layer0_outputs(690)) and (layer0_outputs(11890)));
    outputs(10416) <= not(layer0_outputs(5150));
    outputs(10417) <= layer0_outputs(3512);
    outputs(10418) <= (layer0_outputs(8574)) or (layer0_outputs(3943));
    outputs(10419) <= (layer0_outputs(5516)) or (layer0_outputs(3608));
    outputs(10420) <= (layer0_outputs(6569)) xor (layer0_outputs(505));
    outputs(10421) <= (layer0_outputs(1416)) and not (layer0_outputs(12045));
    outputs(10422) <= not((layer0_outputs(6565)) and (layer0_outputs(7674)));
    outputs(10423) <= (layer0_outputs(2422)) or (layer0_outputs(11985));
    outputs(10424) <= (layer0_outputs(1327)) xor (layer0_outputs(12572));
    outputs(10425) <= not(layer0_outputs(6644)) or (layer0_outputs(11692));
    outputs(10426) <= layer0_outputs(5230);
    outputs(10427) <= not((layer0_outputs(3370)) xor (layer0_outputs(7095)));
    outputs(10428) <= (layer0_outputs(8073)) and not (layer0_outputs(2374));
    outputs(10429) <= layer0_outputs(11991);
    outputs(10430) <= not(layer0_outputs(8055));
    outputs(10431) <= not(layer0_outputs(1217));
    outputs(10432) <= not(layer0_outputs(8167)) or (layer0_outputs(3518));
    outputs(10433) <= not(layer0_outputs(11006));
    outputs(10434) <= (layer0_outputs(8832)) xor (layer0_outputs(318));
    outputs(10435) <= layer0_outputs(3713);
    outputs(10436) <= not((layer0_outputs(500)) xor (layer0_outputs(7206)));
    outputs(10437) <= not((layer0_outputs(7222)) xor (layer0_outputs(8)));
    outputs(10438) <= not((layer0_outputs(9323)) xor (layer0_outputs(2540)));
    outputs(10439) <= (layer0_outputs(12618)) and (layer0_outputs(4343));
    outputs(10440) <= not(layer0_outputs(9859));
    outputs(10441) <= layer0_outputs(790);
    outputs(10442) <= not(layer0_outputs(7942));
    outputs(10443) <= (layer0_outputs(1056)) and (layer0_outputs(6249));
    outputs(10444) <= not(layer0_outputs(10775)) or (layer0_outputs(9267));
    outputs(10445) <= (layer0_outputs(2179)) and not (layer0_outputs(10835));
    outputs(10446) <= (layer0_outputs(2309)) or (layer0_outputs(3101));
    outputs(10447) <= not((layer0_outputs(868)) or (layer0_outputs(11244)));
    outputs(10448) <= (layer0_outputs(4920)) xor (layer0_outputs(4802));
    outputs(10449) <= not(layer0_outputs(7416));
    outputs(10450) <= not(layer0_outputs(12718)) or (layer0_outputs(12081));
    outputs(10451) <= (layer0_outputs(12604)) xor (layer0_outputs(8932));
    outputs(10452) <= not(layer0_outputs(2328));
    outputs(10453) <= (layer0_outputs(9686)) xor (layer0_outputs(11962));
    outputs(10454) <= not((layer0_outputs(10121)) xor (layer0_outputs(2929)));
    outputs(10455) <= (layer0_outputs(12015)) xor (layer0_outputs(7770));
    outputs(10456) <= not(layer0_outputs(3866));
    outputs(10457) <= (layer0_outputs(3848)) or (layer0_outputs(2329));
    outputs(10458) <= not(layer0_outputs(11126)) or (layer0_outputs(1951));
    outputs(10459) <= layer0_outputs(12195);
    outputs(10460) <= layer0_outputs(6435);
    outputs(10461) <= (layer0_outputs(8773)) xor (layer0_outputs(9112));
    outputs(10462) <= (layer0_outputs(2895)) xor (layer0_outputs(9616));
    outputs(10463) <= layer0_outputs(3475);
    outputs(10464) <= not(layer0_outputs(6330)) or (layer0_outputs(5708));
    outputs(10465) <= layer0_outputs(3265);
    outputs(10466) <= layer0_outputs(3108);
    outputs(10467) <= not(layer0_outputs(4208));
    outputs(10468) <= not(layer0_outputs(6342)) or (layer0_outputs(7481));
    outputs(10469) <= not(layer0_outputs(5066)) or (layer0_outputs(1396));
    outputs(10470) <= not((layer0_outputs(11636)) xor (layer0_outputs(9057)));
    outputs(10471) <= not(layer0_outputs(7513)) or (layer0_outputs(10116));
    outputs(10472) <= (layer0_outputs(4619)) xor (layer0_outputs(10783));
    outputs(10473) <= (layer0_outputs(12515)) xor (layer0_outputs(4160));
    outputs(10474) <= not((layer0_outputs(1573)) or (layer0_outputs(312)));
    outputs(10475) <= not(layer0_outputs(5398)) or (layer0_outputs(11948));
    outputs(10476) <= not((layer0_outputs(2609)) xor (layer0_outputs(7944)));
    outputs(10477) <= (layer0_outputs(1219)) xor (layer0_outputs(2995));
    outputs(10478) <= not(layer0_outputs(4196));
    outputs(10479) <= not(layer0_outputs(1282)) or (layer0_outputs(6141));
    outputs(10480) <= not((layer0_outputs(6988)) and (layer0_outputs(684)));
    outputs(10481) <= not((layer0_outputs(4224)) xor (layer0_outputs(4500)));
    outputs(10482) <= (layer0_outputs(1653)) and not (layer0_outputs(12288));
    outputs(10483) <= (layer0_outputs(8572)) xor (layer0_outputs(2448));
    outputs(10484) <= (layer0_outputs(8300)) xor (layer0_outputs(8931));
    outputs(10485) <= not((layer0_outputs(10215)) xor (layer0_outputs(3573)));
    outputs(10486) <= layer0_outputs(9059);
    outputs(10487) <= not(layer0_outputs(6577));
    outputs(10488) <= not((layer0_outputs(12368)) xor (layer0_outputs(12505)));
    outputs(10489) <= (layer0_outputs(9211)) xor (layer0_outputs(2545));
    outputs(10490) <= layer0_outputs(4857);
    outputs(10491) <= not((layer0_outputs(10755)) xor (layer0_outputs(12509)));
    outputs(10492) <= not(layer0_outputs(7414)) or (layer0_outputs(12069));
    outputs(10493) <= layer0_outputs(12717);
    outputs(10494) <= (layer0_outputs(10180)) xor (layer0_outputs(214));
    outputs(10495) <= not(layer0_outputs(11860));
    outputs(10496) <= layer0_outputs(3613);
    outputs(10497) <= layer0_outputs(8568);
    outputs(10498) <= not((layer0_outputs(1736)) xor (layer0_outputs(3328)));
    outputs(10499) <= (layer0_outputs(7518)) or (layer0_outputs(7347));
    outputs(10500) <= not(layer0_outputs(10617));
    outputs(10501) <= (layer0_outputs(12235)) or (layer0_outputs(5159));
    outputs(10502) <= not((layer0_outputs(6567)) and (layer0_outputs(916)));
    outputs(10503) <= (layer0_outputs(11898)) and not (layer0_outputs(424));
    outputs(10504) <= (layer0_outputs(9824)) and (layer0_outputs(3203));
    outputs(10505) <= not((layer0_outputs(12168)) xor (layer0_outputs(8468)));
    outputs(10506) <= not((layer0_outputs(233)) and (layer0_outputs(6573)));
    outputs(10507) <= not(layer0_outputs(2439));
    outputs(10508) <= (layer0_outputs(9792)) xor (layer0_outputs(3187));
    outputs(10509) <= not(layer0_outputs(7737)) or (layer0_outputs(10875));
    outputs(10510) <= layer0_outputs(10493);
    outputs(10511) <= not((layer0_outputs(5270)) and (layer0_outputs(7572)));
    outputs(10512) <= layer0_outputs(5686);
    outputs(10513) <= (layer0_outputs(8506)) xor (layer0_outputs(7776));
    outputs(10514) <= (layer0_outputs(7038)) or (layer0_outputs(12077));
    outputs(10515) <= not(layer0_outputs(9366)) or (layer0_outputs(11046));
    outputs(10516) <= (layer0_outputs(486)) or (layer0_outputs(1621));
    outputs(10517) <= not((layer0_outputs(5207)) or (layer0_outputs(1312)));
    outputs(10518) <= not((layer0_outputs(7534)) and (layer0_outputs(10357)));
    outputs(10519) <= not((layer0_outputs(3574)) xor (layer0_outputs(10332)));
    outputs(10520) <= not((layer0_outputs(2068)) xor (layer0_outputs(173)));
    outputs(10521) <= layer0_outputs(7117);
    outputs(10522) <= layer0_outputs(5329);
    outputs(10523) <= not(layer0_outputs(1560));
    outputs(10524) <= not((layer0_outputs(8842)) xor (layer0_outputs(3964)));
    outputs(10525) <= not(layer0_outputs(4033));
    outputs(10526) <= not(layer0_outputs(10177)) or (layer0_outputs(4517));
    outputs(10527) <= layer0_outputs(7937);
    outputs(10528) <= not(layer0_outputs(7367));
    outputs(10529) <= layer0_outputs(514);
    outputs(10530) <= (layer0_outputs(2950)) xor (layer0_outputs(1112));
    outputs(10531) <= (layer0_outputs(7419)) xor (layer0_outputs(11269));
    outputs(10532) <= not(layer0_outputs(11475));
    outputs(10533) <= not((layer0_outputs(5237)) and (layer0_outputs(11310)));
    outputs(10534) <= (layer0_outputs(2446)) xor (layer0_outputs(10313));
    outputs(10535) <= (layer0_outputs(10202)) xor (layer0_outputs(8946));
    outputs(10536) <= layer0_outputs(7870);
    outputs(10537) <= not((layer0_outputs(11688)) and (layer0_outputs(2001)));
    outputs(10538) <= not((layer0_outputs(3321)) and (layer0_outputs(8425)));
    outputs(10539) <= layer0_outputs(3353);
    outputs(10540) <= layer0_outputs(6102);
    outputs(10541) <= not((layer0_outputs(5701)) xor (layer0_outputs(10954)));
    outputs(10542) <= (layer0_outputs(7012)) xor (layer0_outputs(3864));
    outputs(10543) <= layer0_outputs(11168);
    outputs(10544) <= (layer0_outputs(678)) xor (layer0_outputs(9946));
    outputs(10545) <= not((layer0_outputs(3039)) xor (layer0_outputs(1358)));
    outputs(10546) <= not(layer0_outputs(7205));
    outputs(10547) <= (layer0_outputs(385)) xor (layer0_outputs(6903));
    outputs(10548) <= not((layer0_outputs(5777)) and (layer0_outputs(5745)));
    outputs(10549) <= not(layer0_outputs(7191));
    outputs(10550) <= layer0_outputs(812);
    outputs(10551) <= (layer0_outputs(4519)) xor (layer0_outputs(7049));
    outputs(10552) <= not(layer0_outputs(8963)) or (layer0_outputs(8516));
    outputs(10553) <= not(layer0_outputs(1067));
    outputs(10554) <= not(layer0_outputs(4746)) or (layer0_outputs(12444));
    outputs(10555) <= not(layer0_outputs(907));
    outputs(10556) <= (layer0_outputs(7373)) or (layer0_outputs(3029));
    outputs(10557) <= not((layer0_outputs(11358)) or (layer0_outputs(12749)));
    outputs(10558) <= not(layer0_outputs(866));
    outputs(10559) <= not(layer0_outputs(4783)) or (layer0_outputs(10898));
    outputs(10560) <= (layer0_outputs(2880)) xor (layer0_outputs(4867));
    outputs(10561) <= not(layer0_outputs(4082));
    outputs(10562) <= not(layer0_outputs(10218));
    outputs(10563) <= (layer0_outputs(633)) or (layer0_outputs(9167));
    outputs(10564) <= (layer0_outputs(6444)) xor (layer0_outputs(9573));
    outputs(10565) <= not(layer0_outputs(7543));
    outputs(10566) <= (layer0_outputs(10604)) or (layer0_outputs(3495));
    outputs(10567) <= not(layer0_outputs(5640));
    outputs(10568) <= (layer0_outputs(5814)) xor (layer0_outputs(3388));
    outputs(10569) <= '1';
    outputs(10570) <= not(layer0_outputs(1233)) or (layer0_outputs(12128));
    outputs(10571) <= layer0_outputs(856);
    outputs(10572) <= not(layer0_outputs(12398)) or (layer0_outputs(2252));
    outputs(10573) <= not(layer0_outputs(1372)) or (layer0_outputs(12324));
    outputs(10574) <= not(layer0_outputs(11860));
    outputs(10575) <= not((layer0_outputs(288)) xor (layer0_outputs(2661)));
    outputs(10576) <= not(layer0_outputs(5640));
    outputs(10577) <= not((layer0_outputs(10513)) xor (layer0_outputs(5569)));
    outputs(10578) <= layer0_outputs(12203);
    outputs(10579) <= (layer0_outputs(4017)) xor (layer0_outputs(542));
    outputs(10580) <= not(layer0_outputs(7050)) or (layer0_outputs(7237));
    outputs(10581) <= layer0_outputs(2788);
    outputs(10582) <= (layer0_outputs(2216)) xor (layer0_outputs(5636));
    outputs(10583) <= layer0_outputs(5275);
    outputs(10584) <= (layer0_outputs(12646)) xor (layer0_outputs(12057));
    outputs(10585) <= not((layer0_outputs(12731)) and (layer0_outputs(497)));
    outputs(10586) <= not(layer0_outputs(2202));
    outputs(10587) <= not((layer0_outputs(10863)) and (layer0_outputs(4502)));
    outputs(10588) <= not((layer0_outputs(12244)) xor (layer0_outputs(1326)));
    outputs(10589) <= layer0_outputs(12617);
    outputs(10590) <= not(layer0_outputs(7595));
    outputs(10591) <= '1';
    outputs(10592) <= not((layer0_outputs(10711)) and (layer0_outputs(10132)));
    outputs(10593) <= layer0_outputs(2311);
    outputs(10594) <= layer0_outputs(11709);
    outputs(10595) <= layer0_outputs(1926);
    outputs(10596) <= not(layer0_outputs(5852)) or (layer0_outputs(9390));
    outputs(10597) <= not((layer0_outputs(9808)) and (layer0_outputs(5593)));
    outputs(10598) <= (layer0_outputs(12727)) xor (layer0_outputs(3214));
    outputs(10599) <= not(layer0_outputs(1372));
    outputs(10600) <= layer0_outputs(12207);
    outputs(10601) <= not((layer0_outputs(10053)) xor (layer0_outputs(11519)));
    outputs(10602) <= (layer0_outputs(5509)) xor (layer0_outputs(10769));
    outputs(10603) <= (layer0_outputs(6945)) xor (layer0_outputs(6501));
    outputs(10604) <= not(layer0_outputs(4394));
    outputs(10605) <= not((layer0_outputs(12784)) xor (layer0_outputs(10581)));
    outputs(10606) <= (layer0_outputs(11530)) or (layer0_outputs(7393));
    outputs(10607) <= (layer0_outputs(7258)) xor (layer0_outputs(9514));
    outputs(10608) <= (layer0_outputs(1661)) and not (layer0_outputs(11093));
    outputs(10609) <= not(layer0_outputs(1715)) or (layer0_outputs(6822));
    outputs(10610) <= layer0_outputs(6221);
    outputs(10611) <= not((layer0_outputs(7846)) xor (layer0_outputs(9621)));
    outputs(10612) <= not((layer0_outputs(8928)) xor (layer0_outputs(12737)));
    outputs(10613) <= not((layer0_outputs(3193)) and (layer0_outputs(6772)));
    outputs(10614) <= not((layer0_outputs(9334)) and (layer0_outputs(7338)));
    outputs(10615) <= not(layer0_outputs(12004));
    outputs(10616) <= layer0_outputs(6606);
    outputs(10617) <= not(layer0_outputs(12623));
    outputs(10618) <= (layer0_outputs(8010)) and (layer0_outputs(5526));
    outputs(10619) <= not(layer0_outputs(4076));
    outputs(10620) <= layer0_outputs(477);
    outputs(10621) <= layer0_outputs(4946);
    outputs(10622) <= not(layer0_outputs(267)) or (layer0_outputs(8203));
    outputs(10623) <= layer0_outputs(5082);
    outputs(10624) <= not(layer0_outputs(203));
    outputs(10625) <= not(layer0_outputs(12596));
    outputs(10626) <= not((layer0_outputs(6644)) and (layer0_outputs(12170)));
    outputs(10627) <= not((layer0_outputs(7596)) xor (layer0_outputs(5233)));
    outputs(10628) <= not(layer0_outputs(4869));
    outputs(10629) <= not(layer0_outputs(12574));
    outputs(10630) <= (layer0_outputs(9064)) or (layer0_outputs(3227));
    outputs(10631) <= not((layer0_outputs(10000)) xor (layer0_outputs(12778)));
    outputs(10632) <= (layer0_outputs(8509)) xor (layer0_outputs(1138));
    outputs(10633) <= (layer0_outputs(8839)) or (layer0_outputs(258));
    outputs(10634) <= (layer0_outputs(1713)) xor (layer0_outputs(10338));
    outputs(10635) <= not((layer0_outputs(5626)) or (layer0_outputs(9210)));
    outputs(10636) <= (layer0_outputs(3210)) xor (layer0_outputs(3145));
    outputs(10637) <= not((layer0_outputs(3643)) xor (layer0_outputs(637)));
    outputs(10638) <= not((layer0_outputs(10385)) xor (layer0_outputs(2586)));
    outputs(10639) <= not((layer0_outputs(9142)) xor (layer0_outputs(4911)));
    outputs(10640) <= not((layer0_outputs(2933)) and (layer0_outputs(12165)));
    outputs(10641) <= (layer0_outputs(8709)) and (layer0_outputs(1099));
    outputs(10642) <= '1';
    outputs(10643) <= layer0_outputs(3119);
    outputs(10644) <= not(layer0_outputs(1327));
    outputs(10645) <= (layer0_outputs(5299)) and not (layer0_outputs(4486));
    outputs(10646) <= not((layer0_outputs(11566)) xor (layer0_outputs(4692)));
    outputs(10647) <= not((layer0_outputs(341)) xor (layer0_outputs(6122)));
    outputs(10648) <= not(layer0_outputs(1406));
    outputs(10649) <= not((layer0_outputs(11641)) xor (layer0_outputs(9512)));
    outputs(10650) <= not(layer0_outputs(1408));
    outputs(10651) <= not(layer0_outputs(6160)) or (layer0_outputs(11090));
    outputs(10652) <= layer0_outputs(1490);
    outputs(10653) <= not((layer0_outputs(1389)) and (layer0_outputs(2563)));
    outputs(10654) <= (layer0_outputs(3994)) or (layer0_outputs(5271));
    outputs(10655) <= not(layer0_outputs(8379)) or (layer0_outputs(8822));
    outputs(10656) <= not(layer0_outputs(6340));
    outputs(10657) <= not(layer0_outputs(6468));
    outputs(10658) <= layer0_outputs(12219);
    outputs(10659) <= not(layer0_outputs(2709));
    outputs(10660) <= not((layer0_outputs(11337)) and (layer0_outputs(6144)));
    outputs(10661) <= not(layer0_outputs(830));
    outputs(10662) <= not(layer0_outputs(3920));
    outputs(10663) <= not(layer0_outputs(4118));
    outputs(10664) <= layer0_outputs(8778);
    outputs(10665) <= not(layer0_outputs(5293));
    outputs(10666) <= not(layer0_outputs(5015));
    outputs(10667) <= not(layer0_outputs(12545));
    outputs(10668) <= not((layer0_outputs(5274)) xor (layer0_outputs(1058)));
    outputs(10669) <= not((layer0_outputs(8756)) xor (layer0_outputs(5539)));
    outputs(10670) <= (layer0_outputs(5340)) and (layer0_outputs(9072));
    outputs(10671) <= not((layer0_outputs(2522)) and (layer0_outputs(7934)));
    outputs(10672) <= layer0_outputs(6826);
    outputs(10673) <= not((layer0_outputs(10143)) xor (layer0_outputs(9826)));
    outputs(10674) <= not((layer0_outputs(8239)) or (layer0_outputs(10835)));
    outputs(10675) <= not(layer0_outputs(8474)) or (layer0_outputs(11925));
    outputs(10676) <= not((layer0_outputs(6285)) xor (layer0_outputs(491)));
    outputs(10677) <= (layer0_outputs(12518)) xor (layer0_outputs(11648));
    outputs(10678) <= not(layer0_outputs(3842));
    outputs(10679) <= (layer0_outputs(6914)) xor (layer0_outputs(2048));
    outputs(10680) <= not(layer0_outputs(8221));
    outputs(10681) <= not(layer0_outputs(7099));
    outputs(10682) <= (layer0_outputs(11282)) and (layer0_outputs(8916));
    outputs(10683) <= not((layer0_outputs(1346)) xor (layer0_outputs(1359)));
    outputs(10684) <= not((layer0_outputs(5727)) xor (layer0_outputs(8815)));
    outputs(10685) <= not(layer0_outputs(721)) or (layer0_outputs(2543));
    outputs(10686) <= layer0_outputs(10795);
    outputs(10687) <= not((layer0_outputs(9426)) xor (layer0_outputs(160)));
    outputs(10688) <= not((layer0_outputs(10023)) and (layer0_outputs(9144)));
    outputs(10689) <= (layer0_outputs(7976)) and not (layer0_outputs(1370));
    outputs(10690) <= (layer0_outputs(11345)) xor (layer0_outputs(880));
    outputs(10691) <= not(layer0_outputs(970));
    outputs(10692) <= not((layer0_outputs(9568)) xor (layer0_outputs(404)));
    outputs(10693) <= (layer0_outputs(789)) or (layer0_outputs(11911));
    outputs(10694) <= not((layer0_outputs(5175)) xor (layer0_outputs(5169)));
    outputs(10695) <= not(layer0_outputs(5672));
    outputs(10696) <= (layer0_outputs(8430)) xor (layer0_outputs(3722));
    outputs(10697) <= not((layer0_outputs(6598)) xor (layer0_outputs(5632)));
    outputs(10698) <= layer0_outputs(5122);
    outputs(10699) <= not(layer0_outputs(5513)) or (layer0_outputs(369));
    outputs(10700) <= (layer0_outputs(3018)) and (layer0_outputs(368));
    outputs(10701) <= not((layer0_outputs(12494)) xor (layer0_outputs(4004)));
    outputs(10702) <= layer0_outputs(7693);
    outputs(10703) <= not((layer0_outputs(6551)) xor (layer0_outputs(7481)));
    outputs(10704) <= not((layer0_outputs(5211)) xor (layer0_outputs(2131)));
    outputs(10705) <= layer0_outputs(3133);
    outputs(10706) <= layer0_outputs(8369);
    outputs(10707) <= not((layer0_outputs(11653)) or (layer0_outputs(12243)));
    outputs(10708) <= not(layer0_outputs(11672));
    outputs(10709) <= (layer0_outputs(950)) or (layer0_outputs(6058));
    outputs(10710) <= not((layer0_outputs(4997)) and (layer0_outputs(2869)));
    outputs(10711) <= (layer0_outputs(3420)) and not (layer0_outputs(7479));
    outputs(10712) <= (layer0_outputs(8268)) xor (layer0_outputs(5249));
    outputs(10713) <= not((layer0_outputs(2010)) xor (layer0_outputs(7810)));
    outputs(10714) <= not(layer0_outputs(4594));
    outputs(10715) <= (layer0_outputs(10839)) and not (layer0_outputs(2361));
    outputs(10716) <= not(layer0_outputs(12234));
    outputs(10717) <= layer0_outputs(6983);
    outputs(10718) <= not((layer0_outputs(7282)) xor (layer0_outputs(5186)));
    outputs(10719) <= not(layer0_outputs(890)) or (layer0_outputs(6943));
    outputs(10720) <= not(layer0_outputs(7742));
    outputs(10721) <= not((layer0_outputs(7158)) and (layer0_outputs(4653)));
    outputs(10722) <= not(layer0_outputs(7822)) or (layer0_outputs(239));
    outputs(10723) <= (layer0_outputs(7902)) and not (layer0_outputs(7745));
    outputs(10724) <= '1';
    outputs(10725) <= not((layer0_outputs(11895)) and (layer0_outputs(3074)));
    outputs(10726) <= not(layer0_outputs(1241));
    outputs(10727) <= not((layer0_outputs(5500)) or (layer0_outputs(811)));
    outputs(10728) <= not((layer0_outputs(12597)) xor (layer0_outputs(10422)));
    outputs(10729) <= not((layer0_outputs(11963)) and (layer0_outputs(3957)));
    outputs(10730) <= (layer0_outputs(9338)) or (layer0_outputs(90));
    outputs(10731) <= (layer0_outputs(9129)) and (layer0_outputs(4098));
    outputs(10732) <= not((layer0_outputs(6915)) and (layer0_outputs(12317)));
    outputs(10733) <= not(layer0_outputs(12783));
    outputs(10734) <= (layer0_outputs(11203)) and (layer0_outputs(9882));
    outputs(10735) <= (layer0_outputs(11608)) xor (layer0_outputs(5690));
    outputs(10736) <= not(layer0_outputs(9389)) or (layer0_outputs(12779));
    outputs(10737) <= not(layer0_outputs(10910));
    outputs(10738) <= (layer0_outputs(5512)) or (layer0_outputs(8043));
    outputs(10739) <= not((layer0_outputs(2279)) and (layer0_outputs(628)));
    outputs(10740) <= not(layer0_outputs(1411));
    outputs(10741) <= (layer0_outputs(10208)) xor (layer0_outputs(5506));
    outputs(10742) <= not((layer0_outputs(11167)) and (layer0_outputs(11310)));
    outputs(10743) <= not(layer0_outputs(1322));
    outputs(10744) <= not(layer0_outputs(1678)) or (layer0_outputs(8290));
    outputs(10745) <= (layer0_outputs(5712)) or (layer0_outputs(2888));
    outputs(10746) <= not(layer0_outputs(10627)) or (layer0_outputs(4227));
    outputs(10747) <= not((layer0_outputs(12304)) and (layer0_outputs(9287)));
    outputs(10748) <= layer0_outputs(2634);
    outputs(10749) <= not((layer0_outputs(3460)) xor (layer0_outputs(10281)));
    outputs(10750) <= not((layer0_outputs(9598)) xor (layer0_outputs(6196)));
    outputs(10751) <= not(layer0_outputs(5614));
    outputs(10752) <= not(layer0_outputs(4095)) or (layer0_outputs(12143));
    outputs(10753) <= (layer0_outputs(3826)) or (layer0_outputs(378));
    outputs(10754) <= not(layer0_outputs(9534));
    outputs(10755) <= not((layer0_outputs(1911)) and (layer0_outputs(362)));
    outputs(10756) <= layer0_outputs(8987);
    outputs(10757) <= not((layer0_outputs(4575)) or (layer0_outputs(6447)));
    outputs(10758) <= (layer0_outputs(8478)) or (layer0_outputs(10702));
    outputs(10759) <= not(layer0_outputs(9547)) or (layer0_outputs(2115));
    outputs(10760) <= layer0_outputs(10576);
    outputs(10761) <= not(layer0_outputs(7020));
    outputs(10762) <= not((layer0_outputs(11216)) and (layer0_outputs(5943)));
    outputs(10763) <= layer0_outputs(12096);
    outputs(10764) <= not(layer0_outputs(11045));
    outputs(10765) <= (layer0_outputs(8744)) xor (layer0_outputs(114));
    outputs(10766) <= layer0_outputs(5568);
    outputs(10767) <= not(layer0_outputs(11512)) or (layer0_outputs(3865));
    outputs(10768) <= not(layer0_outputs(3970));
    outputs(10769) <= not(layer0_outputs(8376));
    outputs(10770) <= (layer0_outputs(9774)) and not (layer0_outputs(7073));
    outputs(10771) <= not((layer0_outputs(12001)) and (layer0_outputs(11811)));
    outputs(10772) <= layer0_outputs(11523);
    outputs(10773) <= not((layer0_outputs(5219)) xor (layer0_outputs(7112)));
    outputs(10774) <= (layer0_outputs(1921)) and not (layer0_outputs(7205));
    outputs(10775) <= not((layer0_outputs(3318)) and (layer0_outputs(7408)));
    outputs(10776) <= not(layer0_outputs(5011));
    outputs(10777) <= not((layer0_outputs(6104)) xor (layer0_outputs(2815)));
    outputs(10778) <= not(layer0_outputs(9501));
    outputs(10779) <= (layer0_outputs(9795)) xor (layer0_outputs(5094));
    outputs(10780) <= not((layer0_outputs(5746)) xor (layer0_outputs(12163)));
    outputs(10781) <= layer0_outputs(6839);
    outputs(10782) <= layer0_outputs(422);
    outputs(10783) <= not((layer0_outputs(12344)) xor (layer0_outputs(2867)));
    outputs(10784) <= (layer0_outputs(6274)) and not (layer0_outputs(11145));
    outputs(10785) <= not(layer0_outputs(8386));
    outputs(10786) <= (layer0_outputs(669)) and not (layer0_outputs(1262));
    outputs(10787) <= not(layer0_outputs(6587));
    outputs(10788) <= (layer0_outputs(6936)) and not (layer0_outputs(10445));
    outputs(10789) <= not(layer0_outputs(10353));
    outputs(10790) <= not((layer0_outputs(7660)) xor (layer0_outputs(896)));
    outputs(10791) <= (layer0_outputs(5287)) and not (layer0_outputs(4185));
    outputs(10792) <= layer0_outputs(5366);
    outputs(10793) <= not((layer0_outputs(10419)) xor (layer0_outputs(9030)));
    outputs(10794) <= layer0_outputs(7365);
    outputs(10795) <= not(layer0_outputs(877)) or (layer0_outputs(1686));
    outputs(10796) <= layer0_outputs(1873);
    outputs(10797) <= layer0_outputs(8173);
    outputs(10798) <= layer0_outputs(1463);
    outputs(10799) <= (layer0_outputs(8283)) xor (layer0_outputs(530));
    outputs(10800) <= not((layer0_outputs(12122)) xor (layer0_outputs(3525)));
    outputs(10801) <= (layer0_outputs(1192)) or (layer0_outputs(6703));
    outputs(10802) <= (layer0_outputs(8227)) xor (layer0_outputs(8205));
    outputs(10803) <= (layer0_outputs(2348)) or (layer0_outputs(4624));
    outputs(10804) <= (layer0_outputs(3845)) xor (layer0_outputs(3461));
    outputs(10805) <= not(layer0_outputs(5266));
    outputs(10806) <= not(layer0_outputs(9143));
    outputs(10807) <= (layer0_outputs(5985)) xor (layer0_outputs(5585));
    outputs(10808) <= not(layer0_outputs(3129));
    outputs(10809) <= not(layer0_outputs(4244));
    outputs(10810) <= (layer0_outputs(6316)) xor (layer0_outputs(4192));
    outputs(10811) <= (layer0_outputs(8450)) and not (layer0_outputs(347));
    outputs(10812) <= not(layer0_outputs(4183));
    outputs(10813) <= (layer0_outputs(247)) xor (layer0_outputs(8959));
    outputs(10814) <= not(layer0_outputs(11901)) or (layer0_outputs(8498));
    outputs(10815) <= not((layer0_outputs(11808)) xor (layer0_outputs(8087)));
    outputs(10816) <= not((layer0_outputs(1523)) and (layer0_outputs(10455)));
    outputs(10817) <= not(layer0_outputs(11548));
    outputs(10818) <= not(layer0_outputs(12776)) or (layer0_outputs(5841));
    outputs(10819) <= (layer0_outputs(5655)) and not (layer0_outputs(1263));
    outputs(10820) <= not(layer0_outputs(12641)) or (layer0_outputs(11403));
    outputs(10821) <= layer0_outputs(1781);
    outputs(10822) <= (layer0_outputs(10138)) and not (layer0_outputs(11252));
    outputs(10823) <= not(layer0_outputs(5688));
    outputs(10824) <= not(layer0_outputs(11285));
    outputs(10825) <= not((layer0_outputs(11012)) and (layer0_outputs(8193)));
    outputs(10826) <= (layer0_outputs(11498)) xor (layer0_outputs(6765));
    outputs(10827) <= not(layer0_outputs(1393)) or (layer0_outputs(12582));
    outputs(10828) <= (layer0_outputs(730)) and (layer0_outputs(5495));
    outputs(10829) <= not((layer0_outputs(9343)) or (layer0_outputs(10963)));
    outputs(10830) <= (layer0_outputs(5615)) xor (layer0_outputs(2971));
    outputs(10831) <= not(layer0_outputs(3526));
    outputs(10832) <= layer0_outputs(8893);
    outputs(10833) <= layer0_outputs(8487);
    outputs(10834) <= (layer0_outputs(7851)) or (layer0_outputs(2004));
    outputs(10835) <= not(layer0_outputs(9940));
    outputs(10836) <= not((layer0_outputs(5864)) xor (layer0_outputs(1104)));
    outputs(10837) <= not((layer0_outputs(570)) xor (layer0_outputs(2194)));
    outputs(10838) <= (layer0_outputs(12669)) xor (layer0_outputs(12707));
    outputs(10839) <= (layer0_outputs(4803)) and not (layer0_outputs(7707));
    outputs(10840) <= not(layer0_outputs(548));
    outputs(10841) <= layer0_outputs(8937);
    outputs(10842) <= not((layer0_outputs(9285)) or (layer0_outputs(12018)));
    outputs(10843) <= (layer0_outputs(6879)) and not (layer0_outputs(455));
    outputs(10844) <= not(layer0_outputs(7689));
    outputs(10845) <= not((layer0_outputs(8715)) xor (layer0_outputs(10742)));
    outputs(10846) <= not(layer0_outputs(1601));
    outputs(10847) <= not((layer0_outputs(11646)) xor (layer0_outputs(3737)));
    outputs(10848) <= not(layer0_outputs(9649)) or (layer0_outputs(9667));
    outputs(10849) <= not((layer0_outputs(1520)) and (layer0_outputs(6884)));
    outputs(10850) <= not(layer0_outputs(4842));
    outputs(10851) <= (layer0_outputs(2618)) xor (layer0_outputs(2952));
    outputs(10852) <= (layer0_outputs(566)) xor (layer0_outputs(1425));
    outputs(10853) <= not(layer0_outputs(12661)) or (layer0_outputs(8981));
    outputs(10854) <= not((layer0_outputs(945)) xor (layer0_outputs(10780)));
    outputs(10855) <= layer0_outputs(3539);
    outputs(10856) <= (layer0_outputs(3803)) or (layer0_outputs(12124));
    outputs(10857) <= not(layer0_outputs(5201));
    outputs(10858) <= not(layer0_outputs(191));
    outputs(10859) <= (layer0_outputs(12588)) xor (layer0_outputs(5670));
    outputs(10860) <= not((layer0_outputs(4030)) xor (layer0_outputs(3172)));
    outputs(10861) <= not((layer0_outputs(10957)) or (layer0_outputs(4147)));
    outputs(10862) <= (layer0_outputs(10183)) or (layer0_outputs(600));
    outputs(10863) <= not((layer0_outputs(6318)) or (layer0_outputs(3116)));
    outputs(10864) <= not((layer0_outputs(9748)) xor (layer0_outputs(10816)));
    outputs(10865) <= (layer0_outputs(6145)) and not (layer0_outputs(5184));
    outputs(10866) <= not((layer0_outputs(6300)) xor (layer0_outputs(7292)));
    outputs(10867) <= not(layer0_outputs(195));
    outputs(10868) <= not(layer0_outputs(3882)) or (layer0_outputs(5502));
    outputs(10869) <= (layer0_outputs(3030)) and not (layer0_outputs(5924));
    outputs(10870) <= not((layer0_outputs(2974)) xor (layer0_outputs(9047)));
    outputs(10871) <= not((layer0_outputs(1216)) xor (layer0_outputs(2385)));
    outputs(10872) <= (layer0_outputs(11535)) xor (layer0_outputs(3401));
    outputs(10873) <= not(layer0_outputs(7430)) or (layer0_outputs(3881));
    outputs(10874) <= not(layer0_outputs(6596));
    outputs(10875) <= not(layer0_outputs(5440)) or (layer0_outputs(6310));
    outputs(10876) <= not((layer0_outputs(9309)) xor (layer0_outputs(9668)));
    outputs(10877) <= not((layer0_outputs(782)) xor (layer0_outputs(9113)));
    outputs(10878) <= layer0_outputs(9925);
    outputs(10879) <= (layer0_outputs(6732)) and not (layer0_outputs(10599));
    outputs(10880) <= (layer0_outputs(3685)) or (layer0_outputs(5550));
    outputs(10881) <= not((layer0_outputs(3856)) or (layer0_outputs(3780)));
    outputs(10882) <= not((layer0_outputs(5361)) or (layer0_outputs(592)));
    outputs(10883) <= not(layer0_outputs(9440)) or (layer0_outputs(12262));
    outputs(10884) <= not(layer0_outputs(2170));
    outputs(10885) <= (layer0_outputs(12376)) or (layer0_outputs(10049));
    outputs(10886) <= not((layer0_outputs(4707)) xor (layer0_outputs(6245)));
    outputs(10887) <= not((layer0_outputs(10257)) and (layer0_outputs(6867)));
    outputs(10888) <= (layer0_outputs(11505)) and not (layer0_outputs(9044));
    outputs(10889) <= not(layer0_outputs(7087)) or (layer0_outputs(9034));
    outputs(10890) <= not(layer0_outputs(3612)) or (layer0_outputs(1811));
    outputs(10891) <= (layer0_outputs(7701)) xor (layer0_outputs(8051));
    outputs(10892) <= not((layer0_outputs(5542)) xor (layer0_outputs(3391)));
    outputs(10893) <= not(layer0_outputs(10421)) or (layer0_outputs(10446));
    outputs(10894) <= not(layer0_outputs(6751));
    outputs(10895) <= not(layer0_outputs(7350)) or (layer0_outputs(1013));
    outputs(10896) <= not(layer0_outputs(1727));
    outputs(10897) <= not((layer0_outputs(3451)) xor (layer0_outputs(8784)));
    outputs(10898) <= not((layer0_outputs(7352)) xor (layer0_outputs(9238)));
    outputs(10899) <= not((layer0_outputs(12088)) xor (layer0_outputs(12318)));
    outputs(10900) <= layer0_outputs(11422);
    outputs(10901) <= not(layer0_outputs(8495)) or (layer0_outputs(7351));
    outputs(10902) <= not((layer0_outputs(1095)) xor (layer0_outputs(9414)));
    outputs(10903) <= layer0_outputs(11333);
    outputs(10904) <= (layer0_outputs(1896)) xor (layer0_outputs(7694));
    outputs(10905) <= (layer0_outputs(11077)) xor (layer0_outputs(4008));
    outputs(10906) <= not(layer0_outputs(4408)) or (layer0_outputs(11679));
    outputs(10907) <= not((layer0_outputs(5562)) and (layer0_outputs(10416)));
    outputs(10908) <= not((layer0_outputs(3277)) xor (layer0_outputs(5667)));
    outputs(10909) <= layer0_outputs(4968);
    outputs(10910) <= layer0_outputs(6591);
    outputs(10911) <= (layer0_outputs(2206)) xor (layer0_outputs(11659));
    outputs(10912) <= layer0_outputs(2670);
    outputs(10913) <= (layer0_outputs(12179)) xor (layer0_outputs(8132));
    outputs(10914) <= not((layer0_outputs(2770)) or (layer0_outputs(4939)));
    outputs(10915) <= not(layer0_outputs(3325)) or (layer0_outputs(4276));
    outputs(10916) <= (layer0_outputs(129)) xor (layer0_outputs(12553));
    outputs(10917) <= (layer0_outputs(6407)) and not (layer0_outputs(7016));
    outputs(10918) <= not(layer0_outputs(11889));
    outputs(10919) <= (layer0_outputs(7555)) or (layer0_outputs(11003));
    outputs(10920) <= not(layer0_outputs(8613));
    outputs(10921) <= not(layer0_outputs(12369));
    outputs(10922) <= not((layer0_outputs(1620)) xor (layer0_outputs(5381)));
    outputs(10923) <= (layer0_outputs(8600)) and not (layer0_outputs(12587));
    outputs(10924) <= not(layer0_outputs(9219));
    outputs(10925) <= not(layer0_outputs(12631)) or (layer0_outputs(11782));
    outputs(10926) <= layer0_outputs(11392);
    outputs(10927) <= not(layer0_outputs(6026));
    outputs(10928) <= layer0_outputs(784);
    outputs(10929) <= not(layer0_outputs(8083)) or (layer0_outputs(11908));
    outputs(10930) <= not(layer0_outputs(4071)) or (layer0_outputs(5433));
    outputs(10931) <= (layer0_outputs(9237)) or (layer0_outputs(4514));
    outputs(10932) <= (layer0_outputs(2603)) xor (layer0_outputs(5306));
    outputs(10933) <= (layer0_outputs(10790)) or (layer0_outputs(7353));
    outputs(10934) <= not(layer0_outputs(4057)) or (layer0_outputs(4030));
    outputs(10935) <= layer0_outputs(658);
    outputs(10936) <= not(layer0_outputs(9055)) or (layer0_outputs(3728));
    outputs(10937) <= (layer0_outputs(7227)) xor (layer0_outputs(5766));
    outputs(10938) <= layer0_outputs(10399);
    outputs(10939) <= (layer0_outputs(1157)) xor (layer0_outputs(12741));
    outputs(10940) <= not(layer0_outputs(2786));
    outputs(10941) <= not((layer0_outputs(12451)) and (layer0_outputs(2711)));
    outputs(10942) <= layer0_outputs(1676);
    outputs(10943) <= not((layer0_outputs(7119)) xor (layer0_outputs(8411)));
    outputs(10944) <= layer0_outputs(514);
    outputs(10945) <= layer0_outputs(4455);
    outputs(10946) <= layer0_outputs(9267);
    outputs(10947) <= not((layer0_outputs(12345)) or (layer0_outputs(2486)));
    outputs(10948) <= not((layer0_outputs(5844)) xor (layer0_outputs(5801)));
    outputs(10949) <= (layer0_outputs(12036)) or (layer0_outputs(9817));
    outputs(10950) <= (layer0_outputs(766)) or (layer0_outputs(3941));
    outputs(10951) <= not(layer0_outputs(6380));
    outputs(10952) <= layer0_outputs(6407);
    outputs(10953) <= (layer0_outputs(3397)) xor (layer0_outputs(1377));
    outputs(10954) <= not((layer0_outputs(9074)) xor (layer0_outputs(2892)));
    outputs(10955) <= layer0_outputs(7772);
    outputs(10956) <= not(layer0_outputs(2339)) or (layer0_outputs(9006));
    outputs(10957) <= layer0_outputs(5992);
    outputs(10958) <= not((layer0_outputs(1216)) and (layer0_outputs(9759)));
    outputs(10959) <= not((layer0_outputs(5323)) xor (layer0_outputs(11103)));
    outputs(10960) <= (layer0_outputs(11376)) xor (layer0_outputs(5899));
    outputs(10961) <= not((layer0_outputs(6357)) xor (layer0_outputs(7009)));
    outputs(10962) <= not((layer0_outputs(5405)) and (layer0_outputs(3021)));
    outputs(10963) <= layer0_outputs(12797);
    outputs(10964) <= (layer0_outputs(7295)) xor (layer0_outputs(5437));
    outputs(10965) <= (layer0_outputs(4542)) or (layer0_outputs(6911));
    outputs(10966) <= not(layer0_outputs(10201)) or (layer0_outputs(7687));
    outputs(10967) <= (layer0_outputs(7182)) xor (layer0_outputs(12515));
    outputs(10968) <= not(layer0_outputs(7560));
    outputs(10969) <= layer0_outputs(7103);
    outputs(10970) <= not(layer0_outputs(2569));
    outputs(10971) <= layer0_outputs(11256);
    outputs(10972) <= not((layer0_outputs(278)) xor (layer0_outputs(7232)));
    outputs(10973) <= not(layer0_outputs(315));
    outputs(10974) <= not(layer0_outputs(7291));
    outputs(10975) <= (layer0_outputs(7846)) xor (layer0_outputs(6277));
    outputs(10976) <= not(layer0_outputs(6470)) or (layer0_outputs(1224));
    outputs(10977) <= layer0_outputs(9332);
    outputs(10978) <= not(layer0_outputs(1974));
    outputs(10979) <= not((layer0_outputs(709)) or (layer0_outputs(3679)));
    outputs(10980) <= not(layer0_outputs(8090));
    outputs(10981) <= not(layer0_outputs(3730));
    outputs(10982) <= not(layer0_outputs(12672));
    outputs(10983) <= not(layer0_outputs(2598)) or (layer0_outputs(8820));
    outputs(10984) <= not((layer0_outputs(8289)) or (layer0_outputs(3504)));
    outputs(10985) <= (layer0_outputs(10470)) and (layer0_outputs(1363));
    outputs(10986) <= (layer0_outputs(11597)) xor (layer0_outputs(8291));
    outputs(10987) <= not(layer0_outputs(11371));
    outputs(10988) <= not(layer0_outputs(2898));
    outputs(10989) <= (layer0_outputs(6674)) xor (layer0_outputs(7431));
    outputs(10990) <= layer0_outputs(10791);
    outputs(10991) <= (layer0_outputs(7076)) or (layer0_outputs(2079));
    outputs(10992) <= (layer0_outputs(7832)) and not (layer0_outputs(11088));
    outputs(10993) <= layer0_outputs(7437);
    outputs(10994) <= layer0_outputs(11494);
    outputs(10995) <= layer0_outputs(6864);
    outputs(10996) <= not(layer0_outputs(2147));
    outputs(10997) <= not(layer0_outputs(9163));
    outputs(10998) <= (layer0_outputs(3918)) and not (layer0_outputs(2687));
    outputs(10999) <= not(layer0_outputs(8115));
    outputs(11000) <= not((layer0_outputs(9454)) and (layer0_outputs(4108)));
    outputs(11001) <= not((layer0_outputs(7608)) xor (layer0_outputs(4141)));
    outputs(11002) <= (layer0_outputs(11795)) xor (layer0_outputs(2893));
    outputs(11003) <= not(layer0_outputs(442));
    outputs(11004) <= not((layer0_outputs(3810)) or (layer0_outputs(2611)));
    outputs(11005) <= not((layer0_outputs(9961)) xor (layer0_outputs(10648)));
    outputs(11006) <= (layer0_outputs(2212)) xor (layer0_outputs(9625));
    outputs(11007) <= not(layer0_outputs(7768));
    outputs(11008) <= not(layer0_outputs(6052)) or (layer0_outputs(5187));
    outputs(11009) <= layer0_outputs(1595);
    outputs(11010) <= not(layer0_outputs(3425));
    outputs(11011) <= layer0_outputs(6637);
    outputs(11012) <= (layer0_outputs(8278)) and not (layer0_outputs(12201));
    outputs(11013) <= (layer0_outputs(6246)) xor (layer0_outputs(3880));
    outputs(11014) <= not((layer0_outputs(874)) xor (layer0_outputs(645)));
    outputs(11015) <= not((layer0_outputs(9820)) xor (layer0_outputs(4647)));
    outputs(11016) <= not(layer0_outputs(8280));
    outputs(11017) <= not((layer0_outputs(10258)) and (layer0_outputs(318)));
    outputs(11018) <= not((layer0_outputs(2445)) and (layer0_outputs(4468)));
    outputs(11019) <= not((layer0_outputs(7395)) and (layer0_outputs(209)));
    outputs(11020) <= (layer0_outputs(3800)) xor (layer0_outputs(8879));
    outputs(11021) <= layer0_outputs(8632);
    outputs(11022) <= not((layer0_outputs(9420)) xor (layer0_outputs(12150)));
    outputs(11023) <= (layer0_outputs(1433)) xor (layer0_outputs(6290));
    outputs(11024) <= (layer0_outputs(1024)) xor (layer0_outputs(298));
    outputs(11025) <= (layer0_outputs(6679)) or (layer0_outputs(7494));
    outputs(11026) <= not(layer0_outputs(5227)) or (layer0_outputs(4654));
    outputs(11027) <= not((layer0_outputs(9363)) and (layer0_outputs(3301)));
    outputs(11028) <= not(layer0_outputs(11865));
    outputs(11029) <= not(layer0_outputs(9550));
    outputs(11030) <= not((layer0_outputs(9677)) xor (layer0_outputs(4481)));
    outputs(11031) <= (layer0_outputs(8332)) or (layer0_outputs(8584));
    outputs(11032) <= not(layer0_outputs(10284));
    outputs(11033) <= not(layer0_outputs(8061));
    outputs(11034) <= layer0_outputs(6735);
    outputs(11035) <= not((layer0_outputs(12770)) and (layer0_outputs(6379)));
    outputs(11036) <= not(layer0_outputs(3966)) or (layer0_outputs(6087));
    outputs(11037) <= not(layer0_outputs(10652));
    outputs(11038) <= (layer0_outputs(6366)) or (layer0_outputs(10167));
    outputs(11039) <= layer0_outputs(5282);
    outputs(11040) <= layer0_outputs(11367);
    outputs(11041) <= not(layer0_outputs(9689));
    outputs(11042) <= not(layer0_outputs(10879));
    outputs(11043) <= not((layer0_outputs(1786)) xor (layer0_outputs(27)));
    outputs(11044) <= not((layer0_outputs(5535)) or (layer0_outputs(10468)));
    outputs(11045) <= not((layer0_outputs(4587)) xor (layer0_outputs(9405)));
    outputs(11046) <= not((layer0_outputs(2036)) and (layer0_outputs(11676)));
    outputs(11047) <= not(layer0_outputs(5403));
    outputs(11048) <= not(layer0_outputs(3577));
    outputs(11049) <= '1';
    outputs(11050) <= layer0_outputs(6970);
    outputs(11051) <= layer0_outputs(3040);
    outputs(11052) <= not((layer0_outputs(10426)) and (layer0_outputs(1047)));
    outputs(11053) <= (layer0_outputs(12150)) or (layer0_outputs(9943));
    outputs(11054) <= not((layer0_outputs(1818)) xor (layer0_outputs(8543)));
    outputs(11055) <= not(layer0_outputs(12099));
    outputs(11056) <= not((layer0_outputs(6586)) xor (layer0_outputs(11502)));
    outputs(11057) <= not((layer0_outputs(1901)) and (layer0_outputs(12497)));
    outputs(11058) <= layer0_outputs(9069);
    outputs(11059) <= not((layer0_outputs(5888)) xor (layer0_outputs(7506)));
    outputs(11060) <= '1';
    outputs(11061) <= (layer0_outputs(4679)) xor (layer0_outputs(2128));
    outputs(11062) <= not((layer0_outputs(10693)) and (layer0_outputs(9175)));
    outputs(11063) <= not((layer0_outputs(9020)) xor (layer0_outputs(679)));
    outputs(11064) <= not(layer0_outputs(10535));
    outputs(11065) <= not(layer0_outputs(1918)) or (layer0_outputs(11552));
    outputs(11066) <= layer0_outputs(2889);
    outputs(11067) <= not((layer0_outputs(3868)) xor (layer0_outputs(9845)));
    outputs(11068) <= not((layer0_outputs(6935)) xor (layer0_outputs(1055)));
    outputs(11069) <= (layer0_outputs(6810)) or (layer0_outputs(4521));
    outputs(11070) <= layer0_outputs(4279);
    outputs(11071) <= layer0_outputs(8346);
    outputs(11072) <= not(layer0_outputs(341));
    outputs(11073) <= (layer0_outputs(12266)) or (layer0_outputs(10973));
    outputs(11074) <= (layer0_outputs(1252)) xor (layer0_outputs(512));
    outputs(11075) <= not((layer0_outputs(4730)) xor (layer0_outputs(1206)));
    outputs(11076) <= layer0_outputs(183);
    outputs(11077) <= not(layer0_outputs(2235));
    outputs(11078) <= not(layer0_outputs(2022));
    outputs(11079) <= not(layer0_outputs(10616));
    outputs(11080) <= layer0_outputs(9543);
    outputs(11081) <= (layer0_outputs(12632)) xor (layer0_outputs(5583));
    outputs(11082) <= (layer0_outputs(10895)) xor (layer0_outputs(11882));
    outputs(11083) <= layer0_outputs(538);
    outputs(11084) <= not((layer0_outputs(4792)) or (layer0_outputs(7330)));
    outputs(11085) <= not(layer0_outputs(6293));
    outputs(11086) <= not(layer0_outputs(6580));
    outputs(11087) <= not(layer0_outputs(1186));
    outputs(11088) <= layer0_outputs(7024);
    outputs(11089) <= layer0_outputs(1989);
    outputs(11090) <= (layer0_outputs(1044)) and not (layer0_outputs(1540));
    outputs(11091) <= not(layer0_outputs(7828));
    outputs(11092) <= layer0_outputs(8202);
    outputs(11093) <= not((layer0_outputs(2540)) xor (layer0_outputs(9080)));
    outputs(11094) <= not(layer0_outputs(3416));
    outputs(11095) <= (layer0_outputs(12371)) and (layer0_outputs(12107));
    outputs(11096) <= not(layer0_outputs(1538)) or (layer0_outputs(7808));
    outputs(11097) <= not(layer0_outputs(5438)) or (layer0_outputs(11386));
    outputs(11098) <= not(layer0_outputs(5509)) or (layer0_outputs(872));
    outputs(11099) <= (layer0_outputs(1711)) xor (layer0_outputs(10774));
    outputs(11100) <= not(layer0_outputs(11950));
    outputs(11101) <= (layer0_outputs(12686)) xor (layer0_outputs(6501));
    outputs(11102) <= (layer0_outputs(8782)) xor (layer0_outputs(319));
    outputs(11103) <= (layer0_outputs(79)) or (layer0_outputs(4566));
    outputs(11104) <= not((layer0_outputs(1533)) and (layer0_outputs(4366)));
    outputs(11105) <= (layer0_outputs(1213)) or (layer0_outputs(8232));
    outputs(11106) <= not((layer0_outputs(7965)) and (layer0_outputs(9062)));
    outputs(11107) <= not(layer0_outputs(12512)) or (layer0_outputs(5736));
    outputs(11108) <= layer0_outputs(4748);
    outputs(11109) <= not((layer0_outputs(10641)) xor (layer0_outputs(8858)));
    outputs(11110) <= not(layer0_outputs(2664)) or (layer0_outputs(10903));
    outputs(11111) <= layer0_outputs(6015);
    outputs(11112) <= (layer0_outputs(7331)) xor (layer0_outputs(212));
    outputs(11113) <= (layer0_outputs(6178)) or (layer0_outputs(6654));
    outputs(11114) <= (layer0_outputs(5778)) and not (layer0_outputs(5529));
    outputs(11115) <= not(layer0_outputs(6462));
    outputs(11116) <= layer0_outputs(11294);
    outputs(11117) <= layer0_outputs(2080);
    outputs(11118) <= not((layer0_outputs(2024)) or (layer0_outputs(4704)));
    outputs(11119) <= not(layer0_outputs(2975));
    outputs(11120) <= layer0_outputs(5453);
    outputs(11121) <= not((layer0_outputs(11616)) xor (layer0_outputs(8776)));
    outputs(11122) <= not(layer0_outputs(8179)) or (layer0_outputs(1517));
    outputs(11123) <= not((layer0_outputs(10083)) and (layer0_outputs(2393)));
    outputs(11124) <= (layer0_outputs(1478)) or (layer0_outputs(7283));
    outputs(11125) <= not(layer0_outputs(1406)) or (layer0_outputs(10506));
    outputs(11126) <= (layer0_outputs(2675)) and not (layer0_outputs(10937));
    outputs(11127) <= not((layer0_outputs(12643)) xor (layer0_outputs(1999)));
    outputs(11128) <= not(layer0_outputs(2914)) or (layer0_outputs(3482));
    outputs(11129) <= not((layer0_outputs(4723)) xor (layer0_outputs(3568)));
    outputs(11130) <= (layer0_outputs(1944)) xor (layer0_outputs(408));
    outputs(11131) <= (layer0_outputs(24)) xor (layer0_outputs(1453));
    outputs(11132) <= layer0_outputs(10750);
    outputs(11133) <= not((layer0_outputs(5281)) xor (layer0_outputs(1106)));
    outputs(11134) <= not(layer0_outputs(4571));
    outputs(11135) <= layer0_outputs(6974);
    outputs(11136) <= layer0_outputs(11780);
    outputs(11137) <= layer0_outputs(2903);
    outputs(11138) <= (layer0_outputs(4137)) and (layer0_outputs(5517));
    outputs(11139) <= not((layer0_outputs(7048)) xor (layer0_outputs(5984)));
    outputs(11140) <= layer0_outputs(6710);
    outputs(11141) <= layer0_outputs(1733);
    outputs(11142) <= not((layer0_outputs(8182)) xor (layer0_outputs(8640)));
    outputs(11143) <= not((layer0_outputs(7648)) xor (layer0_outputs(2270)));
    outputs(11144) <= not(layer0_outputs(5710));
    outputs(11145) <= layer0_outputs(3578);
    outputs(11146) <= layer0_outputs(12109);
    outputs(11147) <= layer0_outputs(7013);
    outputs(11148) <= layer0_outputs(11275);
    outputs(11149) <= layer0_outputs(11084);
    outputs(11150) <= not(layer0_outputs(8759));
    outputs(11151) <= layer0_outputs(12123);
    outputs(11152) <= not((layer0_outputs(8207)) xor (layer0_outputs(9239)));
    outputs(11153) <= layer0_outputs(12328);
    outputs(11154) <= not(layer0_outputs(9176));
    outputs(11155) <= not(layer0_outputs(2746));
    outputs(11156) <= layer0_outputs(1334);
    outputs(11157) <= not(layer0_outputs(8774));
    outputs(11158) <= not(layer0_outputs(4706));
    outputs(11159) <= not((layer0_outputs(7375)) or (layer0_outputs(11140)));
    outputs(11160) <= layer0_outputs(1421);
    outputs(11161) <= (layer0_outputs(12459)) and (layer0_outputs(10080));
    outputs(11162) <= (layer0_outputs(4104)) and (layer0_outputs(320));
    outputs(11163) <= (layer0_outputs(8755)) xor (layer0_outputs(1498));
    outputs(11164) <= not(layer0_outputs(10112)) or (layer0_outputs(11627));
    outputs(11165) <= not(layer0_outputs(10910)) or (layer0_outputs(4336));
    outputs(11166) <= not((layer0_outputs(6370)) or (layer0_outputs(12171)));
    outputs(11167) <= not(layer0_outputs(1237));
    outputs(11168) <= not((layer0_outputs(2915)) xor (layer0_outputs(2500)));
    outputs(11169) <= (layer0_outputs(11505)) and not (layer0_outputs(4420));
    outputs(11170) <= (layer0_outputs(522)) xor (layer0_outputs(5980));
    outputs(11171) <= not(layer0_outputs(5537));
    outputs(11172) <= (layer0_outputs(5464)) and not (layer0_outputs(10877));
    outputs(11173) <= not((layer0_outputs(4650)) xor (layer0_outputs(1619)));
    outputs(11174) <= layer0_outputs(5482);
    outputs(11175) <= (layer0_outputs(11682)) xor (layer0_outputs(6023));
    outputs(11176) <= (layer0_outputs(9704)) xor (layer0_outputs(11962));
    outputs(11177) <= not(layer0_outputs(1576));
    outputs(11178) <= layer0_outputs(10297);
    outputs(11179) <= (layer0_outputs(8406)) and (layer0_outputs(2751));
    outputs(11180) <= layer0_outputs(11513);
    outputs(11181) <= not(layer0_outputs(4887));
    outputs(11182) <= (layer0_outputs(12799)) and not (layer0_outputs(9509));
    outputs(11183) <= layer0_outputs(5378);
    outputs(11184) <= not(layer0_outputs(3434)) or (layer0_outputs(8347));
    outputs(11185) <= (layer0_outputs(10613)) or (layer0_outputs(7212));
    outputs(11186) <= not((layer0_outputs(1328)) and (layer0_outputs(11558)));
    outputs(11187) <= layer0_outputs(10518);
    outputs(11188) <= layer0_outputs(6568);
    outputs(11189) <= not(layer0_outputs(10694));
    outputs(11190) <= not((layer0_outputs(9758)) xor (layer0_outputs(4306)));
    outputs(11191) <= not(layer0_outputs(1919));
    outputs(11192) <= not(layer0_outputs(3770)) or (layer0_outputs(10170));
    outputs(11193) <= layer0_outputs(5800);
    outputs(11194) <= (layer0_outputs(2498)) xor (layer0_outputs(4591));
    outputs(11195) <= (layer0_outputs(11599)) xor (layer0_outputs(8240));
    outputs(11196) <= layer0_outputs(5476);
    outputs(11197) <= not(layer0_outputs(4944)) or (layer0_outputs(11797));
    outputs(11198) <= not((layer0_outputs(11645)) and (layer0_outputs(364)));
    outputs(11199) <= not((layer0_outputs(12022)) xor (layer0_outputs(264)));
    outputs(11200) <= layer0_outputs(10160);
    outputs(11201) <= not(layer0_outputs(12369));
    outputs(11202) <= layer0_outputs(2698);
    outputs(11203) <= layer0_outputs(884);
    outputs(11204) <= not((layer0_outputs(3519)) and (layer0_outputs(11042)));
    outputs(11205) <= not(layer0_outputs(10089)) or (layer0_outputs(9296));
    outputs(11206) <= layer0_outputs(4850);
    outputs(11207) <= layer0_outputs(1261);
    outputs(11208) <= not(layer0_outputs(3432)) or (layer0_outputs(7046));
    outputs(11209) <= not(layer0_outputs(9248));
    outputs(11210) <= not((layer0_outputs(2779)) xor (layer0_outputs(11245)));
    outputs(11211) <= layer0_outputs(12671);
    outputs(11212) <= layer0_outputs(7789);
    outputs(11213) <= (layer0_outputs(10577)) xor (layer0_outputs(4249));
    outputs(11214) <= layer0_outputs(10008);
    outputs(11215) <= layer0_outputs(6301);
    outputs(11216) <= not(layer0_outputs(1784)) or (layer0_outputs(3664));
    outputs(11217) <= (layer0_outputs(3117)) xor (layer0_outputs(3366));
    outputs(11218) <= not((layer0_outputs(12263)) xor (layer0_outputs(5046)));
    outputs(11219) <= layer0_outputs(4917);
    outputs(11220) <= layer0_outputs(329);
    outputs(11221) <= (layer0_outputs(10391)) and not (layer0_outputs(9470));
    outputs(11222) <= not((layer0_outputs(10649)) xor (layer0_outputs(1172)));
    outputs(11223) <= not(layer0_outputs(2990));
    outputs(11224) <= (layer0_outputs(12213)) or (layer0_outputs(5565));
    outputs(11225) <= not(layer0_outputs(7172));
    outputs(11226) <= (layer0_outputs(40)) xor (layer0_outputs(1813));
    outputs(11227) <= not(layer0_outputs(6394));
    outputs(11228) <= '1';
    outputs(11229) <= (layer0_outputs(11665)) and not (layer0_outputs(125));
    outputs(11230) <= not(layer0_outputs(3587));
    outputs(11231) <= not(layer0_outputs(10272));
    outputs(11232) <= not(layer0_outputs(12310));
    outputs(11233) <= (layer0_outputs(6383)) and not (layer0_outputs(8965));
    outputs(11234) <= not(layer0_outputs(7030));
    outputs(11235) <= layer0_outputs(5282);
    outputs(11236) <= not(layer0_outputs(11878));
    outputs(11237) <= layer0_outputs(7267);
    outputs(11238) <= (layer0_outputs(3995)) xor (layer0_outputs(2390));
    outputs(11239) <= not((layer0_outputs(11648)) or (layer0_outputs(1519)));
    outputs(11240) <= not((layer0_outputs(6582)) xor (layer0_outputs(4261)));
    outputs(11241) <= not((layer0_outputs(12247)) xor (layer0_outputs(11638)));
    outputs(11242) <= not((layer0_outputs(4684)) xor (layer0_outputs(8504)));
    outputs(11243) <= not(layer0_outputs(4715)) or (layer0_outputs(1933));
    outputs(11244) <= not((layer0_outputs(11500)) or (layer0_outputs(6183)));
    outputs(11245) <= not((layer0_outputs(1347)) and (layer0_outputs(4199)));
    outputs(11246) <= (layer0_outputs(7927)) xor (layer0_outputs(9207));
    outputs(11247) <= not((layer0_outputs(304)) and (layer0_outputs(905)));
    outputs(11248) <= '1';
    outputs(11249) <= not((layer0_outputs(2816)) xor (layer0_outputs(1663)));
    outputs(11250) <= (layer0_outputs(5053)) xor (layer0_outputs(8424));
    outputs(11251) <= (layer0_outputs(447)) xor (layer0_outputs(10860));
    outputs(11252) <= not(layer0_outputs(908));
    outputs(11253) <= not((layer0_outputs(4757)) xor (layer0_outputs(12636)));
    outputs(11254) <= layer0_outputs(12527);
    outputs(11255) <= (layer0_outputs(6638)) or (layer0_outputs(8667));
    outputs(11256) <= (layer0_outputs(7823)) xor (layer0_outputs(12071));
    outputs(11257) <= not((layer0_outputs(7960)) xor (layer0_outputs(131)));
    outputs(11258) <= layer0_outputs(9471);
    outputs(11259) <= (layer0_outputs(4454)) xor (layer0_outputs(9091));
    outputs(11260) <= not(layer0_outputs(4378));
    outputs(11261) <= layer0_outputs(6094);
    outputs(11262) <= not((layer0_outputs(5511)) xor (layer0_outputs(6978)));
    outputs(11263) <= not(layer0_outputs(2308)) or (layer0_outputs(12320));
    outputs(11264) <= layer0_outputs(9050);
    outputs(11265) <= not((layer0_outputs(10196)) xor (layer0_outputs(10826)));
    outputs(11266) <= not(layer0_outputs(109));
    outputs(11267) <= (layer0_outputs(2852)) xor (layer0_outputs(303));
    outputs(11268) <= layer0_outputs(7509);
    outputs(11269) <= not((layer0_outputs(9832)) and (layer0_outputs(8050)));
    outputs(11270) <= (layer0_outputs(1802)) xor (layer0_outputs(12057));
    outputs(11271) <= layer0_outputs(901);
    outputs(11272) <= (layer0_outputs(3495)) or (layer0_outputs(800));
    outputs(11273) <= not((layer0_outputs(4683)) and (layer0_outputs(6900)));
    outputs(11274) <= not(layer0_outputs(1577));
    outputs(11275) <= '0';
    outputs(11276) <= layer0_outputs(1893);
    outputs(11277) <= (layer0_outputs(12513)) and not (layer0_outputs(3783));
    outputs(11278) <= not(layer0_outputs(12243)) or (layer0_outputs(4075));
    outputs(11279) <= not((layer0_outputs(11458)) xor (layer0_outputs(10690)));
    outputs(11280) <= not((layer0_outputs(11987)) and (layer0_outputs(4673)));
    outputs(11281) <= (layer0_outputs(4518)) xor (layer0_outputs(4519));
    outputs(11282) <= (layer0_outputs(2367)) and not (layer0_outputs(7712));
    outputs(11283) <= not(layer0_outputs(10062)) or (layer0_outputs(4202));
    outputs(11284) <= not((layer0_outputs(2520)) and (layer0_outputs(6299)));
    outputs(11285) <= not((layer0_outputs(1971)) xor (layer0_outputs(9553)));
    outputs(11286) <= (layer0_outputs(5989)) xor (layer0_outputs(6802));
    outputs(11287) <= (layer0_outputs(1274)) or (layer0_outputs(10255));
    outputs(11288) <= not(layer0_outputs(10574));
    outputs(11289) <= layer0_outputs(236);
    outputs(11290) <= not(layer0_outputs(1141));
    outputs(11291) <= not(layer0_outputs(8775)) or (layer0_outputs(259));
    outputs(11292) <= (layer0_outputs(428)) and not (layer0_outputs(1524));
    outputs(11293) <= (layer0_outputs(7250)) and not (layer0_outputs(7835));
    outputs(11294) <= layer0_outputs(11582);
    outputs(11295) <= not((layer0_outputs(11136)) or (layer0_outputs(3633)));
    outputs(11296) <= layer0_outputs(6115);
    outputs(11297) <= not(layer0_outputs(10607));
    outputs(11298) <= not(layer0_outputs(8813));
    outputs(11299) <= (layer0_outputs(11658)) and not (layer0_outputs(4858));
    outputs(11300) <= (layer0_outputs(10868)) and not (layer0_outputs(9563));
    outputs(11301) <= (layer0_outputs(1926)) xor (layer0_outputs(7319));
    outputs(11302) <= not(layer0_outputs(7786));
    outputs(11303) <= (layer0_outputs(4799)) xor (layer0_outputs(1853));
    outputs(11304) <= (layer0_outputs(5237)) or (layer0_outputs(8437));
    outputs(11305) <= (layer0_outputs(12360)) or (layer0_outputs(10204));
    outputs(11306) <= layer0_outputs(12757);
    outputs(11307) <= not((layer0_outputs(4018)) and (layer0_outputs(6868)));
    outputs(11308) <= (layer0_outputs(8477)) and not (layer0_outputs(9971));
    outputs(11309) <= not(layer0_outputs(11383));
    outputs(11310) <= (layer0_outputs(11547)) xor (layer0_outputs(3054));
    outputs(11311) <= not(layer0_outputs(10673)) or (layer0_outputs(4212));
    outputs(11312) <= (layer0_outputs(10125)) xor (layer0_outputs(6785));
    outputs(11313) <= not((layer0_outputs(5840)) xor (layer0_outputs(10389)));
    outputs(11314) <= not(layer0_outputs(6665)) or (layer0_outputs(5240));
    outputs(11315) <= (layer0_outputs(7895)) and not (layer0_outputs(5032));
    outputs(11316) <= layer0_outputs(9372);
    outputs(11317) <= (layer0_outputs(12130)) xor (layer0_outputs(5017));
    outputs(11318) <= not(layer0_outputs(4664)) or (layer0_outputs(9386));
    outputs(11319) <= (layer0_outputs(11330)) and not (layer0_outputs(1278));
    outputs(11320) <= not(layer0_outputs(9089));
    outputs(11321) <= (layer0_outputs(1647)) xor (layer0_outputs(8536));
    outputs(11322) <= (layer0_outputs(5197)) and not (layer0_outputs(6228));
    outputs(11323) <= not((layer0_outputs(12497)) xor (layer0_outputs(12393)));
    outputs(11324) <= not((layer0_outputs(7355)) xor (layer0_outputs(4114)));
    outputs(11325) <= layer0_outputs(8085);
    outputs(11326) <= layer0_outputs(639);
    outputs(11327) <= (layer0_outputs(1464)) xor (layer0_outputs(7553));
    outputs(11328) <= (layer0_outputs(6858)) and not (layer0_outputs(8062));
    outputs(11329) <= (layer0_outputs(7554)) and not (layer0_outputs(7304));
    outputs(11330) <= (layer0_outputs(2376)) or (layer0_outputs(12613));
    outputs(11331) <= not((layer0_outputs(1124)) and (layer0_outputs(11881)));
    outputs(11332) <= layer0_outputs(5823);
    outputs(11333) <= layer0_outputs(7249);
    outputs(11334) <= layer0_outputs(3792);
    outputs(11335) <= not((layer0_outputs(4422)) xor (layer0_outputs(10739)));
    outputs(11336) <= (layer0_outputs(825)) or (layer0_outputs(5230));
    outputs(11337) <= not(layer0_outputs(12522));
    outputs(11338) <= not(layer0_outputs(5952));
    outputs(11339) <= (layer0_outputs(2924)) xor (layer0_outputs(5818));
    outputs(11340) <= layer0_outputs(11120);
    outputs(11341) <= not((layer0_outputs(2789)) xor (layer0_outputs(8319)));
    outputs(11342) <= (layer0_outputs(5124)) xor (layer0_outputs(4505));
    outputs(11343) <= (layer0_outputs(6931)) or (layer0_outputs(11345));
    outputs(11344) <= (layer0_outputs(2946)) xor (layer0_outputs(65));
    outputs(11345) <= not(layer0_outputs(7370)) or (layer0_outputs(1037));
    outputs(11346) <= not((layer0_outputs(9910)) and (layer0_outputs(1610)));
    outputs(11347) <= not(layer0_outputs(6262)) or (layer0_outputs(527));
    outputs(11348) <= layer0_outputs(6745);
    outputs(11349) <= layer0_outputs(5764);
    outputs(11350) <= not((layer0_outputs(883)) xor (layer0_outputs(10470)));
    outputs(11351) <= layer0_outputs(353);
    outputs(11352) <= not((layer0_outputs(10373)) xor (layer0_outputs(9871)));
    outputs(11353) <= not(layer0_outputs(9767));
    outputs(11354) <= not(layer0_outputs(9928));
    outputs(11355) <= not(layer0_outputs(8804)) or (layer0_outputs(3973));
    outputs(11356) <= layer0_outputs(787);
    outputs(11357) <= (layer0_outputs(9027)) and (layer0_outputs(5299));
    outputs(11358) <= not((layer0_outputs(10761)) xor (layer0_outputs(1292)));
    outputs(11359) <= (layer0_outputs(3753)) xor (layer0_outputs(7660));
    outputs(11360) <= not(layer0_outputs(2237)) or (layer0_outputs(6441));
    outputs(11361) <= layer0_outputs(4354);
    outputs(11362) <= layer0_outputs(9110);
    outputs(11363) <= not((layer0_outputs(7590)) xor (layer0_outputs(8391)));
    outputs(11364) <= not((layer0_outputs(4124)) xor (layer0_outputs(10187)));
    outputs(11365) <= (layer0_outputs(3889)) and not (layer0_outputs(4495));
    outputs(11366) <= layer0_outputs(8770);
    outputs(11367) <= layer0_outputs(1203);
    outputs(11368) <= not(layer0_outputs(540)) or (layer0_outputs(8288));
    outputs(11369) <= layer0_outputs(2013);
    outputs(11370) <= (layer0_outputs(262)) xor (layer0_outputs(10139));
    outputs(11371) <= not((layer0_outputs(10913)) xor (layer0_outputs(6635)));
    outputs(11372) <= not(layer0_outputs(10293)) or (layer0_outputs(11761));
    outputs(11373) <= not(layer0_outputs(2507)) or (layer0_outputs(5934));
    outputs(11374) <= (layer0_outputs(10146)) or (layer0_outputs(6908));
    outputs(11375) <= not(layer0_outputs(11626));
    outputs(11376) <= not((layer0_outputs(11321)) and (layer0_outputs(6612)));
    outputs(11377) <= not((layer0_outputs(441)) xor (layer0_outputs(4851)));
    outputs(11378) <= (layer0_outputs(2332)) or (layer0_outputs(12585));
    outputs(11379) <= not((layer0_outputs(1624)) xor (layer0_outputs(2659)));
    outputs(11380) <= not(layer0_outputs(11528));
    outputs(11381) <= not((layer0_outputs(2324)) or (layer0_outputs(4121)));
    outputs(11382) <= (layer0_outputs(5744)) xor (layer0_outputs(2045));
    outputs(11383) <= not(layer0_outputs(12503));
    outputs(11384) <= not((layer0_outputs(5)) xor (layer0_outputs(767)));
    outputs(11385) <= (layer0_outputs(5629)) xor (layer0_outputs(7015));
    outputs(11386) <= not(layer0_outputs(6590)) or (layer0_outputs(258));
    outputs(11387) <= (layer0_outputs(9918)) xor (layer0_outputs(1159));
    outputs(11388) <= not(layer0_outputs(10788));
    outputs(11389) <= (layer0_outputs(5148)) xor (layer0_outputs(8071));
    outputs(11390) <= not(layer0_outputs(4570)) or (layer0_outputs(1307));
    outputs(11391) <= not((layer0_outputs(12645)) and (layer0_outputs(12598)));
    outputs(11392) <= not(layer0_outputs(7971)) or (layer0_outputs(11058));
    outputs(11393) <= (layer0_outputs(3368)) xor (layer0_outputs(19));
    outputs(11394) <= not(layer0_outputs(5183)) or (layer0_outputs(7045));
    outputs(11395) <= not((layer0_outputs(6294)) xor (layer0_outputs(1703)));
    outputs(11396) <= (layer0_outputs(2428)) and not (layer0_outputs(10355));
    outputs(11397) <= (layer0_outputs(6861)) xor (layer0_outputs(2323));
    outputs(11398) <= layer0_outputs(5617);
    outputs(11399) <= not((layer0_outputs(1684)) xor (layer0_outputs(7613)));
    outputs(11400) <= not(layer0_outputs(11188));
    outputs(11401) <= not(layer0_outputs(6830)) or (layer0_outputs(12193));
    outputs(11402) <= not(layer0_outputs(12793)) or (layer0_outputs(10415));
    outputs(11403) <= not(layer0_outputs(6434));
    outputs(11404) <= not(layer0_outputs(4175)) or (layer0_outputs(4817));
    outputs(11405) <= (layer0_outputs(7696)) and not (layer0_outputs(10037));
    outputs(11406) <= layer0_outputs(8717);
    outputs(11407) <= (layer0_outputs(1832)) xor (layer0_outputs(11169));
    outputs(11408) <= (layer0_outputs(156)) and (layer0_outputs(9846));
    outputs(11409) <= (layer0_outputs(4497)) xor (layer0_outputs(8377));
    outputs(11410) <= layer0_outputs(3270);
    outputs(11411) <= not(layer0_outputs(1202));
    outputs(11412) <= not(layer0_outputs(671));
    outputs(11413) <= not(layer0_outputs(9030)) or (layer0_outputs(11154));
    outputs(11414) <= (layer0_outputs(3213)) and (layer0_outputs(7864));
    outputs(11415) <= not((layer0_outputs(8644)) and (layer0_outputs(8101)));
    outputs(11416) <= (layer0_outputs(2222)) xor (layer0_outputs(5678));
    outputs(11417) <= layer0_outputs(3935);
    outputs(11418) <= '1';
    outputs(11419) <= (layer0_outputs(7912)) and not (layer0_outputs(11606));
    outputs(11420) <= (layer0_outputs(11903)) xor (layer0_outputs(7966));
    outputs(11421) <= not(layer0_outputs(7325)) or (layer0_outputs(5690));
    outputs(11422) <= layer0_outputs(3664);
    outputs(11423) <= (layer0_outputs(9277)) xor (layer0_outputs(3883));
    outputs(11424) <= (layer0_outputs(3840)) or (layer0_outputs(9531));
    outputs(11425) <= not((layer0_outputs(245)) and (layer0_outputs(8471)));
    outputs(11426) <= (layer0_outputs(7017)) xor (layer0_outputs(5367));
    outputs(11427) <= layer0_outputs(9221);
    outputs(11428) <= (layer0_outputs(427)) xor (layer0_outputs(10145));
    outputs(11429) <= layer0_outputs(3045);
    outputs(11430) <= layer0_outputs(7104);
    outputs(11431) <= not((layer0_outputs(9227)) xor (layer0_outputs(10847)));
    outputs(11432) <= not(layer0_outputs(3387)) or (layer0_outputs(3988));
    outputs(11433) <= not((layer0_outputs(5410)) and (layer0_outputs(8788)));
    outputs(11434) <= not(layer0_outputs(6725));
    outputs(11435) <= (layer0_outputs(10917)) xor (layer0_outputs(12536));
    outputs(11436) <= not((layer0_outputs(4174)) xor (layer0_outputs(985)));
    outputs(11437) <= not(layer0_outputs(436));
    outputs(11438) <= (layer0_outputs(421)) or (layer0_outputs(8711));
    outputs(11439) <= not(layer0_outputs(10200)) or (layer0_outputs(9241));
    outputs(11440) <= (layer0_outputs(665)) and not (layer0_outputs(3472));
    outputs(11441) <= not(layer0_outputs(11238)) or (layer0_outputs(10985));
    outputs(11442) <= (layer0_outputs(10787)) xor (layer0_outputs(8289));
    outputs(11443) <= (layer0_outputs(1399)) xor (layer0_outputs(972));
    outputs(11444) <= (layer0_outputs(715)) and not (layer0_outputs(5280));
    outputs(11445) <= not((layer0_outputs(6766)) xor (layer0_outputs(340)));
    outputs(11446) <= not((layer0_outputs(10176)) xor (layer0_outputs(3474)));
    outputs(11447) <= layer0_outputs(2299);
    outputs(11448) <= (layer0_outputs(3699)) xor (layer0_outputs(2247));
    outputs(11449) <= (layer0_outputs(4361)) xor (layer0_outputs(2219));
    outputs(11450) <= (layer0_outputs(7272)) and not (layer0_outputs(10659));
    outputs(11451) <= not(layer0_outputs(7224)) or (layer0_outputs(11649));
    outputs(11452) <= not(layer0_outputs(11286));
    outputs(11453) <= (layer0_outputs(6431)) xor (layer0_outputs(2359));
    outputs(11454) <= layer0_outputs(2050);
    outputs(11455) <= (layer0_outputs(12359)) and not (layer0_outputs(1640));
    outputs(11456) <= (layer0_outputs(1888)) xor (layer0_outputs(3271));
    outputs(11457) <= (layer0_outputs(9697)) and not (layer0_outputs(3440));
    outputs(11458) <= not(layer0_outputs(3015)) or (layer0_outputs(10668));
    outputs(11459) <= layer0_outputs(7146);
    outputs(11460) <= not(layer0_outputs(2589)) or (layer0_outputs(7847));
    outputs(11461) <= layer0_outputs(7914);
    outputs(11462) <= (layer0_outputs(1783)) xor (layer0_outputs(4134));
    outputs(11463) <= layer0_outputs(6592);
    outputs(11464) <= not(layer0_outputs(4985));
    outputs(11465) <= (layer0_outputs(11556)) and not (layer0_outputs(11387));
    outputs(11466) <= not((layer0_outputs(10734)) xor (layer0_outputs(303)));
    outputs(11467) <= not((layer0_outputs(5915)) and (layer0_outputs(9469)));
    outputs(11468) <= layer0_outputs(4052);
    outputs(11469) <= (layer0_outputs(809)) xor (layer0_outputs(12581));
    outputs(11470) <= not(layer0_outputs(7629));
    outputs(11471) <= layer0_outputs(8780);
    outputs(11472) <= not((layer0_outputs(9234)) xor (layer0_outputs(6534)));
    outputs(11473) <= not((layer0_outputs(10180)) and (layer0_outputs(3809)));
    outputs(11474) <= layer0_outputs(10536);
    outputs(11475) <= not(layer0_outputs(6061));
    outputs(11476) <= not(layer0_outputs(4990));
    outputs(11477) <= not(layer0_outputs(5336)) or (layer0_outputs(5156));
    outputs(11478) <= not((layer0_outputs(4860)) and (layer0_outputs(11787)));
    outputs(11479) <= not((layer0_outputs(3993)) xor (layer0_outputs(5784)));
    outputs(11480) <= layer0_outputs(9970);
    outputs(11481) <= not(layer0_outputs(7354)) or (layer0_outputs(8603));
    outputs(11482) <= not((layer0_outputs(10079)) and (layer0_outputs(7762)));
    outputs(11483) <= (layer0_outputs(10164)) xor (layer0_outputs(3762));
    outputs(11484) <= (layer0_outputs(3423)) xor (layer0_outputs(11289));
    outputs(11485) <= not(layer0_outputs(5669)) or (layer0_outputs(10843));
    outputs(11486) <= not(layer0_outputs(2970));
    outputs(11487) <= not((layer0_outputs(5439)) xor (layer0_outputs(7412)));
    outputs(11488) <= layer0_outputs(6481);
    outputs(11489) <= (layer0_outputs(9589)) or (layer0_outputs(11391));
    outputs(11490) <= not(layer0_outputs(5218));
    outputs(11491) <= not(layer0_outputs(4232));
    outputs(11492) <= not(layer0_outputs(7453));
    outputs(11493) <= (layer0_outputs(6539)) and not (layer0_outputs(7820));
    outputs(11494) <= (layer0_outputs(3732)) xor (layer0_outputs(7664));
    outputs(11495) <= layer0_outputs(9677);
    outputs(11496) <= (layer0_outputs(11176)) xor (layer0_outputs(3084));
    outputs(11497) <= layer0_outputs(3768);
    outputs(11498) <= layer0_outputs(9354);
    outputs(11499) <= (layer0_outputs(1410)) or (layer0_outputs(9382));
    outputs(11500) <= layer0_outputs(8946);
    outputs(11501) <= not(layer0_outputs(12201));
    outputs(11502) <= not(layer0_outputs(6187)) or (layer0_outputs(10194));
    outputs(11503) <= not((layer0_outputs(3010)) and (layer0_outputs(4442)));
    outputs(11504) <= not(layer0_outputs(4667)) or (layer0_outputs(3174));
    outputs(11505) <= not(layer0_outputs(2203));
    outputs(11506) <= not(layer0_outputs(11866));
    outputs(11507) <= not(layer0_outputs(8390)) or (layer0_outputs(9098));
    outputs(11508) <= layer0_outputs(2621);
    outputs(11509) <= (layer0_outputs(4384)) or (layer0_outputs(6856));
    outputs(11510) <= (layer0_outputs(9410)) xor (layer0_outputs(5903));
    outputs(11511) <= layer0_outputs(4543);
    outputs(11512) <= not(layer0_outputs(11306));
    outputs(11513) <= '1';
    outputs(11514) <= not(layer0_outputs(5785));
    outputs(11515) <= not((layer0_outputs(11938)) xor (layer0_outputs(6105)));
    outputs(11516) <= (layer0_outputs(3331)) xor (layer0_outputs(4297));
    outputs(11517) <= not(layer0_outputs(8148));
    outputs(11518) <= (layer0_outputs(567)) or (layer0_outputs(7303));
    outputs(11519) <= not(layer0_outputs(8708)) or (layer0_outputs(12693));
    outputs(11520) <= not(layer0_outputs(3459));
    outputs(11521) <= layer0_outputs(3474);
    outputs(11522) <= (layer0_outputs(3555)) or (layer0_outputs(4635));
    outputs(11523) <= not(layer0_outputs(8358));
    outputs(11524) <= not((layer0_outputs(4451)) and (layer0_outputs(11608)));
    outputs(11525) <= (layer0_outputs(2114)) and not (layer0_outputs(5755));
    outputs(11526) <= layer0_outputs(10178);
    outputs(11527) <= not(layer0_outputs(1117));
    outputs(11528) <= not(layer0_outputs(8984));
    outputs(11529) <= layer0_outputs(7238);
    outputs(11530) <= not(layer0_outputs(3327));
    outputs(11531) <= not(layer0_outputs(2743)) or (layer0_outputs(11254));
    outputs(11532) <= not((layer0_outputs(9122)) or (layer0_outputs(10967)));
    outputs(11533) <= not(layer0_outputs(1243));
    outputs(11534) <= not(layer0_outputs(10030));
    outputs(11535) <= not(layer0_outputs(4979));
    outputs(11536) <= (layer0_outputs(8457)) xor (layer0_outputs(12091));
    outputs(11537) <= layer0_outputs(983);
    outputs(11538) <= not((layer0_outputs(5241)) xor (layer0_outputs(9247)));
    outputs(11539) <= (layer0_outputs(4469)) xor (layer0_outputs(11464));
    outputs(11540) <= not(layer0_outputs(5084));
    outputs(11541) <= not(layer0_outputs(4529));
    outputs(11542) <= not(layer0_outputs(6346)) or (layer0_outputs(11403));
    outputs(11543) <= (layer0_outputs(7790)) or (layer0_outputs(5396));
    outputs(11544) <= layer0_outputs(10956);
    outputs(11545) <= not((layer0_outputs(4890)) xor (layer0_outputs(7765)));
    outputs(11546) <= not((layer0_outputs(7565)) xor (layer0_outputs(1723)));
    outputs(11547) <= (layer0_outputs(10224)) and not (layer0_outputs(8361));
    outputs(11548) <= not(layer0_outputs(12172));
    outputs(11549) <= not(layer0_outputs(3105));
    outputs(11550) <= layer0_outputs(9522);
    outputs(11551) <= layer0_outputs(7266);
    outputs(11552) <= not(layer0_outputs(11303));
    outputs(11553) <= not(layer0_outputs(3588));
    outputs(11554) <= not(layer0_outputs(6828));
    outputs(11555) <= not(layer0_outputs(331));
    outputs(11556) <= (layer0_outputs(8731)) xor (layer0_outputs(6049));
    outputs(11557) <= not((layer0_outputs(12559)) xor (layer0_outputs(6180)));
    outputs(11558) <= (layer0_outputs(7450)) xor (layer0_outputs(12475));
    outputs(11559) <= not(layer0_outputs(4384));
    outputs(11560) <= (layer0_outputs(12694)) or (layer0_outputs(9844));
    outputs(11561) <= (layer0_outputs(5445)) and not (layer0_outputs(6811));
    outputs(11562) <= not((layer0_outputs(1197)) or (layer0_outputs(9991)));
    outputs(11563) <= (layer0_outputs(9461)) and not (layer0_outputs(1905));
    outputs(11564) <= (layer0_outputs(7112)) xor (layer0_outputs(8530));
    outputs(11565) <= not((layer0_outputs(12796)) or (layer0_outputs(490)));
    outputs(11566) <= not(layer0_outputs(4652));
    outputs(11567) <= not((layer0_outputs(725)) xor (layer0_outputs(886)));
    outputs(11568) <= not((layer0_outputs(11108)) xor (layer0_outputs(7193)));
    outputs(11569) <= layer0_outputs(174);
    outputs(11570) <= layer0_outputs(11383);
    outputs(11571) <= (layer0_outputs(9729)) and (layer0_outputs(954));
    outputs(11572) <= not(layer0_outputs(7515));
    outputs(11573) <= not((layer0_outputs(7123)) and (layer0_outputs(11812)));
    outputs(11574) <= (layer0_outputs(9862)) and (layer0_outputs(6086));
    outputs(11575) <= not(layer0_outputs(7854));
    outputs(11576) <= (layer0_outputs(6394)) and (layer0_outputs(6719));
    outputs(11577) <= not((layer0_outputs(3767)) xor (layer0_outputs(1690)));
    outputs(11578) <= not(layer0_outputs(917));
    outputs(11579) <= not((layer0_outputs(7230)) or (layer0_outputs(10798)));
    outputs(11580) <= (layer0_outputs(963)) xor (layer0_outputs(9181));
    outputs(11581) <= (layer0_outputs(12019)) and (layer0_outputs(5139));
    outputs(11582) <= layer0_outputs(5977);
    outputs(11583) <= (layer0_outputs(8404)) and (layer0_outputs(11066));
    outputs(11584) <= not(layer0_outputs(5684));
    outputs(11585) <= (layer0_outputs(3092)) and not (layer0_outputs(7911));
    outputs(11586) <= not((layer0_outputs(8935)) xor (layer0_outputs(3304)));
    outputs(11587) <= layer0_outputs(1978);
    outputs(11588) <= not((layer0_outputs(11348)) xor (layer0_outputs(7646)));
    outputs(11589) <= not((layer0_outputs(556)) or (layer0_outputs(3795)));
    outputs(11590) <= not(layer0_outputs(11181));
    outputs(11591) <= not(layer0_outputs(1946));
    outputs(11592) <= not(layer0_outputs(668)) or (layer0_outputs(6286));
    outputs(11593) <= not((layer0_outputs(9739)) xor (layer0_outputs(2223)));
    outputs(11594) <= (layer0_outputs(11801)) xor (layer0_outputs(11316));
    outputs(11595) <= not(layer0_outputs(3530));
    outputs(11596) <= (layer0_outputs(355)) xor (layer0_outputs(7924));
    outputs(11597) <= not(layer0_outputs(9015));
    outputs(11598) <= (layer0_outputs(4941)) and not (layer0_outputs(3841));
    outputs(11599) <= not(layer0_outputs(1355));
    outputs(11600) <= not(layer0_outputs(10389));
    outputs(11601) <= layer0_outputs(9526);
    outputs(11602) <= not(layer0_outputs(10220));
    outputs(11603) <= (layer0_outputs(11976)) xor (layer0_outputs(2132));
    outputs(11604) <= not((layer0_outputs(2844)) or (layer0_outputs(522)));
    outputs(11605) <= layer0_outputs(9348);
    outputs(11606) <= not(layer0_outputs(4742));
    outputs(11607) <= not(layer0_outputs(8348));
    outputs(11608) <= (layer0_outputs(4152)) and not (layer0_outputs(1254));
    outputs(11609) <= layer0_outputs(10305);
    outputs(11610) <= (layer0_outputs(8951)) or (layer0_outputs(3070));
    outputs(11611) <= not((layer0_outputs(1642)) xor (layer0_outputs(12094)));
    outputs(11612) <= not((layer0_outputs(3615)) xor (layer0_outputs(9172)));
    outputs(11613) <= not((layer0_outputs(8178)) or (layer0_outputs(8387)));
    outputs(11614) <= (layer0_outputs(5527)) xor (layer0_outputs(2353));
    outputs(11615) <= layer0_outputs(10753);
    outputs(11616) <= not(layer0_outputs(12285));
    outputs(11617) <= layer0_outputs(10154);
    outputs(11618) <= (layer0_outputs(10765)) and not (layer0_outputs(5757));
    outputs(11619) <= (layer0_outputs(1427)) xor (layer0_outputs(9374));
    outputs(11620) <= not((layer0_outputs(6096)) or (layer0_outputs(11970)));
    outputs(11621) <= (layer0_outputs(2504)) and not (layer0_outputs(7553));
    outputs(11622) <= (layer0_outputs(8880)) and (layer0_outputs(1272));
    outputs(11623) <= (layer0_outputs(12417)) xor (layer0_outputs(11952));
    outputs(11624) <= (layer0_outputs(6880)) and (layer0_outputs(6897));
    outputs(11625) <= not(layer0_outputs(7983));
    outputs(11626) <= not(layer0_outputs(1449));
    outputs(11627) <= not(layer0_outputs(9974));
    outputs(11628) <= not(layer0_outputs(11365));
    outputs(11629) <= not(layer0_outputs(330)) or (layer0_outputs(9862));
    outputs(11630) <= layer0_outputs(9530);
    outputs(11631) <= not(layer0_outputs(5546));
    outputs(11632) <= not(layer0_outputs(8104));
    outputs(11633) <= (layer0_outputs(9909)) or (layer0_outputs(12323));
    outputs(11634) <= not(layer0_outputs(4674));
    outputs(11635) <= (layer0_outputs(37)) xor (layer0_outputs(9662));
    outputs(11636) <= (layer0_outputs(12457)) and not (layer0_outputs(8434));
    outputs(11637) <= not(layer0_outputs(4233));
    outputs(11638) <= (layer0_outputs(11934)) and not (layer0_outputs(6107));
    outputs(11639) <= not(layer0_outputs(8114));
    outputs(11640) <= not(layer0_outputs(1408));
    outputs(11641) <= layer0_outputs(8305);
    outputs(11642) <= (layer0_outputs(130)) xor (layer0_outputs(7560));
    outputs(11643) <= not(layer0_outputs(3050));
    outputs(11644) <= (layer0_outputs(5316)) xor (layer0_outputs(4140));
    outputs(11645) <= layer0_outputs(1487);
    outputs(11646) <= layer0_outputs(479);
    outputs(11647) <= not(layer0_outputs(12059)) or (layer0_outputs(2204));
    outputs(11648) <= (layer0_outputs(1394)) xor (layer0_outputs(12519));
    outputs(11649) <= not(layer0_outputs(10727)) or (layer0_outputs(6047));
    outputs(11650) <= (layer0_outputs(4622)) and not (layer0_outputs(4050));
    outputs(11651) <= layer0_outputs(1938);
    outputs(11652) <= not(layer0_outputs(594));
    outputs(11653) <= not((layer0_outputs(8314)) or (layer0_outputs(6756)));
    outputs(11654) <= layer0_outputs(6848);
    outputs(11655) <= not(layer0_outputs(7890));
    outputs(11656) <= not(layer0_outputs(7992));
    outputs(11657) <= layer0_outputs(8343);
    outputs(11658) <= layer0_outputs(8411);
    outputs(11659) <= not((layer0_outputs(2434)) xor (layer0_outputs(11984)));
    outputs(11660) <= layer0_outputs(3044);
    outputs(11661) <= layer0_outputs(8712);
    outputs(11662) <= not((layer0_outputs(3008)) or (layer0_outputs(772)));
    outputs(11663) <= layer0_outputs(5044);
    outputs(11664) <= layer0_outputs(4047);
    outputs(11665) <= (layer0_outputs(12478)) and not (layer0_outputs(165));
    outputs(11666) <= not(layer0_outputs(4289));
    outputs(11667) <= not((layer0_outputs(3913)) or (layer0_outputs(2842)));
    outputs(11668) <= layer0_outputs(847);
    outputs(11669) <= (layer0_outputs(2261)) xor (layer0_outputs(12666));
    outputs(11670) <= (layer0_outputs(6214)) or (layer0_outputs(6188));
    outputs(11671) <= not(layer0_outputs(5562)) or (layer0_outputs(1247));
    outputs(11672) <= not(layer0_outputs(5088));
    outputs(11673) <= (layer0_outputs(3483)) and not (layer0_outputs(9090));
    outputs(11674) <= layer0_outputs(11318);
    outputs(11675) <= not(layer0_outputs(5683));
    outputs(11676) <= not(layer0_outputs(3095));
    outputs(11677) <= layer0_outputs(6436);
    outputs(11678) <= layer0_outputs(7159);
    outputs(11679) <= (layer0_outputs(4486)) and (layer0_outputs(7244));
    outputs(11680) <= layer0_outputs(11509);
    outputs(11681) <= not(layer0_outputs(4972));
    outputs(11682) <= not(layer0_outputs(41));
    outputs(11683) <= (layer0_outputs(11679)) and not (layer0_outputs(12528));
    outputs(11684) <= not((layer0_outputs(7230)) xor (layer0_outputs(8608)));
    outputs(11685) <= not((layer0_outputs(1922)) or (layer0_outputs(2002)));
    outputs(11686) <= not((layer0_outputs(2907)) xor (layer0_outputs(12603)));
    outputs(11687) <= not((layer0_outputs(4770)) and (layer0_outputs(2653)));
    outputs(11688) <= (layer0_outputs(10402)) xor (layer0_outputs(6683));
    outputs(11689) <= not((layer0_outputs(11487)) xor (layer0_outputs(5996)));
    outputs(11690) <= (layer0_outputs(10097)) and (layer0_outputs(12042));
    outputs(11691) <= layer0_outputs(2228);
    outputs(11692) <= (layer0_outputs(9436)) and not (layer0_outputs(8483));
    outputs(11693) <= not((layer0_outputs(6562)) and (layer0_outputs(2126)));
    outputs(11694) <= not(layer0_outputs(11329));
    outputs(11695) <= layer0_outputs(2747);
    outputs(11696) <= layer0_outputs(8128);
    outputs(11697) <= layer0_outputs(10890);
    outputs(11698) <= not(layer0_outputs(7954));
    outputs(11699) <= (layer0_outputs(8317)) xor (layer0_outputs(1219));
    outputs(11700) <= (layer0_outputs(76)) and not (layer0_outputs(11126));
    outputs(11701) <= (layer0_outputs(12580)) xor (layer0_outputs(9521));
    outputs(11702) <= (layer0_outputs(854)) and not (layer0_outputs(926));
    outputs(11703) <= (layer0_outputs(2747)) and (layer0_outputs(5197));
    outputs(11704) <= (layer0_outputs(11809)) and not (layer0_outputs(9790));
    outputs(11705) <= (layer0_outputs(7631)) and not (layer0_outputs(5149));
    outputs(11706) <= not(layer0_outputs(8553));
    outputs(11707) <= not(layer0_outputs(2671));
    outputs(11708) <= not((layer0_outputs(8763)) xor (layer0_outputs(9635)));
    outputs(11709) <= not(layer0_outputs(2008)) or (layer0_outputs(10267));
    outputs(11710) <= not((layer0_outputs(3934)) xor (layer0_outputs(2651)));
    outputs(11711) <= not((layer0_outputs(3987)) xor (layer0_outputs(8087)));
    outputs(11712) <= layer0_outputs(12222);
    outputs(11713) <= not(layer0_outputs(2044));
    outputs(11714) <= (layer0_outputs(2963)) and not (layer0_outputs(313));
    outputs(11715) <= layer0_outputs(732);
    outputs(11716) <= not((layer0_outputs(7271)) xor (layer0_outputs(10482)));
    outputs(11717) <= not((layer0_outputs(12048)) xor (layer0_outputs(2365)));
    outputs(11718) <= layer0_outputs(7296);
    outputs(11719) <= not((layer0_outputs(878)) xor (layer0_outputs(4692)));
    outputs(11720) <= (layer0_outputs(6763)) and not (layer0_outputs(3019));
    outputs(11721) <= not(layer0_outputs(4172)) or (layer0_outputs(7838));
    outputs(11722) <= not((layer0_outputs(4032)) xor (layer0_outputs(1560)));
    outputs(11723) <= layer0_outputs(5079);
    outputs(11724) <= not((layer0_outputs(6033)) or (layer0_outputs(953)));
    outputs(11725) <= (layer0_outputs(7327)) and not (layer0_outputs(4766));
    outputs(11726) <= (layer0_outputs(4894)) and (layer0_outputs(11880));
    outputs(11727) <= not((layer0_outputs(11021)) or (layer0_outputs(3224)));
    outputs(11728) <= (layer0_outputs(1746)) xor (layer0_outputs(3637));
    outputs(11729) <= not(layer0_outputs(3995));
    outputs(11730) <= not((layer0_outputs(10636)) or (layer0_outputs(8032)));
    outputs(11731) <= layer0_outputs(5113);
    outputs(11732) <= not((layer0_outputs(12549)) or (layer0_outputs(6443)));
    outputs(11733) <= not(layer0_outputs(2628));
    outputs(11734) <= (layer0_outputs(6318)) and not (layer0_outputs(9727));
    outputs(11735) <= (layer0_outputs(6516)) and (layer0_outputs(7403));
    outputs(11736) <= (layer0_outputs(8449)) and (layer0_outputs(7929));
    outputs(11737) <= not(layer0_outputs(5721)) or (layer0_outputs(8734));
    outputs(11738) <= not((layer0_outputs(6666)) xor (layer0_outputs(8677)));
    outputs(11739) <= layer0_outputs(8407);
    outputs(11740) <= (layer0_outputs(8629)) or (layer0_outputs(8515));
    outputs(11741) <= (layer0_outputs(12562)) and not (layer0_outputs(9182));
    outputs(11742) <= not(layer0_outputs(2498));
    outputs(11743) <= layer0_outputs(12366);
    outputs(11744) <= (layer0_outputs(4987)) and not (layer0_outputs(7655));
    outputs(11745) <= layer0_outputs(9459);
    outputs(11746) <= not((layer0_outputs(10475)) xor (layer0_outputs(593)));
    outputs(11747) <= not((layer0_outputs(11858)) or (layer0_outputs(149)));
    outputs(11748) <= (layer0_outputs(4363)) and not (layer0_outputs(7194));
    outputs(11749) <= layer0_outputs(555);
    outputs(11750) <= (layer0_outputs(10129)) and (layer0_outputs(7068));
    outputs(11751) <= not(layer0_outputs(2524));
    outputs(11752) <= not(layer0_outputs(7273));
    outputs(11753) <= (layer0_outputs(8005)) xor (layer0_outputs(10828));
    outputs(11754) <= (layer0_outputs(11708)) and (layer0_outputs(7454));
    outputs(11755) <= layer0_outputs(8704);
    outputs(11756) <= (layer0_outputs(3733)) and (layer0_outputs(5662));
    outputs(11757) <= (layer0_outputs(2837)) xor (layer0_outputs(439));
    outputs(11758) <= (layer0_outputs(2020)) and not (layer0_outputs(3188));
    outputs(11759) <= layer0_outputs(7326);
    outputs(11760) <= layer0_outputs(706);
    outputs(11761) <= not(layer0_outputs(10357));
    outputs(11762) <= not(layer0_outputs(4076));
    outputs(11763) <= (layer0_outputs(2981)) and not (layer0_outputs(9137));
    outputs(11764) <= not(layer0_outputs(9067));
    outputs(11765) <= not(layer0_outputs(7666));
    outputs(11766) <= layer0_outputs(10508);
    outputs(11767) <= not((layer0_outputs(5791)) xor (layer0_outputs(9852)));
    outputs(11768) <= (layer0_outputs(4889)) xor (layer0_outputs(2386));
    outputs(11769) <= not(layer0_outputs(10311));
    outputs(11770) <= not((layer0_outputs(483)) xor (layer0_outputs(1753)));
    outputs(11771) <= layer0_outputs(3933);
    outputs(11772) <= not(layer0_outputs(184));
    outputs(11773) <= layer0_outputs(6336);
    outputs(11774) <= layer0_outputs(43);
    outputs(11775) <= not(layer0_outputs(1742));
    outputs(11776) <= layer0_outputs(11409);
    outputs(11777) <= not(layer0_outputs(15));
    outputs(11778) <= (layer0_outputs(12781)) xor (layer0_outputs(10474));
    outputs(11779) <= (layer0_outputs(9928)) and not (layer0_outputs(1289));
    outputs(11780) <= not(layer0_outputs(11759));
    outputs(11781) <= (layer0_outputs(7987)) or (layer0_outputs(4546));
    outputs(11782) <= not(layer0_outputs(11501));
    outputs(11783) <= layer0_outputs(5474);
    outputs(11784) <= (layer0_outputs(959)) and not (layer0_outputs(6808));
    outputs(11785) <= not(layer0_outputs(1052));
    outputs(11786) <= (layer0_outputs(7311)) or (layer0_outputs(7015));
    outputs(11787) <= not((layer0_outputs(1352)) xor (layer0_outputs(6161)));
    outputs(11788) <= (layer0_outputs(10064)) and (layer0_outputs(6468));
    outputs(11789) <= not(layer0_outputs(2944)) or (layer0_outputs(7718));
    outputs(11790) <= not((layer0_outputs(2947)) xor (layer0_outputs(3548)));
    outputs(11791) <= layer0_outputs(6457);
    outputs(11792) <= not(layer0_outputs(8508));
    outputs(11793) <= not(layer0_outputs(4280));
    outputs(11794) <= not(layer0_outputs(9195));
    outputs(11795) <= not(layer0_outputs(4744)) or (layer0_outputs(909));
    outputs(11796) <= layer0_outputs(11294);
    outputs(11797) <= '1';
    outputs(11798) <= layer0_outputs(4814);
    outputs(11799) <= not(layer0_outputs(9398));
    outputs(11800) <= not(layer0_outputs(2870));
    outputs(11801) <= layer0_outputs(3698);
    outputs(11802) <= layer0_outputs(9693);
    outputs(11803) <= not(layer0_outputs(3843));
    outputs(11804) <= not(layer0_outputs(8917));
    outputs(11805) <= layer0_outputs(9522);
    outputs(11806) <= not(layer0_outputs(9206));
    outputs(11807) <= (layer0_outputs(12362)) and (layer0_outputs(9024));
    outputs(11808) <= layer0_outputs(226);
    outputs(11809) <= not(layer0_outputs(6218)) or (layer0_outputs(6745));
    outputs(11810) <= not((layer0_outputs(4355)) xor (layer0_outputs(5429)));
    outputs(11811) <= not(layer0_outputs(3923));
    outputs(11812) <= (layer0_outputs(2547)) and not (layer0_outputs(11376));
    outputs(11813) <= (layer0_outputs(1342)) and (layer0_outputs(11661));
    outputs(11814) <= (layer0_outputs(3365)) and not (layer0_outputs(6975));
    outputs(11815) <= layer0_outputs(4935);
    outputs(11816) <= (layer0_outputs(11845)) and not (layer0_outputs(7610));
    outputs(11817) <= layer0_outputs(3888);
    outputs(11818) <= (layer0_outputs(4092)) or (layer0_outputs(312));
    outputs(11819) <= layer0_outputs(8329);
    outputs(11820) <= (layer0_outputs(7816)) xor (layer0_outputs(5760));
    outputs(11821) <= not(layer0_outputs(11609));
    outputs(11822) <= not(layer0_outputs(2922));
    outputs(11823) <= not((layer0_outputs(727)) xor (layer0_outputs(9873)));
    outputs(11824) <= not(layer0_outputs(2906));
    outputs(11825) <= layer0_outputs(3091);
    outputs(11826) <= (layer0_outputs(5986)) xor (layer0_outputs(5176));
    outputs(11827) <= layer0_outputs(3492);
    outputs(11828) <= (layer0_outputs(1356)) and not (layer0_outputs(5107));
    outputs(11829) <= (layer0_outputs(1128)) and not (layer0_outputs(6010));
    outputs(11830) <= not((layer0_outputs(5267)) xor (layer0_outputs(10407)));
    outputs(11831) <= (layer0_outputs(11353)) xor (layer0_outputs(4951));
    outputs(11832) <= not(layer0_outputs(4536));
    outputs(11833) <= not((layer0_outputs(10203)) xor (layer0_outputs(3656)));
    outputs(11834) <= not(layer0_outputs(5431));
    outputs(11835) <= not(layer0_outputs(6905));
    outputs(11836) <= not((layer0_outputs(12517)) or (layer0_outputs(6230)));
    outputs(11837) <= not((layer0_outputs(6105)) xor (layer0_outputs(4736)));
    outputs(11838) <= (layer0_outputs(5739)) and not (layer0_outputs(2874));
    outputs(11839) <= (layer0_outputs(8661)) xor (layer0_outputs(1601));
    outputs(11840) <= not(layer0_outputs(9340));
    outputs(11841) <= not(layer0_outputs(511));
    outputs(11842) <= (layer0_outputs(5717)) and (layer0_outputs(3980));
    outputs(11843) <= not(layer0_outputs(10876));
    outputs(11844) <= (layer0_outputs(11905)) and not (layer0_outputs(1669));
    outputs(11845) <= not((layer0_outputs(6793)) xor (layer0_outputs(10029)));
    outputs(11846) <= (layer0_outputs(12066)) and (layer0_outputs(7757));
    outputs(11847) <= not(layer0_outputs(7376));
    outputs(11848) <= (layer0_outputs(5774)) or (layer0_outputs(2882));
    outputs(11849) <= (layer0_outputs(1712)) xor (layer0_outputs(3369));
    outputs(11850) <= not(layer0_outputs(8719));
    outputs(11851) <= (layer0_outputs(12506)) xor (layer0_outputs(7218));
    outputs(11852) <= not(layer0_outputs(12413));
    outputs(11853) <= not(layer0_outputs(9406)) or (layer0_outputs(10215));
    outputs(11854) <= (layer0_outputs(4379)) and not (layer0_outputs(5134));
    outputs(11855) <= (layer0_outputs(10096)) and not (layer0_outputs(10512));
    outputs(11856) <= layer0_outputs(1979);
    outputs(11857) <= layer0_outputs(1093);
    outputs(11858) <= not(layer0_outputs(11424));
    outputs(11859) <= not(layer0_outputs(9891));
    outputs(11860) <= (layer0_outputs(699)) and (layer0_outputs(10036));
    outputs(11861) <= layer0_outputs(4046);
    outputs(11862) <= not((layer0_outputs(2005)) xor (layer0_outputs(4431)));
    outputs(11863) <= not(layer0_outputs(10041));
    outputs(11864) <= (layer0_outputs(4567)) xor (layer0_outputs(2088));
    outputs(11865) <= not((layer0_outputs(2668)) xor (layer0_outputs(4572)));
    outputs(11866) <= (layer0_outputs(5097)) and not (layer0_outputs(6693));
    outputs(11867) <= layer0_outputs(8310);
    outputs(11868) <= layer0_outputs(1803);
    outputs(11869) <= (layer0_outputs(6657)) xor (layer0_outputs(5764));
    outputs(11870) <= layer0_outputs(4686);
    outputs(11871) <= (layer0_outputs(81)) and not (layer0_outputs(12724));
    outputs(11872) <= not(layer0_outputs(11100));
    outputs(11873) <= (layer0_outputs(520)) or (layer0_outputs(8746));
    outputs(11874) <= not((layer0_outputs(2708)) xor (layer0_outputs(4334)));
    outputs(11875) <= (layer0_outputs(9875)) and not (layer0_outputs(6526));
    outputs(11876) <= not((layer0_outputs(4826)) xor (layer0_outputs(9739)));
    outputs(11877) <= not(layer0_outputs(4313));
    outputs(11878) <= not((layer0_outputs(640)) xor (layer0_outputs(7483)));
    outputs(11879) <= not(layer0_outputs(11452));
    outputs(11880) <= not(layer0_outputs(12794));
    outputs(11881) <= layer0_outputs(3528);
    outputs(11882) <= not((layer0_outputs(7775)) xor (layer0_outputs(10965)));
    outputs(11883) <= (layer0_outputs(7040)) and (layer0_outputs(9036));
    outputs(11884) <= (layer0_outputs(525)) and (layer0_outputs(7411));
    outputs(11885) <= not(layer0_outputs(3189));
    outputs(11886) <= (layer0_outputs(6598)) and not (layer0_outputs(398));
    outputs(11887) <= not(layer0_outputs(12655));
    outputs(11888) <= not((layer0_outputs(10371)) or (layer0_outputs(8811)));
    outputs(11889) <= not((layer0_outputs(12166)) xor (layer0_outputs(3438)));
    outputs(11890) <= (layer0_outputs(8913)) xor (layer0_outputs(3248));
    outputs(11891) <= (layer0_outputs(6068)) and not (layer0_outputs(12061));
    outputs(11892) <= not(layer0_outputs(9657));
    outputs(11893) <= layer0_outputs(9279);
    outputs(11894) <= not((layer0_outputs(11142)) xor (layer0_outputs(6487)));
    outputs(11895) <= (layer0_outputs(11595)) xor (layer0_outputs(3162));
    outputs(11896) <= not((layer0_outputs(8219)) xor (layer0_outputs(5220)));
    outputs(11897) <= not((layer0_outputs(8320)) xor (layer0_outputs(2305)));
    outputs(11898) <= not(layer0_outputs(4434));
    outputs(11899) <= (layer0_outputs(9321)) and not (layer0_outputs(6990));
    outputs(11900) <= not(layer0_outputs(11937));
    outputs(11901) <= (layer0_outputs(9021)) xor (layer0_outputs(11301));
    outputs(11902) <= not((layer0_outputs(6466)) xor (layer0_outputs(7432)));
    outputs(11903) <= (layer0_outputs(6046)) xor (layer0_outputs(2091));
    outputs(11904) <= layer0_outputs(6572);
    outputs(11905) <= not((layer0_outputs(2133)) or (layer0_outputs(4933)));
    outputs(11906) <= (layer0_outputs(11234)) xor (layer0_outputs(8492));
    outputs(11907) <= layer0_outputs(4331);
    outputs(11908) <= not((layer0_outputs(7680)) xor (layer0_outputs(8350)));
    outputs(11909) <= not(layer0_outputs(10732));
    outputs(11910) <= not((layer0_outputs(12691)) xor (layer0_outputs(5415)));
    outputs(11911) <= (layer0_outputs(11304)) xor (layer0_outputs(9813));
    outputs(11912) <= not((layer0_outputs(3703)) xor (layer0_outputs(5316)));
    outputs(11913) <= layer0_outputs(12232);
    outputs(11914) <= layer0_outputs(3655);
    outputs(11915) <= not((layer0_outputs(4511)) xor (layer0_outputs(11095)));
    outputs(11916) <= not(layer0_outputs(1656));
    outputs(11917) <= (layer0_outputs(4819)) and not (layer0_outputs(7305));
    outputs(11918) <= not((layer0_outputs(7593)) xor (layer0_outputs(1491)));
    outputs(11919) <= layer0_outputs(7274);
    outputs(11920) <= (layer0_outputs(532)) xor (layer0_outputs(12756));
    outputs(11921) <= layer0_outputs(10960);
    outputs(11922) <= not(layer0_outputs(10343));
    outputs(11923) <= (layer0_outputs(4815)) xor (layer0_outputs(3804));
    outputs(11924) <= not(layer0_outputs(9327));
    outputs(11925) <= (layer0_outputs(9447)) and not (layer0_outputs(2307));
    outputs(11926) <= (layer0_outputs(11951)) xor (layer0_outputs(5062));
    outputs(11927) <= not(layer0_outputs(3610));
    outputs(11928) <= not(layer0_outputs(10836));
    outputs(11929) <= (layer0_outputs(4733)) xor (layer0_outputs(5029));
    outputs(11930) <= layer0_outputs(7936);
    outputs(11931) <= layer0_outputs(11210);
    outputs(11932) <= (layer0_outputs(6074)) xor (layer0_outputs(5637));
    outputs(11933) <= layer0_outputs(9685);
    outputs(11934) <= not((layer0_outputs(3632)) or (layer0_outputs(8243)));
    outputs(11935) <= not(layer0_outputs(10896));
    outputs(11936) <= (layer0_outputs(5564)) and not (layer0_outputs(7233));
    outputs(11937) <= (layer0_outputs(3790)) and not (layer0_outputs(4488));
    outputs(11938) <= (layer0_outputs(2164)) or (layer0_outputs(10752));
    outputs(11939) <= not(layer0_outputs(3718));
    outputs(11940) <= not((layer0_outputs(8518)) xor (layer0_outputs(6172)));
    outputs(11941) <= not(layer0_outputs(6494));
    outputs(11942) <= not(layer0_outputs(4784)) or (layer0_outputs(11344));
    outputs(11943) <= layer0_outputs(12594);
    outputs(11944) <= not(layer0_outputs(10648)) or (layer0_outputs(10504));
    outputs(11945) <= not(layer0_outputs(11419));
    outputs(11946) <= not(layer0_outputs(3435));
    outputs(11947) <= not(layer0_outputs(716));
    outputs(11948) <= layer0_outputs(1418);
    outputs(11949) <= (layer0_outputs(11146)) and (layer0_outputs(199));
    outputs(11950) <= not((layer0_outputs(9527)) or (layer0_outputs(3138)));
    outputs(11951) <= not(layer0_outputs(4771));
    outputs(11952) <= (layer0_outputs(1443)) xor (layer0_outputs(11128));
    outputs(11953) <= layer0_outputs(11258);
    outputs(11954) <= layer0_outputs(10960);
    outputs(11955) <= not((layer0_outputs(7439)) or (layer0_outputs(3619)));
    outputs(11956) <= not(layer0_outputs(1822));
    outputs(11957) <= not((layer0_outputs(12612)) xor (layer0_outputs(7259)));
    outputs(11958) <= (layer0_outputs(636)) and not (layer0_outputs(9959));
    outputs(11959) <= not(layer0_outputs(9609));
    outputs(11960) <= layer0_outputs(2006);
    outputs(11961) <= layer0_outputs(11640);
    outputs(11962) <= not((layer0_outputs(10220)) or (layer0_outputs(5727)));
    outputs(11963) <= layer0_outputs(11003);
    outputs(11964) <= not((layer0_outputs(7603)) xor (layer0_outputs(10407)));
    outputs(11965) <= not(layer0_outputs(1700));
    outputs(11966) <= not(layer0_outputs(3410)) or (layer0_outputs(9252));
    outputs(11967) <= layer0_outputs(11944);
    outputs(11968) <= not((layer0_outputs(11955)) xor (layer0_outputs(3238)));
    outputs(11969) <= not((layer0_outputs(2853)) or (layer0_outputs(11888)));
    outputs(11970) <= (layer0_outputs(9274)) and not (layer0_outputs(8368));
    outputs(11971) <= not((layer0_outputs(6108)) xor (layer0_outputs(1542)));
    outputs(11972) <= not(layer0_outputs(7148));
    outputs(11973) <= not(layer0_outputs(6633));
    outputs(11974) <= (layer0_outputs(12730)) xor (layer0_outputs(4934));
    outputs(11975) <= (layer0_outputs(6685)) and not (layer0_outputs(5130));
    outputs(11976) <= not(layer0_outputs(1204));
    outputs(11977) <= not((layer0_outputs(1185)) xor (layer0_outputs(11955)));
    outputs(11978) <= not((layer0_outputs(3872)) or (layer0_outputs(761)));
    outputs(11979) <= not(layer0_outputs(8984));
    outputs(11980) <= not(layer0_outputs(11181));
    outputs(11981) <= not(layer0_outputs(221));
    outputs(11982) <= not(layer0_outputs(5221));
    outputs(11983) <= layer0_outputs(3297);
    outputs(11984) <= layer0_outputs(11838);
    outputs(11985) <= (layer0_outputs(4304)) xor (layer0_outputs(7870));
    outputs(11986) <= '0';
    outputs(11987) <= not((layer0_outputs(11274)) xor (layer0_outputs(10730)));
    outputs(11988) <= not(layer0_outputs(10542)) or (layer0_outputs(2290));
    outputs(11989) <= not(layer0_outputs(866));
    outputs(11990) <= not(layer0_outputs(10554));
    outputs(11991) <= layer0_outputs(11210);
    outputs(11992) <= layer0_outputs(825);
    outputs(11993) <= (layer0_outputs(2007)) and not (layer0_outputs(4150));
    outputs(11994) <= not(layer0_outputs(7180));
    outputs(11995) <= (layer0_outputs(8026)) and not (layer0_outputs(11580));
    outputs(11996) <= not((layer0_outputs(1159)) or (layer0_outputs(11036)));
    outputs(11997) <= not(layer0_outputs(2689));
    outputs(11998) <= layer0_outputs(9278);
    outputs(11999) <= layer0_outputs(9096);
    outputs(12000) <= (layer0_outputs(2303)) and (layer0_outputs(8211));
    outputs(12001) <= not((layer0_outputs(2546)) xor (layer0_outputs(1225)));
    outputs(12002) <= (layer0_outputs(2135)) xor (layer0_outputs(4485));
    outputs(12003) <= not(layer0_outputs(10630));
    outputs(12004) <= not(layer0_outputs(8592));
    outputs(12005) <= not((layer0_outputs(3775)) xor (layer0_outputs(2553)));
    outputs(12006) <= (layer0_outputs(641)) and (layer0_outputs(5964));
    outputs(12007) <= (layer0_outputs(7101)) xor (layer0_outputs(1057));
    outputs(12008) <= (layer0_outputs(9161)) xor (layer0_outputs(7439));
    outputs(12009) <= (layer0_outputs(11546)) and not (layer0_outputs(1920));
    outputs(12010) <= (layer0_outputs(4238)) and (layer0_outputs(8562));
    outputs(12011) <= not((layer0_outputs(11800)) xor (layer0_outputs(7644)));
    outputs(12012) <= (layer0_outputs(10716)) and not (layer0_outputs(1660));
    outputs(12013) <= (layer0_outputs(3426)) and (layer0_outputs(3549));
    outputs(12014) <= layer0_outputs(2292);
    outputs(12015) <= layer0_outputs(6641);
    outputs(12016) <= layer0_outputs(7817);
    outputs(12017) <= not((layer0_outputs(5136)) xor (layer0_outputs(5195)));
    outputs(12018) <= not((layer0_outputs(458)) xor (layer0_outputs(2195)));
    outputs(12019) <= not(layer0_outputs(491)) or (layer0_outputs(2189));
    outputs(12020) <= not(layer0_outputs(11741));
    outputs(12021) <= not(layer0_outputs(9848));
    outputs(12022) <= layer0_outputs(1735);
    outputs(12023) <= not((layer0_outputs(4168)) xor (layer0_outputs(10773)));
    outputs(12024) <= (layer0_outputs(2063)) and (layer0_outputs(1791));
    outputs(12025) <= not((layer0_outputs(10513)) xor (layer0_outputs(5946)));
    outputs(12026) <= layer0_outputs(11426);
    outputs(12027) <= not(layer0_outputs(896));
    outputs(12028) <= not((layer0_outputs(1641)) or (layer0_outputs(191)));
    outputs(12029) <= (layer0_outputs(10027)) and not (layer0_outputs(7882));
    outputs(12030) <= (layer0_outputs(9795)) and not (layer0_outputs(4695));
    outputs(12031) <= not(layer0_outputs(5575));
    outputs(12032) <= (layer0_outputs(8098)) xor (layer0_outputs(4528));
    outputs(12033) <= not(layer0_outputs(9771));
    outputs(12034) <= not(layer0_outputs(2987));
    outputs(12035) <= not(layer0_outputs(2509)) or (layer0_outputs(7796));
    outputs(12036) <= not(layer0_outputs(9401));
    outputs(12037) <= layer0_outputs(10238);
    outputs(12038) <= not((layer0_outputs(429)) xor (layer0_outputs(5605)));
    outputs(12039) <= layer0_outputs(7567);
    outputs(12040) <= not(layer0_outputs(7527));
    outputs(12041) <= not((layer0_outputs(5353)) and (layer0_outputs(12220)));
    outputs(12042) <= layer0_outputs(7332);
    outputs(12043) <= not(layer0_outputs(7610));
    outputs(12044) <= not(layer0_outputs(7957));
    outputs(12045) <= (layer0_outputs(12744)) xor (layer0_outputs(4048));
    outputs(12046) <= (layer0_outputs(713)) xor (layer0_outputs(4524));
    outputs(12047) <= (layer0_outputs(6125)) xor (layer0_outputs(3592));
    outputs(12048) <= (layer0_outputs(5251)) and (layer0_outputs(10820));
    outputs(12049) <= layer0_outputs(681);
    outputs(12050) <= not(layer0_outputs(6854));
    outputs(12051) <= not((layer0_outputs(1608)) xor (layer0_outputs(3498)));
    outputs(12052) <= layer0_outputs(6576);
    outputs(12053) <= not(layer0_outputs(247)) or (layer0_outputs(10806));
    outputs(12054) <= not((layer0_outputs(5863)) or (layer0_outputs(9747)));
    outputs(12055) <= (layer0_outputs(12448)) and (layer0_outputs(12739));
    outputs(12056) <= not(layer0_outputs(7302));
    outputs(12057) <= layer0_outputs(17);
    outputs(12058) <= not(layer0_outputs(8705));
    outputs(12059) <= not(layer0_outputs(10268));
    outputs(12060) <= layer0_outputs(319);
    outputs(12061) <= layer0_outputs(7310);
    outputs(12062) <= layer0_outputs(2052);
    outputs(12063) <= (layer0_outputs(4179)) xor (layer0_outputs(4975));
    outputs(12064) <= (layer0_outputs(6360)) and not (layer0_outputs(8525));
    outputs(12065) <= not((layer0_outputs(7464)) xor (layer0_outputs(11730)));
    outputs(12066) <= layer0_outputs(12297);
    outputs(12067) <= not(layer0_outputs(8540));
    outputs(12068) <= not(layer0_outputs(273));
    outputs(12069) <= (layer0_outputs(10398)) xor (layer0_outputs(9867));
    outputs(12070) <= not(layer0_outputs(2379));
    outputs(12071) <= layer0_outputs(10504);
    outputs(12072) <= layer0_outputs(2110);
    outputs(12073) <= not(layer0_outputs(4100));
    outputs(12074) <= not((layer0_outputs(9031)) xor (layer0_outputs(2868)));
    outputs(12075) <= (layer0_outputs(7696)) xor (layer0_outputs(11311));
    outputs(12076) <= not(layer0_outputs(2473));
    outputs(12077) <= (layer0_outputs(7203)) xor (layer0_outputs(106));
    outputs(12078) <= not((layer0_outputs(5597)) xor (layer0_outputs(9541)));
    outputs(12079) <= not(layer0_outputs(11064));
    outputs(12080) <= layer0_outputs(5075);
    outputs(12081) <= not(layer0_outputs(7164));
    outputs(12082) <= (layer0_outputs(2055)) xor (layer0_outputs(4138));
    outputs(12083) <= (layer0_outputs(1065)) xor (layer0_outputs(6490));
    outputs(12084) <= (layer0_outputs(3997)) and not (layer0_outputs(5022));
    outputs(12085) <= (layer0_outputs(1866)) xor (layer0_outputs(2070));
    outputs(12086) <= not((layer0_outputs(11882)) xor (layer0_outputs(1400)));
    outputs(12087) <= not((layer0_outputs(2752)) or (layer0_outputs(5472)));
    outputs(12088) <= (layer0_outputs(3232)) and (layer0_outputs(814));
    outputs(12089) <= not(layer0_outputs(11600)) or (layer0_outputs(11426));
    outputs(12090) <= layer0_outputs(286);
    outputs(12091) <= (layer0_outputs(1173)) and not (layer0_outputs(3284));
    outputs(12092) <= not((layer0_outputs(3093)) and (layer0_outputs(119)));
    outputs(12093) <= not(layer0_outputs(12309));
    outputs(12094) <= layer0_outputs(6360);
    outputs(12095) <= not((layer0_outputs(1002)) and (layer0_outputs(727)));
    outputs(12096) <= (layer0_outputs(5694)) and (layer0_outputs(1328));
    outputs(12097) <= (layer0_outputs(4859)) and not (layer0_outputs(9335));
    outputs(12098) <= (layer0_outputs(8098)) and (layer0_outputs(441));
    outputs(12099) <= (layer0_outputs(7168)) xor (layer0_outputs(8699));
    outputs(12100) <= not((layer0_outputs(6173)) xor (layer0_outputs(6455)));
    outputs(12101) <= layer0_outputs(478);
    outputs(12102) <= not(layer0_outputs(4914));
    outputs(12103) <= not(layer0_outputs(1123));
    outputs(12104) <= (layer0_outputs(2394)) and not (layer0_outputs(12163));
    outputs(12105) <= not((layer0_outputs(3564)) and (layer0_outputs(5317)));
    outputs(12106) <= not((layer0_outputs(1043)) or (layer0_outputs(10289)));
    outputs(12107) <= (layer0_outputs(306)) and (layer0_outputs(4965));
    outputs(12108) <= not((layer0_outputs(731)) xor (layer0_outputs(2554)));
    outputs(12109) <= (layer0_outputs(2273)) and not (layer0_outputs(3401));
    outputs(12110) <= not(layer0_outputs(3831));
    outputs(12111) <= not(layer0_outputs(7821));
    outputs(12112) <= (layer0_outputs(11414)) xor (layer0_outputs(123));
    outputs(12113) <= not(layer0_outputs(7401));
    outputs(12114) <= (layer0_outputs(93)) xor (layer0_outputs(9983));
    outputs(12115) <= layer0_outputs(2165);
    outputs(12116) <= not(layer0_outputs(12648));
    outputs(12117) <= not(layer0_outputs(5836));
    outputs(12118) <= not(layer0_outputs(9025));
    outputs(12119) <= not((layer0_outputs(4854)) xor (layer0_outputs(5918)));
    outputs(12120) <= layer0_outputs(6818);
    outputs(12121) <= not(layer0_outputs(29));
    outputs(12122) <= not(layer0_outputs(9720));
    outputs(12123) <= not((layer0_outputs(12013)) and (layer0_outputs(6705)));
    outputs(12124) <= not(layer0_outputs(4534));
    outputs(12125) <= not(layer0_outputs(6682));
    outputs(12126) <= not((layer0_outputs(3838)) or (layer0_outputs(10056)));
    outputs(12127) <= layer0_outputs(7562);
    outputs(12128) <= not(layer0_outputs(8968));
    outputs(12129) <= not((layer0_outputs(4781)) or (layer0_outputs(10134)));
    outputs(12130) <= not((layer0_outputs(2558)) or (layer0_outputs(1441)));
    outputs(12131) <= not(layer0_outputs(107));
    outputs(12132) <= not(layer0_outputs(11285));
    outputs(12133) <= not(layer0_outputs(196));
    outputs(12134) <= layer0_outputs(12591);
    outputs(12135) <= not((layer0_outputs(12046)) and (layer0_outputs(12286)));
    outputs(12136) <= (layer0_outputs(5321)) and not (layer0_outputs(2794));
    outputs(12137) <= not((layer0_outputs(7065)) xor (layer0_outputs(2484)));
    outputs(12138) <= not((layer0_outputs(746)) xor (layer0_outputs(12157)));
    outputs(12139) <= layer0_outputs(656);
    outputs(12140) <= (layer0_outputs(5488)) xor (layer0_outputs(3185));
    outputs(12141) <= (layer0_outputs(10367)) or (layer0_outputs(6421));
    outputs(12142) <= not(layer0_outputs(7751));
    outputs(12143) <= layer0_outputs(6512);
    outputs(12144) <= (layer0_outputs(10814)) xor (layer0_outputs(6557));
    outputs(12145) <= layer0_outputs(12691);
    outputs(12146) <= not(layer0_outputs(11619));
    outputs(12147) <= not(layer0_outputs(7234));
    outputs(12148) <= not(layer0_outputs(9586));
    outputs(12149) <= (layer0_outputs(12110)) xor (layer0_outputs(11463));
    outputs(12150) <= (layer0_outputs(381)) and not (layer0_outputs(4593));
    outputs(12151) <= (layer0_outputs(7472)) and not (layer0_outputs(9718));
    outputs(12152) <= layer0_outputs(2629);
    outputs(12153) <= (layer0_outputs(3034)) and (layer0_outputs(10087));
    outputs(12154) <= (layer0_outputs(9590)) xor (layer0_outputs(2671));
    outputs(12155) <= not(layer0_outputs(7127));
    outputs(12156) <= not((layer0_outputs(7722)) xor (layer0_outputs(2506)));
    outputs(12157) <= not(layer0_outputs(4));
    outputs(12158) <= (layer0_outputs(5021)) and (layer0_outputs(1939));
    outputs(12159) <= not((layer0_outputs(4874)) xor (layer0_outputs(1858)));
    outputs(12160) <= layer0_outputs(2828);
    outputs(12161) <= not(layer0_outputs(4488));
    outputs(12162) <= not(layer0_outputs(74));
    outputs(12163) <= not(layer0_outputs(9749));
    outputs(12164) <= layer0_outputs(10069);
    outputs(12165) <= (layer0_outputs(1265)) and not (layer0_outputs(5927));
    outputs(12166) <= layer0_outputs(9016);
    outputs(12167) <= layer0_outputs(7241);
    outputs(12168) <= not((layer0_outputs(4264)) xor (layer0_outputs(11643)));
    outputs(12169) <= (layer0_outputs(10427)) and not (layer0_outputs(2655));
    outputs(12170) <= not((layer0_outputs(8915)) or (layer0_outputs(2134)));
    outputs(12171) <= layer0_outputs(11852);
    outputs(12172) <= not(layer0_outputs(9239));
    outputs(12173) <= not(layer0_outputs(5173));
    outputs(12174) <= (layer0_outputs(2419)) xor (layer0_outputs(11541));
    outputs(12175) <= (layer0_outputs(1191)) and (layer0_outputs(3895));
    outputs(12176) <= layer0_outputs(2352);
    outputs(12177) <= not(layer0_outputs(4665));
    outputs(12178) <= (layer0_outputs(1457)) and not (layer0_outputs(8140));
    outputs(12179) <= layer0_outputs(10403);
    outputs(12180) <= (layer0_outputs(12548)) and not (layer0_outputs(10541));
    outputs(12181) <= (layer0_outputs(3618)) xor (layer0_outputs(10436));
    outputs(12182) <= not(layer0_outputs(15));
    outputs(12183) <= (layer0_outputs(12552)) and (layer0_outputs(1705));
    outputs(12184) <= (layer0_outputs(10346)) xor (layer0_outputs(1970));
    outputs(12185) <= layer0_outputs(10631);
    outputs(12186) <= not((layer0_outputs(9847)) xor (layer0_outputs(7284)));
    outputs(12187) <= (layer0_outputs(3264)) and (layer0_outputs(12450));
    outputs(12188) <= layer0_outputs(12086);
    outputs(12189) <= layer0_outputs(1385);
    outputs(12190) <= (layer0_outputs(7097)) xor (layer0_outputs(11867));
    outputs(12191) <= (layer0_outputs(11149)) and (layer0_outputs(9827));
    outputs(12192) <= not((layer0_outputs(9453)) xor (layer0_outputs(11747)));
    outputs(12193) <= (layer0_outputs(3035)) xor (layer0_outputs(3812));
    outputs(12194) <= (layer0_outputs(8912)) xor (layer0_outputs(2067));
    outputs(12195) <= not(layer0_outputs(4292));
    outputs(12196) <= (layer0_outputs(10497)) xor (layer0_outputs(7175));
    outputs(12197) <= not(layer0_outputs(11478));
    outputs(12198) <= not(layer0_outputs(8976));
    outputs(12199) <= not((layer0_outputs(1772)) or (layer0_outputs(1829)));
    outputs(12200) <= (layer0_outputs(7062)) xor (layer0_outputs(8187));
    outputs(12201) <= not((layer0_outputs(7278)) xor (layer0_outputs(3444)));
    outputs(12202) <= not(layer0_outputs(4088));
    outputs(12203) <= layer0_outputs(3545);
    outputs(12204) <= not((layer0_outputs(11504)) xor (layer0_outputs(8929)));
    outputs(12205) <= layer0_outputs(1498);
    outputs(12206) <= not(layer0_outputs(10916));
    outputs(12207) <= not((layer0_outputs(5071)) xor (layer0_outputs(541)));
    outputs(12208) <= (layer0_outputs(12364)) xor (layer0_outputs(11377));
    outputs(12209) <= not(layer0_outputs(7911)) or (layer0_outputs(3934));
    outputs(12210) <= not((layer0_outputs(9546)) or (layer0_outputs(11834)));
    outputs(12211) <= not(layer0_outputs(9567)) or (layer0_outputs(3285));
    outputs(12212) <= (layer0_outputs(271)) and not (layer0_outputs(3532));
    outputs(12213) <= (layer0_outputs(1902)) xor (layer0_outputs(11970));
    outputs(12214) <= not(layer0_outputs(3211));
    outputs(12215) <= layer0_outputs(4152);
    outputs(12216) <= layer0_outputs(5470);
    outputs(12217) <= layer0_outputs(11361);
    outputs(12218) <= (layer0_outputs(12160)) and (layer0_outputs(5569));
    outputs(12219) <= layer0_outputs(3787);
    outputs(12220) <= layer0_outputs(12507);
    outputs(12221) <= not(layer0_outputs(5633));
    outputs(12222) <= (layer0_outputs(1218)) and (layer0_outputs(2754));
    outputs(12223) <= not((layer0_outputs(3705)) or (layer0_outputs(12477)));
    outputs(12224) <= layer0_outputs(12055);
    outputs(12225) <= (layer0_outputs(9519)) xor (layer0_outputs(1489));
    outputs(12226) <= layer0_outputs(5870);
    outputs(12227) <= layer0_outputs(4734);
    outputs(12228) <= not(layer0_outputs(3540));
    outputs(12229) <= (layer0_outputs(10107)) and not (layer0_outputs(7200));
    outputs(12230) <= layer0_outputs(8538);
    outputs(12231) <= (layer0_outputs(9766)) and not (layer0_outputs(4766));
    outputs(12232) <= not((layer0_outputs(8251)) or (layer0_outputs(1966)));
    outputs(12233) <= layer0_outputs(7923);
    outputs(12234) <= not(layer0_outputs(10010));
    outputs(12235) <= layer0_outputs(2083);
    outputs(12236) <= (layer0_outputs(5779)) and (layer0_outputs(10824));
    outputs(12237) <= not(layer0_outputs(4545));
    outputs(12238) <= layer0_outputs(4487);
    outputs(12239) <= (layer0_outputs(3395)) xor (layer0_outputs(12397));
    outputs(12240) <= (layer0_outputs(11327)) xor (layer0_outputs(97));
    outputs(12241) <= (layer0_outputs(12769)) xor (layer0_outputs(4355));
    outputs(12242) <= '0';
    outputs(12243) <= not(layer0_outputs(7080));
    outputs(12244) <= not(layer0_outputs(11456));
    outputs(12245) <= not(layer0_outputs(4696));
    outputs(12246) <= layer0_outputs(10849);
    outputs(12247) <= (layer0_outputs(10720)) xor (layer0_outputs(11903));
    outputs(12248) <= (layer0_outputs(1805)) xor (layer0_outputs(6661));
    outputs(12249) <= not((layer0_outputs(9733)) xor (layer0_outputs(11473)));
    outputs(12250) <= (layer0_outputs(7378)) xor (layer0_outputs(11440));
    outputs(12251) <= not(layer0_outputs(12407)) or (layer0_outputs(11858));
    outputs(12252) <= not((layer0_outputs(7433)) xor (layer0_outputs(6828)));
    outputs(12253) <= not(layer0_outputs(9464));
    outputs(12254) <= not((layer0_outputs(10541)) xor (layer0_outputs(4906)));
    outputs(12255) <= (layer0_outputs(9998)) and not (layer0_outputs(6170));
    outputs(12256) <= not(layer0_outputs(2169));
    outputs(12257) <= not(layer0_outputs(1670));
    outputs(12258) <= not((layer0_outputs(841)) or (layer0_outputs(7192)));
    outputs(12259) <= layer0_outputs(12453);
    outputs(12260) <= not(layer0_outputs(2406));
    outputs(12261) <= layer0_outputs(9996);
    outputs(12262) <= not(layer0_outputs(11507));
    outputs(12263) <= layer0_outputs(3007);
    outputs(12264) <= layer0_outputs(7769);
    outputs(12265) <= not((layer0_outputs(12789)) xor (layer0_outputs(8720)));
    outputs(12266) <= not(layer0_outputs(3795));
    outputs(12267) <= (layer0_outputs(11457)) or (layer0_outputs(8341));
    outputs(12268) <= (layer0_outputs(12371)) and (layer0_outputs(9719));
    outputs(12269) <= not(layer0_outputs(2349));
    outputs(12270) <= not(layer0_outputs(12615));
    outputs(12271) <= not(layer0_outputs(12280));
    outputs(12272) <= not(layer0_outputs(2572));
    outputs(12273) <= not(layer0_outputs(7125));
    outputs(12274) <= not((layer0_outputs(11235)) xor (layer0_outputs(521)));
    outputs(12275) <= (layer0_outputs(5623)) and not (layer0_outputs(4433));
    outputs(12276) <= not((layer0_outputs(5978)) or (layer0_outputs(12381)));
    outputs(12277) <= not(layer0_outputs(7763));
    outputs(12278) <= layer0_outputs(1527);
    outputs(12279) <= (layer0_outputs(9938)) and (layer0_outputs(12356));
    outputs(12280) <= (layer0_outputs(9315)) or (layer0_outputs(5919));
    outputs(12281) <= layer0_outputs(7594);
    outputs(12282) <= (layer0_outputs(9611)) xor (layer0_outputs(10567));
    outputs(12283) <= (layer0_outputs(7781)) and not (layer0_outputs(2186));
    outputs(12284) <= (layer0_outputs(8091)) and not (layer0_outputs(2858));
    outputs(12285) <= not((layer0_outputs(3726)) or (layer0_outputs(5372)));
    outputs(12286) <= layer0_outputs(7415);
    outputs(12287) <= (layer0_outputs(544)) xor (layer0_outputs(2887));
    outputs(12288) <= not(layer0_outputs(6906));
    outputs(12289) <= not(layer0_outputs(5055));
    outputs(12290) <= not((layer0_outputs(10316)) xor (layer0_outputs(1222)));
    outputs(12291) <= not((layer0_outputs(10250)) xor (layer0_outputs(617)));
    outputs(12292) <= layer0_outputs(5515);
    outputs(12293) <= not((layer0_outputs(6712)) and (layer0_outputs(1284)));
    outputs(12294) <= not(layer0_outputs(8536));
    outputs(12295) <= not(layer0_outputs(831));
    outputs(12296) <= not((layer0_outputs(425)) or (layer0_outputs(4156)));
    outputs(12297) <= not(layer0_outputs(9499));
    outputs(12298) <= not(layer0_outputs(5141)) or (layer0_outputs(3339));
    outputs(12299) <= layer0_outputs(5380);
    outputs(12300) <= (layer0_outputs(2787)) and not (layer0_outputs(9825));
    outputs(12301) <= not(layer0_outputs(3721)) or (layer0_outputs(7231));
    outputs(12302) <= (layer0_outputs(3492)) and (layer0_outputs(5810));
    outputs(12303) <= not(layer0_outputs(10831));
    outputs(12304) <= not((layer0_outputs(10857)) or (layer0_outputs(12606)));
    outputs(12305) <= not((layer0_outputs(4789)) xor (layer0_outputs(1153)));
    outputs(12306) <= (layer0_outputs(4939)) and (layer0_outputs(1674));
    outputs(12307) <= layer0_outputs(12225);
    outputs(12308) <= (layer0_outputs(1190)) and (layer0_outputs(5159));
    outputs(12309) <= not(layer0_outputs(8791));
    outputs(12310) <= not(layer0_outputs(8584)) or (layer0_outputs(7408));
    outputs(12311) <= not(layer0_outputs(9518));
    outputs(12312) <= (layer0_outputs(9918)) or (layer0_outputs(10283));
    outputs(12313) <= not(layer0_outputs(99));
    outputs(12314) <= (layer0_outputs(11787)) and not (layer0_outputs(10580));
    outputs(12315) <= layer0_outputs(9599);
    outputs(12316) <= not(layer0_outputs(8655));
    outputs(12317) <= not(layer0_outputs(10684));
    outputs(12318) <= layer0_outputs(4361);
    outputs(12319) <= not((layer0_outputs(5228)) and (layer0_outputs(3631)));
    outputs(12320) <= (layer0_outputs(10643)) or (layer0_outputs(1942));
    outputs(12321) <= (layer0_outputs(9421)) and (layer0_outputs(2963));
    outputs(12322) <= not(layer0_outputs(9680));
    outputs(12323) <= layer0_outputs(2367);
    outputs(12324) <= (layer0_outputs(10376)) xor (layer0_outputs(8624));
    outputs(12325) <= layer0_outputs(12763);
    outputs(12326) <= not(layer0_outputs(9153));
    outputs(12327) <= layer0_outputs(476);
    outputs(12328) <= (layer0_outputs(9029)) and not (layer0_outputs(3014));
    outputs(12329) <= not(layer0_outputs(11264));
    outputs(12330) <= not(layer0_outputs(8397));
    outputs(12331) <= layer0_outputs(8698);
    outputs(12332) <= layer0_outputs(326);
    outputs(12333) <= not((layer0_outputs(2226)) xor (layer0_outputs(8126)));
    outputs(12334) <= layer0_outputs(3834);
    outputs(12335) <= (layer0_outputs(5994)) and (layer0_outputs(6005));
    outputs(12336) <= not(layer0_outputs(453));
    outputs(12337) <= (layer0_outputs(10245)) xor (layer0_outputs(5824));
    outputs(12338) <= not(layer0_outputs(861));
    outputs(12339) <= (layer0_outputs(1048)) xor (layer0_outputs(7915));
    outputs(12340) <= layer0_outputs(4120);
    outputs(12341) <= (layer0_outputs(571)) xor (layer0_outputs(8076));
    outputs(12342) <= layer0_outputs(765);
    outputs(12343) <= not((layer0_outputs(1313)) or (layer0_outputs(11356)));
    outputs(12344) <= layer0_outputs(9197);
    outputs(12345) <= not(layer0_outputs(12705));
    outputs(12346) <= (layer0_outputs(12210)) and not (layer0_outputs(11267));
    outputs(12347) <= (layer0_outputs(4377)) and not (layer0_outputs(644));
    outputs(12348) <= layer0_outputs(3143);
    outputs(12349) <= not((layer0_outputs(5965)) or (layer0_outputs(5420)));
    outputs(12350) <= not(layer0_outputs(4164));
    outputs(12351) <= layer0_outputs(11085);
    outputs(12352) <= not(layer0_outputs(9020));
    outputs(12353) <= not(layer0_outputs(5618));
    outputs(12354) <= layer0_outputs(11015);
    outputs(12355) <= (layer0_outputs(12088)) and (layer0_outputs(8894));
    outputs(12356) <= layer0_outputs(1003);
    outputs(12357) <= not((layer0_outputs(5368)) xor (layer0_outputs(10670)));
    outputs(12358) <= (layer0_outputs(8781)) and (layer0_outputs(394));
    outputs(12359) <= not(layer0_outputs(6339)) or (layer0_outputs(5263));
    outputs(12360) <= not((layer0_outputs(9449)) xor (layer0_outputs(12108)));
    outputs(12361) <= layer0_outputs(6786);
    outputs(12362) <= '0';
    outputs(12363) <= not(layer0_outputs(3510));
    outputs(12364) <= (layer0_outputs(1630)) and not (layer0_outputs(7200));
    outputs(12365) <= not((layer0_outputs(5827)) and (layer0_outputs(3440)));
    outputs(12366) <= layer0_outputs(8841);
    outputs(12367) <= not((layer0_outputs(621)) xor (layer0_outputs(8658)));
    outputs(12368) <= not(layer0_outputs(8122));
    outputs(12369) <= not(layer0_outputs(5944));
    outputs(12370) <= not(layer0_outputs(1959));
    outputs(12371) <= layer0_outputs(1584);
    outputs(12372) <= layer0_outputs(3072);
    outputs(12373) <= layer0_outputs(945);
    outputs(12374) <= not((layer0_outputs(9777)) xor (layer0_outputs(903)));
    outputs(12375) <= layer0_outputs(11584);
    outputs(12376) <= not(layer0_outputs(6256));
    outputs(12377) <= not(layer0_outputs(10123));
    outputs(12378) <= not(layer0_outputs(12458));
    outputs(12379) <= layer0_outputs(6726);
    outputs(12380) <= layer0_outputs(534);
    outputs(12381) <= layer0_outputs(4871);
    outputs(12382) <= not((layer0_outputs(2066)) xor (layer0_outputs(4637)));
    outputs(12383) <= not((layer0_outputs(4191)) or (layer0_outputs(12772)));
    outputs(12384) <= not(layer0_outputs(503));
    outputs(12385) <= not(layer0_outputs(592)) or (layer0_outputs(2074));
    outputs(12386) <= (layer0_outputs(2826)) and (layer0_outputs(11829));
    outputs(12387) <= (layer0_outputs(1579)) xor (layer0_outputs(7085));
    outputs(12388) <= not((layer0_outputs(1422)) xor (layer0_outputs(4853)));
    outputs(12389) <= not(layer0_outputs(5346));
    outputs(12390) <= not((layer0_outputs(704)) or (layer0_outputs(5922)));
    outputs(12391) <= not(layer0_outputs(8917));
    outputs(12392) <= (layer0_outputs(11665)) and (layer0_outputs(779));
    outputs(12393) <= not(layer0_outputs(11963));
    outputs(12394) <= not((layer0_outputs(4825)) xor (layer0_outputs(7221)));
    outputs(12395) <= '0';
    outputs(12396) <= not((layer0_outputs(11028)) or (layer0_outputs(8105)));
    outputs(12397) <= not(layer0_outputs(8676)) or (layer0_outputs(11136));
    outputs(12398) <= layer0_outputs(10071);
    outputs(12399) <= (layer0_outputs(10950)) xor (layer0_outputs(10030));
    outputs(12400) <= (layer0_outputs(11912)) xor (layer0_outputs(4144));
    outputs(12401) <= not((layer0_outputs(9342)) xor (layer0_outputs(5081)));
    outputs(12402) <= layer0_outputs(9540);
    outputs(12403) <= layer0_outputs(4234);
    outputs(12404) <= (layer0_outputs(4679)) and not (layer0_outputs(837));
    outputs(12405) <= not((layer0_outputs(5007)) or (layer0_outputs(1960)));
    outputs(12406) <= layer0_outputs(1454);
    outputs(12407) <= not(layer0_outputs(7996));
    outputs(12408) <= layer0_outputs(4187);
    outputs(12409) <= not(layer0_outputs(12173));
    outputs(12410) <= (layer0_outputs(2263)) xor (layer0_outputs(6132));
    outputs(12411) <= not(layer0_outputs(11610));
    outputs(12412) <= (layer0_outputs(2003)) and (layer0_outputs(11922));
    outputs(12413) <= (layer0_outputs(11496)) and not (layer0_outputs(7634));
    outputs(12414) <= (layer0_outputs(10844)) and not (layer0_outputs(11315));
    outputs(12415) <= not(layer0_outputs(9917));
    outputs(12416) <= (layer0_outputs(9298)) and not (layer0_outputs(3391));
    outputs(12417) <= not(layer0_outputs(4425));
    outputs(12418) <= not((layer0_outputs(84)) or (layer0_outputs(1996)));
    outputs(12419) <= layer0_outputs(6278);
    outputs(12420) <= not((layer0_outputs(10892)) xor (layer0_outputs(7585)));
    outputs(12421) <= not(layer0_outputs(73));
    outputs(12422) <= layer0_outputs(4417);
    outputs(12423) <= not(layer0_outputs(5086));
    outputs(12424) <= (layer0_outputs(11229)) xor (layer0_outputs(1651));
    outputs(12425) <= not((layer0_outputs(8156)) xor (layer0_outputs(3441)));
    outputs(12426) <= not((layer0_outputs(10995)) and (layer0_outputs(8829)));
    outputs(12427) <= layer0_outputs(238);
    outputs(12428) <= not(layer0_outputs(5616)) or (layer0_outputs(4522));
    outputs(12429) <= not((layer0_outputs(7688)) or (layer0_outputs(1626)));
    outputs(12430) <= not((layer0_outputs(3327)) xor (layer0_outputs(6902)));
    outputs(12431) <= not((layer0_outputs(8524)) xor (layer0_outputs(9397)));
    outputs(12432) <= not(layer0_outputs(12549));
    outputs(12433) <= layer0_outputs(8574);
    outputs(12434) <= layer0_outputs(8601);
    outputs(12435) <= layer0_outputs(5439);
    outputs(12436) <= not(layer0_outputs(2696));
    outputs(12437) <= layer0_outputs(7521);
    outputs(12438) <= (layer0_outputs(2208)) xor (layer0_outputs(3754));
    outputs(12439) <= (layer0_outputs(6451)) and (layer0_outputs(5244));
    outputs(12440) <= not(layer0_outputs(6079));
    outputs(12441) <= layer0_outputs(1950);
    outputs(12442) <= (layer0_outputs(6824)) and (layer0_outputs(1208));
    outputs(12443) <= (layer0_outputs(7076)) and not (layer0_outputs(7517));
    outputs(12444) <= (layer0_outputs(1275)) xor (layer0_outputs(3905));
    outputs(12445) <= not((layer0_outputs(5796)) or (layer0_outputs(5174)));
    outputs(12446) <= layer0_outputs(546);
    outputs(12447) <= (layer0_outputs(6217)) or (layer0_outputs(4626));
    outputs(12448) <= layer0_outputs(1332);
    outputs(12449) <= not(layer0_outputs(4892)) or (layer0_outputs(11130));
    outputs(12450) <= (layer0_outputs(8110)) and not (layer0_outputs(10026));
    outputs(12451) <= not(layer0_outputs(10560)) or (layer0_outputs(3965));
    outputs(12452) <= (layer0_outputs(12165)) and (layer0_outputs(9479));
    outputs(12453) <= layer0_outputs(88);
    outputs(12454) <= layer0_outputs(3366);
    outputs(12455) <= layer0_outputs(9388);
    outputs(12456) <= (layer0_outputs(11269)) xor (layer0_outputs(2809));
    outputs(12457) <= not((layer0_outputs(5411)) xor (layer0_outputs(6106)));
    outputs(12458) <= (layer0_outputs(1367)) and not (layer0_outputs(11935));
    outputs(12459) <= not((layer0_outputs(10811)) xor (layer0_outputs(4032)));
    outputs(12460) <= not(layer0_outputs(5156)) or (layer0_outputs(3628));
    outputs(12461) <= (layer0_outputs(6717)) xor (layer0_outputs(11240));
    outputs(12462) <= not((layer0_outputs(11314)) xor (layer0_outputs(7474)));
    outputs(12463) <= not(layer0_outputs(8002));
    outputs(12464) <= (layer0_outputs(7894)) and not (layer0_outputs(3464));
    outputs(12465) <= layer0_outputs(10851);
    outputs(12466) <= not(layer0_outputs(9102));
    outputs(12467) <= (layer0_outputs(11189)) and not (layer0_outputs(8751));
    outputs(12468) <= not((layer0_outputs(6741)) xor (layer0_outputs(11537)));
    outputs(12469) <= (layer0_outputs(2674)) xor (layer0_outputs(7573));
    outputs(12470) <= layer0_outputs(3591);
    outputs(12471) <= layer0_outputs(1288);
    outputs(12472) <= (layer0_outputs(8370)) and not (layer0_outputs(5950));
    outputs(12473) <= not(layer0_outputs(361));
    outputs(12474) <= not(layer0_outputs(871));
    outputs(12475) <= layer0_outputs(10990);
    outputs(12476) <= (layer0_outputs(2040)) and not (layer0_outputs(5914));
    outputs(12477) <= not(layer0_outputs(4501));
    outputs(12478) <= not((layer0_outputs(729)) xor (layer0_outputs(4747)));
    outputs(12479) <= (layer0_outputs(7216)) and not (layer0_outputs(8733));
    outputs(12480) <= not(layer0_outputs(8078));
    outputs(12481) <= not(layer0_outputs(4878));
    outputs(12482) <= not((layer0_outputs(6925)) and (layer0_outputs(2127)));
    outputs(12483) <= layer0_outputs(6870);
    outputs(12484) <= not(layer0_outputs(2117));
    outputs(12485) <= layer0_outputs(10092);
    outputs(12486) <= (layer0_outputs(8928)) and not (layer0_outputs(6409));
    outputs(12487) <= not(layer0_outputs(1413));
    outputs(12488) <= layer0_outputs(9344);
    outputs(12489) <= (layer0_outputs(5693)) and not (layer0_outputs(12438));
    outputs(12490) <= layer0_outputs(9303);
    outputs(12491) <= not(layer0_outputs(5151));
    outputs(12492) <= not((layer0_outputs(9433)) xor (layer0_outputs(3654)));
    outputs(12493) <= layer0_outputs(8962);
    outputs(12494) <= not((layer0_outputs(6731)) xor (layer0_outputs(2301)));
    outputs(12495) <= not(layer0_outputs(5128));
    outputs(12496) <= layer0_outputs(2212);
    outputs(12497) <= (layer0_outputs(9154)) and not (layer0_outputs(751));
    outputs(12498) <= not(layer0_outputs(624)) or (layer0_outputs(7986));
    outputs(12499) <= (layer0_outputs(6479)) xor (layer0_outputs(9997));
    outputs(12500) <= not(layer0_outputs(6006));
    outputs(12501) <= (layer0_outputs(10302)) xor (layer0_outputs(11279));
    outputs(12502) <= (layer0_outputs(12602)) and (layer0_outputs(417));
    outputs(12503) <= not((layer0_outputs(4241)) and (layer0_outputs(10281)));
    outputs(12504) <= (layer0_outputs(1062)) and not (layer0_outputs(8021));
    outputs(12505) <= (layer0_outputs(5571)) xor (layer0_outputs(10720));
    outputs(12506) <= not((layer0_outputs(5413)) or (layer0_outputs(8803)));
    outputs(12507) <= layer0_outputs(2968);
    outputs(12508) <= (layer0_outputs(7771)) xor (layer0_outputs(4756));
    outputs(12509) <= not(layer0_outputs(9346));
    outputs(12510) <= layer0_outputs(8781);
    outputs(12511) <= not(layer0_outputs(178));
    outputs(12512) <= (layer0_outputs(3475)) xor (layer0_outputs(412));
    outputs(12513) <= not(layer0_outputs(1223)) or (layer0_outputs(10832));
    outputs(12514) <= (layer0_outputs(894)) and not (layer0_outputs(5130));
    outputs(12515) <= not((layer0_outputs(927)) or (layer0_outputs(3462)));
    outputs(12516) <= (layer0_outputs(12491)) and not (layer0_outputs(612));
    outputs(12517) <= not(layer0_outputs(9468));
    outputs(12518) <= layer0_outputs(11926);
    outputs(12519) <= (layer0_outputs(2305)) xor (layer0_outputs(9964));
    outputs(12520) <= not((layer0_outputs(5356)) xor (layer0_outputs(3491)));
    outputs(12521) <= not(layer0_outputs(10569));
    outputs(12522) <= layer0_outputs(11447);
    outputs(12523) <= (layer0_outputs(6788)) and not (layer0_outputs(2586));
    outputs(12524) <= not((layer0_outputs(12422)) xor (layer0_outputs(11186)));
    outputs(12525) <= not(layer0_outputs(8665));
    outputs(12526) <= not(layer0_outputs(182));
    outputs(12527) <= layer0_outputs(12725);
    outputs(12528) <= layer0_outputs(2609);
    outputs(12529) <= not((layer0_outputs(6919)) or (layer0_outputs(8004)));
    outputs(12530) <= not(layer0_outputs(1999));
    outputs(12531) <= not((layer0_outputs(12056)) xor (layer0_outputs(498)));
    outputs(12532) <= (layer0_outputs(5199)) and (layer0_outputs(5992));
    outputs(12533) <= (layer0_outputs(1021)) xor (layer0_outputs(2562));
    outputs(12534) <= (layer0_outputs(1985)) xor (layer0_outputs(3273));
    outputs(12535) <= (layer0_outputs(12269)) xor (layer0_outputs(5319));
    outputs(12536) <= not((layer0_outputs(7952)) or (layer0_outputs(11695)));
    outputs(12537) <= not(layer0_outputs(11397));
    outputs(12538) <= not((layer0_outputs(3503)) and (layer0_outputs(4806)));
    outputs(12539) <= not((layer0_outputs(6415)) and (layer0_outputs(9596)));
    outputs(12540) <= (layer0_outputs(2829)) and not (layer0_outputs(1819));
    outputs(12541) <= layer0_outputs(10300);
    outputs(12542) <= not(layer0_outputs(11874));
    outputs(12543) <= (layer0_outputs(5395)) xor (layer0_outputs(7369));
    outputs(12544) <= not(layer0_outputs(315));
    outputs(12545) <= (layer0_outputs(6916)) xor (layer0_outputs(1764));
    outputs(12546) <= (layer0_outputs(11775)) and (layer0_outputs(9272));
    outputs(12547) <= not((layer0_outputs(8008)) xor (layer0_outputs(688)));
    outputs(12548) <= layer0_outputs(8129);
    outputs(12549) <= layer0_outputs(6553);
    outputs(12550) <= layer0_outputs(1940);
    outputs(12551) <= not(layer0_outputs(6000)) or (layer0_outputs(430));
    outputs(12552) <= not(layer0_outputs(6200));
    outputs(12553) <= (layer0_outputs(9029)) and (layer0_outputs(12186));
    outputs(12554) <= not(layer0_outputs(5466));
    outputs(12555) <= layer0_outputs(8402);
    outputs(12556) <= (layer0_outputs(1512)) and not (layer0_outputs(3364));
    outputs(12557) <= not(layer0_outputs(5675));
    outputs(12558) <= not(layer0_outputs(4180));
    outputs(12559) <= (layer0_outputs(6021)) or (layer0_outputs(9275));
    outputs(12560) <= layer0_outputs(6846);
    outputs(12561) <= not((layer0_outputs(12226)) xor (layer0_outputs(11826)));
    outputs(12562) <= (layer0_outputs(9966)) or (layer0_outputs(12488));
    outputs(12563) <= not(layer0_outputs(6488));
    outputs(12564) <= not((layer0_outputs(2524)) or (layer0_outputs(11699)));
    outputs(12565) <= (layer0_outputs(116)) or (layer0_outputs(2387));
    outputs(12566) <= not(layer0_outputs(7497));
    outputs(12567) <= layer0_outputs(209);
    outputs(12568) <= not((layer0_outputs(8595)) or (layer0_outputs(3990)));
    outputs(12569) <= (layer0_outputs(5145)) and not (layer0_outputs(3136));
    outputs(12570) <= not((layer0_outputs(3916)) xor (layer0_outputs(2554)));
    outputs(12571) <= (layer0_outputs(6564)) and (layer0_outputs(10548));
    outputs(12572) <= layer0_outputs(6794);
    outputs(12573) <= layer0_outputs(10315);
    outputs(12574) <= not(layer0_outputs(11723));
    outputs(12575) <= not(layer0_outputs(8966));
    outputs(12576) <= not(layer0_outputs(8956));
    outputs(12577) <= layer0_outputs(5795);
    outputs(12578) <= not((layer0_outputs(1209)) xor (layer0_outputs(202)));
    outputs(12579) <= not((layer0_outputs(5137)) xor (layer0_outputs(10615)));
    outputs(12580) <= (layer0_outputs(5725)) and (layer0_outputs(9215));
    outputs(12581) <= layer0_outputs(10384);
    outputs(12582) <= not((layer0_outputs(12728)) xor (layer0_outputs(2322)));
    outputs(12583) <= not(layer0_outputs(8904));
    outputs(12584) <= (layer0_outputs(5862)) and not (layer0_outputs(2840));
    outputs(12585) <= (layer0_outputs(10614)) xor (layer0_outputs(4177));
    outputs(12586) <= not((layer0_outputs(9864)) xor (layer0_outputs(6807)));
    outputs(12587) <= not(layer0_outputs(6401));
    outputs(12588) <= not((layer0_outputs(8608)) or (layer0_outputs(11129)));
    outputs(12589) <= layer0_outputs(8452);
    outputs(12590) <= not(layer0_outputs(9346));
    outputs(12591) <= layer0_outputs(4277);
    outputs(12592) <= layer0_outputs(11519);
    outputs(12593) <= layer0_outputs(2087);
    outputs(12594) <= not((layer0_outputs(6593)) xor (layer0_outputs(11319)));
    outputs(12595) <= layer0_outputs(3990);
    outputs(12596) <= layer0_outputs(9879);
    outputs(12597) <= not(layer0_outputs(1553));
    outputs(12598) <= not(layer0_outputs(8121)) or (layer0_outputs(1348));
    outputs(12599) <= not(layer0_outputs(6932));
    outputs(12600) <= not((layer0_outputs(527)) xor (layer0_outputs(7581)));
    outputs(12601) <= not(layer0_outputs(7491));
    outputs(12602) <= not((layer0_outputs(1022)) xor (layer0_outputs(3806)));
    outputs(12603) <= not(layer0_outputs(6211)) or (layer0_outputs(2904));
    outputs(12604) <= not((layer0_outputs(8200)) xor (layer0_outputs(10204)));
    outputs(12605) <= layer0_outputs(2632);
    outputs(12606) <= (layer0_outputs(148)) and (layer0_outputs(12349));
    outputs(12607) <= not(layer0_outputs(8921));
    outputs(12608) <= layer0_outputs(954);
    outputs(12609) <= (layer0_outputs(7370)) xor (layer0_outputs(2814));
    outputs(12610) <= layer0_outputs(5858);
    outputs(12611) <= not((layer0_outputs(7600)) xor (layer0_outputs(11883)));
    outputs(12612) <= layer0_outputs(2728);
    outputs(12613) <= layer0_outputs(6715);
    outputs(12614) <= not((layer0_outputs(2465)) and (layer0_outputs(1611)));
    outputs(12615) <= not(layer0_outputs(1993));
    outputs(12616) <= (layer0_outputs(7047)) and not (layer0_outputs(2951));
    outputs(12617) <= not(layer0_outputs(1229));
    outputs(12618) <= not((layer0_outputs(12122)) xor (layer0_outputs(4259)));
    outputs(12619) <= (layer0_outputs(5001)) xor (layer0_outputs(3648));
    outputs(12620) <= layer0_outputs(5160);
    outputs(12621) <= layer0_outputs(5105);
    outputs(12622) <= layer0_outputs(2957);
    outputs(12623) <= (layer0_outputs(781)) xor (layer0_outputs(12547));
    outputs(12624) <= not((layer0_outputs(12030)) xor (layer0_outputs(4340)));
    outputs(12625) <= (layer0_outputs(5900)) or (layer0_outputs(4727));
    outputs(12626) <= layer0_outputs(9659);
    outputs(12627) <= (layer0_outputs(5423)) and (layer0_outputs(5666));
    outputs(12628) <= (layer0_outputs(2543)) and (layer0_outputs(2823));
    outputs(12629) <= (layer0_outputs(3477)) xor (layer0_outputs(10725));
    outputs(12630) <= (layer0_outputs(5645)) and not (layer0_outputs(4));
    outputs(12631) <= (layer0_outputs(8025)) and not (layer0_outputs(10768));
    outputs(12632) <= not(layer0_outputs(9268));
    outputs(12633) <= layer0_outputs(2472);
    outputs(12634) <= (layer0_outputs(8545)) and (layer0_outputs(8129));
    outputs(12635) <= (layer0_outputs(2245)) and not (layer0_outputs(4694));
    outputs(12636) <= (layer0_outputs(11117)) and not (layer0_outputs(6664));
    outputs(12637) <= layer0_outputs(5459);
    outputs(12638) <= not(layer0_outputs(5138));
    outputs(12639) <= not(layer0_outputs(7465));
    outputs(12640) <= not(layer0_outputs(8585));
    outputs(12641) <= not(layer0_outputs(7116));
    outputs(12642) <= (layer0_outputs(1221)) xor (layer0_outputs(7035));
    outputs(12643) <= not((layer0_outputs(11666)) xor (layer0_outputs(21)));
    outputs(12644) <= (layer0_outputs(10219)) and not (layer0_outputs(269));
    outputs(12645) <= not(layer0_outputs(6832));
    outputs(12646) <= (layer0_outputs(11603)) and (layer0_outputs(6124));
    outputs(12647) <= not((layer0_outputs(584)) or (layer0_outputs(2123)));
    outputs(12648) <= not((layer0_outputs(12301)) or (layer0_outputs(4529)));
    outputs(12649) <= (layer0_outputs(10559)) and not (layer0_outputs(10598));
    outputs(12650) <= layer0_outputs(10288);
    outputs(12651) <= layer0_outputs(6395);
    outputs(12652) <= (layer0_outputs(1915)) and not (layer0_outputs(53));
    outputs(12653) <= not(layer0_outputs(3230));
    outputs(12654) <= (layer0_outputs(7631)) and not (layer0_outputs(720));
    outputs(12655) <= '0';
    outputs(12656) <= not((layer0_outputs(11688)) xor (layer0_outputs(1280)));
    outputs(12657) <= (layer0_outputs(4372)) xor (layer0_outputs(1367));
    outputs(12658) <= not(layer0_outputs(1910));
    outputs(12659) <= not((layer0_outputs(4763)) or (layer0_outputs(12085)));
    outputs(12660) <= not(layer0_outputs(3169));
    outputs(12661) <= layer0_outputs(6316);
    outputs(12662) <= not((layer0_outputs(1304)) or (layer0_outputs(473)));
    outputs(12663) <= not((layer0_outputs(11389)) xor (layer0_outputs(7847)));
    outputs(12664) <= not((layer0_outputs(1954)) xor (layer0_outputs(2981)));
    outputs(12665) <= not((layer0_outputs(6206)) or (layer0_outputs(2039)));
    outputs(12666) <= layer0_outputs(719);
    outputs(12667) <= not(layer0_outputs(10344));
    outputs(12668) <= layer0_outputs(4274);
    outputs(12669) <= (layer0_outputs(300)) xor (layer0_outputs(373));
    outputs(12670) <= layer0_outputs(892);
    outputs(12671) <= (layer0_outputs(1298)) xor (layer0_outputs(8436));
    outputs(12672) <= (layer0_outputs(10184)) xor (layer0_outputs(6304));
    outputs(12673) <= not(layer0_outputs(11693));
    outputs(12674) <= (layer0_outputs(918)) and not (layer0_outputs(8344));
    outputs(12675) <= not(layer0_outputs(1023));
    outputs(12676) <= not((layer0_outputs(2346)) xor (layer0_outputs(6980)));
    outputs(12677) <= not(layer0_outputs(2603)) or (layer0_outputs(8494));
    outputs(12678) <= not(layer0_outputs(1899));
    outputs(12679) <= layer0_outputs(12275);
    outputs(12680) <= not(layer0_outputs(10290)) or (layer0_outputs(7732));
    outputs(12681) <= (layer0_outputs(840)) xor (layer0_outputs(297));
    outputs(12682) <= not((layer0_outputs(4490)) xor (layer0_outputs(2330)));
    outputs(12683) <= not(layer0_outputs(8127));
    outputs(12684) <= (layer0_outputs(12123)) and not (layer0_outputs(5147));
    outputs(12685) <= not(layer0_outputs(820));
    outputs(12686) <= layer0_outputs(8143);
    outputs(12687) <= layer0_outputs(11678);
    outputs(12688) <= not(layer0_outputs(12762));
    outputs(12689) <= not(layer0_outputs(10878)) or (layer0_outputs(1352));
    outputs(12690) <= layer0_outputs(6354);
    outputs(12691) <= not(layer0_outputs(11510)) or (layer0_outputs(4828));
    outputs(12692) <= not(layer0_outputs(9105)) or (layer0_outputs(9892));
    outputs(12693) <= not((layer0_outputs(10380)) xor (layer0_outputs(1588)));
    outputs(12694) <= (layer0_outputs(2506)) xor (layer0_outputs(9460));
    outputs(12695) <= (layer0_outputs(5019)) and not (layer0_outputs(12256));
    outputs(12696) <= (layer0_outputs(9215)) xor (layer0_outputs(11499));
    outputs(12697) <= (layer0_outputs(12665)) xor (layer0_outputs(3582));
    outputs(12698) <= not(layer0_outputs(3085));
    outputs(12699) <= (layer0_outputs(9815)) or (layer0_outputs(5926));
    outputs(12700) <= layer0_outputs(9671);
    outputs(12701) <= (layer0_outputs(11159)) or (layer0_outputs(4620));
    outputs(12702) <= not(layer0_outputs(10538));
    outputs(12703) <= (layer0_outputs(12082)) and not (layer0_outputs(6089));
    outputs(12704) <= layer0_outputs(12445);
    outputs(12705) <= (layer0_outputs(10808)) and not (layer0_outputs(717));
    outputs(12706) <= not(layer0_outputs(4709));
    outputs(12707) <= not(layer0_outputs(10552));
    outputs(12708) <= not(layer0_outputs(5154));
    outputs(12709) <= (layer0_outputs(1856)) xor (layer0_outputs(4059));
    outputs(12710) <= (layer0_outputs(1369)) and not (layer0_outputs(10622));
    outputs(12711) <= (layer0_outputs(4441)) and (layer0_outputs(3504));
    outputs(12712) <= not((layer0_outputs(2688)) and (layer0_outputs(2283)));
    outputs(12713) <= not((layer0_outputs(6863)) or (layer0_outputs(9519)));
    outputs(12714) <= (layer0_outputs(8795)) or (layer0_outputs(6173));
    outputs(12715) <= not((layer0_outputs(3028)) or (layer0_outputs(5266)));
    outputs(12716) <= not(layer0_outputs(5107));
    outputs(12717) <= not(layer0_outputs(9895));
    outputs(12718) <= layer0_outputs(4054);
    outputs(12719) <= (layer0_outputs(4719)) and not (layer0_outputs(12156));
    outputs(12720) <= layer0_outputs(10179);
    outputs(12721) <= not(layer0_outputs(157));
    outputs(12722) <= (layer0_outputs(11830)) and (layer0_outputs(6140));
    outputs(12723) <= layer0_outputs(10051);
    outputs(12724) <= (layer0_outputs(6761)) xor (layer0_outputs(8845));
    outputs(12725) <= layer0_outputs(4107);
    outputs(12726) <= not((layer0_outputs(6219)) or (layer0_outputs(5300)));
    outputs(12727) <= not(layer0_outputs(6699));
    outputs(12728) <= not((layer0_outputs(11885)) and (layer0_outputs(9723)));
    outputs(12729) <= not(layer0_outputs(12420));
    outputs(12730) <= (layer0_outputs(10667)) and not (layer0_outputs(7016));
    outputs(12731) <= not(layer0_outputs(3588));
    outputs(12732) <= not(layer0_outputs(9615));
    outputs(12733) <= layer0_outputs(417);
    outputs(12734) <= layer0_outputs(7620);
    outputs(12735) <= (layer0_outputs(4839)) and not (layer0_outputs(1464));
    outputs(12736) <= layer0_outputs(893);
    outputs(12737) <= not((layer0_outputs(1965)) and (layer0_outputs(6223)));
    outputs(12738) <= not(layer0_outputs(10089));
    outputs(12739) <= layer0_outputs(9798);
    outputs(12740) <= (layer0_outputs(10388)) and (layer0_outputs(3996));
    outputs(12741) <= (layer0_outputs(3248)) and not (layer0_outputs(674));
    outputs(12742) <= layer0_outputs(601);
    outputs(12743) <= not((layer0_outputs(5328)) xor (layer0_outputs(10873)));
    outputs(12744) <= (layer0_outputs(11586)) xor (layer0_outputs(12583));
    outputs(12745) <= not(layer0_outputs(2225));
    outputs(12746) <= not(layer0_outputs(3289));
    outputs(12747) <= not(layer0_outputs(4410));
    outputs(12748) <= not((layer0_outputs(5337)) and (layer0_outputs(2414)));
    outputs(12749) <= (layer0_outputs(8636)) and not (layer0_outputs(8315));
    outputs(12750) <= (layer0_outputs(9027)) and not (layer0_outputs(12018));
    outputs(12751) <= (layer0_outputs(3307)) and (layer0_outputs(6701));
    outputs(12752) <= not((layer0_outputs(3830)) or (layer0_outputs(12474)));
    outputs(12753) <= (layer0_outputs(5670)) xor (layer0_outputs(3772));
    outputs(12754) <= not((layer0_outputs(5042)) and (layer0_outputs(7522)));
    outputs(12755) <= not(layer0_outputs(10004));
    outputs(12756) <= (layer0_outputs(2686)) xor (layer0_outputs(10562));
    outputs(12757) <= not(layer0_outputs(11023));
    outputs(12758) <= (layer0_outputs(8365)) and not (layer0_outputs(803));
    outputs(12759) <= not((layer0_outputs(6389)) or (layer0_outputs(4685)));
    outputs(12760) <= layer0_outputs(10964);
    outputs(12761) <= not(layer0_outputs(12777));
    outputs(12762) <= not(layer0_outputs(3204));
    outputs(12763) <= not(layer0_outputs(3255));
    outputs(12764) <= (layer0_outputs(1500)) or (layer0_outputs(891));
    outputs(12765) <= (layer0_outputs(4316)) xor (layer0_outputs(1761));
    outputs(12766) <= (layer0_outputs(360)) and (layer0_outputs(7944));
    outputs(12767) <= layer0_outputs(5199);
    outputs(12768) <= (layer0_outputs(8082)) xor (layer0_outputs(5979));
    outputs(12769) <= not(layer0_outputs(11150));
    outputs(12770) <= not((layer0_outputs(11606)) xor (layer0_outputs(204)));
    outputs(12771) <= not(layer0_outputs(1131));
    outputs(12772) <= not((layer0_outputs(6524)) xor (layer0_outputs(3971)));
    outputs(12773) <= layer0_outputs(6309);
    outputs(12774) <= layer0_outputs(4135);
    outputs(12775) <= (layer0_outputs(7863)) and (layer0_outputs(10304));
    outputs(12776) <= not((layer0_outputs(3263)) or (layer0_outputs(77)));
    outputs(12777) <= not(layer0_outputs(99));
    outputs(12778) <= not(layer0_outputs(8555)) or (layer0_outputs(9639));
    outputs(12779) <= not((layer0_outputs(1554)) or (layer0_outputs(12154)));
    outputs(12780) <= not(layer0_outputs(11031));
    outputs(12781) <= layer0_outputs(4426);
    outputs(12782) <= not(layer0_outputs(5059));
    outputs(12783) <= (layer0_outputs(277)) xor (layer0_outputs(975));
    outputs(12784) <= layer0_outputs(7388);
    outputs(12785) <= not(layer0_outputs(1499));
    outputs(12786) <= not(layer0_outputs(53));
    outputs(12787) <= not(layer0_outputs(12339));
    outputs(12788) <= not(layer0_outputs(5633));
    outputs(12789) <= not((layer0_outputs(9561)) xor (layer0_outputs(914)));
    outputs(12790) <= not((layer0_outputs(11706)) xor (layer0_outputs(9258)));
    outputs(12791) <= (layer0_outputs(9737)) and not (layer0_outputs(4263));
    outputs(12792) <= (layer0_outputs(601)) and not (layer0_outputs(7270));
    outputs(12793) <= not((layer0_outputs(6800)) xor (layer0_outputs(752)));
    outputs(12794) <= not(layer0_outputs(12454)) or (layer0_outputs(11147));
    outputs(12795) <= not(layer0_outputs(7451));
    outputs(12796) <= layer0_outputs(7576);
    outputs(12797) <= layer0_outputs(8450);
    outputs(12798) <= not(layer0_outputs(3644));
    outputs(12799) <= not(layer0_outputs(7055));

end Behavioral;
