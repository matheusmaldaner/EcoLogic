library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(7679 downto 0);
    signal layer1_outputs: std_logic_vector(7679 downto 0);
    signal layer2_outputs: std_logic_vector(7679 downto 0);
    signal layer3_outputs: std_logic_vector(7679 downto 0);
    signal layer4_outputs: std_logic_vector(7679 downto 0);
    signal layer5_outputs: std_logic_vector(7679 downto 0);
    signal layer6_outputs: std_logic_vector(7679 downto 0);
    signal layer7_outputs: std_logic_vector(7679 downto 0);
    signal layer8_outputs: std_logic_vector(7679 downto 0);

begin
    layer0_outputs(0) <= '0';
    layer0_outputs(1) <= b;
    layer0_outputs(2) <= not (a xor b);
    layer0_outputs(3) <= not a;
    layer0_outputs(4) <= not b or a;
    layer0_outputs(5) <= not a or b;
    layer0_outputs(6) <= not a;
    layer0_outputs(7) <= '0';
    layer0_outputs(8) <= b;
    layer0_outputs(9) <= '0';
    layer0_outputs(10) <= not b or a;
    layer0_outputs(11) <= a;
    layer0_outputs(12) <= not a;
    layer0_outputs(13) <= not (a and b);
    layer0_outputs(14) <= not a;
    layer0_outputs(15) <= b and not a;
    layer0_outputs(16) <= b;
    layer0_outputs(17) <= not b;
    layer0_outputs(18) <= '0';
    layer0_outputs(19) <= a;
    layer0_outputs(20) <= not a;
    layer0_outputs(21) <= '0';
    layer0_outputs(22) <= not a or b;
    layer0_outputs(23) <= not (a and b);
    layer0_outputs(24) <= b;
    layer0_outputs(25) <= b;
    layer0_outputs(26) <= not (a xor b);
    layer0_outputs(27) <= a;
    layer0_outputs(28) <= b;
    layer0_outputs(29) <= not b;
    layer0_outputs(30) <= a or b;
    layer0_outputs(31) <= not a;
    layer0_outputs(32) <= not b;
    layer0_outputs(33) <= not (a and b);
    layer0_outputs(34) <= a;
    layer0_outputs(35) <= b;
    layer0_outputs(36) <= a;
    layer0_outputs(37) <= a;
    layer0_outputs(38) <= '1';
    layer0_outputs(39) <= not a or b;
    layer0_outputs(40) <= a xor b;
    layer0_outputs(41) <= b;
    layer0_outputs(42) <= not b;
    layer0_outputs(43) <= '1';
    layer0_outputs(44) <= not (a xor b);
    layer0_outputs(45) <= not (a xor b);
    layer0_outputs(46) <= a or b;
    layer0_outputs(47) <= b;
    layer0_outputs(48) <= not a;
    layer0_outputs(49) <= not a;
    layer0_outputs(50) <= not (a and b);
    layer0_outputs(51) <= b;
    layer0_outputs(52) <= not b;
    layer0_outputs(53) <= '0';
    layer0_outputs(54) <= not (a xor b);
    layer0_outputs(55) <= not b or a;
    layer0_outputs(56) <= a and b;
    layer0_outputs(57) <= not a;
    layer0_outputs(58) <= not (a and b);
    layer0_outputs(59) <= not b;
    layer0_outputs(60) <= a;
    layer0_outputs(61) <= a and not b;
    layer0_outputs(62) <= not (a or b);
    layer0_outputs(63) <= a xor b;
    layer0_outputs(64) <= not a or b;
    layer0_outputs(65) <= not b;
    layer0_outputs(66) <= not (a or b);
    layer0_outputs(67) <= not (a xor b);
    layer0_outputs(68) <= not b or a;
    layer0_outputs(69) <= not b or a;
    layer0_outputs(70) <= not b or a;
    layer0_outputs(71) <= '1';
    layer0_outputs(72) <= '0';
    layer0_outputs(73) <= not a or b;
    layer0_outputs(74) <= b;
    layer0_outputs(75) <= a;
    layer0_outputs(76) <= '0';
    layer0_outputs(77) <= not (a or b);
    layer0_outputs(78) <= a and not b;
    layer0_outputs(79) <= a and not b;
    layer0_outputs(80) <= b and not a;
    layer0_outputs(81) <= not b;
    layer0_outputs(82) <= a or b;
    layer0_outputs(83) <= '1';
    layer0_outputs(84) <= '1';
    layer0_outputs(85) <= not (a xor b);
    layer0_outputs(86) <= a;
    layer0_outputs(87) <= not a or b;
    layer0_outputs(88) <= not (a or b);
    layer0_outputs(89) <= '1';
    layer0_outputs(90) <= not (a xor b);
    layer0_outputs(91) <= not b or a;
    layer0_outputs(92) <= a or b;
    layer0_outputs(93) <= a or b;
    layer0_outputs(94) <= a xor b;
    layer0_outputs(95) <= not b;
    layer0_outputs(96) <= b;
    layer0_outputs(97) <= b and not a;
    layer0_outputs(98) <= not a or b;
    layer0_outputs(99) <= not b;
    layer0_outputs(100) <= not b;
    layer0_outputs(101) <= not (a or b);
    layer0_outputs(102) <= '1';
    layer0_outputs(103) <= not (a xor b);
    layer0_outputs(104) <= not a or b;
    layer0_outputs(105) <= not b or a;
    layer0_outputs(106) <= '1';
    layer0_outputs(107) <= not (a or b);
    layer0_outputs(108) <= '0';
    layer0_outputs(109) <= a;
    layer0_outputs(110) <= not (a and b);
    layer0_outputs(111) <= a or b;
    layer0_outputs(112) <= a and not b;
    layer0_outputs(113) <= a;
    layer0_outputs(114) <= not (a and b);
    layer0_outputs(115) <= b;
    layer0_outputs(116) <= not b;
    layer0_outputs(117) <= not a or b;
    layer0_outputs(118) <= not b;
    layer0_outputs(119) <= not (a or b);
    layer0_outputs(120) <= not (a and b);
    layer0_outputs(121) <= not a;
    layer0_outputs(122) <= a;
    layer0_outputs(123) <= not a;
    layer0_outputs(124) <= not (a and b);
    layer0_outputs(125) <= not b or a;
    layer0_outputs(126) <= not b;
    layer0_outputs(127) <= not a or b;
    layer0_outputs(128) <= not b;
    layer0_outputs(129) <= a xor b;
    layer0_outputs(130) <= not b or a;
    layer0_outputs(131) <= '0';
    layer0_outputs(132) <= not a;
    layer0_outputs(133) <= '0';
    layer0_outputs(134) <= not b;
    layer0_outputs(135) <= a xor b;
    layer0_outputs(136) <= b;
    layer0_outputs(137) <= not (a and b);
    layer0_outputs(138) <= '1';
    layer0_outputs(139) <= a xor b;
    layer0_outputs(140) <= not (a and b);
    layer0_outputs(141) <= not a;
    layer0_outputs(142) <= not (a and b);
    layer0_outputs(143) <= b;
    layer0_outputs(144) <= not b or a;
    layer0_outputs(145) <= not a or b;
    layer0_outputs(146) <= not (a xor b);
    layer0_outputs(147) <= a xor b;
    layer0_outputs(148) <= '0';
    layer0_outputs(149) <= b and not a;
    layer0_outputs(150) <= a or b;
    layer0_outputs(151) <= not (a or b);
    layer0_outputs(152) <= not a or b;
    layer0_outputs(153) <= a and not b;
    layer0_outputs(154) <= a or b;
    layer0_outputs(155) <= a;
    layer0_outputs(156) <= b;
    layer0_outputs(157) <= '1';
    layer0_outputs(158) <= '1';
    layer0_outputs(159) <= '0';
    layer0_outputs(160) <= '0';
    layer0_outputs(161) <= not (a and b);
    layer0_outputs(162) <= not (a and b);
    layer0_outputs(163) <= not b or a;
    layer0_outputs(164) <= a and b;
    layer0_outputs(165) <= a xor b;
    layer0_outputs(166) <= a xor b;
    layer0_outputs(167) <= '0';
    layer0_outputs(168) <= '0';
    layer0_outputs(169) <= a xor b;
    layer0_outputs(170) <= not (a xor b);
    layer0_outputs(171) <= a xor b;
    layer0_outputs(172) <= not (a or b);
    layer0_outputs(173) <= not (a xor b);
    layer0_outputs(174) <= not (a xor b);
    layer0_outputs(175) <= a and b;
    layer0_outputs(176) <= not a;
    layer0_outputs(177) <= a and b;
    layer0_outputs(178) <= not (a or b);
    layer0_outputs(179) <= a or b;
    layer0_outputs(180) <= a;
    layer0_outputs(181) <= b;
    layer0_outputs(182) <= '0';
    layer0_outputs(183) <= a or b;
    layer0_outputs(184) <= not (a and b);
    layer0_outputs(185) <= a and b;
    layer0_outputs(186) <= not a or b;
    layer0_outputs(187) <= not b;
    layer0_outputs(188) <= not (a and b);
    layer0_outputs(189) <= '0';
    layer0_outputs(190) <= b;
    layer0_outputs(191) <= a and b;
    layer0_outputs(192) <= a xor b;
    layer0_outputs(193) <= '0';
    layer0_outputs(194) <= a xor b;
    layer0_outputs(195) <= '1';
    layer0_outputs(196) <= a;
    layer0_outputs(197) <= a;
    layer0_outputs(198) <= b;
    layer0_outputs(199) <= '1';
    layer0_outputs(200) <= b;
    layer0_outputs(201) <= not b;
    layer0_outputs(202) <= a and not b;
    layer0_outputs(203) <= '1';
    layer0_outputs(204) <= not (a or b);
    layer0_outputs(205) <= not (a or b);
    layer0_outputs(206) <= '0';
    layer0_outputs(207) <= b and not a;
    layer0_outputs(208) <= not a;
    layer0_outputs(209) <= not a or b;
    layer0_outputs(210) <= a and not b;
    layer0_outputs(211) <= a;
    layer0_outputs(212) <= a xor b;
    layer0_outputs(213) <= a xor b;
    layer0_outputs(214) <= not b or a;
    layer0_outputs(215) <= '1';
    layer0_outputs(216) <= not (a or b);
    layer0_outputs(217) <= not a;
    layer0_outputs(218) <= '0';
    layer0_outputs(219) <= not (a or b);
    layer0_outputs(220) <= b and not a;
    layer0_outputs(221) <= '0';
    layer0_outputs(222) <= a or b;
    layer0_outputs(223) <= not b or a;
    layer0_outputs(224) <= not b or a;
    layer0_outputs(225) <= a xor b;
    layer0_outputs(226) <= not a;
    layer0_outputs(227) <= not (a xor b);
    layer0_outputs(228) <= not (a or b);
    layer0_outputs(229) <= '0';
    layer0_outputs(230) <= not a;
    layer0_outputs(231) <= a or b;
    layer0_outputs(232) <= a or b;
    layer0_outputs(233) <= not (a and b);
    layer0_outputs(234) <= not b or a;
    layer0_outputs(235) <= '1';
    layer0_outputs(236) <= a or b;
    layer0_outputs(237) <= not b;
    layer0_outputs(238) <= not b or a;
    layer0_outputs(239) <= not b;
    layer0_outputs(240) <= b and not a;
    layer0_outputs(241) <= not (a xor b);
    layer0_outputs(242) <= not a or b;
    layer0_outputs(243) <= a xor b;
    layer0_outputs(244) <= '0';
    layer0_outputs(245) <= a;
    layer0_outputs(246) <= a xor b;
    layer0_outputs(247) <= '0';
    layer0_outputs(248) <= not a or b;
    layer0_outputs(249) <= a xor b;
    layer0_outputs(250) <= '0';
    layer0_outputs(251) <= not (a or b);
    layer0_outputs(252) <= not b;
    layer0_outputs(253) <= '1';
    layer0_outputs(254) <= b and not a;
    layer0_outputs(255) <= not (a or b);
    layer0_outputs(256) <= '1';
    layer0_outputs(257) <= a and b;
    layer0_outputs(258) <= not (a or b);
    layer0_outputs(259) <= a and b;
    layer0_outputs(260) <= a and not b;
    layer0_outputs(261) <= b;
    layer0_outputs(262) <= a and b;
    layer0_outputs(263) <= not a;
    layer0_outputs(264) <= not a or b;
    layer0_outputs(265) <= '0';
    layer0_outputs(266) <= not (a and b);
    layer0_outputs(267) <= '1';
    layer0_outputs(268) <= not b;
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= not b or a;
    layer0_outputs(271) <= not a or b;
    layer0_outputs(272) <= not a or b;
    layer0_outputs(273) <= not a or b;
    layer0_outputs(274) <= a and not b;
    layer0_outputs(275) <= a and b;
    layer0_outputs(276) <= a and not b;
    layer0_outputs(277) <= '1';
    layer0_outputs(278) <= not (a xor b);
    layer0_outputs(279) <= not (a and b);
    layer0_outputs(280) <= a and b;
    layer0_outputs(281) <= not a or b;
    layer0_outputs(282) <= a and b;
    layer0_outputs(283) <= not b;
    layer0_outputs(284) <= a;
    layer0_outputs(285) <= a and b;
    layer0_outputs(286) <= a and b;
    layer0_outputs(287) <= '0';
    layer0_outputs(288) <= not a;
    layer0_outputs(289) <= '1';
    layer0_outputs(290) <= a or b;
    layer0_outputs(291) <= a and b;
    layer0_outputs(292) <= b;
    layer0_outputs(293) <= not a;
    layer0_outputs(294) <= a;
    layer0_outputs(295) <= not (a xor b);
    layer0_outputs(296) <= a or b;
    layer0_outputs(297) <= a and not b;
    layer0_outputs(298) <= not (a xor b);
    layer0_outputs(299) <= not a or b;
    layer0_outputs(300) <= not (a xor b);
    layer0_outputs(301) <= not (a or b);
    layer0_outputs(302) <= a;
    layer0_outputs(303) <= b;
    layer0_outputs(304) <= a;
    layer0_outputs(305) <= a or b;
    layer0_outputs(306) <= a or b;
    layer0_outputs(307) <= a and not b;
    layer0_outputs(308) <= not b;
    layer0_outputs(309) <= not (a and b);
    layer0_outputs(310) <= not (a or b);
    layer0_outputs(311) <= not a or b;
    layer0_outputs(312) <= not b or a;
    layer0_outputs(313) <= a and not b;
    layer0_outputs(314) <= a or b;
    layer0_outputs(315) <= not b;
    layer0_outputs(316) <= a and not b;
    layer0_outputs(317) <= not a or b;
    layer0_outputs(318) <= a;
    layer0_outputs(319) <= a;
    layer0_outputs(320) <= '1';
    layer0_outputs(321) <= b and not a;
    layer0_outputs(322) <= a xor b;
    layer0_outputs(323) <= not (a or b);
    layer0_outputs(324) <= b and not a;
    layer0_outputs(325) <= not (a or b);
    layer0_outputs(326) <= a;
    layer0_outputs(327) <= not a or b;
    layer0_outputs(328) <= a xor b;
    layer0_outputs(329) <= not b;
    layer0_outputs(330) <= not (a or b);
    layer0_outputs(331) <= not (a and b);
    layer0_outputs(332) <= not b;
    layer0_outputs(333) <= '0';
    layer0_outputs(334) <= not b;
    layer0_outputs(335) <= not b or a;
    layer0_outputs(336) <= not (a and b);
    layer0_outputs(337) <= a;
    layer0_outputs(338) <= '1';
    layer0_outputs(339) <= not a or b;
    layer0_outputs(340) <= a or b;
    layer0_outputs(341) <= a;
    layer0_outputs(342) <= b and not a;
    layer0_outputs(343) <= not a;
    layer0_outputs(344) <= not a;
    layer0_outputs(345) <= a and not b;
    layer0_outputs(346) <= '1';
    layer0_outputs(347) <= a and b;
    layer0_outputs(348) <= b and not a;
    layer0_outputs(349) <= not a;
    layer0_outputs(350) <= not (a and b);
    layer0_outputs(351) <= not (a and b);
    layer0_outputs(352) <= a and b;
    layer0_outputs(353) <= not a or b;
    layer0_outputs(354) <= not (a and b);
    layer0_outputs(355) <= a;
    layer0_outputs(356) <= a and b;
    layer0_outputs(357) <= not (a or b);
    layer0_outputs(358) <= not a;
    layer0_outputs(359) <= a;
    layer0_outputs(360) <= a;
    layer0_outputs(361) <= not (a and b);
    layer0_outputs(362) <= not b or a;
    layer0_outputs(363) <= b;
    layer0_outputs(364) <= not a or b;
    layer0_outputs(365) <= not b;
    layer0_outputs(366) <= a or b;
    layer0_outputs(367) <= not (a or b);
    layer0_outputs(368) <= not a;
    layer0_outputs(369) <= not b or a;
    layer0_outputs(370) <= a;
    layer0_outputs(371) <= a and b;
    layer0_outputs(372) <= not (a and b);
    layer0_outputs(373) <= a;
    layer0_outputs(374) <= '1';
    layer0_outputs(375) <= a;
    layer0_outputs(376) <= '0';
    layer0_outputs(377) <= not (a and b);
    layer0_outputs(378) <= not b;
    layer0_outputs(379) <= a;
    layer0_outputs(380) <= not a;
    layer0_outputs(381) <= a and b;
    layer0_outputs(382) <= a and not b;
    layer0_outputs(383) <= not b or a;
    layer0_outputs(384) <= a xor b;
    layer0_outputs(385) <= not b;
    layer0_outputs(386) <= '0';
    layer0_outputs(387) <= a or b;
    layer0_outputs(388) <= b and not a;
    layer0_outputs(389) <= b and not a;
    layer0_outputs(390) <= a and not b;
    layer0_outputs(391) <= not (a xor b);
    layer0_outputs(392) <= not b;
    layer0_outputs(393) <= not (a or b);
    layer0_outputs(394) <= a or b;
    layer0_outputs(395) <= b;
    layer0_outputs(396) <= a and b;
    layer0_outputs(397) <= a and b;
    layer0_outputs(398) <= a;
    layer0_outputs(399) <= a xor b;
    layer0_outputs(400) <= not a;
    layer0_outputs(401) <= a;
    layer0_outputs(402) <= not b or a;
    layer0_outputs(403) <= not (a or b);
    layer0_outputs(404) <= a or b;
    layer0_outputs(405) <= not (a xor b);
    layer0_outputs(406) <= not (a and b);
    layer0_outputs(407) <= not a or b;
    layer0_outputs(408) <= b and not a;
    layer0_outputs(409) <= not b or a;
    layer0_outputs(410) <= '1';
    layer0_outputs(411) <= not b;
    layer0_outputs(412) <= not (a or b);
    layer0_outputs(413) <= not b;
    layer0_outputs(414) <= '0';
    layer0_outputs(415) <= a xor b;
    layer0_outputs(416) <= not b;
    layer0_outputs(417) <= not b or a;
    layer0_outputs(418) <= not (a xor b);
    layer0_outputs(419) <= not a;
    layer0_outputs(420) <= not b;
    layer0_outputs(421) <= not b;
    layer0_outputs(422) <= not a or b;
    layer0_outputs(423) <= not a or b;
    layer0_outputs(424) <= b;
    layer0_outputs(425) <= a or b;
    layer0_outputs(426) <= a;
    layer0_outputs(427) <= not a;
    layer0_outputs(428) <= b;
    layer0_outputs(429) <= not (a xor b);
    layer0_outputs(430) <= a or b;
    layer0_outputs(431) <= '1';
    layer0_outputs(432) <= a;
    layer0_outputs(433) <= not a;
    layer0_outputs(434) <= a xor b;
    layer0_outputs(435) <= not a or b;
    layer0_outputs(436) <= a;
    layer0_outputs(437) <= not a;
    layer0_outputs(438) <= a xor b;
    layer0_outputs(439) <= a xor b;
    layer0_outputs(440) <= a xor b;
    layer0_outputs(441) <= not a or b;
    layer0_outputs(442) <= '1';
    layer0_outputs(443) <= b and not a;
    layer0_outputs(444) <= not (a and b);
    layer0_outputs(445) <= a or b;
    layer0_outputs(446) <= not (a or b);
    layer0_outputs(447) <= not a or b;
    layer0_outputs(448) <= a xor b;
    layer0_outputs(449) <= a and b;
    layer0_outputs(450) <= a and b;
    layer0_outputs(451) <= a and not b;
    layer0_outputs(452) <= a;
    layer0_outputs(453) <= '0';
    layer0_outputs(454) <= a and not b;
    layer0_outputs(455) <= a and not b;
    layer0_outputs(456) <= not a or b;
    layer0_outputs(457) <= b;
    layer0_outputs(458) <= not b or a;
    layer0_outputs(459) <= not b or a;
    layer0_outputs(460) <= not (a or b);
    layer0_outputs(461) <= not a or b;
    layer0_outputs(462) <= not b or a;
    layer0_outputs(463) <= '0';
    layer0_outputs(464) <= a or b;
    layer0_outputs(465) <= not (a xor b);
    layer0_outputs(466) <= a;
    layer0_outputs(467) <= a;
    layer0_outputs(468) <= not a or b;
    layer0_outputs(469) <= '1';
    layer0_outputs(470) <= not b;
    layer0_outputs(471) <= a and not b;
    layer0_outputs(472) <= not a or b;
    layer0_outputs(473) <= not (a or b);
    layer0_outputs(474) <= not (a xor b);
    layer0_outputs(475) <= '1';
    layer0_outputs(476) <= not (a and b);
    layer0_outputs(477) <= a and b;
    layer0_outputs(478) <= not (a xor b);
    layer0_outputs(479) <= a xor b;
    layer0_outputs(480) <= a or b;
    layer0_outputs(481) <= not (a or b);
    layer0_outputs(482) <= not a;
    layer0_outputs(483) <= not a;
    layer0_outputs(484) <= a or b;
    layer0_outputs(485) <= not (a or b);
    layer0_outputs(486) <= a;
    layer0_outputs(487) <= not b;
    layer0_outputs(488) <= a or b;
    layer0_outputs(489) <= not a;
    layer0_outputs(490) <= not a or b;
    layer0_outputs(491) <= b and not a;
    layer0_outputs(492) <= not b;
    layer0_outputs(493) <= not a;
    layer0_outputs(494) <= not b or a;
    layer0_outputs(495) <= a;
    layer0_outputs(496) <= '1';
    layer0_outputs(497) <= '0';
    layer0_outputs(498) <= '1';
    layer0_outputs(499) <= a;
    layer0_outputs(500) <= a xor b;
    layer0_outputs(501) <= not a;
    layer0_outputs(502) <= '0';
    layer0_outputs(503) <= not (a xor b);
    layer0_outputs(504) <= b and not a;
    layer0_outputs(505) <= not b;
    layer0_outputs(506) <= b;
    layer0_outputs(507) <= not a or b;
    layer0_outputs(508) <= a and b;
    layer0_outputs(509) <= b;
    layer0_outputs(510) <= not b;
    layer0_outputs(511) <= not (a xor b);
    layer0_outputs(512) <= '1';
    layer0_outputs(513) <= a and b;
    layer0_outputs(514) <= b and not a;
    layer0_outputs(515) <= '1';
    layer0_outputs(516) <= '0';
    layer0_outputs(517) <= not a or b;
    layer0_outputs(518) <= a or b;
    layer0_outputs(519) <= not b or a;
    layer0_outputs(520) <= not (a and b);
    layer0_outputs(521) <= not b;
    layer0_outputs(522) <= '0';
    layer0_outputs(523) <= a and b;
    layer0_outputs(524) <= b;
    layer0_outputs(525) <= a;
    layer0_outputs(526) <= a and b;
    layer0_outputs(527) <= b and not a;
    layer0_outputs(528) <= a;
    layer0_outputs(529) <= not a or b;
    layer0_outputs(530) <= a;
    layer0_outputs(531) <= a;
    layer0_outputs(532) <= not a or b;
    layer0_outputs(533) <= a;
    layer0_outputs(534) <= '1';
    layer0_outputs(535) <= not b or a;
    layer0_outputs(536) <= a or b;
    layer0_outputs(537) <= b and not a;
    layer0_outputs(538) <= b;
    layer0_outputs(539) <= not (a xor b);
    layer0_outputs(540) <= not (a and b);
    layer0_outputs(541) <= b;
    layer0_outputs(542) <= '1';
    layer0_outputs(543) <= a;
    layer0_outputs(544) <= not a;
    layer0_outputs(545) <= not (a xor b);
    layer0_outputs(546) <= not b;
    layer0_outputs(547) <= '1';
    layer0_outputs(548) <= not a;
    layer0_outputs(549) <= b;
    layer0_outputs(550) <= b and not a;
    layer0_outputs(551) <= not (a or b);
    layer0_outputs(552) <= '0';
    layer0_outputs(553) <= a or b;
    layer0_outputs(554) <= '0';
    layer0_outputs(555) <= not (a xor b);
    layer0_outputs(556) <= b and not a;
    layer0_outputs(557) <= a xor b;
    layer0_outputs(558) <= a and b;
    layer0_outputs(559) <= a or b;
    layer0_outputs(560) <= not b;
    layer0_outputs(561) <= b and not a;
    layer0_outputs(562) <= a or b;
    layer0_outputs(563) <= a and b;
    layer0_outputs(564) <= not b or a;
    layer0_outputs(565) <= not a or b;
    layer0_outputs(566) <= not a;
    layer0_outputs(567) <= b;
    layer0_outputs(568) <= not (a or b);
    layer0_outputs(569) <= a and b;
    layer0_outputs(570) <= not (a or b);
    layer0_outputs(571) <= a or b;
    layer0_outputs(572) <= not (a xor b);
    layer0_outputs(573) <= a and b;
    layer0_outputs(574) <= b;
    layer0_outputs(575) <= not a;
    layer0_outputs(576) <= b;
    layer0_outputs(577) <= b and not a;
    layer0_outputs(578) <= not (a xor b);
    layer0_outputs(579) <= not b;
    layer0_outputs(580) <= not a;
    layer0_outputs(581) <= not a or b;
    layer0_outputs(582) <= a;
    layer0_outputs(583) <= '1';
    layer0_outputs(584) <= '0';
    layer0_outputs(585) <= a xor b;
    layer0_outputs(586) <= not (a or b);
    layer0_outputs(587) <= '0';
    layer0_outputs(588) <= b and not a;
    layer0_outputs(589) <= a or b;
    layer0_outputs(590) <= not b or a;
    layer0_outputs(591) <= not (a or b);
    layer0_outputs(592) <= b;
    layer0_outputs(593) <= not b or a;
    layer0_outputs(594) <= not a;
    layer0_outputs(595) <= not b or a;
    layer0_outputs(596) <= a;
    layer0_outputs(597) <= '0';
    layer0_outputs(598) <= b and not a;
    layer0_outputs(599) <= not (a and b);
    layer0_outputs(600) <= not (a xor b);
    layer0_outputs(601) <= not (a xor b);
    layer0_outputs(602) <= b;
    layer0_outputs(603) <= '1';
    layer0_outputs(604) <= '1';
    layer0_outputs(605) <= not (a or b);
    layer0_outputs(606) <= a;
    layer0_outputs(607) <= a or b;
    layer0_outputs(608) <= '1';
    layer0_outputs(609) <= '0';
    layer0_outputs(610) <= a or b;
    layer0_outputs(611) <= a and b;
    layer0_outputs(612) <= b;
    layer0_outputs(613) <= b;
    layer0_outputs(614) <= not (a and b);
    layer0_outputs(615) <= '1';
    layer0_outputs(616) <= a;
    layer0_outputs(617) <= a and b;
    layer0_outputs(618) <= b and not a;
    layer0_outputs(619) <= not b or a;
    layer0_outputs(620) <= not (a xor b);
    layer0_outputs(621) <= a or b;
    layer0_outputs(622) <= '0';
    layer0_outputs(623) <= a xor b;
    layer0_outputs(624) <= not a;
    layer0_outputs(625) <= '0';
    layer0_outputs(626) <= a xor b;
    layer0_outputs(627) <= a xor b;
    layer0_outputs(628) <= not b or a;
    layer0_outputs(629) <= not b or a;
    layer0_outputs(630) <= not a or b;
    layer0_outputs(631) <= '0';
    layer0_outputs(632) <= a or b;
    layer0_outputs(633) <= b;
    layer0_outputs(634) <= '1';
    layer0_outputs(635) <= not a;
    layer0_outputs(636) <= b;
    layer0_outputs(637) <= b and not a;
    layer0_outputs(638) <= '1';
    layer0_outputs(639) <= a or b;
    layer0_outputs(640) <= '1';
    layer0_outputs(641) <= b and not a;
    layer0_outputs(642) <= '1';
    layer0_outputs(643) <= '0';
    layer0_outputs(644) <= a;
    layer0_outputs(645) <= a;
    layer0_outputs(646) <= '1';
    layer0_outputs(647) <= a;
    layer0_outputs(648) <= a and b;
    layer0_outputs(649) <= '1';
    layer0_outputs(650) <= '0';
    layer0_outputs(651) <= '0';
    layer0_outputs(652) <= b;
    layer0_outputs(653) <= a or b;
    layer0_outputs(654) <= not b;
    layer0_outputs(655) <= a xor b;
    layer0_outputs(656) <= not a;
    layer0_outputs(657) <= b;
    layer0_outputs(658) <= a or b;
    layer0_outputs(659) <= not (a or b);
    layer0_outputs(660) <= a and b;
    layer0_outputs(661) <= not a;
    layer0_outputs(662) <= '1';
    layer0_outputs(663) <= not a or b;
    layer0_outputs(664) <= a;
    layer0_outputs(665) <= '0';
    layer0_outputs(666) <= b and not a;
    layer0_outputs(667) <= a or b;
    layer0_outputs(668) <= not a;
    layer0_outputs(669) <= not (a xor b);
    layer0_outputs(670) <= '0';
    layer0_outputs(671) <= '0';
    layer0_outputs(672) <= '0';
    layer0_outputs(673) <= '1';
    layer0_outputs(674) <= not a or b;
    layer0_outputs(675) <= not b or a;
    layer0_outputs(676) <= not b or a;
    layer0_outputs(677) <= a;
    layer0_outputs(678) <= '1';
    layer0_outputs(679) <= '0';
    layer0_outputs(680) <= not b;
    layer0_outputs(681) <= not a or b;
    layer0_outputs(682) <= b and not a;
    layer0_outputs(683) <= '0';
    layer0_outputs(684) <= a or b;
    layer0_outputs(685) <= a and not b;
    layer0_outputs(686) <= b and not a;
    layer0_outputs(687) <= a xor b;
    layer0_outputs(688) <= a or b;
    layer0_outputs(689) <= a or b;
    layer0_outputs(690) <= '0';
    layer0_outputs(691) <= a and not b;
    layer0_outputs(692) <= not (a xor b);
    layer0_outputs(693) <= a;
    layer0_outputs(694) <= '1';
    layer0_outputs(695) <= not (a and b);
    layer0_outputs(696) <= not (a xor b);
    layer0_outputs(697) <= not a;
    layer0_outputs(698) <= not a;
    layer0_outputs(699) <= not (a or b);
    layer0_outputs(700) <= a;
    layer0_outputs(701) <= '0';
    layer0_outputs(702) <= not (a and b);
    layer0_outputs(703) <= not (a or b);
    layer0_outputs(704) <= not (a xor b);
    layer0_outputs(705) <= not a or b;
    layer0_outputs(706) <= not (a and b);
    layer0_outputs(707) <= not a or b;
    layer0_outputs(708) <= not (a or b);
    layer0_outputs(709) <= not b or a;
    layer0_outputs(710) <= not a or b;
    layer0_outputs(711) <= b and not a;
    layer0_outputs(712) <= not a or b;
    layer0_outputs(713) <= not a or b;
    layer0_outputs(714) <= a and not b;
    layer0_outputs(715) <= a and not b;
    layer0_outputs(716) <= not a;
    layer0_outputs(717) <= not (a or b);
    layer0_outputs(718) <= not b;
    layer0_outputs(719) <= not b or a;
    layer0_outputs(720) <= a and not b;
    layer0_outputs(721) <= not a;
    layer0_outputs(722) <= not b or a;
    layer0_outputs(723) <= b and not a;
    layer0_outputs(724) <= not b or a;
    layer0_outputs(725) <= not (a or b);
    layer0_outputs(726) <= not b or a;
    layer0_outputs(727) <= not (a and b);
    layer0_outputs(728) <= a xor b;
    layer0_outputs(729) <= not a;
    layer0_outputs(730) <= a and not b;
    layer0_outputs(731) <= not (a xor b);
    layer0_outputs(732) <= a or b;
    layer0_outputs(733) <= '0';
    layer0_outputs(734) <= not b or a;
    layer0_outputs(735) <= not a;
    layer0_outputs(736) <= a and b;
    layer0_outputs(737) <= not b or a;
    layer0_outputs(738) <= not a;
    layer0_outputs(739) <= not b;
    layer0_outputs(740) <= a xor b;
    layer0_outputs(741) <= b and not a;
    layer0_outputs(742) <= b and not a;
    layer0_outputs(743) <= not b;
    layer0_outputs(744) <= b and not a;
    layer0_outputs(745) <= not (a or b);
    layer0_outputs(746) <= '1';
    layer0_outputs(747) <= not a;
    layer0_outputs(748) <= b and not a;
    layer0_outputs(749) <= '1';
    layer0_outputs(750) <= not (a or b);
    layer0_outputs(751) <= b and not a;
    layer0_outputs(752) <= b and not a;
    layer0_outputs(753) <= not a or b;
    layer0_outputs(754) <= not (a or b);
    layer0_outputs(755) <= not (a or b);
    layer0_outputs(756) <= not b;
    layer0_outputs(757) <= '0';
    layer0_outputs(758) <= a or b;
    layer0_outputs(759) <= not a or b;
    layer0_outputs(760) <= not (a xor b);
    layer0_outputs(761) <= not (a or b);
    layer0_outputs(762) <= not (a or b);
    layer0_outputs(763) <= not (a and b);
    layer0_outputs(764) <= a or b;
    layer0_outputs(765) <= not b;
    layer0_outputs(766) <= not b;
    layer0_outputs(767) <= not (a or b);
    layer0_outputs(768) <= a and not b;
    layer0_outputs(769) <= not (a and b);
    layer0_outputs(770) <= not b;
    layer0_outputs(771) <= a and not b;
    layer0_outputs(772) <= b;
    layer0_outputs(773) <= a and not b;
    layer0_outputs(774) <= not a;
    layer0_outputs(775) <= a;
    layer0_outputs(776) <= a and b;
    layer0_outputs(777) <= '1';
    layer0_outputs(778) <= not a;
    layer0_outputs(779) <= a or b;
    layer0_outputs(780) <= not a;
    layer0_outputs(781) <= not (a xor b);
    layer0_outputs(782) <= a and not b;
    layer0_outputs(783) <= not (a or b);
    layer0_outputs(784) <= not a;
    layer0_outputs(785) <= a and b;
    layer0_outputs(786) <= b and not a;
    layer0_outputs(787) <= not a or b;
    layer0_outputs(788) <= not b or a;
    layer0_outputs(789) <= a;
    layer0_outputs(790) <= a xor b;
    layer0_outputs(791) <= '0';
    layer0_outputs(792) <= b and not a;
    layer0_outputs(793) <= b and not a;
    layer0_outputs(794) <= '0';
    layer0_outputs(795) <= a or b;
    layer0_outputs(796) <= not (a xor b);
    layer0_outputs(797) <= a xor b;
    layer0_outputs(798) <= not (a and b);
    layer0_outputs(799) <= not a;
    layer0_outputs(800) <= not (a xor b);
    layer0_outputs(801) <= not b or a;
    layer0_outputs(802) <= a and b;
    layer0_outputs(803) <= '1';
    layer0_outputs(804) <= not b;
    layer0_outputs(805) <= '1';
    layer0_outputs(806) <= '1';
    layer0_outputs(807) <= a and not b;
    layer0_outputs(808) <= '0';
    layer0_outputs(809) <= '1';
    layer0_outputs(810) <= a or b;
    layer0_outputs(811) <= a or b;
    layer0_outputs(812) <= not (a or b);
    layer0_outputs(813) <= a and not b;
    layer0_outputs(814) <= a xor b;
    layer0_outputs(815) <= b;
    layer0_outputs(816) <= not (a or b);
    layer0_outputs(817) <= a;
    layer0_outputs(818) <= a;
    layer0_outputs(819) <= not (a xor b);
    layer0_outputs(820) <= b and not a;
    layer0_outputs(821) <= '0';
    layer0_outputs(822) <= not (a and b);
    layer0_outputs(823) <= not (a xor b);
    layer0_outputs(824) <= not b or a;
    layer0_outputs(825) <= b and not a;
    layer0_outputs(826) <= a and b;
    layer0_outputs(827) <= not (a and b);
    layer0_outputs(828) <= not b or a;
    layer0_outputs(829) <= '0';
    layer0_outputs(830) <= not (a or b);
    layer0_outputs(831) <= a and not b;
    layer0_outputs(832) <= not a or b;
    layer0_outputs(833) <= not (a and b);
    layer0_outputs(834) <= '1';
    layer0_outputs(835) <= a and not b;
    layer0_outputs(836) <= not (a or b);
    layer0_outputs(837) <= not a;
    layer0_outputs(838) <= b;
    layer0_outputs(839) <= '0';
    layer0_outputs(840) <= not b or a;
    layer0_outputs(841) <= not a;
    layer0_outputs(842) <= not a or b;
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= not (a or b);
    layer0_outputs(845) <= not (a and b);
    layer0_outputs(846) <= not (a and b);
    layer0_outputs(847) <= not a;
    layer0_outputs(848) <= not (a or b);
    layer0_outputs(849) <= '1';
    layer0_outputs(850) <= not (a and b);
    layer0_outputs(851) <= not a;
    layer0_outputs(852) <= b and not a;
    layer0_outputs(853) <= not (a or b);
    layer0_outputs(854) <= not (a xor b);
    layer0_outputs(855) <= b and not a;
    layer0_outputs(856) <= '0';
    layer0_outputs(857) <= '1';
    layer0_outputs(858) <= a and not b;
    layer0_outputs(859) <= not a;
    layer0_outputs(860) <= not a;
    layer0_outputs(861) <= not (a xor b);
    layer0_outputs(862) <= b and not a;
    layer0_outputs(863) <= a and b;
    layer0_outputs(864) <= b and not a;
    layer0_outputs(865) <= not b or a;
    layer0_outputs(866) <= a;
    layer0_outputs(867) <= '1';
    layer0_outputs(868) <= a xor b;
    layer0_outputs(869) <= not b or a;
    layer0_outputs(870) <= not a or b;
    layer0_outputs(871) <= not b;
    layer0_outputs(872) <= not a;
    layer0_outputs(873) <= '1';
    layer0_outputs(874) <= not b;
    layer0_outputs(875) <= a;
    layer0_outputs(876) <= a or b;
    layer0_outputs(877) <= not (a xor b);
    layer0_outputs(878) <= a;
    layer0_outputs(879) <= not a or b;
    layer0_outputs(880) <= '0';
    layer0_outputs(881) <= b and not a;
    layer0_outputs(882) <= not a;
    layer0_outputs(883) <= a;
    layer0_outputs(884) <= a or b;
    layer0_outputs(885) <= a and b;
    layer0_outputs(886) <= a and b;
    layer0_outputs(887) <= not a or b;
    layer0_outputs(888) <= not a or b;
    layer0_outputs(889) <= '0';
    layer0_outputs(890) <= not b;
    layer0_outputs(891) <= not (a and b);
    layer0_outputs(892) <= b;
    layer0_outputs(893) <= not a;
    layer0_outputs(894) <= a and not b;
    layer0_outputs(895) <= not a or b;
    layer0_outputs(896) <= '1';
    layer0_outputs(897) <= b;
    layer0_outputs(898) <= b;
    layer0_outputs(899) <= not a or b;
    layer0_outputs(900) <= not a or b;
    layer0_outputs(901) <= not (a xor b);
    layer0_outputs(902) <= not a;
    layer0_outputs(903) <= '0';
    layer0_outputs(904) <= b;
    layer0_outputs(905) <= b;
    layer0_outputs(906) <= a or b;
    layer0_outputs(907) <= a and b;
    layer0_outputs(908) <= a and b;
    layer0_outputs(909) <= a and not b;
    layer0_outputs(910) <= b and not a;
    layer0_outputs(911) <= '1';
    layer0_outputs(912) <= not (a or b);
    layer0_outputs(913) <= not (a or b);
    layer0_outputs(914) <= b;
    layer0_outputs(915) <= '0';
    layer0_outputs(916) <= b and not a;
    layer0_outputs(917) <= b;
    layer0_outputs(918) <= not a;
    layer0_outputs(919) <= not (a or b);
    layer0_outputs(920) <= not a or b;
    layer0_outputs(921) <= not a or b;
    layer0_outputs(922) <= b and not a;
    layer0_outputs(923) <= not (a and b);
    layer0_outputs(924) <= not (a or b);
    layer0_outputs(925) <= '0';
    layer0_outputs(926) <= '0';
    layer0_outputs(927) <= a or b;
    layer0_outputs(928) <= not a;
    layer0_outputs(929) <= not (a xor b);
    layer0_outputs(930) <= not a or b;
    layer0_outputs(931) <= not (a and b);
    layer0_outputs(932) <= a and not b;
    layer0_outputs(933) <= not b;
    layer0_outputs(934) <= not b or a;
    layer0_outputs(935) <= a xor b;
    layer0_outputs(936) <= a;
    layer0_outputs(937) <= not a;
    layer0_outputs(938) <= '0';
    layer0_outputs(939) <= a or b;
    layer0_outputs(940) <= not (a xor b);
    layer0_outputs(941) <= not b or a;
    layer0_outputs(942) <= b;
    layer0_outputs(943) <= not (a xor b);
    layer0_outputs(944) <= not a;
    layer0_outputs(945) <= a xor b;
    layer0_outputs(946) <= a and not b;
    layer0_outputs(947) <= not a;
    layer0_outputs(948) <= '1';
    layer0_outputs(949) <= b and not a;
    layer0_outputs(950) <= not (a or b);
    layer0_outputs(951) <= not b or a;
    layer0_outputs(952) <= not a;
    layer0_outputs(953) <= not b;
    layer0_outputs(954) <= '1';
    layer0_outputs(955) <= '0';
    layer0_outputs(956) <= a xor b;
    layer0_outputs(957) <= not (a xor b);
    layer0_outputs(958) <= b;
    layer0_outputs(959) <= not (a or b);
    layer0_outputs(960) <= '0';
    layer0_outputs(961) <= not a;
    layer0_outputs(962) <= not a;
    layer0_outputs(963) <= not (a or b);
    layer0_outputs(964) <= not a;
    layer0_outputs(965) <= a xor b;
    layer0_outputs(966) <= not b or a;
    layer0_outputs(967) <= '0';
    layer0_outputs(968) <= a and not b;
    layer0_outputs(969) <= a;
    layer0_outputs(970) <= b;
    layer0_outputs(971) <= not (a and b);
    layer0_outputs(972) <= a and b;
    layer0_outputs(973) <= '1';
    layer0_outputs(974) <= not b;
    layer0_outputs(975) <= '0';
    layer0_outputs(976) <= not b or a;
    layer0_outputs(977) <= a;
    layer0_outputs(978) <= not (a and b);
    layer0_outputs(979) <= not a;
    layer0_outputs(980) <= a and b;
    layer0_outputs(981) <= b;
    layer0_outputs(982) <= '1';
    layer0_outputs(983) <= a xor b;
    layer0_outputs(984) <= not a or b;
    layer0_outputs(985) <= a and not b;
    layer0_outputs(986) <= a and not b;
    layer0_outputs(987) <= not (a and b);
    layer0_outputs(988) <= a or b;
    layer0_outputs(989) <= '0';
    layer0_outputs(990) <= a and not b;
    layer0_outputs(991) <= a and not b;
    layer0_outputs(992) <= a and b;
    layer0_outputs(993) <= '1';
    layer0_outputs(994) <= a and not b;
    layer0_outputs(995) <= a and b;
    layer0_outputs(996) <= not a or b;
    layer0_outputs(997) <= a and not b;
    layer0_outputs(998) <= b and not a;
    layer0_outputs(999) <= not b;
    layer0_outputs(1000) <= a xor b;
    layer0_outputs(1001) <= a or b;
    layer0_outputs(1002) <= not (a and b);
    layer0_outputs(1003) <= a and not b;
    layer0_outputs(1004) <= a or b;
    layer0_outputs(1005) <= not a;
    layer0_outputs(1006) <= a;
    layer0_outputs(1007) <= '0';
    layer0_outputs(1008) <= a and not b;
    layer0_outputs(1009) <= a xor b;
    layer0_outputs(1010) <= a and not b;
    layer0_outputs(1011) <= a and not b;
    layer0_outputs(1012) <= a and b;
    layer0_outputs(1013) <= '0';
    layer0_outputs(1014) <= not b;
    layer0_outputs(1015) <= a;
    layer0_outputs(1016) <= b and not a;
    layer0_outputs(1017) <= a;
    layer0_outputs(1018) <= not (a or b);
    layer0_outputs(1019) <= a;
    layer0_outputs(1020) <= not (a xor b);
    layer0_outputs(1021) <= '1';
    layer0_outputs(1022) <= not (a and b);
    layer0_outputs(1023) <= a;
    layer0_outputs(1024) <= not a or b;
    layer0_outputs(1025) <= not a or b;
    layer0_outputs(1026) <= not b or a;
    layer0_outputs(1027) <= b;
    layer0_outputs(1028) <= not a or b;
    layer0_outputs(1029) <= not (a or b);
    layer0_outputs(1030) <= b;
    layer0_outputs(1031) <= a and not b;
    layer0_outputs(1032) <= a xor b;
    layer0_outputs(1033) <= b and not a;
    layer0_outputs(1034) <= a xor b;
    layer0_outputs(1035) <= not b or a;
    layer0_outputs(1036) <= not a or b;
    layer0_outputs(1037) <= not a or b;
    layer0_outputs(1038) <= not a;
    layer0_outputs(1039) <= not (a or b);
    layer0_outputs(1040) <= '0';
    layer0_outputs(1041) <= b and not a;
    layer0_outputs(1042) <= '0';
    layer0_outputs(1043) <= a and not b;
    layer0_outputs(1044) <= not (a or b);
    layer0_outputs(1045) <= a xor b;
    layer0_outputs(1046) <= not a;
    layer0_outputs(1047) <= not (a or b);
    layer0_outputs(1048) <= not b or a;
    layer0_outputs(1049) <= not b or a;
    layer0_outputs(1050) <= b;
    layer0_outputs(1051) <= '0';
    layer0_outputs(1052) <= a or b;
    layer0_outputs(1053) <= not a;
    layer0_outputs(1054) <= '0';
    layer0_outputs(1055) <= not a or b;
    layer0_outputs(1056) <= a xor b;
    layer0_outputs(1057) <= not a or b;
    layer0_outputs(1058) <= not a;
    layer0_outputs(1059) <= '1';
    layer0_outputs(1060) <= a and b;
    layer0_outputs(1061) <= not (a or b);
    layer0_outputs(1062) <= not a;
    layer0_outputs(1063) <= not (a xor b);
    layer0_outputs(1064) <= a and b;
    layer0_outputs(1065) <= '0';
    layer0_outputs(1066) <= a xor b;
    layer0_outputs(1067) <= not a;
    layer0_outputs(1068) <= '1';
    layer0_outputs(1069) <= not (a and b);
    layer0_outputs(1070) <= not a or b;
    layer0_outputs(1071) <= '0';
    layer0_outputs(1072) <= '0';
    layer0_outputs(1073) <= a;
    layer0_outputs(1074) <= b and not a;
    layer0_outputs(1075) <= a xor b;
    layer0_outputs(1076) <= b;
    layer0_outputs(1077) <= a or b;
    layer0_outputs(1078) <= not a or b;
    layer0_outputs(1079) <= not (a xor b);
    layer0_outputs(1080) <= '1';
    layer0_outputs(1081) <= a or b;
    layer0_outputs(1082) <= not b or a;
    layer0_outputs(1083) <= not (a xor b);
    layer0_outputs(1084) <= not b;
    layer0_outputs(1085) <= '0';
    layer0_outputs(1086) <= not (a xor b);
    layer0_outputs(1087) <= a xor b;
    layer0_outputs(1088) <= b;
    layer0_outputs(1089) <= a xor b;
    layer0_outputs(1090) <= a xor b;
    layer0_outputs(1091) <= not (a xor b);
    layer0_outputs(1092) <= not b or a;
    layer0_outputs(1093) <= a and not b;
    layer0_outputs(1094) <= '1';
    layer0_outputs(1095) <= a or b;
    layer0_outputs(1096) <= not a or b;
    layer0_outputs(1097) <= '0';
    layer0_outputs(1098) <= not a;
    layer0_outputs(1099) <= '1';
    layer0_outputs(1100) <= a or b;
    layer0_outputs(1101) <= not (a or b);
    layer0_outputs(1102) <= not (a and b);
    layer0_outputs(1103) <= not (a and b);
    layer0_outputs(1104) <= a;
    layer0_outputs(1105) <= '0';
    layer0_outputs(1106) <= a;
    layer0_outputs(1107) <= not a;
    layer0_outputs(1108) <= not (a and b);
    layer0_outputs(1109) <= '1';
    layer0_outputs(1110) <= '1';
    layer0_outputs(1111) <= not a or b;
    layer0_outputs(1112) <= not a;
    layer0_outputs(1113) <= a;
    layer0_outputs(1114) <= a or b;
    layer0_outputs(1115) <= a and not b;
    layer0_outputs(1116) <= a and not b;
    layer0_outputs(1117) <= not (a and b);
    layer0_outputs(1118) <= '1';
    layer0_outputs(1119) <= a xor b;
    layer0_outputs(1120) <= '0';
    layer0_outputs(1121) <= not a;
    layer0_outputs(1122) <= a;
    layer0_outputs(1123) <= not a or b;
    layer0_outputs(1124) <= a and b;
    layer0_outputs(1125) <= not a or b;
    layer0_outputs(1126) <= not (a and b);
    layer0_outputs(1127) <= '0';
    layer0_outputs(1128) <= not (a or b);
    layer0_outputs(1129) <= not a or b;
    layer0_outputs(1130) <= not (a and b);
    layer0_outputs(1131) <= not b or a;
    layer0_outputs(1132) <= a;
    layer0_outputs(1133) <= '0';
    layer0_outputs(1134) <= '1';
    layer0_outputs(1135) <= not a or b;
    layer0_outputs(1136) <= not b or a;
    layer0_outputs(1137) <= not (a xor b);
    layer0_outputs(1138) <= not (a and b);
    layer0_outputs(1139) <= a and not b;
    layer0_outputs(1140) <= b;
    layer0_outputs(1141) <= a and not b;
    layer0_outputs(1142) <= not (a xor b);
    layer0_outputs(1143) <= a;
    layer0_outputs(1144) <= b;
    layer0_outputs(1145) <= a;
    layer0_outputs(1146) <= a and b;
    layer0_outputs(1147) <= not b;
    layer0_outputs(1148) <= '0';
    layer0_outputs(1149) <= '1';
    layer0_outputs(1150) <= a xor b;
    layer0_outputs(1151) <= not (a or b);
    layer0_outputs(1152) <= not b or a;
    layer0_outputs(1153) <= not a;
    layer0_outputs(1154) <= a and b;
    layer0_outputs(1155) <= not b or a;
    layer0_outputs(1156) <= not a;
    layer0_outputs(1157) <= a;
    layer0_outputs(1158) <= a and not b;
    layer0_outputs(1159) <= '0';
    layer0_outputs(1160) <= a xor b;
    layer0_outputs(1161) <= not (a and b);
    layer0_outputs(1162) <= a and b;
    layer0_outputs(1163) <= not b;
    layer0_outputs(1164) <= not (a xor b);
    layer0_outputs(1165) <= not (a or b);
    layer0_outputs(1166) <= not (a xor b);
    layer0_outputs(1167) <= not (a or b);
    layer0_outputs(1168) <= a and not b;
    layer0_outputs(1169) <= not (a xor b);
    layer0_outputs(1170) <= not (a xor b);
    layer0_outputs(1171) <= a;
    layer0_outputs(1172) <= not (a xor b);
    layer0_outputs(1173) <= a or b;
    layer0_outputs(1174) <= not b;
    layer0_outputs(1175) <= a or b;
    layer0_outputs(1176) <= b;
    layer0_outputs(1177) <= a xor b;
    layer0_outputs(1178) <= not b or a;
    layer0_outputs(1179) <= '0';
    layer0_outputs(1180) <= '1';
    layer0_outputs(1181) <= '0';
    layer0_outputs(1182) <= not a;
    layer0_outputs(1183) <= not a;
    layer0_outputs(1184) <= not (a xor b);
    layer0_outputs(1185) <= not (a and b);
    layer0_outputs(1186) <= a or b;
    layer0_outputs(1187) <= not (a and b);
    layer0_outputs(1188) <= '0';
    layer0_outputs(1189) <= a and not b;
    layer0_outputs(1190) <= not a;
    layer0_outputs(1191) <= not a or b;
    layer0_outputs(1192) <= not b;
    layer0_outputs(1193) <= a and b;
    layer0_outputs(1194) <= a xor b;
    layer0_outputs(1195) <= not a or b;
    layer0_outputs(1196) <= a or b;
    layer0_outputs(1197) <= not a or b;
    layer0_outputs(1198) <= not (a or b);
    layer0_outputs(1199) <= '0';
    layer0_outputs(1200) <= a;
    layer0_outputs(1201) <= not a or b;
    layer0_outputs(1202) <= b;
    layer0_outputs(1203) <= not (a or b);
    layer0_outputs(1204) <= a and not b;
    layer0_outputs(1205) <= not (a xor b);
    layer0_outputs(1206) <= not b;
    layer0_outputs(1207) <= not (a and b);
    layer0_outputs(1208) <= '0';
    layer0_outputs(1209) <= a;
    layer0_outputs(1210) <= a xor b;
    layer0_outputs(1211) <= '0';
    layer0_outputs(1212) <= not b;
    layer0_outputs(1213) <= a or b;
    layer0_outputs(1214) <= '1';
    layer0_outputs(1215) <= a and not b;
    layer0_outputs(1216) <= b;
    layer0_outputs(1217) <= not b;
    layer0_outputs(1218) <= not (a xor b);
    layer0_outputs(1219) <= a or b;
    layer0_outputs(1220) <= a or b;
    layer0_outputs(1221) <= not b;
    layer0_outputs(1222) <= not a;
    layer0_outputs(1223) <= a xor b;
    layer0_outputs(1224) <= not b or a;
    layer0_outputs(1225) <= not a or b;
    layer0_outputs(1226) <= a;
    layer0_outputs(1227) <= b;
    layer0_outputs(1228) <= not (a and b);
    layer0_outputs(1229) <= a and not b;
    layer0_outputs(1230) <= a xor b;
    layer0_outputs(1231) <= not b or a;
    layer0_outputs(1232) <= not (a xor b);
    layer0_outputs(1233) <= b and not a;
    layer0_outputs(1234) <= b;
    layer0_outputs(1235) <= a xor b;
    layer0_outputs(1236) <= not (a and b);
    layer0_outputs(1237) <= not (a or b);
    layer0_outputs(1238) <= not a or b;
    layer0_outputs(1239) <= not (a or b);
    layer0_outputs(1240) <= not a or b;
    layer0_outputs(1241) <= not b;
    layer0_outputs(1242) <= a;
    layer0_outputs(1243) <= not a or b;
    layer0_outputs(1244) <= not a or b;
    layer0_outputs(1245) <= a and b;
    layer0_outputs(1246) <= a or b;
    layer0_outputs(1247) <= a;
    layer0_outputs(1248) <= not (a or b);
    layer0_outputs(1249) <= a and not b;
    layer0_outputs(1250) <= a xor b;
    layer0_outputs(1251) <= '0';
    layer0_outputs(1252) <= not (a and b);
    layer0_outputs(1253) <= not b or a;
    layer0_outputs(1254) <= '1';
    layer0_outputs(1255) <= '1';
    layer0_outputs(1256) <= a and not b;
    layer0_outputs(1257) <= a xor b;
    layer0_outputs(1258) <= b and not a;
    layer0_outputs(1259) <= b;
    layer0_outputs(1260) <= not a or b;
    layer0_outputs(1261) <= not b;
    layer0_outputs(1262) <= b and not a;
    layer0_outputs(1263) <= a and not b;
    layer0_outputs(1264) <= b;
    layer0_outputs(1265) <= a and b;
    layer0_outputs(1266) <= not b or a;
    layer0_outputs(1267) <= b;
    layer0_outputs(1268) <= not (a or b);
    layer0_outputs(1269) <= not b;
    layer0_outputs(1270) <= not a;
    layer0_outputs(1271) <= not (a and b);
    layer0_outputs(1272) <= b;
    layer0_outputs(1273) <= a or b;
    layer0_outputs(1274) <= not (a and b);
    layer0_outputs(1275) <= a and b;
    layer0_outputs(1276) <= not a or b;
    layer0_outputs(1277) <= not b;
    layer0_outputs(1278) <= a;
    layer0_outputs(1279) <= b;
    layer0_outputs(1280) <= a or b;
    layer0_outputs(1281) <= '0';
    layer0_outputs(1282) <= '1';
    layer0_outputs(1283) <= '1';
    layer0_outputs(1284) <= not (a and b);
    layer0_outputs(1285) <= not b or a;
    layer0_outputs(1286) <= not (a xor b);
    layer0_outputs(1287) <= not b or a;
    layer0_outputs(1288) <= a xor b;
    layer0_outputs(1289) <= b;
    layer0_outputs(1290) <= not b or a;
    layer0_outputs(1291) <= not b or a;
    layer0_outputs(1292) <= a and b;
    layer0_outputs(1293) <= not (a or b);
    layer0_outputs(1294) <= not (a xor b);
    layer0_outputs(1295) <= a or b;
    layer0_outputs(1296) <= a and not b;
    layer0_outputs(1297) <= not a;
    layer0_outputs(1298) <= a;
    layer0_outputs(1299) <= a xor b;
    layer0_outputs(1300) <= not b;
    layer0_outputs(1301) <= not (a or b);
    layer0_outputs(1302) <= a or b;
    layer0_outputs(1303) <= not a or b;
    layer0_outputs(1304) <= not (a or b);
    layer0_outputs(1305) <= a or b;
    layer0_outputs(1306) <= a and b;
    layer0_outputs(1307) <= not (a and b);
    layer0_outputs(1308) <= '1';
    layer0_outputs(1309) <= '1';
    layer0_outputs(1310) <= not b or a;
    layer0_outputs(1311) <= not a;
    layer0_outputs(1312) <= a xor b;
    layer0_outputs(1313) <= not (a or b);
    layer0_outputs(1314) <= a;
    layer0_outputs(1315) <= b;
    layer0_outputs(1316) <= not b;
    layer0_outputs(1317) <= not (a and b);
    layer0_outputs(1318) <= '1';
    layer0_outputs(1319) <= b;
    layer0_outputs(1320) <= b and not a;
    layer0_outputs(1321) <= a and not b;
    layer0_outputs(1322) <= '0';
    layer0_outputs(1323) <= not a or b;
    layer0_outputs(1324) <= not a or b;
    layer0_outputs(1325) <= b;
    layer0_outputs(1326) <= b and not a;
    layer0_outputs(1327) <= '1';
    layer0_outputs(1328) <= not b;
    layer0_outputs(1329) <= a or b;
    layer0_outputs(1330) <= not b;
    layer0_outputs(1331) <= not (a or b);
    layer0_outputs(1332) <= b and not a;
    layer0_outputs(1333) <= not b;
    layer0_outputs(1334) <= '0';
    layer0_outputs(1335) <= not (a or b);
    layer0_outputs(1336) <= '0';
    layer0_outputs(1337) <= not (a xor b);
    layer0_outputs(1338) <= not b;
    layer0_outputs(1339) <= b and not a;
    layer0_outputs(1340) <= not b or a;
    layer0_outputs(1341) <= '1';
    layer0_outputs(1342) <= not (a and b);
    layer0_outputs(1343) <= a or b;
    layer0_outputs(1344) <= not b;
    layer0_outputs(1345) <= a and not b;
    layer0_outputs(1346) <= '0';
    layer0_outputs(1347) <= not (a xor b);
    layer0_outputs(1348) <= not (a and b);
    layer0_outputs(1349) <= not (a or b);
    layer0_outputs(1350) <= b;
    layer0_outputs(1351) <= '1';
    layer0_outputs(1352) <= not (a and b);
    layer0_outputs(1353) <= a xor b;
    layer0_outputs(1354) <= a and b;
    layer0_outputs(1355) <= not a;
    layer0_outputs(1356) <= not b;
    layer0_outputs(1357) <= '1';
    layer0_outputs(1358) <= not a;
    layer0_outputs(1359) <= '0';
    layer0_outputs(1360) <= not b or a;
    layer0_outputs(1361) <= a or b;
    layer0_outputs(1362) <= '0';
    layer0_outputs(1363) <= not b or a;
    layer0_outputs(1364) <= not a;
    layer0_outputs(1365) <= a or b;
    layer0_outputs(1366) <= not (a or b);
    layer0_outputs(1367) <= a and not b;
    layer0_outputs(1368) <= b and not a;
    layer0_outputs(1369) <= not a;
    layer0_outputs(1370) <= not (a and b);
    layer0_outputs(1371) <= '1';
    layer0_outputs(1372) <= not b;
    layer0_outputs(1373) <= not b or a;
    layer0_outputs(1374) <= not b;
    layer0_outputs(1375) <= '1';
    layer0_outputs(1376) <= a or b;
    layer0_outputs(1377) <= '1';
    layer0_outputs(1378) <= a or b;
    layer0_outputs(1379) <= not (a xor b);
    layer0_outputs(1380) <= not (a or b);
    layer0_outputs(1381) <= b;
    layer0_outputs(1382) <= a;
    layer0_outputs(1383) <= not b;
    layer0_outputs(1384) <= b;
    layer0_outputs(1385) <= a or b;
    layer0_outputs(1386) <= not a;
    layer0_outputs(1387) <= '1';
    layer0_outputs(1388) <= '1';
    layer0_outputs(1389) <= not (a or b);
    layer0_outputs(1390) <= not a;
    layer0_outputs(1391) <= not b or a;
    layer0_outputs(1392) <= not b;
    layer0_outputs(1393) <= not a;
    layer0_outputs(1394) <= not (a or b);
    layer0_outputs(1395) <= '1';
    layer0_outputs(1396) <= not b;
    layer0_outputs(1397) <= not (a xor b);
    layer0_outputs(1398) <= b;
    layer0_outputs(1399) <= not b;
    layer0_outputs(1400) <= a and not b;
    layer0_outputs(1401) <= a and not b;
    layer0_outputs(1402) <= a and not b;
    layer0_outputs(1403) <= a and not b;
    layer0_outputs(1404) <= b and not a;
    layer0_outputs(1405) <= not b;
    layer0_outputs(1406) <= a;
    layer0_outputs(1407) <= b;
    layer0_outputs(1408) <= a and not b;
    layer0_outputs(1409) <= b;
    layer0_outputs(1410) <= a;
    layer0_outputs(1411) <= b and not a;
    layer0_outputs(1412) <= '1';
    layer0_outputs(1413) <= not b;
    layer0_outputs(1414) <= '0';
    layer0_outputs(1415) <= '0';
    layer0_outputs(1416) <= not (a and b);
    layer0_outputs(1417) <= a or b;
    layer0_outputs(1418) <= a or b;
    layer0_outputs(1419) <= b;
    layer0_outputs(1420) <= '1';
    layer0_outputs(1421) <= '0';
    layer0_outputs(1422) <= a;
    layer0_outputs(1423) <= not (a xor b);
    layer0_outputs(1424) <= not a;
    layer0_outputs(1425) <= '0';
    layer0_outputs(1426) <= '1';
    layer0_outputs(1427) <= not b or a;
    layer0_outputs(1428) <= not (a or b);
    layer0_outputs(1429) <= a and not b;
    layer0_outputs(1430) <= a and b;
    layer0_outputs(1431) <= not a or b;
    layer0_outputs(1432) <= b;
    layer0_outputs(1433) <= '0';
    layer0_outputs(1434) <= not a;
    layer0_outputs(1435) <= a;
    layer0_outputs(1436) <= '0';
    layer0_outputs(1437) <= not a or b;
    layer0_outputs(1438) <= not (a and b);
    layer0_outputs(1439) <= '0';
    layer0_outputs(1440) <= b and not a;
    layer0_outputs(1441) <= not (a and b);
    layer0_outputs(1442) <= not a or b;
    layer0_outputs(1443) <= not (a xor b);
    layer0_outputs(1444) <= not b;
    layer0_outputs(1445) <= not a;
    layer0_outputs(1446) <= not b;
    layer0_outputs(1447) <= a;
    layer0_outputs(1448) <= not b or a;
    layer0_outputs(1449) <= not a;
    layer0_outputs(1450) <= a and not b;
    layer0_outputs(1451) <= '1';
    layer0_outputs(1452) <= a and not b;
    layer0_outputs(1453) <= not a;
    layer0_outputs(1454) <= '0';
    layer0_outputs(1455) <= not a or b;
    layer0_outputs(1456) <= a;
    layer0_outputs(1457) <= '1';
    layer0_outputs(1458) <= not (a or b);
    layer0_outputs(1459) <= not b;
    layer0_outputs(1460) <= not (a or b);
    layer0_outputs(1461) <= not a;
    layer0_outputs(1462) <= '1';
    layer0_outputs(1463) <= '0';
    layer0_outputs(1464) <= not (a and b);
    layer0_outputs(1465) <= a;
    layer0_outputs(1466) <= not a;
    layer0_outputs(1467) <= b;
    layer0_outputs(1468) <= b;
    layer0_outputs(1469) <= not (a or b);
    layer0_outputs(1470) <= not a or b;
    layer0_outputs(1471) <= not b;
    layer0_outputs(1472) <= b;
    layer0_outputs(1473) <= a;
    layer0_outputs(1474) <= not b or a;
    layer0_outputs(1475) <= a and b;
    layer0_outputs(1476) <= not (a xor b);
    layer0_outputs(1477) <= a;
    layer0_outputs(1478) <= not (a and b);
    layer0_outputs(1479) <= not a or b;
    layer0_outputs(1480) <= not (a or b);
    layer0_outputs(1481) <= a and b;
    layer0_outputs(1482) <= b and not a;
    layer0_outputs(1483) <= not (a and b);
    layer0_outputs(1484) <= not (a and b);
    layer0_outputs(1485) <= b;
    layer0_outputs(1486) <= b and not a;
    layer0_outputs(1487) <= not (a or b);
    layer0_outputs(1488) <= not (a and b);
    layer0_outputs(1489) <= not b or a;
    layer0_outputs(1490) <= '0';
    layer0_outputs(1491) <= '0';
    layer0_outputs(1492) <= not a or b;
    layer0_outputs(1493) <= a and b;
    layer0_outputs(1494) <= not b or a;
    layer0_outputs(1495) <= a or b;
    layer0_outputs(1496) <= not (a xor b);
    layer0_outputs(1497) <= not (a and b);
    layer0_outputs(1498) <= '0';
    layer0_outputs(1499) <= a and not b;
    layer0_outputs(1500) <= '1';
    layer0_outputs(1501) <= a or b;
    layer0_outputs(1502) <= '1';
    layer0_outputs(1503) <= a or b;
    layer0_outputs(1504) <= a and not b;
    layer0_outputs(1505) <= '0';
    layer0_outputs(1506) <= not b or a;
    layer0_outputs(1507) <= not a;
    layer0_outputs(1508) <= not b or a;
    layer0_outputs(1509) <= b and not a;
    layer0_outputs(1510) <= a and not b;
    layer0_outputs(1511) <= '0';
    layer0_outputs(1512) <= not (a or b);
    layer0_outputs(1513) <= a;
    layer0_outputs(1514) <= not (a and b);
    layer0_outputs(1515) <= a;
    layer0_outputs(1516) <= a and not b;
    layer0_outputs(1517) <= a or b;
    layer0_outputs(1518) <= '1';
    layer0_outputs(1519) <= not (a or b);
    layer0_outputs(1520) <= b;
    layer0_outputs(1521) <= not (a and b);
    layer0_outputs(1522) <= a or b;
    layer0_outputs(1523) <= a or b;
    layer0_outputs(1524) <= not b or a;
    layer0_outputs(1525) <= not b or a;
    layer0_outputs(1526) <= not (a xor b);
    layer0_outputs(1527) <= not b or a;
    layer0_outputs(1528) <= not (a and b);
    layer0_outputs(1529) <= '0';
    layer0_outputs(1530) <= a;
    layer0_outputs(1531) <= not (a or b);
    layer0_outputs(1532) <= '0';
    layer0_outputs(1533) <= a and b;
    layer0_outputs(1534) <= a and b;
    layer0_outputs(1535) <= '1';
    layer0_outputs(1536) <= not (a or b);
    layer0_outputs(1537) <= '1';
    layer0_outputs(1538) <= b and not a;
    layer0_outputs(1539) <= not b;
    layer0_outputs(1540) <= a xor b;
    layer0_outputs(1541) <= not b;
    layer0_outputs(1542) <= not a;
    layer0_outputs(1543) <= '0';
    layer0_outputs(1544) <= '0';
    layer0_outputs(1545) <= not (a and b);
    layer0_outputs(1546) <= not (a and b);
    layer0_outputs(1547) <= '0';
    layer0_outputs(1548) <= not (a or b);
    layer0_outputs(1549) <= a or b;
    layer0_outputs(1550) <= not a or b;
    layer0_outputs(1551) <= a and not b;
    layer0_outputs(1552) <= not b or a;
    layer0_outputs(1553) <= a and not b;
    layer0_outputs(1554) <= not a;
    layer0_outputs(1555) <= a or b;
    layer0_outputs(1556) <= a or b;
    layer0_outputs(1557) <= not a;
    layer0_outputs(1558) <= a xor b;
    layer0_outputs(1559) <= not a;
    layer0_outputs(1560) <= not a;
    layer0_outputs(1561) <= a or b;
    layer0_outputs(1562) <= not b or a;
    layer0_outputs(1563) <= a;
    layer0_outputs(1564) <= a or b;
    layer0_outputs(1565) <= a and not b;
    layer0_outputs(1566) <= '0';
    layer0_outputs(1567) <= not a or b;
    layer0_outputs(1568) <= not (a xor b);
    layer0_outputs(1569) <= a and not b;
    layer0_outputs(1570) <= a xor b;
    layer0_outputs(1571) <= not (a and b);
    layer0_outputs(1572) <= '1';
    layer0_outputs(1573) <= a or b;
    layer0_outputs(1574) <= a;
    layer0_outputs(1575) <= not (a and b);
    layer0_outputs(1576) <= not b;
    layer0_outputs(1577) <= '0';
    layer0_outputs(1578) <= a xor b;
    layer0_outputs(1579) <= a and b;
    layer0_outputs(1580) <= not (a and b);
    layer0_outputs(1581) <= not b or a;
    layer0_outputs(1582) <= b;
    layer0_outputs(1583) <= '1';
    layer0_outputs(1584) <= not (a and b);
    layer0_outputs(1585) <= not b;
    layer0_outputs(1586) <= not (a or b);
    layer0_outputs(1587) <= not a;
    layer0_outputs(1588) <= not a or b;
    layer0_outputs(1589) <= not a or b;
    layer0_outputs(1590) <= a;
    layer0_outputs(1591) <= a xor b;
    layer0_outputs(1592) <= not a;
    layer0_outputs(1593) <= a and not b;
    layer0_outputs(1594) <= b;
    layer0_outputs(1595) <= not (a and b);
    layer0_outputs(1596) <= not a;
    layer0_outputs(1597) <= '0';
    layer0_outputs(1598) <= not (a or b);
    layer0_outputs(1599) <= a xor b;
    layer0_outputs(1600) <= b;
    layer0_outputs(1601) <= '0';
    layer0_outputs(1602) <= not b or a;
    layer0_outputs(1603) <= a xor b;
    layer0_outputs(1604) <= '0';
    layer0_outputs(1605) <= '0';
    layer0_outputs(1606) <= not b;
    layer0_outputs(1607) <= a and not b;
    layer0_outputs(1608) <= '1';
    layer0_outputs(1609) <= '1';
    layer0_outputs(1610) <= not a or b;
    layer0_outputs(1611) <= a xor b;
    layer0_outputs(1612) <= a and not b;
    layer0_outputs(1613) <= not a or b;
    layer0_outputs(1614) <= not b or a;
    layer0_outputs(1615) <= b;
    layer0_outputs(1616) <= a and not b;
    layer0_outputs(1617) <= a;
    layer0_outputs(1618) <= not (a and b);
    layer0_outputs(1619) <= a and not b;
    layer0_outputs(1620) <= '0';
    layer0_outputs(1621) <= a and not b;
    layer0_outputs(1622) <= b;
    layer0_outputs(1623) <= a and not b;
    layer0_outputs(1624) <= '0';
    layer0_outputs(1625) <= b and not a;
    layer0_outputs(1626) <= not a or b;
    layer0_outputs(1627) <= not (a or b);
    layer0_outputs(1628) <= b;
    layer0_outputs(1629) <= not (a and b);
    layer0_outputs(1630) <= not a or b;
    layer0_outputs(1631) <= a and not b;
    layer0_outputs(1632) <= not b or a;
    layer0_outputs(1633) <= not (a or b);
    layer0_outputs(1634) <= not a;
    layer0_outputs(1635) <= a and b;
    layer0_outputs(1636) <= a;
    layer0_outputs(1637) <= not (a or b);
    layer0_outputs(1638) <= b;
    layer0_outputs(1639) <= '0';
    layer0_outputs(1640) <= not (a or b);
    layer0_outputs(1641) <= not a;
    layer0_outputs(1642) <= '1';
    layer0_outputs(1643) <= a or b;
    layer0_outputs(1644) <= not (a and b);
    layer0_outputs(1645) <= a;
    layer0_outputs(1646) <= a and not b;
    layer0_outputs(1647) <= a and not b;
    layer0_outputs(1648) <= a;
    layer0_outputs(1649) <= not (a and b);
    layer0_outputs(1650) <= not b or a;
    layer0_outputs(1651) <= not (a or b);
    layer0_outputs(1652) <= a and not b;
    layer0_outputs(1653) <= b;
    layer0_outputs(1654) <= not (a and b);
    layer0_outputs(1655) <= a or b;
    layer0_outputs(1656) <= a or b;
    layer0_outputs(1657) <= not (a or b);
    layer0_outputs(1658) <= a and not b;
    layer0_outputs(1659) <= '1';
    layer0_outputs(1660) <= not (a or b);
    layer0_outputs(1661) <= not a or b;
    layer0_outputs(1662) <= a and not b;
    layer0_outputs(1663) <= a and not b;
    layer0_outputs(1664) <= a and b;
    layer0_outputs(1665) <= not a or b;
    layer0_outputs(1666) <= not (a and b);
    layer0_outputs(1667) <= a and b;
    layer0_outputs(1668) <= '1';
    layer0_outputs(1669) <= not (a or b);
    layer0_outputs(1670) <= not a or b;
    layer0_outputs(1671) <= '0';
    layer0_outputs(1672) <= not b or a;
    layer0_outputs(1673) <= not b;
    layer0_outputs(1674) <= not (a or b);
    layer0_outputs(1675) <= a or b;
    layer0_outputs(1676) <= not a or b;
    layer0_outputs(1677) <= a and not b;
    layer0_outputs(1678) <= '1';
    layer0_outputs(1679) <= not a;
    layer0_outputs(1680) <= not a or b;
    layer0_outputs(1681) <= '0';
    layer0_outputs(1682) <= b and not a;
    layer0_outputs(1683) <= not (a xor b);
    layer0_outputs(1684) <= not a or b;
    layer0_outputs(1685) <= not (a or b);
    layer0_outputs(1686) <= not (a and b);
    layer0_outputs(1687) <= not (a and b);
    layer0_outputs(1688) <= a or b;
    layer0_outputs(1689) <= not (a and b);
    layer0_outputs(1690) <= '1';
    layer0_outputs(1691) <= '0';
    layer0_outputs(1692) <= not a;
    layer0_outputs(1693) <= a and not b;
    layer0_outputs(1694) <= a or b;
    layer0_outputs(1695) <= not a;
    layer0_outputs(1696) <= not a;
    layer0_outputs(1697) <= b;
    layer0_outputs(1698) <= '1';
    layer0_outputs(1699) <= b and not a;
    layer0_outputs(1700) <= a and not b;
    layer0_outputs(1701) <= a;
    layer0_outputs(1702) <= a and b;
    layer0_outputs(1703) <= '0';
    layer0_outputs(1704) <= a or b;
    layer0_outputs(1705) <= a;
    layer0_outputs(1706) <= not a or b;
    layer0_outputs(1707) <= a;
    layer0_outputs(1708) <= not (a xor b);
    layer0_outputs(1709) <= not b;
    layer0_outputs(1710) <= a;
    layer0_outputs(1711) <= '0';
    layer0_outputs(1712) <= a and b;
    layer0_outputs(1713) <= a or b;
    layer0_outputs(1714) <= not b or a;
    layer0_outputs(1715) <= a;
    layer0_outputs(1716) <= '1';
    layer0_outputs(1717) <= a;
    layer0_outputs(1718) <= b and not a;
    layer0_outputs(1719) <= not a or b;
    layer0_outputs(1720) <= not (a xor b);
    layer0_outputs(1721) <= not (a or b);
    layer0_outputs(1722) <= '1';
    layer0_outputs(1723) <= not a or b;
    layer0_outputs(1724) <= '1';
    layer0_outputs(1725) <= not a;
    layer0_outputs(1726) <= a xor b;
    layer0_outputs(1727) <= b and not a;
    layer0_outputs(1728) <= a xor b;
    layer0_outputs(1729) <= not (a and b);
    layer0_outputs(1730) <= a xor b;
    layer0_outputs(1731) <= b;
    layer0_outputs(1732) <= not b;
    layer0_outputs(1733) <= not (a and b);
    layer0_outputs(1734) <= not b;
    layer0_outputs(1735) <= '1';
    layer0_outputs(1736) <= a and b;
    layer0_outputs(1737) <= a or b;
    layer0_outputs(1738) <= b;
    layer0_outputs(1739) <= a and b;
    layer0_outputs(1740) <= '1';
    layer0_outputs(1741) <= '0';
    layer0_outputs(1742) <= a xor b;
    layer0_outputs(1743) <= a and b;
    layer0_outputs(1744) <= not (a and b);
    layer0_outputs(1745) <= a;
    layer0_outputs(1746) <= not a or b;
    layer0_outputs(1747) <= '1';
    layer0_outputs(1748) <= a;
    layer0_outputs(1749) <= a;
    layer0_outputs(1750) <= not a or b;
    layer0_outputs(1751) <= a and not b;
    layer0_outputs(1752) <= a or b;
    layer0_outputs(1753) <= '1';
    layer0_outputs(1754) <= a;
    layer0_outputs(1755) <= b and not a;
    layer0_outputs(1756) <= '0';
    layer0_outputs(1757) <= a or b;
    layer0_outputs(1758) <= a or b;
    layer0_outputs(1759) <= not a or b;
    layer0_outputs(1760) <= not (a xor b);
    layer0_outputs(1761) <= a or b;
    layer0_outputs(1762) <= not a;
    layer0_outputs(1763) <= a and b;
    layer0_outputs(1764) <= not b;
    layer0_outputs(1765) <= b;
    layer0_outputs(1766) <= not b;
    layer0_outputs(1767) <= a and b;
    layer0_outputs(1768) <= not (a xor b);
    layer0_outputs(1769) <= a and b;
    layer0_outputs(1770) <= not (a and b);
    layer0_outputs(1771) <= a and b;
    layer0_outputs(1772) <= '0';
    layer0_outputs(1773) <= not (a or b);
    layer0_outputs(1774) <= not (a xor b);
    layer0_outputs(1775) <= not b or a;
    layer0_outputs(1776) <= '1';
    layer0_outputs(1777) <= not b or a;
    layer0_outputs(1778) <= a and b;
    layer0_outputs(1779) <= not (a and b);
    layer0_outputs(1780) <= '1';
    layer0_outputs(1781) <= a and not b;
    layer0_outputs(1782) <= '1';
    layer0_outputs(1783) <= not a or b;
    layer0_outputs(1784) <= a or b;
    layer0_outputs(1785) <= '1';
    layer0_outputs(1786) <= not (a or b);
    layer0_outputs(1787) <= not (a and b);
    layer0_outputs(1788) <= a and not b;
    layer0_outputs(1789) <= a and b;
    layer0_outputs(1790) <= a xor b;
    layer0_outputs(1791) <= not (a and b);
    layer0_outputs(1792) <= a and not b;
    layer0_outputs(1793) <= not b;
    layer0_outputs(1794) <= a or b;
    layer0_outputs(1795) <= a xor b;
    layer0_outputs(1796) <= '1';
    layer0_outputs(1797) <= not a or b;
    layer0_outputs(1798) <= a and not b;
    layer0_outputs(1799) <= b;
    layer0_outputs(1800) <= not (a or b);
    layer0_outputs(1801) <= not (a xor b);
    layer0_outputs(1802) <= not (a or b);
    layer0_outputs(1803) <= a and b;
    layer0_outputs(1804) <= a xor b;
    layer0_outputs(1805) <= a;
    layer0_outputs(1806) <= a and not b;
    layer0_outputs(1807) <= a and not b;
    layer0_outputs(1808) <= a xor b;
    layer0_outputs(1809) <= not a or b;
    layer0_outputs(1810) <= a;
    layer0_outputs(1811) <= not a;
    layer0_outputs(1812) <= not b or a;
    layer0_outputs(1813) <= not (a or b);
    layer0_outputs(1814) <= b;
    layer0_outputs(1815) <= '0';
    layer0_outputs(1816) <= b and not a;
    layer0_outputs(1817) <= not b or a;
    layer0_outputs(1818) <= b and not a;
    layer0_outputs(1819) <= '1';
    layer0_outputs(1820) <= '0';
    layer0_outputs(1821) <= not b or a;
    layer0_outputs(1822) <= b;
    layer0_outputs(1823) <= not a;
    layer0_outputs(1824) <= a and b;
    layer0_outputs(1825) <= b and not a;
    layer0_outputs(1826) <= not (a and b);
    layer0_outputs(1827) <= a or b;
    layer0_outputs(1828) <= a and not b;
    layer0_outputs(1829) <= a and not b;
    layer0_outputs(1830) <= b and not a;
    layer0_outputs(1831) <= a and b;
    layer0_outputs(1832) <= not b or a;
    layer0_outputs(1833) <= not b or a;
    layer0_outputs(1834) <= not b or a;
    layer0_outputs(1835) <= a and not b;
    layer0_outputs(1836) <= not a;
    layer0_outputs(1837) <= a xor b;
    layer0_outputs(1838) <= '1';
    layer0_outputs(1839) <= not a or b;
    layer0_outputs(1840) <= b and not a;
    layer0_outputs(1841) <= a or b;
    layer0_outputs(1842) <= not b;
    layer0_outputs(1843) <= '0';
    layer0_outputs(1844) <= a or b;
    layer0_outputs(1845) <= not b or a;
    layer0_outputs(1846) <= a xor b;
    layer0_outputs(1847) <= a or b;
    layer0_outputs(1848) <= '1';
    layer0_outputs(1849) <= '0';
    layer0_outputs(1850) <= b;
    layer0_outputs(1851) <= not a;
    layer0_outputs(1852) <= a and not b;
    layer0_outputs(1853) <= not (a or b);
    layer0_outputs(1854) <= not (a and b);
    layer0_outputs(1855) <= not (a or b);
    layer0_outputs(1856) <= a;
    layer0_outputs(1857) <= b and not a;
    layer0_outputs(1858) <= a and not b;
    layer0_outputs(1859) <= not a or b;
    layer0_outputs(1860) <= a or b;
    layer0_outputs(1861) <= b;
    layer0_outputs(1862) <= not (a and b);
    layer0_outputs(1863) <= not a or b;
    layer0_outputs(1864) <= not a;
    layer0_outputs(1865) <= not (a and b);
    layer0_outputs(1866) <= '0';
    layer0_outputs(1867) <= '1';
    layer0_outputs(1868) <= not (a or b);
    layer0_outputs(1869) <= a and b;
    layer0_outputs(1870) <= not a or b;
    layer0_outputs(1871) <= not b or a;
    layer0_outputs(1872) <= b;
    layer0_outputs(1873) <= a;
    layer0_outputs(1874) <= not (a and b);
    layer0_outputs(1875) <= not (a xor b);
    layer0_outputs(1876) <= a xor b;
    layer0_outputs(1877) <= not a or b;
    layer0_outputs(1878) <= b;
    layer0_outputs(1879) <= b;
    layer0_outputs(1880) <= not (a or b);
    layer0_outputs(1881) <= '0';
    layer0_outputs(1882) <= not b or a;
    layer0_outputs(1883) <= not b;
    layer0_outputs(1884) <= not b;
    layer0_outputs(1885) <= not b;
    layer0_outputs(1886) <= a or b;
    layer0_outputs(1887) <= not (a or b);
    layer0_outputs(1888) <= not (a and b);
    layer0_outputs(1889) <= '1';
    layer0_outputs(1890) <= not a or b;
    layer0_outputs(1891) <= a and b;
    layer0_outputs(1892) <= '1';
    layer0_outputs(1893) <= a and b;
    layer0_outputs(1894) <= a xor b;
    layer0_outputs(1895) <= '0';
    layer0_outputs(1896) <= '1';
    layer0_outputs(1897) <= a and b;
    layer0_outputs(1898) <= a and b;
    layer0_outputs(1899) <= not a or b;
    layer0_outputs(1900) <= not a;
    layer0_outputs(1901) <= '0';
    layer0_outputs(1902) <= a or b;
    layer0_outputs(1903) <= not (a or b);
    layer0_outputs(1904) <= not (a xor b);
    layer0_outputs(1905) <= a and b;
    layer0_outputs(1906) <= not a;
    layer0_outputs(1907) <= not b;
    layer0_outputs(1908) <= a and not b;
    layer0_outputs(1909) <= '1';
    layer0_outputs(1910) <= '1';
    layer0_outputs(1911) <= '0';
    layer0_outputs(1912) <= not (a or b);
    layer0_outputs(1913) <= a xor b;
    layer0_outputs(1914) <= not (a and b);
    layer0_outputs(1915) <= a;
    layer0_outputs(1916) <= not (a or b);
    layer0_outputs(1917) <= not b or a;
    layer0_outputs(1918) <= a and b;
    layer0_outputs(1919) <= not (a and b);
    layer0_outputs(1920) <= '0';
    layer0_outputs(1921) <= not b;
    layer0_outputs(1922) <= not b;
    layer0_outputs(1923) <= b and not a;
    layer0_outputs(1924) <= b and not a;
    layer0_outputs(1925) <= b;
    layer0_outputs(1926) <= '1';
    layer0_outputs(1927) <= b and not a;
    layer0_outputs(1928) <= '1';
    layer0_outputs(1929) <= not a or b;
    layer0_outputs(1930) <= a and b;
    layer0_outputs(1931) <= not b;
    layer0_outputs(1932) <= a;
    layer0_outputs(1933) <= not (a xor b);
    layer0_outputs(1934) <= not b or a;
    layer0_outputs(1935) <= a and b;
    layer0_outputs(1936) <= a and b;
    layer0_outputs(1937) <= a and not b;
    layer0_outputs(1938) <= not b or a;
    layer0_outputs(1939) <= not (a or b);
    layer0_outputs(1940) <= a and b;
    layer0_outputs(1941) <= '1';
    layer0_outputs(1942) <= not b or a;
    layer0_outputs(1943) <= b and not a;
    layer0_outputs(1944) <= a;
    layer0_outputs(1945) <= not b or a;
    layer0_outputs(1946) <= a and b;
    layer0_outputs(1947) <= a;
    layer0_outputs(1948) <= a and not b;
    layer0_outputs(1949) <= not b or a;
    layer0_outputs(1950) <= not (a or b);
    layer0_outputs(1951) <= a;
    layer0_outputs(1952) <= b;
    layer0_outputs(1953) <= not a;
    layer0_outputs(1954) <= not (a and b);
    layer0_outputs(1955) <= a and not b;
    layer0_outputs(1956) <= not a or b;
    layer0_outputs(1957) <= not (a or b);
    layer0_outputs(1958) <= a;
    layer0_outputs(1959) <= b;
    layer0_outputs(1960) <= '1';
    layer0_outputs(1961) <= a and not b;
    layer0_outputs(1962) <= a and not b;
    layer0_outputs(1963) <= '0';
    layer0_outputs(1964) <= not (a or b);
    layer0_outputs(1965) <= a xor b;
    layer0_outputs(1966) <= a or b;
    layer0_outputs(1967) <= a and b;
    layer0_outputs(1968) <= a and b;
    layer0_outputs(1969) <= '0';
    layer0_outputs(1970) <= not a;
    layer0_outputs(1971) <= b and not a;
    layer0_outputs(1972) <= not (a xor b);
    layer0_outputs(1973) <= not b;
    layer0_outputs(1974) <= not (a or b);
    layer0_outputs(1975) <= b;
    layer0_outputs(1976) <= not b;
    layer0_outputs(1977) <= a and b;
    layer0_outputs(1978) <= '1';
    layer0_outputs(1979) <= a and b;
    layer0_outputs(1980) <= '1';
    layer0_outputs(1981) <= not a;
    layer0_outputs(1982) <= not a or b;
    layer0_outputs(1983) <= not a;
    layer0_outputs(1984) <= a;
    layer0_outputs(1985) <= b;
    layer0_outputs(1986) <= b and not a;
    layer0_outputs(1987) <= not (a and b);
    layer0_outputs(1988) <= not (a xor b);
    layer0_outputs(1989) <= not b or a;
    layer0_outputs(1990) <= not b;
    layer0_outputs(1991) <= a;
    layer0_outputs(1992) <= not a or b;
    layer0_outputs(1993) <= not (a xor b);
    layer0_outputs(1994) <= '1';
    layer0_outputs(1995) <= '0';
    layer0_outputs(1996) <= not (a or b);
    layer0_outputs(1997) <= not (a xor b);
    layer0_outputs(1998) <= not (a or b);
    layer0_outputs(1999) <= a;
    layer0_outputs(2000) <= '1';
    layer0_outputs(2001) <= not b or a;
    layer0_outputs(2002) <= not (a xor b);
    layer0_outputs(2003) <= b and not a;
    layer0_outputs(2004) <= '0';
    layer0_outputs(2005) <= not b or a;
    layer0_outputs(2006) <= not a or b;
    layer0_outputs(2007) <= not (a or b);
    layer0_outputs(2008) <= not b;
    layer0_outputs(2009) <= a or b;
    layer0_outputs(2010) <= not b or a;
    layer0_outputs(2011) <= a;
    layer0_outputs(2012) <= not a;
    layer0_outputs(2013) <= not (a xor b);
    layer0_outputs(2014) <= a;
    layer0_outputs(2015) <= not a;
    layer0_outputs(2016) <= a or b;
    layer0_outputs(2017) <= b and not a;
    layer0_outputs(2018) <= b and not a;
    layer0_outputs(2019) <= not b or a;
    layer0_outputs(2020) <= not a or b;
    layer0_outputs(2021) <= a and b;
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= a and not b;
    layer0_outputs(2024) <= '0';
    layer0_outputs(2025) <= b;
    layer0_outputs(2026) <= '1';
    layer0_outputs(2027) <= a and b;
    layer0_outputs(2028) <= a and b;
    layer0_outputs(2029) <= a and b;
    layer0_outputs(2030) <= a xor b;
    layer0_outputs(2031) <= a or b;
    layer0_outputs(2032) <= a;
    layer0_outputs(2033) <= b;
    layer0_outputs(2034) <= not b or a;
    layer0_outputs(2035) <= not (a or b);
    layer0_outputs(2036) <= a;
    layer0_outputs(2037) <= a and b;
    layer0_outputs(2038) <= not b;
    layer0_outputs(2039) <= not a;
    layer0_outputs(2040) <= not (a or b);
    layer0_outputs(2041) <= not b or a;
    layer0_outputs(2042) <= a and b;
    layer0_outputs(2043) <= a or b;
    layer0_outputs(2044) <= not a or b;
    layer0_outputs(2045) <= '1';
    layer0_outputs(2046) <= a or b;
    layer0_outputs(2047) <= '0';
    layer0_outputs(2048) <= a and b;
    layer0_outputs(2049) <= not b or a;
    layer0_outputs(2050) <= a xor b;
    layer0_outputs(2051) <= a and b;
    layer0_outputs(2052) <= a and b;
    layer0_outputs(2053) <= a and b;
    layer0_outputs(2054) <= a or b;
    layer0_outputs(2055) <= a xor b;
    layer0_outputs(2056) <= not (a and b);
    layer0_outputs(2057) <= '0';
    layer0_outputs(2058) <= a and not b;
    layer0_outputs(2059) <= not b;
    layer0_outputs(2060) <= not (a or b);
    layer0_outputs(2061) <= not b or a;
    layer0_outputs(2062) <= not a;
    layer0_outputs(2063) <= not b;
    layer0_outputs(2064) <= a and not b;
    layer0_outputs(2065) <= a xor b;
    layer0_outputs(2066) <= not (a and b);
    layer0_outputs(2067) <= b and not a;
    layer0_outputs(2068) <= not (a and b);
    layer0_outputs(2069) <= not (a or b);
    layer0_outputs(2070) <= a and b;
    layer0_outputs(2071) <= not (a or b);
    layer0_outputs(2072) <= a and b;
    layer0_outputs(2073) <= not (a or b);
    layer0_outputs(2074) <= not (a and b);
    layer0_outputs(2075) <= not b or a;
    layer0_outputs(2076) <= not a;
    layer0_outputs(2077) <= not b;
    layer0_outputs(2078) <= not a or b;
    layer0_outputs(2079) <= '0';
    layer0_outputs(2080) <= a or b;
    layer0_outputs(2081) <= a or b;
    layer0_outputs(2082) <= a and b;
    layer0_outputs(2083) <= b and not a;
    layer0_outputs(2084) <= b and not a;
    layer0_outputs(2085) <= '1';
    layer0_outputs(2086) <= b and not a;
    layer0_outputs(2087) <= not (a and b);
    layer0_outputs(2088) <= b and not a;
    layer0_outputs(2089) <= a or b;
    layer0_outputs(2090) <= not (a xor b);
    layer0_outputs(2091) <= b;
    layer0_outputs(2092) <= not a;
    layer0_outputs(2093) <= not b;
    layer0_outputs(2094) <= b and not a;
    layer0_outputs(2095) <= b and not a;
    layer0_outputs(2096) <= b and not a;
    layer0_outputs(2097) <= a and b;
    layer0_outputs(2098) <= a or b;
    layer0_outputs(2099) <= a or b;
    layer0_outputs(2100) <= a xor b;
    layer0_outputs(2101) <= a and not b;
    layer0_outputs(2102) <= a;
    layer0_outputs(2103) <= a and not b;
    layer0_outputs(2104) <= not a or b;
    layer0_outputs(2105) <= not (a and b);
    layer0_outputs(2106) <= not a;
    layer0_outputs(2107) <= not (a and b);
    layer0_outputs(2108) <= b and not a;
    layer0_outputs(2109) <= not (a and b);
    layer0_outputs(2110) <= not a;
    layer0_outputs(2111) <= not a or b;
    layer0_outputs(2112) <= b;
    layer0_outputs(2113) <= '1';
    layer0_outputs(2114) <= a or b;
    layer0_outputs(2115) <= a xor b;
    layer0_outputs(2116) <= a or b;
    layer0_outputs(2117) <= a and b;
    layer0_outputs(2118) <= not (a xor b);
    layer0_outputs(2119) <= not (a xor b);
    layer0_outputs(2120) <= '1';
    layer0_outputs(2121) <= '0';
    layer0_outputs(2122) <= a and not b;
    layer0_outputs(2123) <= not a or b;
    layer0_outputs(2124) <= not b;
    layer0_outputs(2125) <= not b or a;
    layer0_outputs(2126) <= not b;
    layer0_outputs(2127) <= '1';
    layer0_outputs(2128) <= not (a and b);
    layer0_outputs(2129) <= a or b;
    layer0_outputs(2130) <= a and not b;
    layer0_outputs(2131) <= not (a xor b);
    layer0_outputs(2132) <= b;
    layer0_outputs(2133) <= '1';
    layer0_outputs(2134) <= b;
    layer0_outputs(2135) <= not (a xor b);
    layer0_outputs(2136) <= '1';
    layer0_outputs(2137) <= '0';
    layer0_outputs(2138) <= not (a or b);
    layer0_outputs(2139) <= a xor b;
    layer0_outputs(2140) <= not (a or b);
    layer0_outputs(2141) <= a;
    layer0_outputs(2142) <= not (a xor b);
    layer0_outputs(2143) <= b;
    layer0_outputs(2144) <= a and not b;
    layer0_outputs(2145) <= '0';
    layer0_outputs(2146) <= a or b;
    layer0_outputs(2147) <= not b;
    layer0_outputs(2148) <= b and not a;
    layer0_outputs(2149) <= b;
    layer0_outputs(2150) <= a;
    layer0_outputs(2151) <= not a;
    layer0_outputs(2152) <= '0';
    layer0_outputs(2153) <= not b or a;
    layer0_outputs(2154) <= a or b;
    layer0_outputs(2155) <= a;
    layer0_outputs(2156) <= not (a xor b);
    layer0_outputs(2157) <= a;
    layer0_outputs(2158) <= not a;
    layer0_outputs(2159) <= not (a or b);
    layer0_outputs(2160) <= '0';
    layer0_outputs(2161) <= a or b;
    layer0_outputs(2162) <= not a;
    layer0_outputs(2163) <= a or b;
    layer0_outputs(2164) <= not b;
    layer0_outputs(2165) <= not (a and b);
    layer0_outputs(2166) <= not (a and b);
    layer0_outputs(2167) <= a and not b;
    layer0_outputs(2168) <= not (a xor b);
    layer0_outputs(2169) <= not (a or b);
    layer0_outputs(2170) <= b and not a;
    layer0_outputs(2171) <= b and not a;
    layer0_outputs(2172) <= a and b;
    layer0_outputs(2173) <= a and not b;
    layer0_outputs(2174) <= '1';
    layer0_outputs(2175) <= a and not b;
    layer0_outputs(2176) <= not b or a;
    layer0_outputs(2177) <= not a;
    layer0_outputs(2178) <= not b or a;
    layer0_outputs(2179) <= a;
    layer0_outputs(2180) <= a or b;
    layer0_outputs(2181) <= a and not b;
    layer0_outputs(2182) <= a and not b;
    layer0_outputs(2183) <= a or b;
    layer0_outputs(2184) <= a;
    layer0_outputs(2185) <= not (a or b);
    layer0_outputs(2186) <= not (a and b);
    layer0_outputs(2187) <= not (a xor b);
    layer0_outputs(2188) <= not a;
    layer0_outputs(2189) <= not a or b;
    layer0_outputs(2190) <= not (a xor b);
    layer0_outputs(2191) <= b and not a;
    layer0_outputs(2192) <= not (a or b);
    layer0_outputs(2193) <= '0';
    layer0_outputs(2194) <= not b or a;
    layer0_outputs(2195) <= not a or b;
    layer0_outputs(2196) <= b;
    layer0_outputs(2197) <= not (a xor b);
    layer0_outputs(2198) <= not (a xor b);
    layer0_outputs(2199) <= not (a and b);
    layer0_outputs(2200) <= b;
    layer0_outputs(2201) <= a;
    layer0_outputs(2202) <= '1';
    layer0_outputs(2203) <= a or b;
    layer0_outputs(2204) <= not a or b;
    layer0_outputs(2205) <= not (a xor b);
    layer0_outputs(2206) <= a or b;
    layer0_outputs(2207) <= not (a and b);
    layer0_outputs(2208) <= not (a or b);
    layer0_outputs(2209) <= b;
    layer0_outputs(2210) <= '0';
    layer0_outputs(2211) <= '0';
    layer0_outputs(2212) <= b and not a;
    layer0_outputs(2213) <= not b or a;
    layer0_outputs(2214) <= not a;
    layer0_outputs(2215) <= a;
    layer0_outputs(2216) <= not b or a;
    layer0_outputs(2217) <= not b;
    layer0_outputs(2218) <= '1';
    layer0_outputs(2219) <= a and not b;
    layer0_outputs(2220) <= a and not b;
    layer0_outputs(2221) <= not (a or b);
    layer0_outputs(2222) <= not b or a;
    layer0_outputs(2223) <= not (a and b);
    layer0_outputs(2224) <= '0';
    layer0_outputs(2225) <= not b;
    layer0_outputs(2226) <= not b or a;
    layer0_outputs(2227) <= not a;
    layer0_outputs(2228) <= '1';
    layer0_outputs(2229) <= a or b;
    layer0_outputs(2230) <= a or b;
    layer0_outputs(2231) <= b and not a;
    layer0_outputs(2232) <= not b or a;
    layer0_outputs(2233) <= a xor b;
    layer0_outputs(2234) <= a or b;
    layer0_outputs(2235) <= a and b;
    layer0_outputs(2236) <= not a;
    layer0_outputs(2237) <= not b;
    layer0_outputs(2238) <= not b;
    layer0_outputs(2239) <= a or b;
    layer0_outputs(2240) <= not (a or b);
    layer0_outputs(2241) <= not a;
    layer0_outputs(2242) <= a or b;
    layer0_outputs(2243) <= '0';
    layer0_outputs(2244) <= not b;
    layer0_outputs(2245) <= a xor b;
    layer0_outputs(2246) <= a and not b;
    layer0_outputs(2247) <= not (a or b);
    layer0_outputs(2248) <= not (a and b);
    layer0_outputs(2249) <= not a or b;
    layer0_outputs(2250) <= not a or b;
    layer0_outputs(2251) <= '1';
    layer0_outputs(2252) <= not a;
    layer0_outputs(2253) <= not (a and b);
    layer0_outputs(2254) <= not (a or b);
    layer0_outputs(2255) <= a or b;
    layer0_outputs(2256) <= not (a or b);
    layer0_outputs(2257) <= not a;
    layer0_outputs(2258) <= a and b;
    layer0_outputs(2259) <= not a;
    layer0_outputs(2260) <= not b;
    layer0_outputs(2261) <= not b or a;
    layer0_outputs(2262) <= a;
    layer0_outputs(2263) <= a;
    layer0_outputs(2264) <= '1';
    layer0_outputs(2265) <= b and not a;
    layer0_outputs(2266) <= a and b;
    layer0_outputs(2267) <= a and not b;
    layer0_outputs(2268) <= a;
    layer0_outputs(2269) <= not b or a;
    layer0_outputs(2270) <= a or b;
    layer0_outputs(2271) <= not b or a;
    layer0_outputs(2272) <= not a;
    layer0_outputs(2273) <= a;
    layer0_outputs(2274) <= a and not b;
    layer0_outputs(2275) <= not (a or b);
    layer0_outputs(2276) <= not (a or b);
    layer0_outputs(2277) <= not a;
    layer0_outputs(2278) <= '0';
    layer0_outputs(2279) <= b;
    layer0_outputs(2280) <= a;
    layer0_outputs(2281) <= not a;
    layer0_outputs(2282) <= not (a and b);
    layer0_outputs(2283) <= not (a and b);
    layer0_outputs(2284) <= not b;
    layer0_outputs(2285) <= a or b;
    layer0_outputs(2286) <= not b;
    layer0_outputs(2287) <= not b or a;
    layer0_outputs(2288) <= not b;
    layer0_outputs(2289) <= not (a or b);
    layer0_outputs(2290) <= not b or a;
    layer0_outputs(2291) <= not (a and b);
    layer0_outputs(2292) <= b and not a;
    layer0_outputs(2293) <= b;
    layer0_outputs(2294) <= not (a or b);
    layer0_outputs(2295) <= not a;
    layer0_outputs(2296) <= not b;
    layer0_outputs(2297) <= not a;
    layer0_outputs(2298) <= not (a and b);
    layer0_outputs(2299) <= a or b;
    layer0_outputs(2300) <= not (a and b);
    layer0_outputs(2301) <= not a or b;
    layer0_outputs(2302) <= not a;
    layer0_outputs(2303) <= b;
    layer0_outputs(2304) <= a xor b;
    layer0_outputs(2305) <= not (a xor b);
    layer0_outputs(2306) <= not (a or b);
    layer0_outputs(2307) <= not b or a;
    layer0_outputs(2308) <= not b or a;
    layer0_outputs(2309) <= a and not b;
    layer0_outputs(2310) <= a;
    layer0_outputs(2311) <= '0';
    layer0_outputs(2312) <= not (a xor b);
    layer0_outputs(2313) <= not b;
    layer0_outputs(2314) <= not (a or b);
    layer0_outputs(2315) <= b;
    layer0_outputs(2316) <= not a or b;
    layer0_outputs(2317) <= not (a xor b);
    layer0_outputs(2318) <= not b;
    layer0_outputs(2319) <= not a;
    layer0_outputs(2320) <= not b;
    layer0_outputs(2321) <= a and b;
    layer0_outputs(2322) <= b and not a;
    layer0_outputs(2323) <= not a or b;
    layer0_outputs(2324) <= not (a and b);
    layer0_outputs(2325) <= '1';
    layer0_outputs(2326) <= b;
    layer0_outputs(2327) <= a or b;
    layer0_outputs(2328) <= a or b;
    layer0_outputs(2329) <= not (a or b);
    layer0_outputs(2330) <= a;
    layer0_outputs(2331) <= b;
    layer0_outputs(2332) <= not (a and b);
    layer0_outputs(2333) <= not (a or b);
    layer0_outputs(2334) <= '1';
    layer0_outputs(2335) <= a and not b;
    layer0_outputs(2336) <= a xor b;
    layer0_outputs(2337) <= not (a and b);
    layer0_outputs(2338) <= not b;
    layer0_outputs(2339) <= a or b;
    layer0_outputs(2340) <= not (a xor b);
    layer0_outputs(2341) <= a xor b;
    layer0_outputs(2342) <= not (a xor b);
    layer0_outputs(2343) <= not (a or b);
    layer0_outputs(2344) <= b and not a;
    layer0_outputs(2345) <= '1';
    layer0_outputs(2346) <= not a;
    layer0_outputs(2347) <= b;
    layer0_outputs(2348) <= a and not b;
    layer0_outputs(2349) <= b;
    layer0_outputs(2350) <= not a or b;
    layer0_outputs(2351) <= not b;
    layer0_outputs(2352) <= '1';
    layer0_outputs(2353) <= a and b;
    layer0_outputs(2354) <= b;
    layer0_outputs(2355) <= b and not a;
    layer0_outputs(2356) <= a;
    layer0_outputs(2357) <= '0';
    layer0_outputs(2358) <= '0';
    layer0_outputs(2359) <= b and not a;
    layer0_outputs(2360) <= not a;
    layer0_outputs(2361) <= a;
    layer0_outputs(2362) <= not b;
    layer0_outputs(2363) <= b;
    layer0_outputs(2364) <= not (a or b);
    layer0_outputs(2365) <= a or b;
    layer0_outputs(2366) <= not (a and b);
    layer0_outputs(2367) <= not b;
    layer0_outputs(2368) <= a;
    layer0_outputs(2369) <= '1';
    layer0_outputs(2370) <= b;
    layer0_outputs(2371) <= '1';
    layer0_outputs(2372) <= not b;
    layer0_outputs(2373) <= a xor b;
    layer0_outputs(2374) <= b;
    layer0_outputs(2375) <= not a or b;
    layer0_outputs(2376) <= b and not a;
    layer0_outputs(2377) <= a or b;
    layer0_outputs(2378) <= not (a or b);
    layer0_outputs(2379) <= a or b;
    layer0_outputs(2380) <= not (a and b);
    layer0_outputs(2381) <= not (a xor b);
    layer0_outputs(2382) <= a;
    layer0_outputs(2383) <= b and not a;
    layer0_outputs(2384) <= b;
    layer0_outputs(2385) <= not b;
    layer0_outputs(2386) <= a and not b;
    layer0_outputs(2387) <= '1';
    layer0_outputs(2388) <= not (a or b);
    layer0_outputs(2389) <= not a;
    layer0_outputs(2390) <= a;
    layer0_outputs(2391) <= not (a xor b);
    layer0_outputs(2392) <= a;
    layer0_outputs(2393) <= a and not b;
    layer0_outputs(2394) <= not (a or b);
    layer0_outputs(2395) <= not b or a;
    layer0_outputs(2396) <= '0';
    layer0_outputs(2397) <= a or b;
    layer0_outputs(2398) <= not a;
    layer0_outputs(2399) <= not (a xor b);
    layer0_outputs(2400) <= b;
    layer0_outputs(2401) <= not (a xor b);
    layer0_outputs(2402) <= '1';
    layer0_outputs(2403) <= a;
    layer0_outputs(2404) <= not a;
    layer0_outputs(2405) <= b and not a;
    layer0_outputs(2406) <= not a;
    layer0_outputs(2407) <= b;
    layer0_outputs(2408) <= not (a or b);
    layer0_outputs(2409) <= not a or b;
    layer0_outputs(2410) <= not (a or b);
    layer0_outputs(2411) <= not (a or b);
    layer0_outputs(2412) <= not b or a;
    layer0_outputs(2413) <= not (a and b);
    layer0_outputs(2414) <= not b;
    layer0_outputs(2415) <= not (a xor b);
    layer0_outputs(2416) <= not b or a;
    layer0_outputs(2417) <= not a or b;
    layer0_outputs(2418) <= not (a or b);
    layer0_outputs(2419) <= not (a xor b);
    layer0_outputs(2420) <= a and not b;
    layer0_outputs(2421) <= '0';
    layer0_outputs(2422) <= a or b;
    layer0_outputs(2423) <= not a;
    layer0_outputs(2424) <= b;
    layer0_outputs(2425) <= not a;
    layer0_outputs(2426) <= not (a or b);
    layer0_outputs(2427) <= a xor b;
    layer0_outputs(2428) <= not (a and b);
    layer0_outputs(2429) <= not b;
    layer0_outputs(2430) <= not (a or b);
    layer0_outputs(2431) <= a or b;
    layer0_outputs(2432) <= not (a or b);
    layer0_outputs(2433) <= not b;
    layer0_outputs(2434) <= not a or b;
    layer0_outputs(2435) <= a xor b;
    layer0_outputs(2436) <= not b;
    layer0_outputs(2437) <= a and b;
    layer0_outputs(2438) <= a;
    layer0_outputs(2439) <= not a or b;
    layer0_outputs(2440) <= '0';
    layer0_outputs(2441) <= not (a xor b);
    layer0_outputs(2442) <= '1';
    layer0_outputs(2443) <= a or b;
    layer0_outputs(2444) <= not b;
    layer0_outputs(2445) <= b and not a;
    layer0_outputs(2446) <= '1';
    layer0_outputs(2447) <= not b or a;
    layer0_outputs(2448) <= '1';
    layer0_outputs(2449) <= b and not a;
    layer0_outputs(2450) <= not a;
    layer0_outputs(2451) <= not (a or b);
    layer0_outputs(2452) <= not b or a;
    layer0_outputs(2453) <= not a or b;
    layer0_outputs(2454) <= not b or a;
    layer0_outputs(2455) <= not (a or b);
    layer0_outputs(2456) <= '0';
    layer0_outputs(2457) <= a and not b;
    layer0_outputs(2458) <= a;
    layer0_outputs(2459) <= a or b;
    layer0_outputs(2460) <= a or b;
    layer0_outputs(2461) <= b;
    layer0_outputs(2462) <= b and not a;
    layer0_outputs(2463) <= '0';
    layer0_outputs(2464) <= not (a xor b);
    layer0_outputs(2465) <= not (a xor b);
    layer0_outputs(2466) <= a;
    layer0_outputs(2467) <= b;
    layer0_outputs(2468) <= not b or a;
    layer0_outputs(2469) <= not a or b;
    layer0_outputs(2470) <= not a or b;
    layer0_outputs(2471) <= b and not a;
    layer0_outputs(2472) <= not a or b;
    layer0_outputs(2473) <= a or b;
    layer0_outputs(2474) <= a or b;
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= not b or a;
    layer0_outputs(2477) <= b and not a;
    layer0_outputs(2478) <= a;
    layer0_outputs(2479) <= not a;
    layer0_outputs(2480) <= a;
    layer0_outputs(2481) <= not (a and b);
    layer0_outputs(2482) <= not b;
    layer0_outputs(2483) <= '0';
    layer0_outputs(2484) <= not (a xor b);
    layer0_outputs(2485) <= not a or b;
    layer0_outputs(2486) <= not (a xor b);
    layer0_outputs(2487) <= a and b;
    layer0_outputs(2488) <= not b or a;
    layer0_outputs(2489) <= a xor b;
    layer0_outputs(2490) <= a and not b;
    layer0_outputs(2491) <= '0';
    layer0_outputs(2492) <= b and not a;
    layer0_outputs(2493) <= a or b;
    layer0_outputs(2494) <= a xor b;
    layer0_outputs(2495) <= not b;
    layer0_outputs(2496) <= a xor b;
    layer0_outputs(2497) <= b;
    layer0_outputs(2498) <= a;
    layer0_outputs(2499) <= a;
    layer0_outputs(2500) <= '1';
    layer0_outputs(2501) <= a;
    layer0_outputs(2502) <= not b or a;
    layer0_outputs(2503) <= not a;
    layer0_outputs(2504) <= not b or a;
    layer0_outputs(2505) <= a xor b;
    layer0_outputs(2506) <= not (a and b);
    layer0_outputs(2507) <= not a or b;
    layer0_outputs(2508) <= '0';
    layer0_outputs(2509) <= a xor b;
    layer0_outputs(2510) <= not b or a;
    layer0_outputs(2511) <= not b;
    layer0_outputs(2512) <= a;
    layer0_outputs(2513) <= not (a or b);
    layer0_outputs(2514) <= not (a or b);
    layer0_outputs(2515) <= a and b;
    layer0_outputs(2516) <= a or b;
    layer0_outputs(2517) <= b;
    layer0_outputs(2518) <= '0';
    layer0_outputs(2519) <= not (a or b);
    layer0_outputs(2520) <= not a;
    layer0_outputs(2521) <= a or b;
    layer0_outputs(2522) <= a or b;
    layer0_outputs(2523) <= not a or b;
    layer0_outputs(2524) <= not (a xor b);
    layer0_outputs(2525) <= a;
    layer0_outputs(2526) <= a;
    layer0_outputs(2527) <= a;
    layer0_outputs(2528) <= not a;
    layer0_outputs(2529) <= a and not b;
    layer0_outputs(2530) <= a or b;
    layer0_outputs(2531) <= not (a and b);
    layer0_outputs(2532) <= '1';
    layer0_outputs(2533) <= a or b;
    layer0_outputs(2534) <= not b or a;
    layer0_outputs(2535) <= not a;
    layer0_outputs(2536) <= not a or b;
    layer0_outputs(2537) <= not (a or b);
    layer0_outputs(2538) <= a;
    layer0_outputs(2539) <= not b;
    layer0_outputs(2540) <= '1';
    layer0_outputs(2541) <= a;
    layer0_outputs(2542) <= a or b;
    layer0_outputs(2543) <= not b;
    layer0_outputs(2544) <= not b;
    layer0_outputs(2545) <= not (a or b);
    layer0_outputs(2546) <= not b or a;
    layer0_outputs(2547) <= b and not a;
    layer0_outputs(2548) <= not (a and b);
    layer0_outputs(2549) <= a and not b;
    layer0_outputs(2550) <= b;
    layer0_outputs(2551) <= not a;
    layer0_outputs(2552) <= a or b;
    layer0_outputs(2553) <= a;
    layer0_outputs(2554) <= '1';
    layer0_outputs(2555) <= a;
    layer0_outputs(2556) <= not a or b;
    layer0_outputs(2557) <= a;
    layer0_outputs(2558) <= '0';
    layer0_outputs(2559) <= not (a and b);
    layer0_outputs(2560) <= a or b;
    layer0_outputs(2561) <= a;
    layer0_outputs(2562) <= '0';
    layer0_outputs(2563) <= a and b;
    layer0_outputs(2564) <= a xor b;
    layer0_outputs(2565) <= not (a or b);
    layer0_outputs(2566) <= not b;
    layer0_outputs(2567) <= a;
    layer0_outputs(2568) <= not a or b;
    layer0_outputs(2569) <= a;
    layer0_outputs(2570) <= b;
    layer0_outputs(2571) <= '1';
    layer0_outputs(2572) <= not (a xor b);
    layer0_outputs(2573) <= a;
    layer0_outputs(2574) <= not (a and b);
    layer0_outputs(2575) <= a;
    layer0_outputs(2576) <= b;
    layer0_outputs(2577) <= not b or a;
    layer0_outputs(2578) <= not a;
    layer0_outputs(2579) <= b;
    layer0_outputs(2580) <= a;
    layer0_outputs(2581) <= a and not b;
    layer0_outputs(2582) <= '0';
    layer0_outputs(2583) <= '0';
    layer0_outputs(2584) <= not b;
    layer0_outputs(2585) <= '1';
    layer0_outputs(2586) <= a or b;
    layer0_outputs(2587) <= not (a and b);
    layer0_outputs(2588) <= a and b;
    layer0_outputs(2589) <= not (a and b);
    layer0_outputs(2590) <= not a;
    layer0_outputs(2591) <= '1';
    layer0_outputs(2592) <= not (a and b);
    layer0_outputs(2593) <= a and b;
    layer0_outputs(2594) <= a or b;
    layer0_outputs(2595) <= a and b;
    layer0_outputs(2596) <= not b or a;
    layer0_outputs(2597) <= not a or b;
    layer0_outputs(2598) <= '0';
    layer0_outputs(2599) <= b and not a;
    layer0_outputs(2600) <= not (a or b);
    layer0_outputs(2601) <= a or b;
    layer0_outputs(2602) <= not a or b;
    layer0_outputs(2603) <= '0';
    layer0_outputs(2604) <= '0';
    layer0_outputs(2605) <= '1';
    layer0_outputs(2606) <= not a or b;
    layer0_outputs(2607) <= b;
    layer0_outputs(2608) <= '1';
    layer0_outputs(2609) <= not a or b;
    layer0_outputs(2610) <= '0';
    layer0_outputs(2611) <= b and not a;
    layer0_outputs(2612) <= not (a or b);
    layer0_outputs(2613) <= not b or a;
    layer0_outputs(2614) <= '1';
    layer0_outputs(2615) <= b and not a;
    layer0_outputs(2616) <= not b or a;
    layer0_outputs(2617) <= not a or b;
    layer0_outputs(2618) <= a xor b;
    layer0_outputs(2619) <= a and b;
    layer0_outputs(2620) <= not (a and b);
    layer0_outputs(2621) <= '1';
    layer0_outputs(2622) <= not a;
    layer0_outputs(2623) <= a or b;
    layer0_outputs(2624) <= not (a and b);
    layer0_outputs(2625) <= a;
    layer0_outputs(2626) <= a and not b;
    layer0_outputs(2627) <= a and not b;
    layer0_outputs(2628) <= a or b;
    layer0_outputs(2629) <= not a;
    layer0_outputs(2630) <= not a;
    layer0_outputs(2631) <= not (a or b);
    layer0_outputs(2632) <= not b;
    layer0_outputs(2633) <= a and not b;
    layer0_outputs(2634) <= not (a and b);
    layer0_outputs(2635) <= '1';
    layer0_outputs(2636) <= not (a xor b);
    layer0_outputs(2637) <= a and not b;
    layer0_outputs(2638) <= a xor b;
    layer0_outputs(2639) <= a and b;
    layer0_outputs(2640) <= b and not a;
    layer0_outputs(2641) <= b;
    layer0_outputs(2642) <= not b;
    layer0_outputs(2643) <= not (a xor b);
    layer0_outputs(2644) <= a;
    layer0_outputs(2645) <= b;
    layer0_outputs(2646) <= b and not a;
    layer0_outputs(2647) <= not b;
    layer0_outputs(2648) <= a and b;
    layer0_outputs(2649) <= not b or a;
    layer0_outputs(2650) <= not a or b;
    layer0_outputs(2651) <= not b;
    layer0_outputs(2652) <= not a;
    layer0_outputs(2653) <= a;
    layer0_outputs(2654) <= a and not b;
    layer0_outputs(2655) <= a;
    layer0_outputs(2656) <= not b;
    layer0_outputs(2657) <= b;
    layer0_outputs(2658) <= a and not b;
    layer0_outputs(2659) <= not (a or b);
    layer0_outputs(2660) <= a xor b;
    layer0_outputs(2661) <= b and not a;
    layer0_outputs(2662) <= not (a and b);
    layer0_outputs(2663) <= '0';
    layer0_outputs(2664) <= not a;
    layer0_outputs(2665) <= a and b;
    layer0_outputs(2666) <= a and b;
    layer0_outputs(2667) <= b;
    layer0_outputs(2668) <= '1';
    layer0_outputs(2669) <= a and b;
    layer0_outputs(2670) <= a and not b;
    layer0_outputs(2671) <= not b or a;
    layer0_outputs(2672) <= not (a and b);
    layer0_outputs(2673) <= not a;
    layer0_outputs(2674) <= a or b;
    layer0_outputs(2675) <= a xor b;
    layer0_outputs(2676) <= b and not a;
    layer0_outputs(2677) <= not a;
    layer0_outputs(2678) <= a;
    layer0_outputs(2679) <= '0';
    layer0_outputs(2680) <= not (a and b);
    layer0_outputs(2681) <= not (a and b);
    layer0_outputs(2682) <= '0';
    layer0_outputs(2683) <= a xor b;
    layer0_outputs(2684) <= '1';
    layer0_outputs(2685) <= '1';
    layer0_outputs(2686) <= a;
    layer0_outputs(2687) <= a;
    layer0_outputs(2688) <= a and not b;
    layer0_outputs(2689) <= a or b;
    layer0_outputs(2690) <= a;
    layer0_outputs(2691) <= a;
    layer0_outputs(2692) <= a and not b;
    layer0_outputs(2693) <= a or b;
    layer0_outputs(2694) <= a and not b;
    layer0_outputs(2695) <= a and b;
    layer0_outputs(2696) <= a;
    layer0_outputs(2697) <= not b or a;
    layer0_outputs(2698) <= not a;
    layer0_outputs(2699) <= not b or a;
    layer0_outputs(2700) <= a xor b;
    layer0_outputs(2701) <= not (a or b);
    layer0_outputs(2702) <= not (a or b);
    layer0_outputs(2703) <= '0';
    layer0_outputs(2704) <= not b;
    layer0_outputs(2705) <= '0';
    layer0_outputs(2706) <= a or b;
    layer0_outputs(2707) <= not a;
    layer0_outputs(2708) <= '0';
    layer0_outputs(2709) <= not (a xor b);
    layer0_outputs(2710) <= b and not a;
    layer0_outputs(2711) <= not a or b;
    layer0_outputs(2712) <= '1';
    layer0_outputs(2713) <= not b or a;
    layer0_outputs(2714) <= a or b;
    layer0_outputs(2715) <= a xor b;
    layer0_outputs(2716) <= a or b;
    layer0_outputs(2717) <= not (a and b);
    layer0_outputs(2718) <= a;
    layer0_outputs(2719) <= b;
    layer0_outputs(2720) <= a and b;
    layer0_outputs(2721) <= not a;
    layer0_outputs(2722) <= not b;
    layer0_outputs(2723) <= a and b;
    layer0_outputs(2724) <= a or b;
    layer0_outputs(2725) <= a xor b;
    layer0_outputs(2726) <= not a;
    layer0_outputs(2727) <= '0';
    layer0_outputs(2728) <= not (a or b);
    layer0_outputs(2729) <= not b;
    layer0_outputs(2730) <= not (a or b);
    layer0_outputs(2731) <= a;
    layer0_outputs(2732) <= not a;
    layer0_outputs(2733) <= not a or b;
    layer0_outputs(2734) <= not b;
    layer0_outputs(2735) <= a;
    layer0_outputs(2736) <= '1';
    layer0_outputs(2737) <= a or b;
    layer0_outputs(2738) <= a;
    layer0_outputs(2739) <= not (a and b);
    layer0_outputs(2740) <= a and not b;
    layer0_outputs(2741) <= b and not a;
    layer0_outputs(2742) <= a and not b;
    layer0_outputs(2743) <= a and not b;
    layer0_outputs(2744) <= not (a xor b);
    layer0_outputs(2745) <= a xor b;
    layer0_outputs(2746) <= a or b;
    layer0_outputs(2747) <= b;
    layer0_outputs(2748) <= b;
    layer0_outputs(2749) <= not (a xor b);
    layer0_outputs(2750) <= not b or a;
    layer0_outputs(2751) <= a;
    layer0_outputs(2752) <= not (a and b);
    layer0_outputs(2753) <= not a or b;
    layer0_outputs(2754) <= not (a xor b);
    layer0_outputs(2755) <= not a;
    layer0_outputs(2756) <= not (a and b);
    layer0_outputs(2757) <= b and not a;
    layer0_outputs(2758) <= not (a and b);
    layer0_outputs(2759) <= b;
    layer0_outputs(2760) <= '1';
    layer0_outputs(2761) <= a and b;
    layer0_outputs(2762) <= a and not b;
    layer0_outputs(2763) <= b and not a;
    layer0_outputs(2764) <= not (a and b);
    layer0_outputs(2765) <= a;
    layer0_outputs(2766) <= a;
    layer0_outputs(2767) <= b and not a;
    layer0_outputs(2768) <= not (a and b);
    layer0_outputs(2769) <= a or b;
    layer0_outputs(2770) <= b and not a;
    layer0_outputs(2771) <= not (a or b);
    layer0_outputs(2772) <= not a;
    layer0_outputs(2773) <= '0';
    layer0_outputs(2774) <= not (a and b);
    layer0_outputs(2775) <= a and not b;
    layer0_outputs(2776) <= a or b;
    layer0_outputs(2777) <= a and b;
    layer0_outputs(2778) <= '0';
    layer0_outputs(2779) <= not (a xor b);
    layer0_outputs(2780) <= a or b;
    layer0_outputs(2781) <= not (a and b);
    layer0_outputs(2782) <= a;
    layer0_outputs(2783) <= a xor b;
    layer0_outputs(2784) <= not b or a;
    layer0_outputs(2785) <= not (a and b);
    layer0_outputs(2786) <= not (a or b);
    layer0_outputs(2787) <= b;
    layer0_outputs(2788) <= a;
    layer0_outputs(2789) <= '0';
    layer0_outputs(2790) <= not a or b;
    layer0_outputs(2791) <= not a;
    layer0_outputs(2792) <= a or b;
    layer0_outputs(2793) <= '1';
    layer0_outputs(2794) <= b;
    layer0_outputs(2795) <= a or b;
    layer0_outputs(2796) <= not (a xor b);
    layer0_outputs(2797) <= '0';
    layer0_outputs(2798) <= a or b;
    layer0_outputs(2799) <= not (a xor b);
    layer0_outputs(2800) <= not (a and b);
    layer0_outputs(2801) <= '0';
    layer0_outputs(2802) <= not (a or b);
    layer0_outputs(2803) <= a and b;
    layer0_outputs(2804) <= not (a and b);
    layer0_outputs(2805) <= '0';
    layer0_outputs(2806) <= a and not b;
    layer0_outputs(2807) <= a xor b;
    layer0_outputs(2808) <= not b;
    layer0_outputs(2809) <= not (a and b);
    layer0_outputs(2810) <= '1';
    layer0_outputs(2811) <= b and not a;
    layer0_outputs(2812) <= a or b;
    layer0_outputs(2813) <= '0';
    layer0_outputs(2814) <= not (a and b);
    layer0_outputs(2815) <= not (a or b);
    layer0_outputs(2816) <= a and not b;
    layer0_outputs(2817) <= not (a or b);
    layer0_outputs(2818) <= a and b;
    layer0_outputs(2819) <= not (a or b);
    layer0_outputs(2820) <= b and not a;
    layer0_outputs(2821) <= not b or a;
    layer0_outputs(2822) <= '0';
    layer0_outputs(2823) <= a;
    layer0_outputs(2824) <= not (a and b);
    layer0_outputs(2825) <= b;
    layer0_outputs(2826) <= not (a or b);
    layer0_outputs(2827) <= b;
    layer0_outputs(2828) <= not (a xor b);
    layer0_outputs(2829) <= b and not a;
    layer0_outputs(2830) <= a;
    layer0_outputs(2831) <= a xor b;
    layer0_outputs(2832) <= a xor b;
    layer0_outputs(2833) <= a;
    layer0_outputs(2834) <= a and not b;
    layer0_outputs(2835) <= '0';
    layer0_outputs(2836) <= '0';
    layer0_outputs(2837) <= '0';
    layer0_outputs(2838) <= not a;
    layer0_outputs(2839) <= a;
    layer0_outputs(2840) <= a and b;
    layer0_outputs(2841) <= b;
    layer0_outputs(2842) <= a or b;
    layer0_outputs(2843) <= not b;
    layer0_outputs(2844) <= a and not b;
    layer0_outputs(2845) <= not b or a;
    layer0_outputs(2846) <= b and not a;
    layer0_outputs(2847) <= b;
    layer0_outputs(2848) <= b;
    layer0_outputs(2849) <= a;
    layer0_outputs(2850) <= not (a xor b);
    layer0_outputs(2851) <= not (a xor b);
    layer0_outputs(2852) <= b;
    layer0_outputs(2853) <= not b;
    layer0_outputs(2854) <= '1';
    layer0_outputs(2855) <= a;
    layer0_outputs(2856) <= not b or a;
    layer0_outputs(2857) <= '1';
    layer0_outputs(2858) <= a and not b;
    layer0_outputs(2859) <= a and not b;
    layer0_outputs(2860) <= not a or b;
    layer0_outputs(2861) <= not (a xor b);
    layer0_outputs(2862) <= b and not a;
    layer0_outputs(2863) <= '1';
    layer0_outputs(2864) <= not (a or b);
    layer0_outputs(2865) <= a or b;
    layer0_outputs(2866) <= not (a xor b);
    layer0_outputs(2867) <= '1';
    layer0_outputs(2868) <= not b;
    layer0_outputs(2869) <= not (a and b);
    layer0_outputs(2870) <= a xor b;
    layer0_outputs(2871) <= not b or a;
    layer0_outputs(2872) <= not a or b;
    layer0_outputs(2873) <= a and b;
    layer0_outputs(2874) <= not (a and b);
    layer0_outputs(2875) <= a or b;
    layer0_outputs(2876) <= not a;
    layer0_outputs(2877) <= b;
    layer0_outputs(2878) <= not b or a;
    layer0_outputs(2879) <= not a;
    layer0_outputs(2880) <= not b or a;
    layer0_outputs(2881) <= a;
    layer0_outputs(2882) <= not (a or b);
    layer0_outputs(2883) <= b;
    layer0_outputs(2884) <= b and not a;
    layer0_outputs(2885) <= not (a and b);
    layer0_outputs(2886) <= a;
    layer0_outputs(2887) <= a or b;
    layer0_outputs(2888) <= not a;
    layer0_outputs(2889) <= b and not a;
    layer0_outputs(2890) <= not b;
    layer0_outputs(2891) <= not b or a;
    layer0_outputs(2892) <= b and not a;
    layer0_outputs(2893) <= not b;
    layer0_outputs(2894) <= not a or b;
    layer0_outputs(2895) <= a xor b;
    layer0_outputs(2896) <= not (a or b);
    layer0_outputs(2897) <= a;
    layer0_outputs(2898) <= a or b;
    layer0_outputs(2899) <= not a or b;
    layer0_outputs(2900) <= not b;
    layer0_outputs(2901) <= a xor b;
    layer0_outputs(2902) <= b and not a;
    layer0_outputs(2903) <= b;
    layer0_outputs(2904) <= not b or a;
    layer0_outputs(2905) <= not a;
    layer0_outputs(2906) <= a or b;
    layer0_outputs(2907) <= b;
    layer0_outputs(2908) <= not b or a;
    layer0_outputs(2909) <= b;
    layer0_outputs(2910) <= not b;
    layer0_outputs(2911) <= '1';
    layer0_outputs(2912) <= not (a or b);
    layer0_outputs(2913) <= b;
    layer0_outputs(2914) <= not (a and b);
    layer0_outputs(2915) <= a and b;
    layer0_outputs(2916) <= not a or b;
    layer0_outputs(2917) <= not a;
    layer0_outputs(2918) <= a or b;
    layer0_outputs(2919) <= b;
    layer0_outputs(2920) <= a or b;
    layer0_outputs(2921) <= not b;
    layer0_outputs(2922) <= '1';
    layer0_outputs(2923) <= not a;
    layer0_outputs(2924) <= a or b;
    layer0_outputs(2925) <= '0';
    layer0_outputs(2926) <= b;
    layer0_outputs(2927) <= a or b;
    layer0_outputs(2928) <= not b;
    layer0_outputs(2929) <= not a or b;
    layer0_outputs(2930) <= a or b;
    layer0_outputs(2931) <= a and b;
    layer0_outputs(2932) <= b;
    layer0_outputs(2933) <= a xor b;
    layer0_outputs(2934) <= a or b;
    layer0_outputs(2935) <= not b;
    layer0_outputs(2936) <= b;
    layer0_outputs(2937) <= not b;
    layer0_outputs(2938) <= b;
    layer0_outputs(2939) <= not (a or b);
    layer0_outputs(2940) <= b and not a;
    layer0_outputs(2941) <= b;
    layer0_outputs(2942) <= '0';
    layer0_outputs(2943) <= b;
    layer0_outputs(2944) <= not a or b;
    layer0_outputs(2945) <= a;
    layer0_outputs(2946) <= b and not a;
    layer0_outputs(2947) <= not a or b;
    layer0_outputs(2948) <= not (a or b);
    layer0_outputs(2949) <= not (a and b);
    layer0_outputs(2950) <= a xor b;
    layer0_outputs(2951) <= a;
    layer0_outputs(2952) <= not a or b;
    layer0_outputs(2953) <= a and not b;
    layer0_outputs(2954) <= not a;
    layer0_outputs(2955) <= '0';
    layer0_outputs(2956) <= '0';
    layer0_outputs(2957) <= b;
    layer0_outputs(2958) <= '1';
    layer0_outputs(2959) <= '1';
    layer0_outputs(2960) <= not (a and b);
    layer0_outputs(2961) <= not b or a;
    layer0_outputs(2962) <= not (a xor b);
    layer0_outputs(2963) <= not b or a;
    layer0_outputs(2964) <= a;
    layer0_outputs(2965) <= not b;
    layer0_outputs(2966) <= not b;
    layer0_outputs(2967) <= a and not b;
    layer0_outputs(2968) <= a;
    layer0_outputs(2969) <= '1';
    layer0_outputs(2970) <= not a or b;
    layer0_outputs(2971) <= a;
    layer0_outputs(2972) <= a;
    layer0_outputs(2973) <= not (a xor b);
    layer0_outputs(2974) <= not (a or b);
    layer0_outputs(2975) <= not b;
    layer0_outputs(2976) <= '0';
    layer0_outputs(2977) <= b;
    layer0_outputs(2978) <= not (a xor b);
    layer0_outputs(2979) <= b;
    layer0_outputs(2980) <= a and b;
    layer0_outputs(2981) <= a and b;
    layer0_outputs(2982) <= a or b;
    layer0_outputs(2983) <= a;
    layer0_outputs(2984) <= '0';
    layer0_outputs(2985) <= b and not a;
    layer0_outputs(2986) <= not (a xor b);
    layer0_outputs(2987) <= not (a or b);
    layer0_outputs(2988) <= not (a xor b);
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= a;
    layer0_outputs(2991) <= b;
    layer0_outputs(2992) <= not a or b;
    layer0_outputs(2993) <= a and not b;
    layer0_outputs(2994) <= '1';
    layer0_outputs(2995) <= b;
    layer0_outputs(2996) <= not b;
    layer0_outputs(2997) <= a;
    layer0_outputs(2998) <= not (a and b);
    layer0_outputs(2999) <= '1';
    layer0_outputs(3000) <= not b;
    layer0_outputs(3001) <= a xor b;
    layer0_outputs(3002) <= a xor b;
    layer0_outputs(3003) <= a xor b;
    layer0_outputs(3004) <= not b or a;
    layer0_outputs(3005) <= not (a or b);
    layer0_outputs(3006) <= b;
    layer0_outputs(3007) <= a and b;
    layer0_outputs(3008) <= '1';
    layer0_outputs(3009) <= a and not b;
    layer0_outputs(3010) <= not b;
    layer0_outputs(3011) <= not b;
    layer0_outputs(3012) <= not a;
    layer0_outputs(3013) <= a and not b;
    layer0_outputs(3014) <= not b or a;
    layer0_outputs(3015) <= a or b;
    layer0_outputs(3016) <= '0';
    layer0_outputs(3017) <= not b or a;
    layer0_outputs(3018) <= not (a and b);
    layer0_outputs(3019) <= not a;
    layer0_outputs(3020) <= b;
    layer0_outputs(3021) <= '0';
    layer0_outputs(3022) <= '0';
    layer0_outputs(3023) <= not (a xor b);
    layer0_outputs(3024) <= a;
    layer0_outputs(3025) <= a and not b;
    layer0_outputs(3026) <= a or b;
    layer0_outputs(3027) <= not b or a;
    layer0_outputs(3028) <= b and not a;
    layer0_outputs(3029) <= '1';
    layer0_outputs(3030) <= not (a and b);
    layer0_outputs(3031) <= a and b;
    layer0_outputs(3032) <= a;
    layer0_outputs(3033) <= a xor b;
    layer0_outputs(3034) <= not (a xor b);
    layer0_outputs(3035) <= a xor b;
    layer0_outputs(3036) <= not a;
    layer0_outputs(3037) <= not a;
    layer0_outputs(3038) <= '0';
    layer0_outputs(3039) <= not b or a;
    layer0_outputs(3040) <= not a or b;
    layer0_outputs(3041) <= not (a or b);
    layer0_outputs(3042) <= a or b;
    layer0_outputs(3043) <= a and b;
    layer0_outputs(3044) <= a xor b;
    layer0_outputs(3045) <= a or b;
    layer0_outputs(3046) <= not b;
    layer0_outputs(3047) <= a or b;
    layer0_outputs(3048) <= '0';
    layer0_outputs(3049) <= b and not a;
    layer0_outputs(3050) <= a and b;
    layer0_outputs(3051) <= not a;
    layer0_outputs(3052) <= a and not b;
    layer0_outputs(3053) <= a;
    layer0_outputs(3054) <= a or b;
    layer0_outputs(3055) <= '1';
    layer0_outputs(3056) <= not a or b;
    layer0_outputs(3057) <= not b;
    layer0_outputs(3058) <= not (a and b);
    layer0_outputs(3059) <= a and b;
    layer0_outputs(3060) <= not b;
    layer0_outputs(3061) <= a and b;
    layer0_outputs(3062) <= a and not b;
    layer0_outputs(3063) <= '1';
    layer0_outputs(3064) <= a xor b;
    layer0_outputs(3065) <= a and not b;
    layer0_outputs(3066) <= b and not a;
    layer0_outputs(3067) <= not a;
    layer0_outputs(3068) <= not (a and b);
    layer0_outputs(3069) <= b;
    layer0_outputs(3070) <= not a or b;
    layer0_outputs(3071) <= b;
    layer0_outputs(3072) <= '1';
    layer0_outputs(3073) <= a xor b;
    layer0_outputs(3074) <= not (a and b);
    layer0_outputs(3075) <= a and b;
    layer0_outputs(3076) <= a and not b;
    layer0_outputs(3077) <= b;
    layer0_outputs(3078) <= not b;
    layer0_outputs(3079) <= not b;
    layer0_outputs(3080) <= '0';
    layer0_outputs(3081) <= b and not a;
    layer0_outputs(3082) <= not (a or b);
    layer0_outputs(3083) <= not a;
    layer0_outputs(3084) <= not a;
    layer0_outputs(3085) <= '0';
    layer0_outputs(3086) <= not b;
    layer0_outputs(3087) <= '1';
    layer0_outputs(3088) <= not a;
    layer0_outputs(3089) <= '1';
    layer0_outputs(3090) <= b;
    layer0_outputs(3091) <= not (a and b);
    layer0_outputs(3092) <= not (a or b);
    layer0_outputs(3093) <= '0';
    layer0_outputs(3094) <= not (a and b);
    layer0_outputs(3095) <= a or b;
    layer0_outputs(3096) <= not b;
    layer0_outputs(3097) <= not a or b;
    layer0_outputs(3098) <= not (a or b);
    layer0_outputs(3099) <= a xor b;
    layer0_outputs(3100) <= a;
    layer0_outputs(3101) <= a and not b;
    layer0_outputs(3102) <= not (a or b);
    layer0_outputs(3103) <= a and b;
    layer0_outputs(3104) <= a or b;
    layer0_outputs(3105) <= not a;
    layer0_outputs(3106) <= '0';
    layer0_outputs(3107) <= not (a or b);
    layer0_outputs(3108) <= not b or a;
    layer0_outputs(3109) <= b;
    layer0_outputs(3110) <= a and b;
    layer0_outputs(3111) <= not a;
    layer0_outputs(3112) <= not b;
    layer0_outputs(3113) <= a and b;
    layer0_outputs(3114) <= not a or b;
    layer0_outputs(3115) <= a and b;
    layer0_outputs(3116) <= not b or a;
    layer0_outputs(3117) <= '0';
    layer0_outputs(3118) <= not (a or b);
    layer0_outputs(3119) <= a or b;
    layer0_outputs(3120) <= not a;
    layer0_outputs(3121) <= a;
    layer0_outputs(3122) <= '1';
    layer0_outputs(3123) <= '1';
    layer0_outputs(3124) <= not b;
    layer0_outputs(3125) <= a;
    layer0_outputs(3126) <= a and b;
    layer0_outputs(3127) <= b and not a;
    layer0_outputs(3128) <= a and not b;
    layer0_outputs(3129) <= a and not b;
    layer0_outputs(3130) <= a xor b;
    layer0_outputs(3131) <= a xor b;
    layer0_outputs(3132) <= not a;
    layer0_outputs(3133) <= not b;
    layer0_outputs(3134) <= not b or a;
    layer0_outputs(3135) <= a and b;
    layer0_outputs(3136) <= not (a and b);
    layer0_outputs(3137) <= not (a xor b);
    layer0_outputs(3138) <= a;
    layer0_outputs(3139) <= a xor b;
    layer0_outputs(3140) <= '0';
    layer0_outputs(3141) <= not a;
    layer0_outputs(3142) <= '1';
    layer0_outputs(3143) <= a;
    layer0_outputs(3144) <= not (a and b);
    layer0_outputs(3145) <= '1';
    layer0_outputs(3146) <= '1';
    layer0_outputs(3147) <= '1';
    layer0_outputs(3148) <= a and b;
    layer0_outputs(3149) <= a and b;
    layer0_outputs(3150) <= a xor b;
    layer0_outputs(3151) <= not (a xor b);
    layer0_outputs(3152) <= a xor b;
    layer0_outputs(3153) <= a;
    layer0_outputs(3154) <= b;
    layer0_outputs(3155) <= not (a or b);
    layer0_outputs(3156) <= not a;
    layer0_outputs(3157) <= not b or a;
    layer0_outputs(3158) <= '0';
    layer0_outputs(3159) <= not b;
    layer0_outputs(3160) <= not (a and b);
    layer0_outputs(3161) <= not (a xor b);
    layer0_outputs(3162) <= a xor b;
    layer0_outputs(3163) <= '1';
    layer0_outputs(3164) <= not a;
    layer0_outputs(3165) <= '0';
    layer0_outputs(3166) <= a or b;
    layer0_outputs(3167) <= not a;
    layer0_outputs(3168) <= '1';
    layer0_outputs(3169) <= a and b;
    layer0_outputs(3170) <= a and not b;
    layer0_outputs(3171) <= a;
    layer0_outputs(3172) <= a and not b;
    layer0_outputs(3173) <= not (a and b);
    layer0_outputs(3174) <= not b or a;
    layer0_outputs(3175) <= not (a and b);
    layer0_outputs(3176) <= not (a and b);
    layer0_outputs(3177) <= not a or b;
    layer0_outputs(3178) <= not (a and b);
    layer0_outputs(3179) <= a;
    layer0_outputs(3180) <= a;
    layer0_outputs(3181) <= a and not b;
    layer0_outputs(3182) <= not a;
    layer0_outputs(3183) <= not b;
    layer0_outputs(3184) <= b;
    layer0_outputs(3185) <= a or b;
    layer0_outputs(3186) <= a;
    layer0_outputs(3187) <= not (a or b);
    layer0_outputs(3188) <= not b;
    layer0_outputs(3189) <= not b or a;
    layer0_outputs(3190) <= not b or a;
    layer0_outputs(3191) <= not (a or b);
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= not b;
    layer0_outputs(3194) <= '0';
    layer0_outputs(3195) <= a;
    layer0_outputs(3196) <= not (a xor b);
    layer0_outputs(3197) <= not (a or b);
    layer0_outputs(3198) <= a and b;
    layer0_outputs(3199) <= not (a or b);
    layer0_outputs(3200) <= a;
    layer0_outputs(3201) <= '0';
    layer0_outputs(3202) <= not a;
    layer0_outputs(3203) <= b and not a;
    layer0_outputs(3204) <= a xor b;
    layer0_outputs(3205) <= not (a xor b);
    layer0_outputs(3206) <= not b;
    layer0_outputs(3207) <= not (a or b);
    layer0_outputs(3208) <= not (a or b);
    layer0_outputs(3209) <= not (a or b);
    layer0_outputs(3210) <= not b;
    layer0_outputs(3211) <= not a or b;
    layer0_outputs(3212) <= '0';
    layer0_outputs(3213) <= not b;
    layer0_outputs(3214) <= b;
    layer0_outputs(3215) <= not (a or b);
    layer0_outputs(3216) <= not b or a;
    layer0_outputs(3217) <= not a;
    layer0_outputs(3218) <= a or b;
    layer0_outputs(3219) <= a;
    layer0_outputs(3220) <= '1';
    layer0_outputs(3221) <= '0';
    layer0_outputs(3222) <= not (a or b);
    layer0_outputs(3223) <= not b or a;
    layer0_outputs(3224) <= a;
    layer0_outputs(3225) <= not (a or b);
    layer0_outputs(3226) <= not a;
    layer0_outputs(3227) <= not b;
    layer0_outputs(3228) <= not b or a;
    layer0_outputs(3229) <= not (a xor b);
    layer0_outputs(3230) <= not (a or b);
    layer0_outputs(3231) <= not (a or b);
    layer0_outputs(3232) <= not a or b;
    layer0_outputs(3233) <= a and b;
    layer0_outputs(3234) <= '1';
    layer0_outputs(3235) <= b and not a;
    layer0_outputs(3236) <= b and not a;
    layer0_outputs(3237) <= '1';
    layer0_outputs(3238) <= a and not b;
    layer0_outputs(3239) <= a;
    layer0_outputs(3240) <= '0';
    layer0_outputs(3241) <= not (a xor b);
    layer0_outputs(3242) <= not (a and b);
    layer0_outputs(3243) <= not (a and b);
    layer0_outputs(3244) <= a or b;
    layer0_outputs(3245) <= a;
    layer0_outputs(3246) <= a;
    layer0_outputs(3247) <= a;
    layer0_outputs(3248) <= '0';
    layer0_outputs(3249) <= not a;
    layer0_outputs(3250) <= a or b;
    layer0_outputs(3251) <= not (a xor b);
    layer0_outputs(3252) <= not (a xor b);
    layer0_outputs(3253) <= a or b;
    layer0_outputs(3254) <= not b or a;
    layer0_outputs(3255) <= a or b;
    layer0_outputs(3256) <= a xor b;
    layer0_outputs(3257) <= a xor b;
    layer0_outputs(3258) <= a and not b;
    layer0_outputs(3259) <= '1';
    layer0_outputs(3260) <= not a or b;
    layer0_outputs(3261) <= a or b;
    layer0_outputs(3262) <= b and not a;
    layer0_outputs(3263) <= b and not a;
    layer0_outputs(3264) <= a or b;
    layer0_outputs(3265) <= a and b;
    layer0_outputs(3266) <= not (a and b);
    layer0_outputs(3267) <= a;
    layer0_outputs(3268) <= not a;
    layer0_outputs(3269) <= b;
    layer0_outputs(3270) <= a and b;
    layer0_outputs(3271) <= not (a or b);
    layer0_outputs(3272) <= a;
    layer0_outputs(3273) <= a or b;
    layer0_outputs(3274) <= a and b;
    layer0_outputs(3275) <= not (a xor b);
    layer0_outputs(3276) <= not b or a;
    layer0_outputs(3277) <= a and b;
    layer0_outputs(3278) <= not a or b;
    layer0_outputs(3279) <= a and b;
    layer0_outputs(3280) <= not a;
    layer0_outputs(3281) <= not (a and b);
    layer0_outputs(3282) <= a or b;
    layer0_outputs(3283) <= '0';
    layer0_outputs(3284) <= b and not a;
    layer0_outputs(3285) <= '1';
    layer0_outputs(3286) <= not b or a;
    layer0_outputs(3287) <= a or b;
    layer0_outputs(3288) <= '1';
    layer0_outputs(3289) <= a and b;
    layer0_outputs(3290) <= '1';
    layer0_outputs(3291) <= '1';
    layer0_outputs(3292) <= a or b;
    layer0_outputs(3293) <= not (a xor b);
    layer0_outputs(3294) <= not a or b;
    layer0_outputs(3295) <= '1';
    layer0_outputs(3296) <= b;
    layer0_outputs(3297) <= not b;
    layer0_outputs(3298) <= '1';
    layer0_outputs(3299) <= not a or b;
    layer0_outputs(3300) <= not a or b;
    layer0_outputs(3301) <= a;
    layer0_outputs(3302) <= a and b;
    layer0_outputs(3303) <= '1';
    layer0_outputs(3304) <= '1';
    layer0_outputs(3305) <= not b;
    layer0_outputs(3306) <= not b;
    layer0_outputs(3307) <= '0';
    layer0_outputs(3308) <= not (a or b);
    layer0_outputs(3309) <= a and b;
    layer0_outputs(3310) <= '0';
    layer0_outputs(3311) <= '1';
    layer0_outputs(3312) <= '0';
    layer0_outputs(3313) <= not (a or b);
    layer0_outputs(3314) <= not (a xor b);
    layer0_outputs(3315) <= not (a or b);
    layer0_outputs(3316) <= not (a or b);
    layer0_outputs(3317) <= not (a or b);
    layer0_outputs(3318) <= not (a or b);
    layer0_outputs(3319) <= not b;
    layer0_outputs(3320) <= not (a or b);
    layer0_outputs(3321) <= not a;
    layer0_outputs(3322) <= not b;
    layer0_outputs(3323) <= not b;
    layer0_outputs(3324) <= '0';
    layer0_outputs(3325) <= '0';
    layer0_outputs(3326) <= not a or b;
    layer0_outputs(3327) <= a;
    layer0_outputs(3328) <= '1';
    layer0_outputs(3329) <= a xor b;
    layer0_outputs(3330) <= '1';
    layer0_outputs(3331) <= not (a xor b);
    layer0_outputs(3332) <= '0';
    layer0_outputs(3333) <= not a;
    layer0_outputs(3334) <= '0';
    layer0_outputs(3335) <= not (a and b);
    layer0_outputs(3336) <= b;
    layer0_outputs(3337) <= b;
    layer0_outputs(3338) <= a and b;
    layer0_outputs(3339) <= a;
    layer0_outputs(3340) <= a and b;
    layer0_outputs(3341) <= a and not b;
    layer0_outputs(3342) <= not a or b;
    layer0_outputs(3343) <= not b or a;
    layer0_outputs(3344) <= not a or b;
    layer0_outputs(3345) <= b and not a;
    layer0_outputs(3346) <= not b or a;
    layer0_outputs(3347) <= not (a and b);
    layer0_outputs(3348) <= not (a or b);
    layer0_outputs(3349) <= not a or b;
    layer0_outputs(3350) <= a xor b;
    layer0_outputs(3351) <= a and b;
    layer0_outputs(3352) <= not (a or b);
    layer0_outputs(3353) <= a and b;
    layer0_outputs(3354) <= '1';
    layer0_outputs(3355) <= not b;
    layer0_outputs(3356) <= not (a xor b);
    layer0_outputs(3357) <= b and not a;
    layer0_outputs(3358) <= not b;
    layer0_outputs(3359) <= b;
    layer0_outputs(3360) <= '1';
    layer0_outputs(3361) <= not a or b;
    layer0_outputs(3362) <= not b or a;
    layer0_outputs(3363) <= not a or b;
    layer0_outputs(3364) <= a;
    layer0_outputs(3365) <= not (a and b);
    layer0_outputs(3366) <= not (a or b);
    layer0_outputs(3367) <= a;
    layer0_outputs(3368) <= a;
    layer0_outputs(3369) <= a xor b;
    layer0_outputs(3370) <= a or b;
    layer0_outputs(3371) <= not (a or b);
    layer0_outputs(3372) <= b;
    layer0_outputs(3373) <= '1';
    layer0_outputs(3374) <= not a;
    layer0_outputs(3375) <= not (a or b);
    layer0_outputs(3376) <= not a or b;
    layer0_outputs(3377) <= a or b;
    layer0_outputs(3378) <= '0';
    layer0_outputs(3379) <= a xor b;
    layer0_outputs(3380) <= b;
    layer0_outputs(3381) <= not a or b;
    layer0_outputs(3382) <= '1';
    layer0_outputs(3383) <= not b;
    layer0_outputs(3384) <= '0';
    layer0_outputs(3385) <= a and b;
    layer0_outputs(3386) <= not a or b;
    layer0_outputs(3387) <= not b;
    layer0_outputs(3388) <= b and not a;
    layer0_outputs(3389) <= not a or b;
    layer0_outputs(3390) <= a;
    layer0_outputs(3391) <= not a;
    layer0_outputs(3392) <= b and not a;
    layer0_outputs(3393) <= a xor b;
    layer0_outputs(3394) <= not a;
    layer0_outputs(3395) <= a xor b;
    layer0_outputs(3396) <= a xor b;
    layer0_outputs(3397) <= '0';
    layer0_outputs(3398) <= not b or a;
    layer0_outputs(3399) <= '0';
    layer0_outputs(3400) <= a;
    layer0_outputs(3401) <= b;
    layer0_outputs(3402) <= a;
    layer0_outputs(3403) <= b;
    layer0_outputs(3404) <= not (a and b);
    layer0_outputs(3405) <= a or b;
    layer0_outputs(3406) <= a and not b;
    layer0_outputs(3407) <= '0';
    layer0_outputs(3408) <= a and b;
    layer0_outputs(3409) <= b and not a;
    layer0_outputs(3410) <= a xor b;
    layer0_outputs(3411) <= not a;
    layer0_outputs(3412) <= '1';
    layer0_outputs(3413) <= not b;
    layer0_outputs(3414) <= a or b;
    layer0_outputs(3415) <= a or b;
    layer0_outputs(3416) <= b and not a;
    layer0_outputs(3417) <= not (a or b);
    layer0_outputs(3418) <= a and not b;
    layer0_outputs(3419) <= not b or a;
    layer0_outputs(3420) <= b;
    layer0_outputs(3421) <= a;
    layer0_outputs(3422) <= not (a xor b);
    layer0_outputs(3423) <= not b or a;
    layer0_outputs(3424) <= a and not b;
    layer0_outputs(3425) <= not a or b;
    layer0_outputs(3426) <= b and not a;
    layer0_outputs(3427) <= not (a xor b);
    layer0_outputs(3428) <= a or b;
    layer0_outputs(3429) <= not a;
    layer0_outputs(3430) <= not (a or b);
    layer0_outputs(3431) <= not (a and b);
    layer0_outputs(3432) <= '0';
    layer0_outputs(3433) <= '0';
    layer0_outputs(3434) <= a or b;
    layer0_outputs(3435) <= not b or a;
    layer0_outputs(3436) <= b and not a;
    layer0_outputs(3437) <= '1';
    layer0_outputs(3438) <= a and not b;
    layer0_outputs(3439) <= a and b;
    layer0_outputs(3440) <= a xor b;
    layer0_outputs(3441) <= a or b;
    layer0_outputs(3442) <= b and not a;
    layer0_outputs(3443) <= not (a or b);
    layer0_outputs(3444) <= not (a xor b);
    layer0_outputs(3445) <= b and not a;
    layer0_outputs(3446) <= a and b;
    layer0_outputs(3447) <= not a;
    layer0_outputs(3448) <= '0';
    layer0_outputs(3449) <= not (a xor b);
    layer0_outputs(3450) <= b;
    layer0_outputs(3451) <= not b or a;
    layer0_outputs(3452) <= not (a and b);
    layer0_outputs(3453) <= a xor b;
    layer0_outputs(3454) <= not b or a;
    layer0_outputs(3455) <= '1';
    layer0_outputs(3456) <= a;
    layer0_outputs(3457) <= '0';
    layer0_outputs(3458) <= not (a and b);
    layer0_outputs(3459) <= '0';
    layer0_outputs(3460) <= not b or a;
    layer0_outputs(3461) <= a and b;
    layer0_outputs(3462) <= a and not b;
    layer0_outputs(3463) <= b;
    layer0_outputs(3464) <= not b or a;
    layer0_outputs(3465) <= a;
    layer0_outputs(3466) <= not b or a;
    layer0_outputs(3467) <= a;
    layer0_outputs(3468) <= b;
    layer0_outputs(3469) <= a and not b;
    layer0_outputs(3470) <= a and not b;
    layer0_outputs(3471) <= not (a or b);
    layer0_outputs(3472) <= not (a or b);
    layer0_outputs(3473) <= '0';
    layer0_outputs(3474) <= not b;
    layer0_outputs(3475) <= not a or b;
    layer0_outputs(3476) <= not b or a;
    layer0_outputs(3477) <= '1';
    layer0_outputs(3478) <= a and not b;
    layer0_outputs(3479) <= not b or a;
    layer0_outputs(3480) <= not b;
    layer0_outputs(3481) <= not b or a;
    layer0_outputs(3482) <= a xor b;
    layer0_outputs(3483) <= a;
    layer0_outputs(3484) <= not b or a;
    layer0_outputs(3485) <= a and not b;
    layer0_outputs(3486) <= not b;
    layer0_outputs(3487) <= not (a and b);
    layer0_outputs(3488) <= a xor b;
    layer0_outputs(3489) <= not a;
    layer0_outputs(3490) <= not (a and b);
    layer0_outputs(3491) <= '1';
    layer0_outputs(3492) <= not b;
    layer0_outputs(3493) <= '0';
    layer0_outputs(3494) <= not (a and b);
    layer0_outputs(3495) <= not a or b;
    layer0_outputs(3496) <= not b or a;
    layer0_outputs(3497) <= a xor b;
    layer0_outputs(3498) <= not a or b;
    layer0_outputs(3499) <= a or b;
    layer0_outputs(3500) <= b;
    layer0_outputs(3501) <= not b or a;
    layer0_outputs(3502) <= a or b;
    layer0_outputs(3503) <= a and not b;
    layer0_outputs(3504) <= not (a or b);
    layer0_outputs(3505) <= not (a xor b);
    layer0_outputs(3506) <= not b;
    layer0_outputs(3507) <= b and not a;
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= not (a or b);
    layer0_outputs(3510) <= not (a or b);
    layer0_outputs(3511) <= a and not b;
    layer0_outputs(3512) <= '0';
    layer0_outputs(3513) <= not b or a;
    layer0_outputs(3514) <= '1';
    layer0_outputs(3515) <= not (a or b);
    layer0_outputs(3516) <= a;
    layer0_outputs(3517) <= a and b;
    layer0_outputs(3518) <= not (a or b);
    layer0_outputs(3519) <= a and b;
    layer0_outputs(3520) <= a or b;
    layer0_outputs(3521) <= not (a xor b);
    layer0_outputs(3522) <= '1';
    layer0_outputs(3523) <= not b or a;
    layer0_outputs(3524) <= '0';
    layer0_outputs(3525) <= not b;
    layer0_outputs(3526) <= a xor b;
    layer0_outputs(3527) <= '0';
    layer0_outputs(3528) <= not (a or b);
    layer0_outputs(3529) <= '1';
    layer0_outputs(3530) <= a;
    layer0_outputs(3531) <= not (a xor b);
    layer0_outputs(3532) <= '0';
    layer0_outputs(3533) <= not a or b;
    layer0_outputs(3534) <= a or b;
    layer0_outputs(3535) <= not b or a;
    layer0_outputs(3536) <= not b;
    layer0_outputs(3537) <= not (a xor b);
    layer0_outputs(3538) <= b and not a;
    layer0_outputs(3539) <= not b or a;
    layer0_outputs(3540) <= not b;
    layer0_outputs(3541) <= not b;
    layer0_outputs(3542) <= a and not b;
    layer0_outputs(3543) <= not b;
    layer0_outputs(3544) <= not (a xor b);
    layer0_outputs(3545) <= a or b;
    layer0_outputs(3546) <= not (a or b);
    layer0_outputs(3547) <= b;
    layer0_outputs(3548) <= b and not a;
    layer0_outputs(3549) <= b;
    layer0_outputs(3550) <= not b;
    layer0_outputs(3551) <= not b or a;
    layer0_outputs(3552) <= not (a and b);
    layer0_outputs(3553) <= not (a and b);
    layer0_outputs(3554) <= not b;
    layer0_outputs(3555) <= not (a xor b);
    layer0_outputs(3556) <= not b;
    layer0_outputs(3557) <= not a or b;
    layer0_outputs(3558) <= not b or a;
    layer0_outputs(3559) <= b and not a;
    layer0_outputs(3560) <= b and not a;
    layer0_outputs(3561) <= not b or a;
    layer0_outputs(3562) <= not a or b;
    layer0_outputs(3563) <= not a;
    layer0_outputs(3564) <= not (a or b);
    layer0_outputs(3565) <= not a;
    layer0_outputs(3566) <= a and not b;
    layer0_outputs(3567) <= not b or a;
    layer0_outputs(3568) <= not (a or b);
    layer0_outputs(3569) <= not (a or b);
    layer0_outputs(3570) <= a or b;
    layer0_outputs(3571) <= b and not a;
    layer0_outputs(3572) <= not a;
    layer0_outputs(3573) <= not (a or b);
    layer0_outputs(3574) <= '1';
    layer0_outputs(3575) <= a;
    layer0_outputs(3576) <= not b or a;
    layer0_outputs(3577) <= a or b;
    layer0_outputs(3578) <= not b;
    layer0_outputs(3579) <= a and b;
    layer0_outputs(3580) <= a and not b;
    layer0_outputs(3581) <= not a;
    layer0_outputs(3582) <= not (a or b);
    layer0_outputs(3583) <= '1';
    layer0_outputs(3584) <= not a;
    layer0_outputs(3585) <= '1';
    layer0_outputs(3586) <= a xor b;
    layer0_outputs(3587) <= a;
    layer0_outputs(3588) <= not b;
    layer0_outputs(3589) <= not (a and b);
    layer0_outputs(3590) <= not (a and b);
    layer0_outputs(3591) <= not a or b;
    layer0_outputs(3592) <= '1';
    layer0_outputs(3593) <= a;
    layer0_outputs(3594) <= not a or b;
    layer0_outputs(3595) <= a and b;
    layer0_outputs(3596) <= not b;
    layer0_outputs(3597) <= not (a or b);
    layer0_outputs(3598) <= not a;
    layer0_outputs(3599) <= not (a or b);
    layer0_outputs(3600) <= not (a and b);
    layer0_outputs(3601) <= not a or b;
    layer0_outputs(3602) <= not b or a;
    layer0_outputs(3603) <= '1';
    layer0_outputs(3604) <= '1';
    layer0_outputs(3605) <= a and b;
    layer0_outputs(3606) <= a xor b;
    layer0_outputs(3607) <= not b;
    layer0_outputs(3608) <= a and b;
    layer0_outputs(3609) <= not a;
    layer0_outputs(3610) <= a and not b;
    layer0_outputs(3611) <= not (a and b);
    layer0_outputs(3612) <= a and not b;
    layer0_outputs(3613) <= not (a or b);
    layer0_outputs(3614) <= not a or b;
    layer0_outputs(3615) <= '1';
    layer0_outputs(3616) <= not b or a;
    layer0_outputs(3617) <= b and not a;
    layer0_outputs(3618) <= not b or a;
    layer0_outputs(3619) <= not (a and b);
    layer0_outputs(3620) <= not (a xor b);
    layer0_outputs(3621) <= not b or a;
    layer0_outputs(3622) <= '1';
    layer0_outputs(3623) <= b;
    layer0_outputs(3624) <= '1';
    layer0_outputs(3625) <= b;
    layer0_outputs(3626) <= not a;
    layer0_outputs(3627) <= '1';
    layer0_outputs(3628) <= not a;
    layer0_outputs(3629) <= not (a xor b);
    layer0_outputs(3630) <= b;
    layer0_outputs(3631) <= not a or b;
    layer0_outputs(3632) <= not b;
    layer0_outputs(3633) <= not (a and b);
    layer0_outputs(3634) <= '0';
    layer0_outputs(3635) <= not a or b;
    layer0_outputs(3636) <= not b or a;
    layer0_outputs(3637) <= '1';
    layer0_outputs(3638) <= not a or b;
    layer0_outputs(3639) <= b and not a;
    layer0_outputs(3640) <= a xor b;
    layer0_outputs(3641) <= not a;
    layer0_outputs(3642) <= a and not b;
    layer0_outputs(3643) <= not a;
    layer0_outputs(3644) <= a;
    layer0_outputs(3645) <= '0';
    layer0_outputs(3646) <= not (a and b);
    layer0_outputs(3647) <= b;
    layer0_outputs(3648) <= '1';
    layer0_outputs(3649) <= not (a xor b);
    layer0_outputs(3650) <= b;
    layer0_outputs(3651) <= not (a and b);
    layer0_outputs(3652) <= '0';
    layer0_outputs(3653) <= '0';
    layer0_outputs(3654) <= a or b;
    layer0_outputs(3655) <= a and not b;
    layer0_outputs(3656) <= a or b;
    layer0_outputs(3657) <= not b;
    layer0_outputs(3658) <= a;
    layer0_outputs(3659) <= a or b;
    layer0_outputs(3660) <= '1';
    layer0_outputs(3661) <= not (a and b);
    layer0_outputs(3662) <= a;
    layer0_outputs(3663) <= not b or a;
    layer0_outputs(3664) <= not (a or b);
    layer0_outputs(3665) <= not (a xor b);
    layer0_outputs(3666) <= '0';
    layer0_outputs(3667) <= a;
    layer0_outputs(3668) <= a xor b;
    layer0_outputs(3669) <= a and b;
    layer0_outputs(3670) <= not (a and b);
    layer0_outputs(3671) <= a and b;
    layer0_outputs(3672) <= not a;
    layer0_outputs(3673) <= not b or a;
    layer0_outputs(3674) <= not b or a;
    layer0_outputs(3675) <= not b;
    layer0_outputs(3676) <= a or b;
    layer0_outputs(3677) <= not (a and b);
    layer0_outputs(3678) <= not b;
    layer0_outputs(3679) <= a or b;
    layer0_outputs(3680) <= a and b;
    layer0_outputs(3681) <= b and not a;
    layer0_outputs(3682) <= not a or b;
    layer0_outputs(3683) <= a or b;
    layer0_outputs(3684) <= a;
    layer0_outputs(3685) <= b and not a;
    layer0_outputs(3686) <= '1';
    layer0_outputs(3687) <= b and not a;
    layer0_outputs(3688) <= a or b;
    layer0_outputs(3689) <= not (a or b);
    layer0_outputs(3690) <= b and not a;
    layer0_outputs(3691) <= '0';
    layer0_outputs(3692) <= a;
    layer0_outputs(3693) <= '0';
    layer0_outputs(3694) <= b and not a;
    layer0_outputs(3695) <= '1';
    layer0_outputs(3696) <= '0';
    layer0_outputs(3697) <= not (a or b);
    layer0_outputs(3698) <= a;
    layer0_outputs(3699) <= a xor b;
    layer0_outputs(3700) <= not a or b;
    layer0_outputs(3701) <= a and not b;
    layer0_outputs(3702) <= not b;
    layer0_outputs(3703) <= '1';
    layer0_outputs(3704) <= not (a xor b);
    layer0_outputs(3705) <= not a or b;
    layer0_outputs(3706) <= a and not b;
    layer0_outputs(3707) <= not (a xor b);
    layer0_outputs(3708) <= b;
    layer0_outputs(3709) <= a xor b;
    layer0_outputs(3710) <= b;
    layer0_outputs(3711) <= a;
    layer0_outputs(3712) <= a;
    layer0_outputs(3713) <= b and not a;
    layer0_outputs(3714) <= not a or b;
    layer0_outputs(3715) <= a and not b;
    layer0_outputs(3716) <= not b or a;
    layer0_outputs(3717) <= not (a xor b);
    layer0_outputs(3718) <= a or b;
    layer0_outputs(3719) <= a;
    layer0_outputs(3720) <= not b or a;
    layer0_outputs(3721) <= a and b;
    layer0_outputs(3722) <= not (a or b);
    layer0_outputs(3723) <= b and not a;
    layer0_outputs(3724) <= not (a or b);
    layer0_outputs(3725) <= a xor b;
    layer0_outputs(3726) <= not a;
    layer0_outputs(3727) <= '1';
    layer0_outputs(3728) <= a and not b;
    layer0_outputs(3729) <= '0';
    layer0_outputs(3730) <= a and not b;
    layer0_outputs(3731) <= not a;
    layer0_outputs(3732) <= '1';
    layer0_outputs(3733) <= a;
    layer0_outputs(3734) <= a or b;
    layer0_outputs(3735) <= a and b;
    layer0_outputs(3736) <= a and b;
    layer0_outputs(3737) <= not a or b;
    layer0_outputs(3738) <= not a;
    layer0_outputs(3739) <= a and not b;
    layer0_outputs(3740) <= a;
    layer0_outputs(3741) <= '0';
    layer0_outputs(3742) <= not (a xor b);
    layer0_outputs(3743) <= not b or a;
    layer0_outputs(3744) <= not a;
    layer0_outputs(3745) <= a and b;
    layer0_outputs(3746) <= not (a or b);
    layer0_outputs(3747) <= not b or a;
    layer0_outputs(3748) <= not b or a;
    layer0_outputs(3749) <= not (a or b);
    layer0_outputs(3750) <= b and not a;
    layer0_outputs(3751) <= not (a or b);
    layer0_outputs(3752) <= not b;
    layer0_outputs(3753) <= '0';
    layer0_outputs(3754) <= a and not b;
    layer0_outputs(3755) <= a and b;
    layer0_outputs(3756) <= not (a or b);
    layer0_outputs(3757) <= a and not b;
    layer0_outputs(3758) <= not (a or b);
    layer0_outputs(3759) <= not b;
    layer0_outputs(3760) <= a and not b;
    layer0_outputs(3761) <= '0';
    layer0_outputs(3762) <= '0';
    layer0_outputs(3763) <= not (a or b);
    layer0_outputs(3764) <= a;
    layer0_outputs(3765) <= '0';
    layer0_outputs(3766) <= a or b;
    layer0_outputs(3767) <= not b or a;
    layer0_outputs(3768) <= not b;
    layer0_outputs(3769) <= '0';
    layer0_outputs(3770) <= not b or a;
    layer0_outputs(3771) <= b;
    layer0_outputs(3772) <= not a;
    layer0_outputs(3773) <= not b;
    layer0_outputs(3774) <= '0';
    layer0_outputs(3775) <= '0';
    layer0_outputs(3776) <= b and not a;
    layer0_outputs(3777) <= not a or b;
    layer0_outputs(3778) <= not a or b;
    layer0_outputs(3779) <= a and b;
    layer0_outputs(3780) <= b and not a;
    layer0_outputs(3781) <= not (a or b);
    layer0_outputs(3782) <= a and not b;
    layer0_outputs(3783) <= b;
    layer0_outputs(3784) <= not (a or b);
    layer0_outputs(3785) <= '1';
    layer0_outputs(3786) <= a xor b;
    layer0_outputs(3787) <= '1';
    layer0_outputs(3788) <= b and not a;
    layer0_outputs(3789) <= a and b;
    layer0_outputs(3790) <= a and not b;
    layer0_outputs(3791) <= not (a or b);
    layer0_outputs(3792) <= not b;
    layer0_outputs(3793) <= b;
    layer0_outputs(3794) <= b;
    layer0_outputs(3795) <= '1';
    layer0_outputs(3796) <= a and b;
    layer0_outputs(3797) <= '1';
    layer0_outputs(3798) <= a and not b;
    layer0_outputs(3799) <= not b;
    layer0_outputs(3800) <= not (a xor b);
    layer0_outputs(3801) <= not a;
    layer0_outputs(3802) <= b and not a;
    layer0_outputs(3803) <= a or b;
    layer0_outputs(3804) <= not (a and b);
    layer0_outputs(3805) <= not (a and b);
    layer0_outputs(3806) <= b;
    layer0_outputs(3807) <= not a;
    layer0_outputs(3808) <= not b;
    layer0_outputs(3809) <= not (a and b);
    layer0_outputs(3810) <= b;
    layer0_outputs(3811) <= not a;
    layer0_outputs(3812) <= not b;
    layer0_outputs(3813) <= a xor b;
    layer0_outputs(3814) <= a and b;
    layer0_outputs(3815) <= a and not b;
    layer0_outputs(3816) <= a xor b;
    layer0_outputs(3817) <= a;
    layer0_outputs(3818) <= a and b;
    layer0_outputs(3819) <= not (a and b);
    layer0_outputs(3820) <= b;
    layer0_outputs(3821) <= not (a or b);
    layer0_outputs(3822) <= '1';
    layer0_outputs(3823) <= a and b;
    layer0_outputs(3824) <= '0';
    layer0_outputs(3825) <= a and b;
    layer0_outputs(3826) <= b and not a;
    layer0_outputs(3827) <= a and not b;
    layer0_outputs(3828) <= not b or a;
    layer0_outputs(3829) <= a and not b;
    layer0_outputs(3830) <= not b or a;
    layer0_outputs(3831) <= not (a or b);
    layer0_outputs(3832) <= not (a or b);
    layer0_outputs(3833) <= a and b;
    layer0_outputs(3834) <= a;
    layer0_outputs(3835) <= a or b;
    layer0_outputs(3836) <= not (a and b);
    layer0_outputs(3837) <= not (a or b);
    layer0_outputs(3838) <= not (a and b);
    layer0_outputs(3839) <= a and not b;
    layer0_outputs(3840) <= not b;
    layer0_outputs(3841) <= a and b;
    layer0_outputs(3842) <= a or b;
    layer0_outputs(3843) <= b;
    layer0_outputs(3844) <= not (a and b);
    layer0_outputs(3845) <= not a or b;
    layer0_outputs(3846) <= not a or b;
    layer0_outputs(3847) <= '1';
    layer0_outputs(3848) <= a xor b;
    layer0_outputs(3849) <= b;
    layer0_outputs(3850) <= a xor b;
    layer0_outputs(3851) <= a and b;
    layer0_outputs(3852) <= not a;
    layer0_outputs(3853) <= not b;
    layer0_outputs(3854) <= not b or a;
    layer0_outputs(3855) <= '1';
    layer0_outputs(3856) <= not (a xor b);
    layer0_outputs(3857) <= b;
    layer0_outputs(3858) <= not (a xor b);
    layer0_outputs(3859) <= '0';
    layer0_outputs(3860) <= '0';
    layer0_outputs(3861) <= not a;
    layer0_outputs(3862) <= a and b;
    layer0_outputs(3863) <= b and not a;
    layer0_outputs(3864) <= a or b;
    layer0_outputs(3865) <= not b;
    layer0_outputs(3866) <= not b;
    layer0_outputs(3867) <= not a or b;
    layer0_outputs(3868) <= not a;
    layer0_outputs(3869) <= '1';
    layer0_outputs(3870) <= not b or a;
    layer0_outputs(3871) <= a;
    layer0_outputs(3872) <= a and not b;
    layer0_outputs(3873) <= a and b;
    layer0_outputs(3874) <= not (a and b);
    layer0_outputs(3875) <= not b or a;
    layer0_outputs(3876) <= a and not b;
    layer0_outputs(3877) <= a and not b;
    layer0_outputs(3878) <= a and b;
    layer0_outputs(3879) <= a or b;
    layer0_outputs(3880) <= b;
    layer0_outputs(3881) <= '1';
    layer0_outputs(3882) <= a and b;
    layer0_outputs(3883) <= not (a or b);
    layer0_outputs(3884) <= not a;
    layer0_outputs(3885) <= not (a or b);
    layer0_outputs(3886) <= a xor b;
    layer0_outputs(3887) <= a and b;
    layer0_outputs(3888) <= not a;
    layer0_outputs(3889) <= '0';
    layer0_outputs(3890) <= not b or a;
    layer0_outputs(3891) <= not (a or b);
    layer0_outputs(3892) <= not b;
    layer0_outputs(3893) <= b and not a;
    layer0_outputs(3894) <= not b or a;
    layer0_outputs(3895) <= not a;
    layer0_outputs(3896) <= '0';
    layer0_outputs(3897) <= not (a xor b);
    layer0_outputs(3898) <= a;
    layer0_outputs(3899) <= not (a and b);
    layer0_outputs(3900) <= a and not b;
    layer0_outputs(3901) <= not a;
    layer0_outputs(3902) <= a and b;
    layer0_outputs(3903) <= a and b;
    layer0_outputs(3904) <= not a or b;
    layer0_outputs(3905) <= not a or b;
    layer0_outputs(3906) <= not (a xor b);
    layer0_outputs(3907) <= '1';
    layer0_outputs(3908) <= a xor b;
    layer0_outputs(3909) <= a xor b;
    layer0_outputs(3910) <= a and not b;
    layer0_outputs(3911) <= b;
    layer0_outputs(3912) <= not b or a;
    layer0_outputs(3913) <= not a;
    layer0_outputs(3914) <= not b;
    layer0_outputs(3915) <= not (a or b);
    layer0_outputs(3916) <= a xor b;
    layer0_outputs(3917) <= b and not a;
    layer0_outputs(3918) <= not (a and b);
    layer0_outputs(3919) <= not b or a;
    layer0_outputs(3920) <= b;
    layer0_outputs(3921) <= b and not a;
    layer0_outputs(3922) <= a;
    layer0_outputs(3923) <= not (a xor b);
    layer0_outputs(3924) <= '0';
    layer0_outputs(3925) <= not a;
    layer0_outputs(3926) <= a;
    layer0_outputs(3927) <= not (a or b);
    layer0_outputs(3928) <= '1';
    layer0_outputs(3929) <= not a or b;
    layer0_outputs(3930) <= a xor b;
    layer0_outputs(3931) <= '0';
    layer0_outputs(3932) <= b;
    layer0_outputs(3933) <= not (a or b);
    layer0_outputs(3934) <= not (a or b);
    layer0_outputs(3935) <= not a;
    layer0_outputs(3936) <= '0';
    layer0_outputs(3937) <= not a;
    layer0_outputs(3938) <= a and b;
    layer0_outputs(3939) <= not a or b;
    layer0_outputs(3940) <= not b or a;
    layer0_outputs(3941) <= a;
    layer0_outputs(3942) <= not a or b;
    layer0_outputs(3943) <= not a;
    layer0_outputs(3944) <= not a or b;
    layer0_outputs(3945) <= '1';
    layer0_outputs(3946) <= not b;
    layer0_outputs(3947) <= a or b;
    layer0_outputs(3948) <= '1';
    layer0_outputs(3949) <= not a or b;
    layer0_outputs(3950) <= a and not b;
    layer0_outputs(3951) <= '0';
    layer0_outputs(3952) <= a or b;
    layer0_outputs(3953) <= '0';
    layer0_outputs(3954) <= a;
    layer0_outputs(3955) <= '1';
    layer0_outputs(3956) <= not a;
    layer0_outputs(3957) <= a or b;
    layer0_outputs(3958) <= b and not a;
    layer0_outputs(3959) <= not b;
    layer0_outputs(3960) <= not b;
    layer0_outputs(3961) <= a and b;
    layer0_outputs(3962) <= '0';
    layer0_outputs(3963) <= a and not b;
    layer0_outputs(3964) <= a xor b;
    layer0_outputs(3965) <= not (a or b);
    layer0_outputs(3966) <= not b or a;
    layer0_outputs(3967) <= not (a and b);
    layer0_outputs(3968) <= b;
    layer0_outputs(3969) <= a and b;
    layer0_outputs(3970) <= a or b;
    layer0_outputs(3971) <= not a;
    layer0_outputs(3972) <= b;
    layer0_outputs(3973) <= a and b;
    layer0_outputs(3974) <= not b or a;
    layer0_outputs(3975) <= a or b;
    layer0_outputs(3976) <= not b;
    layer0_outputs(3977) <= not (a and b);
    layer0_outputs(3978) <= b;
    layer0_outputs(3979) <= not a;
    layer0_outputs(3980) <= a and b;
    layer0_outputs(3981) <= a or b;
    layer0_outputs(3982) <= a;
    layer0_outputs(3983) <= not (a xor b);
    layer0_outputs(3984) <= a and not b;
    layer0_outputs(3985) <= not (a and b);
    layer0_outputs(3986) <= not b;
    layer0_outputs(3987) <= '1';
    layer0_outputs(3988) <= '0';
    layer0_outputs(3989) <= not b;
    layer0_outputs(3990) <= not (a and b);
    layer0_outputs(3991) <= a and b;
    layer0_outputs(3992) <= a and not b;
    layer0_outputs(3993) <= '1';
    layer0_outputs(3994) <= b and not a;
    layer0_outputs(3995) <= a;
    layer0_outputs(3996) <= '0';
    layer0_outputs(3997) <= a or b;
    layer0_outputs(3998) <= not a or b;
    layer0_outputs(3999) <= b and not a;
    layer0_outputs(4000) <= not a;
    layer0_outputs(4001) <= b and not a;
    layer0_outputs(4002) <= not b or a;
    layer0_outputs(4003) <= a;
    layer0_outputs(4004) <= not (a and b);
    layer0_outputs(4005) <= not a or b;
    layer0_outputs(4006) <= '0';
    layer0_outputs(4007) <= b;
    layer0_outputs(4008) <= '0';
    layer0_outputs(4009) <= a or b;
    layer0_outputs(4010) <= a;
    layer0_outputs(4011) <= b and not a;
    layer0_outputs(4012) <= not (a and b);
    layer0_outputs(4013) <= not b or a;
    layer0_outputs(4014) <= not a;
    layer0_outputs(4015) <= not (a and b);
    layer0_outputs(4016) <= '0';
    layer0_outputs(4017) <= not (a or b);
    layer0_outputs(4018) <= not (a or b);
    layer0_outputs(4019) <= not a or b;
    layer0_outputs(4020) <= '1';
    layer0_outputs(4021) <= '1';
    layer0_outputs(4022) <= a;
    layer0_outputs(4023) <= a xor b;
    layer0_outputs(4024) <= not a or b;
    layer0_outputs(4025) <= not a;
    layer0_outputs(4026) <= not (a xor b);
    layer0_outputs(4027) <= a or b;
    layer0_outputs(4028) <= a;
    layer0_outputs(4029) <= not (a or b);
    layer0_outputs(4030) <= not (a and b);
    layer0_outputs(4031) <= a or b;
    layer0_outputs(4032) <= a or b;
    layer0_outputs(4033) <= a or b;
    layer0_outputs(4034) <= '1';
    layer0_outputs(4035) <= '1';
    layer0_outputs(4036) <= a xor b;
    layer0_outputs(4037) <= not b or a;
    layer0_outputs(4038) <= not (a xor b);
    layer0_outputs(4039) <= '0';
    layer0_outputs(4040) <= '1';
    layer0_outputs(4041) <= a and b;
    layer0_outputs(4042) <= not b;
    layer0_outputs(4043) <= not a or b;
    layer0_outputs(4044) <= not (a and b);
    layer0_outputs(4045) <= a xor b;
    layer0_outputs(4046) <= not (a xor b);
    layer0_outputs(4047) <= not b or a;
    layer0_outputs(4048) <= a or b;
    layer0_outputs(4049) <= not (a or b);
    layer0_outputs(4050) <= '0';
    layer0_outputs(4051) <= a or b;
    layer0_outputs(4052) <= b;
    layer0_outputs(4053) <= not a;
    layer0_outputs(4054) <= not (a or b);
    layer0_outputs(4055) <= '1';
    layer0_outputs(4056) <= b and not a;
    layer0_outputs(4057) <= b and not a;
    layer0_outputs(4058) <= not a;
    layer0_outputs(4059) <= b;
    layer0_outputs(4060) <= a or b;
    layer0_outputs(4061) <= not (a and b);
    layer0_outputs(4062) <= '1';
    layer0_outputs(4063) <= b and not a;
    layer0_outputs(4064) <= a and not b;
    layer0_outputs(4065) <= a and not b;
    layer0_outputs(4066) <= not (a and b);
    layer0_outputs(4067) <= b;
    layer0_outputs(4068) <= b;
    layer0_outputs(4069) <= a xor b;
    layer0_outputs(4070) <= a;
    layer0_outputs(4071) <= a;
    layer0_outputs(4072) <= not a or b;
    layer0_outputs(4073) <= b;
    layer0_outputs(4074) <= not (a and b);
    layer0_outputs(4075) <= not a;
    layer0_outputs(4076) <= not b or a;
    layer0_outputs(4077) <= b;
    layer0_outputs(4078) <= b and not a;
    layer0_outputs(4079) <= not (a xor b);
    layer0_outputs(4080) <= not (a or b);
    layer0_outputs(4081) <= b;
    layer0_outputs(4082) <= a and not b;
    layer0_outputs(4083) <= not b;
    layer0_outputs(4084) <= not a or b;
    layer0_outputs(4085) <= not b;
    layer0_outputs(4086) <= not b;
    layer0_outputs(4087) <= a or b;
    layer0_outputs(4088) <= not a or b;
    layer0_outputs(4089) <= not (a or b);
    layer0_outputs(4090) <= not (a xor b);
    layer0_outputs(4091) <= a;
    layer0_outputs(4092) <= not a or b;
    layer0_outputs(4093) <= not (a xor b);
    layer0_outputs(4094) <= not b or a;
    layer0_outputs(4095) <= a xor b;
    layer0_outputs(4096) <= a and not b;
    layer0_outputs(4097) <= not a;
    layer0_outputs(4098) <= not (a or b);
    layer0_outputs(4099) <= a and b;
    layer0_outputs(4100) <= a and not b;
    layer0_outputs(4101) <= not a;
    layer0_outputs(4102) <= not a;
    layer0_outputs(4103) <= a or b;
    layer0_outputs(4104) <= b and not a;
    layer0_outputs(4105) <= b;
    layer0_outputs(4106) <= b;
    layer0_outputs(4107) <= '0';
    layer0_outputs(4108) <= a or b;
    layer0_outputs(4109) <= a and not b;
    layer0_outputs(4110) <= not (a xor b);
    layer0_outputs(4111) <= '1';
    layer0_outputs(4112) <= '0';
    layer0_outputs(4113) <= not (a and b);
    layer0_outputs(4114) <= not (a xor b);
    layer0_outputs(4115) <= a;
    layer0_outputs(4116) <= a and b;
    layer0_outputs(4117) <= a and not b;
    layer0_outputs(4118) <= not a;
    layer0_outputs(4119) <= b and not a;
    layer0_outputs(4120) <= a and not b;
    layer0_outputs(4121) <= a and b;
    layer0_outputs(4122) <= not a;
    layer0_outputs(4123) <= a and not b;
    layer0_outputs(4124) <= not b;
    layer0_outputs(4125) <= a xor b;
    layer0_outputs(4126) <= not (a and b);
    layer0_outputs(4127) <= not a or b;
    layer0_outputs(4128) <= '1';
    layer0_outputs(4129) <= not b;
    layer0_outputs(4130) <= not (a and b);
    layer0_outputs(4131) <= '0';
    layer0_outputs(4132) <= not a;
    layer0_outputs(4133) <= a xor b;
    layer0_outputs(4134) <= a or b;
    layer0_outputs(4135) <= not (a or b);
    layer0_outputs(4136) <= a;
    layer0_outputs(4137) <= not (a and b);
    layer0_outputs(4138) <= not a;
    layer0_outputs(4139) <= not (a and b);
    layer0_outputs(4140) <= a and b;
    layer0_outputs(4141) <= b and not a;
    layer0_outputs(4142) <= b and not a;
    layer0_outputs(4143) <= a and not b;
    layer0_outputs(4144) <= not b;
    layer0_outputs(4145) <= not (a xor b);
    layer0_outputs(4146) <= b;
    layer0_outputs(4147) <= not (a and b);
    layer0_outputs(4148) <= not a;
    layer0_outputs(4149) <= a or b;
    layer0_outputs(4150) <= not a;
    layer0_outputs(4151) <= '1';
    layer0_outputs(4152) <= not a or b;
    layer0_outputs(4153) <= not (a and b);
    layer0_outputs(4154) <= '1';
    layer0_outputs(4155) <= not (a xor b);
    layer0_outputs(4156) <= '0';
    layer0_outputs(4157) <= '0';
    layer0_outputs(4158) <= a;
    layer0_outputs(4159) <= a and not b;
    layer0_outputs(4160) <= a or b;
    layer0_outputs(4161) <= b and not a;
    layer0_outputs(4162) <= a xor b;
    layer0_outputs(4163) <= a and not b;
    layer0_outputs(4164) <= a and b;
    layer0_outputs(4165) <= b and not a;
    layer0_outputs(4166) <= '1';
    layer0_outputs(4167) <= not (a and b);
    layer0_outputs(4168) <= '0';
    layer0_outputs(4169) <= not a;
    layer0_outputs(4170) <= '1';
    layer0_outputs(4171) <= a and b;
    layer0_outputs(4172) <= not b;
    layer0_outputs(4173) <= '1';
    layer0_outputs(4174) <= b and not a;
    layer0_outputs(4175) <= '0';
    layer0_outputs(4176) <= a;
    layer0_outputs(4177) <= b and not a;
    layer0_outputs(4178) <= b and not a;
    layer0_outputs(4179) <= a;
    layer0_outputs(4180) <= a and not b;
    layer0_outputs(4181) <= b and not a;
    layer0_outputs(4182) <= not (a and b);
    layer0_outputs(4183) <= a and b;
    layer0_outputs(4184) <= '1';
    layer0_outputs(4185) <= '0';
    layer0_outputs(4186) <= '0';
    layer0_outputs(4187) <= not (a xor b);
    layer0_outputs(4188) <= not b;
    layer0_outputs(4189) <= a and not b;
    layer0_outputs(4190) <= '1';
    layer0_outputs(4191) <= not (a or b);
    layer0_outputs(4192) <= a and b;
    layer0_outputs(4193) <= not (a and b);
    layer0_outputs(4194) <= '1';
    layer0_outputs(4195) <= a or b;
    layer0_outputs(4196) <= '1';
    layer0_outputs(4197) <= b;
    layer0_outputs(4198) <= b;
    layer0_outputs(4199) <= '1';
    layer0_outputs(4200) <= not (a xor b);
    layer0_outputs(4201) <= b;
    layer0_outputs(4202) <= not (a and b);
    layer0_outputs(4203) <= not b or a;
    layer0_outputs(4204) <= not b;
    layer0_outputs(4205) <= a or b;
    layer0_outputs(4206) <= '0';
    layer0_outputs(4207) <= a;
    layer0_outputs(4208) <= a;
    layer0_outputs(4209) <= a and b;
    layer0_outputs(4210) <= not b or a;
    layer0_outputs(4211) <= b and not a;
    layer0_outputs(4212) <= not b;
    layer0_outputs(4213) <= a;
    layer0_outputs(4214) <= '0';
    layer0_outputs(4215) <= not b;
    layer0_outputs(4216) <= a and not b;
    layer0_outputs(4217) <= b;
    layer0_outputs(4218) <= a xor b;
    layer0_outputs(4219) <= '1';
    layer0_outputs(4220) <= '1';
    layer0_outputs(4221) <= a;
    layer0_outputs(4222) <= a and not b;
    layer0_outputs(4223) <= b;
    layer0_outputs(4224) <= not a;
    layer0_outputs(4225) <= not b or a;
    layer0_outputs(4226) <= '1';
    layer0_outputs(4227) <= a xor b;
    layer0_outputs(4228) <= not (a or b);
    layer0_outputs(4229) <= not (a or b);
    layer0_outputs(4230) <= '0';
    layer0_outputs(4231) <= not a or b;
    layer0_outputs(4232) <= b and not a;
    layer0_outputs(4233) <= b;
    layer0_outputs(4234) <= a or b;
    layer0_outputs(4235) <= not b or a;
    layer0_outputs(4236) <= a or b;
    layer0_outputs(4237) <= not (a xor b);
    layer0_outputs(4238) <= b;
    layer0_outputs(4239) <= not a;
    layer0_outputs(4240) <= b and not a;
    layer0_outputs(4241) <= not a or b;
    layer0_outputs(4242) <= not b or a;
    layer0_outputs(4243) <= not a;
    layer0_outputs(4244) <= not (a xor b);
    layer0_outputs(4245) <= not (a xor b);
    layer0_outputs(4246) <= b;
    layer0_outputs(4247) <= not (a or b);
    layer0_outputs(4248) <= '0';
    layer0_outputs(4249) <= not (a and b);
    layer0_outputs(4250) <= not (a or b);
    layer0_outputs(4251) <= b;
    layer0_outputs(4252) <= not b;
    layer0_outputs(4253) <= a;
    layer0_outputs(4254) <= b;
    layer0_outputs(4255) <= a or b;
    layer0_outputs(4256) <= a;
    layer0_outputs(4257) <= '1';
    layer0_outputs(4258) <= not (a xor b);
    layer0_outputs(4259) <= a or b;
    layer0_outputs(4260) <= a;
    layer0_outputs(4261) <= a and not b;
    layer0_outputs(4262) <= b;
    layer0_outputs(4263) <= not (a or b);
    layer0_outputs(4264) <= not (a and b);
    layer0_outputs(4265) <= b;
    layer0_outputs(4266) <= a xor b;
    layer0_outputs(4267) <= not (a and b);
    layer0_outputs(4268) <= not a or b;
    layer0_outputs(4269) <= not (a or b);
    layer0_outputs(4270) <= not (a xor b);
    layer0_outputs(4271) <= a xor b;
    layer0_outputs(4272) <= not b;
    layer0_outputs(4273) <= a;
    layer0_outputs(4274) <= '0';
    layer0_outputs(4275) <= b and not a;
    layer0_outputs(4276) <= a or b;
    layer0_outputs(4277) <= b;
    layer0_outputs(4278) <= a xor b;
    layer0_outputs(4279) <= not (a xor b);
    layer0_outputs(4280) <= not (a xor b);
    layer0_outputs(4281) <= a and not b;
    layer0_outputs(4282) <= '1';
    layer0_outputs(4283) <= not (a and b);
    layer0_outputs(4284) <= a;
    layer0_outputs(4285) <= not a or b;
    layer0_outputs(4286) <= not a;
    layer0_outputs(4287) <= a;
    layer0_outputs(4288) <= b and not a;
    layer0_outputs(4289) <= a;
    layer0_outputs(4290) <= '1';
    layer0_outputs(4291) <= not b or a;
    layer0_outputs(4292) <= '0';
    layer0_outputs(4293) <= a and not b;
    layer0_outputs(4294) <= not a or b;
    layer0_outputs(4295) <= '0';
    layer0_outputs(4296) <= not (a xor b);
    layer0_outputs(4297) <= a and not b;
    layer0_outputs(4298) <= '0';
    layer0_outputs(4299) <= not b or a;
    layer0_outputs(4300) <= not (a and b);
    layer0_outputs(4301) <= a or b;
    layer0_outputs(4302) <= not a;
    layer0_outputs(4303) <= a and b;
    layer0_outputs(4304) <= not a or b;
    layer0_outputs(4305) <= not (a and b);
    layer0_outputs(4306) <= b;
    layer0_outputs(4307) <= a;
    layer0_outputs(4308) <= b;
    layer0_outputs(4309) <= not b;
    layer0_outputs(4310) <= not b or a;
    layer0_outputs(4311) <= a xor b;
    layer0_outputs(4312) <= not b;
    layer0_outputs(4313) <= not (a or b);
    layer0_outputs(4314) <= b;
    layer0_outputs(4315) <= a or b;
    layer0_outputs(4316) <= a or b;
    layer0_outputs(4317) <= not (a or b);
    layer0_outputs(4318) <= a or b;
    layer0_outputs(4319) <= '1';
    layer0_outputs(4320) <= not a;
    layer0_outputs(4321) <= '0';
    layer0_outputs(4322) <= a or b;
    layer0_outputs(4323) <= a and b;
    layer0_outputs(4324) <= '1';
    layer0_outputs(4325) <= not b;
    layer0_outputs(4326) <= not (a xor b);
    layer0_outputs(4327) <= a or b;
    layer0_outputs(4328) <= b;
    layer0_outputs(4329) <= a or b;
    layer0_outputs(4330) <= '1';
    layer0_outputs(4331) <= not (a or b);
    layer0_outputs(4332) <= a and not b;
    layer0_outputs(4333) <= b and not a;
    layer0_outputs(4334) <= not (a or b);
    layer0_outputs(4335) <= a and b;
    layer0_outputs(4336) <= not (a or b);
    layer0_outputs(4337) <= b and not a;
    layer0_outputs(4338) <= not (a or b);
    layer0_outputs(4339) <= not a;
    layer0_outputs(4340) <= a;
    layer0_outputs(4341) <= a and not b;
    layer0_outputs(4342) <= not a or b;
    layer0_outputs(4343) <= not (a and b);
    layer0_outputs(4344) <= b;
    layer0_outputs(4345) <= '0';
    layer0_outputs(4346) <= not b or a;
    layer0_outputs(4347) <= not (a or b);
    layer0_outputs(4348) <= not (a and b);
    layer0_outputs(4349) <= a;
    layer0_outputs(4350) <= '1';
    layer0_outputs(4351) <= a xor b;
    layer0_outputs(4352) <= not (a and b);
    layer0_outputs(4353) <= not (a and b);
    layer0_outputs(4354) <= '1';
    layer0_outputs(4355) <= not b or a;
    layer0_outputs(4356) <= not b;
    layer0_outputs(4357) <= a and b;
    layer0_outputs(4358) <= not (a or b);
    layer0_outputs(4359) <= a and b;
    layer0_outputs(4360) <= a xor b;
    layer0_outputs(4361) <= not (a or b);
    layer0_outputs(4362) <= not b;
    layer0_outputs(4363) <= a and not b;
    layer0_outputs(4364) <= '0';
    layer0_outputs(4365) <= '1';
    layer0_outputs(4366) <= not b or a;
    layer0_outputs(4367) <= not a or b;
    layer0_outputs(4368) <= not (a and b);
    layer0_outputs(4369) <= a and not b;
    layer0_outputs(4370) <= not b or a;
    layer0_outputs(4371) <= b;
    layer0_outputs(4372) <= b;
    layer0_outputs(4373) <= not (a or b);
    layer0_outputs(4374) <= b and not a;
    layer0_outputs(4375) <= '1';
    layer0_outputs(4376) <= '0';
    layer0_outputs(4377) <= '0';
    layer0_outputs(4378) <= a and b;
    layer0_outputs(4379) <= not (a and b);
    layer0_outputs(4380) <= not a or b;
    layer0_outputs(4381) <= not a or b;
    layer0_outputs(4382) <= not (a xor b);
    layer0_outputs(4383) <= a;
    layer0_outputs(4384) <= not a or b;
    layer0_outputs(4385) <= not (a or b);
    layer0_outputs(4386) <= '0';
    layer0_outputs(4387) <= not (a or b);
    layer0_outputs(4388) <= a or b;
    layer0_outputs(4389) <= b and not a;
    layer0_outputs(4390) <= '0';
    layer0_outputs(4391) <= not (a or b);
    layer0_outputs(4392) <= a or b;
    layer0_outputs(4393) <= '0';
    layer0_outputs(4394) <= a or b;
    layer0_outputs(4395) <= not b or a;
    layer0_outputs(4396) <= '0';
    layer0_outputs(4397) <= b;
    layer0_outputs(4398) <= not (a or b);
    layer0_outputs(4399) <= a or b;
    layer0_outputs(4400) <= b;
    layer0_outputs(4401) <= not a;
    layer0_outputs(4402) <= not b or a;
    layer0_outputs(4403) <= a;
    layer0_outputs(4404) <= b and not a;
    layer0_outputs(4405) <= not a;
    layer0_outputs(4406) <= not a;
    layer0_outputs(4407) <= '1';
    layer0_outputs(4408) <= a xor b;
    layer0_outputs(4409) <= not a;
    layer0_outputs(4410) <= '0';
    layer0_outputs(4411) <= a and not b;
    layer0_outputs(4412) <= '0';
    layer0_outputs(4413) <= '0';
    layer0_outputs(4414) <= a and b;
    layer0_outputs(4415) <= not (a and b);
    layer0_outputs(4416) <= not a;
    layer0_outputs(4417) <= '0';
    layer0_outputs(4418) <= b;
    layer0_outputs(4419) <= not a or b;
    layer0_outputs(4420) <= '0';
    layer0_outputs(4421) <= '0';
    layer0_outputs(4422) <= b;
    layer0_outputs(4423) <= b and not a;
    layer0_outputs(4424) <= '0';
    layer0_outputs(4425) <= b and not a;
    layer0_outputs(4426) <= b;
    layer0_outputs(4427) <= b and not a;
    layer0_outputs(4428) <= b and not a;
    layer0_outputs(4429) <= not (a or b);
    layer0_outputs(4430) <= a;
    layer0_outputs(4431) <= not (a or b);
    layer0_outputs(4432) <= not a or b;
    layer0_outputs(4433) <= not (a xor b);
    layer0_outputs(4434) <= not a;
    layer0_outputs(4435) <= b and not a;
    layer0_outputs(4436) <= not (a and b);
    layer0_outputs(4437) <= not a or b;
    layer0_outputs(4438) <= '1';
    layer0_outputs(4439) <= not b or a;
    layer0_outputs(4440) <= not (a and b);
    layer0_outputs(4441) <= a;
    layer0_outputs(4442) <= not b or a;
    layer0_outputs(4443) <= not a or b;
    layer0_outputs(4444) <= a or b;
    layer0_outputs(4445) <= a;
    layer0_outputs(4446) <= a and not b;
    layer0_outputs(4447) <= a and not b;
    layer0_outputs(4448) <= not a;
    layer0_outputs(4449) <= not (a or b);
    layer0_outputs(4450) <= a and not b;
    layer0_outputs(4451) <= not (a and b);
    layer0_outputs(4452) <= a;
    layer0_outputs(4453) <= not b;
    layer0_outputs(4454) <= not a;
    layer0_outputs(4455) <= '1';
    layer0_outputs(4456) <= '1';
    layer0_outputs(4457) <= not a;
    layer0_outputs(4458) <= '0';
    layer0_outputs(4459) <= a xor b;
    layer0_outputs(4460) <= a or b;
    layer0_outputs(4461) <= not (a or b);
    layer0_outputs(4462) <= a and not b;
    layer0_outputs(4463) <= not a or b;
    layer0_outputs(4464) <= not (a or b);
    layer0_outputs(4465) <= not (a xor b);
    layer0_outputs(4466) <= not a;
    layer0_outputs(4467) <= '1';
    layer0_outputs(4468) <= a xor b;
    layer0_outputs(4469) <= not (a or b);
    layer0_outputs(4470) <= '1';
    layer0_outputs(4471) <= not a or b;
    layer0_outputs(4472) <= not (a xor b);
    layer0_outputs(4473) <= not a or b;
    layer0_outputs(4474) <= not (a or b);
    layer0_outputs(4475) <= not b or a;
    layer0_outputs(4476) <= not a;
    layer0_outputs(4477) <= a or b;
    layer0_outputs(4478) <= not b;
    layer0_outputs(4479) <= not a;
    layer0_outputs(4480) <= '1';
    layer0_outputs(4481) <= '1';
    layer0_outputs(4482) <= '1';
    layer0_outputs(4483) <= not b;
    layer0_outputs(4484) <= not (a and b);
    layer0_outputs(4485) <= a;
    layer0_outputs(4486) <= b;
    layer0_outputs(4487) <= not (a or b);
    layer0_outputs(4488) <= not b or a;
    layer0_outputs(4489) <= a xor b;
    layer0_outputs(4490) <= b and not a;
    layer0_outputs(4491) <= a and b;
    layer0_outputs(4492) <= a and not b;
    layer0_outputs(4493) <= not b or a;
    layer0_outputs(4494) <= a and b;
    layer0_outputs(4495) <= a and b;
    layer0_outputs(4496) <= a xor b;
    layer0_outputs(4497) <= a and b;
    layer0_outputs(4498) <= '0';
    layer0_outputs(4499) <= not a;
    layer0_outputs(4500) <= b;
    layer0_outputs(4501) <= not b;
    layer0_outputs(4502) <= not a or b;
    layer0_outputs(4503) <= not b or a;
    layer0_outputs(4504) <= a xor b;
    layer0_outputs(4505) <= b;
    layer0_outputs(4506) <= not b;
    layer0_outputs(4507) <= a;
    layer0_outputs(4508) <= a and b;
    layer0_outputs(4509) <= a;
    layer0_outputs(4510) <= '0';
    layer0_outputs(4511) <= a and not b;
    layer0_outputs(4512) <= '1';
    layer0_outputs(4513) <= a or b;
    layer0_outputs(4514) <= a or b;
    layer0_outputs(4515) <= '0';
    layer0_outputs(4516) <= b;
    layer0_outputs(4517) <= not (a or b);
    layer0_outputs(4518) <= not b;
    layer0_outputs(4519) <= not b;
    layer0_outputs(4520) <= not b or a;
    layer0_outputs(4521) <= a;
    layer0_outputs(4522) <= a and b;
    layer0_outputs(4523) <= b;
    layer0_outputs(4524) <= a xor b;
    layer0_outputs(4525) <= not (a and b);
    layer0_outputs(4526) <= a;
    layer0_outputs(4527) <= '0';
    layer0_outputs(4528) <= not a or b;
    layer0_outputs(4529) <= not (a xor b);
    layer0_outputs(4530) <= not a or b;
    layer0_outputs(4531) <= not a;
    layer0_outputs(4532) <= not (a and b);
    layer0_outputs(4533) <= b and not a;
    layer0_outputs(4534) <= '1';
    layer0_outputs(4535) <= not a;
    layer0_outputs(4536) <= a and b;
    layer0_outputs(4537) <= not a or b;
    layer0_outputs(4538) <= b and not a;
    layer0_outputs(4539) <= '1';
    layer0_outputs(4540) <= a;
    layer0_outputs(4541) <= '1';
    layer0_outputs(4542) <= a;
    layer0_outputs(4543) <= a and not b;
    layer0_outputs(4544) <= a and not b;
    layer0_outputs(4545) <= not b;
    layer0_outputs(4546) <= a xor b;
    layer0_outputs(4547) <= '1';
    layer0_outputs(4548) <= b;
    layer0_outputs(4549) <= b;
    layer0_outputs(4550) <= b;
    layer0_outputs(4551) <= not (a or b);
    layer0_outputs(4552) <= a and b;
    layer0_outputs(4553) <= not b or a;
    layer0_outputs(4554) <= not a;
    layer0_outputs(4555) <= not b;
    layer0_outputs(4556) <= b and not a;
    layer0_outputs(4557) <= not a or b;
    layer0_outputs(4558) <= a xor b;
    layer0_outputs(4559) <= b and not a;
    layer0_outputs(4560) <= not (a or b);
    layer0_outputs(4561) <= b;
    layer0_outputs(4562) <= not b;
    layer0_outputs(4563) <= a and b;
    layer0_outputs(4564) <= not b;
    layer0_outputs(4565) <= a and b;
    layer0_outputs(4566) <= not (a xor b);
    layer0_outputs(4567) <= '1';
    layer0_outputs(4568) <= a and b;
    layer0_outputs(4569) <= '1';
    layer0_outputs(4570) <= not a;
    layer0_outputs(4571) <= '0';
    layer0_outputs(4572) <= not (a and b);
    layer0_outputs(4573) <= '0';
    layer0_outputs(4574) <= a and b;
    layer0_outputs(4575) <= b and not a;
    layer0_outputs(4576) <= not b;
    layer0_outputs(4577) <= a and b;
    layer0_outputs(4578) <= not b;
    layer0_outputs(4579) <= a and b;
    layer0_outputs(4580) <= not (a and b);
    layer0_outputs(4581) <= '1';
    layer0_outputs(4582) <= b;
    layer0_outputs(4583) <= not (a or b);
    layer0_outputs(4584) <= a;
    layer0_outputs(4585) <= b;
    layer0_outputs(4586) <= a or b;
    layer0_outputs(4587) <= '1';
    layer0_outputs(4588) <= a and b;
    layer0_outputs(4589) <= not a or b;
    layer0_outputs(4590) <= a and not b;
    layer0_outputs(4591) <= a and b;
    layer0_outputs(4592) <= not (a and b);
    layer0_outputs(4593) <= not a;
    layer0_outputs(4594) <= '1';
    layer0_outputs(4595) <= b;
    layer0_outputs(4596) <= not a or b;
    layer0_outputs(4597) <= b and not a;
    layer0_outputs(4598) <= a and b;
    layer0_outputs(4599) <= not b;
    layer0_outputs(4600) <= a or b;
    layer0_outputs(4601) <= b and not a;
    layer0_outputs(4602) <= a and b;
    layer0_outputs(4603) <= '1';
    layer0_outputs(4604) <= not (a or b);
    layer0_outputs(4605) <= '0';
    layer0_outputs(4606) <= a;
    layer0_outputs(4607) <= a;
    layer0_outputs(4608) <= a and b;
    layer0_outputs(4609) <= b and not a;
    layer0_outputs(4610) <= b;
    layer0_outputs(4611) <= not a;
    layer0_outputs(4612) <= a and not b;
    layer0_outputs(4613) <= not b;
    layer0_outputs(4614) <= a and b;
    layer0_outputs(4615) <= a and not b;
    layer0_outputs(4616) <= a and not b;
    layer0_outputs(4617) <= a or b;
    layer0_outputs(4618) <= a;
    layer0_outputs(4619) <= not b or a;
    layer0_outputs(4620) <= not a;
    layer0_outputs(4621) <= a xor b;
    layer0_outputs(4622) <= a;
    layer0_outputs(4623) <= a xor b;
    layer0_outputs(4624) <= a or b;
    layer0_outputs(4625) <= a or b;
    layer0_outputs(4626) <= b;
    layer0_outputs(4627) <= not a;
    layer0_outputs(4628) <= a and b;
    layer0_outputs(4629) <= not (a xor b);
    layer0_outputs(4630) <= a or b;
    layer0_outputs(4631) <= a or b;
    layer0_outputs(4632) <= a;
    layer0_outputs(4633) <= a and not b;
    layer0_outputs(4634) <= not a or b;
    layer0_outputs(4635) <= a xor b;
    layer0_outputs(4636) <= a;
    layer0_outputs(4637) <= not a;
    layer0_outputs(4638) <= b;
    layer0_outputs(4639) <= '1';
    layer0_outputs(4640) <= not (a and b);
    layer0_outputs(4641) <= b;
    layer0_outputs(4642) <= b and not a;
    layer0_outputs(4643) <= '0';
    layer0_outputs(4644) <= a and not b;
    layer0_outputs(4645) <= a;
    layer0_outputs(4646) <= a and b;
    layer0_outputs(4647) <= '1';
    layer0_outputs(4648) <= not b;
    layer0_outputs(4649) <= a and not b;
    layer0_outputs(4650) <= a and b;
    layer0_outputs(4651) <= b and not a;
    layer0_outputs(4652) <= not a;
    layer0_outputs(4653) <= not b or a;
    layer0_outputs(4654) <= '0';
    layer0_outputs(4655) <= not (a or b);
    layer0_outputs(4656) <= a or b;
    layer0_outputs(4657) <= not (a xor b);
    layer0_outputs(4658) <= not a;
    layer0_outputs(4659) <= not (a and b);
    layer0_outputs(4660) <= a or b;
    layer0_outputs(4661) <= not (a or b);
    layer0_outputs(4662) <= not b;
    layer0_outputs(4663) <= not b;
    layer0_outputs(4664) <= a xor b;
    layer0_outputs(4665) <= not b or a;
    layer0_outputs(4666) <= a or b;
    layer0_outputs(4667) <= not a;
    layer0_outputs(4668) <= a xor b;
    layer0_outputs(4669) <= b;
    layer0_outputs(4670) <= a and not b;
    layer0_outputs(4671) <= b;
    layer0_outputs(4672) <= a and not b;
    layer0_outputs(4673) <= not a;
    layer0_outputs(4674) <= a;
    layer0_outputs(4675) <= not (a or b);
    layer0_outputs(4676) <= not (a and b);
    layer0_outputs(4677) <= not b or a;
    layer0_outputs(4678) <= not b;
    layer0_outputs(4679) <= b;
    layer0_outputs(4680) <= a and b;
    layer0_outputs(4681) <= not b;
    layer0_outputs(4682) <= '1';
    layer0_outputs(4683) <= a and not b;
    layer0_outputs(4684) <= b;
    layer0_outputs(4685) <= not (a or b);
    layer0_outputs(4686) <= a and b;
    layer0_outputs(4687) <= b;
    layer0_outputs(4688) <= not (a and b);
    layer0_outputs(4689) <= not b;
    layer0_outputs(4690) <= '0';
    layer0_outputs(4691) <= not b;
    layer0_outputs(4692) <= not b;
    layer0_outputs(4693) <= not (a or b);
    layer0_outputs(4694) <= a or b;
    layer0_outputs(4695) <= '0';
    layer0_outputs(4696) <= '1';
    layer0_outputs(4697) <= not (a and b);
    layer0_outputs(4698) <= a and b;
    layer0_outputs(4699) <= '1';
    layer0_outputs(4700) <= not b;
    layer0_outputs(4701) <= a and b;
    layer0_outputs(4702) <= b and not a;
    layer0_outputs(4703) <= not a;
    layer0_outputs(4704) <= a;
    layer0_outputs(4705) <= not b;
    layer0_outputs(4706) <= a or b;
    layer0_outputs(4707) <= a and not b;
    layer0_outputs(4708) <= not a;
    layer0_outputs(4709) <= a;
    layer0_outputs(4710) <= '1';
    layer0_outputs(4711) <= b and not a;
    layer0_outputs(4712) <= a or b;
    layer0_outputs(4713) <= b and not a;
    layer0_outputs(4714) <= '0';
    layer0_outputs(4715) <= not b or a;
    layer0_outputs(4716) <= not (a or b);
    layer0_outputs(4717) <= not b or a;
    layer0_outputs(4718) <= not b or a;
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= b;
    layer0_outputs(4721) <= not b;
    layer0_outputs(4722) <= not a or b;
    layer0_outputs(4723) <= a or b;
    layer0_outputs(4724) <= a and b;
    layer0_outputs(4725) <= not b;
    layer0_outputs(4726) <= a;
    layer0_outputs(4727) <= not (a or b);
    layer0_outputs(4728) <= b;
    layer0_outputs(4729) <= '0';
    layer0_outputs(4730) <= not (a or b);
    layer0_outputs(4731) <= not b or a;
    layer0_outputs(4732) <= not b;
    layer0_outputs(4733) <= a;
    layer0_outputs(4734) <= not b;
    layer0_outputs(4735) <= a and b;
    layer0_outputs(4736) <= a or b;
    layer0_outputs(4737) <= a;
    layer0_outputs(4738) <= a or b;
    layer0_outputs(4739) <= a;
    layer0_outputs(4740) <= b;
    layer0_outputs(4741) <= b and not a;
    layer0_outputs(4742) <= a;
    layer0_outputs(4743) <= '1';
    layer0_outputs(4744) <= b;
    layer0_outputs(4745) <= b and not a;
    layer0_outputs(4746) <= a xor b;
    layer0_outputs(4747) <= not (a xor b);
    layer0_outputs(4748) <= '0';
    layer0_outputs(4749) <= not a;
    layer0_outputs(4750) <= not (a xor b);
    layer0_outputs(4751) <= a and not b;
    layer0_outputs(4752) <= a;
    layer0_outputs(4753) <= a or b;
    layer0_outputs(4754) <= a xor b;
    layer0_outputs(4755) <= a;
    layer0_outputs(4756) <= a;
    layer0_outputs(4757) <= not a;
    layer0_outputs(4758) <= '0';
    layer0_outputs(4759) <= a and not b;
    layer0_outputs(4760) <= b and not a;
    layer0_outputs(4761) <= not a;
    layer0_outputs(4762) <= a and not b;
    layer0_outputs(4763) <= not b or a;
    layer0_outputs(4764) <= a;
    layer0_outputs(4765) <= not (a xor b);
    layer0_outputs(4766) <= not (a and b);
    layer0_outputs(4767) <= a and not b;
    layer0_outputs(4768) <= a and b;
    layer0_outputs(4769) <= '0';
    layer0_outputs(4770) <= not a;
    layer0_outputs(4771) <= '0';
    layer0_outputs(4772) <= not (a xor b);
    layer0_outputs(4773) <= not (a xor b);
    layer0_outputs(4774) <= not (a or b);
    layer0_outputs(4775) <= not b;
    layer0_outputs(4776) <= b and not a;
    layer0_outputs(4777) <= '1';
    layer0_outputs(4778) <= not b;
    layer0_outputs(4779) <= not (a or b);
    layer0_outputs(4780) <= not a;
    layer0_outputs(4781) <= not b;
    layer0_outputs(4782) <= '0';
    layer0_outputs(4783) <= a and b;
    layer0_outputs(4784) <= b and not a;
    layer0_outputs(4785) <= not b or a;
    layer0_outputs(4786) <= b;
    layer0_outputs(4787) <= not a;
    layer0_outputs(4788) <= a and b;
    layer0_outputs(4789) <= not a;
    layer0_outputs(4790) <= not b or a;
    layer0_outputs(4791) <= a or b;
    layer0_outputs(4792) <= '0';
    layer0_outputs(4793) <= not (a or b);
    layer0_outputs(4794) <= b;
    layer0_outputs(4795) <= b;
    layer0_outputs(4796) <= '0';
    layer0_outputs(4797) <= '1';
    layer0_outputs(4798) <= not a;
    layer0_outputs(4799) <= not (a xor b);
    layer0_outputs(4800) <= '1';
    layer0_outputs(4801) <= a xor b;
    layer0_outputs(4802) <= not (a and b);
    layer0_outputs(4803) <= '0';
    layer0_outputs(4804) <= b;
    layer0_outputs(4805) <= not b or a;
    layer0_outputs(4806) <= not (a and b);
    layer0_outputs(4807) <= not (a and b);
    layer0_outputs(4808) <= a;
    layer0_outputs(4809) <= not a or b;
    layer0_outputs(4810) <= not b or a;
    layer0_outputs(4811) <= b and not a;
    layer0_outputs(4812) <= not (a or b);
    layer0_outputs(4813) <= not b or a;
    layer0_outputs(4814) <= not a;
    layer0_outputs(4815) <= not b or a;
    layer0_outputs(4816) <= b;
    layer0_outputs(4817) <= a and b;
    layer0_outputs(4818) <= a;
    layer0_outputs(4819) <= a and not b;
    layer0_outputs(4820) <= not a;
    layer0_outputs(4821) <= not b;
    layer0_outputs(4822) <= b and not a;
    layer0_outputs(4823) <= a;
    layer0_outputs(4824) <= '1';
    layer0_outputs(4825) <= b;
    layer0_outputs(4826) <= b and not a;
    layer0_outputs(4827) <= not (a and b);
    layer0_outputs(4828) <= b;
    layer0_outputs(4829) <= a and b;
    layer0_outputs(4830) <= not b;
    layer0_outputs(4831) <= a and b;
    layer0_outputs(4832) <= not b or a;
    layer0_outputs(4833) <= '0';
    layer0_outputs(4834) <= a or b;
    layer0_outputs(4835) <= not b or a;
    layer0_outputs(4836) <= a and not b;
    layer0_outputs(4837) <= not (a xor b);
    layer0_outputs(4838) <= a xor b;
    layer0_outputs(4839) <= b;
    layer0_outputs(4840) <= a or b;
    layer0_outputs(4841) <= '1';
    layer0_outputs(4842) <= b;
    layer0_outputs(4843) <= a and not b;
    layer0_outputs(4844) <= b;
    layer0_outputs(4845) <= not b;
    layer0_outputs(4846) <= not (a xor b);
    layer0_outputs(4847) <= not b;
    layer0_outputs(4848) <= not a;
    layer0_outputs(4849) <= not b or a;
    layer0_outputs(4850) <= not a;
    layer0_outputs(4851) <= '1';
    layer0_outputs(4852) <= a;
    layer0_outputs(4853) <= b;
    layer0_outputs(4854) <= a and b;
    layer0_outputs(4855) <= not a or b;
    layer0_outputs(4856) <= not (a and b);
    layer0_outputs(4857) <= not b or a;
    layer0_outputs(4858) <= not (a and b);
    layer0_outputs(4859) <= a;
    layer0_outputs(4860) <= not (a xor b);
    layer0_outputs(4861) <= a or b;
    layer0_outputs(4862) <= a xor b;
    layer0_outputs(4863) <= not (a and b);
    layer0_outputs(4864) <= a or b;
    layer0_outputs(4865) <= not a or b;
    layer0_outputs(4866) <= not b;
    layer0_outputs(4867) <= '1';
    layer0_outputs(4868) <= not a or b;
    layer0_outputs(4869) <= not (a or b);
    layer0_outputs(4870) <= '0';
    layer0_outputs(4871) <= not a;
    layer0_outputs(4872) <= '0';
    layer0_outputs(4873) <= b and not a;
    layer0_outputs(4874) <= a;
    layer0_outputs(4875) <= not b or a;
    layer0_outputs(4876) <= b and not a;
    layer0_outputs(4877) <= a and not b;
    layer0_outputs(4878) <= '0';
    layer0_outputs(4879) <= a and not b;
    layer0_outputs(4880) <= a;
    layer0_outputs(4881) <= not b;
    layer0_outputs(4882) <= not (a and b);
    layer0_outputs(4883) <= not a or b;
    layer0_outputs(4884) <= a and not b;
    layer0_outputs(4885) <= '1';
    layer0_outputs(4886) <= '1';
    layer0_outputs(4887) <= '1';
    layer0_outputs(4888) <= not (a or b);
    layer0_outputs(4889) <= a xor b;
    layer0_outputs(4890) <= not b;
    layer0_outputs(4891) <= a and b;
    layer0_outputs(4892) <= b and not a;
    layer0_outputs(4893) <= a xor b;
    layer0_outputs(4894) <= a;
    layer0_outputs(4895) <= not a;
    layer0_outputs(4896) <= not b;
    layer0_outputs(4897) <= not (a and b);
    layer0_outputs(4898) <= b and not a;
    layer0_outputs(4899) <= '0';
    layer0_outputs(4900) <= not (a or b);
    layer0_outputs(4901) <= not (a and b);
    layer0_outputs(4902) <= not (a xor b);
    layer0_outputs(4903) <= a or b;
    layer0_outputs(4904) <= '1';
    layer0_outputs(4905) <= not (a or b);
    layer0_outputs(4906) <= a xor b;
    layer0_outputs(4907) <= '0';
    layer0_outputs(4908) <= a and not b;
    layer0_outputs(4909) <= a or b;
    layer0_outputs(4910) <= '0';
    layer0_outputs(4911) <= a;
    layer0_outputs(4912) <= not (a and b);
    layer0_outputs(4913) <= '1';
    layer0_outputs(4914) <= '1';
    layer0_outputs(4915) <= not (a xor b);
    layer0_outputs(4916) <= a;
    layer0_outputs(4917) <= not (a or b);
    layer0_outputs(4918) <= not (a and b);
    layer0_outputs(4919) <= not (a or b);
    layer0_outputs(4920) <= not b or a;
    layer0_outputs(4921) <= not (a xor b);
    layer0_outputs(4922) <= '1';
    layer0_outputs(4923) <= not a or b;
    layer0_outputs(4924) <= not (a xor b);
    layer0_outputs(4925) <= '1';
    layer0_outputs(4926) <= not a or b;
    layer0_outputs(4927) <= a and b;
    layer0_outputs(4928) <= a;
    layer0_outputs(4929) <= not b;
    layer0_outputs(4930) <= a xor b;
    layer0_outputs(4931) <= not b or a;
    layer0_outputs(4932) <= '1';
    layer0_outputs(4933) <= '0';
    layer0_outputs(4934) <= not (a and b);
    layer0_outputs(4935) <= a;
    layer0_outputs(4936) <= not (a and b);
    layer0_outputs(4937) <= '0';
    layer0_outputs(4938) <= not (a or b);
    layer0_outputs(4939) <= a xor b;
    layer0_outputs(4940) <= not (a and b);
    layer0_outputs(4941) <= a and not b;
    layer0_outputs(4942) <= b;
    layer0_outputs(4943) <= a and not b;
    layer0_outputs(4944) <= b;
    layer0_outputs(4945) <= a or b;
    layer0_outputs(4946) <= not b;
    layer0_outputs(4947) <= not b;
    layer0_outputs(4948) <= b and not a;
    layer0_outputs(4949) <= a and not b;
    layer0_outputs(4950) <= not a;
    layer0_outputs(4951) <= b and not a;
    layer0_outputs(4952) <= not b or a;
    layer0_outputs(4953) <= a or b;
    layer0_outputs(4954) <= a and b;
    layer0_outputs(4955) <= not (a xor b);
    layer0_outputs(4956) <= a or b;
    layer0_outputs(4957) <= '1';
    layer0_outputs(4958) <= not b or a;
    layer0_outputs(4959) <= not b or a;
    layer0_outputs(4960) <= b;
    layer0_outputs(4961) <= not b or a;
    layer0_outputs(4962) <= not b;
    layer0_outputs(4963) <= not (a xor b);
    layer0_outputs(4964) <= not (a and b);
    layer0_outputs(4965) <= not a or b;
    layer0_outputs(4966) <= '0';
    layer0_outputs(4967) <= not a;
    layer0_outputs(4968) <= '1';
    layer0_outputs(4969) <= '0';
    layer0_outputs(4970) <= a xor b;
    layer0_outputs(4971) <= b and not a;
    layer0_outputs(4972) <= a xor b;
    layer0_outputs(4973) <= not a or b;
    layer0_outputs(4974) <= a and not b;
    layer0_outputs(4975) <= a and not b;
    layer0_outputs(4976) <= not (a xor b);
    layer0_outputs(4977) <= '1';
    layer0_outputs(4978) <= not b;
    layer0_outputs(4979) <= a xor b;
    layer0_outputs(4980) <= b and not a;
    layer0_outputs(4981) <= a or b;
    layer0_outputs(4982) <= not a or b;
    layer0_outputs(4983) <= a and b;
    layer0_outputs(4984) <= a and not b;
    layer0_outputs(4985) <= a and not b;
    layer0_outputs(4986) <= '1';
    layer0_outputs(4987) <= a and not b;
    layer0_outputs(4988) <= not (a and b);
    layer0_outputs(4989) <= a and b;
    layer0_outputs(4990) <= not b or a;
    layer0_outputs(4991) <= '1';
    layer0_outputs(4992) <= a xor b;
    layer0_outputs(4993) <= b;
    layer0_outputs(4994) <= not a or b;
    layer0_outputs(4995) <= b and not a;
    layer0_outputs(4996) <= not (a or b);
    layer0_outputs(4997) <= not b or a;
    layer0_outputs(4998) <= not b;
    layer0_outputs(4999) <= not (a and b);
    layer0_outputs(5000) <= b;
    layer0_outputs(5001) <= not (a or b);
    layer0_outputs(5002) <= '1';
    layer0_outputs(5003) <= not (a and b);
    layer0_outputs(5004) <= b and not a;
    layer0_outputs(5005) <= not a or b;
    layer0_outputs(5006) <= '1';
    layer0_outputs(5007) <= not (a or b);
    layer0_outputs(5008) <= not (a and b);
    layer0_outputs(5009) <= not b;
    layer0_outputs(5010) <= '0';
    layer0_outputs(5011) <= not (a xor b);
    layer0_outputs(5012) <= not (a and b);
    layer0_outputs(5013) <= a;
    layer0_outputs(5014) <= a and b;
    layer0_outputs(5015) <= b;
    layer0_outputs(5016) <= not a;
    layer0_outputs(5017) <= '1';
    layer0_outputs(5018) <= a xor b;
    layer0_outputs(5019) <= a;
    layer0_outputs(5020) <= '1';
    layer0_outputs(5021) <= '1';
    layer0_outputs(5022) <= not a;
    layer0_outputs(5023) <= not b;
    layer0_outputs(5024) <= a;
    layer0_outputs(5025) <= a or b;
    layer0_outputs(5026) <= b and not a;
    layer0_outputs(5027) <= '1';
    layer0_outputs(5028) <= not b;
    layer0_outputs(5029) <= b and not a;
    layer0_outputs(5030) <= a;
    layer0_outputs(5031) <= '1';
    layer0_outputs(5032) <= '1';
    layer0_outputs(5033) <= b and not a;
    layer0_outputs(5034) <= '0';
    layer0_outputs(5035) <= not a or b;
    layer0_outputs(5036) <= not (a and b);
    layer0_outputs(5037) <= a;
    layer0_outputs(5038) <= not b or a;
    layer0_outputs(5039) <= not a or b;
    layer0_outputs(5040) <= '0';
    layer0_outputs(5041) <= a and not b;
    layer0_outputs(5042) <= '1';
    layer0_outputs(5043) <= b;
    layer0_outputs(5044) <= '0';
    layer0_outputs(5045) <= not a;
    layer0_outputs(5046) <= a and not b;
    layer0_outputs(5047) <= not b or a;
    layer0_outputs(5048) <= not (a xor b);
    layer0_outputs(5049) <= a xor b;
    layer0_outputs(5050) <= a and not b;
    layer0_outputs(5051) <= a or b;
    layer0_outputs(5052) <= a;
    layer0_outputs(5053) <= b;
    layer0_outputs(5054) <= not (a or b);
    layer0_outputs(5055) <= a;
    layer0_outputs(5056) <= a and b;
    layer0_outputs(5057) <= not a or b;
    layer0_outputs(5058) <= not (a or b);
    layer0_outputs(5059) <= b and not a;
    layer0_outputs(5060) <= a;
    layer0_outputs(5061) <= '0';
    layer0_outputs(5062) <= '1';
    layer0_outputs(5063) <= a and not b;
    layer0_outputs(5064) <= a and not b;
    layer0_outputs(5065) <= a or b;
    layer0_outputs(5066) <= not b;
    layer0_outputs(5067) <= b and not a;
    layer0_outputs(5068) <= a and not b;
    layer0_outputs(5069) <= not a;
    layer0_outputs(5070) <= not (a xor b);
    layer0_outputs(5071) <= b;
    layer0_outputs(5072) <= not (a xor b);
    layer0_outputs(5073) <= a xor b;
    layer0_outputs(5074) <= a xor b;
    layer0_outputs(5075) <= not a;
    layer0_outputs(5076) <= not b;
    layer0_outputs(5077) <= a;
    layer0_outputs(5078) <= a;
    layer0_outputs(5079) <= a;
    layer0_outputs(5080) <= not a;
    layer0_outputs(5081) <= '1';
    layer0_outputs(5082) <= b and not a;
    layer0_outputs(5083) <= not (a or b);
    layer0_outputs(5084) <= a and b;
    layer0_outputs(5085) <= not a or b;
    layer0_outputs(5086) <= b and not a;
    layer0_outputs(5087) <= not (a and b);
    layer0_outputs(5088) <= a and b;
    layer0_outputs(5089) <= a and not b;
    layer0_outputs(5090) <= a or b;
    layer0_outputs(5091) <= a xor b;
    layer0_outputs(5092) <= b and not a;
    layer0_outputs(5093) <= not a or b;
    layer0_outputs(5094) <= not (a xor b);
    layer0_outputs(5095) <= '0';
    layer0_outputs(5096) <= b and not a;
    layer0_outputs(5097) <= '0';
    layer0_outputs(5098) <= '0';
    layer0_outputs(5099) <= not a or b;
    layer0_outputs(5100) <= '1';
    layer0_outputs(5101) <= not (a xor b);
    layer0_outputs(5102) <= not (a or b);
    layer0_outputs(5103) <= '0';
    layer0_outputs(5104) <= not (a xor b);
    layer0_outputs(5105) <= a and not b;
    layer0_outputs(5106) <= not a;
    layer0_outputs(5107) <= a or b;
    layer0_outputs(5108) <= a or b;
    layer0_outputs(5109) <= '0';
    layer0_outputs(5110) <= a and not b;
    layer0_outputs(5111) <= not (a or b);
    layer0_outputs(5112) <= '0';
    layer0_outputs(5113) <= '1';
    layer0_outputs(5114) <= not a or b;
    layer0_outputs(5115) <= a xor b;
    layer0_outputs(5116) <= a;
    layer0_outputs(5117) <= a and not b;
    layer0_outputs(5118) <= not a or b;
    layer0_outputs(5119) <= a and b;
    layer0_outputs(5120) <= a xor b;
    layer0_outputs(5121) <= not (a or b);
    layer0_outputs(5122) <= a xor b;
    layer0_outputs(5123) <= not a or b;
    layer0_outputs(5124) <= not b;
    layer0_outputs(5125) <= not b or a;
    layer0_outputs(5126) <= not (a and b);
    layer0_outputs(5127) <= not (a xor b);
    layer0_outputs(5128) <= '0';
    layer0_outputs(5129) <= not b or a;
    layer0_outputs(5130) <= not b;
    layer0_outputs(5131) <= '1';
    layer0_outputs(5132) <= b;
    layer0_outputs(5133) <= '1';
    layer0_outputs(5134) <= '1';
    layer0_outputs(5135) <= not b or a;
    layer0_outputs(5136) <= b;
    layer0_outputs(5137) <= a and not b;
    layer0_outputs(5138) <= not b;
    layer0_outputs(5139) <= not a or b;
    layer0_outputs(5140) <= not b;
    layer0_outputs(5141) <= not b;
    layer0_outputs(5142) <= '0';
    layer0_outputs(5143) <= not a;
    layer0_outputs(5144) <= not b;
    layer0_outputs(5145) <= not (a or b);
    layer0_outputs(5146) <= '1';
    layer0_outputs(5147) <= a;
    layer0_outputs(5148) <= a or b;
    layer0_outputs(5149) <= not (a and b);
    layer0_outputs(5150) <= '0';
    layer0_outputs(5151) <= b;
    layer0_outputs(5152) <= a or b;
    layer0_outputs(5153) <= a and not b;
    layer0_outputs(5154) <= b and not a;
    layer0_outputs(5155) <= not b or a;
    layer0_outputs(5156) <= not b;
    layer0_outputs(5157) <= a or b;
    layer0_outputs(5158) <= a and b;
    layer0_outputs(5159) <= a;
    layer0_outputs(5160) <= not b;
    layer0_outputs(5161) <= not b;
    layer0_outputs(5162) <= not (a or b);
    layer0_outputs(5163) <= b and not a;
    layer0_outputs(5164) <= not (a or b);
    layer0_outputs(5165) <= b and not a;
    layer0_outputs(5166) <= not a or b;
    layer0_outputs(5167) <= b and not a;
    layer0_outputs(5168) <= b;
    layer0_outputs(5169) <= a and b;
    layer0_outputs(5170) <= not a or b;
    layer0_outputs(5171) <= a;
    layer0_outputs(5172) <= not b or a;
    layer0_outputs(5173) <= '0';
    layer0_outputs(5174) <= '0';
    layer0_outputs(5175) <= a xor b;
    layer0_outputs(5176) <= a;
    layer0_outputs(5177) <= b and not a;
    layer0_outputs(5178) <= not (a or b);
    layer0_outputs(5179) <= not (a and b);
    layer0_outputs(5180) <= not (a or b);
    layer0_outputs(5181) <= not (a xor b);
    layer0_outputs(5182) <= a xor b;
    layer0_outputs(5183) <= not (a or b);
    layer0_outputs(5184) <= a and b;
    layer0_outputs(5185) <= not a;
    layer0_outputs(5186) <= not a;
    layer0_outputs(5187) <= a or b;
    layer0_outputs(5188) <= a xor b;
    layer0_outputs(5189) <= not (a and b);
    layer0_outputs(5190) <= not b;
    layer0_outputs(5191) <= not b;
    layer0_outputs(5192) <= not b or a;
    layer0_outputs(5193) <= b;
    layer0_outputs(5194) <= not a;
    layer0_outputs(5195) <= not b;
    layer0_outputs(5196) <= not a;
    layer0_outputs(5197) <= '1';
    layer0_outputs(5198) <= a or b;
    layer0_outputs(5199) <= not a or b;
    layer0_outputs(5200) <= not a or b;
    layer0_outputs(5201) <= a or b;
    layer0_outputs(5202) <= b;
    layer0_outputs(5203) <= a;
    layer0_outputs(5204) <= a;
    layer0_outputs(5205) <= '0';
    layer0_outputs(5206) <= not a;
    layer0_outputs(5207) <= not (a or b);
    layer0_outputs(5208) <= b and not a;
    layer0_outputs(5209) <= a or b;
    layer0_outputs(5210) <= a or b;
    layer0_outputs(5211) <= not (a or b);
    layer0_outputs(5212) <= not b;
    layer0_outputs(5213) <= not (a or b);
    layer0_outputs(5214) <= not b;
    layer0_outputs(5215) <= b;
    layer0_outputs(5216) <= a xor b;
    layer0_outputs(5217) <= b and not a;
    layer0_outputs(5218) <= not a or b;
    layer0_outputs(5219) <= not (a and b);
    layer0_outputs(5220) <= not (a xor b);
    layer0_outputs(5221) <= not b;
    layer0_outputs(5222) <= not b;
    layer0_outputs(5223) <= a;
    layer0_outputs(5224) <= a and not b;
    layer0_outputs(5225) <= not b or a;
    layer0_outputs(5226) <= a;
    layer0_outputs(5227) <= not a;
    layer0_outputs(5228) <= a;
    layer0_outputs(5229) <= a and not b;
    layer0_outputs(5230) <= a;
    layer0_outputs(5231) <= not (a xor b);
    layer0_outputs(5232) <= not (a or b);
    layer0_outputs(5233) <= '0';
    layer0_outputs(5234) <= not (a or b);
    layer0_outputs(5235) <= a or b;
    layer0_outputs(5236) <= a and b;
    layer0_outputs(5237) <= a;
    layer0_outputs(5238) <= not a or b;
    layer0_outputs(5239) <= b;
    layer0_outputs(5240) <= '0';
    layer0_outputs(5241) <= not a;
    layer0_outputs(5242) <= b;
    layer0_outputs(5243) <= '1';
    layer0_outputs(5244) <= b and not a;
    layer0_outputs(5245) <= '0';
    layer0_outputs(5246) <= '0';
    layer0_outputs(5247) <= a xor b;
    layer0_outputs(5248) <= '1';
    layer0_outputs(5249) <= not (a or b);
    layer0_outputs(5250) <= '1';
    layer0_outputs(5251) <= a xor b;
    layer0_outputs(5252) <= a or b;
    layer0_outputs(5253) <= not a or b;
    layer0_outputs(5254) <= not a or b;
    layer0_outputs(5255) <= a xor b;
    layer0_outputs(5256) <= a and not b;
    layer0_outputs(5257) <= not (a or b);
    layer0_outputs(5258) <= not (a or b);
    layer0_outputs(5259) <= a and not b;
    layer0_outputs(5260) <= b;
    layer0_outputs(5261) <= not a or b;
    layer0_outputs(5262) <= a or b;
    layer0_outputs(5263) <= not a or b;
    layer0_outputs(5264) <= b and not a;
    layer0_outputs(5265) <= a or b;
    layer0_outputs(5266) <= a or b;
    layer0_outputs(5267) <= a or b;
    layer0_outputs(5268) <= b;
    layer0_outputs(5269) <= not a;
    layer0_outputs(5270) <= a and not b;
    layer0_outputs(5271) <= a and b;
    layer0_outputs(5272) <= a xor b;
    layer0_outputs(5273) <= not b;
    layer0_outputs(5274) <= b and not a;
    layer0_outputs(5275) <= a;
    layer0_outputs(5276) <= b;
    layer0_outputs(5277) <= not b;
    layer0_outputs(5278) <= a;
    layer0_outputs(5279) <= b and not a;
    layer0_outputs(5280) <= not b;
    layer0_outputs(5281) <= a and b;
    layer0_outputs(5282) <= a and not b;
    layer0_outputs(5283) <= not a;
    layer0_outputs(5284) <= not a or b;
    layer0_outputs(5285) <= '0';
    layer0_outputs(5286) <= '1';
    layer0_outputs(5287) <= a and not b;
    layer0_outputs(5288) <= '0';
    layer0_outputs(5289) <= a;
    layer0_outputs(5290) <= not b or a;
    layer0_outputs(5291) <= a;
    layer0_outputs(5292) <= a and not b;
    layer0_outputs(5293) <= a;
    layer0_outputs(5294) <= a or b;
    layer0_outputs(5295) <= not (a or b);
    layer0_outputs(5296) <= not (a and b);
    layer0_outputs(5297) <= not b;
    layer0_outputs(5298) <= not (a xor b);
    layer0_outputs(5299) <= a;
    layer0_outputs(5300) <= not (a xor b);
    layer0_outputs(5301) <= not b;
    layer0_outputs(5302) <= a or b;
    layer0_outputs(5303) <= not a or b;
    layer0_outputs(5304) <= a or b;
    layer0_outputs(5305) <= not (a xor b);
    layer0_outputs(5306) <= not (a xor b);
    layer0_outputs(5307) <= b;
    layer0_outputs(5308) <= a;
    layer0_outputs(5309) <= a and b;
    layer0_outputs(5310) <= not (a or b);
    layer0_outputs(5311) <= '1';
    layer0_outputs(5312) <= b;
    layer0_outputs(5313) <= a xor b;
    layer0_outputs(5314) <= not a;
    layer0_outputs(5315) <= a;
    layer0_outputs(5316) <= not b;
    layer0_outputs(5317) <= b;
    layer0_outputs(5318) <= '1';
    layer0_outputs(5319) <= '1';
    layer0_outputs(5320) <= not a;
    layer0_outputs(5321) <= a and b;
    layer0_outputs(5322) <= b;
    layer0_outputs(5323) <= b and not a;
    layer0_outputs(5324) <= '1';
    layer0_outputs(5325) <= a and b;
    layer0_outputs(5326) <= not b;
    layer0_outputs(5327) <= '1';
    layer0_outputs(5328) <= a and not b;
    layer0_outputs(5329) <= a and not b;
    layer0_outputs(5330) <= b;
    layer0_outputs(5331) <= b;
    layer0_outputs(5332) <= '0';
    layer0_outputs(5333) <= a and not b;
    layer0_outputs(5334) <= not b or a;
    layer0_outputs(5335) <= not a or b;
    layer0_outputs(5336) <= a and b;
    layer0_outputs(5337) <= not a or b;
    layer0_outputs(5338) <= not b;
    layer0_outputs(5339) <= not b or a;
    layer0_outputs(5340) <= a or b;
    layer0_outputs(5341) <= a xor b;
    layer0_outputs(5342) <= a;
    layer0_outputs(5343) <= not (a and b);
    layer0_outputs(5344) <= a xor b;
    layer0_outputs(5345) <= '1';
    layer0_outputs(5346) <= a and b;
    layer0_outputs(5347) <= not b;
    layer0_outputs(5348) <= not b or a;
    layer0_outputs(5349) <= b and not a;
    layer0_outputs(5350) <= a and b;
    layer0_outputs(5351) <= '1';
    layer0_outputs(5352) <= a or b;
    layer0_outputs(5353) <= a and not b;
    layer0_outputs(5354) <= not a;
    layer0_outputs(5355) <= a and b;
    layer0_outputs(5356) <= not b;
    layer0_outputs(5357) <= not (a or b);
    layer0_outputs(5358) <= not (a or b);
    layer0_outputs(5359) <= '1';
    layer0_outputs(5360) <= not b;
    layer0_outputs(5361) <= a or b;
    layer0_outputs(5362) <= a or b;
    layer0_outputs(5363) <= a and not b;
    layer0_outputs(5364) <= a or b;
    layer0_outputs(5365) <= a xor b;
    layer0_outputs(5366) <= not a;
    layer0_outputs(5367) <= not (a or b);
    layer0_outputs(5368) <= not a;
    layer0_outputs(5369) <= not a or b;
    layer0_outputs(5370) <= not a;
    layer0_outputs(5371) <= '0';
    layer0_outputs(5372) <= a;
    layer0_outputs(5373) <= not (a and b);
    layer0_outputs(5374) <= a or b;
    layer0_outputs(5375) <= a or b;
    layer0_outputs(5376) <= a xor b;
    layer0_outputs(5377) <= b;
    layer0_outputs(5378) <= b;
    layer0_outputs(5379) <= '0';
    layer0_outputs(5380) <= not (a and b);
    layer0_outputs(5381) <= not b or a;
    layer0_outputs(5382) <= not b;
    layer0_outputs(5383) <= not a or b;
    layer0_outputs(5384) <= b;
    layer0_outputs(5385) <= not (a and b);
    layer0_outputs(5386) <= not a or b;
    layer0_outputs(5387) <= not b or a;
    layer0_outputs(5388) <= not b or a;
    layer0_outputs(5389) <= not (a or b);
    layer0_outputs(5390) <= '1';
    layer0_outputs(5391) <= not (a and b);
    layer0_outputs(5392) <= not (a or b);
    layer0_outputs(5393) <= not a;
    layer0_outputs(5394) <= a or b;
    layer0_outputs(5395) <= '0';
    layer0_outputs(5396) <= a or b;
    layer0_outputs(5397) <= '0';
    layer0_outputs(5398) <= a and not b;
    layer0_outputs(5399) <= b;
    layer0_outputs(5400) <= not (a and b);
    layer0_outputs(5401) <= a xor b;
    layer0_outputs(5402) <= not b or a;
    layer0_outputs(5403) <= a and b;
    layer0_outputs(5404) <= b and not a;
    layer0_outputs(5405) <= a and not b;
    layer0_outputs(5406) <= a and not b;
    layer0_outputs(5407) <= not b;
    layer0_outputs(5408) <= not b;
    layer0_outputs(5409) <= a and not b;
    layer0_outputs(5410) <= a and not b;
    layer0_outputs(5411) <= not (a xor b);
    layer0_outputs(5412) <= a or b;
    layer0_outputs(5413) <= not a or b;
    layer0_outputs(5414) <= not a or b;
    layer0_outputs(5415) <= a and not b;
    layer0_outputs(5416) <= b;
    layer0_outputs(5417) <= '1';
    layer0_outputs(5418) <= '0';
    layer0_outputs(5419) <= not (a or b);
    layer0_outputs(5420) <= not b;
    layer0_outputs(5421) <= b and not a;
    layer0_outputs(5422) <= b and not a;
    layer0_outputs(5423) <= not b;
    layer0_outputs(5424) <= a or b;
    layer0_outputs(5425) <= not a;
    layer0_outputs(5426) <= not a;
    layer0_outputs(5427) <= '0';
    layer0_outputs(5428) <= not a;
    layer0_outputs(5429) <= a or b;
    layer0_outputs(5430) <= b and not a;
    layer0_outputs(5431) <= not b or a;
    layer0_outputs(5432) <= not (a xor b);
    layer0_outputs(5433) <= not a;
    layer0_outputs(5434) <= not b or a;
    layer0_outputs(5435) <= not b;
    layer0_outputs(5436) <= '0';
    layer0_outputs(5437) <= not a or b;
    layer0_outputs(5438) <= a;
    layer0_outputs(5439) <= not (a or b);
    layer0_outputs(5440) <= not b;
    layer0_outputs(5441) <= b and not a;
    layer0_outputs(5442) <= a or b;
    layer0_outputs(5443) <= a xor b;
    layer0_outputs(5444) <= not b or a;
    layer0_outputs(5445) <= '1';
    layer0_outputs(5446) <= not b;
    layer0_outputs(5447) <= a and b;
    layer0_outputs(5448) <= a xor b;
    layer0_outputs(5449) <= a or b;
    layer0_outputs(5450) <= a and not b;
    layer0_outputs(5451) <= not b;
    layer0_outputs(5452) <= a and b;
    layer0_outputs(5453) <= a;
    layer0_outputs(5454) <= a xor b;
    layer0_outputs(5455) <= b and not a;
    layer0_outputs(5456) <= '0';
    layer0_outputs(5457) <= a and not b;
    layer0_outputs(5458) <= not b;
    layer0_outputs(5459) <= not a or b;
    layer0_outputs(5460) <= a or b;
    layer0_outputs(5461) <= '0';
    layer0_outputs(5462) <= not (a and b);
    layer0_outputs(5463) <= '0';
    layer0_outputs(5464) <= not (a or b);
    layer0_outputs(5465) <= not (a xor b);
    layer0_outputs(5466) <= not a or b;
    layer0_outputs(5467) <= not a;
    layer0_outputs(5468) <= a xor b;
    layer0_outputs(5469) <= a or b;
    layer0_outputs(5470) <= '0';
    layer0_outputs(5471) <= a or b;
    layer0_outputs(5472) <= not b or a;
    layer0_outputs(5473) <= not a or b;
    layer0_outputs(5474) <= a or b;
    layer0_outputs(5475) <= '1';
    layer0_outputs(5476) <= not (a or b);
    layer0_outputs(5477) <= not a;
    layer0_outputs(5478) <= b;
    layer0_outputs(5479) <= b and not a;
    layer0_outputs(5480) <= not b;
    layer0_outputs(5481) <= not a or b;
    layer0_outputs(5482) <= a;
    layer0_outputs(5483) <= a and b;
    layer0_outputs(5484) <= a and not b;
    layer0_outputs(5485) <= not a;
    layer0_outputs(5486) <= not a;
    layer0_outputs(5487) <= not a or b;
    layer0_outputs(5488) <= not a;
    layer0_outputs(5489) <= b and not a;
    layer0_outputs(5490) <= not a;
    layer0_outputs(5491) <= not (a and b);
    layer0_outputs(5492) <= not a;
    layer0_outputs(5493) <= b;
    layer0_outputs(5494) <= not a;
    layer0_outputs(5495) <= not b or a;
    layer0_outputs(5496) <= '1';
    layer0_outputs(5497) <= b;
    layer0_outputs(5498) <= b and not a;
    layer0_outputs(5499) <= not b;
    layer0_outputs(5500) <= '1';
    layer0_outputs(5501) <= a xor b;
    layer0_outputs(5502) <= not a;
    layer0_outputs(5503) <= a;
    layer0_outputs(5504) <= a and not b;
    layer0_outputs(5505) <= not b or a;
    layer0_outputs(5506) <= a xor b;
    layer0_outputs(5507) <= a;
    layer0_outputs(5508) <= '1';
    layer0_outputs(5509) <= a and not b;
    layer0_outputs(5510) <= b;
    layer0_outputs(5511) <= '0';
    layer0_outputs(5512) <= b;
    layer0_outputs(5513) <= not (a and b);
    layer0_outputs(5514) <= '0';
    layer0_outputs(5515) <= not (a and b);
    layer0_outputs(5516) <= not (a or b);
    layer0_outputs(5517) <= not (a or b);
    layer0_outputs(5518) <= not (a and b);
    layer0_outputs(5519) <= a and not b;
    layer0_outputs(5520) <= a;
    layer0_outputs(5521) <= a xor b;
    layer0_outputs(5522) <= '0';
    layer0_outputs(5523) <= '1';
    layer0_outputs(5524) <= a xor b;
    layer0_outputs(5525) <= not a;
    layer0_outputs(5526) <= a and not b;
    layer0_outputs(5527) <= not (a xor b);
    layer0_outputs(5528) <= a or b;
    layer0_outputs(5529) <= not b;
    layer0_outputs(5530) <= not (a or b);
    layer0_outputs(5531) <= a and b;
    layer0_outputs(5532) <= a or b;
    layer0_outputs(5533) <= not b;
    layer0_outputs(5534) <= not (a or b);
    layer0_outputs(5535) <= '0';
    layer0_outputs(5536) <= not (a or b);
    layer0_outputs(5537) <= not (a or b);
    layer0_outputs(5538) <= '1';
    layer0_outputs(5539) <= a and b;
    layer0_outputs(5540) <= a and b;
    layer0_outputs(5541) <= not b;
    layer0_outputs(5542) <= '1';
    layer0_outputs(5543) <= not b;
    layer0_outputs(5544) <= not a or b;
    layer0_outputs(5545) <= '1';
    layer0_outputs(5546) <= not a;
    layer0_outputs(5547) <= not (a and b);
    layer0_outputs(5548) <= not (a xor b);
    layer0_outputs(5549) <= not (a or b);
    layer0_outputs(5550) <= '1';
    layer0_outputs(5551) <= a or b;
    layer0_outputs(5552) <= '1';
    layer0_outputs(5553) <= b and not a;
    layer0_outputs(5554) <= not (a and b);
    layer0_outputs(5555) <= a and not b;
    layer0_outputs(5556) <= b and not a;
    layer0_outputs(5557) <= not b or a;
    layer0_outputs(5558) <= not a or b;
    layer0_outputs(5559) <= not a;
    layer0_outputs(5560) <= a xor b;
    layer0_outputs(5561) <= a xor b;
    layer0_outputs(5562) <= a xor b;
    layer0_outputs(5563) <= not a;
    layer0_outputs(5564) <= not b;
    layer0_outputs(5565) <= a and b;
    layer0_outputs(5566) <= not a or b;
    layer0_outputs(5567) <= not (a xor b);
    layer0_outputs(5568) <= '0';
    layer0_outputs(5569) <= not (a xor b);
    layer0_outputs(5570) <= a and not b;
    layer0_outputs(5571) <= not (a xor b);
    layer0_outputs(5572) <= not (a or b);
    layer0_outputs(5573) <= b;
    layer0_outputs(5574) <= a and b;
    layer0_outputs(5575) <= a;
    layer0_outputs(5576) <= '1';
    layer0_outputs(5577) <= not (a xor b);
    layer0_outputs(5578) <= '1';
    layer0_outputs(5579) <= not a;
    layer0_outputs(5580) <= not b or a;
    layer0_outputs(5581) <= not b or a;
    layer0_outputs(5582) <= '1';
    layer0_outputs(5583) <= not a or b;
    layer0_outputs(5584) <= a;
    layer0_outputs(5585) <= b;
    layer0_outputs(5586) <= not (a and b);
    layer0_outputs(5587) <= not (a and b);
    layer0_outputs(5588) <= '0';
    layer0_outputs(5589) <= a;
    layer0_outputs(5590) <= a and not b;
    layer0_outputs(5591) <= b;
    layer0_outputs(5592) <= not a or b;
    layer0_outputs(5593) <= b and not a;
    layer0_outputs(5594) <= not a or b;
    layer0_outputs(5595) <= a and b;
    layer0_outputs(5596) <= not (a and b);
    layer0_outputs(5597) <= not (a xor b);
    layer0_outputs(5598) <= b and not a;
    layer0_outputs(5599) <= not b;
    layer0_outputs(5600) <= not b;
    layer0_outputs(5601) <= not (a and b);
    layer0_outputs(5602) <= not b or a;
    layer0_outputs(5603) <= not (a and b);
    layer0_outputs(5604) <= b;
    layer0_outputs(5605) <= '0';
    layer0_outputs(5606) <= b;
    layer0_outputs(5607) <= not a or b;
    layer0_outputs(5608) <= not (a or b);
    layer0_outputs(5609) <= '1';
    layer0_outputs(5610) <= a;
    layer0_outputs(5611) <= a xor b;
    layer0_outputs(5612) <= a or b;
    layer0_outputs(5613) <= a;
    layer0_outputs(5614) <= a or b;
    layer0_outputs(5615) <= not b;
    layer0_outputs(5616) <= not b or a;
    layer0_outputs(5617) <= not a;
    layer0_outputs(5618) <= not b or a;
    layer0_outputs(5619) <= '0';
    layer0_outputs(5620) <= not (a and b);
    layer0_outputs(5621) <= not (a and b);
    layer0_outputs(5622) <= a;
    layer0_outputs(5623) <= not b;
    layer0_outputs(5624) <= '1';
    layer0_outputs(5625) <= b;
    layer0_outputs(5626) <= a;
    layer0_outputs(5627) <= a;
    layer0_outputs(5628) <= not (a xor b);
    layer0_outputs(5629) <= a;
    layer0_outputs(5630) <= a or b;
    layer0_outputs(5631) <= b and not a;
    layer0_outputs(5632) <= a and b;
    layer0_outputs(5633) <= a or b;
    layer0_outputs(5634) <= not b;
    layer0_outputs(5635) <= not b or a;
    layer0_outputs(5636) <= not b or a;
    layer0_outputs(5637) <= a and not b;
    layer0_outputs(5638) <= not a;
    layer0_outputs(5639) <= b and not a;
    layer0_outputs(5640) <= '1';
    layer0_outputs(5641) <= '0';
    layer0_outputs(5642) <= '0';
    layer0_outputs(5643) <= not b or a;
    layer0_outputs(5644) <= a;
    layer0_outputs(5645) <= not a or b;
    layer0_outputs(5646) <= a and not b;
    layer0_outputs(5647) <= a and not b;
    layer0_outputs(5648) <= not (a xor b);
    layer0_outputs(5649) <= a or b;
    layer0_outputs(5650) <= not (a or b);
    layer0_outputs(5651) <= a;
    layer0_outputs(5652) <= '0';
    layer0_outputs(5653) <= not (a or b);
    layer0_outputs(5654) <= a and b;
    layer0_outputs(5655) <= b;
    layer0_outputs(5656) <= a or b;
    layer0_outputs(5657) <= b;
    layer0_outputs(5658) <= b and not a;
    layer0_outputs(5659) <= not (a or b);
    layer0_outputs(5660) <= a and not b;
    layer0_outputs(5661) <= b and not a;
    layer0_outputs(5662) <= not b;
    layer0_outputs(5663) <= not a;
    layer0_outputs(5664) <= '0';
    layer0_outputs(5665) <= b and not a;
    layer0_outputs(5666) <= b and not a;
    layer0_outputs(5667) <= not (a xor b);
    layer0_outputs(5668) <= not a or b;
    layer0_outputs(5669) <= not b or a;
    layer0_outputs(5670) <= '0';
    layer0_outputs(5671) <= not (a xor b);
    layer0_outputs(5672) <= not a;
    layer0_outputs(5673) <= not (a xor b);
    layer0_outputs(5674) <= not (a or b);
    layer0_outputs(5675) <= not a or b;
    layer0_outputs(5676) <= a or b;
    layer0_outputs(5677) <= not a;
    layer0_outputs(5678) <= not b or a;
    layer0_outputs(5679) <= not a or b;
    layer0_outputs(5680) <= not (a or b);
    layer0_outputs(5681) <= not (a or b);
    layer0_outputs(5682) <= not (a and b);
    layer0_outputs(5683) <= a or b;
    layer0_outputs(5684) <= not b or a;
    layer0_outputs(5685) <= a and not b;
    layer0_outputs(5686) <= a;
    layer0_outputs(5687) <= b;
    layer0_outputs(5688) <= not a or b;
    layer0_outputs(5689) <= b and not a;
    layer0_outputs(5690) <= not (a xor b);
    layer0_outputs(5691) <= not a;
    layer0_outputs(5692) <= not a;
    layer0_outputs(5693) <= b;
    layer0_outputs(5694) <= not (a or b);
    layer0_outputs(5695) <= b;
    layer0_outputs(5696) <= a;
    layer0_outputs(5697) <= a and b;
    layer0_outputs(5698) <= b;
    layer0_outputs(5699) <= a;
    layer0_outputs(5700) <= not a or b;
    layer0_outputs(5701) <= b and not a;
    layer0_outputs(5702) <= a or b;
    layer0_outputs(5703) <= a and b;
    layer0_outputs(5704) <= '0';
    layer0_outputs(5705) <= a and b;
    layer0_outputs(5706) <= not b or a;
    layer0_outputs(5707) <= not b or a;
    layer0_outputs(5708) <= not (a or b);
    layer0_outputs(5709) <= '1';
    layer0_outputs(5710) <= b;
    layer0_outputs(5711) <= not a;
    layer0_outputs(5712) <= a or b;
    layer0_outputs(5713) <= not (a or b);
    layer0_outputs(5714) <= a;
    layer0_outputs(5715) <= not (a or b);
    layer0_outputs(5716) <= '0';
    layer0_outputs(5717) <= not (a and b);
    layer0_outputs(5718) <= not a or b;
    layer0_outputs(5719) <= a;
    layer0_outputs(5720) <= b and not a;
    layer0_outputs(5721) <= a or b;
    layer0_outputs(5722) <= not (a or b);
    layer0_outputs(5723) <= not (a and b);
    layer0_outputs(5724) <= a xor b;
    layer0_outputs(5725) <= a;
    layer0_outputs(5726) <= not b;
    layer0_outputs(5727) <= a or b;
    layer0_outputs(5728) <= a and b;
    layer0_outputs(5729) <= not (a or b);
    layer0_outputs(5730) <= '0';
    layer0_outputs(5731) <= not a;
    layer0_outputs(5732) <= not a;
    layer0_outputs(5733) <= not (a or b);
    layer0_outputs(5734) <= '1';
    layer0_outputs(5735) <= not b;
    layer0_outputs(5736) <= a or b;
    layer0_outputs(5737) <= b;
    layer0_outputs(5738) <= a or b;
    layer0_outputs(5739) <= '1';
    layer0_outputs(5740) <= '1';
    layer0_outputs(5741) <= not (a or b);
    layer0_outputs(5742) <= not b or a;
    layer0_outputs(5743) <= b;
    layer0_outputs(5744) <= a or b;
    layer0_outputs(5745) <= b;
    layer0_outputs(5746) <= not (a and b);
    layer0_outputs(5747) <= not b;
    layer0_outputs(5748) <= a xor b;
    layer0_outputs(5749) <= a;
    layer0_outputs(5750) <= not (a and b);
    layer0_outputs(5751) <= a;
    layer0_outputs(5752) <= not (a xor b);
    layer0_outputs(5753) <= a and b;
    layer0_outputs(5754) <= a;
    layer0_outputs(5755) <= not a or b;
    layer0_outputs(5756) <= not a or b;
    layer0_outputs(5757) <= '1';
    layer0_outputs(5758) <= '0';
    layer0_outputs(5759) <= not b;
    layer0_outputs(5760) <= a or b;
    layer0_outputs(5761) <= a;
    layer0_outputs(5762) <= not b;
    layer0_outputs(5763) <= not b;
    layer0_outputs(5764) <= a;
    layer0_outputs(5765) <= not a or b;
    layer0_outputs(5766) <= not a;
    layer0_outputs(5767) <= not b;
    layer0_outputs(5768) <= '1';
    layer0_outputs(5769) <= not b;
    layer0_outputs(5770) <= '1';
    layer0_outputs(5771) <= not (a or b);
    layer0_outputs(5772) <= not (a xor b);
    layer0_outputs(5773) <= not a or b;
    layer0_outputs(5774) <= not a or b;
    layer0_outputs(5775) <= a and not b;
    layer0_outputs(5776) <= not b;
    layer0_outputs(5777) <= a xor b;
    layer0_outputs(5778) <= a or b;
    layer0_outputs(5779) <= not (a or b);
    layer0_outputs(5780) <= not a;
    layer0_outputs(5781) <= not b or a;
    layer0_outputs(5782) <= not (a xor b);
    layer0_outputs(5783) <= not (a or b);
    layer0_outputs(5784) <= a;
    layer0_outputs(5785) <= a and b;
    layer0_outputs(5786) <= not b;
    layer0_outputs(5787) <= not b or a;
    layer0_outputs(5788) <= not (a and b);
    layer0_outputs(5789) <= not a or b;
    layer0_outputs(5790) <= not a;
    layer0_outputs(5791) <= '1';
    layer0_outputs(5792) <= '0';
    layer0_outputs(5793) <= b;
    layer0_outputs(5794) <= a or b;
    layer0_outputs(5795) <= not (a or b);
    layer0_outputs(5796) <= not b or a;
    layer0_outputs(5797) <= not a or b;
    layer0_outputs(5798) <= a and not b;
    layer0_outputs(5799) <= not (a and b);
    layer0_outputs(5800) <= not (a or b);
    layer0_outputs(5801) <= a;
    layer0_outputs(5802) <= a and not b;
    layer0_outputs(5803) <= '0';
    layer0_outputs(5804) <= a and b;
    layer0_outputs(5805) <= a xor b;
    layer0_outputs(5806) <= a and b;
    layer0_outputs(5807) <= a;
    layer0_outputs(5808) <= b;
    layer0_outputs(5809) <= a and b;
    layer0_outputs(5810) <= '0';
    layer0_outputs(5811) <= a and not b;
    layer0_outputs(5812) <= a or b;
    layer0_outputs(5813) <= a;
    layer0_outputs(5814) <= '1';
    layer0_outputs(5815) <= b;
    layer0_outputs(5816) <= a or b;
    layer0_outputs(5817) <= '1';
    layer0_outputs(5818) <= not (a or b);
    layer0_outputs(5819) <= a and b;
    layer0_outputs(5820) <= b;
    layer0_outputs(5821) <= a or b;
    layer0_outputs(5822) <= b;
    layer0_outputs(5823) <= b;
    layer0_outputs(5824) <= a and b;
    layer0_outputs(5825) <= not a;
    layer0_outputs(5826) <= not b or a;
    layer0_outputs(5827) <= b and not a;
    layer0_outputs(5828) <= not (a or b);
    layer0_outputs(5829) <= not b or a;
    layer0_outputs(5830) <= not a or b;
    layer0_outputs(5831) <= b;
    layer0_outputs(5832) <= not a;
    layer0_outputs(5833) <= not a or b;
    layer0_outputs(5834) <= '0';
    layer0_outputs(5835) <= not (a and b);
    layer0_outputs(5836) <= '1';
    layer0_outputs(5837) <= not b;
    layer0_outputs(5838) <= '1';
    layer0_outputs(5839) <= a or b;
    layer0_outputs(5840) <= not a;
    layer0_outputs(5841) <= '0';
    layer0_outputs(5842) <= a or b;
    layer0_outputs(5843) <= a and b;
    layer0_outputs(5844) <= not a;
    layer0_outputs(5845) <= a or b;
    layer0_outputs(5846) <= not a;
    layer0_outputs(5847) <= not (a xor b);
    layer0_outputs(5848) <= not b;
    layer0_outputs(5849) <= not b;
    layer0_outputs(5850) <= not b;
    layer0_outputs(5851) <= a or b;
    layer0_outputs(5852) <= not (a xor b);
    layer0_outputs(5853) <= not (a or b);
    layer0_outputs(5854) <= not a or b;
    layer0_outputs(5855) <= b;
    layer0_outputs(5856) <= a;
    layer0_outputs(5857) <= not a or b;
    layer0_outputs(5858) <= a or b;
    layer0_outputs(5859) <= not (a xor b);
    layer0_outputs(5860) <= a;
    layer0_outputs(5861) <= not a or b;
    layer0_outputs(5862) <= '0';
    layer0_outputs(5863) <= not a or b;
    layer0_outputs(5864) <= not a or b;
    layer0_outputs(5865) <= not (a and b);
    layer0_outputs(5866) <= a and b;
    layer0_outputs(5867) <= not (a or b);
    layer0_outputs(5868) <= not (a or b);
    layer0_outputs(5869) <= not b or a;
    layer0_outputs(5870) <= a xor b;
    layer0_outputs(5871) <= not b or a;
    layer0_outputs(5872) <= '1';
    layer0_outputs(5873) <= a or b;
    layer0_outputs(5874) <= '1';
    layer0_outputs(5875) <= not a;
    layer0_outputs(5876) <= a and not b;
    layer0_outputs(5877) <= a or b;
    layer0_outputs(5878) <= not a;
    layer0_outputs(5879) <= '0';
    layer0_outputs(5880) <= a;
    layer0_outputs(5881) <= not (a or b);
    layer0_outputs(5882) <= a and not b;
    layer0_outputs(5883) <= not b;
    layer0_outputs(5884) <= not a or b;
    layer0_outputs(5885) <= a or b;
    layer0_outputs(5886) <= b;
    layer0_outputs(5887) <= '0';
    layer0_outputs(5888) <= not b;
    layer0_outputs(5889) <= not (a and b);
    layer0_outputs(5890) <= '1';
    layer0_outputs(5891) <= not b;
    layer0_outputs(5892) <= not a or b;
    layer0_outputs(5893) <= a xor b;
    layer0_outputs(5894) <= '0';
    layer0_outputs(5895) <= not (a xor b);
    layer0_outputs(5896) <= a xor b;
    layer0_outputs(5897) <= not (a xor b);
    layer0_outputs(5898) <= a;
    layer0_outputs(5899) <= b and not a;
    layer0_outputs(5900) <= a;
    layer0_outputs(5901) <= not a;
    layer0_outputs(5902) <= a xor b;
    layer0_outputs(5903) <= not a;
    layer0_outputs(5904) <= a and not b;
    layer0_outputs(5905) <= a xor b;
    layer0_outputs(5906) <= not b or a;
    layer0_outputs(5907) <= b and not a;
    layer0_outputs(5908) <= '1';
    layer0_outputs(5909) <= not (a and b);
    layer0_outputs(5910) <= not b;
    layer0_outputs(5911) <= a xor b;
    layer0_outputs(5912) <= not a or b;
    layer0_outputs(5913) <= '0';
    layer0_outputs(5914) <= not a;
    layer0_outputs(5915) <= a or b;
    layer0_outputs(5916) <= '0';
    layer0_outputs(5917) <= a and b;
    layer0_outputs(5918) <= not (a or b);
    layer0_outputs(5919) <= '1';
    layer0_outputs(5920) <= not a;
    layer0_outputs(5921) <= not a or b;
    layer0_outputs(5922) <= b;
    layer0_outputs(5923) <= b and not a;
    layer0_outputs(5924) <= not (a xor b);
    layer0_outputs(5925) <= '1';
    layer0_outputs(5926) <= not (a and b);
    layer0_outputs(5927) <= b;
    layer0_outputs(5928) <= a or b;
    layer0_outputs(5929) <= not b or a;
    layer0_outputs(5930) <= not b;
    layer0_outputs(5931) <= a;
    layer0_outputs(5932) <= not (a or b);
    layer0_outputs(5933) <= a xor b;
    layer0_outputs(5934) <= a and not b;
    layer0_outputs(5935) <= not (a xor b);
    layer0_outputs(5936) <= b and not a;
    layer0_outputs(5937) <= a;
    layer0_outputs(5938) <= b and not a;
    layer0_outputs(5939) <= '1';
    layer0_outputs(5940) <= a or b;
    layer0_outputs(5941) <= not b;
    layer0_outputs(5942) <= not (a xor b);
    layer0_outputs(5943) <= not (a and b);
    layer0_outputs(5944) <= a and b;
    layer0_outputs(5945) <= b and not a;
    layer0_outputs(5946) <= not a or b;
    layer0_outputs(5947) <= not (a and b);
    layer0_outputs(5948) <= a and b;
    layer0_outputs(5949) <= a and not b;
    layer0_outputs(5950) <= '1';
    layer0_outputs(5951) <= '0';
    layer0_outputs(5952) <= not b or a;
    layer0_outputs(5953) <= a or b;
    layer0_outputs(5954) <= not a;
    layer0_outputs(5955) <= b and not a;
    layer0_outputs(5956) <= not (a and b);
    layer0_outputs(5957) <= a or b;
    layer0_outputs(5958) <= b;
    layer0_outputs(5959) <= '1';
    layer0_outputs(5960) <= a xor b;
    layer0_outputs(5961) <= b and not a;
    layer0_outputs(5962) <= a and not b;
    layer0_outputs(5963) <= not (a and b);
    layer0_outputs(5964) <= a and not b;
    layer0_outputs(5965) <= b;
    layer0_outputs(5966) <= not b;
    layer0_outputs(5967) <= a or b;
    layer0_outputs(5968) <= not (a and b);
    layer0_outputs(5969) <= not b;
    layer0_outputs(5970) <= not (a and b);
    layer0_outputs(5971) <= not a;
    layer0_outputs(5972) <= not a or b;
    layer0_outputs(5973) <= a;
    layer0_outputs(5974) <= a;
    layer0_outputs(5975) <= a or b;
    layer0_outputs(5976) <= a and not b;
    layer0_outputs(5977) <= a or b;
    layer0_outputs(5978) <= b;
    layer0_outputs(5979) <= a;
    layer0_outputs(5980) <= b and not a;
    layer0_outputs(5981) <= '0';
    layer0_outputs(5982) <= a or b;
    layer0_outputs(5983) <= not b;
    layer0_outputs(5984) <= not (a or b);
    layer0_outputs(5985) <= not (a and b);
    layer0_outputs(5986) <= b and not a;
    layer0_outputs(5987) <= a;
    layer0_outputs(5988) <= '0';
    layer0_outputs(5989) <= a or b;
    layer0_outputs(5990) <= not a or b;
    layer0_outputs(5991) <= a or b;
    layer0_outputs(5992) <= not b;
    layer0_outputs(5993) <= not (a and b);
    layer0_outputs(5994) <= not a;
    layer0_outputs(5995) <= a and not b;
    layer0_outputs(5996) <= b;
    layer0_outputs(5997) <= not (a or b);
    layer0_outputs(5998) <= a xor b;
    layer0_outputs(5999) <= not b;
    layer0_outputs(6000) <= a xor b;
    layer0_outputs(6001) <= '0';
    layer0_outputs(6002) <= a or b;
    layer0_outputs(6003) <= not (a xor b);
    layer0_outputs(6004) <= not (a xor b);
    layer0_outputs(6005) <= '0';
    layer0_outputs(6006) <= not b or a;
    layer0_outputs(6007) <= '0';
    layer0_outputs(6008) <= a and b;
    layer0_outputs(6009) <= a and not b;
    layer0_outputs(6010) <= not (a or b);
    layer0_outputs(6011) <= b and not a;
    layer0_outputs(6012) <= '1';
    layer0_outputs(6013) <= a or b;
    layer0_outputs(6014) <= b and not a;
    layer0_outputs(6015) <= '0';
    layer0_outputs(6016) <= a;
    layer0_outputs(6017) <= a and not b;
    layer0_outputs(6018) <= not (a and b);
    layer0_outputs(6019) <= a;
    layer0_outputs(6020) <= b;
    layer0_outputs(6021) <= not (a xor b);
    layer0_outputs(6022) <= not (a or b);
    layer0_outputs(6023) <= a or b;
    layer0_outputs(6024) <= not (a or b);
    layer0_outputs(6025) <= not a;
    layer0_outputs(6026) <= b and not a;
    layer0_outputs(6027) <= a and not b;
    layer0_outputs(6028) <= not a or b;
    layer0_outputs(6029) <= a and b;
    layer0_outputs(6030) <= not (a xor b);
    layer0_outputs(6031) <= '0';
    layer0_outputs(6032) <= b and not a;
    layer0_outputs(6033) <= a or b;
    layer0_outputs(6034) <= not b or a;
    layer0_outputs(6035) <= a xor b;
    layer0_outputs(6036) <= '1';
    layer0_outputs(6037) <= not (a and b);
    layer0_outputs(6038) <= a;
    layer0_outputs(6039) <= b and not a;
    layer0_outputs(6040) <= not a;
    layer0_outputs(6041) <= not a or b;
    layer0_outputs(6042) <= a;
    layer0_outputs(6043) <= not (a and b);
    layer0_outputs(6044) <= not (a and b);
    layer0_outputs(6045) <= a or b;
    layer0_outputs(6046) <= '1';
    layer0_outputs(6047) <= a and b;
    layer0_outputs(6048) <= not b;
    layer0_outputs(6049) <= not b or a;
    layer0_outputs(6050) <= not a or b;
    layer0_outputs(6051) <= not (a and b);
    layer0_outputs(6052) <= '1';
    layer0_outputs(6053) <= a and not b;
    layer0_outputs(6054) <= not b;
    layer0_outputs(6055) <= a xor b;
    layer0_outputs(6056) <= b;
    layer0_outputs(6057) <= b;
    layer0_outputs(6058) <= not b;
    layer0_outputs(6059) <= not b or a;
    layer0_outputs(6060) <= a;
    layer0_outputs(6061) <= a and not b;
    layer0_outputs(6062) <= '1';
    layer0_outputs(6063) <= not b;
    layer0_outputs(6064) <= a and b;
    layer0_outputs(6065) <= not (a or b);
    layer0_outputs(6066) <= a and b;
    layer0_outputs(6067) <= not a or b;
    layer0_outputs(6068) <= a;
    layer0_outputs(6069) <= a and not b;
    layer0_outputs(6070) <= not b or a;
    layer0_outputs(6071) <= not (a or b);
    layer0_outputs(6072) <= not a;
    layer0_outputs(6073) <= b;
    layer0_outputs(6074) <= not a or b;
    layer0_outputs(6075) <= not a or b;
    layer0_outputs(6076) <= '0';
    layer0_outputs(6077) <= '1';
    layer0_outputs(6078) <= '1';
    layer0_outputs(6079) <= not a or b;
    layer0_outputs(6080) <= not (a or b);
    layer0_outputs(6081) <= not a or b;
    layer0_outputs(6082) <= not b;
    layer0_outputs(6083) <= a;
    layer0_outputs(6084) <= '0';
    layer0_outputs(6085) <= '0';
    layer0_outputs(6086) <= a;
    layer0_outputs(6087) <= not a;
    layer0_outputs(6088) <= not b;
    layer0_outputs(6089) <= not (a and b);
    layer0_outputs(6090) <= b and not a;
    layer0_outputs(6091) <= not (a or b);
    layer0_outputs(6092) <= b;
    layer0_outputs(6093) <= not a or b;
    layer0_outputs(6094) <= a and b;
    layer0_outputs(6095) <= not a;
    layer0_outputs(6096) <= not (a or b);
    layer0_outputs(6097) <= '0';
    layer0_outputs(6098) <= a and not b;
    layer0_outputs(6099) <= a;
    layer0_outputs(6100) <= b and not a;
    layer0_outputs(6101) <= not a;
    layer0_outputs(6102) <= not b or a;
    layer0_outputs(6103) <= a and not b;
    layer0_outputs(6104) <= not (a and b);
    layer0_outputs(6105) <= '0';
    layer0_outputs(6106) <= b and not a;
    layer0_outputs(6107) <= not a;
    layer0_outputs(6108) <= a xor b;
    layer0_outputs(6109) <= '1';
    layer0_outputs(6110) <= a xor b;
    layer0_outputs(6111) <= b;
    layer0_outputs(6112) <= not a;
    layer0_outputs(6113) <= not (a xor b);
    layer0_outputs(6114) <= not b or a;
    layer0_outputs(6115) <= not a or b;
    layer0_outputs(6116) <= '0';
    layer0_outputs(6117) <= a and not b;
    layer0_outputs(6118) <= not b or a;
    layer0_outputs(6119) <= '0';
    layer0_outputs(6120) <= a xor b;
    layer0_outputs(6121) <= a or b;
    layer0_outputs(6122) <= not b;
    layer0_outputs(6123) <= '1';
    layer0_outputs(6124) <= b;
    layer0_outputs(6125) <= not b or a;
    layer0_outputs(6126) <= '1';
    layer0_outputs(6127) <= not a or b;
    layer0_outputs(6128) <= a and b;
    layer0_outputs(6129) <= a;
    layer0_outputs(6130) <= not b or a;
    layer0_outputs(6131) <= not b or a;
    layer0_outputs(6132) <= a xor b;
    layer0_outputs(6133) <= b and not a;
    layer0_outputs(6134) <= '0';
    layer0_outputs(6135) <= not a or b;
    layer0_outputs(6136) <= a;
    layer0_outputs(6137) <= b;
    layer0_outputs(6138) <= not (a and b);
    layer0_outputs(6139) <= not b or a;
    layer0_outputs(6140) <= '1';
    layer0_outputs(6141) <= not (a and b);
    layer0_outputs(6142) <= not (a or b);
    layer0_outputs(6143) <= not a;
    layer0_outputs(6144) <= not b;
    layer0_outputs(6145) <= b and not a;
    layer0_outputs(6146) <= a and not b;
    layer0_outputs(6147) <= not (a and b);
    layer0_outputs(6148) <= a or b;
    layer0_outputs(6149) <= not (a or b);
    layer0_outputs(6150) <= a and not b;
    layer0_outputs(6151) <= a;
    layer0_outputs(6152) <= '0';
    layer0_outputs(6153) <= not a;
    layer0_outputs(6154) <= a;
    layer0_outputs(6155) <= not b or a;
    layer0_outputs(6156) <= a xor b;
    layer0_outputs(6157) <= b;
    layer0_outputs(6158) <= a or b;
    layer0_outputs(6159) <= '1';
    layer0_outputs(6160) <= not (a and b);
    layer0_outputs(6161) <= '0';
    layer0_outputs(6162) <= not b;
    layer0_outputs(6163) <= not b or a;
    layer0_outputs(6164) <= not b or a;
    layer0_outputs(6165) <= not b or a;
    layer0_outputs(6166) <= '0';
    layer0_outputs(6167) <= a;
    layer0_outputs(6168) <= not (a xor b);
    layer0_outputs(6169) <= not (a or b);
    layer0_outputs(6170) <= a and b;
    layer0_outputs(6171) <= not a or b;
    layer0_outputs(6172) <= a and b;
    layer0_outputs(6173) <= not (a or b);
    layer0_outputs(6174) <= b;
    layer0_outputs(6175) <= not a or b;
    layer0_outputs(6176) <= not a;
    layer0_outputs(6177) <= a and not b;
    layer0_outputs(6178) <= '0';
    layer0_outputs(6179) <= a and b;
    layer0_outputs(6180) <= not a or b;
    layer0_outputs(6181) <= not b or a;
    layer0_outputs(6182) <= '1';
    layer0_outputs(6183) <= a xor b;
    layer0_outputs(6184) <= a xor b;
    layer0_outputs(6185) <= not (a or b);
    layer0_outputs(6186) <= a;
    layer0_outputs(6187) <= b;
    layer0_outputs(6188) <= a xor b;
    layer0_outputs(6189) <= not (a or b);
    layer0_outputs(6190) <= '0';
    layer0_outputs(6191) <= b;
    layer0_outputs(6192) <= not a;
    layer0_outputs(6193) <= a;
    layer0_outputs(6194) <= '1';
    layer0_outputs(6195) <= a xor b;
    layer0_outputs(6196) <= a;
    layer0_outputs(6197) <= a xor b;
    layer0_outputs(6198) <= not b;
    layer0_outputs(6199) <= not a or b;
    layer0_outputs(6200) <= not (a xor b);
    layer0_outputs(6201) <= a and b;
    layer0_outputs(6202) <= a and b;
    layer0_outputs(6203) <= b;
    layer0_outputs(6204) <= not a;
    layer0_outputs(6205) <= '0';
    layer0_outputs(6206) <= '0';
    layer0_outputs(6207) <= not b or a;
    layer0_outputs(6208) <= b;
    layer0_outputs(6209) <= not (a or b);
    layer0_outputs(6210) <= a and b;
    layer0_outputs(6211) <= a and not b;
    layer0_outputs(6212) <= b;
    layer0_outputs(6213) <= not b;
    layer0_outputs(6214) <= not a;
    layer0_outputs(6215) <= not a;
    layer0_outputs(6216) <= a or b;
    layer0_outputs(6217) <= b and not a;
    layer0_outputs(6218) <= b and not a;
    layer0_outputs(6219) <= not a or b;
    layer0_outputs(6220) <= b and not a;
    layer0_outputs(6221) <= not a or b;
    layer0_outputs(6222) <= a xor b;
    layer0_outputs(6223) <= not a;
    layer0_outputs(6224) <= not b or a;
    layer0_outputs(6225) <= not a or b;
    layer0_outputs(6226) <= '1';
    layer0_outputs(6227) <= a xor b;
    layer0_outputs(6228) <= not b;
    layer0_outputs(6229) <= a or b;
    layer0_outputs(6230) <= a or b;
    layer0_outputs(6231) <= a and b;
    layer0_outputs(6232) <= '1';
    layer0_outputs(6233) <= a;
    layer0_outputs(6234) <= a or b;
    layer0_outputs(6235) <= not b;
    layer0_outputs(6236) <= not a or b;
    layer0_outputs(6237) <= a;
    layer0_outputs(6238) <= a xor b;
    layer0_outputs(6239) <= a xor b;
    layer0_outputs(6240) <= a and b;
    layer0_outputs(6241) <= '1';
    layer0_outputs(6242) <= a or b;
    layer0_outputs(6243) <= not (a and b);
    layer0_outputs(6244) <= not b or a;
    layer0_outputs(6245) <= b and not a;
    layer0_outputs(6246) <= not (a or b);
    layer0_outputs(6247) <= not (a or b);
    layer0_outputs(6248) <= a and b;
    layer0_outputs(6249) <= not b or a;
    layer0_outputs(6250) <= not b;
    layer0_outputs(6251) <= not b;
    layer0_outputs(6252) <= a and not b;
    layer0_outputs(6253) <= a and b;
    layer0_outputs(6254) <= not (a xor b);
    layer0_outputs(6255) <= a xor b;
    layer0_outputs(6256) <= not (a xor b);
    layer0_outputs(6257) <= not a or b;
    layer0_outputs(6258) <= a and b;
    layer0_outputs(6259) <= not a;
    layer0_outputs(6260) <= not a or b;
    layer0_outputs(6261) <= a or b;
    layer0_outputs(6262) <= '1';
    layer0_outputs(6263) <= not a;
    layer0_outputs(6264) <= '0';
    layer0_outputs(6265) <= not (a and b);
    layer0_outputs(6266) <= not (a xor b);
    layer0_outputs(6267) <= not a or b;
    layer0_outputs(6268) <= a or b;
    layer0_outputs(6269) <= a xor b;
    layer0_outputs(6270) <= b;
    layer0_outputs(6271) <= a xor b;
    layer0_outputs(6272) <= b;
    layer0_outputs(6273) <= a and not b;
    layer0_outputs(6274) <= a or b;
    layer0_outputs(6275) <= b and not a;
    layer0_outputs(6276) <= not b or a;
    layer0_outputs(6277) <= not (a xor b);
    layer0_outputs(6278) <= '0';
    layer0_outputs(6279) <= not a;
    layer0_outputs(6280) <= a and b;
    layer0_outputs(6281) <= not (a xor b);
    layer0_outputs(6282) <= not b;
    layer0_outputs(6283) <= a or b;
    layer0_outputs(6284) <= a;
    layer0_outputs(6285) <= a or b;
    layer0_outputs(6286) <= '1';
    layer0_outputs(6287) <= a xor b;
    layer0_outputs(6288) <= not b;
    layer0_outputs(6289) <= not b;
    layer0_outputs(6290) <= not (a xor b);
    layer0_outputs(6291) <= b;
    layer0_outputs(6292) <= '1';
    layer0_outputs(6293) <= not (a and b);
    layer0_outputs(6294) <= a or b;
    layer0_outputs(6295) <= not (a or b);
    layer0_outputs(6296) <= not b or a;
    layer0_outputs(6297) <= not (a or b);
    layer0_outputs(6298) <= b;
    layer0_outputs(6299) <= not a or b;
    layer0_outputs(6300) <= '0';
    layer0_outputs(6301) <= b;
    layer0_outputs(6302) <= not (a xor b);
    layer0_outputs(6303) <= a and not b;
    layer0_outputs(6304) <= a;
    layer0_outputs(6305) <= a and not b;
    layer0_outputs(6306) <= not b or a;
    layer0_outputs(6307) <= not b or a;
    layer0_outputs(6308) <= b and not a;
    layer0_outputs(6309) <= not (a or b);
    layer0_outputs(6310) <= not a or b;
    layer0_outputs(6311) <= '0';
    layer0_outputs(6312) <= a xor b;
    layer0_outputs(6313) <= b;
    layer0_outputs(6314) <= a and b;
    layer0_outputs(6315) <= '0';
    layer0_outputs(6316) <= b and not a;
    layer0_outputs(6317) <= '1';
    layer0_outputs(6318) <= a;
    layer0_outputs(6319) <= a and not b;
    layer0_outputs(6320) <= not a;
    layer0_outputs(6321) <= a and b;
    layer0_outputs(6322) <= not b or a;
    layer0_outputs(6323) <= '0';
    layer0_outputs(6324) <= not b;
    layer0_outputs(6325) <= a xor b;
    layer0_outputs(6326) <= not (a or b);
    layer0_outputs(6327) <= not b or a;
    layer0_outputs(6328) <= not b or a;
    layer0_outputs(6329) <= a or b;
    layer0_outputs(6330) <= a;
    layer0_outputs(6331) <= a xor b;
    layer0_outputs(6332) <= '1';
    layer0_outputs(6333) <= a xor b;
    layer0_outputs(6334) <= a or b;
    layer0_outputs(6335) <= not (a xor b);
    layer0_outputs(6336) <= not (a and b);
    layer0_outputs(6337) <= a and not b;
    layer0_outputs(6338) <= a;
    layer0_outputs(6339) <= '0';
    layer0_outputs(6340) <= not b;
    layer0_outputs(6341) <= a and b;
    layer0_outputs(6342) <= not a;
    layer0_outputs(6343) <= not (a and b);
    layer0_outputs(6344) <= not (a and b);
    layer0_outputs(6345) <= b;
    layer0_outputs(6346) <= a xor b;
    layer0_outputs(6347) <= not a;
    layer0_outputs(6348) <= '0';
    layer0_outputs(6349) <= not (a xor b);
    layer0_outputs(6350) <= not b;
    layer0_outputs(6351) <= b;
    layer0_outputs(6352) <= not b;
    layer0_outputs(6353) <= a xor b;
    layer0_outputs(6354) <= not (a or b);
    layer0_outputs(6355) <= '0';
    layer0_outputs(6356) <= b and not a;
    layer0_outputs(6357) <= '1';
    layer0_outputs(6358) <= '0';
    layer0_outputs(6359) <= a or b;
    layer0_outputs(6360) <= not (a xor b);
    layer0_outputs(6361) <= a and not b;
    layer0_outputs(6362) <= not a;
    layer0_outputs(6363) <= not b or a;
    layer0_outputs(6364) <= not b or a;
    layer0_outputs(6365) <= not a;
    layer0_outputs(6366) <= b and not a;
    layer0_outputs(6367) <= b and not a;
    layer0_outputs(6368) <= a and not b;
    layer0_outputs(6369) <= not (a and b);
    layer0_outputs(6370) <= not (a and b);
    layer0_outputs(6371) <= b and not a;
    layer0_outputs(6372) <= not a or b;
    layer0_outputs(6373) <= a and not b;
    layer0_outputs(6374) <= not (a or b);
    layer0_outputs(6375) <= b;
    layer0_outputs(6376) <= not a or b;
    layer0_outputs(6377) <= a;
    layer0_outputs(6378) <= b and not a;
    layer0_outputs(6379) <= not b or a;
    layer0_outputs(6380) <= a and b;
    layer0_outputs(6381) <= a xor b;
    layer0_outputs(6382) <= not a;
    layer0_outputs(6383) <= b;
    layer0_outputs(6384) <= not (a or b);
    layer0_outputs(6385) <= b and not a;
    layer0_outputs(6386) <= '1';
    layer0_outputs(6387) <= not (a and b);
    layer0_outputs(6388) <= not b;
    layer0_outputs(6389) <= not a or b;
    layer0_outputs(6390) <= a and not b;
    layer0_outputs(6391) <= not a or b;
    layer0_outputs(6392) <= '1';
    layer0_outputs(6393) <= a or b;
    layer0_outputs(6394) <= a xor b;
    layer0_outputs(6395) <= not a or b;
    layer0_outputs(6396) <= b and not a;
    layer0_outputs(6397) <= not a or b;
    layer0_outputs(6398) <= not a or b;
    layer0_outputs(6399) <= not b;
    layer0_outputs(6400) <= not (a or b);
    layer0_outputs(6401) <= a and not b;
    layer0_outputs(6402) <= a and not b;
    layer0_outputs(6403) <= b;
    layer0_outputs(6404) <= not (a xor b);
    layer0_outputs(6405) <= not b;
    layer0_outputs(6406) <= not a or b;
    layer0_outputs(6407) <= b;
    layer0_outputs(6408) <= not (a xor b);
    layer0_outputs(6409) <= '1';
    layer0_outputs(6410) <= not a or b;
    layer0_outputs(6411) <= not (a xor b);
    layer0_outputs(6412) <= '1';
    layer0_outputs(6413) <= not a or b;
    layer0_outputs(6414) <= not a;
    layer0_outputs(6415) <= a and not b;
    layer0_outputs(6416) <= '0';
    layer0_outputs(6417) <= a;
    layer0_outputs(6418) <= b and not a;
    layer0_outputs(6419) <= b and not a;
    layer0_outputs(6420) <= '0';
    layer0_outputs(6421) <= not (a xor b);
    layer0_outputs(6422) <= a and not b;
    layer0_outputs(6423) <= not (a and b);
    layer0_outputs(6424) <= not b or a;
    layer0_outputs(6425) <= '1';
    layer0_outputs(6426) <= a;
    layer0_outputs(6427) <= not a or b;
    layer0_outputs(6428) <= a or b;
    layer0_outputs(6429) <= a;
    layer0_outputs(6430) <= not (a or b);
    layer0_outputs(6431) <= b and not a;
    layer0_outputs(6432) <= a and not b;
    layer0_outputs(6433) <= '0';
    layer0_outputs(6434) <= not (a xor b);
    layer0_outputs(6435) <= not (a xor b);
    layer0_outputs(6436) <= '0';
    layer0_outputs(6437) <= not (a or b);
    layer0_outputs(6438) <= not a;
    layer0_outputs(6439) <= '0';
    layer0_outputs(6440) <= b and not a;
    layer0_outputs(6441) <= a xor b;
    layer0_outputs(6442) <= a;
    layer0_outputs(6443) <= '0';
    layer0_outputs(6444) <= not a;
    layer0_outputs(6445) <= not (a and b);
    layer0_outputs(6446) <= not (a and b);
    layer0_outputs(6447) <= not b;
    layer0_outputs(6448) <= b;
    layer0_outputs(6449) <= not b or a;
    layer0_outputs(6450) <= not b;
    layer0_outputs(6451) <= not (a or b);
    layer0_outputs(6452) <= a or b;
    layer0_outputs(6453) <= a;
    layer0_outputs(6454) <= a and b;
    layer0_outputs(6455) <= not a;
    layer0_outputs(6456) <= '0';
    layer0_outputs(6457) <= a;
    layer0_outputs(6458) <= not (a or b);
    layer0_outputs(6459) <= a and not b;
    layer0_outputs(6460) <= not (a or b);
    layer0_outputs(6461) <= '1';
    layer0_outputs(6462) <= '1';
    layer0_outputs(6463) <= '1';
    layer0_outputs(6464) <= b and not a;
    layer0_outputs(6465) <= not (a and b);
    layer0_outputs(6466) <= b and not a;
    layer0_outputs(6467) <= not (a or b);
    layer0_outputs(6468) <= not (a xor b);
    layer0_outputs(6469) <= not b or a;
    layer0_outputs(6470) <= b and not a;
    layer0_outputs(6471) <= not (a xor b);
    layer0_outputs(6472) <= not b or a;
    layer0_outputs(6473) <= '1';
    layer0_outputs(6474) <= not b or a;
    layer0_outputs(6475) <= not (a or b);
    layer0_outputs(6476) <= a and not b;
    layer0_outputs(6477) <= '0';
    layer0_outputs(6478) <= '1';
    layer0_outputs(6479) <= a and b;
    layer0_outputs(6480) <= a xor b;
    layer0_outputs(6481) <= not (a and b);
    layer0_outputs(6482) <= a and not b;
    layer0_outputs(6483) <= a and b;
    layer0_outputs(6484) <= a xor b;
    layer0_outputs(6485) <= a;
    layer0_outputs(6486) <= a;
    layer0_outputs(6487) <= not b;
    layer0_outputs(6488) <= not (a or b);
    layer0_outputs(6489) <= '1';
    layer0_outputs(6490) <= '1';
    layer0_outputs(6491) <= a and not b;
    layer0_outputs(6492) <= a xor b;
    layer0_outputs(6493) <= b and not a;
    layer0_outputs(6494) <= a and not b;
    layer0_outputs(6495) <= b and not a;
    layer0_outputs(6496) <= not a;
    layer0_outputs(6497) <= a and b;
    layer0_outputs(6498) <= b and not a;
    layer0_outputs(6499) <= not a;
    layer0_outputs(6500) <= not b or a;
    layer0_outputs(6501) <= not a;
    layer0_outputs(6502) <= '1';
    layer0_outputs(6503) <= a and not b;
    layer0_outputs(6504) <= '1';
    layer0_outputs(6505) <= not b or a;
    layer0_outputs(6506) <= a and not b;
    layer0_outputs(6507) <= a and not b;
    layer0_outputs(6508) <= b;
    layer0_outputs(6509) <= not (a xor b);
    layer0_outputs(6510) <= b and not a;
    layer0_outputs(6511) <= not (a or b);
    layer0_outputs(6512) <= a or b;
    layer0_outputs(6513) <= a or b;
    layer0_outputs(6514) <= a xor b;
    layer0_outputs(6515) <= '1';
    layer0_outputs(6516) <= a and not b;
    layer0_outputs(6517) <= not (a or b);
    layer0_outputs(6518) <= not (a xor b);
    layer0_outputs(6519) <= '0';
    layer0_outputs(6520) <= b and not a;
    layer0_outputs(6521) <= a xor b;
    layer0_outputs(6522) <= not (a or b);
    layer0_outputs(6523) <= not b;
    layer0_outputs(6524) <= '1';
    layer0_outputs(6525) <= not b;
    layer0_outputs(6526) <= not a or b;
    layer0_outputs(6527) <= '1';
    layer0_outputs(6528) <= b and not a;
    layer0_outputs(6529) <= not b or a;
    layer0_outputs(6530) <= not (a xor b);
    layer0_outputs(6531) <= a and b;
    layer0_outputs(6532) <= '0';
    layer0_outputs(6533) <= not a;
    layer0_outputs(6534) <= a or b;
    layer0_outputs(6535) <= a xor b;
    layer0_outputs(6536) <= not (a xor b);
    layer0_outputs(6537) <= b;
    layer0_outputs(6538) <= not (a and b);
    layer0_outputs(6539) <= '0';
    layer0_outputs(6540) <= b and not a;
    layer0_outputs(6541) <= b;
    layer0_outputs(6542) <= a and not b;
    layer0_outputs(6543) <= not b;
    layer0_outputs(6544) <= '1';
    layer0_outputs(6545) <= a and b;
    layer0_outputs(6546) <= '0';
    layer0_outputs(6547) <= not a;
    layer0_outputs(6548) <= '0';
    layer0_outputs(6549) <= not a or b;
    layer0_outputs(6550) <= not b;
    layer0_outputs(6551) <= a and not b;
    layer0_outputs(6552) <= a xor b;
    layer0_outputs(6553) <= a xor b;
    layer0_outputs(6554) <= '0';
    layer0_outputs(6555) <= not (a or b);
    layer0_outputs(6556) <= a and not b;
    layer0_outputs(6557) <= a or b;
    layer0_outputs(6558) <= '0';
    layer0_outputs(6559) <= a and not b;
    layer0_outputs(6560) <= not (a or b);
    layer0_outputs(6561) <= a xor b;
    layer0_outputs(6562) <= a;
    layer0_outputs(6563) <= a and not b;
    layer0_outputs(6564) <= not b or a;
    layer0_outputs(6565) <= not b or a;
    layer0_outputs(6566) <= '0';
    layer0_outputs(6567) <= a and not b;
    layer0_outputs(6568) <= not (a xor b);
    layer0_outputs(6569) <= a;
    layer0_outputs(6570) <= not b;
    layer0_outputs(6571) <= a and b;
    layer0_outputs(6572) <= '1';
    layer0_outputs(6573) <= '1';
    layer0_outputs(6574) <= a and not b;
    layer0_outputs(6575) <= not (a or b);
    layer0_outputs(6576) <= not b or a;
    layer0_outputs(6577) <= a or b;
    layer0_outputs(6578) <= a;
    layer0_outputs(6579) <= not (a xor b);
    layer0_outputs(6580) <= not b;
    layer0_outputs(6581) <= a xor b;
    layer0_outputs(6582) <= '1';
    layer0_outputs(6583) <= not b;
    layer0_outputs(6584) <= a and b;
    layer0_outputs(6585) <= '0';
    layer0_outputs(6586) <= a and not b;
    layer0_outputs(6587) <= '1';
    layer0_outputs(6588) <= a and not b;
    layer0_outputs(6589) <= '1';
    layer0_outputs(6590) <= b and not a;
    layer0_outputs(6591) <= not a;
    layer0_outputs(6592) <= a;
    layer0_outputs(6593) <= '0';
    layer0_outputs(6594) <= not a;
    layer0_outputs(6595) <= not a or b;
    layer0_outputs(6596) <= a;
    layer0_outputs(6597) <= b;
    layer0_outputs(6598) <= a or b;
    layer0_outputs(6599) <= '1';
    layer0_outputs(6600) <= not (a xor b);
    layer0_outputs(6601) <= '0';
    layer0_outputs(6602) <= b and not a;
    layer0_outputs(6603) <= not (a and b);
    layer0_outputs(6604) <= '0';
    layer0_outputs(6605) <= not (a xor b);
    layer0_outputs(6606) <= a and b;
    layer0_outputs(6607) <= not (a or b);
    layer0_outputs(6608) <= not (a or b);
    layer0_outputs(6609) <= a xor b;
    layer0_outputs(6610) <= not a;
    layer0_outputs(6611) <= b;
    layer0_outputs(6612) <= a xor b;
    layer0_outputs(6613) <= b and not a;
    layer0_outputs(6614) <= '0';
    layer0_outputs(6615) <= '0';
    layer0_outputs(6616) <= a;
    layer0_outputs(6617) <= b;
    layer0_outputs(6618) <= '1';
    layer0_outputs(6619) <= not b or a;
    layer0_outputs(6620) <= b;
    layer0_outputs(6621) <= a or b;
    layer0_outputs(6622) <= b;
    layer0_outputs(6623) <= a and not b;
    layer0_outputs(6624) <= not (a and b);
    layer0_outputs(6625) <= not b or a;
    layer0_outputs(6626) <= b;
    layer0_outputs(6627) <= not (a or b);
    layer0_outputs(6628) <= not a;
    layer0_outputs(6629) <= a and b;
    layer0_outputs(6630) <= not a or b;
    layer0_outputs(6631) <= a and b;
    layer0_outputs(6632) <= not (a or b);
    layer0_outputs(6633) <= not (a xor b);
    layer0_outputs(6634) <= b;
    layer0_outputs(6635) <= '1';
    layer0_outputs(6636) <= not (a and b);
    layer0_outputs(6637) <= a xor b;
    layer0_outputs(6638) <= a;
    layer0_outputs(6639) <= b;
    layer0_outputs(6640) <= b;
    layer0_outputs(6641) <= a xor b;
    layer0_outputs(6642) <= not a;
    layer0_outputs(6643) <= a or b;
    layer0_outputs(6644) <= not (a and b);
    layer0_outputs(6645) <= not b;
    layer0_outputs(6646) <= a xor b;
    layer0_outputs(6647) <= a and not b;
    layer0_outputs(6648) <= b and not a;
    layer0_outputs(6649) <= not a;
    layer0_outputs(6650) <= not a;
    layer0_outputs(6651) <= not (a and b);
    layer0_outputs(6652) <= b;
    layer0_outputs(6653) <= a and b;
    layer0_outputs(6654) <= a;
    layer0_outputs(6655) <= b and not a;
    layer0_outputs(6656) <= not (a and b);
    layer0_outputs(6657) <= b;
    layer0_outputs(6658) <= '1';
    layer0_outputs(6659) <= a xor b;
    layer0_outputs(6660) <= a or b;
    layer0_outputs(6661) <= a xor b;
    layer0_outputs(6662) <= a and b;
    layer0_outputs(6663) <= b and not a;
    layer0_outputs(6664) <= a and not b;
    layer0_outputs(6665) <= a and b;
    layer0_outputs(6666) <= '0';
    layer0_outputs(6667) <= not a or b;
    layer0_outputs(6668) <= not b;
    layer0_outputs(6669) <= not b;
    layer0_outputs(6670) <= a;
    layer0_outputs(6671) <= a xor b;
    layer0_outputs(6672) <= a xor b;
    layer0_outputs(6673) <= a and b;
    layer0_outputs(6674) <= not (a xor b);
    layer0_outputs(6675) <= not b or a;
    layer0_outputs(6676) <= a xor b;
    layer0_outputs(6677) <= not b or a;
    layer0_outputs(6678) <= a and not b;
    layer0_outputs(6679) <= '0';
    layer0_outputs(6680) <= a or b;
    layer0_outputs(6681) <= a and not b;
    layer0_outputs(6682) <= a;
    layer0_outputs(6683) <= not b;
    layer0_outputs(6684) <= a and not b;
    layer0_outputs(6685) <= b and not a;
    layer0_outputs(6686) <= not b;
    layer0_outputs(6687) <= not a;
    layer0_outputs(6688) <= not a;
    layer0_outputs(6689) <= a and not b;
    layer0_outputs(6690) <= a;
    layer0_outputs(6691) <= '0';
    layer0_outputs(6692) <= not b;
    layer0_outputs(6693) <= not a;
    layer0_outputs(6694) <= a or b;
    layer0_outputs(6695) <= a or b;
    layer0_outputs(6696) <= not b;
    layer0_outputs(6697) <= a and b;
    layer0_outputs(6698) <= b and not a;
    layer0_outputs(6699) <= b and not a;
    layer0_outputs(6700) <= b and not a;
    layer0_outputs(6701) <= '1';
    layer0_outputs(6702) <= a and not b;
    layer0_outputs(6703) <= b;
    layer0_outputs(6704) <= a and b;
    layer0_outputs(6705) <= a;
    layer0_outputs(6706) <= not a or b;
    layer0_outputs(6707) <= not b;
    layer0_outputs(6708) <= a and b;
    layer0_outputs(6709) <= '0';
    layer0_outputs(6710) <= a xor b;
    layer0_outputs(6711) <= b;
    layer0_outputs(6712) <= a xor b;
    layer0_outputs(6713) <= b and not a;
    layer0_outputs(6714) <= b;
    layer0_outputs(6715) <= not a or b;
    layer0_outputs(6716) <= b and not a;
    layer0_outputs(6717) <= not b;
    layer0_outputs(6718) <= '1';
    layer0_outputs(6719) <= a or b;
    layer0_outputs(6720) <= '0';
    layer0_outputs(6721) <= b and not a;
    layer0_outputs(6722) <= a or b;
    layer0_outputs(6723) <= not (a and b);
    layer0_outputs(6724) <= a;
    layer0_outputs(6725) <= not a;
    layer0_outputs(6726) <= not a or b;
    layer0_outputs(6727) <= b and not a;
    layer0_outputs(6728) <= not b or a;
    layer0_outputs(6729) <= '1';
    layer0_outputs(6730) <= '1';
    layer0_outputs(6731) <= b;
    layer0_outputs(6732) <= a and not b;
    layer0_outputs(6733) <= '1';
    layer0_outputs(6734) <= '0';
    layer0_outputs(6735) <= not b;
    layer0_outputs(6736) <= not (a and b);
    layer0_outputs(6737) <= '1';
    layer0_outputs(6738) <= not b or a;
    layer0_outputs(6739) <= '0';
    layer0_outputs(6740) <= not b;
    layer0_outputs(6741) <= '0';
    layer0_outputs(6742) <= a or b;
    layer0_outputs(6743) <= a and b;
    layer0_outputs(6744) <= not b or a;
    layer0_outputs(6745) <= b and not a;
    layer0_outputs(6746) <= not b or a;
    layer0_outputs(6747) <= a;
    layer0_outputs(6748) <= a and b;
    layer0_outputs(6749) <= a and b;
    layer0_outputs(6750) <= not b or a;
    layer0_outputs(6751) <= b and not a;
    layer0_outputs(6752) <= a or b;
    layer0_outputs(6753) <= '0';
    layer0_outputs(6754) <= not (a xor b);
    layer0_outputs(6755) <= '0';
    layer0_outputs(6756) <= '1';
    layer0_outputs(6757) <= not b;
    layer0_outputs(6758) <= a or b;
    layer0_outputs(6759) <= b and not a;
    layer0_outputs(6760) <= not (a and b);
    layer0_outputs(6761) <= a xor b;
    layer0_outputs(6762) <= not b or a;
    layer0_outputs(6763) <= b and not a;
    layer0_outputs(6764) <= a xor b;
    layer0_outputs(6765) <= not (a and b);
    layer0_outputs(6766) <= not a or b;
    layer0_outputs(6767) <= a and b;
    layer0_outputs(6768) <= not b or a;
    layer0_outputs(6769) <= a or b;
    layer0_outputs(6770) <= not (a and b);
    layer0_outputs(6771) <= '1';
    layer0_outputs(6772) <= not a or b;
    layer0_outputs(6773) <= not b or a;
    layer0_outputs(6774) <= '0';
    layer0_outputs(6775) <= not (a and b);
    layer0_outputs(6776) <= not a or b;
    layer0_outputs(6777) <= not (a xor b);
    layer0_outputs(6778) <= a xor b;
    layer0_outputs(6779) <= a and not b;
    layer0_outputs(6780) <= a;
    layer0_outputs(6781) <= a and b;
    layer0_outputs(6782) <= not b;
    layer0_outputs(6783) <= a and not b;
    layer0_outputs(6784) <= a or b;
    layer0_outputs(6785) <= not (a and b);
    layer0_outputs(6786) <= a xor b;
    layer0_outputs(6787) <= a and b;
    layer0_outputs(6788) <= not b or a;
    layer0_outputs(6789) <= not (a and b);
    layer0_outputs(6790) <= b and not a;
    layer0_outputs(6791) <= a;
    layer0_outputs(6792) <= '1';
    layer0_outputs(6793) <= '0';
    layer0_outputs(6794) <= a or b;
    layer0_outputs(6795) <= not (a and b);
    layer0_outputs(6796) <= '1';
    layer0_outputs(6797) <= a or b;
    layer0_outputs(6798) <= not a;
    layer0_outputs(6799) <= b and not a;
    layer0_outputs(6800) <= not b or a;
    layer0_outputs(6801) <= '1';
    layer0_outputs(6802) <= not b or a;
    layer0_outputs(6803) <= a or b;
    layer0_outputs(6804) <= not a or b;
    layer0_outputs(6805) <= a;
    layer0_outputs(6806) <= a and not b;
    layer0_outputs(6807) <= not a or b;
    layer0_outputs(6808) <= not (a xor b);
    layer0_outputs(6809) <= not a or b;
    layer0_outputs(6810) <= not a;
    layer0_outputs(6811) <= a and b;
    layer0_outputs(6812) <= b and not a;
    layer0_outputs(6813) <= b;
    layer0_outputs(6814) <= not (a or b);
    layer0_outputs(6815) <= not (a or b);
    layer0_outputs(6816) <= a;
    layer0_outputs(6817) <= a or b;
    layer0_outputs(6818) <= not (a and b);
    layer0_outputs(6819) <= '1';
    layer0_outputs(6820) <= '1';
    layer0_outputs(6821) <= a;
    layer0_outputs(6822) <= a and b;
    layer0_outputs(6823) <= a;
    layer0_outputs(6824) <= not a;
    layer0_outputs(6825) <= a or b;
    layer0_outputs(6826) <= not (a xor b);
    layer0_outputs(6827) <= not a;
    layer0_outputs(6828) <= b and not a;
    layer0_outputs(6829) <= '0';
    layer0_outputs(6830) <= not a;
    layer0_outputs(6831) <= not b;
    layer0_outputs(6832) <= not a or b;
    layer0_outputs(6833) <= a and not b;
    layer0_outputs(6834) <= '1';
    layer0_outputs(6835) <= not a or b;
    layer0_outputs(6836) <= a or b;
    layer0_outputs(6837) <= not b;
    layer0_outputs(6838) <= a and not b;
    layer0_outputs(6839) <= a or b;
    layer0_outputs(6840) <= not b or a;
    layer0_outputs(6841) <= not (a xor b);
    layer0_outputs(6842) <= a or b;
    layer0_outputs(6843) <= b;
    layer0_outputs(6844) <= not a or b;
    layer0_outputs(6845) <= not a;
    layer0_outputs(6846) <= a and b;
    layer0_outputs(6847) <= a and b;
    layer0_outputs(6848) <= a and not b;
    layer0_outputs(6849) <= a;
    layer0_outputs(6850) <= not b;
    layer0_outputs(6851) <= '0';
    layer0_outputs(6852) <= '0';
    layer0_outputs(6853) <= a;
    layer0_outputs(6854) <= a;
    layer0_outputs(6855) <= not (a or b);
    layer0_outputs(6856) <= a and not b;
    layer0_outputs(6857) <= a or b;
    layer0_outputs(6858) <= not (a or b);
    layer0_outputs(6859) <= a and b;
    layer0_outputs(6860) <= not a;
    layer0_outputs(6861) <= b;
    layer0_outputs(6862) <= a and b;
    layer0_outputs(6863) <= not (a and b);
    layer0_outputs(6864) <= b and not a;
    layer0_outputs(6865) <= not b or a;
    layer0_outputs(6866) <= not (a and b);
    layer0_outputs(6867) <= not b;
    layer0_outputs(6868) <= '1';
    layer0_outputs(6869) <= not (a or b);
    layer0_outputs(6870) <= not (a and b);
    layer0_outputs(6871) <= not (a or b);
    layer0_outputs(6872) <= a;
    layer0_outputs(6873) <= not (a or b);
    layer0_outputs(6874) <= a or b;
    layer0_outputs(6875) <= b and not a;
    layer0_outputs(6876) <= '1';
    layer0_outputs(6877) <= not b;
    layer0_outputs(6878) <= not a or b;
    layer0_outputs(6879) <= not (a or b);
    layer0_outputs(6880) <= a and not b;
    layer0_outputs(6881) <= not (a and b);
    layer0_outputs(6882) <= a xor b;
    layer0_outputs(6883) <= a and b;
    layer0_outputs(6884) <= not a or b;
    layer0_outputs(6885) <= not a or b;
    layer0_outputs(6886) <= not (a xor b);
    layer0_outputs(6887) <= b and not a;
    layer0_outputs(6888) <= not a or b;
    layer0_outputs(6889) <= a and not b;
    layer0_outputs(6890) <= b;
    layer0_outputs(6891) <= a and b;
    layer0_outputs(6892) <= a xor b;
    layer0_outputs(6893) <= not a;
    layer0_outputs(6894) <= a or b;
    layer0_outputs(6895) <= not b or a;
    layer0_outputs(6896) <= a;
    layer0_outputs(6897) <= a or b;
    layer0_outputs(6898) <= not b or a;
    layer0_outputs(6899) <= a;
    layer0_outputs(6900) <= not (a or b);
    layer0_outputs(6901) <= not (a or b);
    layer0_outputs(6902) <= not a or b;
    layer0_outputs(6903) <= not (a and b);
    layer0_outputs(6904) <= b;
    layer0_outputs(6905) <= '1';
    layer0_outputs(6906) <= a or b;
    layer0_outputs(6907) <= a or b;
    layer0_outputs(6908) <= not (a and b);
    layer0_outputs(6909) <= a and b;
    layer0_outputs(6910) <= not (a and b);
    layer0_outputs(6911) <= not a or b;
    layer0_outputs(6912) <= b;
    layer0_outputs(6913) <= not a;
    layer0_outputs(6914) <= not b or a;
    layer0_outputs(6915) <= a and b;
    layer0_outputs(6916) <= not a;
    layer0_outputs(6917) <= not a or b;
    layer0_outputs(6918) <= a or b;
    layer0_outputs(6919) <= not b;
    layer0_outputs(6920) <= not b;
    layer0_outputs(6921) <= not b or a;
    layer0_outputs(6922) <= b;
    layer0_outputs(6923) <= a or b;
    layer0_outputs(6924) <= a and not b;
    layer0_outputs(6925) <= a and b;
    layer0_outputs(6926) <= '0';
    layer0_outputs(6927) <= not (a and b);
    layer0_outputs(6928) <= not (a and b);
    layer0_outputs(6929) <= a and b;
    layer0_outputs(6930) <= '1';
    layer0_outputs(6931) <= a and not b;
    layer0_outputs(6932) <= a and b;
    layer0_outputs(6933) <= not (a or b);
    layer0_outputs(6934) <= a or b;
    layer0_outputs(6935) <= '0';
    layer0_outputs(6936) <= not (a and b);
    layer0_outputs(6937) <= not (a or b);
    layer0_outputs(6938) <= '1';
    layer0_outputs(6939) <= not a;
    layer0_outputs(6940) <= not (a xor b);
    layer0_outputs(6941) <= not (a xor b);
    layer0_outputs(6942) <= a;
    layer0_outputs(6943) <= b and not a;
    layer0_outputs(6944) <= a or b;
    layer0_outputs(6945) <= not (a xor b);
    layer0_outputs(6946) <= '1';
    layer0_outputs(6947) <= not (a xor b);
    layer0_outputs(6948) <= a and b;
    layer0_outputs(6949) <= '0';
    layer0_outputs(6950) <= not b;
    layer0_outputs(6951) <= '1';
    layer0_outputs(6952) <= not a or b;
    layer0_outputs(6953) <= not a;
    layer0_outputs(6954) <= b and not a;
    layer0_outputs(6955) <= a and b;
    layer0_outputs(6956) <= not (a or b);
    layer0_outputs(6957) <= '0';
    layer0_outputs(6958) <= not b or a;
    layer0_outputs(6959) <= not b;
    layer0_outputs(6960) <= not (a or b);
    layer0_outputs(6961) <= '1';
    layer0_outputs(6962) <= not (a and b);
    layer0_outputs(6963) <= not a;
    layer0_outputs(6964) <= a and not b;
    layer0_outputs(6965) <= a and b;
    layer0_outputs(6966) <= a or b;
    layer0_outputs(6967) <= a or b;
    layer0_outputs(6968) <= a;
    layer0_outputs(6969) <= not (a or b);
    layer0_outputs(6970) <= not b;
    layer0_outputs(6971) <= not a;
    layer0_outputs(6972) <= not a;
    layer0_outputs(6973) <= a or b;
    layer0_outputs(6974) <= a and b;
    layer0_outputs(6975) <= a and b;
    layer0_outputs(6976) <= not a;
    layer0_outputs(6977) <= a xor b;
    layer0_outputs(6978) <= not a;
    layer0_outputs(6979) <= not (a and b);
    layer0_outputs(6980) <= b;
    layer0_outputs(6981) <= not b;
    layer0_outputs(6982) <= a and not b;
    layer0_outputs(6983) <= '0';
    layer0_outputs(6984) <= '1';
    layer0_outputs(6985) <= not a;
    layer0_outputs(6986) <= a or b;
    layer0_outputs(6987) <= a xor b;
    layer0_outputs(6988) <= not b;
    layer0_outputs(6989) <= '1';
    layer0_outputs(6990) <= not a;
    layer0_outputs(6991) <= not b or a;
    layer0_outputs(6992) <= a and b;
    layer0_outputs(6993) <= '0';
    layer0_outputs(6994) <= a xor b;
    layer0_outputs(6995) <= a or b;
    layer0_outputs(6996) <= b;
    layer0_outputs(6997) <= not (a xor b);
    layer0_outputs(6998) <= not (a and b);
    layer0_outputs(6999) <= not a or b;
    layer0_outputs(7000) <= a;
    layer0_outputs(7001) <= not b;
    layer0_outputs(7002) <= a;
    layer0_outputs(7003) <= a;
    layer0_outputs(7004) <= a and b;
    layer0_outputs(7005) <= not (a and b);
    layer0_outputs(7006) <= not (a or b);
    layer0_outputs(7007) <= b and not a;
    layer0_outputs(7008) <= not a;
    layer0_outputs(7009) <= a and b;
    layer0_outputs(7010) <= not a;
    layer0_outputs(7011) <= not b;
    layer0_outputs(7012) <= a or b;
    layer0_outputs(7013) <= a and not b;
    layer0_outputs(7014) <= not b or a;
    layer0_outputs(7015) <= not a;
    layer0_outputs(7016) <= not (a and b);
    layer0_outputs(7017) <= not b or a;
    layer0_outputs(7018) <= a;
    layer0_outputs(7019) <= a and not b;
    layer0_outputs(7020) <= not (a xor b);
    layer0_outputs(7021) <= not a or b;
    layer0_outputs(7022) <= not (a or b);
    layer0_outputs(7023) <= b;
    layer0_outputs(7024) <= a and b;
    layer0_outputs(7025) <= not a or b;
    layer0_outputs(7026) <= not a;
    layer0_outputs(7027) <= a or b;
    layer0_outputs(7028) <= b and not a;
    layer0_outputs(7029) <= '0';
    layer0_outputs(7030) <= '0';
    layer0_outputs(7031) <= a and not b;
    layer0_outputs(7032) <= b;
    layer0_outputs(7033) <= not (a and b);
    layer0_outputs(7034) <= b;
    layer0_outputs(7035) <= b and not a;
    layer0_outputs(7036) <= not b;
    layer0_outputs(7037) <= not a;
    layer0_outputs(7038) <= not (a or b);
    layer0_outputs(7039) <= not a;
    layer0_outputs(7040) <= a or b;
    layer0_outputs(7041) <= b;
    layer0_outputs(7042) <= '1';
    layer0_outputs(7043) <= not b;
    layer0_outputs(7044) <= not (a or b);
    layer0_outputs(7045) <= not (a or b);
    layer0_outputs(7046) <= a;
    layer0_outputs(7047) <= a;
    layer0_outputs(7048) <= a or b;
    layer0_outputs(7049) <= not (a or b);
    layer0_outputs(7050) <= a or b;
    layer0_outputs(7051) <= b;
    layer0_outputs(7052) <= not (a or b);
    layer0_outputs(7053) <= a and not b;
    layer0_outputs(7054) <= b and not a;
    layer0_outputs(7055) <= a and not b;
    layer0_outputs(7056) <= not b;
    layer0_outputs(7057) <= '0';
    layer0_outputs(7058) <= a;
    layer0_outputs(7059) <= not b;
    layer0_outputs(7060) <= b and not a;
    layer0_outputs(7061) <= '0';
    layer0_outputs(7062) <= not a or b;
    layer0_outputs(7063) <= not b;
    layer0_outputs(7064) <= '0';
    layer0_outputs(7065) <= not (a and b);
    layer0_outputs(7066) <= a;
    layer0_outputs(7067) <= a and b;
    layer0_outputs(7068) <= not a;
    layer0_outputs(7069) <= not (a xor b);
    layer0_outputs(7070) <= not (a and b);
    layer0_outputs(7071) <= not a;
    layer0_outputs(7072) <= a and not b;
    layer0_outputs(7073) <= b and not a;
    layer0_outputs(7074) <= not (a xor b);
    layer0_outputs(7075) <= not (a xor b);
    layer0_outputs(7076) <= not (a and b);
    layer0_outputs(7077) <= b;
    layer0_outputs(7078) <= not b or a;
    layer0_outputs(7079) <= a and b;
    layer0_outputs(7080) <= not a or b;
    layer0_outputs(7081) <= '1';
    layer0_outputs(7082) <= a;
    layer0_outputs(7083) <= a;
    layer0_outputs(7084) <= a or b;
    layer0_outputs(7085) <= not b or a;
    layer0_outputs(7086) <= not b or a;
    layer0_outputs(7087) <= not a or b;
    layer0_outputs(7088) <= not b;
    layer0_outputs(7089) <= a and b;
    layer0_outputs(7090) <= not (a or b);
    layer0_outputs(7091) <= not b or a;
    layer0_outputs(7092) <= '0';
    layer0_outputs(7093) <= a;
    layer0_outputs(7094) <= a and not b;
    layer0_outputs(7095) <= not a;
    layer0_outputs(7096) <= not (a and b);
    layer0_outputs(7097) <= a and b;
    layer0_outputs(7098) <= not b or a;
    layer0_outputs(7099) <= not (a and b);
    layer0_outputs(7100) <= a xor b;
    layer0_outputs(7101) <= a and b;
    layer0_outputs(7102) <= not b or a;
    layer0_outputs(7103) <= b;
    layer0_outputs(7104) <= a;
    layer0_outputs(7105) <= not (a or b);
    layer0_outputs(7106) <= not b or a;
    layer0_outputs(7107) <= '1';
    layer0_outputs(7108) <= '1';
    layer0_outputs(7109) <= not a or b;
    layer0_outputs(7110) <= not (a or b);
    layer0_outputs(7111) <= a or b;
    layer0_outputs(7112) <= a and b;
    layer0_outputs(7113) <= a;
    layer0_outputs(7114) <= '0';
    layer0_outputs(7115) <= not b;
    layer0_outputs(7116) <= not a or b;
    layer0_outputs(7117) <= a and not b;
    layer0_outputs(7118) <= not (a xor b);
    layer0_outputs(7119) <= not b;
    layer0_outputs(7120) <= b;
    layer0_outputs(7121) <= not (a and b);
    layer0_outputs(7122) <= not b;
    layer0_outputs(7123) <= not (a and b);
    layer0_outputs(7124) <= a xor b;
    layer0_outputs(7125) <= a and not b;
    layer0_outputs(7126) <= not a or b;
    layer0_outputs(7127) <= b;
    layer0_outputs(7128) <= not b;
    layer0_outputs(7129) <= not (a xor b);
    layer0_outputs(7130) <= a and b;
    layer0_outputs(7131) <= not (a or b);
    layer0_outputs(7132) <= not b or a;
    layer0_outputs(7133) <= not (a and b);
    layer0_outputs(7134) <= a;
    layer0_outputs(7135) <= '1';
    layer0_outputs(7136) <= '0';
    layer0_outputs(7137) <= b and not a;
    layer0_outputs(7138) <= not (a xor b);
    layer0_outputs(7139) <= a;
    layer0_outputs(7140) <= a or b;
    layer0_outputs(7141) <= a or b;
    layer0_outputs(7142) <= a;
    layer0_outputs(7143) <= a and b;
    layer0_outputs(7144) <= not b;
    layer0_outputs(7145) <= a;
    layer0_outputs(7146) <= not (a or b);
    layer0_outputs(7147) <= not a or b;
    layer0_outputs(7148) <= '1';
    layer0_outputs(7149) <= b;
    layer0_outputs(7150) <= '1';
    layer0_outputs(7151) <= a or b;
    layer0_outputs(7152) <= not (a and b);
    layer0_outputs(7153) <= '0';
    layer0_outputs(7154) <= '1';
    layer0_outputs(7155) <= not a or b;
    layer0_outputs(7156) <= not a or b;
    layer0_outputs(7157) <= a;
    layer0_outputs(7158) <= not a or b;
    layer0_outputs(7159) <= not b;
    layer0_outputs(7160) <= b and not a;
    layer0_outputs(7161) <= a;
    layer0_outputs(7162) <= not a;
    layer0_outputs(7163) <= a xor b;
    layer0_outputs(7164) <= b and not a;
    layer0_outputs(7165) <= '1';
    layer0_outputs(7166) <= not b;
    layer0_outputs(7167) <= a xor b;
    layer0_outputs(7168) <= a and not b;
    layer0_outputs(7169) <= '1';
    layer0_outputs(7170) <= '1';
    layer0_outputs(7171) <= not (a and b);
    layer0_outputs(7172) <= b;
    layer0_outputs(7173) <= not a or b;
    layer0_outputs(7174) <= not a or b;
    layer0_outputs(7175) <= not b;
    layer0_outputs(7176) <= not b or a;
    layer0_outputs(7177) <= b and not a;
    layer0_outputs(7178) <= not a or b;
    layer0_outputs(7179) <= a and b;
    layer0_outputs(7180) <= not a;
    layer0_outputs(7181) <= not (a and b);
    layer0_outputs(7182) <= not (a xor b);
    layer0_outputs(7183) <= b and not a;
    layer0_outputs(7184) <= a and b;
    layer0_outputs(7185) <= '0';
    layer0_outputs(7186) <= not b or a;
    layer0_outputs(7187) <= not a;
    layer0_outputs(7188) <= not b;
    layer0_outputs(7189) <= a or b;
    layer0_outputs(7190) <= a or b;
    layer0_outputs(7191) <= a;
    layer0_outputs(7192) <= not b;
    layer0_outputs(7193) <= not a;
    layer0_outputs(7194) <= '1';
    layer0_outputs(7195) <= not (a and b);
    layer0_outputs(7196) <= b;
    layer0_outputs(7197) <= not (a and b);
    layer0_outputs(7198) <= '0';
    layer0_outputs(7199) <= a and not b;
    layer0_outputs(7200) <= a and not b;
    layer0_outputs(7201) <= not b;
    layer0_outputs(7202) <= a and not b;
    layer0_outputs(7203) <= '1';
    layer0_outputs(7204) <= not (a or b);
    layer0_outputs(7205) <= not (a xor b);
    layer0_outputs(7206) <= a;
    layer0_outputs(7207) <= not (a or b);
    layer0_outputs(7208) <= a and b;
    layer0_outputs(7209) <= a and not b;
    layer0_outputs(7210) <= a and not b;
    layer0_outputs(7211) <= b and not a;
    layer0_outputs(7212) <= '1';
    layer0_outputs(7213) <= not (a and b);
    layer0_outputs(7214) <= '1';
    layer0_outputs(7215) <= not b;
    layer0_outputs(7216) <= not (a xor b);
    layer0_outputs(7217) <= '1';
    layer0_outputs(7218) <= a and b;
    layer0_outputs(7219) <= not a or b;
    layer0_outputs(7220) <= a;
    layer0_outputs(7221) <= not (a and b);
    layer0_outputs(7222) <= not a;
    layer0_outputs(7223) <= a xor b;
    layer0_outputs(7224) <= not a;
    layer0_outputs(7225) <= a xor b;
    layer0_outputs(7226) <= a and not b;
    layer0_outputs(7227) <= not a or b;
    layer0_outputs(7228) <= a;
    layer0_outputs(7229) <= not b or a;
    layer0_outputs(7230) <= a xor b;
    layer0_outputs(7231) <= not b or a;
    layer0_outputs(7232) <= b and not a;
    layer0_outputs(7233) <= a and b;
    layer0_outputs(7234) <= a and not b;
    layer0_outputs(7235) <= b and not a;
    layer0_outputs(7236) <= not (a and b);
    layer0_outputs(7237) <= not b or a;
    layer0_outputs(7238) <= not a or b;
    layer0_outputs(7239) <= not b;
    layer0_outputs(7240) <= a;
    layer0_outputs(7241) <= a;
    layer0_outputs(7242) <= not (a and b);
    layer0_outputs(7243) <= not b;
    layer0_outputs(7244) <= a;
    layer0_outputs(7245) <= not a;
    layer0_outputs(7246) <= not a;
    layer0_outputs(7247) <= b and not a;
    layer0_outputs(7248) <= not a;
    layer0_outputs(7249) <= a;
    layer0_outputs(7250) <= a xor b;
    layer0_outputs(7251) <= a;
    layer0_outputs(7252) <= b;
    layer0_outputs(7253) <= a and b;
    layer0_outputs(7254) <= a;
    layer0_outputs(7255) <= '1';
    layer0_outputs(7256) <= not a or b;
    layer0_outputs(7257) <= a xor b;
    layer0_outputs(7258) <= b;
    layer0_outputs(7259) <= not b or a;
    layer0_outputs(7260) <= '1';
    layer0_outputs(7261) <= '0';
    layer0_outputs(7262) <= '0';
    layer0_outputs(7263) <= not (a and b);
    layer0_outputs(7264) <= '0';
    layer0_outputs(7265) <= not a or b;
    layer0_outputs(7266) <= a;
    layer0_outputs(7267) <= not (a and b);
    layer0_outputs(7268) <= not a or b;
    layer0_outputs(7269) <= not (a xor b);
    layer0_outputs(7270) <= '0';
    layer0_outputs(7271) <= not a;
    layer0_outputs(7272) <= not a or b;
    layer0_outputs(7273) <= not (a or b);
    layer0_outputs(7274) <= not a or b;
    layer0_outputs(7275) <= not b;
    layer0_outputs(7276) <= a;
    layer0_outputs(7277) <= not b or a;
    layer0_outputs(7278) <= not (a or b);
    layer0_outputs(7279) <= not b;
    layer0_outputs(7280) <= a;
    layer0_outputs(7281) <= '0';
    layer0_outputs(7282) <= b;
    layer0_outputs(7283) <= not b;
    layer0_outputs(7284) <= b and not a;
    layer0_outputs(7285) <= '0';
    layer0_outputs(7286) <= not a;
    layer0_outputs(7287) <= not a or b;
    layer0_outputs(7288) <= not (a xor b);
    layer0_outputs(7289) <= '1';
    layer0_outputs(7290) <= b and not a;
    layer0_outputs(7291) <= not a;
    layer0_outputs(7292) <= a and b;
    layer0_outputs(7293) <= '1';
    layer0_outputs(7294) <= not (a or b);
    layer0_outputs(7295) <= a or b;
    layer0_outputs(7296) <= a or b;
    layer0_outputs(7297) <= not a or b;
    layer0_outputs(7298) <= not (a or b);
    layer0_outputs(7299) <= b and not a;
    layer0_outputs(7300) <= not (a or b);
    layer0_outputs(7301) <= not (a xor b);
    layer0_outputs(7302) <= '0';
    layer0_outputs(7303) <= not b;
    layer0_outputs(7304) <= b and not a;
    layer0_outputs(7305) <= b;
    layer0_outputs(7306) <= not (a or b);
    layer0_outputs(7307) <= a and not b;
    layer0_outputs(7308) <= a and b;
    layer0_outputs(7309) <= a and not b;
    layer0_outputs(7310) <= a and not b;
    layer0_outputs(7311) <= not (a or b);
    layer0_outputs(7312) <= '0';
    layer0_outputs(7313) <= '1';
    layer0_outputs(7314) <= '0';
    layer0_outputs(7315) <= a;
    layer0_outputs(7316) <= a or b;
    layer0_outputs(7317) <= not (a or b);
    layer0_outputs(7318) <= a or b;
    layer0_outputs(7319) <= not (a and b);
    layer0_outputs(7320) <= not a;
    layer0_outputs(7321) <= not b;
    layer0_outputs(7322) <= not a or b;
    layer0_outputs(7323) <= a or b;
    layer0_outputs(7324) <= b;
    layer0_outputs(7325) <= not (a or b);
    layer0_outputs(7326) <= not a;
    layer0_outputs(7327) <= not (a or b);
    layer0_outputs(7328) <= not a or b;
    layer0_outputs(7329) <= a and b;
    layer0_outputs(7330) <= a;
    layer0_outputs(7331) <= a and b;
    layer0_outputs(7332) <= '1';
    layer0_outputs(7333) <= a and b;
    layer0_outputs(7334) <= b and not a;
    layer0_outputs(7335) <= b and not a;
    layer0_outputs(7336) <= a;
    layer0_outputs(7337) <= not a;
    layer0_outputs(7338) <= not a;
    layer0_outputs(7339) <= '0';
    layer0_outputs(7340) <= a;
    layer0_outputs(7341) <= a;
    layer0_outputs(7342) <= a or b;
    layer0_outputs(7343) <= a xor b;
    layer0_outputs(7344) <= a and b;
    layer0_outputs(7345) <= b;
    layer0_outputs(7346) <= not b or a;
    layer0_outputs(7347) <= '0';
    layer0_outputs(7348) <= not a or b;
    layer0_outputs(7349) <= a and b;
    layer0_outputs(7350) <= not a or b;
    layer0_outputs(7351) <= not b;
    layer0_outputs(7352) <= not (a or b);
    layer0_outputs(7353) <= not a or b;
    layer0_outputs(7354) <= '0';
    layer0_outputs(7355) <= not b;
    layer0_outputs(7356) <= a and b;
    layer0_outputs(7357) <= a;
    layer0_outputs(7358) <= a;
    layer0_outputs(7359) <= not (a or b);
    layer0_outputs(7360) <= '0';
    layer0_outputs(7361) <= b and not a;
    layer0_outputs(7362) <= a xor b;
    layer0_outputs(7363) <= a;
    layer0_outputs(7364) <= not b or a;
    layer0_outputs(7365) <= '0';
    layer0_outputs(7366) <= not b or a;
    layer0_outputs(7367) <= not a or b;
    layer0_outputs(7368) <= not b;
    layer0_outputs(7369) <= '0';
    layer0_outputs(7370) <= b and not a;
    layer0_outputs(7371) <= '1';
    layer0_outputs(7372) <= a;
    layer0_outputs(7373) <= '1';
    layer0_outputs(7374) <= a or b;
    layer0_outputs(7375) <= b;
    layer0_outputs(7376) <= not b;
    layer0_outputs(7377) <= a and not b;
    layer0_outputs(7378) <= '1';
    layer0_outputs(7379) <= not b;
    layer0_outputs(7380) <= a;
    layer0_outputs(7381) <= not (a and b);
    layer0_outputs(7382) <= '0';
    layer0_outputs(7383) <= a and not b;
    layer0_outputs(7384) <= a;
    layer0_outputs(7385) <= not (a xor b);
    layer0_outputs(7386) <= not b or a;
    layer0_outputs(7387) <= not b;
    layer0_outputs(7388) <= a;
    layer0_outputs(7389) <= b;
    layer0_outputs(7390) <= not (a or b);
    layer0_outputs(7391) <= not a or b;
    layer0_outputs(7392) <= '1';
    layer0_outputs(7393) <= a or b;
    layer0_outputs(7394) <= not a or b;
    layer0_outputs(7395) <= a and b;
    layer0_outputs(7396) <= a and b;
    layer0_outputs(7397) <= not (a and b);
    layer0_outputs(7398) <= a;
    layer0_outputs(7399) <= not a;
    layer0_outputs(7400) <= not a or b;
    layer0_outputs(7401) <= a;
    layer0_outputs(7402) <= b;
    layer0_outputs(7403) <= a and not b;
    layer0_outputs(7404) <= not (a xor b);
    layer0_outputs(7405) <= not (a or b);
    layer0_outputs(7406) <= not b;
    layer0_outputs(7407) <= not a or b;
    layer0_outputs(7408) <= '0';
    layer0_outputs(7409) <= a or b;
    layer0_outputs(7410) <= a and not b;
    layer0_outputs(7411) <= a and b;
    layer0_outputs(7412) <= not a;
    layer0_outputs(7413) <= a and not b;
    layer0_outputs(7414) <= not (a or b);
    layer0_outputs(7415) <= '1';
    layer0_outputs(7416) <= not (a xor b);
    layer0_outputs(7417) <= b;
    layer0_outputs(7418) <= '1';
    layer0_outputs(7419) <= a;
    layer0_outputs(7420) <= not b;
    layer0_outputs(7421) <= not (a or b);
    layer0_outputs(7422) <= b and not a;
    layer0_outputs(7423) <= not a;
    layer0_outputs(7424) <= '1';
    layer0_outputs(7425) <= not (a or b);
    layer0_outputs(7426) <= not a;
    layer0_outputs(7427) <= a and not b;
    layer0_outputs(7428) <= not a or b;
    layer0_outputs(7429) <= '1';
    layer0_outputs(7430) <= a xor b;
    layer0_outputs(7431) <= a xor b;
    layer0_outputs(7432) <= '1';
    layer0_outputs(7433) <= '0';
    layer0_outputs(7434) <= '0';
    layer0_outputs(7435) <= not b or a;
    layer0_outputs(7436) <= a or b;
    layer0_outputs(7437) <= a;
    layer0_outputs(7438) <= '0';
    layer0_outputs(7439) <= a or b;
    layer0_outputs(7440) <= b;
    layer0_outputs(7441) <= a xor b;
    layer0_outputs(7442) <= '1';
    layer0_outputs(7443) <= not a or b;
    layer0_outputs(7444) <= a and b;
    layer0_outputs(7445) <= not b;
    layer0_outputs(7446) <= '1';
    layer0_outputs(7447) <= a and b;
    layer0_outputs(7448) <= not (a or b);
    layer0_outputs(7449) <= a;
    layer0_outputs(7450) <= '1';
    layer0_outputs(7451) <= b;
    layer0_outputs(7452) <= not b;
    layer0_outputs(7453) <= not b;
    layer0_outputs(7454) <= a and b;
    layer0_outputs(7455) <= a and b;
    layer0_outputs(7456) <= b and not a;
    layer0_outputs(7457) <= a;
    layer0_outputs(7458) <= b and not a;
    layer0_outputs(7459) <= not b;
    layer0_outputs(7460) <= b and not a;
    layer0_outputs(7461) <= a;
    layer0_outputs(7462) <= b;
    layer0_outputs(7463) <= not (a xor b);
    layer0_outputs(7464) <= b and not a;
    layer0_outputs(7465) <= '0';
    layer0_outputs(7466) <= a or b;
    layer0_outputs(7467) <= a and b;
    layer0_outputs(7468) <= a or b;
    layer0_outputs(7469) <= a xor b;
    layer0_outputs(7470) <= not (a or b);
    layer0_outputs(7471) <= not (a or b);
    layer0_outputs(7472) <= '0';
    layer0_outputs(7473) <= not b;
    layer0_outputs(7474) <= '0';
    layer0_outputs(7475) <= b and not a;
    layer0_outputs(7476) <= a and b;
    layer0_outputs(7477) <= b;
    layer0_outputs(7478) <= not (a or b);
    layer0_outputs(7479) <= not (a and b);
    layer0_outputs(7480) <= a;
    layer0_outputs(7481) <= not a;
    layer0_outputs(7482) <= b;
    layer0_outputs(7483) <= not b;
    layer0_outputs(7484) <= not (a or b);
    layer0_outputs(7485) <= b;
    layer0_outputs(7486) <= a;
    layer0_outputs(7487) <= not b or a;
    layer0_outputs(7488) <= not (a and b);
    layer0_outputs(7489) <= b;
    layer0_outputs(7490) <= not b or a;
    layer0_outputs(7491) <= not (a or b);
    layer0_outputs(7492) <= not a or b;
    layer0_outputs(7493) <= not a or b;
    layer0_outputs(7494) <= not b;
    layer0_outputs(7495) <= not (a and b);
    layer0_outputs(7496) <= a and b;
    layer0_outputs(7497) <= not b;
    layer0_outputs(7498) <= a or b;
    layer0_outputs(7499) <= a and b;
    layer0_outputs(7500) <= a;
    layer0_outputs(7501) <= b and not a;
    layer0_outputs(7502) <= a;
    layer0_outputs(7503) <= '1';
    layer0_outputs(7504) <= a or b;
    layer0_outputs(7505) <= '1';
    layer0_outputs(7506) <= '1';
    layer0_outputs(7507) <= a or b;
    layer0_outputs(7508) <= not b;
    layer0_outputs(7509) <= a xor b;
    layer0_outputs(7510) <= '1';
    layer0_outputs(7511) <= not a or b;
    layer0_outputs(7512) <= not b or a;
    layer0_outputs(7513) <= not a;
    layer0_outputs(7514) <= a and not b;
    layer0_outputs(7515) <= '1';
    layer0_outputs(7516) <= not a or b;
    layer0_outputs(7517) <= b and not a;
    layer0_outputs(7518) <= b and not a;
    layer0_outputs(7519) <= '1';
    layer0_outputs(7520) <= b and not a;
    layer0_outputs(7521) <= a or b;
    layer0_outputs(7522) <= a xor b;
    layer0_outputs(7523) <= '1';
    layer0_outputs(7524) <= not a;
    layer0_outputs(7525) <= a or b;
    layer0_outputs(7526) <= not a;
    layer0_outputs(7527) <= '0';
    layer0_outputs(7528) <= not (a xor b);
    layer0_outputs(7529) <= '0';
    layer0_outputs(7530) <= not b;
    layer0_outputs(7531) <= not (a or b);
    layer0_outputs(7532) <= '1';
    layer0_outputs(7533) <= not a;
    layer0_outputs(7534) <= not (a and b);
    layer0_outputs(7535) <= not (a or b);
    layer0_outputs(7536) <= a or b;
    layer0_outputs(7537) <= b and not a;
    layer0_outputs(7538) <= not a;
    layer0_outputs(7539) <= not (a or b);
    layer0_outputs(7540) <= b;
    layer0_outputs(7541) <= not a;
    layer0_outputs(7542) <= a and not b;
    layer0_outputs(7543) <= '1';
    layer0_outputs(7544) <= a and not b;
    layer0_outputs(7545) <= b;
    layer0_outputs(7546) <= not (a xor b);
    layer0_outputs(7547) <= a or b;
    layer0_outputs(7548) <= a and not b;
    layer0_outputs(7549) <= not b or a;
    layer0_outputs(7550) <= '0';
    layer0_outputs(7551) <= a;
    layer0_outputs(7552) <= not (a and b);
    layer0_outputs(7553) <= a and not b;
    layer0_outputs(7554) <= b and not a;
    layer0_outputs(7555) <= a;
    layer0_outputs(7556) <= not a;
    layer0_outputs(7557) <= not (a xor b);
    layer0_outputs(7558) <= not (a or b);
    layer0_outputs(7559) <= b and not a;
    layer0_outputs(7560) <= '1';
    layer0_outputs(7561) <= a and not b;
    layer0_outputs(7562) <= not a;
    layer0_outputs(7563) <= not a or b;
    layer0_outputs(7564) <= '0';
    layer0_outputs(7565) <= '0';
    layer0_outputs(7566) <= a and not b;
    layer0_outputs(7567) <= '0';
    layer0_outputs(7568) <= not (a and b);
    layer0_outputs(7569) <= '1';
    layer0_outputs(7570) <= b and not a;
    layer0_outputs(7571) <= not b;
    layer0_outputs(7572) <= not a;
    layer0_outputs(7573) <= not a;
    layer0_outputs(7574) <= not b;
    layer0_outputs(7575) <= not (a xor b);
    layer0_outputs(7576) <= a and b;
    layer0_outputs(7577) <= a or b;
    layer0_outputs(7578) <= a or b;
    layer0_outputs(7579) <= '0';
    layer0_outputs(7580) <= a and not b;
    layer0_outputs(7581) <= a xor b;
    layer0_outputs(7582) <= not (a xor b);
    layer0_outputs(7583) <= not b or a;
    layer0_outputs(7584) <= b and not a;
    layer0_outputs(7585) <= not b;
    layer0_outputs(7586) <= not (a or b);
    layer0_outputs(7587) <= not b or a;
    layer0_outputs(7588) <= a or b;
    layer0_outputs(7589) <= b and not a;
    layer0_outputs(7590) <= not (a xor b);
    layer0_outputs(7591) <= '1';
    layer0_outputs(7592) <= not a or b;
    layer0_outputs(7593) <= a and not b;
    layer0_outputs(7594) <= b;
    layer0_outputs(7595) <= a and not b;
    layer0_outputs(7596) <= a;
    layer0_outputs(7597) <= not b;
    layer0_outputs(7598) <= a xor b;
    layer0_outputs(7599) <= not b;
    layer0_outputs(7600) <= a and b;
    layer0_outputs(7601) <= a;
    layer0_outputs(7602) <= a or b;
    layer0_outputs(7603) <= not a or b;
    layer0_outputs(7604) <= b;
    layer0_outputs(7605) <= not a;
    layer0_outputs(7606) <= not a or b;
    layer0_outputs(7607) <= b and not a;
    layer0_outputs(7608) <= '1';
    layer0_outputs(7609) <= not (a or b);
    layer0_outputs(7610) <= not (a or b);
    layer0_outputs(7611) <= not (a xor b);
    layer0_outputs(7612) <= not a;
    layer0_outputs(7613) <= b;
    layer0_outputs(7614) <= a;
    layer0_outputs(7615) <= not (a and b);
    layer0_outputs(7616) <= not b;
    layer0_outputs(7617) <= b;
    layer0_outputs(7618) <= a and not b;
    layer0_outputs(7619) <= not (a and b);
    layer0_outputs(7620) <= a xor b;
    layer0_outputs(7621) <= a or b;
    layer0_outputs(7622) <= not a;
    layer0_outputs(7623) <= not b;
    layer0_outputs(7624) <= a;
    layer0_outputs(7625) <= not a or b;
    layer0_outputs(7626) <= not (a and b);
    layer0_outputs(7627) <= a and not b;
    layer0_outputs(7628) <= '1';
    layer0_outputs(7629) <= b;
    layer0_outputs(7630) <= not (a and b);
    layer0_outputs(7631) <= a or b;
    layer0_outputs(7632) <= not b or a;
    layer0_outputs(7633) <= a and b;
    layer0_outputs(7634) <= not (a or b);
    layer0_outputs(7635) <= b;
    layer0_outputs(7636) <= b and not a;
    layer0_outputs(7637) <= a and not b;
    layer0_outputs(7638) <= not a or b;
    layer0_outputs(7639) <= not (a xor b);
    layer0_outputs(7640) <= not b or a;
    layer0_outputs(7641) <= not (a and b);
    layer0_outputs(7642) <= a xor b;
    layer0_outputs(7643) <= '1';
    layer0_outputs(7644) <= '1';
    layer0_outputs(7645) <= b;
    layer0_outputs(7646) <= a and not b;
    layer0_outputs(7647) <= not b;
    layer0_outputs(7648) <= b and not a;
    layer0_outputs(7649) <= not (a and b);
    layer0_outputs(7650) <= not a;
    layer0_outputs(7651) <= '0';
    layer0_outputs(7652) <= not b or a;
    layer0_outputs(7653) <= not a or b;
    layer0_outputs(7654) <= '0';
    layer0_outputs(7655) <= not (a or b);
    layer0_outputs(7656) <= not b;
    layer0_outputs(7657) <= a and not b;
    layer0_outputs(7658) <= b;
    layer0_outputs(7659) <= '0';
    layer0_outputs(7660) <= a;
    layer0_outputs(7661) <= a and b;
    layer0_outputs(7662) <= a xor b;
    layer0_outputs(7663) <= not a;
    layer0_outputs(7664) <= not (a and b);
    layer0_outputs(7665) <= a or b;
    layer0_outputs(7666) <= '0';
    layer0_outputs(7667) <= a and b;
    layer0_outputs(7668) <= b and not a;
    layer0_outputs(7669) <= not a;
    layer0_outputs(7670) <= not b;
    layer0_outputs(7671) <= not (a and b);
    layer0_outputs(7672) <= a or b;
    layer0_outputs(7673) <= not b;
    layer0_outputs(7674) <= not a or b;
    layer0_outputs(7675) <= a xor b;
    layer0_outputs(7676) <= a and b;
    layer0_outputs(7677) <= '1';
    layer0_outputs(7678) <= '1';
    layer0_outputs(7679) <= a and not b;
    layer1_outputs(0) <= a;
    layer1_outputs(1) <= not (a or b);
    layer1_outputs(2) <= b and not a;
    layer1_outputs(3) <= a and b;
    layer1_outputs(4) <= a or b;
    layer1_outputs(5) <= '0';
    layer1_outputs(6) <= not b;
    layer1_outputs(7) <= b and not a;
    layer1_outputs(8) <= '0';
    layer1_outputs(9) <= b;
    layer1_outputs(10) <= not (a or b);
    layer1_outputs(11) <= b and not a;
    layer1_outputs(12) <= '1';
    layer1_outputs(13) <= '1';
    layer1_outputs(14) <= not (a or b);
    layer1_outputs(15) <= a and not b;
    layer1_outputs(16) <= not (a or b);
    layer1_outputs(17) <= a and not b;
    layer1_outputs(18) <= not a;
    layer1_outputs(19) <= a and b;
    layer1_outputs(20) <= a;
    layer1_outputs(21) <= not (a or b);
    layer1_outputs(22) <= '1';
    layer1_outputs(23) <= not (a or b);
    layer1_outputs(24) <= b and not a;
    layer1_outputs(25) <= not a;
    layer1_outputs(26) <= a or b;
    layer1_outputs(27) <= not b or a;
    layer1_outputs(28) <= a or b;
    layer1_outputs(29) <= a or b;
    layer1_outputs(30) <= a;
    layer1_outputs(31) <= '0';
    layer1_outputs(32) <= b and not a;
    layer1_outputs(33) <= not (a or b);
    layer1_outputs(34) <= not b or a;
    layer1_outputs(35) <= a;
    layer1_outputs(36) <= a and b;
    layer1_outputs(37) <= a and not b;
    layer1_outputs(38) <= b and not a;
    layer1_outputs(39) <= not a or b;
    layer1_outputs(40) <= '1';
    layer1_outputs(41) <= not (a or b);
    layer1_outputs(42) <= not b or a;
    layer1_outputs(43) <= a and b;
    layer1_outputs(44) <= '1';
    layer1_outputs(45) <= not (a and b);
    layer1_outputs(46) <= not (a xor b);
    layer1_outputs(47) <= a or b;
    layer1_outputs(48) <= not (a and b);
    layer1_outputs(49) <= a and not b;
    layer1_outputs(50) <= '1';
    layer1_outputs(51) <= not b;
    layer1_outputs(52) <= a;
    layer1_outputs(53) <= a;
    layer1_outputs(54) <= not b;
    layer1_outputs(55) <= not a;
    layer1_outputs(56) <= a xor b;
    layer1_outputs(57) <= b and not a;
    layer1_outputs(58) <= a xor b;
    layer1_outputs(59) <= a xor b;
    layer1_outputs(60) <= b and not a;
    layer1_outputs(61) <= a and b;
    layer1_outputs(62) <= not (a or b);
    layer1_outputs(63) <= not a;
    layer1_outputs(64) <= b;
    layer1_outputs(65) <= not a;
    layer1_outputs(66) <= b;
    layer1_outputs(67) <= not b;
    layer1_outputs(68) <= not a or b;
    layer1_outputs(69) <= not a;
    layer1_outputs(70) <= a and b;
    layer1_outputs(71) <= '0';
    layer1_outputs(72) <= '0';
    layer1_outputs(73) <= not b or a;
    layer1_outputs(74) <= not (a or b);
    layer1_outputs(75) <= '0';
    layer1_outputs(76) <= not (a and b);
    layer1_outputs(77) <= b;
    layer1_outputs(78) <= a and not b;
    layer1_outputs(79) <= not a or b;
    layer1_outputs(80) <= a and b;
    layer1_outputs(81) <= a or b;
    layer1_outputs(82) <= '1';
    layer1_outputs(83) <= not (a and b);
    layer1_outputs(84) <= not a or b;
    layer1_outputs(85) <= not b;
    layer1_outputs(86) <= '0';
    layer1_outputs(87) <= '1';
    layer1_outputs(88) <= b and not a;
    layer1_outputs(89) <= not (a or b);
    layer1_outputs(90) <= a and b;
    layer1_outputs(91) <= b;
    layer1_outputs(92) <= not (a xor b);
    layer1_outputs(93) <= a and b;
    layer1_outputs(94) <= b;
    layer1_outputs(95) <= not b;
    layer1_outputs(96) <= b and not a;
    layer1_outputs(97) <= not b;
    layer1_outputs(98) <= a and not b;
    layer1_outputs(99) <= not b or a;
    layer1_outputs(100) <= a or b;
    layer1_outputs(101) <= b;
    layer1_outputs(102) <= not a or b;
    layer1_outputs(103) <= a and b;
    layer1_outputs(104) <= not a or b;
    layer1_outputs(105) <= not b or a;
    layer1_outputs(106) <= not a or b;
    layer1_outputs(107) <= not a or b;
    layer1_outputs(108) <= a xor b;
    layer1_outputs(109) <= '1';
    layer1_outputs(110) <= a and b;
    layer1_outputs(111) <= '1';
    layer1_outputs(112) <= not (a or b);
    layer1_outputs(113) <= b and not a;
    layer1_outputs(114) <= b and not a;
    layer1_outputs(115) <= not b or a;
    layer1_outputs(116) <= b;
    layer1_outputs(117) <= b;
    layer1_outputs(118) <= b and not a;
    layer1_outputs(119) <= '1';
    layer1_outputs(120) <= a and b;
    layer1_outputs(121) <= not b or a;
    layer1_outputs(122) <= not (a or b);
    layer1_outputs(123) <= not a;
    layer1_outputs(124) <= b and not a;
    layer1_outputs(125) <= b;
    layer1_outputs(126) <= a and not b;
    layer1_outputs(127) <= not a;
    layer1_outputs(128) <= a and not b;
    layer1_outputs(129) <= b and not a;
    layer1_outputs(130) <= b;
    layer1_outputs(131) <= not (a xor b);
    layer1_outputs(132) <= not a;
    layer1_outputs(133) <= not (a and b);
    layer1_outputs(134) <= a xor b;
    layer1_outputs(135) <= not (a and b);
    layer1_outputs(136) <= '0';
    layer1_outputs(137) <= a and b;
    layer1_outputs(138) <= '1';
    layer1_outputs(139) <= not a or b;
    layer1_outputs(140) <= not (a or b);
    layer1_outputs(141) <= not (a or b);
    layer1_outputs(142) <= '0';
    layer1_outputs(143) <= '1';
    layer1_outputs(144) <= not b;
    layer1_outputs(145) <= a;
    layer1_outputs(146) <= '1';
    layer1_outputs(147) <= not (a or b);
    layer1_outputs(148) <= not a;
    layer1_outputs(149) <= b;
    layer1_outputs(150) <= a or b;
    layer1_outputs(151) <= not b or a;
    layer1_outputs(152) <= b;
    layer1_outputs(153) <= not (a and b);
    layer1_outputs(154) <= not b or a;
    layer1_outputs(155) <= a and not b;
    layer1_outputs(156) <= not (a and b);
    layer1_outputs(157) <= a;
    layer1_outputs(158) <= a or b;
    layer1_outputs(159) <= a and not b;
    layer1_outputs(160) <= not b or a;
    layer1_outputs(161) <= '1';
    layer1_outputs(162) <= not a or b;
    layer1_outputs(163) <= a and b;
    layer1_outputs(164) <= not (a and b);
    layer1_outputs(165) <= not (a and b);
    layer1_outputs(166) <= a or b;
    layer1_outputs(167) <= '1';
    layer1_outputs(168) <= not a;
    layer1_outputs(169) <= b and not a;
    layer1_outputs(170) <= a and not b;
    layer1_outputs(171) <= b;
    layer1_outputs(172) <= a xor b;
    layer1_outputs(173) <= not b or a;
    layer1_outputs(174) <= '0';
    layer1_outputs(175) <= a xor b;
    layer1_outputs(176) <= not a;
    layer1_outputs(177) <= a;
    layer1_outputs(178) <= a or b;
    layer1_outputs(179) <= not (a and b);
    layer1_outputs(180) <= a and not b;
    layer1_outputs(181) <= a or b;
    layer1_outputs(182) <= not b;
    layer1_outputs(183) <= a xor b;
    layer1_outputs(184) <= b;
    layer1_outputs(185) <= a or b;
    layer1_outputs(186) <= not a;
    layer1_outputs(187) <= not a;
    layer1_outputs(188) <= not b;
    layer1_outputs(189) <= not (a and b);
    layer1_outputs(190) <= not (a and b);
    layer1_outputs(191) <= not (a and b);
    layer1_outputs(192) <= b and not a;
    layer1_outputs(193) <= a;
    layer1_outputs(194) <= '0';
    layer1_outputs(195) <= not b or a;
    layer1_outputs(196) <= not (a xor b);
    layer1_outputs(197) <= not (a or b);
    layer1_outputs(198) <= b and not a;
    layer1_outputs(199) <= not b;
    layer1_outputs(200) <= not (a and b);
    layer1_outputs(201) <= a or b;
    layer1_outputs(202) <= not (a and b);
    layer1_outputs(203) <= not a;
    layer1_outputs(204) <= not a or b;
    layer1_outputs(205) <= not b or a;
    layer1_outputs(206) <= not b or a;
    layer1_outputs(207) <= b;
    layer1_outputs(208) <= a xor b;
    layer1_outputs(209) <= not a;
    layer1_outputs(210) <= not a or b;
    layer1_outputs(211) <= a or b;
    layer1_outputs(212) <= '1';
    layer1_outputs(213) <= a;
    layer1_outputs(214) <= b;
    layer1_outputs(215) <= b;
    layer1_outputs(216) <= not a or b;
    layer1_outputs(217) <= a and b;
    layer1_outputs(218) <= b and not a;
    layer1_outputs(219) <= '0';
    layer1_outputs(220) <= a and not b;
    layer1_outputs(221) <= not (a and b);
    layer1_outputs(222) <= a;
    layer1_outputs(223) <= not (a and b);
    layer1_outputs(224) <= a;
    layer1_outputs(225) <= not a;
    layer1_outputs(226) <= b and not a;
    layer1_outputs(227) <= a and not b;
    layer1_outputs(228) <= b;
    layer1_outputs(229) <= not (a and b);
    layer1_outputs(230) <= b;
    layer1_outputs(231) <= not b;
    layer1_outputs(232) <= b and not a;
    layer1_outputs(233) <= not (a xor b);
    layer1_outputs(234) <= '0';
    layer1_outputs(235) <= not b;
    layer1_outputs(236) <= not a;
    layer1_outputs(237) <= not b;
    layer1_outputs(238) <= not b or a;
    layer1_outputs(239) <= not (a and b);
    layer1_outputs(240) <= not b;
    layer1_outputs(241) <= b and not a;
    layer1_outputs(242) <= not (a xor b);
    layer1_outputs(243) <= not b;
    layer1_outputs(244) <= not a;
    layer1_outputs(245) <= not b;
    layer1_outputs(246) <= not b;
    layer1_outputs(247) <= not a;
    layer1_outputs(248) <= not (a and b);
    layer1_outputs(249) <= a and not b;
    layer1_outputs(250) <= '0';
    layer1_outputs(251) <= a;
    layer1_outputs(252) <= b;
    layer1_outputs(253) <= not a;
    layer1_outputs(254) <= not (a and b);
    layer1_outputs(255) <= b and not a;
    layer1_outputs(256) <= b and not a;
    layer1_outputs(257) <= '0';
    layer1_outputs(258) <= '1';
    layer1_outputs(259) <= b and not a;
    layer1_outputs(260) <= not b;
    layer1_outputs(261) <= '1';
    layer1_outputs(262) <= a and not b;
    layer1_outputs(263) <= '0';
    layer1_outputs(264) <= a or b;
    layer1_outputs(265) <= b;
    layer1_outputs(266) <= '0';
    layer1_outputs(267) <= a;
    layer1_outputs(268) <= not (a or b);
    layer1_outputs(269) <= not a;
    layer1_outputs(270) <= not (a xor b);
    layer1_outputs(271) <= b;
    layer1_outputs(272) <= b;
    layer1_outputs(273) <= not (a or b);
    layer1_outputs(274) <= a;
    layer1_outputs(275) <= a or b;
    layer1_outputs(276) <= '0';
    layer1_outputs(277) <= b and not a;
    layer1_outputs(278) <= not b;
    layer1_outputs(279) <= a and b;
    layer1_outputs(280) <= '0';
    layer1_outputs(281) <= '1';
    layer1_outputs(282) <= a and not b;
    layer1_outputs(283) <= a;
    layer1_outputs(284) <= not a or b;
    layer1_outputs(285) <= a and not b;
    layer1_outputs(286) <= not (a or b);
    layer1_outputs(287) <= a and not b;
    layer1_outputs(288) <= not b;
    layer1_outputs(289) <= not a;
    layer1_outputs(290) <= a;
    layer1_outputs(291) <= '0';
    layer1_outputs(292) <= not (a xor b);
    layer1_outputs(293) <= not (a or b);
    layer1_outputs(294) <= not (a and b);
    layer1_outputs(295) <= '0';
    layer1_outputs(296) <= not b or a;
    layer1_outputs(297) <= b;
    layer1_outputs(298) <= not a;
    layer1_outputs(299) <= not (a xor b);
    layer1_outputs(300) <= '1';
    layer1_outputs(301) <= not (a and b);
    layer1_outputs(302) <= '0';
    layer1_outputs(303) <= not a;
    layer1_outputs(304) <= b and not a;
    layer1_outputs(305) <= a and b;
    layer1_outputs(306) <= not a or b;
    layer1_outputs(307) <= not (a or b);
    layer1_outputs(308) <= a and b;
    layer1_outputs(309) <= a and b;
    layer1_outputs(310) <= not (a and b);
    layer1_outputs(311) <= a;
    layer1_outputs(312) <= not (a or b);
    layer1_outputs(313) <= '0';
    layer1_outputs(314) <= not (a and b);
    layer1_outputs(315) <= a;
    layer1_outputs(316) <= a or b;
    layer1_outputs(317) <= not a;
    layer1_outputs(318) <= not a;
    layer1_outputs(319) <= a and not b;
    layer1_outputs(320) <= '1';
    layer1_outputs(321) <= not (a or b);
    layer1_outputs(322) <= a xor b;
    layer1_outputs(323) <= not b;
    layer1_outputs(324) <= not b or a;
    layer1_outputs(325) <= not (a and b);
    layer1_outputs(326) <= a;
    layer1_outputs(327) <= a or b;
    layer1_outputs(328) <= a and not b;
    layer1_outputs(329) <= a and not b;
    layer1_outputs(330) <= a;
    layer1_outputs(331) <= not (a and b);
    layer1_outputs(332) <= a xor b;
    layer1_outputs(333) <= a;
    layer1_outputs(334) <= not a;
    layer1_outputs(335) <= '1';
    layer1_outputs(336) <= a or b;
    layer1_outputs(337) <= '0';
    layer1_outputs(338) <= '1';
    layer1_outputs(339) <= b and not a;
    layer1_outputs(340) <= b;
    layer1_outputs(341) <= a and not b;
    layer1_outputs(342) <= not b;
    layer1_outputs(343) <= b;
    layer1_outputs(344) <= not b or a;
    layer1_outputs(345) <= a xor b;
    layer1_outputs(346) <= not (a and b);
    layer1_outputs(347) <= a or b;
    layer1_outputs(348) <= a and not b;
    layer1_outputs(349) <= not (a or b);
    layer1_outputs(350) <= '0';
    layer1_outputs(351) <= a and b;
    layer1_outputs(352) <= not a or b;
    layer1_outputs(353) <= '0';
    layer1_outputs(354) <= not (a or b);
    layer1_outputs(355) <= not (a and b);
    layer1_outputs(356) <= a xor b;
    layer1_outputs(357) <= not a;
    layer1_outputs(358) <= a xor b;
    layer1_outputs(359) <= a or b;
    layer1_outputs(360) <= '1';
    layer1_outputs(361) <= not (a and b);
    layer1_outputs(362) <= b and not a;
    layer1_outputs(363) <= not b or a;
    layer1_outputs(364) <= '1';
    layer1_outputs(365) <= not (a xor b);
    layer1_outputs(366) <= not a or b;
    layer1_outputs(367) <= b;
    layer1_outputs(368) <= b and not a;
    layer1_outputs(369) <= '1';
    layer1_outputs(370) <= '0';
    layer1_outputs(371) <= not (a or b);
    layer1_outputs(372) <= a or b;
    layer1_outputs(373) <= not (a xor b);
    layer1_outputs(374) <= a;
    layer1_outputs(375) <= b;
    layer1_outputs(376) <= b and not a;
    layer1_outputs(377) <= a or b;
    layer1_outputs(378) <= a or b;
    layer1_outputs(379) <= not a or b;
    layer1_outputs(380) <= not (a or b);
    layer1_outputs(381) <= not b or a;
    layer1_outputs(382) <= a and not b;
    layer1_outputs(383) <= a or b;
    layer1_outputs(384) <= b;
    layer1_outputs(385) <= not (a or b);
    layer1_outputs(386) <= not b;
    layer1_outputs(387) <= b;
    layer1_outputs(388) <= not (a or b);
    layer1_outputs(389) <= a xor b;
    layer1_outputs(390) <= '1';
    layer1_outputs(391) <= '0';
    layer1_outputs(392) <= '0';
    layer1_outputs(393) <= a or b;
    layer1_outputs(394) <= not a or b;
    layer1_outputs(395) <= not (a and b);
    layer1_outputs(396) <= b;
    layer1_outputs(397) <= '0';
    layer1_outputs(398) <= a or b;
    layer1_outputs(399) <= a and b;
    layer1_outputs(400) <= b and not a;
    layer1_outputs(401) <= not b;
    layer1_outputs(402) <= not (a or b);
    layer1_outputs(403) <= '1';
    layer1_outputs(404) <= a xor b;
    layer1_outputs(405) <= '0';
    layer1_outputs(406) <= not b;
    layer1_outputs(407) <= not (a xor b);
    layer1_outputs(408) <= a and not b;
    layer1_outputs(409) <= b;
    layer1_outputs(410) <= a or b;
    layer1_outputs(411) <= not (a or b);
    layer1_outputs(412) <= not (a or b);
    layer1_outputs(413) <= a;
    layer1_outputs(414) <= not a or b;
    layer1_outputs(415) <= a and not b;
    layer1_outputs(416) <= not b;
    layer1_outputs(417) <= '0';
    layer1_outputs(418) <= b;
    layer1_outputs(419) <= not (a and b);
    layer1_outputs(420) <= not (a xor b);
    layer1_outputs(421) <= not (a or b);
    layer1_outputs(422) <= '0';
    layer1_outputs(423) <= b and not a;
    layer1_outputs(424) <= b;
    layer1_outputs(425) <= a and not b;
    layer1_outputs(426) <= b;
    layer1_outputs(427) <= a;
    layer1_outputs(428) <= not (a or b);
    layer1_outputs(429) <= not b;
    layer1_outputs(430) <= not a;
    layer1_outputs(431) <= b and not a;
    layer1_outputs(432) <= '1';
    layer1_outputs(433) <= b and not a;
    layer1_outputs(434) <= b and not a;
    layer1_outputs(435) <= not a;
    layer1_outputs(436) <= not a;
    layer1_outputs(437) <= not (a and b);
    layer1_outputs(438) <= a;
    layer1_outputs(439) <= a or b;
    layer1_outputs(440) <= not a or b;
    layer1_outputs(441) <= '0';
    layer1_outputs(442) <= not a;
    layer1_outputs(443) <= not a;
    layer1_outputs(444) <= a or b;
    layer1_outputs(445) <= b;
    layer1_outputs(446) <= b;
    layer1_outputs(447) <= not b;
    layer1_outputs(448) <= '1';
    layer1_outputs(449) <= not a;
    layer1_outputs(450) <= b;
    layer1_outputs(451) <= a or b;
    layer1_outputs(452) <= not a or b;
    layer1_outputs(453) <= not a;
    layer1_outputs(454) <= not a or b;
    layer1_outputs(455) <= b and not a;
    layer1_outputs(456) <= '1';
    layer1_outputs(457) <= b and not a;
    layer1_outputs(458) <= b;
    layer1_outputs(459) <= '0';
    layer1_outputs(460) <= '1';
    layer1_outputs(461) <= '0';
    layer1_outputs(462) <= not (a and b);
    layer1_outputs(463) <= not a or b;
    layer1_outputs(464) <= not b;
    layer1_outputs(465) <= not a or b;
    layer1_outputs(466) <= not (a or b);
    layer1_outputs(467) <= '0';
    layer1_outputs(468) <= not b or a;
    layer1_outputs(469) <= not (a xor b);
    layer1_outputs(470) <= b and not a;
    layer1_outputs(471) <= a or b;
    layer1_outputs(472) <= not a or b;
    layer1_outputs(473) <= b;
    layer1_outputs(474) <= not (a or b);
    layer1_outputs(475) <= b;
    layer1_outputs(476) <= not a;
    layer1_outputs(477) <= not (a and b);
    layer1_outputs(478) <= '1';
    layer1_outputs(479) <= '1';
    layer1_outputs(480) <= '0';
    layer1_outputs(481) <= not a;
    layer1_outputs(482) <= not (a and b);
    layer1_outputs(483) <= '0';
    layer1_outputs(484) <= b;
    layer1_outputs(485) <= b;
    layer1_outputs(486) <= a and not b;
    layer1_outputs(487) <= a and not b;
    layer1_outputs(488) <= b and not a;
    layer1_outputs(489) <= a or b;
    layer1_outputs(490) <= '0';
    layer1_outputs(491) <= not a or b;
    layer1_outputs(492) <= not a or b;
    layer1_outputs(493) <= '1';
    layer1_outputs(494) <= a and b;
    layer1_outputs(495) <= a and not b;
    layer1_outputs(496) <= a xor b;
    layer1_outputs(497) <= '1';
    layer1_outputs(498) <= not (a or b);
    layer1_outputs(499) <= a and not b;
    layer1_outputs(500) <= not (a and b);
    layer1_outputs(501) <= not (a and b);
    layer1_outputs(502) <= b;
    layer1_outputs(503) <= not b or a;
    layer1_outputs(504) <= a;
    layer1_outputs(505) <= '0';
    layer1_outputs(506) <= not a or b;
    layer1_outputs(507) <= a and not b;
    layer1_outputs(508) <= not b or a;
    layer1_outputs(509) <= not b or a;
    layer1_outputs(510) <= not b;
    layer1_outputs(511) <= a and not b;
    layer1_outputs(512) <= not a;
    layer1_outputs(513) <= b;
    layer1_outputs(514) <= not (a xor b);
    layer1_outputs(515) <= '0';
    layer1_outputs(516) <= a;
    layer1_outputs(517) <= '0';
    layer1_outputs(518) <= not a;
    layer1_outputs(519) <= not a or b;
    layer1_outputs(520) <= not (a or b);
    layer1_outputs(521) <= a or b;
    layer1_outputs(522) <= '1';
    layer1_outputs(523) <= b and not a;
    layer1_outputs(524) <= not (a and b);
    layer1_outputs(525) <= not b;
    layer1_outputs(526) <= not b;
    layer1_outputs(527) <= a;
    layer1_outputs(528) <= not b or a;
    layer1_outputs(529) <= a and b;
    layer1_outputs(530) <= b and not a;
    layer1_outputs(531) <= not (a or b);
    layer1_outputs(532) <= b;
    layer1_outputs(533) <= not a or b;
    layer1_outputs(534) <= a and b;
    layer1_outputs(535) <= not (a and b);
    layer1_outputs(536) <= not (a and b);
    layer1_outputs(537) <= b;
    layer1_outputs(538) <= not a;
    layer1_outputs(539) <= b and not a;
    layer1_outputs(540) <= b and not a;
    layer1_outputs(541) <= '0';
    layer1_outputs(542) <= not b or a;
    layer1_outputs(543) <= not b;
    layer1_outputs(544) <= not (a and b);
    layer1_outputs(545) <= b and not a;
    layer1_outputs(546) <= b;
    layer1_outputs(547) <= not b;
    layer1_outputs(548) <= '0';
    layer1_outputs(549) <= not (a or b);
    layer1_outputs(550) <= not (a xor b);
    layer1_outputs(551) <= not (a or b);
    layer1_outputs(552) <= not a;
    layer1_outputs(553) <= not (a xor b);
    layer1_outputs(554) <= b and not a;
    layer1_outputs(555) <= b and not a;
    layer1_outputs(556) <= not (a xor b);
    layer1_outputs(557) <= not (a xor b);
    layer1_outputs(558) <= '0';
    layer1_outputs(559) <= not a;
    layer1_outputs(560) <= b and not a;
    layer1_outputs(561) <= not b;
    layer1_outputs(562) <= not b;
    layer1_outputs(563) <= '0';
    layer1_outputs(564) <= a or b;
    layer1_outputs(565) <= not a;
    layer1_outputs(566) <= not (a xor b);
    layer1_outputs(567) <= '0';
    layer1_outputs(568) <= not b or a;
    layer1_outputs(569) <= a and b;
    layer1_outputs(570) <= a and b;
    layer1_outputs(571) <= '1';
    layer1_outputs(572) <= a and b;
    layer1_outputs(573) <= b;
    layer1_outputs(574) <= a and not b;
    layer1_outputs(575) <= '1';
    layer1_outputs(576) <= not a or b;
    layer1_outputs(577) <= '0';
    layer1_outputs(578) <= not b;
    layer1_outputs(579) <= '0';
    layer1_outputs(580) <= not a or b;
    layer1_outputs(581) <= not (a xor b);
    layer1_outputs(582) <= not a or b;
    layer1_outputs(583) <= a;
    layer1_outputs(584) <= '1';
    layer1_outputs(585) <= not (a and b);
    layer1_outputs(586) <= not a;
    layer1_outputs(587) <= not a or b;
    layer1_outputs(588) <= not b;
    layer1_outputs(589) <= not b;
    layer1_outputs(590) <= '1';
    layer1_outputs(591) <= not (a or b);
    layer1_outputs(592) <= not b;
    layer1_outputs(593) <= a;
    layer1_outputs(594) <= not b or a;
    layer1_outputs(595) <= not b;
    layer1_outputs(596) <= '1';
    layer1_outputs(597) <= a;
    layer1_outputs(598) <= a and b;
    layer1_outputs(599) <= not b;
    layer1_outputs(600) <= not a;
    layer1_outputs(601) <= a and b;
    layer1_outputs(602) <= not a;
    layer1_outputs(603) <= not b or a;
    layer1_outputs(604) <= not a or b;
    layer1_outputs(605) <= b;
    layer1_outputs(606) <= not b or a;
    layer1_outputs(607) <= not (a and b);
    layer1_outputs(608) <= not b;
    layer1_outputs(609) <= a and not b;
    layer1_outputs(610) <= not b or a;
    layer1_outputs(611) <= a or b;
    layer1_outputs(612) <= a and b;
    layer1_outputs(613) <= not b;
    layer1_outputs(614) <= '1';
    layer1_outputs(615) <= '1';
    layer1_outputs(616) <= a;
    layer1_outputs(617) <= a and not b;
    layer1_outputs(618) <= b and not a;
    layer1_outputs(619) <= not b or a;
    layer1_outputs(620) <= not a or b;
    layer1_outputs(621) <= a and not b;
    layer1_outputs(622) <= b and not a;
    layer1_outputs(623) <= b and not a;
    layer1_outputs(624) <= not a or b;
    layer1_outputs(625) <= a or b;
    layer1_outputs(626) <= not (a or b);
    layer1_outputs(627) <= not (a or b);
    layer1_outputs(628) <= a and b;
    layer1_outputs(629) <= b and not a;
    layer1_outputs(630) <= not b or a;
    layer1_outputs(631) <= not a;
    layer1_outputs(632) <= not a;
    layer1_outputs(633) <= '0';
    layer1_outputs(634) <= a and not b;
    layer1_outputs(635) <= a or b;
    layer1_outputs(636) <= b and not a;
    layer1_outputs(637) <= not (a xor b);
    layer1_outputs(638) <= b;
    layer1_outputs(639) <= not a or b;
    layer1_outputs(640) <= '0';
    layer1_outputs(641) <= not b;
    layer1_outputs(642) <= a or b;
    layer1_outputs(643) <= b and not a;
    layer1_outputs(644) <= a xor b;
    layer1_outputs(645) <= b and not a;
    layer1_outputs(646) <= '0';
    layer1_outputs(647) <= not b;
    layer1_outputs(648) <= a and not b;
    layer1_outputs(649) <= a and b;
    layer1_outputs(650) <= not (a or b);
    layer1_outputs(651) <= not (a or b);
    layer1_outputs(652) <= not (a and b);
    layer1_outputs(653) <= '1';
    layer1_outputs(654) <= not b or a;
    layer1_outputs(655) <= not a or b;
    layer1_outputs(656) <= a;
    layer1_outputs(657) <= a xor b;
    layer1_outputs(658) <= not a;
    layer1_outputs(659) <= '0';
    layer1_outputs(660) <= not b;
    layer1_outputs(661) <= a;
    layer1_outputs(662) <= a and not b;
    layer1_outputs(663) <= not a;
    layer1_outputs(664) <= a xor b;
    layer1_outputs(665) <= not (a and b);
    layer1_outputs(666) <= a or b;
    layer1_outputs(667) <= '0';
    layer1_outputs(668) <= '1';
    layer1_outputs(669) <= not b;
    layer1_outputs(670) <= not a or b;
    layer1_outputs(671) <= b and not a;
    layer1_outputs(672) <= '1';
    layer1_outputs(673) <= not (a and b);
    layer1_outputs(674) <= not (a xor b);
    layer1_outputs(675) <= not (a xor b);
    layer1_outputs(676) <= not (a xor b);
    layer1_outputs(677) <= not (a xor b);
    layer1_outputs(678) <= '0';
    layer1_outputs(679) <= not b or a;
    layer1_outputs(680) <= not (a or b);
    layer1_outputs(681) <= not (a or b);
    layer1_outputs(682) <= not b or a;
    layer1_outputs(683) <= a or b;
    layer1_outputs(684) <= not (a or b);
    layer1_outputs(685) <= a xor b;
    layer1_outputs(686) <= not b;
    layer1_outputs(687) <= b;
    layer1_outputs(688) <= not b;
    layer1_outputs(689) <= not (a or b);
    layer1_outputs(690) <= not (a or b);
    layer1_outputs(691) <= b;
    layer1_outputs(692) <= '0';
    layer1_outputs(693) <= '0';
    layer1_outputs(694) <= '0';
    layer1_outputs(695) <= a and b;
    layer1_outputs(696) <= '0';
    layer1_outputs(697) <= '1';
    layer1_outputs(698) <= b;
    layer1_outputs(699) <= not b or a;
    layer1_outputs(700) <= not (a and b);
    layer1_outputs(701) <= not b or a;
    layer1_outputs(702) <= not b;
    layer1_outputs(703) <= b and not a;
    layer1_outputs(704) <= not a;
    layer1_outputs(705) <= not b;
    layer1_outputs(706) <= not (a xor b);
    layer1_outputs(707) <= '0';
    layer1_outputs(708) <= b and not a;
    layer1_outputs(709) <= not b or a;
    layer1_outputs(710) <= '0';
    layer1_outputs(711) <= not b;
    layer1_outputs(712) <= a and not b;
    layer1_outputs(713) <= b;
    layer1_outputs(714) <= '1';
    layer1_outputs(715) <= '0';
    layer1_outputs(716) <= b;
    layer1_outputs(717) <= not (a xor b);
    layer1_outputs(718) <= a and b;
    layer1_outputs(719) <= not a or b;
    layer1_outputs(720) <= not a or b;
    layer1_outputs(721) <= '1';
    layer1_outputs(722) <= a or b;
    layer1_outputs(723) <= not (a xor b);
    layer1_outputs(724) <= not b or a;
    layer1_outputs(725) <= '0';
    layer1_outputs(726) <= a;
    layer1_outputs(727) <= b and not a;
    layer1_outputs(728) <= '0';
    layer1_outputs(729) <= not (a and b);
    layer1_outputs(730) <= not a or b;
    layer1_outputs(731) <= not b;
    layer1_outputs(732) <= not (a and b);
    layer1_outputs(733) <= a;
    layer1_outputs(734) <= a;
    layer1_outputs(735) <= not (a or b);
    layer1_outputs(736) <= not (a or b);
    layer1_outputs(737) <= a or b;
    layer1_outputs(738) <= not a;
    layer1_outputs(739) <= a and b;
    layer1_outputs(740) <= not a or b;
    layer1_outputs(741) <= not b;
    layer1_outputs(742) <= a or b;
    layer1_outputs(743) <= b;
    layer1_outputs(744) <= '0';
    layer1_outputs(745) <= not a;
    layer1_outputs(746) <= not a;
    layer1_outputs(747) <= not b;
    layer1_outputs(748) <= not a or b;
    layer1_outputs(749) <= a and b;
    layer1_outputs(750) <= b and not a;
    layer1_outputs(751) <= not a;
    layer1_outputs(752) <= '1';
    layer1_outputs(753) <= a or b;
    layer1_outputs(754) <= b and not a;
    layer1_outputs(755) <= a xor b;
    layer1_outputs(756) <= not (a xor b);
    layer1_outputs(757) <= not a;
    layer1_outputs(758) <= not a or b;
    layer1_outputs(759) <= not (a and b);
    layer1_outputs(760) <= not b;
    layer1_outputs(761) <= a;
    layer1_outputs(762) <= not b or a;
    layer1_outputs(763) <= not b or a;
    layer1_outputs(764) <= not a or b;
    layer1_outputs(765) <= a;
    layer1_outputs(766) <= not (a and b);
    layer1_outputs(767) <= a;
    layer1_outputs(768) <= not b;
    layer1_outputs(769) <= b and not a;
    layer1_outputs(770) <= '0';
    layer1_outputs(771) <= not (a and b);
    layer1_outputs(772) <= a;
    layer1_outputs(773) <= not a;
    layer1_outputs(774) <= a;
    layer1_outputs(775) <= not (a and b);
    layer1_outputs(776) <= '1';
    layer1_outputs(777) <= not a or b;
    layer1_outputs(778) <= not b;
    layer1_outputs(779) <= a or b;
    layer1_outputs(780) <= not (a or b);
    layer1_outputs(781) <= not a;
    layer1_outputs(782) <= b and not a;
    layer1_outputs(783) <= not (a and b);
    layer1_outputs(784) <= b and not a;
    layer1_outputs(785) <= not a;
    layer1_outputs(786) <= not a;
    layer1_outputs(787) <= '1';
    layer1_outputs(788) <= not (a and b);
    layer1_outputs(789) <= b;
    layer1_outputs(790) <= a xor b;
    layer1_outputs(791) <= b and not a;
    layer1_outputs(792) <= not a or b;
    layer1_outputs(793) <= '1';
    layer1_outputs(794) <= b;
    layer1_outputs(795) <= not a;
    layer1_outputs(796) <= not a;
    layer1_outputs(797) <= a;
    layer1_outputs(798) <= b and not a;
    layer1_outputs(799) <= not (a or b);
    layer1_outputs(800) <= b;
    layer1_outputs(801) <= not a;
    layer1_outputs(802) <= a xor b;
    layer1_outputs(803) <= not a;
    layer1_outputs(804) <= not (a or b);
    layer1_outputs(805) <= '0';
    layer1_outputs(806) <= not b or a;
    layer1_outputs(807) <= a and not b;
    layer1_outputs(808) <= a or b;
    layer1_outputs(809) <= not b;
    layer1_outputs(810) <= not b;
    layer1_outputs(811) <= not (a xor b);
    layer1_outputs(812) <= '1';
    layer1_outputs(813) <= not a or b;
    layer1_outputs(814) <= b and not a;
    layer1_outputs(815) <= a and not b;
    layer1_outputs(816) <= not (a and b);
    layer1_outputs(817) <= a xor b;
    layer1_outputs(818) <= not a;
    layer1_outputs(819) <= b;
    layer1_outputs(820) <= not (a and b);
    layer1_outputs(821) <= '1';
    layer1_outputs(822) <= b and not a;
    layer1_outputs(823) <= not a or b;
    layer1_outputs(824) <= b and not a;
    layer1_outputs(825) <= a and not b;
    layer1_outputs(826) <= not a;
    layer1_outputs(827) <= not a or b;
    layer1_outputs(828) <= not a;
    layer1_outputs(829) <= not a or b;
    layer1_outputs(830) <= not b;
    layer1_outputs(831) <= '0';
    layer1_outputs(832) <= '1';
    layer1_outputs(833) <= '0';
    layer1_outputs(834) <= not a;
    layer1_outputs(835) <= a or b;
    layer1_outputs(836) <= b;
    layer1_outputs(837) <= not b or a;
    layer1_outputs(838) <= not a or b;
    layer1_outputs(839) <= a;
    layer1_outputs(840) <= '1';
    layer1_outputs(841) <= not (a xor b);
    layer1_outputs(842) <= not a or b;
    layer1_outputs(843) <= a and b;
    layer1_outputs(844) <= not a;
    layer1_outputs(845) <= a and not b;
    layer1_outputs(846) <= '0';
    layer1_outputs(847) <= a and b;
    layer1_outputs(848) <= a or b;
    layer1_outputs(849) <= a or b;
    layer1_outputs(850) <= '0';
    layer1_outputs(851) <= a and not b;
    layer1_outputs(852) <= a and not b;
    layer1_outputs(853) <= a and not b;
    layer1_outputs(854) <= '0';
    layer1_outputs(855) <= b;
    layer1_outputs(856) <= not (a or b);
    layer1_outputs(857) <= '1';
    layer1_outputs(858) <= b and not a;
    layer1_outputs(859) <= not b or a;
    layer1_outputs(860) <= a and not b;
    layer1_outputs(861) <= not b or a;
    layer1_outputs(862) <= not (a and b);
    layer1_outputs(863) <= a and b;
    layer1_outputs(864) <= a and b;
    layer1_outputs(865) <= a and b;
    layer1_outputs(866) <= a;
    layer1_outputs(867) <= a and not b;
    layer1_outputs(868) <= b and not a;
    layer1_outputs(869) <= b;
    layer1_outputs(870) <= a and b;
    layer1_outputs(871) <= not b or a;
    layer1_outputs(872) <= '1';
    layer1_outputs(873) <= '0';
    layer1_outputs(874) <= a and b;
    layer1_outputs(875) <= not b or a;
    layer1_outputs(876) <= a and b;
    layer1_outputs(877) <= not (a and b);
    layer1_outputs(878) <= not a or b;
    layer1_outputs(879) <= b and not a;
    layer1_outputs(880) <= '1';
    layer1_outputs(881) <= '0';
    layer1_outputs(882) <= a or b;
    layer1_outputs(883) <= a or b;
    layer1_outputs(884) <= a and b;
    layer1_outputs(885) <= b and not a;
    layer1_outputs(886) <= a and b;
    layer1_outputs(887) <= not a or b;
    layer1_outputs(888) <= not b or a;
    layer1_outputs(889) <= not b or a;
    layer1_outputs(890) <= not a or b;
    layer1_outputs(891) <= a and not b;
    layer1_outputs(892) <= a or b;
    layer1_outputs(893) <= not a or b;
    layer1_outputs(894) <= a and not b;
    layer1_outputs(895) <= not b;
    layer1_outputs(896) <= not a;
    layer1_outputs(897) <= not (a xor b);
    layer1_outputs(898) <= not b;
    layer1_outputs(899) <= not (a or b);
    layer1_outputs(900) <= not a;
    layer1_outputs(901) <= a and b;
    layer1_outputs(902) <= a and not b;
    layer1_outputs(903) <= not a;
    layer1_outputs(904) <= a or b;
    layer1_outputs(905) <= a or b;
    layer1_outputs(906) <= not a;
    layer1_outputs(907) <= not b or a;
    layer1_outputs(908) <= not b or a;
    layer1_outputs(909) <= a and not b;
    layer1_outputs(910) <= '1';
    layer1_outputs(911) <= not (a or b);
    layer1_outputs(912) <= a and not b;
    layer1_outputs(913) <= not b or a;
    layer1_outputs(914) <= '0';
    layer1_outputs(915) <= a and b;
    layer1_outputs(916) <= a and b;
    layer1_outputs(917) <= a or b;
    layer1_outputs(918) <= not b;
    layer1_outputs(919) <= b;
    layer1_outputs(920) <= not b or a;
    layer1_outputs(921) <= not a or b;
    layer1_outputs(922) <= a and not b;
    layer1_outputs(923) <= not a;
    layer1_outputs(924) <= not a or b;
    layer1_outputs(925) <= b;
    layer1_outputs(926) <= not a or b;
    layer1_outputs(927) <= not (a or b);
    layer1_outputs(928) <= not (a and b);
    layer1_outputs(929) <= a xor b;
    layer1_outputs(930) <= not (a and b);
    layer1_outputs(931) <= a;
    layer1_outputs(932) <= not b;
    layer1_outputs(933) <= a or b;
    layer1_outputs(934) <= b;
    layer1_outputs(935) <= not (a or b);
    layer1_outputs(936) <= not b;
    layer1_outputs(937) <= a and not b;
    layer1_outputs(938) <= '0';
    layer1_outputs(939) <= not b;
    layer1_outputs(940) <= not b or a;
    layer1_outputs(941) <= a;
    layer1_outputs(942) <= not a;
    layer1_outputs(943) <= not (a or b);
    layer1_outputs(944) <= not (a or b);
    layer1_outputs(945) <= a xor b;
    layer1_outputs(946) <= not (a and b);
    layer1_outputs(947) <= not a;
    layer1_outputs(948) <= a or b;
    layer1_outputs(949) <= a or b;
    layer1_outputs(950) <= a and not b;
    layer1_outputs(951) <= not b;
    layer1_outputs(952) <= not b or a;
    layer1_outputs(953) <= '1';
    layer1_outputs(954) <= b;
    layer1_outputs(955) <= not a or b;
    layer1_outputs(956) <= a;
    layer1_outputs(957) <= '1';
    layer1_outputs(958) <= a and not b;
    layer1_outputs(959) <= not b;
    layer1_outputs(960) <= not (a or b);
    layer1_outputs(961) <= '1';
    layer1_outputs(962) <= '1';
    layer1_outputs(963) <= a and b;
    layer1_outputs(964) <= not b;
    layer1_outputs(965) <= not (a xor b);
    layer1_outputs(966) <= not (a or b);
    layer1_outputs(967) <= not a or b;
    layer1_outputs(968) <= b and not a;
    layer1_outputs(969) <= not (a xor b);
    layer1_outputs(970) <= not a or b;
    layer1_outputs(971) <= not (a and b);
    layer1_outputs(972) <= not (a and b);
    layer1_outputs(973) <= b;
    layer1_outputs(974) <= not (a and b);
    layer1_outputs(975) <= a;
    layer1_outputs(976) <= b and not a;
    layer1_outputs(977) <= not a;
    layer1_outputs(978) <= a;
    layer1_outputs(979) <= '0';
    layer1_outputs(980) <= a;
    layer1_outputs(981) <= not b or a;
    layer1_outputs(982) <= a;
    layer1_outputs(983) <= b;
    layer1_outputs(984) <= not (a xor b);
    layer1_outputs(985) <= b;
    layer1_outputs(986) <= not a or b;
    layer1_outputs(987) <= a and not b;
    layer1_outputs(988) <= not (a or b);
    layer1_outputs(989) <= '0';
    layer1_outputs(990) <= not b;
    layer1_outputs(991) <= '0';
    layer1_outputs(992) <= not (a and b);
    layer1_outputs(993) <= a and not b;
    layer1_outputs(994) <= a and b;
    layer1_outputs(995) <= a and not b;
    layer1_outputs(996) <= not a;
    layer1_outputs(997) <= b;
    layer1_outputs(998) <= not a or b;
    layer1_outputs(999) <= not a;
    layer1_outputs(1000) <= a and b;
    layer1_outputs(1001) <= b and not a;
    layer1_outputs(1002) <= not (a or b);
    layer1_outputs(1003) <= a and b;
    layer1_outputs(1004) <= not (a or b);
    layer1_outputs(1005) <= '1';
    layer1_outputs(1006) <= b;
    layer1_outputs(1007) <= a;
    layer1_outputs(1008) <= a xor b;
    layer1_outputs(1009) <= a and not b;
    layer1_outputs(1010) <= not b or a;
    layer1_outputs(1011) <= '1';
    layer1_outputs(1012) <= b;
    layer1_outputs(1013) <= '0';
    layer1_outputs(1014) <= not a or b;
    layer1_outputs(1015) <= not b;
    layer1_outputs(1016) <= a;
    layer1_outputs(1017) <= not b;
    layer1_outputs(1018) <= b and not a;
    layer1_outputs(1019) <= b and not a;
    layer1_outputs(1020) <= not (a or b);
    layer1_outputs(1021) <= a or b;
    layer1_outputs(1022) <= not a or b;
    layer1_outputs(1023) <= not b or a;
    layer1_outputs(1024) <= b;
    layer1_outputs(1025) <= not a;
    layer1_outputs(1026) <= not a;
    layer1_outputs(1027) <= a and not b;
    layer1_outputs(1028) <= '1';
    layer1_outputs(1029) <= a or b;
    layer1_outputs(1030) <= not (a or b);
    layer1_outputs(1031) <= not (a xor b);
    layer1_outputs(1032) <= a xor b;
    layer1_outputs(1033) <= a and b;
    layer1_outputs(1034) <= a and not b;
    layer1_outputs(1035) <= not b or a;
    layer1_outputs(1036) <= '1';
    layer1_outputs(1037) <= a and b;
    layer1_outputs(1038) <= a or b;
    layer1_outputs(1039) <= a;
    layer1_outputs(1040) <= a;
    layer1_outputs(1041) <= a and b;
    layer1_outputs(1042) <= a;
    layer1_outputs(1043) <= not b or a;
    layer1_outputs(1044) <= not (a or b);
    layer1_outputs(1045) <= '1';
    layer1_outputs(1046) <= b and not a;
    layer1_outputs(1047) <= not (a or b);
    layer1_outputs(1048) <= a and b;
    layer1_outputs(1049) <= b and not a;
    layer1_outputs(1050) <= a;
    layer1_outputs(1051) <= '1';
    layer1_outputs(1052) <= not (a and b);
    layer1_outputs(1053) <= a;
    layer1_outputs(1054) <= '0';
    layer1_outputs(1055) <= not a or b;
    layer1_outputs(1056) <= not b;
    layer1_outputs(1057) <= not a;
    layer1_outputs(1058) <= a;
    layer1_outputs(1059) <= not (a and b);
    layer1_outputs(1060) <= '1';
    layer1_outputs(1061) <= '0';
    layer1_outputs(1062) <= a;
    layer1_outputs(1063) <= not a or b;
    layer1_outputs(1064) <= '0';
    layer1_outputs(1065) <= a or b;
    layer1_outputs(1066) <= not (a and b);
    layer1_outputs(1067) <= '1';
    layer1_outputs(1068) <= not (a xor b);
    layer1_outputs(1069) <= b;
    layer1_outputs(1070) <= b;
    layer1_outputs(1071) <= not a or b;
    layer1_outputs(1072) <= not a;
    layer1_outputs(1073) <= a and b;
    layer1_outputs(1074) <= not (a or b);
    layer1_outputs(1075) <= '1';
    layer1_outputs(1076) <= a and not b;
    layer1_outputs(1077) <= not (a or b);
    layer1_outputs(1078) <= '0';
    layer1_outputs(1079) <= not (a and b);
    layer1_outputs(1080) <= b;
    layer1_outputs(1081) <= not (a xor b);
    layer1_outputs(1082) <= a or b;
    layer1_outputs(1083) <= '0';
    layer1_outputs(1084) <= not b;
    layer1_outputs(1085) <= not (a and b);
    layer1_outputs(1086) <= not a;
    layer1_outputs(1087) <= a or b;
    layer1_outputs(1088) <= a;
    layer1_outputs(1089) <= not (a xor b);
    layer1_outputs(1090) <= a;
    layer1_outputs(1091) <= a;
    layer1_outputs(1092) <= a;
    layer1_outputs(1093) <= not (a or b);
    layer1_outputs(1094) <= not a;
    layer1_outputs(1095) <= not b or a;
    layer1_outputs(1096) <= not (a or b);
    layer1_outputs(1097) <= '0';
    layer1_outputs(1098) <= not a;
    layer1_outputs(1099) <= not b or a;
    layer1_outputs(1100) <= a and not b;
    layer1_outputs(1101) <= not (a or b);
    layer1_outputs(1102) <= not (a and b);
    layer1_outputs(1103) <= not (a or b);
    layer1_outputs(1104) <= b;
    layer1_outputs(1105) <= '0';
    layer1_outputs(1106) <= '1';
    layer1_outputs(1107) <= b and not a;
    layer1_outputs(1108) <= '0';
    layer1_outputs(1109) <= '0';
    layer1_outputs(1110) <= not a;
    layer1_outputs(1111) <= a and b;
    layer1_outputs(1112) <= not b or a;
    layer1_outputs(1113) <= b;
    layer1_outputs(1114) <= not a;
    layer1_outputs(1115) <= b;
    layer1_outputs(1116) <= a and not b;
    layer1_outputs(1117) <= '0';
    layer1_outputs(1118) <= not a;
    layer1_outputs(1119) <= not (a and b);
    layer1_outputs(1120) <= a and b;
    layer1_outputs(1121) <= not a;
    layer1_outputs(1122) <= not b or a;
    layer1_outputs(1123) <= a;
    layer1_outputs(1124) <= a and not b;
    layer1_outputs(1125) <= a and b;
    layer1_outputs(1126) <= a or b;
    layer1_outputs(1127) <= not b;
    layer1_outputs(1128) <= a and not b;
    layer1_outputs(1129) <= a and b;
    layer1_outputs(1130) <= '0';
    layer1_outputs(1131) <= '1';
    layer1_outputs(1132) <= a and b;
    layer1_outputs(1133) <= '1';
    layer1_outputs(1134) <= a xor b;
    layer1_outputs(1135) <= a or b;
    layer1_outputs(1136) <= not (a and b);
    layer1_outputs(1137) <= not (a or b);
    layer1_outputs(1138) <= a and b;
    layer1_outputs(1139) <= not b;
    layer1_outputs(1140) <= '1';
    layer1_outputs(1141) <= not b or a;
    layer1_outputs(1142) <= a or b;
    layer1_outputs(1143) <= not a;
    layer1_outputs(1144) <= a and b;
    layer1_outputs(1145) <= a and b;
    layer1_outputs(1146) <= '0';
    layer1_outputs(1147) <= not (a and b);
    layer1_outputs(1148) <= not (a xor b);
    layer1_outputs(1149) <= not (a or b);
    layer1_outputs(1150) <= '0';
    layer1_outputs(1151) <= b and not a;
    layer1_outputs(1152) <= not (a or b);
    layer1_outputs(1153) <= '0';
    layer1_outputs(1154) <= not (a or b);
    layer1_outputs(1155) <= not (a xor b);
    layer1_outputs(1156) <= a and b;
    layer1_outputs(1157) <= '0';
    layer1_outputs(1158) <= not a or b;
    layer1_outputs(1159) <= a or b;
    layer1_outputs(1160) <= '0';
    layer1_outputs(1161) <= not b or a;
    layer1_outputs(1162) <= a and not b;
    layer1_outputs(1163) <= b and not a;
    layer1_outputs(1164) <= b;
    layer1_outputs(1165) <= not a or b;
    layer1_outputs(1166) <= '1';
    layer1_outputs(1167) <= a and not b;
    layer1_outputs(1168) <= not b or a;
    layer1_outputs(1169) <= not b;
    layer1_outputs(1170) <= not a;
    layer1_outputs(1171) <= a and not b;
    layer1_outputs(1172) <= a or b;
    layer1_outputs(1173) <= b;
    layer1_outputs(1174) <= b and not a;
    layer1_outputs(1175) <= '1';
    layer1_outputs(1176) <= a;
    layer1_outputs(1177) <= a and not b;
    layer1_outputs(1178) <= a or b;
    layer1_outputs(1179) <= a or b;
    layer1_outputs(1180) <= a;
    layer1_outputs(1181) <= a and not b;
    layer1_outputs(1182) <= not a or b;
    layer1_outputs(1183) <= b and not a;
    layer1_outputs(1184) <= not a;
    layer1_outputs(1185) <= not b;
    layer1_outputs(1186) <= not a or b;
    layer1_outputs(1187) <= a and not b;
    layer1_outputs(1188) <= not b or a;
    layer1_outputs(1189) <= not (a or b);
    layer1_outputs(1190) <= not b;
    layer1_outputs(1191) <= '0';
    layer1_outputs(1192) <= a;
    layer1_outputs(1193) <= '0';
    layer1_outputs(1194) <= not a;
    layer1_outputs(1195) <= a;
    layer1_outputs(1196) <= b;
    layer1_outputs(1197) <= a;
    layer1_outputs(1198) <= not a or b;
    layer1_outputs(1199) <= not (a xor b);
    layer1_outputs(1200) <= not (a and b);
    layer1_outputs(1201) <= b;
    layer1_outputs(1202) <= not (a xor b);
    layer1_outputs(1203) <= '0';
    layer1_outputs(1204) <= a or b;
    layer1_outputs(1205) <= b;
    layer1_outputs(1206) <= b;
    layer1_outputs(1207) <= '0';
    layer1_outputs(1208) <= not b;
    layer1_outputs(1209) <= a;
    layer1_outputs(1210) <= '1';
    layer1_outputs(1211) <= not (a xor b);
    layer1_outputs(1212) <= b;
    layer1_outputs(1213) <= not b or a;
    layer1_outputs(1214) <= not (a and b);
    layer1_outputs(1215) <= '0';
    layer1_outputs(1216) <= not (a and b);
    layer1_outputs(1217) <= a and b;
    layer1_outputs(1218) <= b and not a;
    layer1_outputs(1219) <= a or b;
    layer1_outputs(1220) <= '0';
    layer1_outputs(1221) <= '0';
    layer1_outputs(1222) <= not (a or b);
    layer1_outputs(1223) <= not a;
    layer1_outputs(1224) <= not a or b;
    layer1_outputs(1225) <= a;
    layer1_outputs(1226) <= not (a or b);
    layer1_outputs(1227) <= not (a and b);
    layer1_outputs(1228) <= a or b;
    layer1_outputs(1229) <= not (a or b);
    layer1_outputs(1230) <= not (a and b);
    layer1_outputs(1231) <= '0';
    layer1_outputs(1232) <= not a;
    layer1_outputs(1233) <= a and b;
    layer1_outputs(1234) <= a or b;
    layer1_outputs(1235) <= not b or a;
    layer1_outputs(1236) <= not a or b;
    layer1_outputs(1237) <= not b or a;
    layer1_outputs(1238) <= not a;
    layer1_outputs(1239) <= not a or b;
    layer1_outputs(1240) <= b;
    layer1_outputs(1241) <= not (a and b);
    layer1_outputs(1242) <= not a or b;
    layer1_outputs(1243) <= a and b;
    layer1_outputs(1244) <= not b or a;
    layer1_outputs(1245) <= not a;
    layer1_outputs(1246) <= not (a and b);
    layer1_outputs(1247) <= not b or a;
    layer1_outputs(1248) <= '0';
    layer1_outputs(1249) <= not a or b;
    layer1_outputs(1250) <= a or b;
    layer1_outputs(1251) <= not b;
    layer1_outputs(1252) <= a xor b;
    layer1_outputs(1253) <= not b;
    layer1_outputs(1254) <= not a;
    layer1_outputs(1255) <= not (a and b);
    layer1_outputs(1256) <= '0';
    layer1_outputs(1257) <= not (a or b);
    layer1_outputs(1258) <= a and not b;
    layer1_outputs(1259) <= a and not b;
    layer1_outputs(1260) <= not (a and b);
    layer1_outputs(1261) <= b;
    layer1_outputs(1262) <= a and b;
    layer1_outputs(1263) <= b;
    layer1_outputs(1264) <= '1';
    layer1_outputs(1265) <= '1';
    layer1_outputs(1266) <= a;
    layer1_outputs(1267) <= not b or a;
    layer1_outputs(1268) <= '1';
    layer1_outputs(1269) <= '0';
    layer1_outputs(1270) <= a xor b;
    layer1_outputs(1271) <= not a;
    layer1_outputs(1272) <= a and b;
    layer1_outputs(1273) <= '0';
    layer1_outputs(1274) <= not a or b;
    layer1_outputs(1275) <= not b or a;
    layer1_outputs(1276) <= b;
    layer1_outputs(1277) <= '0';
    layer1_outputs(1278) <= not b;
    layer1_outputs(1279) <= '0';
    layer1_outputs(1280) <= a or b;
    layer1_outputs(1281) <= not (a and b);
    layer1_outputs(1282) <= not b or a;
    layer1_outputs(1283) <= a;
    layer1_outputs(1284) <= a;
    layer1_outputs(1285) <= not (a xor b);
    layer1_outputs(1286) <= b;
    layer1_outputs(1287) <= a and b;
    layer1_outputs(1288) <= not b or a;
    layer1_outputs(1289) <= '1';
    layer1_outputs(1290) <= not a or b;
    layer1_outputs(1291) <= a and b;
    layer1_outputs(1292) <= a and not b;
    layer1_outputs(1293) <= '0';
    layer1_outputs(1294) <= not (a and b);
    layer1_outputs(1295) <= not (a and b);
    layer1_outputs(1296) <= not a or b;
    layer1_outputs(1297) <= not b;
    layer1_outputs(1298) <= b;
    layer1_outputs(1299) <= a;
    layer1_outputs(1300) <= not a or b;
    layer1_outputs(1301) <= a and b;
    layer1_outputs(1302) <= b;
    layer1_outputs(1303) <= a and b;
    layer1_outputs(1304) <= '1';
    layer1_outputs(1305) <= b and not a;
    layer1_outputs(1306) <= b and not a;
    layer1_outputs(1307) <= not b or a;
    layer1_outputs(1308) <= b;
    layer1_outputs(1309) <= a and not b;
    layer1_outputs(1310) <= not b or a;
    layer1_outputs(1311) <= not (a and b);
    layer1_outputs(1312) <= b;
    layer1_outputs(1313) <= '1';
    layer1_outputs(1314) <= not a or b;
    layer1_outputs(1315) <= a;
    layer1_outputs(1316) <= a and b;
    layer1_outputs(1317) <= a or b;
    layer1_outputs(1318) <= a xor b;
    layer1_outputs(1319) <= '0';
    layer1_outputs(1320) <= b;
    layer1_outputs(1321) <= a xor b;
    layer1_outputs(1322) <= a and b;
    layer1_outputs(1323) <= '0';
    layer1_outputs(1324) <= '1';
    layer1_outputs(1325) <= not a or b;
    layer1_outputs(1326) <= a xor b;
    layer1_outputs(1327) <= not b;
    layer1_outputs(1328) <= a and not b;
    layer1_outputs(1329) <= not b;
    layer1_outputs(1330) <= '0';
    layer1_outputs(1331) <= a or b;
    layer1_outputs(1332) <= '1';
    layer1_outputs(1333) <= not (a or b);
    layer1_outputs(1334) <= not b or a;
    layer1_outputs(1335) <= b;
    layer1_outputs(1336) <= a;
    layer1_outputs(1337) <= a and not b;
    layer1_outputs(1338) <= '0';
    layer1_outputs(1339) <= b and not a;
    layer1_outputs(1340) <= not b or a;
    layer1_outputs(1341) <= not a or b;
    layer1_outputs(1342) <= a;
    layer1_outputs(1343) <= a and b;
    layer1_outputs(1344) <= b;
    layer1_outputs(1345) <= '1';
    layer1_outputs(1346) <= not (a xor b);
    layer1_outputs(1347) <= a and b;
    layer1_outputs(1348) <= not a;
    layer1_outputs(1349) <= a or b;
    layer1_outputs(1350) <= not (a and b);
    layer1_outputs(1351) <= not (a and b);
    layer1_outputs(1352) <= not (a and b);
    layer1_outputs(1353) <= not a or b;
    layer1_outputs(1354) <= not (a or b);
    layer1_outputs(1355) <= not b or a;
    layer1_outputs(1356) <= a xor b;
    layer1_outputs(1357) <= a or b;
    layer1_outputs(1358) <= not b;
    layer1_outputs(1359) <= not a or b;
    layer1_outputs(1360) <= not a or b;
    layer1_outputs(1361) <= a;
    layer1_outputs(1362) <= b;
    layer1_outputs(1363) <= a or b;
    layer1_outputs(1364) <= b;
    layer1_outputs(1365) <= a;
    layer1_outputs(1366) <= a and b;
    layer1_outputs(1367) <= '1';
    layer1_outputs(1368) <= '0';
    layer1_outputs(1369) <= '0';
    layer1_outputs(1370) <= b;
    layer1_outputs(1371) <= a and b;
    layer1_outputs(1372) <= b;
    layer1_outputs(1373) <= b;
    layer1_outputs(1374) <= b;
    layer1_outputs(1375) <= not (a or b);
    layer1_outputs(1376) <= a or b;
    layer1_outputs(1377) <= a;
    layer1_outputs(1378) <= b and not a;
    layer1_outputs(1379) <= a and not b;
    layer1_outputs(1380) <= a or b;
    layer1_outputs(1381) <= not a or b;
    layer1_outputs(1382) <= not b;
    layer1_outputs(1383) <= a and not b;
    layer1_outputs(1384) <= a and b;
    layer1_outputs(1385) <= a;
    layer1_outputs(1386) <= b and not a;
    layer1_outputs(1387) <= not b;
    layer1_outputs(1388) <= a and not b;
    layer1_outputs(1389) <= not a;
    layer1_outputs(1390) <= not (a xor b);
    layer1_outputs(1391) <= a and not b;
    layer1_outputs(1392) <= a xor b;
    layer1_outputs(1393) <= not (a or b);
    layer1_outputs(1394) <= not (a or b);
    layer1_outputs(1395) <= not b;
    layer1_outputs(1396) <= not b;
    layer1_outputs(1397) <= a and b;
    layer1_outputs(1398) <= not a;
    layer1_outputs(1399) <= '0';
    layer1_outputs(1400) <= not b;
    layer1_outputs(1401) <= a or b;
    layer1_outputs(1402) <= a;
    layer1_outputs(1403) <= not (a and b);
    layer1_outputs(1404) <= not a;
    layer1_outputs(1405) <= b;
    layer1_outputs(1406) <= a and b;
    layer1_outputs(1407) <= not (a xor b);
    layer1_outputs(1408) <= a or b;
    layer1_outputs(1409) <= b and not a;
    layer1_outputs(1410) <= '1';
    layer1_outputs(1411) <= a;
    layer1_outputs(1412) <= not a;
    layer1_outputs(1413) <= b and not a;
    layer1_outputs(1414) <= not (a or b);
    layer1_outputs(1415) <= '0';
    layer1_outputs(1416) <= b and not a;
    layer1_outputs(1417) <= not (a and b);
    layer1_outputs(1418) <= not b or a;
    layer1_outputs(1419) <= b and not a;
    layer1_outputs(1420) <= not b or a;
    layer1_outputs(1421) <= not b;
    layer1_outputs(1422) <= b;
    layer1_outputs(1423) <= not (a or b);
    layer1_outputs(1424) <= b and not a;
    layer1_outputs(1425) <= a and not b;
    layer1_outputs(1426) <= a;
    layer1_outputs(1427) <= a and b;
    layer1_outputs(1428) <= not a or b;
    layer1_outputs(1429) <= not (a or b);
    layer1_outputs(1430) <= '1';
    layer1_outputs(1431) <= a and b;
    layer1_outputs(1432) <= a and not b;
    layer1_outputs(1433) <= '0';
    layer1_outputs(1434) <= a xor b;
    layer1_outputs(1435) <= a or b;
    layer1_outputs(1436) <= a and b;
    layer1_outputs(1437) <= not (a and b);
    layer1_outputs(1438) <= not b;
    layer1_outputs(1439) <= not (a or b);
    layer1_outputs(1440) <= not b;
    layer1_outputs(1441) <= b and not a;
    layer1_outputs(1442) <= a;
    layer1_outputs(1443) <= a and not b;
    layer1_outputs(1444) <= not b;
    layer1_outputs(1445) <= '0';
    layer1_outputs(1446) <= a or b;
    layer1_outputs(1447) <= a xor b;
    layer1_outputs(1448) <= not (a or b);
    layer1_outputs(1449) <= '1';
    layer1_outputs(1450) <= not b or a;
    layer1_outputs(1451) <= not (a or b);
    layer1_outputs(1452) <= a;
    layer1_outputs(1453) <= not (a or b);
    layer1_outputs(1454) <= b;
    layer1_outputs(1455) <= '1';
    layer1_outputs(1456) <= a and not b;
    layer1_outputs(1457) <= b;
    layer1_outputs(1458) <= '0';
    layer1_outputs(1459) <= not b or a;
    layer1_outputs(1460) <= a or b;
    layer1_outputs(1461) <= not b or a;
    layer1_outputs(1462) <= b and not a;
    layer1_outputs(1463) <= not b or a;
    layer1_outputs(1464) <= a or b;
    layer1_outputs(1465) <= not (a or b);
    layer1_outputs(1466) <= not b;
    layer1_outputs(1467) <= '0';
    layer1_outputs(1468) <= '1';
    layer1_outputs(1469) <= b and not a;
    layer1_outputs(1470) <= a;
    layer1_outputs(1471) <= a or b;
    layer1_outputs(1472) <= a and not b;
    layer1_outputs(1473) <= not b or a;
    layer1_outputs(1474) <= a or b;
    layer1_outputs(1475) <= '1';
    layer1_outputs(1476) <= a xor b;
    layer1_outputs(1477) <= b;
    layer1_outputs(1478) <= not (a and b);
    layer1_outputs(1479) <= a or b;
    layer1_outputs(1480) <= b;
    layer1_outputs(1481) <= '1';
    layer1_outputs(1482) <= not (a or b);
    layer1_outputs(1483) <= not b;
    layer1_outputs(1484) <= not a or b;
    layer1_outputs(1485) <= not b;
    layer1_outputs(1486) <= '0';
    layer1_outputs(1487) <= a;
    layer1_outputs(1488) <= '1';
    layer1_outputs(1489) <= not (a xor b);
    layer1_outputs(1490) <= not (a xor b);
    layer1_outputs(1491) <= '0';
    layer1_outputs(1492) <= a and not b;
    layer1_outputs(1493) <= not a;
    layer1_outputs(1494) <= not b;
    layer1_outputs(1495) <= a xor b;
    layer1_outputs(1496) <= not b;
    layer1_outputs(1497) <= not b or a;
    layer1_outputs(1498) <= not b;
    layer1_outputs(1499) <= not b;
    layer1_outputs(1500) <= '1';
    layer1_outputs(1501) <= '0';
    layer1_outputs(1502) <= '0';
    layer1_outputs(1503) <= not b or a;
    layer1_outputs(1504) <= b;
    layer1_outputs(1505) <= '1';
    layer1_outputs(1506) <= not b;
    layer1_outputs(1507) <= not (a and b);
    layer1_outputs(1508) <= not a or b;
    layer1_outputs(1509) <= not b or a;
    layer1_outputs(1510) <= a xor b;
    layer1_outputs(1511) <= not (a or b);
    layer1_outputs(1512) <= not (a and b);
    layer1_outputs(1513) <= not (a and b);
    layer1_outputs(1514) <= not b or a;
    layer1_outputs(1515) <= not a or b;
    layer1_outputs(1516) <= b and not a;
    layer1_outputs(1517) <= a and not b;
    layer1_outputs(1518) <= '0';
    layer1_outputs(1519) <= '1';
    layer1_outputs(1520) <= '1';
    layer1_outputs(1521) <= a and b;
    layer1_outputs(1522) <= not (a or b);
    layer1_outputs(1523) <= '0';
    layer1_outputs(1524) <= '0';
    layer1_outputs(1525) <= not a;
    layer1_outputs(1526) <= not (a and b);
    layer1_outputs(1527) <= not (a and b);
    layer1_outputs(1528) <= a or b;
    layer1_outputs(1529) <= not (a or b);
    layer1_outputs(1530) <= not (a and b);
    layer1_outputs(1531) <= not (a and b);
    layer1_outputs(1532) <= not b or a;
    layer1_outputs(1533) <= not (a or b);
    layer1_outputs(1534) <= '1';
    layer1_outputs(1535) <= '1';
    layer1_outputs(1536) <= a and not b;
    layer1_outputs(1537) <= a and b;
    layer1_outputs(1538) <= '0';
    layer1_outputs(1539) <= '0';
    layer1_outputs(1540) <= a and not b;
    layer1_outputs(1541) <= not b or a;
    layer1_outputs(1542) <= '0';
    layer1_outputs(1543) <= a and not b;
    layer1_outputs(1544) <= not a;
    layer1_outputs(1545) <= not (a or b);
    layer1_outputs(1546) <= not (a or b);
    layer1_outputs(1547) <= '0';
    layer1_outputs(1548) <= not a or b;
    layer1_outputs(1549) <= a and not b;
    layer1_outputs(1550) <= b and not a;
    layer1_outputs(1551) <= a and b;
    layer1_outputs(1552) <= a and not b;
    layer1_outputs(1553) <= '0';
    layer1_outputs(1554) <= '1';
    layer1_outputs(1555) <= a and not b;
    layer1_outputs(1556) <= b;
    layer1_outputs(1557) <= not a;
    layer1_outputs(1558) <= a or b;
    layer1_outputs(1559) <= a or b;
    layer1_outputs(1560) <= not (a or b);
    layer1_outputs(1561) <= not b;
    layer1_outputs(1562) <= not a;
    layer1_outputs(1563) <= not a;
    layer1_outputs(1564) <= not a;
    layer1_outputs(1565) <= not (a and b);
    layer1_outputs(1566) <= '0';
    layer1_outputs(1567) <= not a or b;
    layer1_outputs(1568) <= '1';
    layer1_outputs(1569) <= not b;
    layer1_outputs(1570) <= not b or a;
    layer1_outputs(1571) <= '0';
    layer1_outputs(1572) <= a;
    layer1_outputs(1573) <= not a or b;
    layer1_outputs(1574) <= a or b;
    layer1_outputs(1575) <= not a;
    layer1_outputs(1576) <= not b or a;
    layer1_outputs(1577) <= a;
    layer1_outputs(1578) <= a or b;
    layer1_outputs(1579) <= '1';
    layer1_outputs(1580) <= b and not a;
    layer1_outputs(1581) <= not (a and b);
    layer1_outputs(1582) <= '0';
    layer1_outputs(1583) <= a and not b;
    layer1_outputs(1584) <= not (a and b);
    layer1_outputs(1585) <= '1';
    layer1_outputs(1586) <= not (a or b);
    layer1_outputs(1587) <= b;
    layer1_outputs(1588) <= not a or b;
    layer1_outputs(1589) <= a or b;
    layer1_outputs(1590) <= '1';
    layer1_outputs(1591) <= a and b;
    layer1_outputs(1592) <= b;
    layer1_outputs(1593) <= a and not b;
    layer1_outputs(1594) <= a;
    layer1_outputs(1595) <= not a;
    layer1_outputs(1596) <= '1';
    layer1_outputs(1597) <= a or b;
    layer1_outputs(1598) <= b and not a;
    layer1_outputs(1599) <= '1';
    layer1_outputs(1600) <= not (a and b);
    layer1_outputs(1601) <= a and b;
    layer1_outputs(1602) <= b and not a;
    layer1_outputs(1603) <= a or b;
    layer1_outputs(1604) <= not a or b;
    layer1_outputs(1605) <= '0';
    layer1_outputs(1606) <= '1';
    layer1_outputs(1607) <= b and not a;
    layer1_outputs(1608) <= not b or a;
    layer1_outputs(1609) <= b and not a;
    layer1_outputs(1610) <= a and not b;
    layer1_outputs(1611) <= b;
    layer1_outputs(1612) <= a xor b;
    layer1_outputs(1613) <= not b;
    layer1_outputs(1614) <= not a or b;
    layer1_outputs(1615) <= not (a and b);
    layer1_outputs(1616) <= a and not b;
    layer1_outputs(1617) <= '1';
    layer1_outputs(1618) <= a or b;
    layer1_outputs(1619) <= not (a and b);
    layer1_outputs(1620) <= not b;
    layer1_outputs(1621) <= not (a or b);
    layer1_outputs(1622) <= not (a and b);
    layer1_outputs(1623) <= a and not b;
    layer1_outputs(1624) <= a;
    layer1_outputs(1625) <= '1';
    layer1_outputs(1626) <= not (a xor b);
    layer1_outputs(1627) <= '0';
    layer1_outputs(1628) <= a and b;
    layer1_outputs(1629) <= '1';
    layer1_outputs(1630) <= a or b;
    layer1_outputs(1631) <= not a or b;
    layer1_outputs(1632) <= a and not b;
    layer1_outputs(1633) <= not a;
    layer1_outputs(1634) <= not a or b;
    layer1_outputs(1635) <= not b;
    layer1_outputs(1636) <= a or b;
    layer1_outputs(1637) <= not b or a;
    layer1_outputs(1638) <= not b;
    layer1_outputs(1639) <= a and not b;
    layer1_outputs(1640) <= not (a xor b);
    layer1_outputs(1641) <= not (a or b);
    layer1_outputs(1642) <= not b;
    layer1_outputs(1643) <= not (a and b);
    layer1_outputs(1644) <= a and b;
    layer1_outputs(1645) <= b;
    layer1_outputs(1646) <= a or b;
    layer1_outputs(1647) <= '1';
    layer1_outputs(1648) <= b and not a;
    layer1_outputs(1649) <= b and not a;
    layer1_outputs(1650) <= '0';
    layer1_outputs(1651) <= not a;
    layer1_outputs(1652) <= not b;
    layer1_outputs(1653) <= not a or b;
    layer1_outputs(1654) <= '1';
    layer1_outputs(1655) <= not (a or b);
    layer1_outputs(1656) <= a or b;
    layer1_outputs(1657) <= a;
    layer1_outputs(1658) <= a or b;
    layer1_outputs(1659) <= '0';
    layer1_outputs(1660) <= not a or b;
    layer1_outputs(1661) <= not (a or b);
    layer1_outputs(1662) <= '1';
    layer1_outputs(1663) <= '0';
    layer1_outputs(1664) <= not (a or b);
    layer1_outputs(1665) <= a and b;
    layer1_outputs(1666) <= not (a and b);
    layer1_outputs(1667) <= a;
    layer1_outputs(1668) <= b and not a;
    layer1_outputs(1669) <= not a or b;
    layer1_outputs(1670) <= b;
    layer1_outputs(1671) <= a or b;
    layer1_outputs(1672) <= not (a xor b);
    layer1_outputs(1673) <= '0';
    layer1_outputs(1674) <= a;
    layer1_outputs(1675) <= '1';
    layer1_outputs(1676) <= a;
    layer1_outputs(1677) <= not a;
    layer1_outputs(1678) <= '0';
    layer1_outputs(1679) <= '1';
    layer1_outputs(1680) <= not (a xor b);
    layer1_outputs(1681) <= a xor b;
    layer1_outputs(1682) <= not (a or b);
    layer1_outputs(1683) <= not b;
    layer1_outputs(1684) <= not a or b;
    layer1_outputs(1685) <= '1';
    layer1_outputs(1686) <= a or b;
    layer1_outputs(1687) <= not b or a;
    layer1_outputs(1688) <= not (a or b);
    layer1_outputs(1689) <= b and not a;
    layer1_outputs(1690) <= not b;
    layer1_outputs(1691) <= a and b;
    layer1_outputs(1692) <= a and b;
    layer1_outputs(1693) <= b and not a;
    layer1_outputs(1694) <= '1';
    layer1_outputs(1695) <= a;
    layer1_outputs(1696) <= a or b;
    layer1_outputs(1697) <= not a or b;
    layer1_outputs(1698) <= a and b;
    layer1_outputs(1699) <= a or b;
    layer1_outputs(1700) <= a;
    layer1_outputs(1701) <= a and not b;
    layer1_outputs(1702) <= '1';
    layer1_outputs(1703) <= a or b;
    layer1_outputs(1704) <= not a;
    layer1_outputs(1705) <= not a or b;
    layer1_outputs(1706) <= not a;
    layer1_outputs(1707) <= a;
    layer1_outputs(1708) <= not a or b;
    layer1_outputs(1709) <= not b or a;
    layer1_outputs(1710) <= a and not b;
    layer1_outputs(1711) <= a and not b;
    layer1_outputs(1712) <= not (a and b);
    layer1_outputs(1713) <= a and not b;
    layer1_outputs(1714) <= not (a or b);
    layer1_outputs(1715) <= b;
    layer1_outputs(1716) <= not a or b;
    layer1_outputs(1717) <= not a or b;
    layer1_outputs(1718) <= not (a xor b);
    layer1_outputs(1719) <= not (a and b);
    layer1_outputs(1720) <= a or b;
    layer1_outputs(1721) <= '1';
    layer1_outputs(1722) <= '0';
    layer1_outputs(1723) <= b;
    layer1_outputs(1724) <= a or b;
    layer1_outputs(1725) <= a and not b;
    layer1_outputs(1726) <= a and b;
    layer1_outputs(1727) <= b and not a;
    layer1_outputs(1728) <= a and not b;
    layer1_outputs(1729) <= not b;
    layer1_outputs(1730) <= not a or b;
    layer1_outputs(1731) <= not (a xor b);
    layer1_outputs(1732) <= not (a or b);
    layer1_outputs(1733) <= a and not b;
    layer1_outputs(1734) <= '0';
    layer1_outputs(1735) <= a and not b;
    layer1_outputs(1736) <= not a;
    layer1_outputs(1737) <= b and not a;
    layer1_outputs(1738) <= '0';
    layer1_outputs(1739) <= a and not b;
    layer1_outputs(1740) <= '0';
    layer1_outputs(1741) <= not b;
    layer1_outputs(1742) <= '1';
    layer1_outputs(1743) <= not (a xor b);
    layer1_outputs(1744) <= '1';
    layer1_outputs(1745) <= a;
    layer1_outputs(1746) <= '0';
    layer1_outputs(1747) <= not (a or b);
    layer1_outputs(1748) <= not b;
    layer1_outputs(1749) <= b and not a;
    layer1_outputs(1750) <= not b;
    layer1_outputs(1751) <= not (a and b);
    layer1_outputs(1752) <= '0';
    layer1_outputs(1753) <= b and not a;
    layer1_outputs(1754) <= not a;
    layer1_outputs(1755) <= not (a or b);
    layer1_outputs(1756) <= not (a and b);
    layer1_outputs(1757) <= b and not a;
    layer1_outputs(1758) <= not a or b;
    layer1_outputs(1759) <= b;
    layer1_outputs(1760) <= not b;
    layer1_outputs(1761) <= not b or a;
    layer1_outputs(1762) <= not b or a;
    layer1_outputs(1763) <= a;
    layer1_outputs(1764) <= b and not a;
    layer1_outputs(1765) <= b;
    layer1_outputs(1766) <= not a;
    layer1_outputs(1767) <= a and b;
    layer1_outputs(1768) <= b and not a;
    layer1_outputs(1769) <= not a or b;
    layer1_outputs(1770) <= not (a xor b);
    layer1_outputs(1771) <= a and b;
    layer1_outputs(1772) <= b;
    layer1_outputs(1773) <= b;
    layer1_outputs(1774) <= b and not a;
    layer1_outputs(1775) <= not a or b;
    layer1_outputs(1776) <= a and b;
    layer1_outputs(1777) <= a or b;
    layer1_outputs(1778) <= '0';
    layer1_outputs(1779) <= a xor b;
    layer1_outputs(1780) <= a;
    layer1_outputs(1781) <= a and not b;
    layer1_outputs(1782) <= a;
    layer1_outputs(1783) <= a or b;
    layer1_outputs(1784) <= not a or b;
    layer1_outputs(1785) <= b;
    layer1_outputs(1786) <= a;
    layer1_outputs(1787) <= a and b;
    layer1_outputs(1788) <= '1';
    layer1_outputs(1789) <= not a;
    layer1_outputs(1790) <= not a or b;
    layer1_outputs(1791) <= b and not a;
    layer1_outputs(1792) <= '0';
    layer1_outputs(1793) <= a and not b;
    layer1_outputs(1794) <= b and not a;
    layer1_outputs(1795) <= b and not a;
    layer1_outputs(1796) <= not (a xor b);
    layer1_outputs(1797) <= '0';
    layer1_outputs(1798) <= '0';
    layer1_outputs(1799) <= not a;
    layer1_outputs(1800) <= '0';
    layer1_outputs(1801) <= b;
    layer1_outputs(1802) <= a and not b;
    layer1_outputs(1803) <= not a or b;
    layer1_outputs(1804) <= a;
    layer1_outputs(1805) <= b;
    layer1_outputs(1806) <= '1';
    layer1_outputs(1807) <= a or b;
    layer1_outputs(1808) <= a or b;
    layer1_outputs(1809) <= a;
    layer1_outputs(1810) <= not a;
    layer1_outputs(1811) <= not b;
    layer1_outputs(1812) <= a and b;
    layer1_outputs(1813) <= not a;
    layer1_outputs(1814) <= a and not b;
    layer1_outputs(1815) <= not a;
    layer1_outputs(1816) <= a and b;
    layer1_outputs(1817) <= not a;
    layer1_outputs(1818) <= b;
    layer1_outputs(1819) <= '1';
    layer1_outputs(1820) <= not (a xor b);
    layer1_outputs(1821) <= not a or b;
    layer1_outputs(1822) <= not a or b;
    layer1_outputs(1823) <= not b;
    layer1_outputs(1824) <= '0';
    layer1_outputs(1825) <= a;
    layer1_outputs(1826) <= not (a and b);
    layer1_outputs(1827) <= not b;
    layer1_outputs(1828) <= not b or a;
    layer1_outputs(1829) <= not a or b;
    layer1_outputs(1830) <= a xor b;
    layer1_outputs(1831) <= '0';
    layer1_outputs(1832) <= a and b;
    layer1_outputs(1833) <= a and not b;
    layer1_outputs(1834) <= not (a and b);
    layer1_outputs(1835) <= not (a or b);
    layer1_outputs(1836) <= a and not b;
    layer1_outputs(1837) <= a;
    layer1_outputs(1838) <= a;
    layer1_outputs(1839) <= not a or b;
    layer1_outputs(1840) <= '1';
    layer1_outputs(1841) <= b;
    layer1_outputs(1842) <= '1';
    layer1_outputs(1843) <= not (a xor b);
    layer1_outputs(1844) <= '0';
    layer1_outputs(1845) <= not a;
    layer1_outputs(1846) <= a or b;
    layer1_outputs(1847) <= a and not b;
    layer1_outputs(1848) <= a and not b;
    layer1_outputs(1849) <= a;
    layer1_outputs(1850) <= a or b;
    layer1_outputs(1851) <= a;
    layer1_outputs(1852) <= '1';
    layer1_outputs(1853) <= a;
    layer1_outputs(1854) <= not b;
    layer1_outputs(1855) <= not a;
    layer1_outputs(1856) <= a and b;
    layer1_outputs(1857) <= not (a or b);
    layer1_outputs(1858) <= a or b;
    layer1_outputs(1859) <= a and b;
    layer1_outputs(1860) <= b;
    layer1_outputs(1861) <= not a;
    layer1_outputs(1862) <= not b;
    layer1_outputs(1863) <= '1';
    layer1_outputs(1864) <= not (a and b);
    layer1_outputs(1865) <= a or b;
    layer1_outputs(1866) <= not (a xor b);
    layer1_outputs(1867) <= not (a or b);
    layer1_outputs(1868) <= not a;
    layer1_outputs(1869) <= a and b;
    layer1_outputs(1870) <= a or b;
    layer1_outputs(1871) <= '0';
    layer1_outputs(1872) <= not (a or b);
    layer1_outputs(1873) <= not a;
    layer1_outputs(1874) <= not b;
    layer1_outputs(1875) <= '1';
    layer1_outputs(1876) <= '1';
    layer1_outputs(1877) <= b and not a;
    layer1_outputs(1878) <= '0';
    layer1_outputs(1879) <= a;
    layer1_outputs(1880) <= a and b;
    layer1_outputs(1881) <= not (a or b);
    layer1_outputs(1882) <= not a or b;
    layer1_outputs(1883) <= not (a or b);
    layer1_outputs(1884) <= not a;
    layer1_outputs(1885) <= not b or a;
    layer1_outputs(1886) <= a xor b;
    layer1_outputs(1887) <= b;
    layer1_outputs(1888) <= b and not a;
    layer1_outputs(1889) <= a or b;
    layer1_outputs(1890) <= not (a and b);
    layer1_outputs(1891) <= b and not a;
    layer1_outputs(1892) <= '1';
    layer1_outputs(1893) <= b and not a;
    layer1_outputs(1894) <= not (a or b);
    layer1_outputs(1895) <= not b;
    layer1_outputs(1896) <= a and not b;
    layer1_outputs(1897) <= a and b;
    layer1_outputs(1898) <= '1';
    layer1_outputs(1899) <= b;
    layer1_outputs(1900) <= not (a or b);
    layer1_outputs(1901) <= '0';
    layer1_outputs(1902) <= not a or b;
    layer1_outputs(1903) <= not (a or b);
    layer1_outputs(1904) <= not b;
    layer1_outputs(1905) <= not (a or b);
    layer1_outputs(1906) <= not a or b;
    layer1_outputs(1907) <= '0';
    layer1_outputs(1908) <= not a;
    layer1_outputs(1909) <= not (a xor b);
    layer1_outputs(1910) <= a xor b;
    layer1_outputs(1911) <= not a;
    layer1_outputs(1912) <= not b;
    layer1_outputs(1913) <= not a or b;
    layer1_outputs(1914) <= not (a or b);
    layer1_outputs(1915) <= not a or b;
    layer1_outputs(1916) <= a and not b;
    layer1_outputs(1917) <= not b or a;
    layer1_outputs(1918) <= '1';
    layer1_outputs(1919) <= not a or b;
    layer1_outputs(1920) <= a and not b;
    layer1_outputs(1921) <= not (a or b);
    layer1_outputs(1922) <= a;
    layer1_outputs(1923) <= '0';
    layer1_outputs(1924) <= a or b;
    layer1_outputs(1925) <= not b or a;
    layer1_outputs(1926) <= '1';
    layer1_outputs(1927) <= not (a and b);
    layer1_outputs(1928) <= not (a or b);
    layer1_outputs(1929) <= '1';
    layer1_outputs(1930) <= not a;
    layer1_outputs(1931) <= a;
    layer1_outputs(1932) <= '0';
    layer1_outputs(1933) <= not b;
    layer1_outputs(1934) <= b and not a;
    layer1_outputs(1935) <= '1';
    layer1_outputs(1936) <= not (a and b);
    layer1_outputs(1937) <= not (a or b);
    layer1_outputs(1938) <= '1';
    layer1_outputs(1939) <= b;
    layer1_outputs(1940) <= not (a or b);
    layer1_outputs(1941) <= not a or b;
    layer1_outputs(1942) <= '1';
    layer1_outputs(1943) <= not a;
    layer1_outputs(1944) <= not b;
    layer1_outputs(1945) <= not a;
    layer1_outputs(1946) <= not (a and b);
    layer1_outputs(1947) <= '1';
    layer1_outputs(1948) <= not (a and b);
    layer1_outputs(1949) <= b and not a;
    layer1_outputs(1950) <= not a;
    layer1_outputs(1951) <= '1';
    layer1_outputs(1952) <= a and not b;
    layer1_outputs(1953) <= '0';
    layer1_outputs(1954) <= '1';
    layer1_outputs(1955) <= not a or b;
    layer1_outputs(1956) <= a and not b;
    layer1_outputs(1957) <= a;
    layer1_outputs(1958) <= not b or a;
    layer1_outputs(1959) <= b and not a;
    layer1_outputs(1960) <= a;
    layer1_outputs(1961) <= a;
    layer1_outputs(1962) <= not (a and b);
    layer1_outputs(1963) <= b;
    layer1_outputs(1964) <= a;
    layer1_outputs(1965) <= a;
    layer1_outputs(1966) <= a and b;
    layer1_outputs(1967) <= not a;
    layer1_outputs(1968) <= b;
    layer1_outputs(1969) <= not a or b;
    layer1_outputs(1970) <= '0';
    layer1_outputs(1971) <= not b;
    layer1_outputs(1972) <= b and not a;
    layer1_outputs(1973) <= '0';
    layer1_outputs(1974) <= not a or b;
    layer1_outputs(1975) <= not a or b;
    layer1_outputs(1976) <= '0';
    layer1_outputs(1977) <= not a;
    layer1_outputs(1978) <= not (a or b);
    layer1_outputs(1979) <= a;
    layer1_outputs(1980) <= a;
    layer1_outputs(1981) <= '0';
    layer1_outputs(1982) <= not a;
    layer1_outputs(1983) <= '1';
    layer1_outputs(1984) <= a and b;
    layer1_outputs(1985) <= not b or a;
    layer1_outputs(1986) <= a;
    layer1_outputs(1987) <= a;
    layer1_outputs(1988) <= '0';
    layer1_outputs(1989) <= '1';
    layer1_outputs(1990) <= not (a or b);
    layer1_outputs(1991) <= not (a or b);
    layer1_outputs(1992) <= not (a xor b);
    layer1_outputs(1993) <= b and not a;
    layer1_outputs(1994) <= '0';
    layer1_outputs(1995) <= not b or a;
    layer1_outputs(1996) <= a;
    layer1_outputs(1997) <= b;
    layer1_outputs(1998) <= not (a or b);
    layer1_outputs(1999) <= a and b;
    layer1_outputs(2000) <= not (a or b);
    layer1_outputs(2001) <= not (a or b);
    layer1_outputs(2002) <= not b;
    layer1_outputs(2003) <= not b;
    layer1_outputs(2004) <= not (a or b);
    layer1_outputs(2005) <= a or b;
    layer1_outputs(2006) <= not a;
    layer1_outputs(2007) <= a and not b;
    layer1_outputs(2008) <= '0';
    layer1_outputs(2009) <= not b or a;
    layer1_outputs(2010) <= not b or a;
    layer1_outputs(2011) <= b and not a;
    layer1_outputs(2012) <= not b or a;
    layer1_outputs(2013) <= a xor b;
    layer1_outputs(2014) <= '0';
    layer1_outputs(2015) <= a or b;
    layer1_outputs(2016) <= a or b;
    layer1_outputs(2017) <= a xor b;
    layer1_outputs(2018) <= not (a or b);
    layer1_outputs(2019) <= not (a and b);
    layer1_outputs(2020) <= not (a or b);
    layer1_outputs(2021) <= b and not a;
    layer1_outputs(2022) <= '1';
    layer1_outputs(2023) <= b;
    layer1_outputs(2024) <= not a or b;
    layer1_outputs(2025) <= '0';
    layer1_outputs(2026) <= not a or b;
    layer1_outputs(2027) <= not (a or b);
    layer1_outputs(2028) <= a or b;
    layer1_outputs(2029) <= '0';
    layer1_outputs(2030) <= not a;
    layer1_outputs(2031) <= '0';
    layer1_outputs(2032) <= '1';
    layer1_outputs(2033) <= not b or a;
    layer1_outputs(2034) <= a;
    layer1_outputs(2035) <= not b or a;
    layer1_outputs(2036) <= not (a and b);
    layer1_outputs(2037) <= not b or a;
    layer1_outputs(2038) <= not (a and b);
    layer1_outputs(2039) <= a and b;
    layer1_outputs(2040) <= '0';
    layer1_outputs(2041) <= not a or b;
    layer1_outputs(2042) <= '0';
    layer1_outputs(2043) <= '0';
    layer1_outputs(2044) <= not (a xor b);
    layer1_outputs(2045) <= '1';
    layer1_outputs(2046) <= b;
    layer1_outputs(2047) <= '1';
    layer1_outputs(2048) <= not a;
    layer1_outputs(2049) <= a;
    layer1_outputs(2050) <= a and not b;
    layer1_outputs(2051) <= not b or a;
    layer1_outputs(2052) <= not (a and b);
    layer1_outputs(2053) <= a and b;
    layer1_outputs(2054) <= '0';
    layer1_outputs(2055) <= not (a or b);
    layer1_outputs(2056) <= not (a or b);
    layer1_outputs(2057) <= a xor b;
    layer1_outputs(2058) <= not b;
    layer1_outputs(2059) <= not b;
    layer1_outputs(2060) <= '1';
    layer1_outputs(2061) <= '1';
    layer1_outputs(2062) <= not b or a;
    layer1_outputs(2063) <= a or b;
    layer1_outputs(2064) <= a and not b;
    layer1_outputs(2065) <= not (a or b);
    layer1_outputs(2066) <= a and not b;
    layer1_outputs(2067) <= not (a or b);
    layer1_outputs(2068) <= not b or a;
    layer1_outputs(2069) <= not (a or b);
    layer1_outputs(2070) <= '0';
    layer1_outputs(2071) <= a;
    layer1_outputs(2072) <= a or b;
    layer1_outputs(2073) <= not (a and b);
    layer1_outputs(2074) <= not a;
    layer1_outputs(2075) <= not (a or b);
    layer1_outputs(2076) <= a and not b;
    layer1_outputs(2077) <= '1';
    layer1_outputs(2078) <= a or b;
    layer1_outputs(2079) <= a;
    layer1_outputs(2080) <= a or b;
    layer1_outputs(2081) <= b and not a;
    layer1_outputs(2082) <= not (a xor b);
    layer1_outputs(2083) <= not b;
    layer1_outputs(2084) <= not a or b;
    layer1_outputs(2085) <= a or b;
    layer1_outputs(2086) <= b;
    layer1_outputs(2087) <= a or b;
    layer1_outputs(2088) <= not (a and b);
    layer1_outputs(2089) <= not a or b;
    layer1_outputs(2090) <= not b or a;
    layer1_outputs(2091) <= a and b;
    layer1_outputs(2092) <= not a or b;
    layer1_outputs(2093) <= a xor b;
    layer1_outputs(2094) <= not b or a;
    layer1_outputs(2095) <= not b or a;
    layer1_outputs(2096) <= a and not b;
    layer1_outputs(2097) <= not b;
    layer1_outputs(2098) <= '0';
    layer1_outputs(2099) <= b and not a;
    layer1_outputs(2100) <= '0';
    layer1_outputs(2101) <= a and b;
    layer1_outputs(2102) <= not b;
    layer1_outputs(2103) <= '0';
    layer1_outputs(2104) <= b and not a;
    layer1_outputs(2105) <= not b;
    layer1_outputs(2106) <= a and not b;
    layer1_outputs(2107) <= not b;
    layer1_outputs(2108) <= not (a or b);
    layer1_outputs(2109) <= not a or b;
    layer1_outputs(2110) <= not (a and b);
    layer1_outputs(2111) <= a;
    layer1_outputs(2112) <= a or b;
    layer1_outputs(2113) <= a and b;
    layer1_outputs(2114) <= '1';
    layer1_outputs(2115) <= not (a or b);
    layer1_outputs(2116) <= not b;
    layer1_outputs(2117) <= not b or a;
    layer1_outputs(2118) <= a and not b;
    layer1_outputs(2119) <= a and not b;
    layer1_outputs(2120) <= a or b;
    layer1_outputs(2121) <= a and b;
    layer1_outputs(2122) <= '1';
    layer1_outputs(2123) <= not a;
    layer1_outputs(2124) <= not a;
    layer1_outputs(2125) <= a;
    layer1_outputs(2126) <= a and b;
    layer1_outputs(2127) <= '1';
    layer1_outputs(2128) <= not b or a;
    layer1_outputs(2129) <= a and not b;
    layer1_outputs(2130) <= not a;
    layer1_outputs(2131) <= '1';
    layer1_outputs(2132) <= not a;
    layer1_outputs(2133) <= not b or a;
    layer1_outputs(2134) <= b and not a;
    layer1_outputs(2135) <= b;
    layer1_outputs(2136) <= '1';
    layer1_outputs(2137) <= '0';
    layer1_outputs(2138) <= not b or a;
    layer1_outputs(2139) <= '0';
    layer1_outputs(2140) <= not a;
    layer1_outputs(2141) <= not a or b;
    layer1_outputs(2142) <= a and b;
    layer1_outputs(2143) <= '0';
    layer1_outputs(2144) <= not (a or b);
    layer1_outputs(2145) <= not b or a;
    layer1_outputs(2146) <= not a;
    layer1_outputs(2147) <= a and b;
    layer1_outputs(2148) <= b and not a;
    layer1_outputs(2149) <= '1';
    layer1_outputs(2150) <= not (a and b);
    layer1_outputs(2151) <= not b;
    layer1_outputs(2152) <= b;
    layer1_outputs(2153) <= not b;
    layer1_outputs(2154) <= '0';
    layer1_outputs(2155) <= not (a or b);
    layer1_outputs(2156) <= not a;
    layer1_outputs(2157) <= not b;
    layer1_outputs(2158) <= not a;
    layer1_outputs(2159) <= not (a and b);
    layer1_outputs(2160) <= '1';
    layer1_outputs(2161) <= not (a or b);
    layer1_outputs(2162) <= not b or a;
    layer1_outputs(2163) <= not b or a;
    layer1_outputs(2164) <= not b or a;
    layer1_outputs(2165) <= a xor b;
    layer1_outputs(2166) <= not a or b;
    layer1_outputs(2167) <= a or b;
    layer1_outputs(2168) <= not b;
    layer1_outputs(2169) <= '1';
    layer1_outputs(2170) <= not b or a;
    layer1_outputs(2171) <= a and b;
    layer1_outputs(2172) <= not (a or b);
    layer1_outputs(2173) <= not (a or b);
    layer1_outputs(2174) <= b;
    layer1_outputs(2175) <= a and not b;
    layer1_outputs(2176) <= not b or a;
    layer1_outputs(2177) <= not (a or b);
    layer1_outputs(2178) <= a;
    layer1_outputs(2179) <= '0';
    layer1_outputs(2180) <= '0';
    layer1_outputs(2181) <= b;
    layer1_outputs(2182) <= '1';
    layer1_outputs(2183) <= a xor b;
    layer1_outputs(2184) <= '1';
    layer1_outputs(2185) <= '0';
    layer1_outputs(2186) <= a;
    layer1_outputs(2187) <= not b or a;
    layer1_outputs(2188) <= a;
    layer1_outputs(2189) <= not (a xor b);
    layer1_outputs(2190) <= not a;
    layer1_outputs(2191) <= not b or a;
    layer1_outputs(2192) <= '1';
    layer1_outputs(2193) <= not (a and b);
    layer1_outputs(2194) <= b;
    layer1_outputs(2195) <= '0';
    layer1_outputs(2196) <= b;
    layer1_outputs(2197) <= not b;
    layer1_outputs(2198) <= not b;
    layer1_outputs(2199) <= a and b;
    layer1_outputs(2200) <= not a or b;
    layer1_outputs(2201) <= b;
    layer1_outputs(2202) <= not a or b;
    layer1_outputs(2203) <= a and not b;
    layer1_outputs(2204) <= a;
    layer1_outputs(2205) <= '0';
    layer1_outputs(2206) <= not b;
    layer1_outputs(2207) <= a and b;
    layer1_outputs(2208) <= '0';
    layer1_outputs(2209) <= '0';
    layer1_outputs(2210) <= not (a or b);
    layer1_outputs(2211) <= a;
    layer1_outputs(2212) <= a or b;
    layer1_outputs(2213) <= b;
    layer1_outputs(2214) <= a and not b;
    layer1_outputs(2215) <= not b or a;
    layer1_outputs(2216) <= not b or a;
    layer1_outputs(2217) <= a or b;
    layer1_outputs(2218) <= not a or b;
    layer1_outputs(2219) <= '0';
    layer1_outputs(2220) <= not (a or b);
    layer1_outputs(2221) <= '0';
    layer1_outputs(2222) <= a or b;
    layer1_outputs(2223) <= not b or a;
    layer1_outputs(2224) <= not (a xor b);
    layer1_outputs(2225) <= '1';
    layer1_outputs(2226) <= b and not a;
    layer1_outputs(2227) <= not a;
    layer1_outputs(2228) <= not (a and b);
    layer1_outputs(2229) <= not b;
    layer1_outputs(2230) <= not (a and b);
    layer1_outputs(2231) <= '0';
    layer1_outputs(2232) <= '0';
    layer1_outputs(2233) <= not (a or b);
    layer1_outputs(2234) <= not (a or b);
    layer1_outputs(2235) <= '1';
    layer1_outputs(2236) <= a;
    layer1_outputs(2237) <= b and not a;
    layer1_outputs(2238) <= not a;
    layer1_outputs(2239) <= not (a and b);
    layer1_outputs(2240) <= not b or a;
    layer1_outputs(2241) <= a xor b;
    layer1_outputs(2242) <= '0';
    layer1_outputs(2243) <= b;
    layer1_outputs(2244) <= '1';
    layer1_outputs(2245) <= not b or a;
    layer1_outputs(2246) <= '1';
    layer1_outputs(2247) <= not b;
    layer1_outputs(2248) <= not a or b;
    layer1_outputs(2249) <= not (a xor b);
    layer1_outputs(2250) <= a and b;
    layer1_outputs(2251) <= '0';
    layer1_outputs(2252) <= not (a and b);
    layer1_outputs(2253) <= '1';
    layer1_outputs(2254) <= not b;
    layer1_outputs(2255) <= b;
    layer1_outputs(2256) <= not b;
    layer1_outputs(2257) <= a and b;
    layer1_outputs(2258) <= '1';
    layer1_outputs(2259) <= not (a or b);
    layer1_outputs(2260) <= not (a or b);
    layer1_outputs(2261) <= a and not b;
    layer1_outputs(2262) <= a;
    layer1_outputs(2263) <= not b or a;
    layer1_outputs(2264) <= b and not a;
    layer1_outputs(2265) <= not a;
    layer1_outputs(2266) <= not (a or b);
    layer1_outputs(2267) <= a or b;
    layer1_outputs(2268) <= a;
    layer1_outputs(2269) <= not a or b;
    layer1_outputs(2270) <= a;
    layer1_outputs(2271) <= b and not a;
    layer1_outputs(2272) <= b and not a;
    layer1_outputs(2273) <= '1';
    layer1_outputs(2274) <= '0';
    layer1_outputs(2275) <= not a;
    layer1_outputs(2276) <= not a;
    layer1_outputs(2277) <= '0';
    layer1_outputs(2278) <= a xor b;
    layer1_outputs(2279) <= a and b;
    layer1_outputs(2280) <= a and b;
    layer1_outputs(2281) <= a or b;
    layer1_outputs(2282) <= not b or a;
    layer1_outputs(2283) <= a xor b;
    layer1_outputs(2284) <= a or b;
    layer1_outputs(2285) <= not a or b;
    layer1_outputs(2286) <= not a;
    layer1_outputs(2287) <= not (a and b);
    layer1_outputs(2288) <= a and b;
    layer1_outputs(2289) <= not a or b;
    layer1_outputs(2290) <= a;
    layer1_outputs(2291) <= '1';
    layer1_outputs(2292) <= b;
    layer1_outputs(2293) <= a and not b;
    layer1_outputs(2294) <= not b or a;
    layer1_outputs(2295) <= b;
    layer1_outputs(2296) <= not b or a;
    layer1_outputs(2297) <= not b or a;
    layer1_outputs(2298) <= b and not a;
    layer1_outputs(2299) <= a and b;
    layer1_outputs(2300) <= '0';
    layer1_outputs(2301) <= not b or a;
    layer1_outputs(2302) <= b and not a;
    layer1_outputs(2303) <= not b or a;
    layer1_outputs(2304) <= a and b;
    layer1_outputs(2305) <= b and not a;
    layer1_outputs(2306) <= b;
    layer1_outputs(2307) <= '1';
    layer1_outputs(2308) <= a and not b;
    layer1_outputs(2309) <= '0';
    layer1_outputs(2310) <= '0';
    layer1_outputs(2311) <= b and not a;
    layer1_outputs(2312) <= not a or b;
    layer1_outputs(2313) <= not (a xor b);
    layer1_outputs(2314) <= not (a and b);
    layer1_outputs(2315) <= not b;
    layer1_outputs(2316) <= '0';
    layer1_outputs(2317) <= b and not a;
    layer1_outputs(2318) <= a or b;
    layer1_outputs(2319) <= a and not b;
    layer1_outputs(2320) <= a and b;
    layer1_outputs(2321) <= not a or b;
    layer1_outputs(2322) <= not a or b;
    layer1_outputs(2323) <= not (a xor b);
    layer1_outputs(2324) <= '0';
    layer1_outputs(2325) <= '1';
    layer1_outputs(2326) <= '0';
    layer1_outputs(2327) <= not a or b;
    layer1_outputs(2328) <= a and b;
    layer1_outputs(2329) <= b;
    layer1_outputs(2330) <= not (a and b);
    layer1_outputs(2331) <= '1';
    layer1_outputs(2332) <= not b or a;
    layer1_outputs(2333) <= b and not a;
    layer1_outputs(2334) <= '1';
    layer1_outputs(2335) <= not a or b;
    layer1_outputs(2336) <= not b or a;
    layer1_outputs(2337) <= not (a or b);
    layer1_outputs(2338) <= a and b;
    layer1_outputs(2339) <= not a or b;
    layer1_outputs(2340) <= not b or a;
    layer1_outputs(2341) <= a or b;
    layer1_outputs(2342) <= '0';
    layer1_outputs(2343) <= a;
    layer1_outputs(2344) <= '0';
    layer1_outputs(2345) <= not (a and b);
    layer1_outputs(2346) <= '1';
    layer1_outputs(2347) <= a;
    layer1_outputs(2348) <= not b;
    layer1_outputs(2349) <= '1';
    layer1_outputs(2350) <= not b;
    layer1_outputs(2351) <= b and not a;
    layer1_outputs(2352) <= a and b;
    layer1_outputs(2353) <= b;
    layer1_outputs(2354) <= not (a or b);
    layer1_outputs(2355) <= '1';
    layer1_outputs(2356) <= not b or a;
    layer1_outputs(2357) <= a;
    layer1_outputs(2358) <= a;
    layer1_outputs(2359) <= a and not b;
    layer1_outputs(2360) <= a and b;
    layer1_outputs(2361) <= not (a xor b);
    layer1_outputs(2362) <= a and b;
    layer1_outputs(2363) <= a or b;
    layer1_outputs(2364) <= not (a and b);
    layer1_outputs(2365) <= b;
    layer1_outputs(2366) <= not a;
    layer1_outputs(2367) <= '0';
    layer1_outputs(2368) <= b;
    layer1_outputs(2369) <= not (a or b);
    layer1_outputs(2370) <= a and not b;
    layer1_outputs(2371) <= not (a or b);
    layer1_outputs(2372) <= a and b;
    layer1_outputs(2373) <= '0';
    layer1_outputs(2374) <= not a or b;
    layer1_outputs(2375) <= a or b;
    layer1_outputs(2376) <= not (a or b);
    layer1_outputs(2377) <= not a or b;
    layer1_outputs(2378) <= b;
    layer1_outputs(2379) <= '1';
    layer1_outputs(2380) <= not (a or b);
    layer1_outputs(2381) <= a and not b;
    layer1_outputs(2382) <= not (a and b);
    layer1_outputs(2383) <= '1';
    layer1_outputs(2384) <= b and not a;
    layer1_outputs(2385) <= not a;
    layer1_outputs(2386) <= not b or a;
    layer1_outputs(2387) <= '0';
    layer1_outputs(2388) <= b and not a;
    layer1_outputs(2389) <= not (a and b);
    layer1_outputs(2390) <= '0';
    layer1_outputs(2391) <= b;
    layer1_outputs(2392) <= not b or a;
    layer1_outputs(2393) <= not b or a;
    layer1_outputs(2394) <= a;
    layer1_outputs(2395) <= not (a or b);
    layer1_outputs(2396) <= not b;
    layer1_outputs(2397) <= '1';
    layer1_outputs(2398) <= '1';
    layer1_outputs(2399) <= a and b;
    layer1_outputs(2400) <= not b or a;
    layer1_outputs(2401) <= not a;
    layer1_outputs(2402) <= not b or a;
    layer1_outputs(2403) <= not a;
    layer1_outputs(2404) <= not a or b;
    layer1_outputs(2405) <= a and not b;
    layer1_outputs(2406) <= a and not b;
    layer1_outputs(2407) <= not (a and b);
    layer1_outputs(2408) <= '0';
    layer1_outputs(2409) <= not a or b;
    layer1_outputs(2410) <= b;
    layer1_outputs(2411) <= b;
    layer1_outputs(2412) <= a or b;
    layer1_outputs(2413) <= '0';
    layer1_outputs(2414) <= not a;
    layer1_outputs(2415) <= a and not b;
    layer1_outputs(2416) <= a and b;
    layer1_outputs(2417) <= a or b;
    layer1_outputs(2418) <= a or b;
    layer1_outputs(2419) <= '1';
    layer1_outputs(2420) <= not a or b;
    layer1_outputs(2421) <= not b or a;
    layer1_outputs(2422) <= '1';
    layer1_outputs(2423) <= '0';
    layer1_outputs(2424) <= not (a xor b);
    layer1_outputs(2425) <= b and not a;
    layer1_outputs(2426) <= '1';
    layer1_outputs(2427) <= not (a and b);
    layer1_outputs(2428) <= b;
    layer1_outputs(2429) <= a;
    layer1_outputs(2430) <= a and b;
    layer1_outputs(2431) <= not (a and b);
    layer1_outputs(2432) <= '1';
    layer1_outputs(2433) <= '1';
    layer1_outputs(2434) <= '0';
    layer1_outputs(2435) <= not b or a;
    layer1_outputs(2436) <= a or b;
    layer1_outputs(2437) <= not b or a;
    layer1_outputs(2438) <= b;
    layer1_outputs(2439) <= not b;
    layer1_outputs(2440) <= not (a xor b);
    layer1_outputs(2441) <= not (a or b);
    layer1_outputs(2442) <= not a or b;
    layer1_outputs(2443) <= '0';
    layer1_outputs(2444) <= not b;
    layer1_outputs(2445) <= b;
    layer1_outputs(2446) <= not b;
    layer1_outputs(2447) <= a;
    layer1_outputs(2448) <= b and not a;
    layer1_outputs(2449) <= a and b;
    layer1_outputs(2450) <= a and not b;
    layer1_outputs(2451) <= not (a or b);
    layer1_outputs(2452) <= b and not a;
    layer1_outputs(2453) <= '1';
    layer1_outputs(2454) <= '1';
    layer1_outputs(2455) <= a and not b;
    layer1_outputs(2456) <= b;
    layer1_outputs(2457) <= b and not a;
    layer1_outputs(2458) <= not b;
    layer1_outputs(2459) <= not (a and b);
    layer1_outputs(2460) <= '0';
    layer1_outputs(2461) <= not (a or b);
    layer1_outputs(2462) <= '0';
    layer1_outputs(2463) <= a or b;
    layer1_outputs(2464) <= a or b;
    layer1_outputs(2465) <= a and not b;
    layer1_outputs(2466) <= '1';
    layer1_outputs(2467) <= not b;
    layer1_outputs(2468) <= b and not a;
    layer1_outputs(2469) <= a and b;
    layer1_outputs(2470) <= a and b;
    layer1_outputs(2471) <= a and not b;
    layer1_outputs(2472) <= b and not a;
    layer1_outputs(2473) <= not a;
    layer1_outputs(2474) <= b;
    layer1_outputs(2475) <= not b or a;
    layer1_outputs(2476) <= b and not a;
    layer1_outputs(2477) <= not b or a;
    layer1_outputs(2478) <= not a or b;
    layer1_outputs(2479) <= not (a and b);
    layer1_outputs(2480) <= '0';
    layer1_outputs(2481) <= b and not a;
    layer1_outputs(2482) <= a or b;
    layer1_outputs(2483) <= not (a or b);
    layer1_outputs(2484) <= a xor b;
    layer1_outputs(2485) <= '0';
    layer1_outputs(2486) <= not a;
    layer1_outputs(2487) <= a and b;
    layer1_outputs(2488) <= not (a xor b);
    layer1_outputs(2489) <= not (a and b);
    layer1_outputs(2490) <= b;
    layer1_outputs(2491) <= not (a or b);
    layer1_outputs(2492) <= not a or b;
    layer1_outputs(2493) <= not (a and b);
    layer1_outputs(2494) <= a xor b;
    layer1_outputs(2495) <= '1';
    layer1_outputs(2496) <= a or b;
    layer1_outputs(2497) <= b and not a;
    layer1_outputs(2498) <= b and not a;
    layer1_outputs(2499) <= a and not b;
    layer1_outputs(2500) <= b;
    layer1_outputs(2501) <= a;
    layer1_outputs(2502) <= '1';
    layer1_outputs(2503) <= not (a and b);
    layer1_outputs(2504) <= a or b;
    layer1_outputs(2505) <= '0';
    layer1_outputs(2506) <= not (a or b);
    layer1_outputs(2507) <= not (a or b);
    layer1_outputs(2508) <= not b;
    layer1_outputs(2509) <= not (a or b);
    layer1_outputs(2510) <= a;
    layer1_outputs(2511) <= '1';
    layer1_outputs(2512) <= '1';
    layer1_outputs(2513) <= a;
    layer1_outputs(2514) <= b;
    layer1_outputs(2515) <= not (a and b);
    layer1_outputs(2516) <= '1';
    layer1_outputs(2517) <= not (a and b);
    layer1_outputs(2518) <= not (a and b);
    layer1_outputs(2519) <= a and b;
    layer1_outputs(2520) <= '1';
    layer1_outputs(2521) <= b and not a;
    layer1_outputs(2522) <= b and not a;
    layer1_outputs(2523) <= not b or a;
    layer1_outputs(2524) <= a xor b;
    layer1_outputs(2525) <= not (a or b);
    layer1_outputs(2526) <= '1';
    layer1_outputs(2527) <= a;
    layer1_outputs(2528) <= '0';
    layer1_outputs(2529) <= b and not a;
    layer1_outputs(2530) <= a and b;
    layer1_outputs(2531) <= not b;
    layer1_outputs(2532) <= not a;
    layer1_outputs(2533) <= b and not a;
    layer1_outputs(2534) <= not (a and b);
    layer1_outputs(2535) <= not b;
    layer1_outputs(2536) <= a or b;
    layer1_outputs(2537) <= not b or a;
    layer1_outputs(2538) <= a;
    layer1_outputs(2539) <= not a or b;
    layer1_outputs(2540) <= not a or b;
    layer1_outputs(2541) <= not b or a;
    layer1_outputs(2542) <= b;
    layer1_outputs(2543) <= '0';
    layer1_outputs(2544) <= b and not a;
    layer1_outputs(2545) <= a;
    layer1_outputs(2546) <= b;
    layer1_outputs(2547) <= not b or a;
    layer1_outputs(2548) <= a or b;
    layer1_outputs(2549) <= not (a and b);
    layer1_outputs(2550) <= not a;
    layer1_outputs(2551) <= '1';
    layer1_outputs(2552) <= '0';
    layer1_outputs(2553) <= a or b;
    layer1_outputs(2554) <= a;
    layer1_outputs(2555) <= not b or a;
    layer1_outputs(2556) <= b and not a;
    layer1_outputs(2557) <= '1';
    layer1_outputs(2558) <= b and not a;
    layer1_outputs(2559) <= b;
    layer1_outputs(2560) <= '1';
    layer1_outputs(2561) <= not a;
    layer1_outputs(2562) <= b and not a;
    layer1_outputs(2563) <= not (a or b);
    layer1_outputs(2564) <= not a;
    layer1_outputs(2565) <= a or b;
    layer1_outputs(2566) <= a or b;
    layer1_outputs(2567) <= a;
    layer1_outputs(2568) <= b and not a;
    layer1_outputs(2569) <= not (a or b);
    layer1_outputs(2570) <= '1';
    layer1_outputs(2571) <= a or b;
    layer1_outputs(2572) <= '1';
    layer1_outputs(2573) <= a and b;
    layer1_outputs(2574) <= '0';
    layer1_outputs(2575) <= a;
    layer1_outputs(2576) <= a;
    layer1_outputs(2577) <= '1';
    layer1_outputs(2578) <= not b;
    layer1_outputs(2579) <= not b;
    layer1_outputs(2580) <= a and b;
    layer1_outputs(2581) <= not b;
    layer1_outputs(2582) <= '1';
    layer1_outputs(2583) <= '1';
    layer1_outputs(2584) <= '1';
    layer1_outputs(2585) <= a or b;
    layer1_outputs(2586) <= not a or b;
    layer1_outputs(2587) <= not a;
    layer1_outputs(2588) <= not a;
    layer1_outputs(2589) <= a;
    layer1_outputs(2590) <= not b;
    layer1_outputs(2591) <= '1';
    layer1_outputs(2592) <= not (a and b);
    layer1_outputs(2593) <= '1';
    layer1_outputs(2594) <= not b;
    layer1_outputs(2595) <= '0';
    layer1_outputs(2596) <= '1';
    layer1_outputs(2597) <= not b;
    layer1_outputs(2598) <= '0';
    layer1_outputs(2599) <= a and not b;
    layer1_outputs(2600) <= not a or b;
    layer1_outputs(2601) <= '1';
    layer1_outputs(2602) <= not a;
    layer1_outputs(2603) <= not b;
    layer1_outputs(2604) <= a and not b;
    layer1_outputs(2605) <= a and not b;
    layer1_outputs(2606) <= '1';
    layer1_outputs(2607) <= '0';
    layer1_outputs(2608) <= not (a and b);
    layer1_outputs(2609) <= not a or b;
    layer1_outputs(2610) <= a and b;
    layer1_outputs(2611) <= b and not a;
    layer1_outputs(2612) <= a or b;
    layer1_outputs(2613) <= b and not a;
    layer1_outputs(2614) <= not b or a;
    layer1_outputs(2615) <= '0';
    layer1_outputs(2616) <= a and not b;
    layer1_outputs(2617) <= a;
    layer1_outputs(2618) <= not (a and b);
    layer1_outputs(2619) <= a xor b;
    layer1_outputs(2620) <= a and b;
    layer1_outputs(2621) <= '1';
    layer1_outputs(2622) <= a and not b;
    layer1_outputs(2623) <= not (a or b);
    layer1_outputs(2624) <= not a or b;
    layer1_outputs(2625) <= a and b;
    layer1_outputs(2626) <= a and not b;
    layer1_outputs(2627) <= not b;
    layer1_outputs(2628) <= not a or b;
    layer1_outputs(2629) <= '1';
    layer1_outputs(2630) <= b;
    layer1_outputs(2631) <= not a or b;
    layer1_outputs(2632) <= a xor b;
    layer1_outputs(2633) <= '1';
    layer1_outputs(2634) <= not b or a;
    layer1_outputs(2635) <= '1';
    layer1_outputs(2636) <= not (a xor b);
    layer1_outputs(2637) <= a and b;
    layer1_outputs(2638) <= '0';
    layer1_outputs(2639) <= not b or a;
    layer1_outputs(2640) <= a or b;
    layer1_outputs(2641) <= '0';
    layer1_outputs(2642) <= a;
    layer1_outputs(2643) <= not a or b;
    layer1_outputs(2644) <= not a;
    layer1_outputs(2645) <= '0';
    layer1_outputs(2646) <= not b;
    layer1_outputs(2647) <= a and not b;
    layer1_outputs(2648) <= a and not b;
    layer1_outputs(2649) <= not (a and b);
    layer1_outputs(2650) <= not b;
    layer1_outputs(2651) <= not a or b;
    layer1_outputs(2652) <= not (a and b);
    layer1_outputs(2653) <= not a;
    layer1_outputs(2654) <= '0';
    layer1_outputs(2655) <= '0';
    layer1_outputs(2656) <= '0';
    layer1_outputs(2657) <= not b or a;
    layer1_outputs(2658) <= '0';
    layer1_outputs(2659) <= '1';
    layer1_outputs(2660) <= not b;
    layer1_outputs(2661) <= '0';
    layer1_outputs(2662) <= b;
    layer1_outputs(2663) <= not (a and b);
    layer1_outputs(2664) <= a xor b;
    layer1_outputs(2665) <= not a or b;
    layer1_outputs(2666) <= not b;
    layer1_outputs(2667) <= a or b;
    layer1_outputs(2668) <= not b or a;
    layer1_outputs(2669) <= not a or b;
    layer1_outputs(2670) <= not (a and b);
    layer1_outputs(2671) <= a xor b;
    layer1_outputs(2672) <= a or b;
    layer1_outputs(2673) <= '1';
    layer1_outputs(2674) <= not a or b;
    layer1_outputs(2675) <= b and not a;
    layer1_outputs(2676) <= a and not b;
    layer1_outputs(2677) <= not a;
    layer1_outputs(2678) <= '1';
    layer1_outputs(2679) <= not a or b;
    layer1_outputs(2680) <= not (a or b);
    layer1_outputs(2681) <= not a or b;
    layer1_outputs(2682) <= not b or a;
    layer1_outputs(2683) <= '0';
    layer1_outputs(2684) <= not a;
    layer1_outputs(2685) <= '0';
    layer1_outputs(2686) <= not (a or b);
    layer1_outputs(2687) <= a or b;
    layer1_outputs(2688) <= not b or a;
    layer1_outputs(2689) <= b and not a;
    layer1_outputs(2690) <= a and not b;
    layer1_outputs(2691) <= not a or b;
    layer1_outputs(2692) <= b;
    layer1_outputs(2693) <= not (a and b);
    layer1_outputs(2694) <= '0';
    layer1_outputs(2695) <= b;
    layer1_outputs(2696) <= a and b;
    layer1_outputs(2697) <= a and b;
    layer1_outputs(2698) <= not a;
    layer1_outputs(2699) <= not (a xor b);
    layer1_outputs(2700) <= not (a or b);
    layer1_outputs(2701) <= not b or a;
    layer1_outputs(2702) <= not (a and b);
    layer1_outputs(2703) <= b and not a;
    layer1_outputs(2704) <= b and not a;
    layer1_outputs(2705) <= a and not b;
    layer1_outputs(2706) <= a and not b;
    layer1_outputs(2707) <= b;
    layer1_outputs(2708) <= not a or b;
    layer1_outputs(2709) <= not b or a;
    layer1_outputs(2710) <= not b;
    layer1_outputs(2711) <= a or b;
    layer1_outputs(2712) <= a and not b;
    layer1_outputs(2713) <= not a or b;
    layer1_outputs(2714) <= not a or b;
    layer1_outputs(2715) <= '1';
    layer1_outputs(2716) <= not (a xor b);
    layer1_outputs(2717) <= '0';
    layer1_outputs(2718) <= not b or a;
    layer1_outputs(2719) <= b and not a;
    layer1_outputs(2720) <= a and not b;
    layer1_outputs(2721) <= not (a xor b);
    layer1_outputs(2722) <= not b or a;
    layer1_outputs(2723) <= a and b;
    layer1_outputs(2724) <= b;
    layer1_outputs(2725) <= not a;
    layer1_outputs(2726) <= a xor b;
    layer1_outputs(2727) <= not (a or b);
    layer1_outputs(2728) <= a and not b;
    layer1_outputs(2729) <= a or b;
    layer1_outputs(2730) <= a and not b;
    layer1_outputs(2731) <= not (a and b);
    layer1_outputs(2732) <= a and b;
    layer1_outputs(2733) <= a and not b;
    layer1_outputs(2734) <= a;
    layer1_outputs(2735) <= '0';
    layer1_outputs(2736) <= not a;
    layer1_outputs(2737) <= a and b;
    layer1_outputs(2738) <= a and not b;
    layer1_outputs(2739) <= a;
    layer1_outputs(2740) <= not (a or b);
    layer1_outputs(2741) <= not a;
    layer1_outputs(2742) <= not (a or b);
    layer1_outputs(2743) <= a or b;
    layer1_outputs(2744) <= b and not a;
    layer1_outputs(2745) <= not a;
    layer1_outputs(2746) <= b and not a;
    layer1_outputs(2747) <= not b;
    layer1_outputs(2748) <= '1';
    layer1_outputs(2749) <= not b;
    layer1_outputs(2750) <= '1';
    layer1_outputs(2751) <= '1';
    layer1_outputs(2752) <= not b or a;
    layer1_outputs(2753) <= '1';
    layer1_outputs(2754) <= not (a or b);
    layer1_outputs(2755) <= not (a xor b);
    layer1_outputs(2756) <= '1';
    layer1_outputs(2757) <= a or b;
    layer1_outputs(2758) <= a and not b;
    layer1_outputs(2759) <= not (a and b);
    layer1_outputs(2760) <= not b;
    layer1_outputs(2761) <= not b or a;
    layer1_outputs(2762) <= '1';
    layer1_outputs(2763) <= not (a and b);
    layer1_outputs(2764) <= '1';
    layer1_outputs(2765) <= not b;
    layer1_outputs(2766) <= '0';
    layer1_outputs(2767) <= not b;
    layer1_outputs(2768) <= not b or a;
    layer1_outputs(2769) <= a or b;
    layer1_outputs(2770) <= not (a or b);
    layer1_outputs(2771) <= not (a or b);
    layer1_outputs(2772) <= '0';
    layer1_outputs(2773) <= b and not a;
    layer1_outputs(2774) <= b;
    layer1_outputs(2775) <= '0';
    layer1_outputs(2776) <= not a;
    layer1_outputs(2777) <= '0';
    layer1_outputs(2778) <= not b or a;
    layer1_outputs(2779) <= a and not b;
    layer1_outputs(2780) <= '1';
    layer1_outputs(2781) <= not b or a;
    layer1_outputs(2782) <= a or b;
    layer1_outputs(2783) <= not a;
    layer1_outputs(2784) <= '0';
    layer1_outputs(2785) <= b and not a;
    layer1_outputs(2786) <= '1';
    layer1_outputs(2787) <= a;
    layer1_outputs(2788) <= b and not a;
    layer1_outputs(2789) <= a or b;
    layer1_outputs(2790) <= not b;
    layer1_outputs(2791) <= '0';
    layer1_outputs(2792) <= a and b;
    layer1_outputs(2793) <= a xor b;
    layer1_outputs(2794) <= not (a or b);
    layer1_outputs(2795) <= a;
    layer1_outputs(2796) <= not (a or b);
    layer1_outputs(2797) <= b and not a;
    layer1_outputs(2798) <= not a;
    layer1_outputs(2799) <= a;
    layer1_outputs(2800) <= a xor b;
    layer1_outputs(2801) <= not a or b;
    layer1_outputs(2802) <= b and not a;
    layer1_outputs(2803) <= b and not a;
    layer1_outputs(2804) <= '0';
    layer1_outputs(2805) <= not (a and b);
    layer1_outputs(2806) <= '1';
    layer1_outputs(2807) <= a or b;
    layer1_outputs(2808) <= not b;
    layer1_outputs(2809) <= not b;
    layer1_outputs(2810) <= a and b;
    layer1_outputs(2811) <= b and not a;
    layer1_outputs(2812) <= not b or a;
    layer1_outputs(2813) <= '1';
    layer1_outputs(2814) <= a and b;
    layer1_outputs(2815) <= not a or b;
    layer1_outputs(2816) <= a;
    layer1_outputs(2817) <= a;
    layer1_outputs(2818) <= not b;
    layer1_outputs(2819) <= '1';
    layer1_outputs(2820) <= '0';
    layer1_outputs(2821) <= not a or b;
    layer1_outputs(2822) <= '0';
    layer1_outputs(2823) <= not b or a;
    layer1_outputs(2824) <= '1';
    layer1_outputs(2825) <= a and b;
    layer1_outputs(2826) <= '0';
    layer1_outputs(2827) <= '0';
    layer1_outputs(2828) <= not a;
    layer1_outputs(2829) <= b;
    layer1_outputs(2830) <= not a;
    layer1_outputs(2831) <= a or b;
    layer1_outputs(2832) <= '0';
    layer1_outputs(2833) <= a and b;
    layer1_outputs(2834) <= not (a xor b);
    layer1_outputs(2835) <= not a;
    layer1_outputs(2836) <= not a;
    layer1_outputs(2837) <= a xor b;
    layer1_outputs(2838) <= '0';
    layer1_outputs(2839) <= not (a and b);
    layer1_outputs(2840) <= a;
    layer1_outputs(2841) <= not b or a;
    layer1_outputs(2842) <= '1';
    layer1_outputs(2843) <= b;
    layer1_outputs(2844) <= not (a or b);
    layer1_outputs(2845) <= not (a or b);
    layer1_outputs(2846) <= a and not b;
    layer1_outputs(2847) <= not (a xor b);
    layer1_outputs(2848) <= not (a xor b);
    layer1_outputs(2849) <= a xor b;
    layer1_outputs(2850) <= a xor b;
    layer1_outputs(2851) <= not b;
    layer1_outputs(2852) <= not b;
    layer1_outputs(2853) <= b;
    layer1_outputs(2854) <= not (a and b);
    layer1_outputs(2855) <= '0';
    layer1_outputs(2856) <= b and not a;
    layer1_outputs(2857) <= not (a or b);
    layer1_outputs(2858) <= a xor b;
    layer1_outputs(2859) <= not a;
    layer1_outputs(2860) <= b;
    layer1_outputs(2861) <= '1';
    layer1_outputs(2862) <= not a or b;
    layer1_outputs(2863) <= a and b;
    layer1_outputs(2864) <= a and b;
    layer1_outputs(2865) <= not (a or b);
    layer1_outputs(2866) <= b;
    layer1_outputs(2867) <= a or b;
    layer1_outputs(2868) <= '0';
    layer1_outputs(2869) <= b and not a;
    layer1_outputs(2870) <= '1';
    layer1_outputs(2871) <= a xor b;
    layer1_outputs(2872) <= a;
    layer1_outputs(2873) <= '1';
    layer1_outputs(2874) <= not (a or b);
    layer1_outputs(2875) <= b;
    layer1_outputs(2876) <= not (a xor b);
    layer1_outputs(2877) <= not b;
    layer1_outputs(2878) <= not b or a;
    layer1_outputs(2879) <= not a or b;
    layer1_outputs(2880) <= not a or b;
    layer1_outputs(2881) <= b;
    layer1_outputs(2882) <= a and not b;
    layer1_outputs(2883) <= '1';
    layer1_outputs(2884) <= a or b;
    layer1_outputs(2885) <= a xor b;
    layer1_outputs(2886) <= not (a and b);
    layer1_outputs(2887) <= a and b;
    layer1_outputs(2888) <= not (a xor b);
    layer1_outputs(2889) <= '1';
    layer1_outputs(2890) <= not b or a;
    layer1_outputs(2891) <= '1';
    layer1_outputs(2892) <= b;
    layer1_outputs(2893) <= a and not b;
    layer1_outputs(2894) <= b;
    layer1_outputs(2895) <= not (a xor b);
    layer1_outputs(2896) <= b and not a;
    layer1_outputs(2897) <= not b or a;
    layer1_outputs(2898) <= '1';
    layer1_outputs(2899) <= a or b;
    layer1_outputs(2900) <= not (a and b);
    layer1_outputs(2901) <= not a or b;
    layer1_outputs(2902) <= '0';
    layer1_outputs(2903) <= b and not a;
    layer1_outputs(2904) <= not (a xor b);
    layer1_outputs(2905) <= a and not b;
    layer1_outputs(2906) <= b and not a;
    layer1_outputs(2907) <= not a or b;
    layer1_outputs(2908) <= '1';
    layer1_outputs(2909) <= not (a or b);
    layer1_outputs(2910) <= not b or a;
    layer1_outputs(2911) <= not a or b;
    layer1_outputs(2912) <= a;
    layer1_outputs(2913) <= '1';
    layer1_outputs(2914) <= a and not b;
    layer1_outputs(2915) <= a or b;
    layer1_outputs(2916) <= not (a or b);
    layer1_outputs(2917) <= b;
    layer1_outputs(2918) <= a or b;
    layer1_outputs(2919) <= '1';
    layer1_outputs(2920) <= b;
    layer1_outputs(2921) <= not (a and b);
    layer1_outputs(2922) <= not a;
    layer1_outputs(2923) <= not (a and b);
    layer1_outputs(2924) <= not b or a;
    layer1_outputs(2925) <= not a;
    layer1_outputs(2926) <= not b or a;
    layer1_outputs(2927) <= not b or a;
    layer1_outputs(2928) <= a and not b;
    layer1_outputs(2929) <= not a;
    layer1_outputs(2930) <= '0';
    layer1_outputs(2931) <= '1';
    layer1_outputs(2932) <= a and b;
    layer1_outputs(2933) <= not a;
    layer1_outputs(2934) <= '1';
    layer1_outputs(2935) <= not a;
    layer1_outputs(2936) <= a or b;
    layer1_outputs(2937) <= a;
    layer1_outputs(2938) <= a;
    layer1_outputs(2939) <= '0';
    layer1_outputs(2940) <= not (a and b);
    layer1_outputs(2941) <= not (a and b);
    layer1_outputs(2942) <= a or b;
    layer1_outputs(2943) <= a or b;
    layer1_outputs(2944) <= not b or a;
    layer1_outputs(2945) <= not a;
    layer1_outputs(2946) <= '1';
    layer1_outputs(2947) <= not b or a;
    layer1_outputs(2948) <= b;
    layer1_outputs(2949) <= '1';
    layer1_outputs(2950) <= not a;
    layer1_outputs(2951) <= not (a and b);
    layer1_outputs(2952) <= not b;
    layer1_outputs(2953) <= not a;
    layer1_outputs(2954) <= a and not b;
    layer1_outputs(2955) <= not b;
    layer1_outputs(2956) <= not a or b;
    layer1_outputs(2957) <= a and b;
    layer1_outputs(2958) <= not b or a;
    layer1_outputs(2959) <= not (a xor b);
    layer1_outputs(2960) <= not b;
    layer1_outputs(2961) <= a;
    layer1_outputs(2962) <= a or b;
    layer1_outputs(2963) <= '1';
    layer1_outputs(2964) <= not b or a;
    layer1_outputs(2965) <= not b or a;
    layer1_outputs(2966) <= '1';
    layer1_outputs(2967) <= a or b;
    layer1_outputs(2968) <= '1';
    layer1_outputs(2969) <= b;
    layer1_outputs(2970) <= b and not a;
    layer1_outputs(2971) <= '0';
    layer1_outputs(2972) <= not a or b;
    layer1_outputs(2973) <= '0';
    layer1_outputs(2974) <= a or b;
    layer1_outputs(2975) <= a and not b;
    layer1_outputs(2976) <= '1';
    layer1_outputs(2977) <= not b or a;
    layer1_outputs(2978) <= a and not b;
    layer1_outputs(2979) <= not (a and b);
    layer1_outputs(2980) <= not b;
    layer1_outputs(2981) <= a;
    layer1_outputs(2982) <= not b;
    layer1_outputs(2983) <= not (a and b);
    layer1_outputs(2984) <= not a or b;
    layer1_outputs(2985) <= a;
    layer1_outputs(2986) <= a;
    layer1_outputs(2987) <= not (a and b);
    layer1_outputs(2988) <= '1';
    layer1_outputs(2989) <= not (a or b);
    layer1_outputs(2990) <= not b or a;
    layer1_outputs(2991) <= a;
    layer1_outputs(2992) <= not b;
    layer1_outputs(2993) <= not (a or b);
    layer1_outputs(2994) <= not (a or b);
    layer1_outputs(2995) <= a and b;
    layer1_outputs(2996) <= '0';
    layer1_outputs(2997) <= a;
    layer1_outputs(2998) <= b and not a;
    layer1_outputs(2999) <= not b;
    layer1_outputs(3000) <= '1';
    layer1_outputs(3001) <= '0';
    layer1_outputs(3002) <= not a or b;
    layer1_outputs(3003) <= b;
    layer1_outputs(3004) <= not b;
    layer1_outputs(3005) <= not (a and b);
    layer1_outputs(3006) <= a and b;
    layer1_outputs(3007) <= not (a or b);
    layer1_outputs(3008) <= '1';
    layer1_outputs(3009) <= not a or b;
    layer1_outputs(3010) <= a;
    layer1_outputs(3011) <= '0';
    layer1_outputs(3012) <= a and b;
    layer1_outputs(3013) <= not (a or b);
    layer1_outputs(3014) <= not a;
    layer1_outputs(3015) <= not a or b;
    layer1_outputs(3016) <= not (a and b);
    layer1_outputs(3017) <= a or b;
    layer1_outputs(3018) <= b and not a;
    layer1_outputs(3019) <= not (a or b);
    layer1_outputs(3020) <= not a or b;
    layer1_outputs(3021) <= b;
    layer1_outputs(3022) <= '0';
    layer1_outputs(3023) <= not b;
    layer1_outputs(3024) <= not a or b;
    layer1_outputs(3025) <= a and not b;
    layer1_outputs(3026) <= b and not a;
    layer1_outputs(3027) <= a or b;
    layer1_outputs(3028) <= a xor b;
    layer1_outputs(3029) <= b;
    layer1_outputs(3030) <= not b or a;
    layer1_outputs(3031) <= not (a and b);
    layer1_outputs(3032) <= a and b;
    layer1_outputs(3033) <= not (a and b);
    layer1_outputs(3034) <= not b or a;
    layer1_outputs(3035) <= a or b;
    layer1_outputs(3036) <= a and not b;
    layer1_outputs(3037) <= '1';
    layer1_outputs(3038) <= not a;
    layer1_outputs(3039) <= a;
    layer1_outputs(3040) <= a;
    layer1_outputs(3041) <= b and not a;
    layer1_outputs(3042) <= a or b;
    layer1_outputs(3043) <= '1';
    layer1_outputs(3044) <= '1';
    layer1_outputs(3045) <= a and not b;
    layer1_outputs(3046) <= b;
    layer1_outputs(3047) <= '1';
    layer1_outputs(3048) <= b;
    layer1_outputs(3049) <= '0';
    layer1_outputs(3050) <= b and not a;
    layer1_outputs(3051) <= a and b;
    layer1_outputs(3052) <= not (a or b);
    layer1_outputs(3053) <= not (a or b);
    layer1_outputs(3054) <= a and b;
    layer1_outputs(3055) <= b and not a;
    layer1_outputs(3056) <= not b;
    layer1_outputs(3057) <= not b;
    layer1_outputs(3058) <= b;
    layer1_outputs(3059) <= b and not a;
    layer1_outputs(3060) <= not b;
    layer1_outputs(3061) <= a or b;
    layer1_outputs(3062) <= a and b;
    layer1_outputs(3063) <= b and not a;
    layer1_outputs(3064) <= '1';
    layer1_outputs(3065) <= not b;
    layer1_outputs(3066) <= a and not b;
    layer1_outputs(3067) <= b;
    layer1_outputs(3068) <= a and not b;
    layer1_outputs(3069) <= a;
    layer1_outputs(3070) <= not (a and b);
    layer1_outputs(3071) <= not a;
    layer1_outputs(3072) <= not b;
    layer1_outputs(3073) <= b;
    layer1_outputs(3074) <= not b or a;
    layer1_outputs(3075) <= '0';
    layer1_outputs(3076) <= b and not a;
    layer1_outputs(3077) <= not a or b;
    layer1_outputs(3078) <= not (a and b);
    layer1_outputs(3079) <= not a;
    layer1_outputs(3080) <= a;
    layer1_outputs(3081) <= b;
    layer1_outputs(3082) <= '1';
    layer1_outputs(3083) <= not b;
    layer1_outputs(3084) <= a and not b;
    layer1_outputs(3085) <= '1';
    layer1_outputs(3086) <= not a;
    layer1_outputs(3087) <= not b;
    layer1_outputs(3088) <= not a;
    layer1_outputs(3089) <= b and not a;
    layer1_outputs(3090) <= '1';
    layer1_outputs(3091) <= a;
    layer1_outputs(3092) <= a or b;
    layer1_outputs(3093) <= b;
    layer1_outputs(3094) <= not (a or b);
    layer1_outputs(3095) <= '1';
    layer1_outputs(3096) <= a and not b;
    layer1_outputs(3097) <= not (a and b);
    layer1_outputs(3098) <= a and b;
    layer1_outputs(3099) <= not (a or b);
    layer1_outputs(3100) <= '1';
    layer1_outputs(3101) <= '0';
    layer1_outputs(3102) <= not (a or b);
    layer1_outputs(3103) <= '0';
    layer1_outputs(3104) <= not (a and b);
    layer1_outputs(3105) <= not a;
    layer1_outputs(3106) <= a and b;
    layer1_outputs(3107) <= not b or a;
    layer1_outputs(3108) <= '0';
    layer1_outputs(3109) <= b and not a;
    layer1_outputs(3110) <= '1';
    layer1_outputs(3111) <= a and not b;
    layer1_outputs(3112) <= not (a and b);
    layer1_outputs(3113) <= not (a and b);
    layer1_outputs(3114) <= not a or b;
    layer1_outputs(3115) <= b;
    layer1_outputs(3116) <= a;
    layer1_outputs(3117) <= not a or b;
    layer1_outputs(3118) <= a and b;
    layer1_outputs(3119) <= a or b;
    layer1_outputs(3120) <= not b or a;
    layer1_outputs(3121) <= not (a and b);
    layer1_outputs(3122) <= a and not b;
    layer1_outputs(3123) <= not (a or b);
    layer1_outputs(3124) <= '1';
    layer1_outputs(3125) <= a or b;
    layer1_outputs(3126) <= not (a and b);
    layer1_outputs(3127) <= not a;
    layer1_outputs(3128) <= '1';
    layer1_outputs(3129) <= a or b;
    layer1_outputs(3130) <= '0';
    layer1_outputs(3131) <= b;
    layer1_outputs(3132) <= not (a and b);
    layer1_outputs(3133) <= b and not a;
    layer1_outputs(3134) <= a and not b;
    layer1_outputs(3135) <= not b;
    layer1_outputs(3136) <= not b;
    layer1_outputs(3137) <= not a;
    layer1_outputs(3138) <= b;
    layer1_outputs(3139) <= a and b;
    layer1_outputs(3140) <= a and b;
    layer1_outputs(3141) <= '1';
    layer1_outputs(3142) <= a or b;
    layer1_outputs(3143) <= '0';
    layer1_outputs(3144) <= not a or b;
    layer1_outputs(3145) <= '0';
    layer1_outputs(3146) <= not b or a;
    layer1_outputs(3147) <= not a or b;
    layer1_outputs(3148) <= a and not b;
    layer1_outputs(3149) <= not a or b;
    layer1_outputs(3150) <= a and b;
    layer1_outputs(3151) <= '1';
    layer1_outputs(3152) <= '0';
    layer1_outputs(3153) <= a and not b;
    layer1_outputs(3154) <= '0';
    layer1_outputs(3155) <= a or b;
    layer1_outputs(3156) <= not (a or b);
    layer1_outputs(3157) <= not a or b;
    layer1_outputs(3158) <= not (a or b);
    layer1_outputs(3159) <= '0';
    layer1_outputs(3160) <= not b;
    layer1_outputs(3161) <= '1';
    layer1_outputs(3162) <= not (a and b);
    layer1_outputs(3163) <= '0';
    layer1_outputs(3164) <= '1';
    layer1_outputs(3165) <= not (a and b);
    layer1_outputs(3166) <= a or b;
    layer1_outputs(3167) <= a and b;
    layer1_outputs(3168) <= not a or b;
    layer1_outputs(3169) <= not b or a;
    layer1_outputs(3170) <= not b;
    layer1_outputs(3171) <= not (a or b);
    layer1_outputs(3172) <= '1';
    layer1_outputs(3173) <= a;
    layer1_outputs(3174) <= not (a or b);
    layer1_outputs(3175) <= not b or a;
    layer1_outputs(3176) <= '0';
    layer1_outputs(3177) <= not b or a;
    layer1_outputs(3178) <= not a;
    layer1_outputs(3179) <= not (a or b);
    layer1_outputs(3180) <= a or b;
    layer1_outputs(3181) <= not (a or b);
    layer1_outputs(3182) <= not a or b;
    layer1_outputs(3183) <= '0';
    layer1_outputs(3184) <= not a or b;
    layer1_outputs(3185) <= not b;
    layer1_outputs(3186) <= not (a or b);
    layer1_outputs(3187) <= not (a and b);
    layer1_outputs(3188) <= not (a and b);
    layer1_outputs(3189) <= b;
    layer1_outputs(3190) <= b and not a;
    layer1_outputs(3191) <= not (a xor b);
    layer1_outputs(3192) <= not b or a;
    layer1_outputs(3193) <= a and not b;
    layer1_outputs(3194) <= not b or a;
    layer1_outputs(3195) <= not b;
    layer1_outputs(3196) <= not b or a;
    layer1_outputs(3197) <= '1';
    layer1_outputs(3198) <= a and not b;
    layer1_outputs(3199) <= a;
    layer1_outputs(3200) <= not (a or b);
    layer1_outputs(3201) <= a or b;
    layer1_outputs(3202) <= a or b;
    layer1_outputs(3203) <= '0';
    layer1_outputs(3204) <= a;
    layer1_outputs(3205) <= b and not a;
    layer1_outputs(3206) <= b and not a;
    layer1_outputs(3207) <= a and b;
    layer1_outputs(3208) <= not (a or b);
    layer1_outputs(3209) <= a or b;
    layer1_outputs(3210) <= not b or a;
    layer1_outputs(3211) <= a and not b;
    layer1_outputs(3212) <= b;
    layer1_outputs(3213) <= '0';
    layer1_outputs(3214) <= b and not a;
    layer1_outputs(3215) <= b;
    layer1_outputs(3216) <= a or b;
    layer1_outputs(3217) <= '0';
    layer1_outputs(3218) <= a and not b;
    layer1_outputs(3219) <= not (a and b);
    layer1_outputs(3220) <= '0';
    layer1_outputs(3221) <= not a or b;
    layer1_outputs(3222) <= a or b;
    layer1_outputs(3223) <= not (a or b);
    layer1_outputs(3224) <= not (a xor b);
    layer1_outputs(3225) <= not (a and b);
    layer1_outputs(3226) <= '1';
    layer1_outputs(3227) <= not (a and b);
    layer1_outputs(3228) <= '1';
    layer1_outputs(3229) <= not (a or b);
    layer1_outputs(3230) <= not (a and b);
    layer1_outputs(3231) <= '1';
    layer1_outputs(3232) <= not (a or b);
    layer1_outputs(3233) <= '1';
    layer1_outputs(3234) <= not a;
    layer1_outputs(3235) <= not a or b;
    layer1_outputs(3236) <= not (a or b);
    layer1_outputs(3237) <= not a;
    layer1_outputs(3238) <= b;
    layer1_outputs(3239) <= a and b;
    layer1_outputs(3240) <= a;
    layer1_outputs(3241) <= b;
    layer1_outputs(3242) <= a xor b;
    layer1_outputs(3243) <= '0';
    layer1_outputs(3244) <= b;
    layer1_outputs(3245) <= not b or a;
    layer1_outputs(3246) <= '0';
    layer1_outputs(3247) <= not b;
    layer1_outputs(3248) <= a or b;
    layer1_outputs(3249) <= a and not b;
    layer1_outputs(3250) <= b and not a;
    layer1_outputs(3251) <= not b;
    layer1_outputs(3252) <= '0';
    layer1_outputs(3253) <= not (a and b);
    layer1_outputs(3254) <= b;
    layer1_outputs(3255) <= b and not a;
    layer1_outputs(3256) <= '1';
    layer1_outputs(3257) <= not b or a;
    layer1_outputs(3258) <= not b or a;
    layer1_outputs(3259) <= not (a or b);
    layer1_outputs(3260) <= '0';
    layer1_outputs(3261) <= not a or b;
    layer1_outputs(3262) <= '0';
    layer1_outputs(3263) <= a and b;
    layer1_outputs(3264) <= '0';
    layer1_outputs(3265) <= a;
    layer1_outputs(3266) <= a and b;
    layer1_outputs(3267) <= '0';
    layer1_outputs(3268) <= a or b;
    layer1_outputs(3269) <= a and b;
    layer1_outputs(3270) <= b and not a;
    layer1_outputs(3271) <= a and not b;
    layer1_outputs(3272) <= b;
    layer1_outputs(3273) <= not (a and b);
    layer1_outputs(3274) <= not b;
    layer1_outputs(3275) <= not a or b;
    layer1_outputs(3276) <= a;
    layer1_outputs(3277) <= not b or a;
    layer1_outputs(3278) <= not (a xor b);
    layer1_outputs(3279) <= '0';
    layer1_outputs(3280) <= not (a or b);
    layer1_outputs(3281) <= not a or b;
    layer1_outputs(3282) <= not b or a;
    layer1_outputs(3283) <= not a;
    layer1_outputs(3284) <= not (a and b);
    layer1_outputs(3285) <= a or b;
    layer1_outputs(3286) <= b;
    layer1_outputs(3287) <= '1';
    layer1_outputs(3288) <= not b;
    layer1_outputs(3289) <= '1';
    layer1_outputs(3290) <= b and not a;
    layer1_outputs(3291) <= not a or b;
    layer1_outputs(3292) <= a;
    layer1_outputs(3293) <= '1';
    layer1_outputs(3294) <= a;
    layer1_outputs(3295) <= not a or b;
    layer1_outputs(3296) <= a;
    layer1_outputs(3297) <= a and not b;
    layer1_outputs(3298) <= not b or a;
    layer1_outputs(3299) <= a and not b;
    layer1_outputs(3300) <= '0';
    layer1_outputs(3301) <= not (a or b);
    layer1_outputs(3302) <= a or b;
    layer1_outputs(3303) <= '1';
    layer1_outputs(3304) <= not (a xor b);
    layer1_outputs(3305) <= '1';
    layer1_outputs(3306) <= not b;
    layer1_outputs(3307) <= b and not a;
    layer1_outputs(3308) <= not (a or b);
    layer1_outputs(3309) <= not a or b;
    layer1_outputs(3310) <= not (a or b);
    layer1_outputs(3311) <= not (a xor b);
    layer1_outputs(3312) <= '0';
    layer1_outputs(3313) <= not (a or b);
    layer1_outputs(3314) <= not (a and b);
    layer1_outputs(3315) <= not a;
    layer1_outputs(3316) <= not (a or b);
    layer1_outputs(3317) <= not a;
    layer1_outputs(3318) <= b;
    layer1_outputs(3319) <= a or b;
    layer1_outputs(3320) <= a and b;
    layer1_outputs(3321) <= a;
    layer1_outputs(3322) <= a or b;
    layer1_outputs(3323) <= b and not a;
    layer1_outputs(3324) <= not (a or b);
    layer1_outputs(3325) <= not b or a;
    layer1_outputs(3326) <= not b;
    layer1_outputs(3327) <= not a;
    layer1_outputs(3328) <= a;
    layer1_outputs(3329) <= '0';
    layer1_outputs(3330) <= not (a or b);
    layer1_outputs(3331) <= b and not a;
    layer1_outputs(3332) <= a and not b;
    layer1_outputs(3333) <= not b or a;
    layer1_outputs(3334) <= b;
    layer1_outputs(3335) <= a and not b;
    layer1_outputs(3336) <= '1';
    layer1_outputs(3337) <= a or b;
    layer1_outputs(3338) <= a and not b;
    layer1_outputs(3339) <= b;
    layer1_outputs(3340) <= not (a and b);
    layer1_outputs(3341) <= a and b;
    layer1_outputs(3342) <= not (a or b);
    layer1_outputs(3343) <= not a;
    layer1_outputs(3344) <= not a;
    layer1_outputs(3345) <= a;
    layer1_outputs(3346) <= a;
    layer1_outputs(3347) <= '0';
    layer1_outputs(3348) <= not (a and b);
    layer1_outputs(3349) <= '0';
    layer1_outputs(3350) <= a or b;
    layer1_outputs(3351) <= not b or a;
    layer1_outputs(3352) <= b;
    layer1_outputs(3353) <= a and not b;
    layer1_outputs(3354) <= not b;
    layer1_outputs(3355) <= not (a or b);
    layer1_outputs(3356) <= a;
    layer1_outputs(3357) <= not a;
    layer1_outputs(3358) <= not b or a;
    layer1_outputs(3359) <= a or b;
    layer1_outputs(3360) <= '1';
    layer1_outputs(3361) <= '0';
    layer1_outputs(3362) <= b and not a;
    layer1_outputs(3363) <= '1';
    layer1_outputs(3364) <= a and b;
    layer1_outputs(3365) <= '1';
    layer1_outputs(3366) <= not a or b;
    layer1_outputs(3367) <= not (a xor b);
    layer1_outputs(3368) <= not (a xor b);
    layer1_outputs(3369) <= not (a and b);
    layer1_outputs(3370) <= not b;
    layer1_outputs(3371) <= a or b;
    layer1_outputs(3372) <= not a or b;
    layer1_outputs(3373) <= a;
    layer1_outputs(3374) <= a;
    layer1_outputs(3375) <= a or b;
    layer1_outputs(3376) <= not b or a;
    layer1_outputs(3377) <= a and b;
    layer1_outputs(3378) <= not (a or b);
    layer1_outputs(3379) <= not (a and b);
    layer1_outputs(3380) <= '0';
    layer1_outputs(3381) <= b and not a;
    layer1_outputs(3382) <= '0';
    layer1_outputs(3383) <= '0';
    layer1_outputs(3384) <= a or b;
    layer1_outputs(3385) <= b and not a;
    layer1_outputs(3386) <= not (a or b);
    layer1_outputs(3387) <= a xor b;
    layer1_outputs(3388) <= not b or a;
    layer1_outputs(3389) <= '1';
    layer1_outputs(3390) <= '1';
    layer1_outputs(3391) <= '1';
    layer1_outputs(3392) <= '0';
    layer1_outputs(3393) <= a or b;
    layer1_outputs(3394) <= a;
    layer1_outputs(3395) <= not (a and b);
    layer1_outputs(3396) <= '0';
    layer1_outputs(3397) <= '1';
    layer1_outputs(3398) <= b;
    layer1_outputs(3399) <= not a or b;
    layer1_outputs(3400) <= not (a and b);
    layer1_outputs(3401) <= not b or a;
    layer1_outputs(3402) <= '0';
    layer1_outputs(3403) <= not (a xor b);
    layer1_outputs(3404) <= not a;
    layer1_outputs(3405) <= a and not b;
    layer1_outputs(3406) <= b;
    layer1_outputs(3407) <= not a or b;
    layer1_outputs(3408) <= '1';
    layer1_outputs(3409) <= not (a and b);
    layer1_outputs(3410) <= not (a and b);
    layer1_outputs(3411) <= not (a xor b);
    layer1_outputs(3412) <= not a or b;
    layer1_outputs(3413) <= '1';
    layer1_outputs(3414) <= not (a and b);
    layer1_outputs(3415) <= '1';
    layer1_outputs(3416) <= a and b;
    layer1_outputs(3417) <= '0';
    layer1_outputs(3418) <= not (a and b);
    layer1_outputs(3419) <= not b or a;
    layer1_outputs(3420) <= not (a and b);
    layer1_outputs(3421) <= not b;
    layer1_outputs(3422) <= '0';
    layer1_outputs(3423) <= not (a or b);
    layer1_outputs(3424) <= not b or a;
    layer1_outputs(3425) <= not a;
    layer1_outputs(3426) <= not b or a;
    layer1_outputs(3427) <= '1';
    layer1_outputs(3428) <= not (a or b);
    layer1_outputs(3429) <= a xor b;
    layer1_outputs(3430) <= not (a and b);
    layer1_outputs(3431) <= not b or a;
    layer1_outputs(3432) <= '1';
    layer1_outputs(3433) <= not a;
    layer1_outputs(3434) <= a and not b;
    layer1_outputs(3435) <= not a;
    layer1_outputs(3436) <= a or b;
    layer1_outputs(3437) <= not b or a;
    layer1_outputs(3438) <= b;
    layer1_outputs(3439) <= '0';
    layer1_outputs(3440) <= b;
    layer1_outputs(3441) <= not a;
    layer1_outputs(3442) <= a and not b;
    layer1_outputs(3443) <= '1';
    layer1_outputs(3444) <= a and b;
    layer1_outputs(3445) <= not (a and b);
    layer1_outputs(3446) <= not b;
    layer1_outputs(3447) <= '0';
    layer1_outputs(3448) <= a;
    layer1_outputs(3449) <= not (a xor b);
    layer1_outputs(3450) <= b;
    layer1_outputs(3451) <= b and not a;
    layer1_outputs(3452) <= not a or b;
    layer1_outputs(3453) <= a;
    layer1_outputs(3454) <= '0';
    layer1_outputs(3455) <= '1';
    layer1_outputs(3456) <= a;
    layer1_outputs(3457) <= '1';
    layer1_outputs(3458) <= a or b;
    layer1_outputs(3459) <= not a;
    layer1_outputs(3460) <= b and not a;
    layer1_outputs(3461) <= not (a and b);
    layer1_outputs(3462) <= a;
    layer1_outputs(3463) <= not a or b;
    layer1_outputs(3464) <= a or b;
    layer1_outputs(3465) <= not a;
    layer1_outputs(3466) <= not b;
    layer1_outputs(3467) <= not a or b;
    layer1_outputs(3468) <= not a or b;
    layer1_outputs(3469) <= not (a or b);
    layer1_outputs(3470) <= b;
    layer1_outputs(3471) <= '0';
    layer1_outputs(3472) <= b;
    layer1_outputs(3473) <= not b or a;
    layer1_outputs(3474) <= not a or b;
    layer1_outputs(3475) <= not (a and b);
    layer1_outputs(3476) <= a or b;
    layer1_outputs(3477) <= a;
    layer1_outputs(3478) <= a or b;
    layer1_outputs(3479) <= a and not b;
    layer1_outputs(3480) <= '1';
    layer1_outputs(3481) <= not (a and b);
    layer1_outputs(3482) <= not (a or b);
    layer1_outputs(3483) <= not a or b;
    layer1_outputs(3484) <= '1';
    layer1_outputs(3485) <= b and not a;
    layer1_outputs(3486) <= a xor b;
    layer1_outputs(3487) <= '1';
    layer1_outputs(3488) <= a and b;
    layer1_outputs(3489) <= not b;
    layer1_outputs(3490) <= not b;
    layer1_outputs(3491) <= a and b;
    layer1_outputs(3492) <= not (a or b);
    layer1_outputs(3493) <= not b or a;
    layer1_outputs(3494) <= not b;
    layer1_outputs(3495) <= a or b;
    layer1_outputs(3496) <= not (a or b);
    layer1_outputs(3497) <= a and b;
    layer1_outputs(3498) <= not a;
    layer1_outputs(3499) <= '1';
    layer1_outputs(3500) <= not a or b;
    layer1_outputs(3501) <= not (a or b);
    layer1_outputs(3502) <= not a;
    layer1_outputs(3503) <= not a or b;
    layer1_outputs(3504) <= not (a xor b);
    layer1_outputs(3505) <= a and not b;
    layer1_outputs(3506) <= not a;
    layer1_outputs(3507) <= a or b;
    layer1_outputs(3508) <= not (a and b);
    layer1_outputs(3509) <= not (a and b);
    layer1_outputs(3510) <= not a or b;
    layer1_outputs(3511) <= not (a and b);
    layer1_outputs(3512) <= b and not a;
    layer1_outputs(3513) <= b and not a;
    layer1_outputs(3514) <= '0';
    layer1_outputs(3515) <= not (a or b);
    layer1_outputs(3516) <= b;
    layer1_outputs(3517) <= not b;
    layer1_outputs(3518) <= not (a and b);
    layer1_outputs(3519) <= b and not a;
    layer1_outputs(3520) <= b;
    layer1_outputs(3521) <= not (a or b);
    layer1_outputs(3522) <= a and not b;
    layer1_outputs(3523) <= not b;
    layer1_outputs(3524) <= not a or b;
    layer1_outputs(3525) <= b;
    layer1_outputs(3526) <= a and b;
    layer1_outputs(3527) <= '1';
    layer1_outputs(3528) <= not a;
    layer1_outputs(3529) <= not (a or b);
    layer1_outputs(3530) <= a;
    layer1_outputs(3531) <= not b or a;
    layer1_outputs(3532) <= not a;
    layer1_outputs(3533) <= a and b;
    layer1_outputs(3534) <= not a;
    layer1_outputs(3535) <= a xor b;
    layer1_outputs(3536) <= not (a and b);
    layer1_outputs(3537) <= a;
    layer1_outputs(3538) <= not b or a;
    layer1_outputs(3539) <= a or b;
    layer1_outputs(3540) <= '0';
    layer1_outputs(3541) <= '1';
    layer1_outputs(3542) <= '0';
    layer1_outputs(3543) <= a;
    layer1_outputs(3544) <= a and not b;
    layer1_outputs(3545) <= a or b;
    layer1_outputs(3546) <= a xor b;
    layer1_outputs(3547) <= a or b;
    layer1_outputs(3548) <= a or b;
    layer1_outputs(3549) <= not b;
    layer1_outputs(3550) <= not a;
    layer1_outputs(3551) <= not b or a;
    layer1_outputs(3552) <= a and not b;
    layer1_outputs(3553) <= '0';
    layer1_outputs(3554) <= '0';
    layer1_outputs(3555) <= '0';
    layer1_outputs(3556) <= not b or a;
    layer1_outputs(3557) <= not b;
    layer1_outputs(3558) <= not b;
    layer1_outputs(3559) <= not a or b;
    layer1_outputs(3560) <= not b;
    layer1_outputs(3561) <= b;
    layer1_outputs(3562) <= not b or a;
    layer1_outputs(3563) <= not (a and b);
    layer1_outputs(3564) <= '1';
    layer1_outputs(3565) <= not a;
    layer1_outputs(3566) <= b and not a;
    layer1_outputs(3567) <= a;
    layer1_outputs(3568) <= '0';
    layer1_outputs(3569) <= b and not a;
    layer1_outputs(3570) <= '1';
    layer1_outputs(3571) <= '1';
    layer1_outputs(3572) <= b and not a;
    layer1_outputs(3573) <= not a;
    layer1_outputs(3574) <= a and not b;
    layer1_outputs(3575) <= '0';
    layer1_outputs(3576) <= a and not b;
    layer1_outputs(3577) <= '1';
    layer1_outputs(3578) <= b;
    layer1_outputs(3579) <= a and b;
    layer1_outputs(3580) <= not a or b;
    layer1_outputs(3581) <= '0';
    layer1_outputs(3582) <= not (a or b);
    layer1_outputs(3583) <= b and not a;
    layer1_outputs(3584) <= b;
    layer1_outputs(3585) <= '0';
    layer1_outputs(3586) <= a and not b;
    layer1_outputs(3587) <= a;
    layer1_outputs(3588) <= a and b;
    layer1_outputs(3589) <= not b or a;
    layer1_outputs(3590) <= '1';
    layer1_outputs(3591) <= '1';
    layer1_outputs(3592) <= b;
    layer1_outputs(3593) <= '0';
    layer1_outputs(3594) <= b and not a;
    layer1_outputs(3595) <= not b or a;
    layer1_outputs(3596) <= b;
    layer1_outputs(3597) <= b;
    layer1_outputs(3598) <= not b or a;
    layer1_outputs(3599) <= not (a or b);
    layer1_outputs(3600) <= not (a or b);
    layer1_outputs(3601) <= a xor b;
    layer1_outputs(3602) <= not (a or b);
    layer1_outputs(3603) <= b and not a;
    layer1_outputs(3604) <= b and not a;
    layer1_outputs(3605) <= b and not a;
    layer1_outputs(3606) <= b and not a;
    layer1_outputs(3607) <= '1';
    layer1_outputs(3608) <= not a;
    layer1_outputs(3609) <= a and b;
    layer1_outputs(3610) <= b and not a;
    layer1_outputs(3611) <= not b or a;
    layer1_outputs(3612) <= '1';
    layer1_outputs(3613) <= '0';
    layer1_outputs(3614) <= not (a and b);
    layer1_outputs(3615) <= '1';
    layer1_outputs(3616) <= not b;
    layer1_outputs(3617) <= a and not b;
    layer1_outputs(3618) <= b;
    layer1_outputs(3619) <= a and b;
    layer1_outputs(3620) <= not b or a;
    layer1_outputs(3621) <= not (a or b);
    layer1_outputs(3622) <= '0';
    layer1_outputs(3623) <= a;
    layer1_outputs(3624) <= not (a and b);
    layer1_outputs(3625) <= not (a or b);
    layer1_outputs(3626) <= not (a and b);
    layer1_outputs(3627) <= b;
    layer1_outputs(3628) <= b;
    layer1_outputs(3629) <= a and not b;
    layer1_outputs(3630) <= a and not b;
    layer1_outputs(3631) <= a and not b;
    layer1_outputs(3632) <= a and b;
    layer1_outputs(3633) <= b and not a;
    layer1_outputs(3634) <= '1';
    layer1_outputs(3635) <= not b or a;
    layer1_outputs(3636) <= b and not a;
    layer1_outputs(3637) <= a and b;
    layer1_outputs(3638) <= a;
    layer1_outputs(3639) <= '1';
    layer1_outputs(3640) <= a;
    layer1_outputs(3641) <= a xor b;
    layer1_outputs(3642) <= not (a and b);
    layer1_outputs(3643) <= not (a or b);
    layer1_outputs(3644) <= a;
    layer1_outputs(3645) <= '1';
    layer1_outputs(3646) <= a;
    layer1_outputs(3647) <= not a or b;
    layer1_outputs(3648) <= b;
    layer1_outputs(3649) <= '0';
    layer1_outputs(3650) <= b;
    layer1_outputs(3651) <= not (a or b);
    layer1_outputs(3652) <= b;
    layer1_outputs(3653) <= b;
    layer1_outputs(3654) <= '0';
    layer1_outputs(3655) <= b;
    layer1_outputs(3656) <= not a or b;
    layer1_outputs(3657) <= not b;
    layer1_outputs(3658) <= b and not a;
    layer1_outputs(3659) <= b and not a;
    layer1_outputs(3660) <= '0';
    layer1_outputs(3661) <= a or b;
    layer1_outputs(3662) <= a or b;
    layer1_outputs(3663) <= not b or a;
    layer1_outputs(3664) <= a;
    layer1_outputs(3665) <= a and b;
    layer1_outputs(3666) <= '1';
    layer1_outputs(3667) <= a or b;
    layer1_outputs(3668) <= not (a xor b);
    layer1_outputs(3669) <= b;
    layer1_outputs(3670) <= not a or b;
    layer1_outputs(3671) <= not a or b;
    layer1_outputs(3672) <= '1';
    layer1_outputs(3673) <= not b or a;
    layer1_outputs(3674) <= b;
    layer1_outputs(3675) <= b and not a;
    layer1_outputs(3676) <= not (a or b);
    layer1_outputs(3677) <= '0';
    layer1_outputs(3678) <= '0';
    layer1_outputs(3679) <= a;
    layer1_outputs(3680) <= a;
    layer1_outputs(3681) <= a and b;
    layer1_outputs(3682) <= a;
    layer1_outputs(3683) <= not a or b;
    layer1_outputs(3684) <= a or b;
    layer1_outputs(3685) <= '1';
    layer1_outputs(3686) <= not (a and b);
    layer1_outputs(3687) <= not a;
    layer1_outputs(3688) <= not (a xor b);
    layer1_outputs(3689) <= b;
    layer1_outputs(3690) <= b and not a;
    layer1_outputs(3691) <= b and not a;
    layer1_outputs(3692) <= not b;
    layer1_outputs(3693) <= a or b;
    layer1_outputs(3694) <= '0';
    layer1_outputs(3695) <= '0';
    layer1_outputs(3696) <= not a;
    layer1_outputs(3697) <= b and not a;
    layer1_outputs(3698) <= b;
    layer1_outputs(3699) <= '0';
    layer1_outputs(3700) <= not a;
    layer1_outputs(3701) <= a and not b;
    layer1_outputs(3702) <= a xor b;
    layer1_outputs(3703) <= '1';
    layer1_outputs(3704) <= b;
    layer1_outputs(3705) <= not b or a;
    layer1_outputs(3706) <= a or b;
    layer1_outputs(3707) <= '0';
    layer1_outputs(3708) <= not a;
    layer1_outputs(3709) <= a or b;
    layer1_outputs(3710) <= b;
    layer1_outputs(3711) <= not (a or b);
    layer1_outputs(3712) <= not b or a;
    layer1_outputs(3713) <= '1';
    layer1_outputs(3714) <= '0';
    layer1_outputs(3715) <= not b;
    layer1_outputs(3716) <= not a or b;
    layer1_outputs(3717) <= not (a or b);
    layer1_outputs(3718) <= not a or b;
    layer1_outputs(3719) <= not b;
    layer1_outputs(3720) <= a and b;
    layer1_outputs(3721) <= '1';
    layer1_outputs(3722) <= a xor b;
    layer1_outputs(3723) <= a;
    layer1_outputs(3724) <= not a;
    layer1_outputs(3725) <= not b or a;
    layer1_outputs(3726) <= a or b;
    layer1_outputs(3727) <= not a;
    layer1_outputs(3728) <= not a or b;
    layer1_outputs(3729) <= not b or a;
    layer1_outputs(3730) <= a and not b;
    layer1_outputs(3731) <= not (a and b);
    layer1_outputs(3732) <= not b;
    layer1_outputs(3733) <= b and not a;
    layer1_outputs(3734) <= not b or a;
    layer1_outputs(3735) <= '1';
    layer1_outputs(3736) <= '1';
    layer1_outputs(3737) <= b;
    layer1_outputs(3738) <= a and b;
    layer1_outputs(3739) <= a and b;
    layer1_outputs(3740) <= '0';
    layer1_outputs(3741) <= not b;
    layer1_outputs(3742) <= a;
    layer1_outputs(3743) <= not b;
    layer1_outputs(3744) <= not a;
    layer1_outputs(3745) <= not b;
    layer1_outputs(3746) <= not b;
    layer1_outputs(3747) <= not b or a;
    layer1_outputs(3748) <= not b or a;
    layer1_outputs(3749) <= not a;
    layer1_outputs(3750) <= '0';
    layer1_outputs(3751) <= a;
    layer1_outputs(3752) <= not b or a;
    layer1_outputs(3753) <= not (a xor b);
    layer1_outputs(3754) <= b and not a;
    layer1_outputs(3755) <= not a or b;
    layer1_outputs(3756) <= not a;
    layer1_outputs(3757) <= not b or a;
    layer1_outputs(3758) <= a or b;
    layer1_outputs(3759) <= b and not a;
    layer1_outputs(3760) <= not b;
    layer1_outputs(3761) <= not a;
    layer1_outputs(3762) <= not b;
    layer1_outputs(3763) <= not (a and b);
    layer1_outputs(3764) <= '0';
    layer1_outputs(3765) <= '0';
    layer1_outputs(3766) <= b and not a;
    layer1_outputs(3767) <= '1';
    layer1_outputs(3768) <= not (a or b);
    layer1_outputs(3769) <= a or b;
    layer1_outputs(3770) <= a and b;
    layer1_outputs(3771) <= not b;
    layer1_outputs(3772) <= not (a and b);
    layer1_outputs(3773) <= not a;
    layer1_outputs(3774) <= not b;
    layer1_outputs(3775) <= '0';
    layer1_outputs(3776) <= b and not a;
    layer1_outputs(3777) <= not a or b;
    layer1_outputs(3778) <= a;
    layer1_outputs(3779) <= not b;
    layer1_outputs(3780) <= '1';
    layer1_outputs(3781) <= '1';
    layer1_outputs(3782) <= '1';
    layer1_outputs(3783) <= not (a xor b);
    layer1_outputs(3784) <= a and not b;
    layer1_outputs(3785) <= not a;
    layer1_outputs(3786) <= b and not a;
    layer1_outputs(3787) <= not (a and b);
    layer1_outputs(3788) <= b;
    layer1_outputs(3789) <= a;
    layer1_outputs(3790) <= not b;
    layer1_outputs(3791) <= b;
    layer1_outputs(3792) <= a;
    layer1_outputs(3793) <= not b;
    layer1_outputs(3794) <= a or b;
    layer1_outputs(3795) <= not (a or b);
    layer1_outputs(3796) <= b;
    layer1_outputs(3797) <= b and not a;
    layer1_outputs(3798) <= a or b;
    layer1_outputs(3799) <= b;
    layer1_outputs(3800) <= '0';
    layer1_outputs(3801) <= b and not a;
    layer1_outputs(3802) <= a and not b;
    layer1_outputs(3803) <= '0';
    layer1_outputs(3804) <= a and b;
    layer1_outputs(3805) <= not a;
    layer1_outputs(3806) <= '0';
    layer1_outputs(3807) <= not (a and b);
    layer1_outputs(3808) <= not a or b;
    layer1_outputs(3809) <= b and not a;
    layer1_outputs(3810) <= '0';
    layer1_outputs(3811) <= not a;
    layer1_outputs(3812) <= not a or b;
    layer1_outputs(3813) <= not (a or b);
    layer1_outputs(3814) <= '1';
    layer1_outputs(3815) <= a;
    layer1_outputs(3816) <= '1';
    layer1_outputs(3817) <= '1';
    layer1_outputs(3818) <= '1';
    layer1_outputs(3819) <= not a;
    layer1_outputs(3820) <= b;
    layer1_outputs(3821) <= '1';
    layer1_outputs(3822) <= not (a or b);
    layer1_outputs(3823) <= not b;
    layer1_outputs(3824) <= not (a or b);
    layer1_outputs(3825) <= a and not b;
    layer1_outputs(3826) <= not (a or b);
    layer1_outputs(3827) <= not a;
    layer1_outputs(3828) <= not (a and b);
    layer1_outputs(3829) <= not (a or b);
    layer1_outputs(3830) <= '0';
    layer1_outputs(3831) <= b and not a;
    layer1_outputs(3832) <= a or b;
    layer1_outputs(3833) <= not (a or b);
    layer1_outputs(3834) <= '1';
    layer1_outputs(3835) <= a;
    layer1_outputs(3836) <= not (a or b);
    layer1_outputs(3837) <= not b or a;
    layer1_outputs(3838) <= not b or a;
    layer1_outputs(3839) <= b and not a;
    layer1_outputs(3840) <= not b;
    layer1_outputs(3841) <= a and b;
    layer1_outputs(3842) <= '0';
    layer1_outputs(3843) <= b and not a;
    layer1_outputs(3844) <= '1';
    layer1_outputs(3845) <= not a;
    layer1_outputs(3846) <= a or b;
    layer1_outputs(3847) <= not a or b;
    layer1_outputs(3848) <= a;
    layer1_outputs(3849) <= not (a or b);
    layer1_outputs(3850) <= not (a and b);
    layer1_outputs(3851) <= not b or a;
    layer1_outputs(3852) <= b;
    layer1_outputs(3853) <= a and b;
    layer1_outputs(3854) <= a and b;
    layer1_outputs(3855) <= not a or b;
    layer1_outputs(3856) <= b and not a;
    layer1_outputs(3857) <= '0';
    layer1_outputs(3858) <= not a or b;
    layer1_outputs(3859) <= a and b;
    layer1_outputs(3860) <= a or b;
    layer1_outputs(3861) <= '1';
    layer1_outputs(3862) <= not (a and b);
    layer1_outputs(3863) <= not (a or b);
    layer1_outputs(3864) <= not (a and b);
    layer1_outputs(3865) <= not a or b;
    layer1_outputs(3866) <= not (a and b);
    layer1_outputs(3867) <= not b or a;
    layer1_outputs(3868) <= not b or a;
    layer1_outputs(3869) <= not a;
    layer1_outputs(3870) <= a or b;
    layer1_outputs(3871) <= a xor b;
    layer1_outputs(3872) <= b and not a;
    layer1_outputs(3873) <= a xor b;
    layer1_outputs(3874) <= '0';
    layer1_outputs(3875) <= not (a and b);
    layer1_outputs(3876) <= a xor b;
    layer1_outputs(3877) <= not b;
    layer1_outputs(3878) <= '1';
    layer1_outputs(3879) <= b;
    layer1_outputs(3880) <= '0';
    layer1_outputs(3881) <= '0';
    layer1_outputs(3882) <= not (a and b);
    layer1_outputs(3883) <= a;
    layer1_outputs(3884) <= a;
    layer1_outputs(3885) <= not a or b;
    layer1_outputs(3886) <= '1';
    layer1_outputs(3887) <= not a or b;
    layer1_outputs(3888) <= b;
    layer1_outputs(3889) <= a or b;
    layer1_outputs(3890) <= a or b;
    layer1_outputs(3891) <= not a;
    layer1_outputs(3892) <= '1';
    layer1_outputs(3893) <= not a;
    layer1_outputs(3894) <= a and b;
    layer1_outputs(3895) <= '1';
    layer1_outputs(3896) <= not (a and b);
    layer1_outputs(3897) <= a and b;
    layer1_outputs(3898) <= not a;
    layer1_outputs(3899) <= a and not b;
    layer1_outputs(3900) <= b and not a;
    layer1_outputs(3901) <= a and not b;
    layer1_outputs(3902) <= '1';
    layer1_outputs(3903) <= a and b;
    layer1_outputs(3904) <= not a;
    layer1_outputs(3905) <= not a;
    layer1_outputs(3906) <= '1';
    layer1_outputs(3907) <= a or b;
    layer1_outputs(3908) <= a xor b;
    layer1_outputs(3909) <= not b;
    layer1_outputs(3910) <= not (a and b);
    layer1_outputs(3911) <= a or b;
    layer1_outputs(3912) <= not b;
    layer1_outputs(3913) <= b;
    layer1_outputs(3914) <= not a or b;
    layer1_outputs(3915) <= not (a or b);
    layer1_outputs(3916) <= a or b;
    layer1_outputs(3917) <= '0';
    layer1_outputs(3918) <= a;
    layer1_outputs(3919) <= '1';
    layer1_outputs(3920) <= not b;
    layer1_outputs(3921) <= a or b;
    layer1_outputs(3922) <= not (a and b);
    layer1_outputs(3923) <= '1';
    layer1_outputs(3924) <= not (a and b);
    layer1_outputs(3925) <= a or b;
    layer1_outputs(3926) <= '0';
    layer1_outputs(3927) <= a;
    layer1_outputs(3928) <= not a;
    layer1_outputs(3929) <= '0';
    layer1_outputs(3930) <= not a or b;
    layer1_outputs(3931) <= a and b;
    layer1_outputs(3932) <= '1';
    layer1_outputs(3933) <= a and not b;
    layer1_outputs(3934) <= not a;
    layer1_outputs(3935) <= '1';
    layer1_outputs(3936) <= not a;
    layer1_outputs(3937) <= not a;
    layer1_outputs(3938) <= a and not b;
    layer1_outputs(3939) <= a and b;
    layer1_outputs(3940) <= not a;
    layer1_outputs(3941) <= a;
    layer1_outputs(3942) <= not b;
    layer1_outputs(3943) <= b and not a;
    layer1_outputs(3944) <= not b or a;
    layer1_outputs(3945) <= a or b;
    layer1_outputs(3946) <= not (a and b);
    layer1_outputs(3947) <= '0';
    layer1_outputs(3948) <= not (a or b);
    layer1_outputs(3949) <= '1';
    layer1_outputs(3950) <= not (a or b);
    layer1_outputs(3951) <= a;
    layer1_outputs(3952) <= not (a and b);
    layer1_outputs(3953) <= b and not a;
    layer1_outputs(3954) <= a;
    layer1_outputs(3955) <= b and not a;
    layer1_outputs(3956) <= a xor b;
    layer1_outputs(3957) <= b;
    layer1_outputs(3958) <= not b or a;
    layer1_outputs(3959) <= b and not a;
    layer1_outputs(3960) <= a and b;
    layer1_outputs(3961) <= '0';
    layer1_outputs(3962) <= a;
    layer1_outputs(3963) <= not (a or b);
    layer1_outputs(3964) <= a or b;
    layer1_outputs(3965) <= '1';
    layer1_outputs(3966) <= not (a xor b);
    layer1_outputs(3967) <= not a;
    layer1_outputs(3968) <= '0';
    layer1_outputs(3969) <= '1';
    layer1_outputs(3970) <= not (a and b);
    layer1_outputs(3971) <= '1';
    layer1_outputs(3972) <= not a or b;
    layer1_outputs(3973) <= not b or a;
    layer1_outputs(3974) <= a and b;
    layer1_outputs(3975) <= a or b;
    layer1_outputs(3976) <= not a or b;
    layer1_outputs(3977) <= a and b;
    layer1_outputs(3978) <= not b;
    layer1_outputs(3979) <= '0';
    layer1_outputs(3980) <= not (a and b);
    layer1_outputs(3981) <= '1';
    layer1_outputs(3982) <= a and not b;
    layer1_outputs(3983) <= not b;
    layer1_outputs(3984) <= b and not a;
    layer1_outputs(3985) <= a;
    layer1_outputs(3986) <= a;
    layer1_outputs(3987) <= a and not b;
    layer1_outputs(3988) <= b and not a;
    layer1_outputs(3989) <= b;
    layer1_outputs(3990) <= not (a or b);
    layer1_outputs(3991) <= not (a or b);
    layer1_outputs(3992) <= not b or a;
    layer1_outputs(3993) <= a and b;
    layer1_outputs(3994) <= not b or a;
    layer1_outputs(3995) <= not (a or b);
    layer1_outputs(3996) <= not b;
    layer1_outputs(3997) <= b;
    layer1_outputs(3998) <= not a;
    layer1_outputs(3999) <= a and b;
    layer1_outputs(4000) <= b;
    layer1_outputs(4001) <= b and not a;
    layer1_outputs(4002) <= a and not b;
    layer1_outputs(4003) <= not (a or b);
    layer1_outputs(4004) <= not (a or b);
    layer1_outputs(4005) <= '1';
    layer1_outputs(4006) <= not b or a;
    layer1_outputs(4007) <= not (a and b);
    layer1_outputs(4008) <= '1';
    layer1_outputs(4009) <= not (a and b);
    layer1_outputs(4010) <= a;
    layer1_outputs(4011) <= a and not b;
    layer1_outputs(4012) <= a and not b;
    layer1_outputs(4013) <= a and not b;
    layer1_outputs(4014) <= a;
    layer1_outputs(4015) <= not (a and b);
    layer1_outputs(4016) <= not (a or b);
    layer1_outputs(4017) <= not b;
    layer1_outputs(4018) <= b and not a;
    layer1_outputs(4019) <= a xor b;
    layer1_outputs(4020) <= not b or a;
    layer1_outputs(4021) <= '1';
    layer1_outputs(4022) <= a;
    layer1_outputs(4023) <= a or b;
    layer1_outputs(4024) <= not (a or b);
    layer1_outputs(4025) <= '1';
    layer1_outputs(4026) <= '0';
    layer1_outputs(4027) <= a and not b;
    layer1_outputs(4028) <= b;
    layer1_outputs(4029) <= a or b;
    layer1_outputs(4030) <= b;
    layer1_outputs(4031) <= not b;
    layer1_outputs(4032) <= b;
    layer1_outputs(4033) <= a and b;
    layer1_outputs(4034) <= not (a and b);
    layer1_outputs(4035) <= not a;
    layer1_outputs(4036) <= not a;
    layer1_outputs(4037) <= a and not b;
    layer1_outputs(4038) <= a and b;
    layer1_outputs(4039) <= not a;
    layer1_outputs(4040) <= '0';
    layer1_outputs(4041) <= b and not a;
    layer1_outputs(4042) <= '0';
    layer1_outputs(4043) <= not a or b;
    layer1_outputs(4044) <= b and not a;
    layer1_outputs(4045) <= a and b;
    layer1_outputs(4046) <= a and not b;
    layer1_outputs(4047) <= not a or b;
    layer1_outputs(4048) <= not (a and b);
    layer1_outputs(4049) <= '0';
    layer1_outputs(4050) <= not b or a;
    layer1_outputs(4051) <= not (a or b);
    layer1_outputs(4052) <= not (a and b);
    layer1_outputs(4053) <= b and not a;
    layer1_outputs(4054) <= '1';
    layer1_outputs(4055) <= '1';
    layer1_outputs(4056) <= not a or b;
    layer1_outputs(4057) <= a;
    layer1_outputs(4058) <= b and not a;
    layer1_outputs(4059) <= a or b;
    layer1_outputs(4060) <= '0';
    layer1_outputs(4061) <= a or b;
    layer1_outputs(4062) <= b and not a;
    layer1_outputs(4063) <= b;
    layer1_outputs(4064) <= b and not a;
    layer1_outputs(4065) <= a and not b;
    layer1_outputs(4066) <= not (a or b);
    layer1_outputs(4067) <= '1';
    layer1_outputs(4068) <= not (a and b);
    layer1_outputs(4069) <= not b;
    layer1_outputs(4070) <= b;
    layer1_outputs(4071) <= not (a and b);
    layer1_outputs(4072) <= not (a and b);
    layer1_outputs(4073) <= b;
    layer1_outputs(4074) <= b;
    layer1_outputs(4075) <= b and not a;
    layer1_outputs(4076) <= a;
    layer1_outputs(4077) <= '1';
    layer1_outputs(4078) <= b;
    layer1_outputs(4079) <= a or b;
    layer1_outputs(4080) <= not b or a;
    layer1_outputs(4081) <= '1';
    layer1_outputs(4082) <= a or b;
    layer1_outputs(4083) <= b and not a;
    layer1_outputs(4084) <= b and not a;
    layer1_outputs(4085) <= not b or a;
    layer1_outputs(4086) <= not (a and b);
    layer1_outputs(4087) <= not a or b;
    layer1_outputs(4088) <= a xor b;
    layer1_outputs(4089) <= '1';
    layer1_outputs(4090) <= '0';
    layer1_outputs(4091) <= '1';
    layer1_outputs(4092) <= a or b;
    layer1_outputs(4093) <= a xor b;
    layer1_outputs(4094) <= b and not a;
    layer1_outputs(4095) <= a and not b;
    layer1_outputs(4096) <= not b or a;
    layer1_outputs(4097) <= '1';
    layer1_outputs(4098) <= '0';
    layer1_outputs(4099) <= b;
    layer1_outputs(4100) <= not b or a;
    layer1_outputs(4101) <= a and not b;
    layer1_outputs(4102) <= not (a and b);
    layer1_outputs(4103) <= a;
    layer1_outputs(4104) <= not b;
    layer1_outputs(4105) <= '0';
    layer1_outputs(4106) <= a xor b;
    layer1_outputs(4107) <= not a;
    layer1_outputs(4108) <= not (a or b);
    layer1_outputs(4109) <= not a or b;
    layer1_outputs(4110) <= not (a and b);
    layer1_outputs(4111) <= not b;
    layer1_outputs(4112) <= not b;
    layer1_outputs(4113) <= a or b;
    layer1_outputs(4114) <= a xor b;
    layer1_outputs(4115) <= not (a or b);
    layer1_outputs(4116) <= b and not a;
    layer1_outputs(4117) <= a or b;
    layer1_outputs(4118) <= not a;
    layer1_outputs(4119) <= not (a and b);
    layer1_outputs(4120) <= not (a and b);
    layer1_outputs(4121) <= not b or a;
    layer1_outputs(4122) <= '1';
    layer1_outputs(4123) <= not b or a;
    layer1_outputs(4124) <= not b or a;
    layer1_outputs(4125) <= not b;
    layer1_outputs(4126) <= a or b;
    layer1_outputs(4127) <= a or b;
    layer1_outputs(4128) <= a and not b;
    layer1_outputs(4129) <= a and not b;
    layer1_outputs(4130) <= not (a or b);
    layer1_outputs(4131) <= a xor b;
    layer1_outputs(4132) <= a and b;
    layer1_outputs(4133) <= '1';
    layer1_outputs(4134) <= a xor b;
    layer1_outputs(4135) <= a or b;
    layer1_outputs(4136) <= '0';
    layer1_outputs(4137) <= a or b;
    layer1_outputs(4138) <= not b;
    layer1_outputs(4139) <= not b;
    layer1_outputs(4140) <= not a or b;
    layer1_outputs(4141) <= b and not a;
    layer1_outputs(4142) <= not a or b;
    layer1_outputs(4143) <= a and b;
    layer1_outputs(4144) <= '1';
    layer1_outputs(4145) <= '1';
    layer1_outputs(4146) <= '0';
    layer1_outputs(4147) <= b and not a;
    layer1_outputs(4148) <= not (a or b);
    layer1_outputs(4149) <= '1';
    layer1_outputs(4150) <= '0';
    layer1_outputs(4151) <= not (a and b);
    layer1_outputs(4152) <= a or b;
    layer1_outputs(4153) <= not a;
    layer1_outputs(4154) <= not a;
    layer1_outputs(4155) <= a;
    layer1_outputs(4156) <= not a or b;
    layer1_outputs(4157) <= not b;
    layer1_outputs(4158) <= b;
    layer1_outputs(4159) <= b and not a;
    layer1_outputs(4160) <= not (a and b);
    layer1_outputs(4161) <= a and b;
    layer1_outputs(4162) <= not a;
    layer1_outputs(4163) <= '0';
    layer1_outputs(4164) <= a and not b;
    layer1_outputs(4165) <= not b;
    layer1_outputs(4166) <= b;
    layer1_outputs(4167) <= b and not a;
    layer1_outputs(4168) <= not (a xor b);
    layer1_outputs(4169) <= '0';
    layer1_outputs(4170) <= '0';
    layer1_outputs(4171) <= not b or a;
    layer1_outputs(4172) <= not b;
    layer1_outputs(4173) <= not a or b;
    layer1_outputs(4174) <= not (a and b);
    layer1_outputs(4175) <= not a;
    layer1_outputs(4176) <= not b;
    layer1_outputs(4177) <= not (a or b);
    layer1_outputs(4178) <= not b or a;
    layer1_outputs(4179) <= a or b;
    layer1_outputs(4180) <= not (a and b);
    layer1_outputs(4181) <= a or b;
    layer1_outputs(4182) <= not a;
    layer1_outputs(4183) <= a and not b;
    layer1_outputs(4184) <= not b or a;
    layer1_outputs(4185) <= a and not b;
    layer1_outputs(4186) <= not (a or b);
    layer1_outputs(4187) <= '1';
    layer1_outputs(4188) <= '1';
    layer1_outputs(4189) <= a xor b;
    layer1_outputs(4190) <= not (a and b);
    layer1_outputs(4191) <= '1';
    layer1_outputs(4192) <= not a;
    layer1_outputs(4193) <= '0';
    layer1_outputs(4194) <= b and not a;
    layer1_outputs(4195) <= not (a or b);
    layer1_outputs(4196) <= a or b;
    layer1_outputs(4197) <= a xor b;
    layer1_outputs(4198) <= not b;
    layer1_outputs(4199) <= not a or b;
    layer1_outputs(4200) <= a or b;
    layer1_outputs(4201) <= not (a and b);
    layer1_outputs(4202) <= not b or a;
    layer1_outputs(4203) <= a xor b;
    layer1_outputs(4204) <= b and not a;
    layer1_outputs(4205) <= a or b;
    layer1_outputs(4206) <= a and b;
    layer1_outputs(4207) <= not b;
    layer1_outputs(4208) <= not b;
    layer1_outputs(4209) <= a and not b;
    layer1_outputs(4210) <= b;
    layer1_outputs(4211) <= a;
    layer1_outputs(4212) <= not a or b;
    layer1_outputs(4213) <= '0';
    layer1_outputs(4214) <= a or b;
    layer1_outputs(4215) <= not (a and b);
    layer1_outputs(4216) <= not (a and b);
    layer1_outputs(4217) <= not (a and b);
    layer1_outputs(4218) <= b and not a;
    layer1_outputs(4219) <= a and not b;
    layer1_outputs(4220) <= b and not a;
    layer1_outputs(4221) <= not a or b;
    layer1_outputs(4222) <= a and b;
    layer1_outputs(4223) <= not (a or b);
    layer1_outputs(4224) <= '1';
    layer1_outputs(4225) <= not b;
    layer1_outputs(4226) <= a;
    layer1_outputs(4227) <= a;
    layer1_outputs(4228) <= not b;
    layer1_outputs(4229) <= '1';
    layer1_outputs(4230) <= not b or a;
    layer1_outputs(4231) <= a and not b;
    layer1_outputs(4232) <= not (a and b);
    layer1_outputs(4233) <= '0';
    layer1_outputs(4234) <= not b or a;
    layer1_outputs(4235) <= b and not a;
    layer1_outputs(4236) <= a and b;
    layer1_outputs(4237) <= a and not b;
    layer1_outputs(4238) <= not (a xor b);
    layer1_outputs(4239) <= not (a xor b);
    layer1_outputs(4240) <= '0';
    layer1_outputs(4241) <= '1';
    layer1_outputs(4242) <= not a;
    layer1_outputs(4243) <= not a or b;
    layer1_outputs(4244) <= b;
    layer1_outputs(4245) <= a;
    layer1_outputs(4246) <= a xor b;
    layer1_outputs(4247) <= not (a and b);
    layer1_outputs(4248) <= not b;
    layer1_outputs(4249) <= not a;
    layer1_outputs(4250) <= '0';
    layer1_outputs(4251) <= b;
    layer1_outputs(4252) <= '0';
    layer1_outputs(4253) <= a;
    layer1_outputs(4254) <= a and not b;
    layer1_outputs(4255) <= not (a and b);
    layer1_outputs(4256) <= not (a and b);
    layer1_outputs(4257) <= a or b;
    layer1_outputs(4258) <= a;
    layer1_outputs(4259) <= b;
    layer1_outputs(4260) <= '0';
    layer1_outputs(4261) <= a and b;
    layer1_outputs(4262) <= not b or a;
    layer1_outputs(4263) <= a or b;
    layer1_outputs(4264) <= a and not b;
    layer1_outputs(4265) <= '1';
    layer1_outputs(4266) <= a;
    layer1_outputs(4267) <= not b;
    layer1_outputs(4268) <= not (a or b);
    layer1_outputs(4269) <= '1';
    layer1_outputs(4270) <= not b;
    layer1_outputs(4271) <= not (a and b);
    layer1_outputs(4272) <= a and b;
    layer1_outputs(4273) <= b and not a;
    layer1_outputs(4274) <= b;
    layer1_outputs(4275) <= not b or a;
    layer1_outputs(4276) <= a or b;
    layer1_outputs(4277) <= not (a or b);
    layer1_outputs(4278) <= b and not a;
    layer1_outputs(4279) <= a and b;
    layer1_outputs(4280) <= '1';
    layer1_outputs(4281) <= a;
    layer1_outputs(4282) <= not a;
    layer1_outputs(4283) <= a xor b;
    layer1_outputs(4284) <= '0';
    layer1_outputs(4285) <= not a;
    layer1_outputs(4286) <= b;
    layer1_outputs(4287) <= a and b;
    layer1_outputs(4288) <= not a;
    layer1_outputs(4289) <= '1';
    layer1_outputs(4290) <= b;
    layer1_outputs(4291) <= a and not b;
    layer1_outputs(4292) <= not (a xor b);
    layer1_outputs(4293) <= a or b;
    layer1_outputs(4294) <= not a or b;
    layer1_outputs(4295) <= a and b;
    layer1_outputs(4296) <= not (a xor b);
    layer1_outputs(4297) <= a and not b;
    layer1_outputs(4298) <= b;
    layer1_outputs(4299) <= not a or b;
    layer1_outputs(4300) <= b and not a;
    layer1_outputs(4301) <= '1';
    layer1_outputs(4302) <= a;
    layer1_outputs(4303) <= a;
    layer1_outputs(4304) <= b and not a;
    layer1_outputs(4305) <= a or b;
    layer1_outputs(4306) <= not (a or b);
    layer1_outputs(4307) <= a;
    layer1_outputs(4308) <= b;
    layer1_outputs(4309) <= b;
    layer1_outputs(4310) <= not b or a;
    layer1_outputs(4311) <= b and not a;
    layer1_outputs(4312) <= '0';
    layer1_outputs(4313) <= not a or b;
    layer1_outputs(4314) <= not b;
    layer1_outputs(4315) <= a and not b;
    layer1_outputs(4316) <= not (a or b);
    layer1_outputs(4317) <= not a;
    layer1_outputs(4318) <= a and b;
    layer1_outputs(4319) <= a and b;
    layer1_outputs(4320) <= b and not a;
    layer1_outputs(4321) <= not b;
    layer1_outputs(4322) <= not (a and b);
    layer1_outputs(4323) <= a and b;
    layer1_outputs(4324) <= not a or b;
    layer1_outputs(4325) <= not b or a;
    layer1_outputs(4326) <= '1';
    layer1_outputs(4327) <= a;
    layer1_outputs(4328) <= a or b;
    layer1_outputs(4329) <= b;
    layer1_outputs(4330) <= b;
    layer1_outputs(4331) <= '0';
    layer1_outputs(4332) <= a or b;
    layer1_outputs(4333) <= a or b;
    layer1_outputs(4334) <= a xor b;
    layer1_outputs(4335) <= not (a or b);
    layer1_outputs(4336) <= b;
    layer1_outputs(4337) <= not a or b;
    layer1_outputs(4338) <= not a;
    layer1_outputs(4339) <= not (a and b);
    layer1_outputs(4340) <= '1';
    layer1_outputs(4341) <= b and not a;
    layer1_outputs(4342) <= not (a or b);
    layer1_outputs(4343) <= a xor b;
    layer1_outputs(4344) <= a or b;
    layer1_outputs(4345) <= not (a xor b);
    layer1_outputs(4346) <= not (a xor b);
    layer1_outputs(4347) <= not (a or b);
    layer1_outputs(4348) <= not (a and b);
    layer1_outputs(4349) <= not b;
    layer1_outputs(4350) <= a and b;
    layer1_outputs(4351) <= not a;
    layer1_outputs(4352) <= not a;
    layer1_outputs(4353) <= not b or a;
    layer1_outputs(4354) <= '0';
    layer1_outputs(4355) <= b and not a;
    layer1_outputs(4356) <= not (a and b);
    layer1_outputs(4357) <= b and not a;
    layer1_outputs(4358) <= a or b;
    layer1_outputs(4359) <= b;
    layer1_outputs(4360) <= not (a xor b);
    layer1_outputs(4361) <= a;
    layer1_outputs(4362) <= not (a or b);
    layer1_outputs(4363) <= not b or a;
    layer1_outputs(4364) <= a and not b;
    layer1_outputs(4365) <= '0';
    layer1_outputs(4366) <= not (a or b);
    layer1_outputs(4367) <= not a or b;
    layer1_outputs(4368) <= not (a and b);
    layer1_outputs(4369) <= a and not b;
    layer1_outputs(4370) <= not (a or b);
    layer1_outputs(4371) <= b;
    layer1_outputs(4372) <= '0';
    layer1_outputs(4373) <= not b or a;
    layer1_outputs(4374) <= not b;
    layer1_outputs(4375) <= a;
    layer1_outputs(4376) <= not b or a;
    layer1_outputs(4377) <= '0';
    layer1_outputs(4378) <= not a;
    layer1_outputs(4379) <= '1';
    layer1_outputs(4380) <= not (a xor b);
    layer1_outputs(4381) <= '1';
    layer1_outputs(4382) <= not (a xor b);
    layer1_outputs(4383) <= '0';
    layer1_outputs(4384) <= not (a and b);
    layer1_outputs(4385) <= a;
    layer1_outputs(4386) <= not (a or b);
    layer1_outputs(4387) <= b and not a;
    layer1_outputs(4388) <= b and not a;
    layer1_outputs(4389) <= not a;
    layer1_outputs(4390) <= a and b;
    layer1_outputs(4391) <= a or b;
    layer1_outputs(4392) <= not a;
    layer1_outputs(4393) <= a and not b;
    layer1_outputs(4394) <= b and not a;
    layer1_outputs(4395) <= a and not b;
    layer1_outputs(4396) <= '0';
    layer1_outputs(4397) <= '0';
    layer1_outputs(4398) <= '1';
    layer1_outputs(4399) <= not (a or b);
    layer1_outputs(4400) <= b;
    layer1_outputs(4401) <= not a;
    layer1_outputs(4402) <= a;
    layer1_outputs(4403) <= not b or a;
    layer1_outputs(4404) <= not a or b;
    layer1_outputs(4405) <= a or b;
    layer1_outputs(4406) <= not (a xor b);
    layer1_outputs(4407) <= a;
    layer1_outputs(4408) <= not (a and b);
    layer1_outputs(4409) <= not b or a;
    layer1_outputs(4410) <= not a or b;
    layer1_outputs(4411) <= a or b;
    layer1_outputs(4412) <= not (a or b);
    layer1_outputs(4413) <= not (a and b);
    layer1_outputs(4414) <= a or b;
    layer1_outputs(4415) <= not b;
    layer1_outputs(4416) <= '1';
    layer1_outputs(4417) <= a or b;
    layer1_outputs(4418) <= not (a xor b);
    layer1_outputs(4419) <= not a;
    layer1_outputs(4420) <= not b;
    layer1_outputs(4421) <= a or b;
    layer1_outputs(4422) <= not (a and b);
    layer1_outputs(4423) <= not a or b;
    layer1_outputs(4424) <= not (a and b);
    layer1_outputs(4425) <= b;
    layer1_outputs(4426) <= '1';
    layer1_outputs(4427) <= b and not a;
    layer1_outputs(4428) <= b and not a;
    layer1_outputs(4429) <= not (a or b);
    layer1_outputs(4430) <= not b or a;
    layer1_outputs(4431) <= a;
    layer1_outputs(4432) <= not b or a;
    layer1_outputs(4433) <= not a;
    layer1_outputs(4434) <= not (a and b);
    layer1_outputs(4435) <= '1';
    layer1_outputs(4436) <= a or b;
    layer1_outputs(4437) <= not b;
    layer1_outputs(4438) <= not a;
    layer1_outputs(4439) <= not a or b;
    layer1_outputs(4440) <= '0';
    layer1_outputs(4441) <= not a or b;
    layer1_outputs(4442) <= not (a or b);
    layer1_outputs(4443) <= '0';
    layer1_outputs(4444) <= a and b;
    layer1_outputs(4445) <= b and not a;
    layer1_outputs(4446) <= b;
    layer1_outputs(4447) <= a or b;
    layer1_outputs(4448) <= not a or b;
    layer1_outputs(4449) <= not a or b;
    layer1_outputs(4450) <= a xor b;
    layer1_outputs(4451) <= a and b;
    layer1_outputs(4452) <= a;
    layer1_outputs(4453) <= b;
    layer1_outputs(4454) <= a and b;
    layer1_outputs(4455) <= b;
    layer1_outputs(4456) <= not (a or b);
    layer1_outputs(4457) <= a xor b;
    layer1_outputs(4458) <= a and not b;
    layer1_outputs(4459) <= a and b;
    layer1_outputs(4460) <= a;
    layer1_outputs(4461) <= b;
    layer1_outputs(4462) <= '1';
    layer1_outputs(4463) <= not (a and b);
    layer1_outputs(4464) <= not a or b;
    layer1_outputs(4465) <= a and b;
    layer1_outputs(4466) <= not a or b;
    layer1_outputs(4467) <= a;
    layer1_outputs(4468) <= not b or a;
    layer1_outputs(4469) <= '1';
    layer1_outputs(4470) <= not a or b;
    layer1_outputs(4471) <= '0';
    layer1_outputs(4472) <= '1';
    layer1_outputs(4473) <= a or b;
    layer1_outputs(4474) <= '1';
    layer1_outputs(4475) <= a and b;
    layer1_outputs(4476) <= not (a and b);
    layer1_outputs(4477) <= not (a or b);
    layer1_outputs(4478) <= not (a xor b);
    layer1_outputs(4479) <= not (a or b);
    layer1_outputs(4480) <= a xor b;
    layer1_outputs(4481) <= not a or b;
    layer1_outputs(4482) <= b and not a;
    layer1_outputs(4483) <= a or b;
    layer1_outputs(4484) <= not b or a;
    layer1_outputs(4485) <= not (a or b);
    layer1_outputs(4486) <= not a;
    layer1_outputs(4487) <= b and not a;
    layer1_outputs(4488) <= not (a xor b);
    layer1_outputs(4489) <= not a;
    layer1_outputs(4490) <= '0';
    layer1_outputs(4491) <= a and b;
    layer1_outputs(4492) <= '1';
    layer1_outputs(4493) <= '1';
    layer1_outputs(4494) <= a and not b;
    layer1_outputs(4495) <= not a;
    layer1_outputs(4496) <= not (a xor b);
    layer1_outputs(4497) <= a;
    layer1_outputs(4498) <= not (a or b);
    layer1_outputs(4499) <= a xor b;
    layer1_outputs(4500) <= '0';
    layer1_outputs(4501) <= not a or b;
    layer1_outputs(4502) <= not (a or b);
    layer1_outputs(4503) <= not b;
    layer1_outputs(4504) <= not a;
    layer1_outputs(4505) <= not b;
    layer1_outputs(4506) <= not b or a;
    layer1_outputs(4507) <= not b or a;
    layer1_outputs(4508) <= not b or a;
    layer1_outputs(4509) <= not b;
    layer1_outputs(4510) <= b and not a;
    layer1_outputs(4511) <= '1';
    layer1_outputs(4512) <= a and not b;
    layer1_outputs(4513) <= not b;
    layer1_outputs(4514) <= b;
    layer1_outputs(4515) <= not b;
    layer1_outputs(4516) <= not a or b;
    layer1_outputs(4517) <= a and b;
    layer1_outputs(4518) <= not a or b;
    layer1_outputs(4519) <= a;
    layer1_outputs(4520) <= a xor b;
    layer1_outputs(4521) <= b;
    layer1_outputs(4522) <= not b or a;
    layer1_outputs(4523) <= not a;
    layer1_outputs(4524) <= a xor b;
    layer1_outputs(4525) <= a and not b;
    layer1_outputs(4526) <= not a or b;
    layer1_outputs(4527) <= b and not a;
    layer1_outputs(4528) <= a xor b;
    layer1_outputs(4529) <= not b;
    layer1_outputs(4530) <= not b or a;
    layer1_outputs(4531) <= a and b;
    layer1_outputs(4532) <= a xor b;
    layer1_outputs(4533) <= not (a or b);
    layer1_outputs(4534) <= not (a or b);
    layer1_outputs(4535) <= a and b;
    layer1_outputs(4536) <= '1';
    layer1_outputs(4537) <= a xor b;
    layer1_outputs(4538) <= a and not b;
    layer1_outputs(4539) <= not b;
    layer1_outputs(4540) <= not (a and b);
    layer1_outputs(4541) <= b and not a;
    layer1_outputs(4542) <= '1';
    layer1_outputs(4543) <= '0';
    layer1_outputs(4544) <= not (a and b);
    layer1_outputs(4545) <= b and not a;
    layer1_outputs(4546) <= '1';
    layer1_outputs(4547) <= b and not a;
    layer1_outputs(4548) <= '0';
    layer1_outputs(4549) <= a or b;
    layer1_outputs(4550) <= b;
    layer1_outputs(4551) <= not a;
    layer1_outputs(4552) <= not (a or b);
    layer1_outputs(4553) <= not (a and b);
    layer1_outputs(4554) <= a;
    layer1_outputs(4555) <= a and not b;
    layer1_outputs(4556) <= '0';
    layer1_outputs(4557) <= not (a or b);
    layer1_outputs(4558) <= '1';
    layer1_outputs(4559) <= b and not a;
    layer1_outputs(4560) <= not a;
    layer1_outputs(4561) <= a or b;
    layer1_outputs(4562) <= not b or a;
    layer1_outputs(4563) <= a;
    layer1_outputs(4564) <= a and not b;
    layer1_outputs(4565) <= a xor b;
    layer1_outputs(4566) <= not (a and b);
    layer1_outputs(4567) <= not a or b;
    layer1_outputs(4568) <= '1';
    layer1_outputs(4569) <= b and not a;
    layer1_outputs(4570) <= '0';
    layer1_outputs(4571) <= not b;
    layer1_outputs(4572) <= not (a and b);
    layer1_outputs(4573) <= a or b;
    layer1_outputs(4574) <= not b or a;
    layer1_outputs(4575) <= not (a and b);
    layer1_outputs(4576) <= not (a and b);
    layer1_outputs(4577) <= '1';
    layer1_outputs(4578) <= a and not b;
    layer1_outputs(4579) <= b and not a;
    layer1_outputs(4580) <= not b;
    layer1_outputs(4581) <= not (a and b);
    layer1_outputs(4582) <= not a or b;
    layer1_outputs(4583) <= not (a xor b);
    layer1_outputs(4584) <= not (a or b);
    layer1_outputs(4585) <= not (a xor b);
    layer1_outputs(4586) <= '0';
    layer1_outputs(4587) <= a and not b;
    layer1_outputs(4588) <= not (a and b);
    layer1_outputs(4589) <= not a;
    layer1_outputs(4590) <= a or b;
    layer1_outputs(4591) <= not (a xor b);
    layer1_outputs(4592) <= not (a or b);
    layer1_outputs(4593) <= '1';
    layer1_outputs(4594) <= a and not b;
    layer1_outputs(4595) <= a;
    layer1_outputs(4596) <= '0';
    layer1_outputs(4597) <= '1';
    layer1_outputs(4598) <= not a;
    layer1_outputs(4599) <= a;
    layer1_outputs(4600) <= not a;
    layer1_outputs(4601) <= '1';
    layer1_outputs(4602) <= not (a or b);
    layer1_outputs(4603) <= a xor b;
    layer1_outputs(4604) <= '0';
    layer1_outputs(4605) <= not a;
    layer1_outputs(4606) <= '1';
    layer1_outputs(4607) <= b and not a;
    layer1_outputs(4608) <= not b or a;
    layer1_outputs(4609) <= b and not a;
    layer1_outputs(4610) <= not (a and b);
    layer1_outputs(4611) <= b and not a;
    layer1_outputs(4612) <= not (a or b);
    layer1_outputs(4613) <= '1';
    layer1_outputs(4614) <= b and not a;
    layer1_outputs(4615) <= a or b;
    layer1_outputs(4616) <= b and not a;
    layer1_outputs(4617) <= a xor b;
    layer1_outputs(4618) <= not b;
    layer1_outputs(4619) <= a and not b;
    layer1_outputs(4620) <= '0';
    layer1_outputs(4621) <= a and b;
    layer1_outputs(4622) <= '0';
    layer1_outputs(4623) <= not (a or b);
    layer1_outputs(4624) <= b;
    layer1_outputs(4625) <= not (a xor b);
    layer1_outputs(4626) <= not (a or b);
    layer1_outputs(4627) <= not (a or b);
    layer1_outputs(4628) <= not b or a;
    layer1_outputs(4629) <= a or b;
    layer1_outputs(4630) <= not (a or b);
    layer1_outputs(4631) <= a and not b;
    layer1_outputs(4632) <= '0';
    layer1_outputs(4633) <= '0';
    layer1_outputs(4634) <= not b or a;
    layer1_outputs(4635) <= not b;
    layer1_outputs(4636) <= b;
    layer1_outputs(4637) <= a xor b;
    layer1_outputs(4638) <= '0';
    layer1_outputs(4639) <= '0';
    layer1_outputs(4640) <= not (a and b);
    layer1_outputs(4641) <= a or b;
    layer1_outputs(4642) <= a and not b;
    layer1_outputs(4643) <= a and not b;
    layer1_outputs(4644) <= not b;
    layer1_outputs(4645) <= a or b;
    layer1_outputs(4646) <= not a;
    layer1_outputs(4647) <= a;
    layer1_outputs(4648) <= '0';
    layer1_outputs(4649) <= not (a and b);
    layer1_outputs(4650) <= a;
    layer1_outputs(4651) <= b and not a;
    layer1_outputs(4652) <= b;
    layer1_outputs(4653) <= a xor b;
    layer1_outputs(4654) <= '1';
    layer1_outputs(4655) <= '0';
    layer1_outputs(4656) <= a and b;
    layer1_outputs(4657) <= a or b;
    layer1_outputs(4658) <= not (a xor b);
    layer1_outputs(4659) <= b and not a;
    layer1_outputs(4660) <= a and b;
    layer1_outputs(4661) <= not (a and b);
    layer1_outputs(4662) <= not a;
    layer1_outputs(4663) <= a;
    layer1_outputs(4664) <= a or b;
    layer1_outputs(4665) <= not (a and b);
    layer1_outputs(4666) <= a or b;
    layer1_outputs(4667) <= not a or b;
    layer1_outputs(4668) <= not (a and b);
    layer1_outputs(4669) <= '1';
    layer1_outputs(4670) <= not a;
    layer1_outputs(4671) <= not b;
    layer1_outputs(4672) <= not a or b;
    layer1_outputs(4673) <= '0';
    layer1_outputs(4674) <= a;
    layer1_outputs(4675) <= not b or a;
    layer1_outputs(4676) <= not (a or b);
    layer1_outputs(4677) <= a;
    layer1_outputs(4678) <= not a or b;
    layer1_outputs(4679) <= not a or b;
    layer1_outputs(4680) <= b and not a;
    layer1_outputs(4681) <= not a or b;
    layer1_outputs(4682) <= not (a and b);
    layer1_outputs(4683) <= not b or a;
    layer1_outputs(4684) <= not (a and b);
    layer1_outputs(4685) <= not b;
    layer1_outputs(4686) <= a;
    layer1_outputs(4687) <= a;
    layer1_outputs(4688) <= '0';
    layer1_outputs(4689) <= not a;
    layer1_outputs(4690) <= not (a or b);
    layer1_outputs(4691) <= a;
    layer1_outputs(4692) <= a xor b;
    layer1_outputs(4693) <= not b;
    layer1_outputs(4694) <= b and not a;
    layer1_outputs(4695) <= not (a xor b);
    layer1_outputs(4696) <= b and not a;
    layer1_outputs(4697) <= '1';
    layer1_outputs(4698) <= not (a and b);
    layer1_outputs(4699) <= a;
    layer1_outputs(4700) <= '0';
    layer1_outputs(4701) <= b and not a;
    layer1_outputs(4702) <= not b or a;
    layer1_outputs(4703) <= not (a xor b);
    layer1_outputs(4704) <= '0';
    layer1_outputs(4705) <= a or b;
    layer1_outputs(4706) <= a and b;
    layer1_outputs(4707) <= '0';
    layer1_outputs(4708) <= not b or a;
    layer1_outputs(4709) <= '0';
    layer1_outputs(4710) <= a;
    layer1_outputs(4711) <= not (a or b);
    layer1_outputs(4712) <= not (a xor b);
    layer1_outputs(4713) <= a and not b;
    layer1_outputs(4714) <= a and not b;
    layer1_outputs(4715) <= not b;
    layer1_outputs(4716) <= a and not b;
    layer1_outputs(4717) <= a or b;
    layer1_outputs(4718) <= a and b;
    layer1_outputs(4719) <= b and not a;
    layer1_outputs(4720) <= '1';
    layer1_outputs(4721) <= not (a or b);
    layer1_outputs(4722) <= not b;
    layer1_outputs(4723) <= b and not a;
    layer1_outputs(4724) <= not (a xor b);
    layer1_outputs(4725) <= b and not a;
    layer1_outputs(4726) <= '1';
    layer1_outputs(4727) <= '1';
    layer1_outputs(4728) <= not b or a;
    layer1_outputs(4729) <= a and b;
    layer1_outputs(4730) <= not (a xor b);
    layer1_outputs(4731) <= '1';
    layer1_outputs(4732) <= not b;
    layer1_outputs(4733) <= not a or b;
    layer1_outputs(4734) <= a;
    layer1_outputs(4735) <= b and not a;
    layer1_outputs(4736) <= not b;
    layer1_outputs(4737) <= a;
    layer1_outputs(4738) <= b and not a;
    layer1_outputs(4739) <= '1';
    layer1_outputs(4740) <= not (a and b);
    layer1_outputs(4741) <= a or b;
    layer1_outputs(4742) <= '1';
    layer1_outputs(4743) <= b;
    layer1_outputs(4744) <= a or b;
    layer1_outputs(4745) <= '0';
    layer1_outputs(4746) <= a or b;
    layer1_outputs(4747) <= not b or a;
    layer1_outputs(4748) <= not a or b;
    layer1_outputs(4749) <= '0';
    layer1_outputs(4750) <= b and not a;
    layer1_outputs(4751) <= b and not a;
    layer1_outputs(4752) <= a and b;
    layer1_outputs(4753) <= b and not a;
    layer1_outputs(4754) <= a and b;
    layer1_outputs(4755) <= not (a and b);
    layer1_outputs(4756) <= not (a or b);
    layer1_outputs(4757) <= '0';
    layer1_outputs(4758) <= not a or b;
    layer1_outputs(4759) <= a and not b;
    layer1_outputs(4760) <= not b or a;
    layer1_outputs(4761) <= '1';
    layer1_outputs(4762) <= '1';
    layer1_outputs(4763) <= not (a or b);
    layer1_outputs(4764) <= not (a and b);
    layer1_outputs(4765) <= not a or b;
    layer1_outputs(4766) <= '1';
    layer1_outputs(4767) <= not (a or b);
    layer1_outputs(4768) <= a or b;
    layer1_outputs(4769) <= a and not b;
    layer1_outputs(4770) <= a or b;
    layer1_outputs(4771) <= '1';
    layer1_outputs(4772) <= a or b;
    layer1_outputs(4773) <= a or b;
    layer1_outputs(4774) <= a;
    layer1_outputs(4775) <= a;
    layer1_outputs(4776) <= b and not a;
    layer1_outputs(4777) <= not (a and b);
    layer1_outputs(4778) <= a and not b;
    layer1_outputs(4779) <= '0';
    layer1_outputs(4780) <= '0';
    layer1_outputs(4781) <= a;
    layer1_outputs(4782) <= not b;
    layer1_outputs(4783) <= not (a and b);
    layer1_outputs(4784) <= '0';
    layer1_outputs(4785) <= a and not b;
    layer1_outputs(4786) <= a;
    layer1_outputs(4787) <= a;
    layer1_outputs(4788) <= not a or b;
    layer1_outputs(4789) <= '0';
    layer1_outputs(4790) <= a;
    layer1_outputs(4791) <= b and not a;
    layer1_outputs(4792) <= not b;
    layer1_outputs(4793) <= a and b;
    layer1_outputs(4794) <= not a or b;
    layer1_outputs(4795) <= a and not b;
    layer1_outputs(4796) <= '1';
    layer1_outputs(4797) <= not (a or b);
    layer1_outputs(4798) <= '1';
    layer1_outputs(4799) <= a;
    layer1_outputs(4800) <= b and not a;
    layer1_outputs(4801) <= a or b;
    layer1_outputs(4802) <= b;
    layer1_outputs(4803) <= '0';
    layer1_outputs(4804) <= not (a xor b);
    layer1_outputs(4805) <= a and not b;
    layer1_outputs(4806) <= a and b;
    layer1_outputs(4807) <= a;
    layer1_outputs(4808) <= a;
    layer1_outputs(4809) <= '0';
    layer1_outputs(4810) <= '0';
    layer1_outputs(4811) <= a and not b;
    layer1_outputs(4812) <= a;
    layer1_outputs(4813) <= a and b;
    layer1_outputs(4814) <= not b or a;
    layer1_outputs(4815) <= not b or a;
    layer1_outputs(4816) <= a or b;
    layer1_outputs(4817) <= b;
    layer1_outputs(4818) <= a xor b;
    layer1_outputs(4819) <= not a or b;
    layer1_outputs(4820) <= not b or a;
    layer1_outputs(4821) <= not a;
    layer1_outputs(4822) <= '0';
    layer1_outputs(4823) <= '1';
    layer1_outputs(4824) <= '0';
    layer1_outputs(4825) <= '1';
    layer1_outputs(4826) <= a and not b;
    layer1_outputs(4827) <= b and not a;
    layer1_outputs(4828) <= a and not b;
    layer1_outputs(4829) <= not (a and b);
    layer1_outputs(4830) <= a and b;
    layer1_outputs(4831) <= '1';
    layer1_outputs(4832) <= not a;
    layer1_outputs(4833) <= not a or b;
    layer1_outputs(4834) <= a;
    layer1_outputs(4835) <= b;
    layer1_outputs(4836) <= a;
    layer1_outputs(4837) <= not (a and b);
    layer1_outputs(4838) <= b and not a;
    layer1_outputs(4839) <= not (a and b);
    layer1_outputs(4840) <= '0';
    layer1_outputs(4841) <= not a or b;
    layer1_outputs(4842) <= not a;
    layer1_outputs(4843) <= a and b;
    layer1_outputs(4844) <= a;
    layer1_outputs(4845) <= not (a or b);
    layer1_outputs(4846) <= not (a and b);
    layer1_outputs(4847) <= b and not a;
    layer1_outputs(4848) <= a and b;
    layer1_outputs(4849) <= not (a xor b);
    layer1_outputs(4850) <= not (a xor b);
    layer1_outputs(4851) <= a and not b;
    layer1_outputs(4852) <= '1';
    layer1_outputs(4853) <= a and b;
    layer1_outputs(4854) <= '1';
    layer1_outputs(4855) <= a and b;
    layer1_outputs(4856) <= not a or b;
    layer1_outputs(4857) <= a;
    layer1_outputs(4858) <= '1';
    layer1_outputs(4859) <= '0';
    layer1_outputs(4860) <= b;
    layer1_outputs(4861) <= not b or a;
    layer1_outputs(4862) <= '1';
    layer1_outputs(4863) <= a or b;
    layer1_outputs(4864) <= '0';
    layer1_outputs(4865) <= '1';
    layer1_outputs(4866) <= b and not a;
    layer1_outputs(4867) <= b and not a;
    layer1_outputs(4868) <= not b or a;
    layer1_outputs(4869) <= not (a or b);
    layer1_outputs(4870) <= b and not a;
    layer1_outputs(4871) <= not (a xor b);
    layer1_outputs(4872) <= not b or a;
    layer1_outputs(4873) <= not (a and b);
    layer1_outputs(4874) <= not a;
    layer1_outputs(4875) <= b and not a;
    layer1_outputs(4876) <= not b;
    layer1_outputs(4877) <= '1';
    layer1_outputs(4878) <= b;
    layer1_outputs(4879) <= '1';
    layer1_outputs(4880) <= a and b;
    layer1_outputs(4881) <= not b or a;
    layer1_outputs(4882) <= not a;
    layer1_outputs(4883) <= not (a or b);
    layer1_outputs(4884) <= not a;
    layer1_outputs(4885) <= not (a and b);
    layer1_outputs(4886) <= not b;
    layer1_outputs(4887) <= not (a and b);
    layer1_outputs(4888) <= a xor b;
    layer1_outputs(4889) <= not a or b;
    layer1_outputs(4890) <= a and not b;
    layer1_outputs(4891) <= a or b;
    layer1_outputs(4892) <= not b;
    layer1_outputs(4893) <= b;
    layer1_outputs(4894) <= a or b;
    layer1_outputs(4895) <= a and not b;
    layer1_outputs(4896) <= not (a or b);
    layer1_outputs(4897) <= a or b;
    layer1_outputs(4898) <= b;
    layer1_outputs(4899) <= '1';
    layer1_outputs(4900) <= not (a xor b);
    layer1_outputs(4901) <= not a;
    layer1_outputs(4902) <= a and b;
    layer1_outputs(4903) <= '0';
    layer1_outputs(4904) <= not b;
    layer1_outputs(4905) <= not a or b;
    layer1_outputs(4906) <= b;
    layer1_outputs(4907) <= not (a or b);
    layer1_outputs(4908) <= a;
    layer1_outputs(4909) <= a or b;
    layer1_outputs(4910) <= not b or a;
    layer1_outputs(4911) <= not (a or b);
    layer1_outputs(4912) <= not b or a;
    layer1_outputs(4913) <= '0';
    layer1_outputs(4914) <= not b or a;
    layer1_outputs(4915) <= not (a or b);
    layer1_outputs(4916) <= not b;
    layer1_outputs(4917) <= b and not a;
    layer1_outputs(4918) <= not a;
    layer1_outputs(4919) <= a and b;
    layer1_outputs(4920) <= a and b;
    layer1_outputs(4921) <= not a;
    layer1_outputs(4922) <= '1';
    layer1_outputs(4923) <= a xor b;
    layer1_outputs(4924) <= not b;
    layer1_outputs(4925) <= not b or a;
    layer1_outputs(4926) <= '0';
    layer1_outputs(4927) <= not (a and b);
    layer1_outputs(4928) <= not b or a;
    layer1_outputs(4929) <= '1';
    layer1_outputs(4930) <= a and not b;
    layer1_outputs(4931) <= '1';
    layer1_outputs(4932) <= not b or a;
    layer1_outputs(4933) <= b and not a;
    layer1_outputs(4934) <= not (a and b);
    layer1_outputs(4935) <= not b or a;
    layer1_outputs(4936) <= '0';
    layer1_outputs(4937) <= not a or b;
    layer1_outputs(4938) <= not b;
    layer1_outputs(4939) <= a and b;
    layer1_outputs(4940) <= a and b;
    layer1_outputs(4941) <= not b;
    layer1_outputs(4942) <= not (a or b);
    layer1_outputs(4943) <= not b or a;
    layer1_outputs(4944) <= not (a or b);
    layer1_outputs(4945) <= not a or b;
    layer1_outputs(4946) <= '1';
    layer1_outputs(4947) <= b;
    layer1_outputs(4948) <= not b or a;
    layer1_outputs(4949) <= not b;
    layer1_outputs(4950) <= not (a xor b);
    layer1_outputs(4951) <= not (a or b);
    layer1_outputs(4952) <= not a or b;
    layer1_outputs(4953) <= not a or b;
    layer1_outputs(4954) <= not a or b;
    layer1_outputs(4955) <= not a or b;
    layer1_outputs(4956) <= b and not a;
    layer1_outputs(4957) <= a;
    layer1_outputs(4958) <= b and not a;
    layer1_outputs(4959) <= a;
    layer1_outputs(4960) <= a or b;
    layer1_outputs(4961) <= '0';
    layer1_outputs(4962) <= '1';
    layer1_outputs(4963) <= a xor b;
    layer1_outputs(4964) <= not b or a;
    layer1_outputs(4965) <= not (a or b);
    layer1_outputs(4966) <= b and not a;
    layer1_outputs(4967) <= b and not a;
    layer1_outputs(4968) <= not a;
    layer1_outputs(4969) <= not (a and b);
    layer1_outputs(4970) <= not b or a;
    layer1_outputs(4971) <= b and not a;
    layer1_outputs(4972) <= b;
    layer1_outputs(4973) <= a and not b;
    layer1_outputs(4974) <= '0';
    layer1_outputs(4975) <= a xor b;
    layer1_outputs(4976) <= '1';
    layer1_outputs(4977) <= not b or a;
    layer1_outputs(4978) <= not (a and b);
    layer1_outputs(4979) <= a;
    layer1_outputs(4980) <= not (a and b);
    layer1_outputs(4981) <= '0';
    layer1_outputs(4982) <= a and not b;
    layer1_outputs(4983) <= not a;
    layer1_outputs(4984) <= '0';
    layer1_outputs(4985) <= '1';
    layer1_outputs(4986) <= a and not b;
    layer1_outputs(4987) <= not a or b;
    layer1_outputs(4988) <= not b;
    layer1_outputs(4989) <= b and not a;
    layer1_outputs(4990) <= not (a or b);
    layer1_outputs(4991) <= not b;
    layer1_outputs(4992) <= '1';
    layer1_outputs(4993) <= '0';
    layer1_outputs(4994) <= not b or a;
    layer1_outputs(4995) <= a or b;
    layer1_outputs(4996) <= a or b;
    layer1_outputs(4997) <= '0';
    layer1_outputs(4998) <= a;
    layer1_outputs(4999) <= not (a or b);
    layer1_outputs(5000) <= a or b;
    layer1_outputs(5001) <= b and not a;
    layer1_outputs(5002) <= not b;
    layer1_outputs(5003) <= a and b;
    layer1_outputs(5004) <= not b or a;
    layer1_outputs(5005) <= a and b;
    layer1_outputs(5006) <= '0';
    layer1_outputs(5007) <= not a;
    layer1_outputs(5008) <= '1';
    layer1_outputs(5009) <= a or b;
    layer1_outputs(5010) <= '1';
    layer1_outputs(5011) <= not (a or b);
    layer1_outputs(5012) <= not (a xor b);
    layer1_outputs(5013) <= b;
    layer1_outputs(5014) <= not (a or b);
    layer1_outputs(5015) <= not b;
    layer1_outputs(5016) <= b and not a;
    layer1_outputs(5017) <= not (a and b);
    layer1_outputs(5018) <= not (a or b);
    layer1_outputs(5019) <= not (a xor b);
    layer1_outputs(5020) <= not b or a;
    layer1_outputs(5021) <= a and not b;
    layer1_outputs(5022) <= '1';
    layer1_outputs(5023) <= '1';
    layer1_outputs(5024) <= not b;
    layer1_outputs(5025) <= a;
    layer1_outputs(5026) <= '1';
    layer1_outputs(5027) <= '0';
    layer1_outputs(5028) <= '0';
    layer1_outputs(5029) <= not b;
    layer1_outputs(5030) <= a and b;
    layer1_outputs(5031) <= a;
    layer1_outputs(5032) <= not a;
    layer1_outputs(5033) <= not a;
    layer1_outputs(5034) <= not a;
    layer1_outputs(5035) <= '1';
    layer1_outputs(5036) <= not (a or b);
    layer1_outputs(5037) <= b and not a;
    layer1_outputs(5038) <= '1';
    layer1_outputs(5039) <= a and not b;
    layer1_outputs(5040) <= '0';
    layer1_outputs(5041) <= b and not a;
    layer1_outputs(5042) <= a;
    layer1_outputs(5043) <= a and b;
    layer1_outputs(5044) <= not b;
    layer1_outputs(5045) <= not a;
    layer1_outputs(5046) <= not (a and b);
    layer1_outputs(5047) <= not a or b;
    layer1_outputs(5048) <= not (a and b);
    layer1_outputs(5049) <= '0';
    layer1_outputs(5050) <= '0';
    layer1_outputs(5051) <= a and b;
    layer1_outputs(5052) <= b and not a;
    layer1_outputs(5053) <= not (a or b);
    layer1_outputs(5054) <= a or b;
    layer1_outputs(5055) <= not a or b;
    layer1_outputs(5056) <= '1';
    layer1_outputs(5057) <= '0';
    layer1_outputs(5058) <= not b or a;
    layer1_outputs(5059) <= not b or a;
    layer1_outputs(5060) <= b;
    layer1_outputs(5061) <= '1';
    layer1_outputs(5062) <= not (a and b);
    layer1_outputs(5063) <= a and not b;
    layer1_outputs(5064) <= a and not b;
    layer1_outputs(5065) <= not (a or b);
    layer1_outputs(5066) <= b and not a;
    layer1_outputs(5067) <= '0';
    layer1_outputs(5068) <= not a;
    layer1_outputs(5069) <= '0';
    layer1_outputs(5070) <= not (a xor b);
    layer1_outputs(5071) <= not a;
    layer1_outputs(5072) <= '1';
    layer1_outputs(5073) <= not (a xor b);
    layer1_outputs(5074) <= a;
    layer1_outputs(5075) <= not (a or b);
    layer1_outputs(5076) <= '1';
    layer1_outputs(5077) <= not b or a;
    layer1_outputs(5078) <= not (a or b);
    layer1_outputs(5079) <= '1';
    layer1_outputs(5080) <= b and not a;
    layer1_outputs(5081) <= not a;
    layer1_outputs(5082) <= not a or b;
    layer1_outputs(5083) <= not (a and b);
    layer1_outputs(5084) <= a and not b;
    layer1_outputs(5085) <= '0';
    layer1_outputs(5086) <= a and b;
    layer1_outputs(5087) <= not a or b;
    layer1_outputs(5088) <= not (a or b);
    layer1_outputs(5089) <= not (a and b);
    layer1_outputs(5090) <= a and b;
    layer1_outputs(5091) <= b;
    layer1_outputs(5092) <= a and not b;
    layer1_outputs(5093) <= not b;
    layer1_outputs(5094) <= not a or b;
    layer1_outputs(5095) <= b and not a;
    layer1_outputs(5096) <= not b;
    layer1_outputs(5097) <= a or b;
    layer1_outputs(5098) <= not a;
    layer1_outputs(5099) <= not a or b;
    layer1_outputs(5100) <= a and b;
    layer1_outputs(5101) <= not (a xor b);
    layer1_outputs(5102) <= a xor b;
    layer1_outputs(5103) <= not (a or b);
    layer1_outputs(5104) <= not a or b;
    layer1_outputs(5105) <= a and not b;
    layer1_outputs(5106) <= '1';
    layer1_outputs(5107) <= a;
    layer1_outputs(5108) <= a and not b;
    layer1_outputs(5109) <= not b;
    layer1_outputs(5110) <= not b;
    layer1_outputs(5111) <= a;
    layer1_outputs(5112) <= '1';
    layer1_outputs(5113) <= not b;
    layer1_outputs(5114) <= '0';
    layer1_outputs(5115) <= '1';
    layer1_outputs(5116) <= not (a xor b);
    layer1_outputs(5117) <= b and not a;
    layer1_outputs(5118) <= not a;
    layer1_outputs(5119) <= not a;
    layer1_outputs(5120) <= b and not a;
    layer1_outputs(5121) <= not a or b;
    layer1_outputs(5122) <= a and b;
    layer1_outputs(5123) <= not (a and b);
    layer1_outputs(5124) <= not b;
    layer1_outputs(5125) <= '0';
    layer1_outputs(5126) <= not (a and b);
    layer1_outputs(5127) <= not b or a;
    layer1_outputs(5128) <= not a or b;
    layer1_outputs(5129) <= '1';
    layer1_outputs(5130) <= a and b;
    layer1_outputs(5131) <= not b or a;
    layer1_outputs(5132) <= a xor b;
    layer1_outputs(5133) <= not b;
    layer1_outputs(5134) <= '1';
    layer1_outputs(5135) <= not a;
    layer1_outputs(5136) <= '0';
    layer1_outputs(5137) <= not (a or b);
    layer1_outputs(5138) <= not (a or b);
    layer1_outputs(5139) <= b and not a;
    layer1_outputs(5140) <= a and not b;
    layer1_outputs(5141) <= b;
    layer1_outputs(5142) <= a;
    layer1_outputs(5143) <= a and b;
    layer1_outputs(5144) <= not a or b;
    layer1_outputs(5145) <= a and not b;
    layer1_outputs(5146) <= b;
    layer1_outputs(5147) <= a and not b;
    layer1_outputs(5148) <= not (a xor b);
    layer1_outputs(5149) <= not b or a;
    layer1_outputs(5150) <= '0';
    layer1_outputs(5151) <= not (a or b);
    layer1_outputs(5152) <= not (a and b);
    layer1_outputs(5153) <= a xor b;
    layer1_outputs(5154) <= b;
    layer1_outputs(5155) <= '0';
    layer1_outputs(5156) <= not a;
    layer1_outputs(5157) <= b and not a;
    layer1_outputs(5158) <= a and not b;
    layer1_outputs(5159) <= not (a or b);
    layer1_outputs(5160) <= '0';
    layer1_outputs(5161) <= a or b;
    layer1_outputs(5162) <= '0';
    layer1_outputs(5163) <= '0';
    layer1_outputs(5164) <= b;
    layer1_outputs(5165) <= not b;
    layer1_outputs(5166) <= b;
    layer1_outputs(5167) <= a or b;
    layer1_outputs(5168) <= '0';
    layer1_outputs(5169) <= '0';
    layer1_outputs(5170) <= not a or b;
    layer1_outputs(5171) <= a xor b;
    layer1_outputs(5172) <= '0';
    layer1_outputs(5173) <= a and not b;
    layer1_outputs(5174) <= b;
    layer1_outputs(5175) <= not a or b;
    layer1_outputs(5176) <= not a or b;
    layer1_outputs(5177) <= '0';
    layer1_outputs(5178) <= not b;
    layer1_outputs(5179) <= not a;
    layer1_outputs(5180) <= a or b;
    layer1_outputs(5181) <= not b;
    layer1_outputs(5182) <= a;
    layer1_outputs(5183) <= b and not a;
    layer1_outputs(5184) <= '1';
    layer1_outputs(5185) <= not (a or b);
    layer1_outputs(5186) <= a and not b;
    layer1_outputs(5187) <= not b;
    layer1_outputs(5188) <= a and not b;
    layer1_outputs(5189) <= not (a or b);
    layer1_outputs(5190) <= a or b;
    layer1_outputs(5191) <= a and not b;
    layer1_outputs(5192) <= '1';
    layer1_outputs(5193) <= not a or b;
    layer1_outputs(5194) <= not a;
    layer1_outputs(5195) <= b and not a;
    layer1_outputs(5196) <= b;
    layer1_outputs(5197) <= a and not b;
    layer1_outputs(5198) <= a xor b;
    layer1_outputs(5199) <= b;
    layer1_outputs(5200) <= not a or b;
    layer1_outputs(5201) <= a and b;
    layer1_outputs(5202) <= not (a and b);
    layer1_outputs(5203) <= a;
    layer1_outputs(5204) <= not b;
    layer1_outputs(5205) <= '1';
    layer1_outputs(5206) <= a and not b;
    layer1_outputs(5207) <= not a or b;
    layer1_outputs(5208) <= a and b;
    layer1_outputs(5209) <= not a;
    layer1_outputs(5210) <= '0';
    layer1_outputs(5211) <= a and b;
    layer1_outputs(5212) <= not (a or b);
    layer1_outputs(5213) <= b;
    layer1_outputs(5214) <= not a or b;
    layer1_outputs(5215) <= a;
    layer1_outputs(5216) <= not a;
    layer1_outputs(5217) <= a;
    layer1_outputs(5218) <= not b;
    layer1_outputs(5219) <= a and not b;
    layer1_outputs(5220) <= '0';
    layer1_outputs(5221) <= not b;
    layer1_outputs(5222) <= a and b;
    layer1_outputs(5223) <= not a or b;
    layer1_outputs(5224) <= a;
    layer1_outputs(5225) <= a or b;
    layer1_outputs(5226) <= a;
    layer1_outputs(5227) <= a and not b;
    layer1_outputs(5228) <= a and b;
    layer1_outputs(5229) <= not (a and b);
    layer1_outputs(5230) <= not (a or b);
    layer1_outputs(5231) <= not (a or b);
    layer1_outputs(5232) <= b and not a;
    layer1_outputs(5233) <= a and b;
    layer1_outputs(5234) <= '0';
    layer1_outputs(5235) <= b;
    layer1_outputs(5236) <= a or b;
    layer1_outputs(5237) <= not b;
    layer1_outputs(5238) <= b and not a;
    layer1_outputs(5239) <= a and not b;
    layer1_outputs(5240) <= a or b;
    layer1_outputs(5241) <= a and b;
    layer1_outputs(5242) <= not (a or b);
    layer1_outputs(5243) <= b;
    layer1_outputs(5244) <= not (a or b);
    layer1_outputs(5245) <= b and not a;
    layer1_outputs(5246) <= a or b;
    layer1_outputs(5247) <= not a;
    layer1_outputs(5248) <= a and b;
    layer1_outputs(5249) <= not (a and b);
    layer1_outputs(5250) <= '0';
    layer1_outputs(5251) <= '1';
    layer1_outputs(5252) <= '0';
    layer1_outputs(5253) <= not b or a;
    layer1_outputs(5254) <= '1';
    layer1_outputs(5255) <= a or b;
    layer1_outputs(5256) <= a;
    layer1_outputs(5257) <= not (a and b);
    layer1_outputs(5258) <= b and not a;
    layer1_outputs(5259) <= not a or b;
    layer1_outputs(5260) <= not b;
    layer1_outputs(5261) <= not b;
    layer1_outputs(5262) <= '1';
    layer1_outputs(5263) <= '0';
    layer1_outputs(5264) <= '0';
    layer1_outputs(5265) <= '1';
    layer1_outputs(5266) <= a and not b;
    layer1_outputs(5267) <= not a or b;
    layer1_outputs(5268) <= a and not b;
    layer1_outputs(5269) <= not (a and b);
    layer1_outputs(5270) <= a;
    layer1_outputs(5271) <= b and not a;
    layer1_outputs(5272) <= a and not b;
    layer1_outputs(5273) <= not b or a;
    layer1_outputs(5274) <= '1';
    layer1_outputs(5275) <= a or b;
    layer1_outputs(5276) <= not a;
    layer1_outputs(5277) <= a xor b;
    layer1_outputs(5278) <= not (a or b);
    layer1_outputs(5279) <= a;
    layer1_outputs(5280) <= a;
    layer1_outputs(5281) <= b;
    layer1_outputs(5282) <= not b;
    layer1_outputs(5283) <= a or b;
    layer1_outputs(5284) <= a;
    layer1_outputs(5285) <= '1';
    layer1_outputs(5286) <= a;
    layer1_outputs(5287) <= not a or b;
    layer1_outputs(5288) <= b and not a;
    layer1_outputs(5289) <= not b or a;
    layer1_outputs(5290) <= a or b;
    layer1_outputs(5291) <= not b;
    layer1_outputs(5292) <= a;
    layer1_outputs(5293) <= '1';
    layer1_outputs(5294) <= a and not b;
    layer1_outputs(5295) <= '1';
    layer1_outputs(5296) <= a and not b;
    layer1_outputs(5297) <= not (a and b);
    layer1_outputs(5298) <= b and not a;
    layer1_outputs(5299) <= a and b;
    layer1_outputs(5300) <= b;
    layer1_outputs(5301) <= a or b;
    layer1_outputs(5302) <= a and b;
    layer1_outputs(5303) <= not b or a;
    layer1_outputs(5304) <= not a;
    layer1_outputs(5305) <= not a;
    layer1_outputs(5306) <= a xor b;
    layer1_outputs(5307) <= not (a or b);
    layer1_outputs(5308) <= a and not b;
    layer1_outputs(5309) <= a and b;
    layer1_outputs(5310) <= not (a or b);
    layer1_outputs(5311) <= not a or b;
    layer1_outputs(5312) <= '1';
    layer1_outputs(5313) <= '0';
    layer1_outputs(5314) <= a;
    layer1_outputs(5315) <= a or b;
    layer1_outputs(5316) <= a;
    layer1_outputs(5317) <= b;
    layer1_outputs(5318) <= '1';
    layer1_outputs(5319) <= b and not a;
    layer1_outputs(5320) <= a or b;
    layer1_outputs(5321) <= a and b;
    layer1_outputs(5322) <= b and not a;
    layer1_outputs(5323) <= not a;
    layer1_outputs(5324) <= '0';
    layer1_outputs(5325) <= not b or a;
    layer1_outputs(5326) <= not (a and b);
    layer1_outputs(5327) <= not b;
    layer1_outputs(5328) <= '1';
    layer1_outputs(5329) <= a and not b;
    layer1_outputs(5330) <= not b;
    layer1_outputs(5331) <= not (a and b);
    layer1_outputs(5332) <= a or b;
    layer1_outputs(5333) <= not (a and b);
    layer1_outputs(5334) <= not b;
    layer1_outputs(5335) <= b and not a;
    layer1_outputs(5336) <= not a or b;
    layer1_outputs(5337) <= not b or a;
    layer1_outputs(5338) <= a;
    layer1_outputs(5339) <= '1';
    layer1_outputs(5340) <= not a;
    layer1_outputs(5341) <= not b;
    layer1_outputs(5342) <= a or b;
    layer1_outputs(5343) <= not (a xor b);
    layer1_outputs(5344) <= not b;
    layer1_outputs(5345) <= not a;
    layer1_outputs(5346) <= b and not a;
    layer1_outputs(5347) <= b;
    layer1_outputs(5348) <= not a or b;
    layer1_outputs(5349) <= a and b;
    layer1_outputs(5350) <= not (a or b);
    layer1_outputs(5351) <= a and b;
    layer1_outputs(5352) <= b;
    layer1_outputs(5353) <= not a or b;
    layer1_outputs(5354) <= '0';
    layer1_outputs(5355) <= a;
    layer1_outputs(5356) <= not a;
    layer1_outputs(5357) <= '1';
    layer1_outputs(5358) <= not a or b;
    layer1_outputs(5359) <= not b or a;
    layer1_outputs(5360) <= not a;
    layer1_outputs(5361) <= b and not a;
    layer1_outputs(5362) <= a and not b;
    layer1_outputs(5363) <= '0';
    layer1_outputs(5364) <= '1';
    layer1_outputs(5365) <= b and not a;
    layer1_outputs(5366) <= not a;
    layer1_outputs(5367) <= a or b;
    layer1_outputs(5368) <= not (a and b);
    layer1_outputs(5369) <= not b;
    layer1_outputs(5370) <= a or b;
    layer1_outputs(5371) <= '1';
    layer1_outputs(5372) <= not (a xor b);
    layer1_outputs(5373) <= not a or b;
    layer1_outputs(5374) <= a xor b;
    layer1_outputs(5375) <= not a or b;
    layer1_outputs(5376) <= not a or b;
    layer1_outputs(5377) <= not b or a;
    layer1_outputs(5378) <= '1';
    layer1_outputs(5379) <= not a or b;
    layer1_outputs(5380) <= not (a and b);
    layer1_outputs(5381) <= a or b;
    layer1_outputs(5382) <= not (a and b);
    layer1_outputs(5383) <= b;
    layer1_outputs(5384) <= '1';
    layer1_outputs(5385) <= not (a and b);
    layer1_outputs(5386) <= not (a and b);
    layer1_outputs(5387) <= b and not a;
    layer1_outputs(5388) <= a and not b;
    layer1_outputs(5389) <= not b or a;
    layer1_outputs(5390) <= a or b;
    layer1_outputs(5391) <= a xor b;
    layer1_outputs(5392) <= b and not a;
    layer1_outputs(5393) <= not (a xor b);
    layer1_outputs(5394) <= b;
    layer1_outputs(5395) <= '1';
    layer1_outputs(5396) <= not (a xor b);
    layer1_outputs(5397) <= not a or b;
    layer1_outputs(5398) <= not (a or b);
    layer1_outputs(5399) <= a and b;
    layer1_outputs(5400) <= not a or b;
    layer1_outputs(5401) <= not b or a;
    layer1_outputs(5402) <= not (a or b);
    layer1_outputs(5403) <= not b;
    layer1_outputs(5404) <= a xor b;
    layer1_outputs(5405) <= '0';
    layer1_outputs(5406) <= not (a xor b);
    layer1_outputs(5407) <= a;
    layer1_outputs(5408) <= not (a and b);
    layer1_outputs(5409) <= a and b;
    layer1_outputs(5410) <= not b;
    layer1_outputs(5411) <= not b or a;
    layer1_outputs(5412) <= not (a xor b);
    layer1_outputs(5413) <= not (a or b);
    layer1_outputs(5414) <= a and b;
    layer1_outputs(5415) <= a;
    layer1_outputs(5416) <= not (a xor b);
    layer1_outputs(5417) <= '1';
    layer1_outputs(5418) <= not b or a;
    layer1_outputs(5419) <= a xor b;
    layer1_outputs(5420) <= not (a and b);
    layer1_outputs(5421) <= '1';
    layer1_outputs(5422) <= not (a or b);
    layer1_outputs(5423) <= a and not b;
    layer1_outputs(5424) <= a and b;
    layer1_outputs(5425) <= '1';
    layer1_outputs(5426) <= '0';
    layer1_outputs(5427) <= '1';
    layer1_outputs(5428) <= not b or a;
    layer1_outputs(5429) <= '0';
    layer1_outputs(5430) <= not (a xor b);
    layer1_outputs(5431) <= b;
    layer1_outputs(5432) <= not (a and b);
    layer1_outputs(5433) <= b and not a;
    layer1_outputs(5434) <= '1';
    layer1_outputs(5435) <= not (a xor b);
    layer1_outputs(5436) <= '1';
    layer1_outputs(5437) <= '0';
    layer1_outputs(5438) <= not b;
    layer1_outputs(5439) <= '1';
    layer1_outputs(5440) <= b;
    layer1_outputs(5441) <= not b;
    layer1_outputs(5442) <= not a;
    layer1_outputs(5443) <= b and not a;
    layer1_outputs(5444) <= not a;
    layer1_outputs(5445) <= a and not b;
    layer1_outputs(5446) <= a;
    layer1_outputs(5447) <= a or b;
    layer1_outputs(5448) <= b and not a;
    layer1_outputs(5449) <= a and b;
    layer1_outputs(5450) <= a;
    layer1_outputs(5451) <= not a;
    layer1_outputs(5452) <= not b;
    layer1_outputs(5453) <= a;
    layer1_outputs(5454) <= a and not b;
    layer1_outputs(5455) <= a;
    layer1_outputs(5456) <= not a;
    layer1_outputs(5457) <= not (a and b);
    layer1_outputs(5458) <= '1';
    layer1_outputs(5459) <= b;
    layer1_outputs(5460) <= '0';
    layer1_outputs(5461) <= not b;
    layer1_outputs(5462) <= a and not b;
    layer1_outputs(5463) <= not a;
    layer1_outputs(5464) <= not b;
    layer1_outputs(5465) <= a and not b;
    layer1_outputs(5466) <= not (a and b);
    layer1_outputs(5467) <= not b or a;
    layer1_outputs(5468) <= not a;
    layer1_outputs(5469) <= b;
    layer1_outputs(5470) <= b and not a;
    layer1_outputs(5471) <= '1';
    layer1_outputs(5472) <= not a;
    layer1_outputs(5473) <= not a;
    layer1_outputs(5474) <= a and b;
    layer1_outputs(5475) <= a or b;
    layer1_outputs(5476) <= not b or a;
    layer1_outputs(5477) <= not a;
    layer1_outputs(5478) <= not a or b;
    layer1_outputs(5479) <= a or b;
    layer1_outputs(5480) <= '0';
    layer1_outputs(5481) <= not b;
    layer1_outputs(5482) <= a xor b;
    layer1_outputs(5483) <= not (a or b);
    layer1_outputs(5484) <= b and not a;
    layer1_outputs(5485) <= not b;
    layer1_outputs(5486) <= not b;
    layer1_outputs(5487) <= not b;
    layer1_outputs(5488) <= '1';
    layer1_outputs(5489) <= b and not a;
    layer1_outputs(5490) <= a and b;
    layer1_outputs(5491) <= '0';
    layer1_outputs(5492) <= not b;
    layer1_outputs(5493) <= not (a or b);
    layer1_outputs(5494) <= a and b;
    layer1_outputs(5495) <= not (a and b);
    layer1_outputs(5496) <= '1';
    layer1_outputs(5497) <= a;
    layer1_outputs(5498) <= b and not a;
    layer1_outputs(5499) <= '1';
    layer1_outputs(5500) <= not b;
    layer1_outputs(5501) <= not (a and b);
    layer1_outputs(5502) <= a or b;
    layer1_outputs(5503) <= not a or b;
    layer1_outputs(5504) <= not a;
    layer1_outputs(5505) <= '1';
    layer1_outputs(5506) <= a and not b;
    layer1_outputs(5507) <= '0';
    layer1_outputs(5508) <= b and not a;
    layer1_outputs(5509) <= not a;
    layer1_outputs(5510) <= not a;
    layer1_outputs(5511) <= not b;
    layer1_outputs(5512) <= b and not a;
    layer1_outputs(5513) <= a and b;
    layer1_outputs(5514) <= a and not b;
    layer1_outputs(5515) <= not (a and b);
    layer1_outputs(5516) <= not b;
    layer1_outputs(5517) <= '0';
    layer1_outputs(5518) <= b and not a;
    layer1_outputs(5519) <= b;
    layer1_outputs(5520) <= not b;
    layer1_outputs(5521) <= a xor b;
    layer1_outputs(5522) <= a or b;
    layer1_outputs(5523) <= a and b;
    layer1_outputs(5524) <= not a;
    layer1_outputs(5525) <= '1';
    layer1_outputs(5526) <= '1';
    layer1_outputs(5527) <= b and not a;
    layer1_outputs(5528) <= a and b;
    layer1_outputs(5529) <= b;
    layer1_outputs(5530) <= not (a and b);
    layer1_outputs(5531) <= b and not a;
    layer1_outputs(5532) <= '0';
    layer1_outputs(5533) <= not (a xor b);
    layer1_outputs(5534) <= a and b;
    layer1_outputs(5535) <= '0';
    layer1_outputs(5536) <= b;
    layer1_outputs(5537) <= b and not a;
    layer1_outputs(5538) <= '1';
    layer1_outputs(5539) <= not b;
    layer1_outputs(5540) <= not a or b;
    layer1_outputs(5541) <= not (a xor b);
    layer1_outputs(5542) <= b;
    layer1_outputs(5543) <= b;
    layer1_outputs(5544) <= b and not a;
    layer1_outputs(5545) <= '1';
    layer1_outputs(5546) <= not a or b;
    layer1_outputs(5547) <= a or b;
    layer1_outputs(5548) <= not (a or b);
    layer1_outputs(5549) <= b and not a;
    layer1_outputs(5550) <= not b;
    layer1_outputs(5551) <= not b or a;
    layer1_outputs(5552) <= not b;
    layer1_outputs(5553) <= '0';
    layer1_outputs(5554) <= a xor b;
    layer1_outputs(5555) <= not a or b;
    layer1_outputs(5556) <= '0';
    layer1_outputs(5557) <= not b;
    layer1_outputs(5558) <= not a;
    layer1_outputs(5559) <= '0';
    layer1_outputs(5560) <= '0';
    layer1_outputs(5561) <= '1';
    layer1_outputs(5562) <= not a or b;
    layer1_outputs(5563) <= a xor b;
    layer1_outputs(5564) <= not b;
    layer1_outputs(5565) <= not b;
    layer1_outputs(5566) <= not (a or b);
    layer1_outputs(5567) <= a;
    layer1_outputs(5568) <= b;
    layer1_outputs(5569) <= a or b;
    layer1_outputs(5570) <= not (a xor b);
    layer1_outputs(5571) <= not (a and b);
    layer1_outputs(5572) <= b and not a;
    layer1_outputs(5573) <= '0';
    layer1_outputs(5574) <= not a or b;
    layer1_outputs(5575) <= b;
    layer1_outputs(5576) <= b and not a;
    layer1_outputs(5577) <= not a or b;
    layer1_outputs(5578) <= b and not a;
    layer1_outputs(5579) <= a or b;
    layer1_outputs(5580) <= not a or b;
    layer1_outputs(5581) <= b;
    layer1_outputs(5582) <= a and b;
    layer1_outputs(5583) <= not a;
    layer1_outputs(5584) <= a or b;
    layer1_outputs(5585) <= '0';
    layer1_outputs(5586) <= '0';
    layer1_outputs(5587) <= '1';
    layer1_outputs(5588) <= a and b;
    layer1_outputs(5589) <= not (a or b);
    layer1_outputs(5590) <= '1';
    layer1_outputs(5591) <= not (a xor b);
    layer1_outputs(5592) <= not a or b;
    layer1_outputs(5593) <= not (a or b);
    layer1_outputs(5594) <= not (a and b);
    layer1_outputs(5595) <= a and not b;
    layer1_outputs(5596) <= a;
    layer1_outputs(5597) <= not a or b;
    layer1_outputs(5598) <= not a or b;
    layer1_outputs(5599) <= not (a or b);
    layer1_outputs(5600) <= not a;
    layer1_outputs(5601) <= a and b;
    layer1_outputs(5602) <= not a or b;
    layer1_outputs(5603) <= a or b;
    layer1_outputs(5604) <= not a;
    layer1_outputs(5605) <= a or b;
    layer1_outputs(5606) <= b and not a;
    layer1_outputs(5607) <= a and not b;
    layer1_outputs(5608) <= a;
    layer1_outputs(5609) <= not a or b;
    layer1_outputs(5610) <= not (a xor b);
    layer1_outputs(5611) <= a or b;
    layer1_outputs(5612) <= not b or a;
    layer1_outputs(5613) <= a and not b;
    layer1_outputs(5614) <= a or b;
    layer1_outputs(5615) <= not a;
    layer1_outputs(5616) <= not a or b;
    layer1_outputs(5617) <= a and b;
    layer1_outputs(5618) <= a;
    layer1_outputs(5619) <= not a;
    layer1_outputs(5620) <= a and not b;
    layer1_outputs(5621) <= a and not b;
    layer1_outputs(5622) <= a xor b;
    layer1_outputs(5623) <= '0';
    layer1_outputs(5624) <= b;
    layer1_outputs(5625) <= a;
    layer1_outputs(5626) <= not b;
    layer1_outputs(5627) <= not (a or b);
    layer1_outputs(5628) <= a or b;
    layer1_outputs(5629) <= '0';
    layer1_outputs(5630) <= a or b;
    layer1_outputs(5631) <= not a;
    layer1_outputs(5632) <= not (a and b);
    layer1_outputs(5633) <= not b;
    layer1_outputs(5634) <= not a or b;
    layer1_outputs(5635) <= not (a and b);
    layer1_outputs(5636) <= not a or b;
    layer1_outputs(5637) <= a or b;
    layer1_outputs(5638) <= not (a and b);
    layer1_outputs(5639) <= b;
    layer1_outputs(5640) <= '0';
    layer1_outputs(5641) <= not (a and b);
    layer1_outputs(5642) <= a and b;
    layer1_outputs(5643) <= not (a or b);
    layer1_outputs(5644) <= not (a xor b);
    layer1_outputs(5645) <= a or b;
    layer1_outputs(5646) <= not b or a;
    layer1_outputs(5647) <= b and not a;
    layer1_outputs(5648) <= '1';
    layer1_outputs(5649) <= not b;
    layer1_outputs(5650) <= not (a and b);
    layer1_outputs(5651) <= a;
    layer1_outputs(5652) <= a or b;
    layer1_outputs(5653) <= '0';
    layer1_outputs(5654) <= not b or a;
    layer1_outputs(5655) <= '1';
    layer1_outputs(5656) <= not (a and b);
    layer1_outputs(5657) <= not b;
    layer1_outputs(5658) <= '0';
    layer1_outputs(5659) <= '0';
    layer1_outputs(5660) <= not a;
    layer1_outputs(5661) <= a;
    layer1_outputs(5662) <= b;
    layer1_outputs(5663) <= not a;
    layer1_outputs(5664) <= a or b;
    layer1_outputs(5665) <= not a or b;
    layer1_outputs(5666) <= b and not a;
    layer1_outputs(5667) <= not a;
    layer1_outputs(5668) <= not a;
    layer1_outputs(5669) <= not b or a;
    layer1_outputs(5670) <= not a;
    layer1_outputs(5671) <= not b;
    layer1_outputs(5672) <= '0';
    layer1_outputs(5673) <= a and not b;
    layer1_outputs(5674) <= a;
    layer1_outputs(5675) <= a and b;
    layer1_outputs(5676) <= not b;
    layer1_outputs(5677) <= b and not a;
    layer1_outputs(5678) <= not (a or b);
    layer1_outputs(5679) <= '0';
    layer1_outputs(5680) <= b;
    layer1_outputs(5681) <= b;
    layer1_outputs(5682) <= b and not a;
    layer1_outputs(5683) <= b and not a;
    layer1_outputs(5684) <= not (a or b);
    layer1_outputs(5685) <= a xor b;
    layer1_outputs(5686) <= not b or a;
    layer1_outputs(5687) <= b and not a;
    layer1_outputs(5688) <= not (a or b);
    layer1_outputs(5689) <= '0';
    layer1_outputs(5690) <= not b or a;
    layer1_outputs(5691) <= not (a or b);
    layer1_outputs(5692) <= a;
    layer1_outputs(5693) <= b;
    layer1_outputs(5694) <= not (a or b);
    layer1_outputs(5695) <= b;
    layer1_outputs(5696) <= '1';
    layer1_outputs(5697) <= not b or a;
    layer1_outputs(5698) <= b;
    layer1_outputs(5699) <= a;
    layer1_outputs(5700) <= not a;
    layer1_outputs(5701) <= a and b;
    layer1_outputs(5702) <= not b;
    layer1_outputs(5703) <= a;
    layer1_outputs(5704) <= not b;
    layer1_outputs(5705) <= '0';
    layer1_outputs(5706) <= not (a or b);
    layer1_outputs(5707) <= '1';
    layer1_outputs(5708) <= not b;
    layer1_outputs(5709) <= b and not a;
    layer1_outputs(5710) <= not b;
    layer1_outputs(5711) <= not b;
    layer1_outputs(5712) <= a xor b;
    layer1_outputs(5713) <= a;
    layer1_outputs(5714) <= b;
    layer1_outputs(5715) <= a;
    layer1_outputs(5716) <= not a;
    layer1_outputs(5717) <= not (a or b);
    layer1_outputs(5718) <= '0';
    layer1_outputs(5719) <= '0';
    layer1_outputs(5720) <= not (a and b);
    layer1_outputs(5721) <= not b;
    layer1_outputs(5722) <= not b;
    layer1_outputs(5723) <= b;
    layer1_outputs(5724) <= b;
    layer1_outputs(5725) <= not (a or b);
    layer1_outputs(5726) <= b;
    layer1_outputs(5727) <= a and b;
    layer1_outputs(5728) <= a or b;
    layer1_outputs(5729) <= not (a or b);
    layer1_outputs(5730) <= not (a or b);
    layer1_outputs(5731) <= b and not a;
    layer1_outputs(5732) <= a and b;
    layer1_outputs(5733) <= a and b;
    layer1_outputs(5734) <= '1';
    layer1_outputs(5735) <= not (a or b);
    layer1_outputs(5736) <= not (a xor b);
    layer1_outputs(5737) <= not b or a;
    layer1_outputs(5738) <= not a;
    layer1_outputs(5739) <= a and not b;
    layer1_outputs(5740) <= not (a xor b);
    layer1_outputs(5741) <= '0';
    layer1_outputs(5742) <= not (a xor b);
    layer1_outputs(5743) <= a;
    layer1_outputs(5744) <= a;
    layer1_outputs(5745) <= not (a and b);
    layer1_outputs(5746) <= '0';
    layer1_outputs(5747) <= not a or b;
    layer1_outputs(5748) <= not b or a;
    layer1_outputs(5749) <= not b;
    layer1_outputs(5750) <= not (a and b);
    layer1_outputs(5751) <= a and b;
    layer1_outputs(5752) <= not (a and b);
    layer1_outputs(5753) <= b and not a;
    layer1_outputs(5754) <= a xor b;
    layer1_outputs(5755) <= a and b;
    layer1_outputs(5756) <= b and not a;
    layer1_outputs(5757) <= not b;
    layer1_outputs(5758) <= not a;
    layer1_outputs(5759) <= not a or b;
    layer1_outputs(5760) <= not (a and b);
    layer1_outputs(5761) <= '0';
    layer1_outputs(5762) <= '1';
    layer1_outputs(5763) <= not (a and b);
    layer1_outputs(5764) <= a and b;
    layer1_outputs(5765) <= a and b;
    layer1_outputs(5766) <= '1';
    layer1_outputs(5767) <= a and b;
    layer1_outputs(5768) <= '1';
    layer1_outputs(5769) <= not a or b;
    layer1_outputs(5770) <= not (a or b);
    layer1_outputs(5771) <= not b or a;
    layer1_outputs(5772) <= '1';
    layer1_outputs(5773) <= b;
    layer1_outputs(5774) <= b;
    layer1_outputs(5775) <= not b;
    layer1_outputs(5776) <= a;
    layer1_outputs(5777) <= not a or b;
    layer1_outputs(5778) <= a and not b;
    layer1_outputs(5779) <= a and b;
    layer1_outputs(5780) <= b;
    layer1_outputs(5781) <= not a;
    layer1_outputs(5782) <= not (a and b);
    layer1_outputs(5783) <= a;
    layer1_outputs(5784) <= not b or a;
    layer1_outputs(5785) <= not (a and b);
    layer1_outputs(5786) <= not a;
    layer1_outputs(5787) <= a or b;
    layer1_outputs(5788) <= a and b;
    layer1_outputs(5789) <= a and b;
    layer1_outputs(5790) <= a or b;
    layer1_outputs(5791) <= a or b;
    layer1_outputs(5792) <= '0';
    layer1_outputs(5793) <= '1';
    layer1_outputs(5794) <= not a or b;
    layer1_outputs(5795) <= '1';
    layer1_outputs(5796) <= not (a and b);
    layer1_outputs(5797) <= not a;
    layer1_outputs(5798) <= a and b;
    layer1_outputs(5799) <= b and not a;
    layer1_outputs(5800) <= not (a or b);
    layer1_outputs(5801) <= b and not a;
    layer1_outputs(5802) <= b and not a;
    layer1_outputs(5803) <= not a;
    layer1_outputs(5804) <= not (a or b);
    layer1_outputs(5805) <= '1';
    layer1_outputs(5806) <= b and not a;
    layer1_outputs(5807) <= a and not b;
    layer1_outputs(5808) <= not a;
    layer1_outputs(5809) <= a and b;
    layer1_outputs(5810) <= not a;
    layer1_outputs(5811) <= '1';
    layer1_outputs(5812) <= not (a or b);
    layer1_outputs(5813) <= a;
    layer1_outputs(5814) <= not (a or b);
    layer1_outputs(5815) <= a;
    layer1_outputs(5816) <= not a;
    layer1_outputs(5817) <= not (a or b);
    layer1_outputs(5818) <= '1';
    layer1_outputs(5819) <= '1';
    layer1_outputs(5820) <= a and b;
    layer1_outputs(5821) <= '0';
    layer1_outputs(5822) <= a;
    layer1_outputs(5823) <= '0';
    layer1_outputs(5824) <= not (a or b);
    layer1_outputs(5825) <= a;
    layer1_outputs(5826) <= a and b;
    layer1_outputs(5827) <= b and not a;
    layer1_outputs(5828) <= not b;
    layer1_outputs(5829) <= '0';
    layer1_outputs(5830) <= a;
    layer1_outputs(5831) <= '0';
    layer1_outputs(5832) <= not b or a;
    layer1_outputs(5833) <= '1';
    layer1_outputs(5834) <= not b;
    layer1_outputs(5835) <= not (a or b);
    layer1_outputs(5836) <= not b;
    layer1_outputs(5837) <= '0';
    layer1_outputs(5838) <= not a or b;
    layer1_outputs(5839) <= a and b;
    layer1_outputs(5840) <= b;
    layer1_outputs(5841) <= a;
    layer1_outputs(5842) <= not a or b;
    layer1_outputs(5843) <= b and not a;
    layer1_outputs(5844) <= b;
    layer1_outputs(5845) <= a xor b;
    layer1_outputs(5846) <= not b;
    layer1_outputs(5847) <= a and b;
    layer1_outputs(5848) <= '1';
    layer1_outputs(5849) <= not a or b;
    layer1_outputs(5850) <= b;
    layer1_outputs(5851) <= not b;
    layer1_outputs(5852) <= not b;
    layer1_outputs(5853) <= not a;
    layer1_outputs(5854) <= a xor b;
    layer1_outputs(5855) <= '0';
    layer1_outputs(5856) <= '1';
    layer1_outputs(5857) <= b and not a;
    layer1_outputs(5858) <= a or b;
    layer1_outputs(5859) <= '0';
    layer1_outputs(5860) <= '0';
    layer1_outputs(5861) <= a;
    layer1_outputs(5862) <= not a;
    layer1_outputs(5863) <= a and not b;
    layer1_outputs(5864) <= '1';
    layer1_outputs(5865) <= a;
    layer1_outputs(5866) <= not b;
    layer1_outputs(5867) <= '0';
    layer1_outputs(5868) <= a;
    layer1_outputs(5869) <= '0';
    layer1_outputs(5870) <= a and not b;
    layer1_outputs(5871) <= not a or b;
    layer1_outputs(5872) <= a;
    layer1_outputs(5873) <= '0';
    layer1_outputs(5874) <= a;
    layer1_outputs(5875) <= b;
    layer1_outputs(5876) <= a;
    layer1_outputs(5877) <= b and not a;
    layer1_outputs(5878) <= a;
    layer1_outputs(5879) <= not a;
    layer1_outputs(5880) <= a and not b;
    layer1_outputs(5881) <= a;
    layer1_outputs(5882) <= '0';
    layer1_outputs(5883) <= '1';
    layer1_outputs(5884) <= not (a or b);
    layer1_outputs(5885) <= b and not a;
    layer1_outputs(5886) <= '0';
    layer1_outputs(5887) <= not b;
    layer1_outputs(5888) <= b;
    layer1_outputs(5889) <= b and not a;
    layer1_outputs(5890) <= a or b;
    layer1_outputs(5891) <= not b or a;
    layer1_outputs(5892) <= '1';
    layer1_outputs(5893) <= not b or a;
    layer1_outputs(5894) <= not b or a;
    layer1_outputs(5895) <= not b or a;
    layer1_outputs(5896) <= a;
    layer1_outputs(5897) <= '1';
    layer1_outputs(5898) <= a;
    layer1_outputs(5899) <= not (a and b);
    layer1_outputs(5900) <= a;
    layer1_outputs(5901) <= b and not a;
    layer1_outputs(5902) <= not (a and b);
    layer1_outputs(5903) <= not (a or b);
    layer1_outputs(5904) <= a or b;
    layer1_outputs(5905) <= b;
    layer1_outputs(5906) <= '1';
    layer1_outputs(5907) <= not a or b;
    layer1_outputs(5908) <= '1';
    layer1_outputs(5909) <= b;
    layer1_outputs(5910) <= not a;
    layer1_outputs(5911) <= not (a xor b);
    layer1_outputs(5912) <= not (a and b);
    layer1_outputs(5913) <= a or b;
    layer1_outputs(5914) <= b;
    layer1_outputs(5915) <= not b;
    layer1_outputs(5916) <= '1';
    layer1_outputs(5917) <= not (a and b);
    layer1_outputs(5918) <= a or b;
    layer1_outputs(5919) <= a and b;
    layer1_outputs(5920) <= a and b;
    layer1_outputs(5921) <= a;
    layer1_outputs(5922) <= not a or b;
    layer1_outputs(5923) <= not (a or b);
    layer1_outputs(5924) <= a and b;
    layer1_outputs(5925) <= '0';
    layer1_outputs(5926) <= a and not b;
    layer1_outputs(5927) <= a and b;
    layer1_outputs(5928) <= not a or b;
    layer1_outputs(5929) <= b and not a;
    layer1_outputs(5930) <= '1';
    layer1_outputs(5931) <= '1';
    layer1_outputs(5932) <= a;
    layer1_outputs(5933) <= '0';
    layer1_outputs(5934) <= a xor b;
    layer1_outputs(5935) <= '0';
    layer1_outputs(5936) <= a;
    layer1_outputs(5937) <= not (a or b);
    layer1_outputs(5938) <= not (a and b);
    layer1_outputs(5939) <= b and not a;
    layer1_outputs(5940) <= a and not b;
    layer1_outputs(5941) <= not b or a;
    layer1_outputs(5942) <= '0';
    layer1_outputs(5943) <= '0';
    layer1_outputs(5944) <= b;
    layer1_outputs(5945) <= not a;
    layer1_outputs(5946) <= '1';
    layer1_outputs(5947) <= a and b;
    layer1_outputs(5948) <= a and b;
    layer1_outputs(5949) <= not (a and b);
    layer1_outputs(5950) <= '1';
    layer1_outputs(5951) <= a xor b;
    layer1_outputs(5952) <= not a;
    layer1_outputs(5953) <= not b or a;
    layer1_outputs(5954) <= b and not a;
    layer1_outputs(5955) <= not b;
    layer1_outputs(5956) <= not a or b;
    layer1_outputs(5957) <= b and not a;
    layer1_outputs(5958) <= b;
    layer1_outputs(5959) <= not a;
    layer1_outputs(5960) <= a;
    layer1_outputs(5961) <= not a or b;
    layer1_outputs(5962) <= not b;
    layer1_outputs(5963) <= not a or b;
    layer1_outputs(5964) <= not (a or b);
    layer1_outputs(5965) <= a xor b;
    layer1_outputs(5966) <= a and not b;
    layer1_outputs(5967) <= a or b;
    layer1_outputs(5968) <= '0';
    layer1_outputs(5969) <= a and not b;
    layer1_outputs(5970) <= a or b;
    layer1_outputs(5971) <= not (a or b);
    layer1_outputs(5972) <= not (a xor b);
    layer1_outputs(5973) <= not (a xor b);
    layer1_outputs(5974) <= '1';
    layer1_outputs(5975) <= not b or a;
    layer1_outputs(5976) <= not (a and b);
    layer1_outputs(5977) <= a xor b;
    layer1_outputs(5978) <= not a;
    layer1_outputs(5979) <= not b or a;
    layer1_outputs(5980) <= not a or b;
    layer1_outputs(5981) <= '1';
    layer1_outputs(5982) <= not a or b;
    layer1_outputs(5983) <= a or b;
    layer1_outputs(5984) <= b and not a;
    layer1_outputs(5985) <= not a or b;
    layer1_outputs(5986) <= '0';
    layer1_outputs(5987) <= a and not b;
    layer1_outputs(5988) <= b and not a;
    layer1_outputs(5989) <= not b or a;
    layer1_outputs(5990) <= not a or b;
    layer1_outputs(5991) <= b;
    layer1_outputs(5992) <= not a;
    layer1_outputs(5993) <= not (a or b);
    layer1_outputs(5994) <= a and b;
    layer1_outputs(5995) <= a and not b;
    layer1_outputs(5996) <= not (a or b);
    layer1_outputs(5997) <= not a;
    layer1_outputs(5998) <= not b;
    layer1_outputs(5999) <= '1';
    layer1_outputs(6000) <= '0';
    layer1_outputs(6001) <= '1';
    layer1_outputs(6002) <= '0';
    layer1_outputs(6003) <= a;
    layer1_outputs(6004) <= a xor b;
    layer1_outputs(6005) <= '1';
    layer1_outputs(6006) <= b and not a;
    layer1_outputs(6007) <= b and not a;
    layer1_outputs(6008) <= not a or b;
    layer1_outputs(6009) <= a xor b;
    layer1_outputs(6010) <= a and b;
    layer1_outputs(6011) <= a and not b;
    layer1_outputs(6012) <= b and not a;
    layer1_outputs(6013) <= not b or a;
    layer1_outputs(6014) <= not (a or b);
    layer1_outputs(6015) <= b;
    layer1_outputs(6016) <= a and not b;
    layer1_outputs(6017) <= not a;
    layer1_outputs(6018) <= '0';
    layer1_outputs(6019) <= a;
    layer1_outputs(6020) <= not (a and b);
    layer1_outputs(6021) <= a and not b;
    layer1_outputs(6022) <= b;
    layer1_outputs(6023) <= a;
    layer1_outputs(6024) <= '1';
    layer1_outputs(6025) <= a and b;
    layer1_outputs(6026) <= not (a or b);
    layer1_outputs(6027) <= a and not b;
    layer1_outputs(6028) <= a and b;
    layer1_outputs(6029) <= a;
    layer1_outputs(6030) <= not b;
    layer1_outputs(6031) <= b;
    layer1_outputs(6032) <= not b or a;
    layer1_outputs(6033) <= '0';
    layer1_outputs(6034) <= b;
    layer1_outputs(6035) <= not a or b;
    layer1_outputs(6036) <= not a or b;
    layer1_outputs(6037) <= a or b;
    layer1_outputs(6038) <= b and not a;
    layer1_outputs(6039) <= a or b;
    layer1_outputs(6040) <= not b or a;
    layer1_outputs(6041) <= a and not b;
    layer1_outputs(6042) <= a or b;
    layer1_outputs(6043) <= '0';
    layer1_outputs(6044) <= '0';
    layer1_outputs(6045) <= '0';
    layer1_outputs(6046) <= a and b;
    layer1_outputs(6047) <= '0';
    layer1_outputs(6048) <= not (a and b);
    layer1_outputs(6049) <= a xor b;
    layer1_outputs(6050) <= b;
    layer1_outputs(6051) <= not (a or b);
    layer1_outputs(6052) <= b and not a;
    layer1_outputs(6053) <= a;
    layer1_outputs(6054) <= b;
    layer1_outputs(6055) <= '1';
    layer1_outputs(6056) <= a or b;
    layer1_outputs(6057) <= not (a and b);
    layer1_outputs(6058) <= a and b;
    layer1_outputs(6059) <= not a;
    layer1_outputs(6060) <= not b;
    layer1_outputs(6061) <= b and not a;
    layer1_outputs(6062) <= '0';
    layer1_outputs(6063) <= not (a xor b);
    layer1_outputs(6064) <= a and b;
    layer1_outputs(6065) <= b and not a;
    layer1_outputs(6066) <= not a;
    layer1_outputs(6067) <= not a or b;
    layer1_outputs(6068) <= a or b;
    layer1_outputs(6069) <= not (a and b);
    layer1_outputs(6070) <= not (a or b);
    layer1_outputs(6071) <= a and b;
    layer1_outputs(6072) <= a and not b;
    layer1_outputs(6073) <= not b or a;
    layer1_outputs(6074) <= a xor b;
    layer1_outputs(6075) <= not (a and b);
    layer1_outputs(6076) <= not (a and b);
    layer1_outputs(6077) <= '1';
    layer1_outputs(6078) <= not a;
    layer1_outputs(6079) <= not (a and b);
    layer1_outputs(6080) <= not (a and b);
    layer1_outputs(6081) <= not b;
    layer1_outputs(6082) <= not (a or b);
    layer1_outputs(6083) <= '0';
    layer1_outputs(6084) <= b and not a;
    layer1_outputs(6085) <= not (a or b);
    layer1_outputs(6086) <= b;
    layer1_outputs(6087) <= b and not a;
    layer1_outputs(6088) <= '0';
    layer1_outputs(6089) <= b;
    layer1_outputs(6090) <= '0';
    layer1_outputs(6091) <= not a or b;
    layer1_outputs(6092) <= '1';
    layer1_outputs(6093) <= b and not a;
    layer1_outputs(6094) <= b;
    layer1_outputs(6095) <= b and not a;
    layer1_outputs(6096) <= a xor b;
    layer1_outputs(6097) <= not a or b;
    layer1_outputs(6098) <= '0';
    layer1_outputs(6099) <= not a or b;
    layer1_outputs(6100) <= not (a or b);
    layer1_outputs(6101) <= '1';
    layer1_outputs(6102) <= not (a xor b);
    layer1_outputs(6103) <= not a or b;
    layer1_outputs(6104) <= '1';
    layer1_outputs(6105) <= '0';
    layer1_outputs(6106) <= not b;
    layer1_outputs(6107) <= not (a or b);
    layer1_outputs(6108) <= not b or a;
    layer1_outputs(6109) <= b and not a;
    layer1_outputs(6110) <= a or b;
    layer1_outputs(6111) <= not a or b;
    layer1_outputs(6112) <= not (a or b);
    layer1_outputs(6113) <= not b or a;
    layer1_outputs(6114) <= not b or a;
    layer1_outputs(6115) <= a or b;
    layer1_outputs(6116) <= not a or b;
    layer1_outputs(6117) <= not (a or b);
    layer1_outputs(6118) <= a and b;
    layer1_outputs(6119) <= not a or b;
    layer1_outputs(6120) <= a and b;
    layer1_outputs(6121) <= b and not a;
    layer1_outputs(6122) <= b and not a;
    layer1_outputs(6123) <= b and not a;
    layer1_outputs(6124) <= not a or b;
    layer1_outputs(6125) <= a or b;
    layer1_outputs(6126) <= not a or b;
    layer1_outputs(6127) <= b;
    layer1_outputs(6128) <= a and b;
    layer1_outputs(6129) <= not (a xor b);
    layer1_outputs(6130) <= b;
    layer1_outputs(6131) <= b and not a;
    layer1_outputs(6132) <= not a;
    layer1_outputs(6133) <= not (a and b);
    layer1_outputs(6134) <= not a;
    layer1_outputs(6135) <= a;
    layer1_outputs(6136) <= not a or b;
    layer1_outputs(6137) <= not (a xor b);
    layer1_outputs(6138) <= not (a and b);
    layer1_outputs(6139) <= '0';
    layer1_outputs(6140) <= not (a xor b);
    layer1_outputs(6141) <= not (a or b);
    layer1_outputs(6142) <= a or b;
    layer1_outputs(6143) <= not a;
    layer1_outputs(6144) <= not (a or b);
    layer1_outputs(6145) <= not a;
    layer1_outputs(6146) <= not b or a;
    layer1_outputs(6147) <= not b or a;
    layer1_outputs(6148) <= '0';
    layer1_outputs(6149) <= b and not a;
    layer1_outputs(6150) <= a xor b;
    layer1_outputs(6151) <= not a or b;
    layer1_outputs(6152) <= '1';
    layer1_outputs(6153) <= not a;
    layer1_outputs(6154) <= b and not a;
    layer1_outputs(6155) <= not (a xor b);
    layer1_outputs(6156) <= not b or a;
    layer1_outputs(6157) <= a or b;
    layer1_outputs(6158) <= a xor b;
    layer1_outputs(6159) <= b;
    layer1_outputs(6160) <= not a;
    layer1_outputs(6161) <= a and not b;
    layer1_outputs(6162) <= not a or b;
    layer1_outputs(6163) <= b and not a;
    layer1_outputs(6164) <= a;
    layer1_outputs(6165) <= not b or a;
    layer1_outputs(6166) <= not b or a;
    layer1_outputs(6167) <= b;
    layer1_outputs(6168) <= not (a and b);
    layer1_outputs(6169) <= a and not b;
    layer1_outputs(6170) <= b and not a;
    layer1_outputs(6171) <= b;
    layer1_outputs(6172) <= '0';
    layer1_outputs(6173) <= not b;
    layer1_outputs(6174) <= b;
    layer1_outputs(6175) <= '0';
    layer1_outputs(6176) <= '1';
    layer1_outputs(6177) <= a and not b;
    layer1_outputs(6178) <= not (a and b);
    layer1_outputs(6179) <= not a or b;
    layer1_outputs(6180) <= a;
    layer1_outputs(6181) <= a and b;
    layer1_outputs(6182) <= a or b;
    layer1_outputs(6183) <= not a or b;
    layer1_outputs(6184) <= not b;
    layer1_outputs(6185) <= a or b;
    layer1_outputs(6186) <= b;
    layer1_outputs(6187) <= not a;
    layer1_outputs(6188) <= a and b;
    layer1_outputs(6189) <= a and not b;
    layer1_outputs(6190) <= a and b;
    layer1_outputs(6191) <= not b or a;
    layer1_outputs(6192) <= not a or b;
    layer1_outputs(6193) <= '1';
    layer1_outputs(6194) <= '0';
    layer1_outputs(6195) <= not (a or b);
    layer1_outputs(6196) <= a or b;
    layer1_outputs(6197) <= '0';
    layer1_outputs(6198) <= a xor b;
    layer1_outputs(6199) <= b;
    layer1_outputs(6200) <= b;
    layer1_outputs(6201) <= b and not a;
    layer1_outputs(6202) <= b and not a;
    layer1_outputs(6203) <= not b;
    layer1_outputs(6204) <= not (a and b);
    layer1_outputs(6205) <= a xor b;
    layer1_outputs(6206) <= b;
    layer1_outputs(6207) <= not b;
    layer1_outputs(6208) <= a and not b;
    layer1_outputs(6209) <= a;
    layer1_outputs(6210) <= a and b;
    layer1_outputs(6211) <= not b;
    layer1_outputs(6212) <= not (a or b);
    layer1_outputs(6213) <= b;
    layer1_outputs(6214) <= '1';
    layer1_outputs(6215) <= not (a or b);
    layer1_outputs(6216) <= b;
    layer1_outputs(6217) <= a or b;
    layer1_outputs(6218) <= not (a and b);
    layer1_outputs(6219) <= '1';
    layer1_outputs(6220) <= '0';
    layer1_outputs(6221) <= '0';
    layer1_outputs(6222) <= b;
    layer1_outputs(6223) <= not (a and b);
    layer1_outputs(6224) <= a and b;
    layer1_outputs(6225) <= b and not a;
    layer1_outputs(6226) <= not a or b;
    layer1_outputs(6227) <= '0';
    layer1_outputs(6228) <= not (a and b);
    layer1_outputs(6229) <= not b;
    layer1_outputs(6230) <= not b or a;
    layer1_outputs(6231) <= a and not b;
    layer1_outputs(6232) <= a xor b;
    layer1_outputs(6233) <= '1';
    layer1_outputs(6234) <= '0';
    layer1_outputs(6235) <= a or b;
    layer1_outputs(6236) <= not a;
    layer1_outputs(6237) <= not b;
    layer1_outputs(6238) <= b;
    layer1_outputs(6239) <= '0';
    layer1_outputs(6240) <= a and b;
    layer1_outputs(6241) <= a;
    layer1_outputs(6242) <= not b;
    layer1_outputs(6243) <= not (a or b);
    layer1_outputs(6244) <= a and b;
    layer1_outputs(6245) <= not a;
    layer1_outputs(6246) <= not (a and b);
    layer1_outputs(6247) <= not b;
    layer1_outputs(6248) <= '0';
    layer1_outputs(6249) <= '1';
    layer1_outputs(6250) <= a and b;
    layer1_outputs(6251) <= not a or b;
    layer1_outputs(6252) <= not b or a;
    layer1_outputs(6253) <= not (a or b);
    layer1_outputs(6254) <= a;
    layer1_outputs(6255) <= a xor b;
    layer1_outputs(6256) <= '1';
    layer1_outputs(6257) <= not a;
    layer1_outputs(6258) <= a and not b;
    layer1_outputs(6259) <= not b;
    layer1_outputs(6260) <= '0';
    layer1_outputs(6261) <= b;
    layer1_outputs(6262) <= not (a and b);
    layer1_outputs(6263) <= not b or a;
    layer1_outputs(6264) <= a and not b;
    layer1_outputs(6265) <= not b;
    layer1_outputs(6266) <= a and b;
    layer1_outputs(6267) <= not b;
    layer1_outputs(6268) <= a and not b;
    layer1_outputs(6269) <= '1';
    layer1_outputs(6270) <= not b or a;
    layer1_outputs(6271) <= '1';
    layer1_outputs(6272) <= not b;
    layer1_outputs(6273) <= not b;
    layer1_outputs(6274) <= '1';
    layer1_outputs(6275) <= not a;
    layer1_outputs(6276) <= '0';
    layer1_outputs(6277) <= not b or a;
    layer1_outputs(6278) <= not (a or b);
    layer1_outputs(6279) <= b and not a;
    layer1_outputs(6280) <= not a;
    layer1_outputs(6281) <= a and not b;
    layer1_outputs(6282) <= '0';
    layer1_outputs(6283) <= not (a xor b);
    layer1_outputs(6284) <= '1';
    layer1_outputs(6285) <= not (a and b);
    layer1_outputs(6286) <= not a;
    layer1_outputs(6287) <= a or b;
    layer1_outputs(6288) <= not (a xor b);
    layer1_outputs(6289) <= a and not b;
    layer1_outputs(6290) <= not (a and b);
    layer1_outputs(6291) <= b and not a;
    layer1_outputs(6292) <= not (a or b);
    layer1_outputs(6293) <= '1';
    layer1_outputs(6294) <= not b;
    layer1_outputs(6295) <= a or b;
    layer1_outputs(6296) <= not (a or b);
    layer1_outputs(6297) <= not (a or b);
    layer1_outputs(6298) <= a xor b;
    layer1_outputs(6299) <= not b or a;
    layer1_outputs(6300) <= b;
    layer1_outputs(6301) <= not (a and b);
    layer1_outputs(6302) <= a and b;
    layer1_outputs(6303) <= not (a or b);
    layer1_outputs(6304) <= not a;
    layer1_outputs(6305) <= b and not a;
    layer1_outputs(6306) <= '1';
    layer1_outputs(6307) <= a or b;
    layer1_outputs(6308) <= not (a xor b);
    layer1_outputs(6309) <= a and not b;
    layer1_outputs(6310) <= b;
    layer1_outputs(6311) <= not (a and b);
    layer1_outputs(6312) <= '0';
    layer1_outputs(6313) <= not a;
    layer1_outputs(6314) <= a and not b;
    layer1_outputs(6315) <= not (a or b);
    layer1_outputs(6316) <= not (a xor b);
    layer1_outputs(6317) <= not (a or b);
    layer1_outputs(6318) <= a and b;
    layer1_outputs(6319) <= '1';
    layer1_outputs(6320) <= b;
    layer1_outputs(6321) <= b and not a;
    layer1_outputs(6322) <= not a or b;
    layer1_outputs(6323) <= '0';
    layer1_outputs(6324) <= b;
    layer1_outputs(6325) <= not (a and b);
    layer1_outputs(6326) <= not (a or b);
    layer1_outputs(6327) <= a and not b;
    layer1_outputs(6328) <= not a;
    layer1_outputs(6329) <= not a;
    layer1_outputs(6330) <= '1';
    layer1_outputs(6331) <= '1';
    layer1_outputs(6332) <= a and b;
    layer1_outputs(6333) <= b;
    layer1_outputs(6334) <= a;
    layer1_outputs(6335) <= not a;
    layer1_outputs(6336) <= a and not b;
    layer1_outputs(6337) <= '1';
    layer1_outputs(6338) <= '0';
    layer1_outputs(6339) <= not (a or b);
    layer1_outputs(6340) <= not (a and b);
    layer1_outputs(6341) <= not b or a;
    layer1_outputs(6342) <= a and b;
    layer1_outputs(6343) <= not (a and b);
    layer1_outputs(6344) <= b and not a;
    layer1_outputs(6345) <= b and not a;
    layer1_outputs(6346) <= not b or a;
    layer1_outputs(6347) <= a and not b;
    layer1_outputs(6348) <= a or b;
    layer1_outputs(6349) <= not b or a;
    layer1_outputs(6350) <= not (a and b);
    layer1_outputs(6351) <= b and not a;
    layer1_outputs(6352) <= b;
    layer1_outputs(6353) <= a and b;
    layer1_outputs(6354) <= not (a or b);
    layer1_outputs(6355) <= not b;
    layer1_outputs(6356) <= '0';
    layer1_outputs(6357) <= a and b;
    layer1_outputs(6358) <= '0';
    layer1_outputs(6359) <= a and not b;
    layer1_outputs(6360) <= not (a and b);
    layer1_outputs(6361) <= '0';
    layer1_outputs(6362) <= not (a xor b);
    layer1_outputs(6363) <= '1';
    layer1_outputs(6364) <= not a;
    layer1_outputs(6365) <= a and not b;
    layer1_outputs(6366) <= not (a and b);
    layer1_outputs(6367) <= a or b;
    layer1_outputs(6368) <= not a or b;
    layer1_outputs(6369) <= a and b;
    layer1_outputs(6370) <= not (a and b);
    layer1_outputs(6371) <= a;
    layer1_outputs(6372) <= not b;
    layer1_outputs(6373) <= a and b;
    layer1_outputs(6374) <= b and not a;
    layer1_outputs(6375) <= '0';
    layer1_outputs(6376) <= b;
    layer1_outputs(6377) <= a and b;
    layer1_outputs(6378) <= not b;
    layer1_outputs(6379) <= not (a or b);
    layer1_outputs(6380) <= not (a or b);
    layer1_outputs(6381) <= '0';
    layer1_outputs(6382) <= '1';
    layer1_outputs(6383) <= not b or a;
    layer1_outputs(6384) <= a or b;
    layer1_outputs(6385) <= b;
    layer1_outputs(6386) <= not b or a;
    layer1_outputs(6387) <= b;
    layer1_outputs(6388) <= not b or a;
    layer1_outputs(6389) <= a and b;
    layer1_outputs(6390) <= not b or a;
    layer1_outputs(6391) <= not a;
    layer1_outputs(6392) <= a or b;
    layer1_outputs(6393) <= '1';
    layer1_outputs(6394) <= a and b;
    layer1_outputs(6395) <= not a or b;
    layer1_outputs(6396) <= not b or a;
    layer1_outputs(6397) <= not (a or b);
    layer1_outputs(6398) <= not (a and b);
    layer1_outputs(6399) <= '1';
    layer1_outputs(6400) <= not a or b;
    layer1_outputs(6401) <= a or b;
    layer1_outputs(6402) <= not b or a;
    layer1_outputs(6403) <= a and b;
    layer1_outputs(6404) <= a;
    layer1_outputs(6405) <= not (a xor b);
    layer1_outputs(6406) <= '0';
    layer1_outputs(6407) <= not b or a;
    layer1_outputs(6408) <= not (a and b);
    layer1_outputs(6409) <= a;
    layer1_outputs(6410) <= '1';
    layer1_outputs(6411) <= not (a or b);
    layer1_outputs(6412) <= '1';
    layer1_outputs(6413) <= not (a and b);
    layer1_outputs(6414) <= a xor b;
    layer1_outputs(6415) <= not a or b;
    layer1_outputs(6416) <= a or b;
    layer1_outputs(6417) <= not b;
    layer1_outputs(6418) <= b and not a;
    layer1_outputs(6419) <= not b or a;
    layer1_outputs(6420) <= '0';
    layer1_outputs(6421) <= '0';
    layer1_outputs(6422) <= a xor b;
    layer1_outputs(6423) <= a or b;
    layer1_outputs(6424) <= a xor b;
    layer1_outputs(6425) <= not b or a;
    layer1_outputs(6426) <= a and not b;
    layer1_outputs(6427) <= b and not a;
    layer1_outputs(6428) <= a and b;
    layer1_outputs(6429) <= not (a or b);
    layer1_outputs(6430) <= a and b;
    layer1_outputs(6431) <= not (a or b);
    layer1_outputs(6432) <= a and not b;
    layer1_outputs(6433) <= '1';
    layer1_outputs(6434) <= not a;
    layer1_outputs(6435) <= a or b;
    layer1_outputs(6436) <= not b or a;
    layer1_outputs(6437) <= not (a and b);
    layer1_outputs(6438) <= b and not a;
    layer1_outputs(6439) <= a and b;
    layer1_outputs(6440) <= a xor b;
    layer1_outputs(6441) <= '0';
    layer1_outputs(6442) <= a or b;
    layer1_outputs(6443) <= a;
    layer1_outputs(6444) <= a and not b;
    layer1_outputs(6445) <= b;
    layer1_outputs(6446) <= a or b;
    layer1_outputs(6447) <= a;
    layer1_outputs(6448) <= not (a or b);
    layer1_outputs(6449) <= a and b;
    layer1_outputs(6450) <= not b or a;
    layer1_outputs(6451) <= not (a xor b);
    layer1_outputs(6452) <= a and b;
    layer1_outputs(6453) <= b and not a;
    layer1_outputs(6454) <= a and not b;
    layer1_outputs(6455) <= a and b;
    layer1_outputs(6456) <= a xor b;
    layer1_outputs(6457) <= not a;
    layer1_outputs(6458) <= a or b;
    layer1_outputs(6459) <= not (a or b);
    layer1_outputs(6460) <= '0';
    layer1_outputs(6461) <= '1';
    layer1_outputs(6462) <= '1';
    layer1_outputs(6463) <= not b or a;
    layer1_outputs(6464) <= a and not b;
    layer1_outputs(6465) <= a and b;
    layer1_outputs(6466) <= not b;
    layer1_outputs(6467) <= a and b;
    layer1_outputs(6468) <= a and not b;
    layer1_outputs(6469) <= not b;
    layer1_outputs(6470) <= not a;
    layer1_outputs(6471) <= a;
    layer1_outputs(6472) <= '1';
    layer1_outputs(6473) <= not b or a;
    layer1_outputs(6474) <= a or b;
    layer1_outputs(6475) <= not b;
    layer1_outputs(6476) <= '1';
    layer1_outputs(6477) <= a or b;
    layer1_outputs(6478) <= '0';
    layer1_outputs(6479) <= b;
    layer1_outputs(6480) <= b and not a;
    layer1_outputs(6481) <= a and not b;
    layer1_outputs(6482) <= a and not b;
    layer1_outputs(6483) <= a and b;
    layer1_outputs(6484) <= '1';
    layer1_outputs(6485) <= '0';
    layer1_outputs(6486) <= not a;
    layer1_outputs(6487) <= a and not b;
    layer1_outputs(6488) <= b and not a;
    layer1_outputs(6489) <= not a;
    layer1_outputs(6490) <= not b or a;
    layer1_outputs(6491) <= not (a and b);
    layer1_outputs(6492) <= not b or a;
    layer1_outputs(6493) <= '1';
    layer1_outputs(6494) <= a or b;
    layer1_outputs(6495) <= not (a and b);
    layer1_outputs(6496) <= not a or b;
    layer1_outputs(6497) <= not b;
    layer1_outputs(6498) <= b and not a;
    layer1_outputs(6499) <= a or b;
    layer1_outputs(6500) <= a and b;
    layer1_outputs(6501) <= a;
    layer1_outputs(6502) <= b and not a;
    layer1_outputs(6503) <= a and not b;
    layer1_outputs(6504) <= not a;
    layer1_outputs(6505) <= a;
    layer1_outputs(6506) <= b and not a;
    layer1_outputs(6507) <= a xor b;
    layer1_outputs(6508) <= b and not a;
    layer1_outputs(6509) <= '0';
    layer1_outputs(6510) <= not (a and b);
    layer1_outputs(6511) <= not (a and b);
    layer1_outputs(6512) <= a;
    layer1_outputs(6513) <= a or b;
    layer1_outputs(6514) <= b;
    layer1_outputs(6515) <= a and b;
    layer1_outputs(6516) <= b;
    layer1_outputs(6517) <= not (a or b);
    layer1_outputs(6518) <= not b;
    layer1_outputs(6519) <= b;
    layer1_outputs(6520) <= not (a or b);
    layer1_outputs(6521) <= not b;
    layer1_outputs(6522) <= a or b;
    layer1_outputs(6523) <= not b;
    layer1_outputs(6524) <= '1';
    layer1_outputs(6525) <= b and not a;
    layer1_outputs(6526) <= not a;
    layer1_outputs(6527) <= b;
    layer1_outputs(6528) <= not a or b;
    layer1_outputs(6529) <= b;
    layer1_outputs(6530) <= not (a or b);
    layer1_outputs(6531) <= '0';
    layer1_outputs(6532) <= not a;
    layer1_outputs(6533) <= a and not b;
    layer1_outputs(6534) <= not a;
    layer1_outputs(6535) <= '1';
    layer1_outputs(6536) <= b and not a;
    layer1_outputs(6537) <= not (a and b);
    layer1_outputs(6538) <= b;
    layer1_outputs(6539) <= not a or b;
    layer1_outputs(6540) <= not (a and b);
    layer1_outputs(6541) <= a;
    layer1_outputs(6542) <= not (a and b);
    layer1_outputs(6543) <= a and not b;
    layer1_outputs(6544) <= not b or a;
    layer1_outputs(6545) <= '1';
    layer1_outputs(6546) <= not b or a;
    layer1_outputs(6547) <= a or b;
    layer1_outputs(6548) <= '1';
    layer1_outputs(6549) <= not a or b;
    layer1_outputs(6550) <= not b or a;
    layer1_outputs(6551) <= not b;
    layer1_outputs(6552) <= a and not b;
    layer1_outputs(6553) <= a and b;
    layer1_outputs(6554) <= not a or b;
    layer1_outputs(6555) <= not b or a;
    layer1_outputs(6556) <= not b or a;
    layer1_outputs(6557) <= not b or a;
    layer1_outputs(6558) <= '1';
    layer1_outputs(6559) <= a and not b;
    layer1_outputs(6560) <= '1';
    layer1_outputs(6561) <= a or b;
    layer1_outputs(6562) <= a;
    layer1_outputs(6563) <= '1';
    layer1_outputs(6564) <= not (a and b);
    layer1_outputs(6565) <= '1';
    layer1_outputs(6566) <= a and b;
    layer1_outputs(6567) <= not a or b;
    layer1_outputs(6568) <= not a or b;
    layer1_outputs(6569) <= b;
    layer1_outputs(6570) <= b;
    layer1_outputs(6571) <= a;
    layer1_outputs(6572) <= not a or b;
    layer1_outputs(6573) <= a and not b;
    layer1_outputs(6574) <= not b;
    layer1_outputs(6575) <= b;
    layer1_outputs(6576) <= not (a or b);
    layer1_outputs(6577) <= not (a and b);
    layer1_outputs(6578) <= '1';
    layer1_outputs(6579) <= not b;
    layer1_outputs(6580) <= a or b;
    layer1_outputs(6581) <= '0';
    layer1_outputs(6582) <= not (a or b);
    layer1_outputs(6583) <= not a or b;
    layer1_outputs(6584) <= not (a and b);
    layer1_outputs(6585) <= '0';
    layer1_outputs(6586) <= a;
    layer1_outputs(6587) <= a and b;
    layer1_outputs(6588) <= a xor b;
    layer1_outputs(6589) <= b and not a;
    layer1_outputs(6590) <= not a or b;
    layer1_outputs(6591) <= a or b;
    layer1_outputs(6592) <= b;
    layer1_outputs(6593) <= not b;
    layer1_outputs(6594) <= not a or b;
    layer1_outputs(6595) <= '1';
    layer1_outputs(6596) <= a and not b;
    layer1_outputs(6597) <= not (a or b);
    layer1_outputs(6598) <= b and not a;
    layer1_outputs(6599) <= not a or b;
    layer1_outputs(6600) <= b and not a;
    layer1_outputs(6601) <= '1';
    layer1_outputs(6602) <= a and b;
    layer1_outputs(6603) <= b and not a;
    layer1_outputs(6604) <= a xor b;
    layer1_outputs(6605) <= not (a and b);
    layer1_outputs(6606) <= b;
    layer1_outputs(6607) <= '0';
    layer1_outputs(6608) <= not (a and b);
    layer1_outputs(6609) <= not (a and b);
    layer1_outputs(6610) <= not a;
    layer1_outputs(6611) <= a;
    layer1_outputs(6612) <= not (a or b);
    layer1_outputs(6613) <= b;
    layer1_outputs(6614) <= not b or a;
    layer1_outputs(6615) <= '1';
    layer1_outputs(6616) <= a xor b;
    layer1_outputs(6617) <= a and not b;
    layer1_outputs(6618) <= a and b;
    layer1_outputs(6619) <= '0';
    layer1_outputs(6620) <= a xor b;
    layer1_outputs(6621) <= a;
    layer1_outputs(6622) <= not b;
    layer1_outputs(6623) <= not a or b;
    layer1_outputs(6624) <= not (a and b);
    layer1_outputs(6625) <= not a or b;
    layer1_outputs(6626) <= b;
    layer1_outputs(6627) <= a;
    layer1_outputs(6628) <= not (a and b);
    layer1_outputs(6629) <= not (a and b);
    layer1_outputs(6630) <= not (a and b);
    layer1_outputs(6631) <= b and not a;
    layer1_outputs(6632) <= not b;
    layer1_outputs(6633) <= not b;
    layer1_outputs(6634) <= not b or a;
    layer1_outputs(6635) <= not (a and b);
    layer1_outputs(6636) <= a and b;
    layer1_outputs(6637) <= b and not a;
    layer1_outputs(6638) <= not a;
    layer1_outputs(6639) <= not a or b;
    layer1_outputs(6640) <= '1';
    layer1_outputs(6641) <= not b or a;
    layer1_outputs(6642) <= not a;
    layer1_outputs(6643) <= not b or a;
    layer1_outputs(6644) <= not b or a;
    layer1_outputs(6645) <= a and not b;
    layer1_outputs(6646) <= a;
    layer1_outputs(6647) <= a or b;
    layer1_outputs(6648) <= a and not b;
    layer1_outputs(6649) <= a or b;
    layer1_outputs(6650) <= not (a and b);
    layer1_outputs(6651) <= '0';
    layer1_outputs(6652) <= a and b;
    layer1_outputs(6653) <= a xor b;
    layer1_outputs(6654) <= '1';
    layer1_outputs(6655) <= b;
    layer1_outputs(6656) <= not b or a;
    layer1_outputs(6657) <= not b or a;
    layer1_outputs(6658) <= '0';
    layer1_outputs(6659) <= a and b;
    layer1_outputs(6660) <= '0';
    layer1_outputs(6661) <= '0';
    layer1_outputs(6662) <= a xor b;
    layer1_outputs(6663) <= '0';
    layer1_outputs(6664) <= b and not a;
    layer1_outputs(6665) <= '1';
    layer1_outputs(6666) <= not a or b;
    layer1_outputs(6667) <= '0';
    layer1_outputs(6668) <= not a;
    layer1_outputs(6669) <= not a or b;
    layer1_outputs(6670) <= not b;
    layer1_outputs(6671) <= not (a or b);
    layer1_outputs(6672) <= a and not b;
    layer1_outputs(6673) <= not b or a;
    layer1_outputs(6674) <= a and not b;
    layer1_outputs(6675) <= b;
    layer1_outputs(6676) <= b and not a;
    layer1_outputs(6677) <= b;
    layer1_outputs(6678) <= '0';
    layer1_outputs(6679) <= not b or a;
    layer1_outputs(6680) <= a and not b;
    layer1_outputs(6681) <= a or b;
    layer1_outputs(6682) <= not a or b;
    layer1_outputs(6683) <= not b;
    layer1_outputs(6684) <= not a;
    layer1_outputs(6685) <= '1';
    layer1_outputs(6686) <= '1';
    layer1_outputs(6687) <= not a or b;
    layer1_outputs(6688) <= not b;
    layer1_outputs(6689) <= b;
    layer1_outputs(6690) <= a or b;
    layer1_outputs(6691) <= a and not b;
    layer1_outputs(6692) <= a or b;
    layer1_outputs(6693) <= '0';
    layer1_outputs(6694) <= not (a and b);
    layer1_outputs(6695) <= a and b;
    layer1_outputs(6696) <= '1';
    layer1_outputs(6697) <= not a or b;
    layer1_outputs(6698) <= b and not a;
    layer1_outputs(6699) <= not b;
    layer1_outputs(6700) <= a or b;
    layer1_outputs(6701) <= '1';
    layer1_outputs(6702) <= not b or a;
    layer1_outputs(6703) <= b and not a;
    layer1_outputs(6704) <= a and not b;
    layer1_outputs(6705) <= not (a or b);
    layer1_outputs(6706) <= not a or b;
    layer1_outputs(6707) <= a or b;
    layer1_outputs(6708) <= '1';
    layer1_outputs(6709) <= a xor b;
    layer1_outputs(6710) <= b and not a;
    layer1_outputs(6711) <= a or b;
    layer1_outputs(6712) <= b and not a;
    layer1_outputs(6713) <= '1';
    layer1_outputs(6714) <= not b;
    layer1_outputs(6715) <= a and not b;
    layer1_outputs(6716) <= b and not a;
    layer1_outputs(6717) <= not a or b;
    layer1_outputs(6718) <= '0';
    layer1_outputs(6719) <= a and not b;
    layer1_outputs(6720) <= not b;
    layer1_outputs(6721) <= not b;
    layer1_outputs(6722) <= not b;
    layer1_outputs(6723) <= '1';
    layer1_outputs(6724) <= not a or b;
    layer1_outputs(6725) <= not a;
    layer1_outputs(6726) <= not b or a;
    layer1_outputs(6727) <= not b;
    layer1_outputs(6728) <= a;
    layer1_outputs(6729) <= not a or b;
    layer1_outputs(6730) <= not b;
    layer1_outputs(6731) <= b;
    layer1_outputs(6732) <= '0';
    layer1_outputs(6733) <= a and b;
    layer1_outputs(6734) <= not a;
    layer1_outputs(6735) <= not a;
    layer1_outputs(6736) <= '1';
    layer1_outputs(6737) <= not b or a;
    layer1_outputs(6738) <= a and not b;
    layer1_outputs(6739) <= a and not b;
    layer1_outputs(6740) <= a and not b;
    layer1_outputs(6741) <= not a;
    layer1_outputs(6742) <= not (a xor b);
    layer1_outputs(6743) <= '1';
    layer1_outputs(6744) <= b;
    layer1_outputs(6745) <= not (a or b);
    layer1_outputs(6746) <= '1';
    layer1_outputs(6747) <= b;
    layer1_outputs(6748) <= a and not b;
    layer1_outputs(6749) <= '0';
    layer1_outputs(6750) <= b;
    layer1_outputs(6751) <= b;
    layer1_outputs(6752) <= a and not b;
    layer1_outputs(6753) <= a;
    layer1_outputs(6754) <= b and not a;
    layer1_outputs(6755) <= not (a and b);
    layer1_outputs(6756) <= not (a xor b);
    layer1_outputs(6757) <= a and b;
    layer1_outputs(6758) <= a and b;
    layer1_outputs(6759) <= not (a or b);
    layer1_outputs(6760) <= not a;
    layer1_outputs(6761) <= b;
    layer1_outputs(6762) <= a or b;
    layer1_outputs(6763) <= b;
    layer1_outputs(6764) <= a and not b;
    layer1_outputs(6765) <= not a or b;
    layer1_outputs(6766) <= not b;
    layer1_outputs(6767) <= not b;
    layer1_outputs(6768) <= a;
    layer1_outputs(6769) <= a and b;
    layer1_outputs(6770) <= a and b;
    layer1_outputs(6771) <= a or b;
    layer1_outputs(6772) <= '1';
    layer1_outputs(6773) <= b;
    layer1_outputs(6774) <= a;
    layer1_outputs(6775) <= b;
    layer1_outputs(6776) <= a;
    layer1_outputs(6777) <= a and b;
    layer1_outputs(6778) <= '0';
    layer1_outputs(6779) <= b;
    layer1_outputs(6780) <= '1';
    layer1_outputs(6781) <= b;
    layer1_outputs(6782) <= a;
    layer1_outputs(6783) <= '0';
    layer1_outputs(6784) <= '0';
    layer1_outputs(6785) <= not a or b;
    layer1_outputs(6786) <= not b;
    layer1_outputs(6787) <= not a;
    layer1_outputs(6788) <= '1';
    layer1_outputs(6789) <= a;
    layer1_outputs(6790) <= a and b;
    layer1_outputs(6791) <= not b;
    layer1_outputs(6792) <= a xor b;
    layer1_outputs(6793) <= b;
    layer1_outputs(6794) <= a xor b;
    layer1_outputs(6795) <= not (a or b);
    layer1_outputs(6796) <= a;
    layer1_outputs(6797) <= not (a and b);
    layer1_outputs(6798) <= '0';
    layer1_outputs(6799) <= a and not b;
    layer1_outputs(6800) <= a and b;
    layer1_outputs(6801) <= not (a or b);
    layer1_outputs(6802) <= not a;
    layer1_outputs(6803) <= b and not a;
    layer1_outputs(6804) <= a and not b;
    layer1_outputs(6805) <= a or b;
    layer1_outputs(6806) <= a;
    layer1_outputs(6807) <= a or b;
    layer1_outputs(6808) <= not a or b;
    layer1_outputs(6809) <= not a or b;
    layer1_outputs(6810) <= '1';
    layer1_outputs(6811) <= not b;
    layer1_outputs(6812) <= not a or b;
    layer1_outputs(6813) <= '1';
    layer1_outputs(6814) <= not b;
    layer1_outputs(6815) <= a or b;
    layer1_outputs(6816) <= b and not a;
    layer1_outputs(6817) <= a or b;
    layer1_outputs(6818) <= not (a or b);
    layer1_outputs(6819) <= not a;
    layer1_outputs(6820) <= not (a and b);
    layer1_outputs(6821) <= not a or b;
    layer1_outputs(6822) <= a and b;
    layer1_outputs(6823) <= '1';
    layer1_outputs(6824) <= '1';
    layer1_outputs(6825) <= '0';
    layer1_outputs(6826) <= a or b;
    layer1_outputs(6827) <= not a or b;
    layer1_outputs(6828) <= a or b;
    layer1_outputs(6829) <= '0';
    layer1_outputs(6830) <= a and not b;
    layer1_outputs(6831) <= a;
    layer1_outputs(6832) <= not a or b;
    layer1_outputs(6833) <= '1';
    layer1_outputs(6834) <= '0';
    layer1_outputs(6835) <= b and not a;
    layer1_outputs(6836) <= not (a or b);
    layer1_outputs(6837) <= not (a and b);
    layer1_outputs(6838) <= not (a or b);
    layer1_outputs(6839) <= a;
    layer1_outputs(6840) <= a and b;
    layer1_outputs(6841) <= not (a and b);
    layer1_outputs(6842) <= not b;
    layer1_outputs(6843) <= not a or b;
    layer1_outputs(6844) <= b and not a;
    layer1_outputs(6845) <= b;
    layer1_outputs(6846) <= '0';
    layer1_outputs(6847) <= not a;
    layer1_outputs(6848) <= b;
    layer1_outputs(6849) <= a and b;
    layer1_outputs(6850) <= not (a and b);
    layer1_outputs(6851) <= a and b;
    layer1_outputs(6852) <= a and b;
    layer1_outputs(6853) <= b and not a;
    layer1_outputs(6854) <= a and b;
    layer1_outputs(6855) <= '0';
    layer1_outputs(6856) <= '0';
    layer1_outputs(6857) <= a;
    layer1_outputs(6858) <= not b or a;
    layer1_outputs(6859) <= not (a and b);
    layer1_outputs(6860) <= not (a and b);
    layer1_outputs(6861) <= a and not b;
    layer1_outputs(6862) <= not (a or b);
    layer1_outputs(6863) <= not (a or b);
    layer1_outputs(6864) <= not a;
    layer1_outputs(6865) <= a xor b;
    layer1_outputs(6866) <= not b or a;
    layer1_outputs(6867) <= a xor b;
    layer1_outputs(6868) <= not b;
    layer1_outputs(6869) <= not a or b;
    layer1_outputs(6870) <= not (a and b);
    layer1_outputs(6871) <= not b or a;
    layer1_outputs(6872) <= b and not a;
    layer1_outputs(6873) <= a or b;
    layer1_outputs(6874) <= a and b;
    layer1_outputs(6875) <= '1';
    layer1_outputs(6876) <= a and not b;
    layer1_outputs(6877) <= not b;
    layer1_outputs(6878) <= b and not a;
    layer1_outputs(6879) <= b and not a;
    layer1_outputs(6880) <= a;
    layer1_outputs(6881) <= '0';
    layer1_outputs(6882) <= a or b;
    layer1_outputs(6883) <= not b;
    layer1_outputs(6884) <= a;
    layer1_outputs(6885) <= a or b;
    layer1_outputs(6886) <= not a or b;
    layer1_outputs(6887) <= not a;
    layer1_outputs(6888) <= not (a or b);
    layer1_outputs(6889) <= a and b;
    layer1_outputs(6890) <= not a;
    layer1_outputs(6891) <= '0';
    layer1_outputs(6892) <= b;
    layer1_outputs(6893) <= a;
    layer1_outputs(6894) <= not a;
    layer1_outputs(6895) <= a and not b;
    layer1_outputs(6896) <= not a;
    layer1_outputs(6897) <= '1';
    layer1_outputs(6898) <= b;
    layer1_outputs(6899) <= a and not b;
    layer1_outputs(6900) <= not (a and b);
    layer1_outputs(6901) <= '1';
    layer1_outputs(6902) <= a and not b;
    layer1_outputs(6903) <= b;
    layer1_outputs(6904) <= a;
    layer1_outputs(6905) <= a and b;
    layer1_outputs(6906) <= not a or b;
    layer1_outputs(6907) <= a and not b;
    layer1_outputs(6908) <= a and b;
    layer1_outputs(6909) <= '0';
    layer1_outputs(6910) <= a;
    layer1_outputs(6911) <= not (a or b);
    layer1_outputs(6912) <= '0';
    layer1_outputs(6913) <= a and not b;
    layer1_outputs(6914) <= b;
    layer1_outputs(6915) <= a and not b;
    layer1_outputs(6916) <= not (a and b);
    layer1_outputs(6917) <= '1';
    layer1_outputs(6918) <= a or b;
    layer1_outputs(6919) <= a and not b;
    layer1_outputs(6920) <= a;
    layer1_outputs(6921) <= not b or a;
    layer1_outputs(6922) <= a;
    layer1_outputs(6923) <= not a;
    layer1_outputs(6924) <= b;
    layer1_outputs(6925) <= not b or a;
    layer1_outputs(6926) <= '0';
    layer1_outputs(6927) <= not b or a;
    layer1_outputs(6928) <= not (a or b);
    layer1_outputs(6929) <= not (a or b);
    layer1_outputs(6930) <= b and not a;
    layer1_outputs(6931) <= not a;
    layer1_outputs(6932) <= not (a or b);
    layer1_outputs(6933) <= '0';
    layer1_outputs(6934) <= not b or a;
    layer1_outputs(6935) <= a and not b;
    layer1_outputs(6936) <= '1';
    layer1_outputs(6937) <= not (a or b);
    layer1_outputs(6938) <= a;
    layer1_outputs(6939) <= '0';
    layer1_outputs(6940) <= '1';
    layer1_outputs(6941) <= '1';
    layer1_outputs(6942) <= '0';
    layer1_outputs(6943) <= '1';
    layer1_outputs(6944) <= b;
    layer1_outputs(6945) <= '0';
    layer1_outputs(6946) <= '1';
    layer1_outputs(6947) <= a xor b;
    layer1_outputs(6948) <= not (a and b);
    layer1_outputs(6949) <= b;
    layer1_outputs(6950) <= a and not b;
    layer1_outputs(6951) <= '0';
    layer1_outputs(6952) <= not b or a;
    layer1_outputs(6953) <= b;
    layer1_outputs(6954) <= b;
    layer1_outputs(6955) <= a xor b;
    layer1_outputs(6956) <= a and b;
    layer1_outputs(6957) <= b and not a;
    layer1_outputs(6958) <= '0';
    layer1_outputs(6959) <= a xor b;
    layer1_outputs(6960) <= a and not b;
    layer1_outputs(6961) <= a and b;
    layer1_outputs(6962) <= not a or b;
    layer1_outputs(6963) <= not a;
    layer1_outputs(6964) <= '0';
    layer1_outputs(6965) <= not (a xor b);
    layer1_outputs(6966) <= not b or a;
    layer1_outputs(6967) <= '1';
    layer1_outputs(6968) <= not a or b;
    layer1_outputs(6969) <= '1';
    layer1_outputs(6970) <= not b;
    layer1_outputs(6971) <= '0';
    layer1_outputs(6972) <= a;
    layer1_outputs(6973) <= not (a or b);
    layer1_outputs(6974) <= not b;
    layer1_outputs(6975) <= not (a or b);
    layer1_outputs(6976) <= '1';
    layer1_outputs(6977) <= b and not a;
    layer1_outputs(6978) <= not a;
    layer1_outputs(6979) <= not b;
    layer1_outputs(6980) <= '0';
    layer1_outputs(6981) <= not (a or b);
    layer1_outputs(6982) <= not b or a;
    layer1_outputs(6983) <= b;
    layer1_outputs(6984) <= a and b;
    layer1_outputs(6985) <= not b or a;
    layer1_outputs(6986) <= '0';
    layer1_outputs(6987) <= not a;
    layer1_outputs(6988) <= a;
    layer1_outputs(6989) <= '1';
    layer1_outputs(6990) <= not (a and b);
    layer1_outputs(6991) <= not (a and b);
    layer1_outputs(6992) <= not b or a;
    layer1_outputs(6993) <= b and not a;
    layer1_outputs(6994) <= not (a or b);
    layer1_outputs(6995) <= not b;
    layer1_outputs(6996) <= not a;
    layer1_outputs(6997) <= '1';
    layer1_outputs(6998) <= '0';
    layer1_outputs(6999) <= a;
    layer1_outputs(7000) <= a;
    layer1_outputs(7001) <= a or b;
    layer1_outputs(7002) <= '0';
    layer1_outputs(7003) <= a;
    layer1_outputs(7004) <= not b or a;
    layer1_outputs(7005) <= not b;
    layer1_outputs(7006) <= '0';
    layer1_outputs(7007) <= a and b;
    layer1_outputs(7008) <= b and not a;
    layer1_outputs(7009) <= a;
    layer1_outputs(7010) <= a and b;
    layer1_outputs(7011) <= not a;
    layer1_outputs(7012) <= not b;
    layer1_outputs(7013) <= '1';
    layer1_outputs(7014) <= b and not a;
    layer1_outputs(7015) <= not (a and b);
    layer1_outputs(7016) <= not a or b;
    layer1_outputs(7017) <= b and not a;
    layer1_outputs(7018) <= not (a xor b);
    layer1_outputs(7019) <= '1';
    layer1_outputs(7020) <= '0';
    layer1_outputs(7021) <= a or b;
    layer1_outputs(7022) <= not (a and b);
    layer1_outputs(7023) <= a;
    layer1_outputs(7024) <= a and not b;
    layer1_outputs(7025) <= b and not a;
    layer1_outputs(7026) <= not b;
    layer1_outputs(7027) <= not a;
    layer1_outputs(7028) <= '0';
    layer1_outputs(7029) <= '1';
    layer1_outputs(7030) <= not b or a;
    layer1_outputs(7031) <= a and b;
    layer1_outputs(7032) <= not a or b;
    layer1_outputs(7033) <= not a or b;
    layer1_outputs(7034) <= '1';
    layer1_outputs(7035) <= not (a or b);
    layer1_outputs(7036) <= '1';
    layer1_outputs(7037) <= a and not b;
    layer1_outputs(7038) <= a or b;
    layer1_outputs(7039) <= not b;
    layer1_outputs(7040) <= b and not a;
    layer1_outputs(7041) <= b and not a;
    layer1_outputs(7042) <= '1';
    layer1_outputs(7043) <= '1';
    layer1_outputs(7044) <= b and not a;
    layer1_outputs(7045) <= not b;
    layer1_outputs(7046) <= not b or a;
    layer1_outputs(7047) <= a;
    layer1_outputs(7048) <= a and b;
    layer1_outputs(7049) <= not b or a;
    layer1_outputs(7050) <= not (a or b);
    layer1_outputs(7051) <= a and b;
    layer1_outputs(7052) <= not b or a;
    layer1_outputs(7053) <= a xor b;
    layer1_outputs(7054) <= not a or b;
    layer1_outputs(7055) <= not (a or b);
    layer1_outputs(7056) <= not a;
    layer1_outputs(7057) <= a;
    layer1_outputs(7058) <= b;
    layer1_outputs(7059) <= '0';
    layer1_outputs(7060) <= not a;
    layer1_outputs(7061) <= not (a or b);
    layer1_outputs(7062) <= not (a and b);
    layer1_outputs(7063) <= not a or b;
    layer1_outputs(7064) <= not (a or b);
    layer1_outputs(7065) <= '1';
    layer1_outputs(7066) <= not (a or b);
    layer1_outputs(7067) <= not (a or b);
    layer1_outputs(7068) <= a;
    layer1_outputs(7069) <= not (a xor b);
    layer1_outputs(7070) <= a or b;
    layer1_outputs(7071) <= not (a or b);
    layer1_outputs(7072) <= a or b;
    layer1_outputs(7073) <= a;
    layer1_outputs(7074) <= a and b;
    layer1_outputs(7075) <= a and not b;
    layer1_outputs(7076) <= not (a or b);
    layer1_outputs(7077) <= not (a and b);
    layer1_outputs(7078) <= b;
    layer1_outputs(7079) <= not a;
    layer1_outputs(7080) <= not a or b;
    layer1_outputs(7081) <= a xor b;
    layer1_outputs(7082) <= b;
    layer1_outputs(7083) <= a;
    layer1_outputs(7084) <= not a;
    layer1_outputs(7085) <= b;
    layer1_outputs(7086) <= not b;
    layer1_outputs(7087) <= '0';
    layer1_outputs(7088) <= not (a and b);
    layer1_outputs(7089) <= b and not a;
    layer1_outputs(7090) <= '0';
    layer1_outputs(7091) <= b;
    layer1_outputs(7092) <= a or b;
    layer1_outputs(7093) <= not a or b;
    layer1_outputs(7094) <= a;
    layer1_outputs(7095) <= not b;
    layer1_outputs(7096) <= not b;
    layer1_outputs(7097) <= b and not a;
    layer1_outputs(7098) <= not b or a;
    layer1_outputs(7099) <= a;
    layer1_outputs(7100) <= not a or b;
    layer1_outputs(7101) <= not (a xor b);
    layer1_outputs(7102) <= a or b;
    layer1_outputs(7103) <= b;
    layer1_outputs(7104) <= b and not a;
    layer1_outputs(7105) <= not a;
    layer1_outputs(7106) <= b and not a;
    layer1_outputs(7107) <= '1';
    layer1_outputs(7108) <= '1';
    layer1_outputs(7109) <= not (a or b);
    layer1_outputs(7110) <= not (a xor b);
    layer1_outputs(7111) <= not b or a;
    layer1_outputs(7112) <= a and b;
    layer1_outputs(7113) <= not b;
    layer1_outputs(7114) <= '0';
    layer1_outputs(7115) <= not (a xor b);
    layer1_outputs(7116) <= not b or a;
    layer1_outputs(7117) <= not b or a;
    layer1_outputs(7118) <= b;
    layer1_outputs(7119) <= not (a or b);
    layer1_outputs(7120) <= a or b;
    layer1_outputs(7121) <= '1';
    layer1_outputs(7122) <= not (a or b);
    layer1_outputs(7123) <= a or b;
    layer1_outputs(7124) <= '0';
    layer1_outputs(7125) <= not a or b;
    layer1_outputs(7126) <= a and not b;
    layer1_outputs(7127) <= not (a and b);
    layer1_outputs(7128) <= a;
    layer1_outputs(7129) <= a xor b;
    layer1_outputs(7130) <= not a or b;
    layer1_outputs(7131) <= not a or b;
    layer1_outputs(7132) <= b and not a;
    layer1_outputs(7133) <= '1';
    layer1_outputs(7134) <= a xor b;
    layer1_outputs(7135) <= '1';
    layer1_outputs(7136) <= a and b;
    layer1_outputs(7137) <= a or b;
    layer1_outputs(7138) <= not (a and b);
    layer1_outputs(7139) <= not b or a;
    layer1_outputs(7140) <= b;
    layer1_outputs(7141) <= '0';
    layer1_outputs(7142) <= '0';
    layer1_outputs(7143) <= a and b;
    layer1_outputs(7144) <= not a or b;
    layer1_outputs(7145) <= '0';
    layer1_outputs(7146) <= not a;
    layer1_outputs(7147) <= not b or a;
    layer1_outputs(7148) <= not (a or b);
    layer1_outputs(7149) <= a or b;
    layer1_outputs(7150) <= not a or b;
    layer1_outputs(7151) <= not a;
    layer1_outputs(7152) <= '0';
    layer1_outputs(7153) <= not (a and b);
    layer1_outputs(7154) <= not b or a;
    layer1_outputs(7155) <= a and not b;
    layer1_outputs(7156) <= not (a xor b);
    layer1_outputs(7157) <= not (a xor b);
    layer1_outputs(7158) <= a;
    layer1_outputs(7159) <= not (a or b);
    layer1_outputs(7160) <= a or b;
    layer1_outputs(7161) <= not b;
    layer1_outputs(7162) <= b;
    layer1_outputs(7163) <= a;
    layer1_outputs(7164) <= '1';
    layer1_outputs(7165) <= not b or a;
    layer1_outputs(7166) <= a xor b;
    layer1_outputs(7167) <= not b;
    layer1_outputs(7168) <= a and b;
    layer1_outputs(7169) <= not b or a;
    layer1_outputs(7170) <= '1';
    layer1_outputs(7171) <= a and not b;
    layer1_outputs(7172) <= '1';
    layer1_outputs(7173) <= b and not a;
    layer1_outputs(7174) <= a or b;
    layer1_outputs(7175) <= not b or a;
    layer1_outputs(7176) <= a or b;
    layer1_outputs(7177) <= a and b;
    layer1_outputs(7178) <= not (a xor b);
    layer1_outputs(7179) <= not b;
    layer1_outputs(7180) <= '1';
    layer1_outputs(7181) <= '1';
    layer1_outputs(7182) <= not (a or b);
    layer1_outputs(7183) <= b and not a;
    layer1_outputs(7184) <= b;
    layer1_outputs(7185) <= b;
    layer1_outputs(7186) <= '1';
    layer1_outputs(7187) <= a or b;
    layer1_outputs(7188) <= not a or b;
    layer1_outputs(7189) <= '1';
    layer1_outputs(7190) <= not b;
    layer1_outputs(7191) <= a and b;
    layer1_outputs(7192) <= '0';
    layer1_outputs(7193) <= b and not a;
    layer1_outputs(7194) <= not (a or b);
    layer1_outputs(7195) <= a or b;
    layer1_outputs(7196) <= '1';
    layer1_outputs(7197) <= a and not b;
    layer1_outputs(7198) <= not a or b;
    layer1_outputs(7199) <= not a or b;
    layer1_outputs(7200) <= b and not a;
    layer1_outputs(7201) <= not (a xor b);
    layer1_outputs(7202) <= '0';
    layer1_outputs(7203) <= not (a or b);
    layer1_outputs(7204) <= a and not b;
    layer1_outputs(7205) <= '1';
    layer1_outputs(7206) <= b and not a;
    layer1_outputs(7207) <= not b;
    layer1_outputs(7208) <= a or b;
    layer1_outputs(7209) <= not (a and b);
    layer1_outputs(7210) <= a and b;
    layer1_outputs(7211) <= a and not b;
    layer1_outputs(7212) <= b and not a;
    layer1_outputs(7213) <= a;
    layer1_outputs(7214) <= '0';
    layer1_outputs(7215) <= a or b;
    layer1_outputs(7216) <= b and not a;
    layer1_outputs(7217) <= '1';
    layer1_outputs(7218) <= '1';
    layer1_outputs(7219) <= b and not a;
    layer1_outputs(7220) <= not a or b;
    layer1_outputs(7221) <= not b;
    layer1_outputs(7222) <= '0';
    layer1_outputs(7223) <= not a or b;
    layer1_outputs(7224) <= not a or b;
    layer1_outputs(7225) <= '1';
    layer1_outputs(7226) <= a;
    layer1_outputs(7227) <= not b;
    layer1_outputs(7228) <= not a or b;
    layer1_outputs(7229) <= a or b;
    layer1_outputs(7230) <= b;
    layer1_outputs(7231) <= not b or a;
    layer1_outputs(7232) <= b;
    layer1_outputs(7233) <= not b;
    layer1_outputs(7234) <= not (a or b);
    layer1_outputs(7235) <= not (a and b);
    layer1_outputs(7236) <= not a;
    layer1_outputs(7237) <= a and b;
    layer1_outputs(7238) <= '1';
    layer1_outputs(7239) <= a;
    layer1_outputs(7240) <= not (a or b);
    layer1_outputs(7241) <= a;
    layer1_outputs(7242) <= '1';
    layer1_outputs(7243) <= not (a or b);
    layer1_outputs(7244) <= '0';
    layer1_outputs(7245) <= a or b;
    layer1_outputs(7246) <= b;
    layer1_outputs(7247) <= a and b;
    layer1_outputs(7248) <= b and not a;
    layer1_outputs(7249) <= not (a xor b);
    layer1_outputs(7250) <= not (a xor b);
    layer1_outputs(7251) <= not b or a;
    layer1_outputs(7252) <= a and b;
    layer1_outputs(7253) <= b and not a;
    layer1_outputs(7254) <= not a or b;
    layer1_outputs(7255) <= a and not b;
    layer1_outputs(7256) <= not b or a;
    layer1_outputs(7257) <= a or b;
    layer1_outputs(7258) <= a;
    layer1_outputs(7259) <= b;
    layer1_outputs(7260) <= '1';
    layer1_outputs(7261) <= b and not a;
    layer1_outputs(7262) <= not a or b;
    layer1_outputs(7263) <= a and b;
    layer1_outputs(7264) <= not b;
    layer1_outputs(7265) <= '0';
    layer1_outputs(7266) <= b and not a;
    layer1_outputs(7267) <= not (a or b);
    layer1_outputs(7268) <= not (a and b);
    layer1_outputs(7269) <= not b or a;
    layer1_outputs(7270) <= not b;
    layer1_outputs(7271) <= '0';
    layer1_outputs(7272) <= '1';
    layer1_outputs(7273) <= not a;
    layer1_outputs(7274) <= not a;
    layer1_outputs(7275) <= b;
    layer1_outputs(7276) <= '1';
    layer1_outputs(7277) <= b;
    layer1_outputs(7278) <= not (a xor b);
    layer1_outputs(7279) <= not (a or b);
    layer1_outputs(7280) <= not (a and b);
    layer1_outputs(7281) <= a and not b;
    layer1_outputs(7282) <= not b;
    layer1_outputs(7283) <= a and not b;
    layer1_outputs(7284) <= not b;
    layer1_outputs(7285) <= b and not a;
    layer1_outputs(7286) <= '1';
    layer1_outputs(7287) <= not (a and b);
    layer1_outputs(7288) <= a and b;
    layer1_outputs(7289) <= '0';
    layer1_outputs(7290) <= b;
    layer1_outputs(7291) <= not (a or b);
    layer1_outputs(7292) <= not a;
    layer1_outputs(7293) <= not b or a;
    layer1_outputs(7294) <= '0';
    layer1_outputs(7295) <= not (a and b);
    layer1_outputs(7296) <= b;
    layer1_outputs(7297) <= not b or a;
    layer1_outputs(7298) <= a and b;
    layer1_outputs(7299) <= not a;
    layer1_outputs(7300) <= a;
    layer1_outputs(7301) <= a and not b;
    layer1_outputs(7302) <= a or b;
    layer1_outputs(7303) <= a;
    layer1_outputs(7304) <= not (a or b);
    layer1_outputs(7305) <= b and not a;
    layer1_outputs(7306) <= a and not b;
    layer1_outputs(7307) <= not b or a;
    layer1_outputs(7308) <= a xor b;
    layer1_outputs(7309) <= b;
    layer1_outputs(7310) <= b;
    layer1_outputs(7311) <= a;
    layer1_outputs(7312) <= a;
    layer1_outputs(7313) <= a;
    layer1_outputs(7314) <= not a or b;
    layer1_outputs(7315) <= not b or a;
    layer1_outputs(7316) <= a or b;
    layer1_outputs(7317) <= not a;
    layer1_outputs(7318) <= '0';
    layer1_outputs(7319) <= not (a xor b);
    layer1_outputs(7320) <= not (a and b);
    layer1_outputs(7321) <= not a or b;
    layer1_outputs(7322) <= not a or b;
    layer1_outputs(7323) <= a;
    layer1_outputs(7324) <= b;
    layer1_outputs(7325) <= not b;
    layer1_outputs(7326) <= not b;
    layer1_outputs(7327) <= '0';
    layer1_outputs(7328) <= not (a xor b);
    layer1_outputs(7329) <= not b or a;
    layer1_outputs(7330) <= not (a and b);
    layer1_outputs(7331) <= not a;
    layer1_outputs(7332) <= a or b;
    layer1_outputs(7333) <= not b;
    layer1_outputs(7334) <= not (a or b);
    layer1_outputs(7335) <= a;
    layer1_outputs(7336) <= a;
    layer1_outputs(7337) <= a and not b;
    layer1_outputs(7338) <= a or b;
    layer1_outputs(7339) <= a and b;
    layer1_outputs(7340) <= b;
    layer1_outputs(7341) <= '0';
    layer1_outputs(7342) <= b;
    layer1_outputs(7343) <= '1';
    layer1_outputs(7344) <= a and not b;
    layer1_outputs(7345) <= b and not a;
    layer1_outputs(7346) <= '0';
    layer1_outputs(7347) <= not (a or b);
    layer1_outputs(7348) <= b;
    layer1_outputs(7349) <= '1';
    layer1_outputs(7350) <= '1';
    layer1_outputs(7351) <= a and not b;
    layer1_outputs(7352) <= not b or a;
    layer1_outputs(7353) <= '0';
    layer1_outputs(7354) <= not (a and b);
    layer1_outputs(7355) <= '0';
    layer1_outputs(7356) <= a;
    layer1_outputs(7357) <= not (a xor b);
    layer1_outputs(7358) <= a;
    layer1_outputs(7359) <= not (a or b);
    layer1_outputs(7360) <= a and b;
    layer1_outputs(7361) <= not a;
    layer1_outputs(7362) <= b;
    layer1_outputs(7363) <= not (a or b);
    layer1_outputs(7364) <= not a;
    layer1_outputs(7365) <= not b or a;
    layer1_outputs(7366) <= a;
    layer1_outputs(7367) <= not (a and b);
    layer1_outputs(7368) <= not (a and b);
    layer1_outputs(7369) <= a xor b;
    layer1_outputs(7370) <= '0';
    layer1_outputs(7371) <= not (a or b);
    layer1_outputs(7372) <= not a or b;
    layer1_outputs(7373) <= '0';
    layer1_outputs(7374) <= '0';
    layer1_outputs(7375) <= a and b;
    layer1_outputs(7376) <= a or b;
    layer1_outputs(7377) <= not b or a;
    layer1_outputs(7378) <= '0';
    layer1_outputs(7379) <= not a;
    layer1_outputs(7380) <= a or b;
    layer1_outputs(7381) <= '0';
    layer1_outputs(7382) <= b;
    layer1_outputs(7383) <= a and b;
    layer1_outputs(7384) <= not (a or b);
    layer1_outputs(7385) <= not (a xor b);
    layer1_outputs(7386) <= not b;
    layer1_outputs(7387) <= a or b;
    layer1_outputs(7388) <= b;
    layer1_outputs(7389) <= a;
    layer1_outputs(7390) <= a or b;
    layer1_outputs(7391) <= a or b;
    layer1_outputs(7392) <= not (a and b);
    layer1_outputs(7393) <= not b or a;
    layer1_outputs(7394) <= a;
    layer1_outputs(7395) <= '1';
    layer1_outputs(7396) <= '1';
    layer1_outputs(7397) <= not b;
    layer1_outputs(7398) <= not (a or b);
    layer1_outputs(7399) <= not a or b;
    layer1_outputs(7400) <= '0';
    layer1_outputs(7401) <= a and not b;
    layer1_outputs(7402) <= '1';
    layer1_outputs(7403) <= not a or b;
    layer1_outputs(7404) <= '0';
    layer1_outputs(7405) <= not (a or b);
    layer1_outputs(7406) <= a xor b;
    layer1_outputs(7407) <= not a or b;
    layer1_outputs(7408) <= a and not b;
    layer1_outputs(7409) <= '0';
    layer1_outputs(7410) <= a or b;
    layer1_outputs(7411) <= '1';
    layer1_outputs(7412) <= b and not a;
    layer1_outputs(7413) <= b and not a;
    layer1_outputs(7414) <= '0';
    layer1_outputs(7415) <= not b;
    layer1_outputs(7416) <= a and not b;
    layer1_outputs(7417) <= a or b;
    layer1_outputs(7418) <= not a;
    layer1_outputs(7419) <= '1';
    layer1_outputs(7420) <= a or b;
    layer1_outputs(7421) <= a;
    layer1_outputs(7422) <= b and not a;
    layer1_outputs(7423) <= a and not b;
    layer1_outputs(7424) <= b and not a;
    layer1_outputs(7425) <= a and not b;
    layer1_outputs(7426) <= not a or b;
    layer1_outputs(7427) <= '1';
    layer1_outputs(7428) <= not (a or b);
    layer1_outputs(7429) <= b and not a;
    layer1_outputs(7430) <= '0';
    layer1_outputs(7431) <= not a or b;
    layer1_outputs(7432) <= '0';
    layer1_outputs(7433) <= a and not b;
    layer1_outputs(7434) <= b;
    layer1_outputs(7435) <= a and b;
    layer1_outputs(7436) <= '1';
    layer1_outputs(7437) <= not a or b;
    layer1_outputs(7438) <= '0';
    layer1_outputs(7439) <= '0';
    layer1_outputs(7440) <= not (a or b);
    layer1_outputs(7441) <= '1';
    layer1_outputs(7442) <= not a or b;
    layer1_outputs(7443) <= not b;
    layer1_outputs(7444) <= '0';
    layer1_outputs(7445) <= not (a or b);
    layer1_outputs(7446) <= a or b;
    layer1_outputs(7447) <= not a or b;
    layer1_outputs(7448) <= not a;
    layer1_outputs(7449) <= a or b;
    layer1_outputs(7450) <= not a;
    layer1_outputs(7451) <= b and not a;
    layer1_outputs(7452) <= not a;
    layer1_outputs(7453) <= a or b;
    layer1_outputs(7454) <= '0';
    layer1_outputs(7455) <= b and not a;
    layer1_outputs(7456) <= not a or b;
    layer1_outputs(7457) <= a and b;
    layer1_outputs(7458) <= b and not a;
    layer1_outputs(7459) <= '0';
    layer1_outputs(7460) <= a or b;
    layer1_outputs(7461) <= b and not a;
    layer1_outputs(7462) <= not (a and b);
    layer1_outputs(7463) <= b and not a;
    layer1_outputs(7464) <= not b;
    layer1_outputs(7465) <= not (a or b);
    layer1_outputs(7466) <= a;
    layer1_outputs(7467) <= a;
    layer1_outputs(7468) <= not a;
    layer1_outputs(7469) <= a and not b;
    layer1_outputs(7470) <= a or b;
    layer1_outputs(7471) <= not b or a;
    layer1_outputs(7472) <= a;
    layer1_outputs(7473) <= a;
    layer1_outputs(7474) <= not (a or b);
    layer1_outputs(7475) <= a and b;
    layer1_outputs(7476) <= '0';
    layer1_outputs(7477) <= '0';
    layer1_outputs(7478) <= b;
    layer1_outputs(7479) <= not b;
    layer1_outputs(7480) <= not (a and b);
    layer1_outputs(7481) <= a;
    layer1_outputs(7482) <= b;
    layer1_outputs(7483) <= b and not a;
    layer1_outputs(7484) <= a and b;
    layer1_outputs(7485) <= b and not a;
    layer1_outputs(7486) <= not b or a;
    layer1_outputs(7487) <= not b or a;
    layer1_outputs(7488) <= not a or b;
    layer1_outputs(7489) <= a and not b;
    layer1_outputs(7490) <= not a or b;
    layer1_outputs(7491) <= not a;
    layer1_outputs(7492) <= a or b;
    layer1_outputs(7493) <= a;
    layer1_outputs(7494) <= a xor b;
    layer1_outputs(7495) <= a or b;
    layer1_outputs(7496) <= a or b;
    layer1_outputs(7497) <= '0';
    layer1_outputs(7498) <= not (a or b);
    layer1_outputs(7499) <= a and not b;
    layer1_outputs(7500) <= not b;
    layer1_outputs(7501) <= a and b;
    layer1_outputs(7502) <= b;
    layer1_outputs(7503) <= b and not a;
    layer1_outputs(7504) <= not b;
    layer1_outputs(7505) <= not b or a;
    layer1_outputs(7506) <= a;
    layer1_outputs(7507) <= not (a or b);
    layer1_outputs(7508) <= '1';
    layer1_outputs(7509) <= '1';
    layer1_outputs(7510) <= not a;
    layer1_outputs(7511) <= b;
    layer1_outputs(7512) <= not a or b;
    layer1_outputs(7513) <= not a;
    layer1_outputs(7514) <= not b;
    layer1_outputs(7515) <= not (a and b);
    layer1_outputs(7516) <= not b or a;
    layer1_outputs(7517) <= not b or a;
    layer1_outputs(7518) <= '1';
    layer1_outputs(7519) <= not b or a;
    layer1_outputs(7520) <= b and not a;
    layer1_outputs(7521) <= '1';
    layer1_outputs(7522) <= a and not b;
    layer1_outputs(7523) <= not b;
    layer1_outputs(7524) <= not a;
    layer1_outputs(7525) <= b and not a;
    layer1_outputs(7526) <= not a;
    layer1_outputs(7527) <= a or b;
    layer1_outputs(7528) <= not (a or b);
    layer1_outputs(7529) <= not b or a;
    layer1_outputs(7530) <= not (a or b);
    layer1_outputs(7531) <= '0';
    layer1_outputs(7532) <= a and not b;
    layer1_outputs(7533) <= not (a and b);
    layer1_outputs(7534) <= a or b;
    layer1_outputs(7535) <= not b;
    layer1_outputs(7536) <= a and b;
    layer1_outputs(7537) <= not a;
    layer1_outputs(7538) <= '1';
    layer1_outputs(7539) <= not a or b;
    layer1_outputs(7540) <= a and b;
    layer1_outputs(7541) <= b;
    layer1_outputs(7542) <= a;
    layer1_outputs(7543) <= not a or b;
    layer1_outputs(7544) <= a xor b;
    layer1_outputs(7545) <= a and b;
    layer1_outputs(7546) <= '0';
    layer1_outputs(7547) <= not (a or b);
    layer1_outputs(7548) <= not (a xor b);
    layer1_outputs(7549) <= b;
    layer1_outputs(7550) <= b;
    layer1_outputs(7551) <= not (a or b);
    layer1_outputs(7552) <= not (a or b);
    layer1_outputs(7553) <= '1';
    layer1_outputs(7554) <= b and not a;
    layer1_outputs(7555) <= b and not a;
    layer1_outputs(7556) <= not a or b;
    layer1_outputs(7557) <= not (a and b);
    layer1_outputs(7558) <= a;
    layer1_outputs(7559) <= '0';
    layer1_outputs(7560) <= a or b;
    layer1_outputs(7561) <= '0';
    layer1_outputs(7562) <= not (a and b);
    layer1_outputs(7563) <= '1';
    layer1_outputs(7564) <= '1';
    layer1_outputs(7565) <= a and b;
    layer1_outputs(7566) <= not (a xor b);
    layer1_outputs(7567) <= not a;
    layer1_outputs(7568) <= not b or a;
    layer1_outputs(7569) <= b and not a;
    layer1_outputs(7570) <= not a or b;
    layer1_outputs(7571) <= not (a and b);
    layer1_outputs(7572) <= not (a xor b);
    layer1_outputs(7573) <= a;
    layer1_outputs(7574) <= a;
    layer1_outputs(7575) <= a and not b;
    layer1_outputs(7576) <= not b or a;
    layer1_outputs(7577) <= '1';
    layer1_outputs(7578) <= not b or a;
    layer1_outputs(7579) <= not (a and b);
    layer1_outputs(7580) <= '1';
    layer1_outputs(7581) <= not a;
    layer1_outputs(7582) <= a;
    layer1_outputs(7583) <= '1';
    layer1_outputs(7584) <= '1';
    layer1_outputs(7585) <= not b or a;
    layer1_outputs(7586) <= a or b;
    layer1_outputs(7587) <= not a;
    layer1_outputs(7588) <= b and not a;
    layer1_outputs(7589) <= not b or a;
    layer1_outputs(7590) <= b;
    layer1_outputs(7591) <= not (a and b);
    layer1_outputs(7592) <= a;
    layer1_outputs(7593) <= not b or a;
    layer1_outputs(7594) <= not a;
    layer1_outputs(7595) <= not a or b;
    layer1_outputs(7596) <= b and not a;
    layer1_outputs(7597) <= a and b;
    layer1_outputs(7598) <= a and not b;
    layer1_outputs(7599) <= a or b;
    layer1_outputs(7600) <= not (a xor b);
    layer1_outputs(7601) <= not a;
    layer1_outputs(7602) <= not b;
    layer1_outputs(7603) <= a or b;
    layer1_outputs(7604) <= b;
    layer1_outputs(7605) <= a or b;
    layer1_outputs(7606) <= a xor b;
    layer1_outputs(7607) <= not (a xor b);
    layer1_outputs(7608) <= a and b;
    layer1_outputs(7609) <= a and not b;
    layer1_outputs(7610) <= a and b;
    layer1_outputs(7611) <= not (a or b);
    layer1_outputs(7612) <= '1';
    layer1_outputs(7613) <= not b or a;
    layer1_outputs(7614) <= '0';
    layer1_outputs(7615) <= not b or a;
    layer1_outputs(7616) <= not b;
    layer1_outputs(7617) <= not a;
    layer1_outputs(7618) <= not b or a;
    layer1_outputs(7619) <= not b;
    layer1_outputs(7620) <= a and b;
    layer1_outputs(7621) <= '1';
    layer1_outputs(7622) <= a and b;
    layer1_outputs(7623) <= not b or a;
    layer1_outputs(7624) <= b and not a;
    layer1_outputs(7625) <= not a or b;
    layer1_outputs(7626) <= '0';
    layer1_outputs(7627) <= b and not a;
    layer1_outputs(7628) <= a and not b;
    layer1_outputs(7629) <= not b or a;
    layer1_outputs(7630) <= not b or a;
    layer1_outputs(7631) <= a or b;
    layer1_outputs(7632) <= not b or a;
    layer1_outputs(7633) <= '0';
    layer1_outputs(7634) <= not (a and b);
    layer1_outputs(7635) <= a;
    layer1_outputs(7636) <= a;
    layer1_outputs(7637) <= not a or b;
    layer1_outputs(7638) <= '1';
    layer1_outputs(7639) <= a or b;
    layer1_outputs(7640) <= a and b;
    layer1_outputs(7641) <= not a;
    layer1_outputs(7642) <= not a or b;
    layer1_outputs(7643) <= b and not a;
    layer1_outputs(7644) <= a or b;
    layer1_outputs(7645) <= '0';
    layer1_outputs(7646) <= '0';
    layer1_outputs(7647) <= not (a or b);
    layer1_outputs(7648) <= b;
    layer1_outputs(7649) <= not b;
    layer1_outputs(7650) <= not a or b;
    layer1_outputs(7651) <= a or b;
    layer1_outputs(7652) <= a or b;
    layer1_outputs(7653) <= not (a and b);
    layer1_outputs(7654) <= not a or b;
    layer1_outputs(7655) <= not (a xor b);
    layer1_outputs(7656) <= a or b;
    layer1_outputs(7657) <= '0';
    layer1_outputs(7658) <= not a;
    layer1_outputs(7659) <= not (a or b);
    layer1_outputs(7660) <= not b or a;
    layer1_outputs(7661) <= not (a and b);
    layer1_outputs(7662) <= '1';
    layer1_outputs(7663) <= a and b;
    layer1_outputs(7664) <= not b or a;
    layer1_outputs(7665) <= '1';
    layer1_outputs(7666) <= a or b;
    layer1_outputs(7667) <= not (a and b);
    layer1_outputs(7668) <= a and not b;
    layer1_outputs(7669) <= a;
    layer1_outputs(7670) <= '1';
    layer1_outputs(7671) <= b;
    layer1_outputs(7672) <= not b or a;
    layer1_outputs(7673) <= '0';
    layer1_outputs(7674) <= not (a and b);
    layer1_outputs(7675) <= not b;
    layer1_outputs(7676) <= b;
    layer1_outputs(7677) <= not a or b;
    layer1_outputs(7678) <= not a;
    layer1_outputs(7679) <= a;
    layer2_outputs(0) <= not b or a;
    layer2_outputs(1) <= a and b;
    layer2_outputs(2) <= b;
    layer2_outputs(3) <= not b;
    layer2_outputs(4) <= a;
    layer2_outputs(5) <= not (a and b);
    layer2_outputs(6) <= not (a xor b);
    layer2_outputs(7) <= a;
    layer2_outputs(8) <= b;
    layer2_outputs(9) <= a;
    layer2_outputs(10) <= b and not a;
    layer2_outputs(11) <= '0';
    layer2_outputs(12) <= a;
    layer2_outputs(13) <= not a;
    layer2_outputs(14) <= not a;
    layer2_outputs(15) <= '1';
    layer2_outputs(16) <= not (a and b);
    layer2_outputs(17) <= not a or b;
    layer2_outputs(18) <= b;
    layer2_outputs(19) <= b;
    layer2_outputs(20) <= not a;
    layer2_outputs(21) <= a xor b;
    layer2_outputs(22) <= b and not a;
    layer2_outputs(23) <= '0';
    layer2_outputs(24) <= b and not a;
    layer2_outputs(25) <= a or b;
    layer2_outputs(26) <= a;
    layer2_outputs(27) <= '0';
    layer2_outputs(28) <= b and not a;
    layer2_outputs(29) <= a and not b;
    layer2_outputs(30) <= b and not a;
    layer2_outputs(31) <= '0';
    layer2_outputs(32) <= '0';
    layer2_outputs(33) <= a;
    layer2_outputs(34) <= b and not a;
    layer2_outputs(35) <= b;
    layer2_outputs(36) <= not (a or b);
    layer2_outputs(37) <= not b or a;
    layer2_outputs(38) <= '1';
    layer2_outputs(39) <= '1';
    layer2_outputs(40) <= '1';
    layer2_outputs(41) <= b;
    layer2_outputs(42) <= a;
    layer2_outputs(43) <= not a;
    layer2_outputs(44) <= not b or a;
    layer2_outputs(45) <= not b;
    layer2_outputs(46) <= not a or b;
    layer2_outputs(47) <= a and not b;
    layer2_outputs(48) <= a;
    layer2_outputs(49) <= a;
    layer2_outputs(50) <= not (a or b);
    layer2_outputs(51) <= not a or b;
    layer2_outputs(52) <= a and not b;
    layer2_outputs(53) <= b;
    layer2_outputs(54) <= b;
    layer2_outputs(55) <= not a or b;
    layer2_outputs(56) <= a;
    layer2_outputs(57) <= a and not b;
    layer2_outputs(58) <= b and not a;
    layer2_outputs(59) <= a;
    layer2_outputs(60) <= b and not a;
    layer2_outputs(61) <= not b or a;
    layer2_outputs(62) <= not b;
    layer2_outputs(63) <= a or b;
    layer2_outputs(64) <= a or b;
    layer2_outputs(65) <= b;
    layer2_outputs(66) <= '0';
    layer2_outputs(67) <= not a;
    layer2_outputs(68) <= not (a or b);
    layer2_outputs(69) <= '0';
    layer2_outputs(70) <= b;
    layer2_outputs(71) <= not (a and b);
    layer2_outputs(72) <= not (a or b);
    layer2_outputs(73) <= not (a xor b);
    layer2_outputs(74) <= not b;
    layer2_outputs(75) <= not a;
    layer2_outputs(76) <= not b;
    layer2_outputs(77) <= not a;
    layer2_outputs(78) <= a;
    layer2_outputs(79) <= not (a and b);
    layer2_outputs(80) <= a;
    layer2_outputs(81) <= not (a or b);
    layer2_outputs(82) <= a and not b;
    layer2_outputs(83) <= not a or b;
    layer2_outputs(84) <= not b or a;
    layer2_outputs(85) <= a and not b;
    layer2_outputs(86) <= not (a and b);
    layer2_outputs(87) <= not a or b;
    layer2_outputs(88) <= b;
    layer2_outputs(89) <= b;
    layer2_outputs(90) <= '1';
    layer2_outputs(91) <= a;
    layer2_outputs(92) <= '1';
    layer2_outputs(93) <= not (a or b);
    layer2_outputs(94) <= not b or a;
    layer2_outputs(95) <= not b;
    layer2_outputs(96) <= '0';
    layer2_outputs(97) <= '1';
    layer2_outputs(98) <= b;
    layer2_outputs(99) <= not a or b;
    layer2_outputs(100) <= a and not b;
    layer2_outputs(101) <= a and b;
    layer2_outputs(102) <= b and not a;
    layer2_outputs(103) <= a;
    layer2_outputs(104) <= not (a or b);
    layer2_outputs(105) <= not b or a;
    layer2_outputs(106) <= '1';
    layer2_outputs(107) <= not b or a;
    layer2_outputs(108) <= a and b;
    layer2_outputs(109) <= b;
    layer2_outputs(110) <= not a or b;
    layer2_outputs(111) <= not a or b;
    layer2_outputs(112) <= a and b;
    layer2_outputs(113) <= not (a or b);
    layer2_outputs(114) <= a or b;
    layer2_outputs(115) <= not (a and b);
    layer2_outputs(116) <= not a;
    layer2_outputs(117) <= not b or a;
    layer2_outputs(118) <= not (a and b);
    layer2_outputs(119) <= not a;
    layer2_outputs(120) <= not b or a;
    layer2_outputs(121) <= not a or b;
    layer2_outputs(122) <= not (a and b);
    layer2_outputs(123) <= '0';
    layer2_outputs(124) <= a or b;
    layer2_outputs(125) <= a and b;
    layer2_outputs(126) <= not (a and b);
    layer2_outputs(127) <= not b or a;
    layer2_outputs(128) <= a and not b;
    layer2_outputs(129) <= '1';
    layer2_outputs(130) <= '1';
    layer2_outputs(131) <= b;
    layer2_outputs(132) <= a and b;
    layer2_outputs(133) <= not (a and b);
    layer2_outputs(134) <= a and not b;
    layer2_outputs(135) <= b;
    layer2_outputs(136) <= a and b;
    layer2_outputs(137) <= '0';
    layer2_outputs(138) <= a;
    layer2_outputs(139) <= '1';
    layer2_outputs(140) <= a or b;
    layer2_outputs(141) <= '1';
    layer2_outputs(142) <= a;
    layer2_outputs(143) <= not (a xor b);
    layer2_outputs(144) <= a and b;
    layer2_outputs(145) <= a xor b;
    layer2_outputs(146) <= b and not a;
    layer2_outputs(147) <= not (a and b);
    layer2_outputs(148) <= b;
    layer2_outputs(149) <= a or b;
    layer2_outputs(150) <= a or b;
    layer2_outputs(151) <= not (a or b);
    layer2_outputs(152) <= a;
    layer2_outputs(153) <= not (a or b);
    layer2_outputs(154) <= b and not a;
    layer2_outputs(155) <= a and b;
    layer2_outputs(156) <= not b;
    layer2_outputs(157) <= '0';
    layer2_outputs(158) <= a or b;
    layer2_outputs(159) <= not a or b;
    layer2_outputs(160) <= a and not b;
    layer2_outputs(161) <= b and not a;
    layer2_outputs(162) <= a and b;
    layer2_outputs(163) <= a and b;
    layer2_outputs(164) <= a;
    layer2_outputs(165) <= a or b;
    layer2_outputs(166) <= not b;
    layer2_outputs(167) <= '0';
    layer2_outputs(168) <= a and b;
    layer2_outputs(169) <= not a or b;
    layer2_outputs(170) <= b and not a;
    layer2_outputs(171) <= not a or b;
    layer2_outputs(172) <= not a;
    layer2_outputs(173) <= '1';
    layer2_outputs(174) <= a and not b;
    layer2_outputs(175) <= not (a and b);
    layer2_outputs(176) <= b;
    layer2_outputs(177) <= a and b;
    layer2_outputs(178) <= a xor b;
    layer2_outputs(179) <= not (a and b);
    layer2_outputs(180) <= not b;
    layer2_outputs(181) <= not a or b;
    layer2_outputs(182) <= a xor b;
    layer2_outputs(183) <= a and not b;
    layer2_outputs(184) <= not b;
    layer2_outputs(185) <= not a;
    layer2_outputs(186) <= a xor b;
    layer2_outputs(187) <= not b;
    layer2_outputs(188) <= not (a and b);
    layer2_outputs(189) <= not (a or b);
    layer2_outputs(190) <= b;
    layer2_outputs(191) <= a and b;
    layer2_outputs(192) <= not a;
    layer2_outputs(193) <= b and not a;
    layer2_outputs(194) <= not a;
    layer2_outputs(195) <= b;
    layer2_outputs(196) <= '0';
    layer2_outputs(197) <= '1';
    layer2_outputs(198) <= a or b;
    layer2_outputs(199) <= a and not b;
    layer2_outputs(200) <= not (a or b);
    layer2_outputs(201) <= not a;
    layer2_outputs(202) <= not (a xor b);
    layer2_outputs(203) <= not a or b;
    layer2_outputs(204) <= b;
    layer2_outputs(205) <= not b;
    layer2_outputs(206) <= not b or a;
    layer2_outputs(207) <= '1';
    layer2_outputs(208) <= '1';
    layer2_outputs(209) <= not b or a;
    layer2_outputs(210) <= '1';
    layer2_outputs(211) <= a;
    layer2_outputs(212) <= '0';
    layer2_outputs(213) <= not a or b;
    layer2_outputs(214) <= not (a or b);
    layer2_outputs(215) <= a or b;
    layer2_outputs(216) <= b;
    layer2_outputs(217) <= a and not b;
    layer2_outputs(218) <= a;
    layer2_outputs(219) <= not a or b;
    layer2_outputs(220) <= b and not a;
    layer2_outputs(221) <= b and not a;
    layer2_outputs(222) <= a;
    layer2_outputs(223) <= not a or b;
    layer2_outputs(224) <= a xor b;
    layer2_outputs(225) <= a and not b;
    layer2_outputs(226) <= a and not b;
    layer2_outputs(227) <= not b;
    layer2_outputs(228) <= b and not a;
    layer2_outputs(229) <= not a;
    layer2_outputs(230) <= a or b;
    layer2_outputs(231) <= a xor b;
    layer2_outputs(232) <= not b;
    layer2_outputs(233) <= a;
    layer2_outputs(234) <= not b;
    layer2_outputs(235) <= a and b;
    layer2_outputs(236) <= a or b;
    layer2_outputs(237) <= not (a xor b);
    layer2_outputs(238) <= not (a xor b);
    layer2_outputs(239) <= a or b;
    layer2_outputs(240) <= a or b;
    layer2_outputs(241) <= b and not a;
    layer2_outputs(242) <= a xor b;
    layer2_outputs(243) <= '0';
    layer2_outputs(244) <= a and b;
    layer2_outputs(245) <= '1';
    layer2_outputs(246) <= not (a or b);
    layer2_outputs(247) <= not b or a;
    layer2_outputs(248) <= not b or a;
    layer2_outputs(249) <= not (a or b);
    layer2_outputs(250) <= not b or a;
    layer2_outputs(251) <= b;
    layer2_outputs(252) <= a and not b;
    layer2_outputs(253) <= not b;
    layer2_outputs(254) <= not (a or b);
    layer2_outputs(255) <= not a;
    layer2_outputs(256) <= '1';
    layer2_outputs(257) <= b;
    layer2_outputs(258) <= not (a or b);
    layer2_outputs(259) <= not b;
    layer2_outputs(260) <= not (a and b);
    layer2_outputs(261) <= b and not a;
    layer2_outputs(262) <= a and b;
    layer2_outputs(263) <= b and not a;
    layer2_outputs(264) <= not (a or b);
    layer2_outputs(265) <= a and not b;
    layer2_outputs(266) <= a or b;
    layer2_outputs(267) <= not (a and b);
    layer2_outputs(268) <= b;
    layer2_outputs(269) <= b and not a;
    layer2_outputs(270) <= a or b;
    layer2_outputs(271) <= '0';
    layer2_outputs(272) <= not a;
    layer2_outputs(273) <= b and not a;
    layer2_outputs(274) <= not a or b;
    layer2_outputs(275) <= a;
    layer2_outputs(276) <= not b;
    layer2_outputs(277) <= not b or a;
    layer2_outputs(278) <= a and not b;
    layer2_outputs(279) <= '1';
    layer2_outputs(280) <= not (a or b);
    layer2_outputs(281) <= not a;
    layer2_outputs(282) <= a or b;
    layer2_outputs(283) <= not (a and b);
    layer2_outputs(284) <= not (a and b);
    layer2_outputs(285) <= '0';
    layer2_outputs(286) <= not a;
    layer2_outputs(287) <= not b or a;
    layer2_outputs(288) <= not b or a;
    layer2_outputs(289) <= b and not a;
    layer2_outputs(290) <= not b;
    layer2_outputs(291) <= a and b;
    layer2_outputs(292) <= not a or b;
    layer2_outputs(293) <= a;
    layer2_outputs(294) <= '1';
    layer2_outputs(295) <= a and not b;
    layer2_outputs(296) <= not (a and b);
    layer2_outputs(297) <= a;
    layer2_outputs(298) <= a and b;
    layer2_outputs(299) <= a and not b;
    layer2_outputs(300) <= not a;
    layer2_outputs(301) <= b and not a;
    layer2_outputs(302) <= a and b;
    layer2_outputs(303) <= not (a or b);
    layer2_outputs(304) <= b and not a;
    layer2_outputs(305) <= '1';
    layer2_outputs(306) <= not (a and b);
    layer2_outputs(307) <= not a or b;
    layer2_outputs(308) <= b and not a;
    layer2_outputs(309) <= b;
    layer2_outputs(310) <= '0';
    layer2_outputs(311) <= b and not a;
    layer2_outputs(312) <= not b or a;
    layer2_outputs(313) <= '1';
    layer2_outputs(314) <= '0';
    layer2_outputs(315) <= a or b;
    layer2_outputs(316) <= a;
    layer2_outputs(317) <= b and not a;
    layer2_outputs(318) <= '1';
    layer2_outputs(319) <= a and b;
    layer2_outputs(320) <= a and not b;
    layer2_outputs(321) <= '1';
    layer2_outputs(322) <= '0';
    layer2_outputs(323) <= '0';
    layer2_outputs(324) <= b;
    layer2_outputs(325) <= not b or a;
    layer2_outputs(326) <= '0';
    layer2_outputs(327) <= a;
    layer2_outputs(328) <= '1';
    layer2_outputs(329) <= not b;
    layer2_outputs(330) <= a and not b;
    layer2_outputs(331) <= b;
    layer2_outputs(332) <= b and not a;
    layer2_outputs(333) <= not b;
    layer2_outputs(334) <= not (a and b);
    layer2_outputs(335) <= not b;
    layer2_outputs(336) <= not (a and b);
    layer2_outputs(337) <= not b;
    layer2_outputs(338) <= not a;
    layer2_outputs(339) <= not b;
    layer2_outputs(340) <= '1';
    layer2_outputs(341) <= b;
    layer2_outputs(342) <= a and b;
    layer2_outputs(343) <= not b;
    layer2_outputs(344) <= '1';
    layer2_outputs(345) <= '0';
    layer2_outputs(346) <= '0';
    layer2_outputs(347) <= a and b;
    layer2_outputs(348) <= b and not a;
    layer2_outputs(349) <= a and not b;
    layer2_outputs(350) <= a and b;
    layer2_outputs(351) <= not (a and b);
    layer2_outputs(352) <= '0';
    layer2_outputs(353) <= '1';
    layer2_outputs(354) <= not (a or b);
    layer2_outputs(355) <= not a;
    layer2_outputs(356) <= b;
    layer2_outputs(357) <= not a;
    layer2_outputs(358) <= a and not b;
    layer2_outputs(359) <= not a or b;
    layer2_outputs(360) <= '0';
    layer2_outputs(361) <= '0';
    layer2_outputs(362) <= a and b;
    layer2_outputs(363) <= b and not a;
    layer2_outputs(364) <= a and not b;
    layer2_outputs(365) <= not b or a;
    layer2_outputs(366) <= '0';
    layer2_outputs(367) <= '1';
    layer2_outputs(368) <= a or b;
    layer2_outputs(369) <= not a or b;
    layer2_outputs(370) <= a;
    layer2_outputs(371) <= a;
    layer2_outputs(372) <= not a;
    layer2_outputs(373) <= not (a xor b);
    layer2_outputs(374) <= a and b;
    layer2_outputs(375) <= not (a or b);
    layer2_outputs(376) <= '0';
    layer2_outputs(377) <= '0';
    layer2_outputs(378) <= '0';
    layer2_outputs(379) <= not (a and b);
    layer2_outputs(380) <= not (a or b);
    layer2_outputs(381) <= not a;
    layer2_outputs(382) <= '0';
    layer2_outputs(383) <= a and not b;
    layer2_outputs(384) <= not a;
    layer2_outputs(385) <= not b or a;
    layer2_outputs(386) <= not b or a;
    layer2_outputs(387) <= '0';
    layer2_outputs(388) <= not a or b;
    layer2_outputs(389) <= not a;
    layer2_outputs(390) <= '0';
    layer2_outputs(391) <= '1';
    layer2_outputs(392) <= '1';
    layer2_outputs(393) <= b;
    layer2_outputs(394) <= '0';
    layer2_outputs(395) <= not b or a;
    layer2_outputs(396) <= a and b;
    layer2_outputs(397) <= not a or b;
    layer2_outputs(398) <= a and b;
    layer2_outputs(399) <= '1';
    layer2_outputs(400) <= not (a and b);
    layer2_outputs(401) <= b and not a;
    layer2_outputs(402) <= a or b;
    layer2_outputs(403) <= '1';
    layer2_outputs(404) <= a and b;
    layer2_outputs(405) <= not a or b;
    layer2_outputs(406) <= '1';
    layer2_outputs(407) <= '1';
    layer2_outputs(408) <= not (a and b);
    layer2_outputs(409) <= a and b;
    layer2_outputs(410) <= '1';
    layer2_outputs(411) <= not a or b;
    layer2_outputs(412) <= not (a xor b);
    layer2_outputs(413) <= a xor b;
    layer2_outputs(414) <= a and not b;
    layer2_outputs(415) <= '1';
    layer2_outputs(416) <= a and b;
    layer2_outputs(417) <= '0';
    layer2_outputs(418) <= a;
    layer2_outputs(419) <= not b;
    layer2_outputs(420) <= a;
    layer2_outputs(421) <= not (a and b);
    layer2_outputs(422) <= b and not a;
    layer2_outputs(423) <= b;
    layer2_outputs(424) <= not a;
    layer2_outputs(425) <= not (a or b);
    layer2_outputs(426) <= not b;
    layer2_outputs(427) <= b and not a;
    layer2_outputs(428) <= '1';
    layer2_outputs(429) <= not b or a;
    layer2_outputs(430) <= a;
    layer2_outputs(431) <= '0';
    layer2_outputs(432) <= not a;
    layer2_outputs(433) <= a and not b;
    layer2_outputs(434) <= b and not a;
    layer2_outputs(435) <= not a;
    layer2_outputs(436) <= '1';
    layer2_outputs(437) <= b;
    layer2_outputs(438) <= '1';
    layer2_outputs(439) <= b and not a;
    layer2_outputs(440) <= not (a xor b);
    layer2_outputs(441) <= a and not b;
    layer2_outputs(442) <= b;
    layer2_outputs(443) <= a and not b;
    layer2_outputs(444) <= not (a or b);
    layer2_outputs(445) <= not b;
    layer2_outputs(446) <= a and b;
    layer2_outputs(447) <= not b or a;
    layer2_outputs(448) <= not a;
    layer2_outputs(449) <= a xor b;
    layer2_outputs(450) <= b;
    layer2_outputs(451) <= b;
    layer2_outputs(452) <= a or b;
    layer2_outputs(453) <= '1';
    layer2_outputs(454) <= b;
    layer2_outputs(455) <= a and b;
    layer2_outputs(456) <= not (a or b);
    layer2_outputs(457) <= '0';
    layer2_outputs(458) <= a;
    layer2_outputs(459) <= not b or a;
    layer2_outputs(460) <= '1';
    layer2_outputs(461) <= b;
    layer2_outputs(462) <= a and not b;
    layer2_outputs(463) <= a and b;
    layer2_outputs(464) <= '0';
    layer2_outputs(465) <= a and b;
    layer2_outputs(466) <= not (a xor b);
    layer2_outputs(467) <= not (a and b);
    layer2_outputs(468) <= not b;
    layer2_outputs(469) <= b;
    layer2_outputs(470) <= not a;
    layer2_outputs(471) <= a and not b;
    layer2_outputs(472) <= a and not b;
    layer2_outputs(473) <= not (a and b);
    layer2_outputs(474) <= '0';
    layer2_outputs(475) <= not b or a;
    layer2_outputs(476) <= '0';
    layer2_outputs(477) <= a and b;
    layer2_outputs(478) <= a xor b;
    layer2_outputs(479) <= a and b;
    layer2_outputs(480) <= a and not b;
    layer2_outputs(481) <= not a or b;
    layer2_outputs(482) <= a or b;
    layer2_outputs(483) <= not (a and b);
    layer2_outputs(484) <= a and b;
    layer2_outputs(485) <= not (a or b);
    layer2_outputs(486) <= not (a and b);
    layer2_outputs(487) <= not b;
    layer2_outputs(488) <= a;
    layer2_outputs(489) <= not a;
    layer2_outputs(490) <= '1';
    layer2_outputs(491) <= a;
    layer2_outputs(492) <= not a;
    layer2_outputs(493) <= a or b;
    layer2_outputs(494) <= a or b;
    layer2_outputs(495) <= '0';
    layer2_outputs(496) <= not (a and b);
    layer2_outputs(497) <= not b;
    layer2_outputs(498) <= not a;
    layer2_outputs(499) <= not a;
    layer2_outputs(500) <= a and not b;
    layer2_outputs(501) <= b and not a;
    layer2_outputs(502) <= not a;
    layer2_outputs(503) <= a xor b;
    layer2_outputs(504) <= a;
    layer2_outputs(505) <= not b;
    layer2_outputs(506) <= not a or b;
    layer2_outputs(507) <= not b;
    layer2_outputs(508) <= not (a and b);
    layer2_outputs(509) <= not a or b;
    layer2_outputs(510) <= not a or b;
    layer2_outputs(511) <= not (a and b);
    layer2_outputs(512) <= b and not a;
    layer2_outputs(513) <= '0';
    layer2_outputs(514) <= a or b;
    layer2_outputs(515) <= a xor b;
    layer2_outputs(516) <= not (a or b);
    layer2_outputs(517) <= '1';
    layer2_outputs(518) <= not (a or b);
    layer2_outputs(519) <= a and not b;
    layer2_outputs(520) <= a;
    layer2_outputs(521) <= not b;
    layer2_outputs(522) <= b and not a;
    layer2_outputs(523) <= b;
    layer2_outputs(524) <= not a;
    layer2_outputs(525) <= not b or a;
    layer2_outputs(526) <= a or b;
    layer2_outputs(527) <= a and not b;
    layer2_outputs(528) <= not a or b;
    layer2_outputs(529) <= not b or a;
    layer2_outputs(530) <= not a or b;
    layer2_outputs(531) <= '0';
    layer2_outputs(532) <= not (a or b);
    layer2_outputs(533) <= '1';
    layer2_outputs(534) <= not a or b;
    layer2_outputs(535) <= a;
    layer2_outputs(536) <= not (a or b);
    layer2_outputs(537) <= '1';
    layer2_outputs(538) <= not (a and b);
    layer2_outputs(539) <= '0';
    layer2_outputs(540) <= a or b;
    layer2_outputs(541) <= a or b;
    layer2_outputs(542) <= not (a and b);
    layer2_outputs(543) <= '0';
    layer2_outputs(544) <= a and b;
    layer2_outputs(545) <= not a or b;
    layer2_outputs(546) <= b and not a;
    layer2_outputs(547) <= b and not a;
    layer2_outputs(548) <= a or b;
    layer2_outputs(549) <= a and not b;
    layer2_outputs(550) <= '1';
    layer2_outputs(551) <= a and not b;
    layer2_outputs(552) <= b and not a;
    layer2_outputs(553) <= a or b;
    layer2_outputs(554) <= a xor b;
    layer2_outputs(555) <= b and not a;
    layer2_outputs(556) <= a;
    layer2_outputs(557) <= not (a xor b);
    layer2_outputs(558) <= a and b;
    layer2_outputs(559) <= '0';
    layer2_outputs(560) <= not (a and b);
    layer2_outputs(561) <= not (a and b);
    layer2_outputs(562) <= a or b;
    layer2_outputs(563) <= b and not a;
    layer2_outputs(564) <= not (a or b);
    layer2_outputs(565) <= b;
    layer2_outputs(566) <= b;
    layer2_outputs(567) <= not a;
    layer2_outputs(568) <= not b or a;
    layer2_outputs(569) <= not a;
    layer2_outputs(570) <= b and not a;
    layer2_outputs(571) <= a and b;
    layer2_outputs(572) <= not a;
    layer2_outputs(573) <= not a;
    layer2_outputs(574) <= a;
    layer2_outputs(575) <= b and not a;
    layer2_outputs(576) <= '1';
    layer2_outputs(577) <= not a or b;
    layer2_outputs(578) <= '1';
    layer2_outputs(579) <= a and b;
    layer2_outputs(580) <= a and not b;
    layer2_outputs(581) <= '1';
    layer2_outputs(582) <= not a;
    layer2_outputs(583) <= not (a and b);
    layer2_outputs(584) <= a or b;
    layer2_outputs(585) <= not a;
    layer2_outputs(586) <= '0';
    layer2_outputs(587) <= a or b;
    layer2_outputs(588) <= a and not b;
    layer2_outputs(589) <= b;
    layer2_outputs(590) <= not b;
    layer2_outputs(591) <= not b;
    layer2_outputs(592) <= a and b;
    layer2_outputs(593) <= a;
    layer2_outputs(594) <= not a;
    layer2_outputs(595) <= a;
    layer2_outputs(596) <= not a or b;
    layer2_outputs(597) <= not b;
    layer2_outputs(598) <= not a or b;
    layer2_outputs(599) <= not a;
    layer2_outputs(600) <= a and not b;
    layer2_outputs(601) <= a and b;
    layer2_outputs(602) <= not (a or b);
    layer2_outputs(603) <= a and b;
    layer2_outputs(604) <= not b or a;
    layer2_outputs(605) <= '0';
    layer2_outputs(606) <= not a;
    layer2_outputs(607) <= a;
    layer2_outputs(608) <= a and not b;
    layer2_outputs(609) <= '0';
    layer2_outputs(610) <= not (a xor b);
    layer2_outputs(611) <= a;
    layer2_outputs(612) <= not (a xor b);
    layer2_outputs(613) <= '0';
    layer2_outputs(614) <= b;
    layer2_outputs(615) <= a xor b;
    layer2_outputs(616) <= '0';
    layer2_outputs(617) <= not b;
    layer2_outputs(618) <= not a;
    layer2_outputs(619) <= b;
    layer2_outputs(620) <= not a or b;
    layer2_outputs(621) <= b;
    layer2_outputs(622) <= a or b;
    layer2_outputs(623) <= not b or a;
    layer2_outputs(624) <= a;
    layer2_outputs(625) <= not b or a;
    layer2_outputs(626) <= not (a and b);
    layer2_outputs(627) <= not (a or b);
    layer2_outputs(628) <= not (a and b);
    layer2_outputs(629) <= b;
    layer2_outputs(630) <= a and b;
    layer2_outputs(631) <= '0';
    layer2_outputs(632) <= '0';
    layer2_outputs(633) <= not (a or b);
    layer2_outputs(634) <= not a;
    layer2_outputs(635) <= not b;
    layer2_outputs(636) <= a xor b;
    layer2_outputs(637) <= b;
    layer2_outputs(638) <= not a or b;
    layer2_outputs(639) <= not a or b;
    layer2_outputs(640) <= a and not b;
    layer2_outputs(641) <= not (a and b);
    layer2_outputs(642) <= not (a and b);
    layer2_outputs(643) <= not b;
    layer2_outputs(644) <= b;
    layer2_outputs(645) <= '1';
    layer2_outputs(646) <= b;
    layer2_outputs(647) <= not (a or b);
    layer2_outputs(648) <= not b;
    layer2_outputs(649) <= not a or b;
    layer2_outputs(650) <= not a or b;
    layer2_outputs(651) <= '1';
    layer2_outputs(652) <= a;
    layer2_outputs(653) <= a and not b;
    layer2_outputs(654) <= not b;
    layer2_outputs(655) <= not (a and b);
    layer2_outputs(656) <= a and not b;
    layer2_outputs(657) <= not a or b;
    layer2_outputs(658) <= b;
    layer2_outputs(659) <= a and not b;
    layer2_outputs(660) <= a and b;
    layer2_outputs(661) <= not (a or b);
    layer2_outputs(662) <= not b or a;
    layer2_outputs(663) <= '0';
    layer2_outputs(664) <= not (a xor b);
    layer2_outputs(665) <= a or b;
    layer2_outputs(666) <= a and not b;
    layer2_outputs(667) <= a or b;
    layer2_outputs(668) <= a and b;
    layer2_outputs(669) <= a;
    layer2_outputs(670) <= a and b;
    layer2_outputs(671) <= not b or a;
    layer2_outputs(672) <= not (a xor b);
    layer2_outputs(673) <= not (a or b);
    layer2_outputs(674) <= '0';
    layer2_outputs(675) <= a;
    layer2_outputs(676) <= a and not b;
    layer2_outputs(677) <= '0';
    layer2_outputs(678) <= '0';
    layer2_outputs(679) <= not a or b;
    layer2_outputs(680) <= not (a or b);
    layer2_outputs(681) <= b;
    layer2_outputs(682) <= not b;
    layer2_outputs(683) <= '0';
    layer2_outputs(684) <= not b or a;
    layer2_outputs(685) <= a and not b;
    layer2_outputs(686) <= a or b;
    layer2_outputs(687) <= b;
    layer2_outputs(688) <= not (a or b);
    layer2_outputs(689) <= b and not a;
    layer2_outputs(690) <= a and b;
    layer2_outputs(691) <= not b or a;
    layer2_outputs(692) <= not a;
    layer2_outputs(693) <= a and b;
    layer2_outputs(694) <= not (a or b);
    layer2_outputs(695) <= '0';
    layer2_outputs(696) <= b;
    layer2_outputs(697) <= '0';
    layer2_outputs(698) <= not a;
    layer2_outputs(699) <= a or b;
    layer2_outputs(700) <= a and not b;
    layer2_outputs(701) <= a and b;
    layer2_outputs(702) <= a and not b;
    layer2_outputs(703) <= not (a and b);
    layer2_outputs(704) <= b and not a;
    layer2_outputs(705) <= '1';
    layer2_outputs(706) <= '1';
    layer2_outputs(707) <= b and not a;
    layer2_outputs(708) <= a and b;
    layer2_outputs(709) <= not b;
    layer2_outputs(710) <= not b or a;
    layer2_outputs(711) <= '0';
    layer2_outputs(712) <= '1';
    layer2_outputs(713) <= '0';
    layer2_outputs(714) <= a and b;
    layer2_outputs(715) <= not a;
    layer2_outputs(716) <= b and not a;
    layer2_outputs(717) <= not (a and b);
    layer2_outputs(718) <= not a;
    layer2_outputs(719) <= not b or a;
    layer2_outputs(720) <= a;
    layer2_outputs(721) <= a;
    layer2_outputs(722) <= not b or a;
    layer2_outputs(723) <= '0';
    layer2_outputs(724) <= '0';
    layer2_outputs(725) <= not (a or b);
    layer2_outputs(726) <= not a;
    layer2_outputs(727) <= b;
    layer2_outputs(728) <= '1';
    layer2_outputs(729) <= not b or a;
    layer2_outputs(730) <= a xor b;
    layer2_outputs(731) <= '0';
    layer2_outputs(732) <= not a or b;
    layer2_outputs(733) <= not a;
    layer2_outputs(734) <= a and not b;
    layer2_outputs(735) <= a xor b;
    layer2_outputs(736) <= b and not a;
    layer2_outputs(737) <= not b or a;
    layer2_outputs(738) <= not a;
    layer2_outputs(739) <= a;
    layer2_outputs(740) <= '1';
    layer2_outputs(741) <= not a or b;
    layer2_outputs(742) <= not a;
    layer2_outputs(743) <= a;
    layer2_outputs(744) <= '0';
    layer2_outputs(745) <= '0';
    layer2_outputs(746) <= not (a and b);
    layer2_outputs(747) <= b and not a;
    layer2_outputs(748) <= a;
    layer2_outputs(749) <= '1';
    layer2_outputs(750) <= not a;
    layer2_outputs(751) <= not (a xor b);
    layer2_outputs(752) <= not (a or b);
    layer2_outputs(753) <= not a or b;
    layer2_outputs(754) <= not a;
    layer2_outputs(755) <= a;
    layer2_outputs(756) <= a and b;
    layer2_outputs(757) <= a;
    layer2_outputs(758) <= a;
    layer2_outputs(759) <= a or b;
    layer2_outputs(760) <= a;
    layer2_outputs(761) <= a xor b;
    layer2_outputs(762) <= b;
    layer2_outputs(763) <= a and b;
    layer2_outputs(764) <= a and b;
    layer2_outputs(765) <= not a;
    layer2_outputs(766) <= not (a or b);
    layer2_outputs(767) <= a or b;
    layer2_outputs(768) <= a or b;
    layer2_outputs(769) <= '0';
    layer2_outputs(770) <= not a;
    layer2_outputs(771) <= not (a and b);
    layer2_outputs(772) <= a and b;
    layer2_outputs(773) <= not (a or b);
    layer2_outputs(774) <= b and not a;
    layer2_outputs(775) <= not b or a;
    layer2_outputs(776) <= '0';
    layer2_outputs(777) <= not a;
    layer2_outputs(778) <= '1';
    layer2_outputs(779) <= not (a or b);
    layer2_outputs(780) <= not b or a;
    layer2_outputs(781) <= a and not b;
    layer2_outputs(782) <= a and not b;
    layer2_outputs(783) <= a and b;
    layer2_outputs(784) <= a xor b;
    layer2_outputs(785) <= a;
    layer2_outputs(786) <= b and not a;
    layer2_outputs(787) <= a;
    layer2_outputs(788) <= '1';
    layer2_outputs(789) <= not (a or b);
    layer2_outputs(790) <= not a or b;
    layer2_outputs(791) <= b and not a;
    layer2_outputs(792) <= not a;
    layer2_outputs(793) <= not a or b;
    layer2_outputs(794) <= not a or b;
    layer2_outputs(795) <= a;
    layer2_outputs(796) <= b;
    layer2_outputs(797) <= not b;
    layer2_outputs(798) <= a;
    layer2_outputs(799) <= not (a and b);
    layer2_outputs(800) <= '1';
    layer2_outputs(801) <= '1';
    layer2_outputs(802) <= not (a or b);
    layer2_outputs(803) <= a;
    layer2_outputs(804) <= a or b;
    layer2_outputs(805) <= not b or a;
    layer2_outputs(806) <= '0';
    layer2_outputs(807) <= a and not b;
    layer2_outputs(808) <= not (a and b);
    layer2_outputs(809) <= not b or a;
    layer2_outputs(810) <= a;
    layer2_outputs(811) <= not b or a;
    layer2_outputs(812) <= a;
    layer2_outputs(813) <= b;
    layer2_outputs(814) <= not b;
    layer2_outputs(815) <= not b;
    layer2_outputs(816) <= not (a and b);
    layer2_outputs(817) <= a and not b;
    layer2_outputs(818) <= '0';
    layer2_outputs(819) <= not a;
    layer2_outputs(820) <= not (a or b);
    layer2_outputs(821) <= not b or a;
    layer2_outputs(822) <= '0';
    layer2_outputs(823) <= b and not a;
    layer2_outputs(824) <= not a;
    layer2_outputs(825) <= not b;
    layer2_outputs(826) <= not (a or b);
    layer2_outputs(827) <= not a;
    layer2_outputs(828) <= a and b;
    layer2_outputs(829) <= a;
    layer2_outputs(830) <= b;
    layer2_outputs(831) <= not b or a;
    layer2_outputs(832) <= not b;
    layer2_outputs(833) <= a and b;
    layer2_outputs(834) <= not a or b;
    layer2_outputs(835) <= a and not b;
    layer2_outputs(836) <= a and b;
    layer2_outputs(837) <= a or b;
    layer2_outputs(838) <= a and not b;
    layer2_outputs(839) <= a or b;
    layer2_outputs(840) <= not b;
    layer2_outputs(841) <= a and not b;
    layer2_outputs(842) <= not (a xor b);
    layer2_outputs(843) <= a;
    layer2_outputs(844) <= '0';
    layer2_outputs(845) <= a and b;
    layer2_outputs(846) <= not (a or b);
    layer2_outputs(847) <= b;
    layer2_outputs(848) <= a and b;
    layer2_outputs(849) <= a or b;
    layer2_outputs(850) <= not a or b;
    layer2_outputs(851) <= not a;
    layer2_outputs(852) <= a or b;
    layer2_outputs(853) <= not a or b;
    layer2_outputs(854) <= a and b;
    layer2_outputs(855) <= not (a or b);
    layer2_outputs(856) <= not b or a;
    layer2_outputs(857) <= not a;
    layer2_outputs(858) <= a or b;
    layer2_outputs(859) <= a or b;
    layer2_outputs(860) <= a and b;
    layer2_outputs(861) <= a;
    layer2_outputs(862) <= not a;
    layer2_outputs(863) <= a and b;
    layer2_outputs(864) <= b and not a;
    layer2_outputs(865) <= '1';
    layer2_outputs(866) <= not (a and b);
    layer2_outputs(867) <= '1';
    layer2_outputs(868) <= '1';
    layer2_outputs(869) <= '1';
    layer2_outputs(870) <= '1';
    layer2_outputs(871) <= a and not b;
    layer2_outputs(872) <= not (a and b);
    layer2_outputs(873) <= not (a xor b);
    layer2_outputs(874) <= a;
    layer2_outputs(875) <= not b or a;
    layer2_outputs(876) <= not (a or b);
    layer2_outputs(877) <= not a or b;
    layer2_outputs(878) <= b and not a;
    layer2_outputs(879) <= '0';
    layer2_outputs(880) <= '1';
    layer2_outputs(881) <= '0';
    layer2_outputs(882) <= not b or a;
    layer2_outputs(883) <= a;
    layer2_outputs(884) <= a and not b;
    layer2_outputs(885) <= not (a and b);
    layer2_outputs(886) <= not (a and b);
    layer2_outputs(887) <= not b or a;
    layer2_outputs(888) <= not a;
    layer2_outputs(889) <= '1';
    layer2_outputs(890) <= '1';
    layer2_outputs(891) <= a and not b;
    layer2_outputs(892) <= '1';
    layer2_outputs(893) <= a or b;
    layer2_outputs(894) <= not b or a;
    layer2_outputs(895) <= not b;
    layer2_outputs(896) <= not a or b;
    layer2_outputs(897) <= '0';
    layer2_outputs(898) <= not a;
    layer2_outputs(899) <= not b or a;
    layer2_outputs(900) <= a or b;
    layer2_outputs(901) <= not a;
    layer2_outputs(902) <= '1';
    layer2_outputs(903) <= not (a xor b);
    layer2_outputs(904) <= a and not b;
    layer2_outputs(905) <= not b or a;
    layer2_outputs(906) <= a xor b;
    layer2_outputs(907) <= '1';
    layer2_outputs(908) <= a xor b;
    layer2_outputs(909) <= a xor b;
    layer2_outputs(910) <= not b or a;
    layer2_outputs(911) <= b and not a;
    layer2_outputs(912) <= a and b;
    layer2_outputs(913) <= '1';
    layer2_outputs(914) <= a or b;
    layer2_outputs(915) <= not a;
    layer2_outputs(916) <= not (a or b);
    layer2_outputs(917) <= '1';
    layer2_outputs(918) <= not (a or b);
    layer2_outputs(919) <= a or b;
    layer2_outputs(920) <= a and b;
    layer2_outputs(921) <= b and not a;
    layer2_outputs(922) <= not a;
    layer2_outputs(923) <= a;
    layer2_outputs(924) <= not b or a;
    layer2_outputs(925) <= not a or b;
    layer2_outputs(926) <= not b;
    layer2_outputs(927) <= not b or a;
    layer2_outputs(928) <= a and b;
    layer2_outputs(929) <= not (a and b);
    layer2_outputs(930) <= '0';
    layer2_outputs(931) <= '0';
    layer2_outputs(932) <= not b or a;
    layer2_outputs(933) <= a and b;
    layer2_outputs(934) <= a and b;
    layer2_outputs(935) <= a or b;
    layer2_outputs(936) <= b and not a;
    layer2_outputs(937) <= not b;
    layer2_outputs(938) <= a;
    layer2_outputs(939) <= not (a or b);
    layer2_outputs(940) <= a and b;
    layer2_outputs(941) <= a or b;
    layer2_outputs(942) <= not a;
    layer2_outputs(943) <= not b;
    layer2_outputs(944) <= not (a and b);
    layer2_outputs(945) <= a or b;
    layer2_outputs(946) <= not (a and b);
    layer2_outputs(947) <= a or b;
    layer2_outputs(948) <= b and not a;
    layer2_outputs(949) <= '0';
    layer2_outputs(950) <= not a;
    layer2_outputs(951) <= not (a or b);
    layer2_outputs(952) <= not b or a;
    layer2_outputs(953) <= a and b;
    layer2_outputs(954) <= a;
    layer2_outputs(955) <= not b;
    layer2_outputs(956) <= a and b;
    layer2_outputs(957) <= a or b;
    layer2_outputs(958) <= a and not b;
    layer2_outputs(959) <= a or b;
    layer2_outputs(960) <= b;
    layer2_outputs(961) <= not a or b;
    layer2_outputs(962) <= b;
    layer2_outputs(963) <= not a;
    layer2_outputs(964) <= not (a and b);
    layer2_outputs(965) <= a and not b;
    layer2_outputs(966) <= not a or b;
    layer2_outputs(967) <= a or b;
    layer2_outputs(968) <= not a;
    layer2_outputs(969) <= b;
    layer2_outputs(970) <= not a;
    layer2_outputs(971) <= a and b;
    layer2_outputs(972) <= not b;
    layer2_outputs(973) <= a and b;
    layer2_outputs(974) <= not (a and b);
    layer2_outputs(975) <= not b;
    layer2_outputs(976) <= a and not b;
    layer2_outputs(977) <= not a or b;
    layer2_outputs(978) <= a or b;
    layer2_outputs(979) <= '0';
    layer2_outputs(980) <= b and not a;
    layer2_outputs(981) <= a or b;
    layer2_outputs(982) <= a and not b;
    layer2_outputs(983) <= '0';
    layer2_outputs(984) <= not a;
    layer2_outputs(985) <= not (a or b);
    layer2_outputs(986) <= '1';
    layer2_outputs(987) <= not (a and b);
    layer2_outputs(988) <= a and b;
    layer2_outputs(989) <= '0';
    layer2_outputs(990) <= '0';
    layer2_outputs(991) <= '1';
    layer2_outputs(992) <= a and b;
    layer2_outputs(993) <= not a;
    layer2_outputs(994) <= not (a and b);
    layer2_outputs(995) <= b and not a;
    layer2_outputs(996) <= b and not a;
    layer2_outputs(997) <= a and b;
    layer2_outputs(998) <= not a;
    layer2_outputs(999) <= not a;
    layer2_outputs(1000) <= a and b;
    layer2_outputs(1001) <= not (a xor b);
    layer2_outputs(1002) <= not (a or b);
    layer2_outputs(1003) <= b and not a;
    layer2_outputs(1004) <= b;
    layer2_outputs(1005) <= not b;
    layer2_outputs(1006) <= not (a and b);
    layer2_outputs(1007) <= a;
    layer2_outputs(1008) <= '1';
    layer2_outputs(1009) <= '1';
    layer2_outputs(1010) <= not b;
    layer2_outputs(1011) <= a;
    layer2_outputs(1012) <= '0';
    layer2_outputs(1013) <= not (a xor b);
    layer2_outputs(1014) <= b;
    layer2_outputs(1015) <= not a;
    layer2_outputs(1016) <= a and not b;
    layer2_outputs(1017) <= not (a and b);
    layer2_outputs(1018) <= a or b;
    layer2_outputs(1019) <= not b;
    layer2_outputs(1020) <= not a or b;
    layer2_outputs(1021) <= not a;
    layer2_outputs(1022) <= '1';
    layer2_outputs(1023) <= '0';
    layer2_outputs(1024) <= not (a and b);
    layer2_outputs(1025) <= b and not a;
    layer2_outputs(1026) <= not b or a;
    layer2_outputs(1027) <= not a or b;
    layer2_outputs(1028) <= not b or a;
    layer2_outputs(1029) <= b;
    layer2_outputs(1030) <= not a or b;
    layer2_outputs(1031) <= not (a xor b);
    layer2_outputs(1032) <= '0';
    layer2_outputs(1033) <= a or b;
    layer2_outputs(1034) <= a;
    layer2_outputs(1035) <= not b or a;
    layer2_outputs(1036) <= not b or a;
    layer2_outputs(1037) <= not a;
    layer2_outputs(1038) <= '0';
    layer2_outputs(1039) <= not b or a;
    layer2_outputs(1040) <= '1';
    layer2_outputs(1041) <= not b or a;
    layer2_outputs(1042) <= a and b;
    layer2_outputs(1043) <= a or b;
    layer2_outputs(1044) <= not (a or b);
    layer2_outputs(1045) <= b and not a;
    layer2_outputs(1046) <= b and not a;
    layer2_outputs(1047) <= b;
    layer2_outputs(1048) <= not a or b;
    layer2_outputs(1049) <= not b or a;
    layer2_outputs(1050) <= a and b;
    layer2_outputs(1051) <= b;
    layer2_outputs(1052) <= not a or b;
    layer2_outputs(1053) <= not b;
    layer2_outputs(1054) <= not b;
    layer2_outputs(1055) <= not (a or b);
    layer2_outputs(1056) <= not b;
    layer2_outputs(1057) <= not (a xor b);
    layer2_outputs(1058) <= not (a and b);
    layer2_outputs(1059) <= '0';
    layer2_outputs(1060) <= b and not a;
    layer2_outputs(1061) <= a and b;
    layer2_outputs(1062) <= b;
    layer2_outputs(1063) <= '1';
    layer2_outputs(1064) <= b and not a;
    layer2_outputs(1065) <= b;
    layer2_outputs(1066) <= not (a or b);
    layer2_outputs(1067) <= b;
    layer2_outputs(1068) <= not (a and b);
    layer2_outputs(1069) <= not b;
    layer2_outputs(1070) <= a or b;
    layer2_outputs(1071) <= a xor b;
    layer2_outputs(1072) <= a and not b;
    layer2_outputs(1073) <= a xor b;
    layer2_outputs(1074) <= '0';
    layer2_outputs(1075) <= not a or b;
    layer2_outputs(1076) <= a xor b;
    layer2_outputs(1077) <= a and not b;
    layer2_outputs(1078) <= not b or a;
    layer2_outputs(1079) <= '0';
    layer2_outputs(1080) <= not a;
    layer2_outputs(1081) <= a and b;
    layer2_outputs(1082) <= a and not b;
    layer2_outputs(1083) <= a and b;
    layer2_outputs(1084) <= not a;
    layer2_outputs(1085) <= b and not a;
    layer2_outputs(1086) <= b;
    layer2_outputs(1087) <= a and not b;
    layer2_outputs(1088) <= not b;
    layer2_outputs(1089) <= not (a xor b);
    layer2_outputs(1090) <= '0';
    layer2_outputs(1091) <= b and not a;
    layer2_outputs(1092) <= a;
    layer2_outputs(1093) <= not (a or b);
    layer2_outputs(1094) <= not (a or b);
    layer2_outputs(1095) <= a and b;
    layer2_outputs(1096) <= '0';
    layer2_outputs(1097) <= '1';
    layer2_outputs(1098) <= '0';
    layer2_outputs(1099) <= not b;
    layer2_outputs(1100) <= a and not b;
    layer2_outputs(1101) <= b;
    layer2_outputs(1102) <= a or b;
    layer2_outputs(1103) <= not b;
    layer2_outputs(1104) <= b;
    layer2_outputs(1105) <= not b;
    layer2_outputs(1106) <= not (a or b);
    layer2_outputs(1107) <= a and not b;
    layer2_outputs(1108) <= not a or b;
    layer2_outputs(1109) <= not (a or b);
    layer2_outputs(1110) <= not (a or b);
    layer2_outputs(1111) <= a;
    layer2_outputs(1112) <= b and not a;
    layer2_outputs(1113) <= '1';
    layer2_outputs(1114) <= '0';
    layer2_outputs(1115) <= a;
    layer2_outputs(1116) <= not a;
    layer2_outputs(1117) <= a and not b;
    layer2_outputs(1118) <= not (a and b);
    layer2_outputs(1119) <= '0';
    layer2_outputs(1120) <= b;
    layer2_outputs(1121) <= not (a and b);
    layer2_outputs(1122) <= b and not a;
    layer2_outputs(1123) <= b;
    layer2_outputs(1124) <= a and not b;
    layer2_outputs(1125) <= b and not a;
    layer2_outputs(1126) <= not a or b;
    layer2_outputs(1127) <= '1';
    layer2_outputs(1128) <= '1';
    layer2_outputs(1129) <= not (a or b);
    layer2_outputs(1130) <= a or b;
    layer2_outputs(1131) <= b;
    layer2_outputs(1132) <= not b or a;
    layer2_outputs(1133) <= '1';
    layer2_outputs(1134) <= a xor b;
    layer2_outputs(1135) <= a and b;
    layer2_outputs(1136) <= not b or a;
    layer2_outputs(1137) <= b and not a;
    layer2_outputs(1138) <= a or b;
    layer2_outputs(1139) <= not a or b;
    layer2_outputs(1140) <= not (a and b);
    layer2_outputs(1141) <= a and b;
    layer2_outputs(1142) <= a and b;
    layer2_outputs(1143) <= not a or b;
    layer2_outputs(1144) <= not a;
    layer2_outputs(1145) <= a and b;
    layer2_outputs(1146) <= not (a xor b);
    layer2_outputs(1147) <= not (a or b);
    layer2_outputs(1148) <= a or b;
    layer2_outputs(1149) <= a and b;
    layer2_outputs(1150) <= '0';
    layer2_outputs(1151) <= a and b;
    layer2_outputs(1152) <= '0';
    layer2_outputs(1153) <= b and not a;
    layer2_outputs(1154) <= not a or b;
    layer2_outputs(1155) <= a or b;
    layer2_outputs(1156) <= a and not b;
    layer2_outputs(1157) <= a;
    layer2_outputs(1158) <= '1';
    layer2_outputs(1159) <= not (a and b);
    layer2_outputs(1160) <= b;
    layer2_outputs(1161) <= not a;
    layer2_outputs(1162) <= b and not a;
    layer2_outputs(1163) <= not a or b;
    layer2_outputs(1164) <= not (a and b);
    layer2_outputs(1165) <= not (a or b);
    layer2_outputs(1166) <= '1';
    layer2_outputs(1167) <= a and b;
    layer2_outputs(1168) <= a or b;
    layer2_outputs(1169) <= a and b;
    layer2_outputs(1170) <= not b or a;
    layer2_outputs(1171) <= '1';
    layer2_outputs(1172) <= not b;
    layer2_outputs(1173) <= a or b;
    layer2_outputs(1174) <= not b;
    layer2_outputs(1175) <= not (a xor b);
    layer2_outputs(1176) <= a and not b;
    layer2_outputs(1177) <= not (a or b);
    layer2_outputs(1178) <= not (a or b);
    layer2_outputs(1179) <= b;
    layer2_outputs(1180) <= not (a xor b);
    layer2_outputs(1181) <= not (a or b);
    layer2_outputs(1182) <= not b or a;
    layer2_outputs(1183) <= a and not b;
    layer2_outputs(1184) <= '0';
    layer2_outputs(1185) <= '0';
    layer2_outputs(1186) <= '0';
    layer2_outputs(1187) <= not a or b;
    layer2_outputs(1188) <= not (a or b);
    layer2_outputs(1189) <= not a or b;
    layer2_outputs(1190) <= a or b;
    layer2_outputs(1191) <= b and not a;
    layer2_outputs(1192) <= b and not a;
    layer2_outputs(1193) <= a;
    layer2_outputs(1194) <= a;
    layer2_outputs(1195) <= not b or a;
    layer2_outputs(1196) <= '0';
    layer2_outputs(1197) <= '1';
    layer2_outputs(1198) <= a and not b;
    layer2_outputs(1199) <= b and not a;
    layer2_outputs(1200) <= not (a and b);
    layer2_outputs(1201) <= not a;
    layer2_outputs(1202) <= a xor b;
    layer2_outputs(1203) <= a or b;
    layer2_outputs(1204) <= a;
    layer2_outputs(1205) <= a;
    layer2_outputs(1206) <= not b;
    layer2_outputs(1207) <= a and not b;
    layer2_outputs(1208) <= not a or b;
    layer2_outputs(1209) <= '1';
    layer2_outputs(1210) <= a;
    layer2_outputs(1211) <= not (a or b);
    layer2_outputs(1212) <= a;
    layer2_outputs(1213) <= a;
    layer2_outputs(1214) <= '1';
    layer2_outputs(1215) <= a;
    layer2_outputs(1216) <= b;
    layer2_outputs(1217) <= not a or b;
    layer2_outputs(1218) <= a and not b;
    layer2_outputs(1219) <= a or b;
    layer2_outputs(1220) <= '1';
    layer2_outputs(1221) <= a;
    layer2_outputs(1222) <= '0';
    layer2_outputs(1223) <= not b or a;
    layer2_outputs(1224) <= a and not b;
    layer2_outputs(1225) <= not a or b;
    layer2_outputs(1226) <= not (a or b);
    layer2_outputs(1227) <= a;
    layer2_outputs(1228) <= a or b;
    layer2_outputs(1229) <= '1';
    layer2_outputs(1230) <= not (a xor b);
    layer2_outputs(1231) <= not b or a;
    layer2_outputs(1232) <= not b or a;
    layer2_outputs(1233) <= a and not b;
    layer2_outputs(1234) <= a xor b;
    layer2_outputs(1235) <= not a;
    layer2_outputs(1236) <= '0';
    layer2_outputs(1237) <= '1';
    layer2_outputs(1238) <= a or b;
    layer2_outputs(1239) <= '0';
    layer2_outputs(1240) <= not a;
    layer2_outputs(1241) <= not b;
    layer2_outputs(1242) <= not (a and b);
    layer2_outputs(1243) <= not a or b;
    layer2_outputs(1244) <= a and not b;
    layer2_outputs(1245) <= not b or a;
    layer2_outputs(1246) <= '0';
    layer2_outputs(1247) <= '1';
    layer2_outputs(1248) <= not b or a;
    layer2_outputs(1249) <= b;
    layer2_outputs(1250) <= a or b;
    layer2_outputs(1251) <= not (a and b);
    layer2_outputs(1252) <= b;
    layer2_outputs(1253) <= a and b;
    layer2_outputs(1254) <= a;
    layer2_outputs(1255) <= not b or a;
    layer2_outputs(1256) <= not (a and b);
    layer2_outputs(1257) <= b;
    layer2_outputs(1258) <= a or b;
    layer2_outputs(1259) <= a or b;
    layer2_outputs(1260) <= a;
    layer2_outputs(1261) <= a;
    layer2_outputs(1262) <= '1';
    layer2_outputs(1263) <= b and not a;
    layer2_outputs(1264) <= '1';
    layer2_outputs(1265) <= not (a and b);
    layer2_outputs(1266) <= not b or a;
    layer2_outputs(1267) <= not (a or b);
    layer2_outputs(1268) <= a or b;
    layer2_outputs(1269) <= a and not b;
    layer2_outputs(1270) <= a or b;
    layer2_outputs(1271) <= not (a or b);
    layer2_outputs(1272) <= a and not b;
    layer2_outputs(1273) <= b and not a;
    layer2_outputs(1274) <= not b or a;
    layer2_outputs(1275) <= not (a or b);
    layer2_outputs(1276) <= not a or b;
    layer2_outputs(1277) <= not b or a;
    layer2_outputs(1278) <= a xor b;
    layer2_outputs(1279) <= b and not a;
    layer2_outputs(1280) <= a;
    layer2_outputs(1281) <= a and not b;
    layer2_outputs(1282) <= not a;
    layer2_outputs(1283) <= not a or b;
    layer2_outputs(1284) <= '1';
    layer2_outputs(1285) <= not a;
    layer2_outputs(1286) <= not b;
    layer2_outputs(1287) <= b and not a;
    layer2_outputs(1288) <= a;
    layer2_outputs(1289) <= a and b;
    layer2_outputs(1290) <= not (a and b);
    layer2_outputs(1291) <= not (a and b);
    layer2_outputs(1292) <= not (a and b);
    layer2_outputs(1293) <= b and not a;
    layer2_outputs(1294) <= '0';
    layer2_outputs(1295) <= '0';
    layer2_outputs(1296) <= a and b;
    layer2_outputs(1297) <= not (a or b);
    layer2_outputs(1298) <= a or b;
    layer2_outputs(1299) <= not (a and b);
    layer2_outputs(1300) <= not a or b;
    layer2_outputs(1301) <= b;
    layer2_outputs(1302) <= b and not a;
    layer2_outputs(1303) <= '0';
    layer2_outputs(1304) <= a and not b;
    layer2_outputs(1305) <= not b;
    layer2_outputs(1306) <= a or b;
    layer2_outputs(1307) <= not (a or b);
    layer2_outputs(1308) <= '0';
    layer2_outputs(1309) <= not a;
    layer2_outputs(1310) <= a;
    layer2_outputs(1311) <= not (a or b);
    layer2_outputs(1312) <= not a or b;
    layer2_outputs(1313) <= a or b;
    layer2_outputs(1314) <= not a or b;
    layer2_outputs(1315) <= not (a and b);
    layer2_outputs(1316) <= not a or b;
    layer2_outputs(1317) <= a or b;
    layer2_outputs(1318) <= b;
    layer2_outputs(1319) <= not (a and b);
    layer2_outputs(1320) <= '0';
    layer2_outputs(1321) <= not a or b;
    layer2_outputs(1322) <= not a or b;
    layer2_outputs(1323) <= a;
    layer2_outputs(1324) <= '0';
    layer2_outputs(1325) <= not (a or b);
    layer2_outputs(1326) <= '1';
    layer2_outputs(1327) <= '1';
    layer2_outputs(1328) <= not a or b;
    layer2_outputs(1329) <= '1';
    layer2_outputs(1330) <= a or b;
    layer2_outputs(1331) <= not (a and b);
    layer2_outputs(1332) <= not a or b;
    layer2_outputs(1333) <= not (a or b);
    layer2_outputs(1334) <= not (a or b);
    layer2_outputs(1335) <= not b;
    layer2_outputs(1336) <= b;
    layer2_outputs(1337) <= a and b;
    layer2_outputs(1338) <= a or b;
    layer2_outputs(1339) <= a or b;
    layer2_outputs(1340) <= a;
    layer2_outputs(1341) <= not a;
    layer2_outputs(1342) <= a;
    layer2_outputs(1343) <= '1';
    layer2_outputs(1344) <= a and not b;
    layer2_outputs(1345) <= a;
    layer2_outputs(1346) <= a and not b;
    layer2_outputs(1347) <= not a or b;
    layer2_outputs(1348) <= a or b;
    layer2_outputs(1349) <= not a or b;
    layer2_outputs(1350) <= not a or b;
    layer2_outputs(1351) <= b and not a;
    layer2_outputs(1352) <= '1';
    layer2_outputs(1353) <= '1';
    layer2_outputs(1354) <= a or b;
    layer2_outputs(1355) <= not a;
    layer2_outputs(1356) <= not (a and b);
    layer2_outputs(1357) <= a and b;
    layer2_outputs(1358) <= a and not b;
    layer2_outputs(1359) <= b and not a;
    layer2_outputs(1360) <= a or b;
    layer2_outputs(1361) <= '0';
    layer2_outputs(1362) <= a;
    layer2_outputs(1363) <= '1';
    layer2_outputs(1364) <= a and not b;
    layer2_outputs(1365) <= a and b;
    layer2_outputs(1366) <= not a;
    layer2_outputs(1367) <= not b;
    layer2_outputs(1368) <= not (a or b);
    layer2_outputs(1369) <= not (a and b);
    layer2_outputs(1370) <= not b or a;
    layer2_outputs(1371) <= not a or b;
    layer2_outputs(1372) <= '0';
    layer2_outputs(1373) <= not b;
    layer2_outputs(1374) <= not a or b;
    layer2_outputs(1375) <= '1';
    layer2_outputs(1376) <= not (a and b);
    layer2_outputs(1377) <= a;
    layer2_outputs(1378) <= a or b;
    layer2_outputs(1379) <= a and b;
    layer2_outputs(1380) <= a or b;
    layer2_outputs(1381) <= a and not b;
    layer2_outputs(1382) <= b;
    layer2_outputs(1383) <= a and not b;
    layer2_outputs(1384) <= '1';
    layer2_outputs(1385) <= not (a xor b);
    layer2_outputs(1386) <= '1';
    layer2_outputs(1387) <= b;
    layer2_outputs(1388) <= a;
    layer2_outputs(1389) <= b and not a;
    layer2_outputs(1390) <= '0';
    layer2_outputs(1391) <= '1';
    layer2_outputs(1392) <= not b or a;
    layer2_outputs(1393) <= b and not a;
    layer2_outputs(1394) <= b and not a;
    layer2_outputs(1395) <= a and b;
    layer2_outputs(1396) <= a;
    layer2_outputs(1397) <= not b or a;
    layer2_outputs(1398) <= a and not b;
    layer2_outputs(1399) <= not a;
    layer2_outputs(1400) <= not (a and b);
    layer2_outputs(1401) <= '0';
    layer2_outputs(1402) <= a or b;
    layer2_outputs(1403) <= not a;
    layer2_outputs(1404) <= not (a and b);
    layer2_outputs(1405) <= not a;
    layer2_outputs(1406) <= a;
    layer2_outputs(1407) <= not a;
    layer2_outputs(1408) <= a and not b;
    layer2_outputs(1409) <= not a;
    layer2_outputs(1410) <= '1';
    layer2_outputs(1411) <= not a;
    layer2_outputs(1412) <= '1';
    layer2_outputs(1413) <= b;
    layer2_outputs(1414) <= a and not b;
    layer2_outputs(1415) <= not a;
    layer2_outputs(1416) <= b;
    layer2_outputs(1417) <= '0';
    layer2_outputs(1418) <= not b;
    layer2_outputs(1419) <= '1';
    layer2_outputs(1420) <= not a;
    layer2_outputs(1421) <= not a or b;
    layer2_outputs(1422) <= not a;
    layer2_outputs(1423) <= not a;
    layer2_outputs(1424) <= not b;
    layer2_outputs(1425) <= not (a and b);
    layer2_outputs(1426) <= '0';
    layer2_outputs(1427) <= a and not b;
    layer2_outputs(1428) <= '0';
    layer2_outputs(1429) <= '0';
    layer2_outputs(1430) <= '1';
    layer2_outputs(1431) <= not (a or b);
    layer2_outputs(1432) <= '1';
    layer2_outputs(1433) <= not a;
    layer2_outputs(1434) <= not (a or b);
    layer2_outputs(1435) <= a;
    layer2_outputs(1436) <= b;
    layer2_outputs(1437) <= b;
    layer2_outputs(1438) <= not b or a;
    layer2_outputs(1439) <= not (a xor b);
    layer2_outputs(1440) <= not b;
    layer2_outputs(1441) <= b and not a;
    layer2_outputs(1442) <= a or b;
    layer2_outputs(1443) <= b;
    layer2_outputs(1444) <= '1';
    layer2_outputs(1445) <= not a or b;
    layer2_outputs(1446) <= not b;
    layer2_outputs(1447) <= '1';
    layer2_outputs(1448) <= a or b;
    layer2_outputs(1449) <= not (a and b);
    layer2_outputs(1450) <= a and not b;
    layer2_outputs(1451) <= not (a or b);
    layer2_outputs(1452) <= not (a or b);
    layer2_outputs(1453) <= a or b;
    layer2_outputs(1454) <= not (a and b);
    layer2_outputs(1455) <= not a;
    layer2_outputs(1456) <= a and b;
    layer2_outputs(1457) <= a or b;
    layer2_outputs(1458) <= '0';
    layer2_outputs(1459) <= b;
    layer2_outputs(1460) <= not b;
    layer2_outputs(1461) <= '1';
    layer2_outputs(1462) <= a and b;
    layer2_outputs(1463) <= a;
    layer2_outputs(1464) <= a or b;
    layer2_outputs(1465) <= '1';
    layer2_outputs(1466) <= not (a and b);
    layer2_outputs(1467) <= '1';
    layer2_outputs(1468) <= '0';
    layer2_outputs(1469) <= a or b;
    layer2_outputs(1470) <= '0';
    layer2_outputs(1471) <= a and b;
    layer2_outputs(1472) <= not b;
    layer2_outputs(1473) <= '1';
    layer2_outputs(1474) <= '1';
    layer2_outputs(1475) <= a;
    layer2_outputs(1476) <= not a or b;
    layer2_outputs(1477) <= '1';
    layer2_outputs(1478) <= not a;
    layer2_outputs(1479) <= a;
    layer2_outputs(1480) <= not a or b;
    layer2_outputs(1481) <= '0';
    layer2_outputs(1482) <= a;
    layer2_outputs(1483) <= b and not a;
    layer2_outputs(1484) <= a and b;
    layer2_outputs(1485) <= not b or a;
    layer2_outputs(1486) <= not a;
    layer2_outputs(1487) <= a and not b;
    layer2_outputs(1488) <= not a;
    layer2_outputs(1489) <= not (a and b);
    layer2_outputs(1490) <= b and not a;
    layer2_outputs(1491) <= not (a or b);
    layer2_outputs(1492) <= '1';
    layer2_outputs(1493) <= a and not b;
    layer2_outputs(1494) <= not a;
    layer2_outputs(1495) <= a and not b;
    layer2_outputs(1496) <= not (a and b);
    layer2_outputs(1497) <= not b;
    layer2_outputs(1498) <= b;
    layer2_outputs(1499) <= '1';
    layer2_outputs(1500) <= a;
    layer2_outputs(1501) <= a;
    layer2_outputs(1502) <= not (a xor b);
    layer2_outputs(1503) <= not b;
    layer2_outputs(1504) <= not a;
    layer2_outputs(1505) <= a;
    layer2_outputs(1506) <= a and b;
    layer2_outputs(1507) <= '1';
    layer2_outputs(1508) <= not (a and b);
    layer2_outputs(1509) <= not (a and b);
    layer2_outputs(1510) <= '1';
    layer2_outputs(1511) <= '1';
    layer2_outputs(1512) <= not b;
    layer2_outputs(1513) <= not a;
    layer2_outputs(1514) <= b and not a;
    layer2_outputs(1515) <= not b;
    layer2_outputs(1516) <= not b or a;
    layer2_outputs(1517) <= not b;
    layer2_outputs(1518) <= not b or a;
    layer2_outputs(1519) <= '0';
    layer2_outputs(1520) <= '0';
    layer2_outputs(1521) <= a or b;
    layer2_outputs(1522) <= a or b;
    layer2_outputs(1523) <= a;
    layer2_outputs(1524) <= not b or a;
    layer2_outputs(1525) <= a and b;
    layer2_outputs(1526) <= not a or b;
    layer2_outputs(1527) <= a or b;
    layer2_outputs(1528) <= a and not b;
    layer2_outputs(1529) <= b;
    layer2_outputs(1530) <= not (a and b);
    layer2_outputs(1531) <= not b or a;
    layer2_outputs(1532) <= not a;
    layer2_outputs(1533) <= not (a and b);
    layer2_outputs(1534) <= not b or a;
    layer2_outputs(1535) <= not a;
    layer2_outputs(1536) <= '0';
    layer2_outputs(1537) <= a and b;
    layer2_outputs(1538) <= '0';
    layer2_outputs(1539) <= not (a and b);
    layer2_outputs(1540) <= not (a xor b);
    layer2_outputs(1541) <= not b or a;
    layer2_outputs(1542) <= not (a and b);
    layer2_outputs(1543) <= a;
    layer2_outputs(1544) <= not b or a;
    layer2_outputs(1545) <= not (a or b);
    layer2_outputs(1546) <= not b;
    layer2_outputs(1547) <= '0';
    layer2_outputs(1548) <= a xor b;
    layer2_outputs(1549) <= b and not a;
    layer2_outputs(1550) <= a and b;
    layer2_outputs(1551) <= a xor b;
    layer2_outputs(1552) <= not a;
    layer2_outputs(1553) <= not (a xor b);
    layer2_outputs(1554) <= not b or a;
    layer2_outputs(1555) <= not a or b;
    layer2_outputs(1556) <= not (a and b);
    layer2_outputs(1557) <= not a;
    layer2_outputs(1558) <= not (a or b);
    layer2_outputs(1559) <= '0';
    layer2_outputs(1560) <= '0';
    layer2_outputs(1561) <= a;
    layer2_outputs(1562) <= '0';
    layer2_outputs(1563) <= a and b;
    layer2_outputs(1564) <= not (a and b);
    layer2_outputs(1565) <= b;
    layer2_outputs(1566) <= not b;
    layer2_outputs(1567) <= b and not a;
    layer2_outputs(1568) <= '1';
    layer2_outputs(1569) <= a;
    layer2_outputs(1570) <= a;
    layer2_outputs(1571) <= b;
    layer2_outputs(1572) <= not b or a;
    layer2_outputs(1573) <= not a;
    layer2_outputs(1574) <= not b;
    layer2_outputs(1575) <= not a or b;
    layer2_outputs(1576) <= b;
    layer2_outputs(1577) <= a and b;
    layer2_outputs(1578) <= b;
    layer2_outputs(1579) <= b;
    layer2_outputs(1580) <= a and b;
    layer2_outputs(1581) <= a or b;
    layer2_outputs(1582) <= not b;
    layer2_outputs(1583) <= not a or b;
    layer2_outputs(1584) <= not b or a;
    layer2_outputs(1585) <= not (a and b);
    layer2_outputs(1586) <= '0';
    layer2_outputs(1587) <= a xor b;
    layer2_outputs(1588) <= a and b;
    layer2_outputs(1589) <= '1';
    layer2_outputs(1590) <= not (a or b);
    layer2_outputs(1591) <= a or b;
    layer2_outputs(1592) <= not (a or b);
    layer2_outputs(1593) <= not a or b;
    layer2_outputs(1594) <= b;
    layer2_outputs(1595) <= b and not a;
    layer2_outputs(1596) <= a;
    layer2_outputs(1597) <= not (a or b);
    layer2_outputs(1598) <= a and b;
    layer2_outputs(1599) <= '1';
    layer2_outputs(1600) <= not b;
    layer2_outputs(1601) <= a xor b;
    layer2_outputs(1602) <= not b;
    layer2_outputs(1603) <= not (a or b);
    layer2_outputs(1604) <= a;
    layer2_outputs(1605) <= a and not b;
    layer2_outputs(1606) <= not b or a;
    layer2_outputs(1607) <= '1';
    layer2_outputs(1608) <= a;
    layer2_outputs(1609) <= not (a and b);
    layer2_outputs(1610) <= b and not a;
    layer2_outputs(1611) <= '1';
    layer2_outputs(1612) <= b;
    layer2_outputs(1613) <= not a or b;
    layer2_outputs(1614) <= not a;
    layer2_outputs(1615) <= not (a or b);
    layer2_outputs(1616) <= not a;
    layer2_outputs(1617) <= not b or a;
    layer2_outputs(1618) <= not (a and b);
    layer2_outputs(1619) <= a;
    layer2_outputs(1620) <= a and b;
    layer2_outputs(1621) <= a;
    layer2_outputs(1622) <= '0';
    layer2_outputs(1623) <= a and not b;
    layer2_outputs(1624) <= not a or b;
    layer2_outputs(1625) <= b;
    layer2_outputs(1626) <= not (a or b);
    layer2_outputs(1627) <= '1';
    layer2_outputs(1628) <= a;
    layer2_outputs(1629) <= a or b;
    layer2_outputs(1630) <= a;
    layer2_outputs(1631) <= not a or b;
    layer2_outputs(1632) <= a or b;
    layer2_outputs(1633) <= b and not a;
    layer2_outputs(1634) <= not (a or b);
    layer2_outputs(1635) <= not b or a;
    layer2_outputs(1636) <= a;
    layer2_outputs(1637) <= a or b;
    layer2_outputs(1638) <= '1';
    layer2_outputs(1639) <= b and not a;
    layer2_outputs(1640) <= a and b;
    layer2_outputs(1641) <= '1';
    layer2_outputs(1642) <= '1';
    layer2_outputs(1643) <= b;
    layer2_outputs(1644) <= a and b;
    layer2_outputs(1645) <= a and not b;
    layer2_outputs(1646) <= a and b;
    layer2_outputs(1647) <= a or b;
    layer2_outputs(1648) <= not b or a;
    layer2_outputs(1649) <= b and not a;
    layer2_outputs(1650) <= not a or b;
    layer2_outputs(1651) <= b and not a;
    layer2_outputs(1652) <= not (a xor b);
    layer2_outputs(1653) <= not a;
    layer2_outputs(1654) <= not b;
    layer2_outputs(1655) <= not a or b;
    layer2_outputs(1656) <= a and not b;
    layer2_outputs(1657) <= '1';
    layer2_outputs(1658) <= not b or a;
    layer2_outputs(1659) <= '1';
    layer2_outputs(1660) <= not b;
    layer2_outputs(1661) <= not b or a;
    layer2_outputs(1662) <= a and not b;
    layer2_outputs(1663) <= a;
    layer2_outputs(1664) <= b and not a;
    layer2_outputs(1665) <= a or b;
    layer2_outputs(1666) <= not b;
    layer2_outputs(1667) <= b and not a;
    layer2_outputs(1668) <= a and b;
    layer2_outputs(1669) <= a;
    layer2_outputs(1670) <= not (a or b);
    layer2_outputs(1671) <= not (a or b);
    layer2_outputs(1672) <= '0';
    layer2_outputs(1673) <= not (a or b);
    layer2_outputs(1674) <= not a;
    layer2_outputs(1675) <= a and not b;
    layer2_outputs(1676) <= a xor b;
    layer2_outputs(1677) <= a or b;
    layer2_outputs(1678) <= not (a and b);
    layer2_outputs(1679) <= not b or a;
    layer2_outputs(1680) <= not (a or b);
    layer2_outputs(1681) <= a or b;
    layer2_outputs(1682) <= b and not a;
    layer2_outputs(1683) <= not b;
    layer2_outputs(1684) <= a and b;
    layer2_outputs(1685) <= not b;
    layer2_outputs(1686) <= '0';
    layer2_outputs(1687) <= not b or a;
    layer2_outputs(1688) <= a or b;
    layer2_outputs(1689) <= not b or a;
    layer2_outputs(1690) <= not a or b;
    layer2_outputs(1691) <= b;
    layer2_outputs(1692) <= a or b;
    layer2_outputs(1693) <= a;
    layer2_outputs(1694) <= '1';
    layer2_outputs(1695) <= not (a or b);
    layer2_outputs(1696) <= not (a and b);
    layer2_outputs(1697) <= not (a or b);
    layer2_outputs(1698) <= not a;
    layer2_outputs(1699) <= '1';
    layer2_outputs(1700) <= b;
    layer2_outputs(1701) <= not b;
    layer2_outputs(1702) <= not b;
    layer2_outputs(1703) <= b;
    layer2_outputs(1704) <= a or b;
    layer2_outputs(1705) <= a and b;
    layer2_outputs(1706) <= '1';
    layer2_outputs(1707) <= not b;
    layer2_outputs(1708) <= not a or b;
    layer2_outputs(1709) <= not a;
    layer2_outputs(1710) <= not a;
    layer2_outputs(1711) <= not a;
    layer2_outputs(1712) <= not a or b;
    layer2_outputs(1713) <= a and b;
    layer2_outputs(1714) <= b;
    layer2_outputs(1715) <= a and b;
    layer2_outputs(1716) <= a;
    layer2_outputs(1717) <= not b or a;
    layer2_outputs(1718) <= a or b;
    layer2_outputs(1719) <= not (a and b);
    layer2_outputs(1720) <= '1';
    layer2_outputs(1721) <= not (a and b);
    layer2_outputs(1722) <= a;
    layer2_outputs(1723) <= a;
    layer2_outputs(1724) <= '1';
    layer2_outputs(1725) <= a and b;
    layer2_outputs(1726) <= not (a xor b);
    layer2_outputs(1727) <= not (a or b);
    layer2_outputs(1728) <= b;
    layer2_outputs(1729) <= a and not b;
    layer2_outputs(1730) <= b and not a;
    layer2_outputs(1731) <= not (a and b);
    layer2_outputs(1732) <= not a;
    layer2_outputs(1733) <= a;
    layer2_outputs(1734) <= a;
    layer2_outputs(1735) <= a and not b;
    layer2_outputs(1736) <= '0';
    layer2_outputs(1737) <= a and b;
    layer2_outputs(1738) <= a;
    layer2_outputs(1739) <= '0';
    layer2_outputs(1740) <= '0';
    layer2_outputs(1741) <= not a;
    layer2_outputs(1742) <= not (a and b);
    layer2_outputs(1743) <= not a or b;
    layer2_outputs(1744) <= b and not a;
    layer2_outputs(1745) <= not b or a;
    layer2_outputs(1746) <= a xor b;
    layer2_outputs(1747) <= '0';
    layer2_outputs(1748) <= '1';
    layer2_outputs(1749) <= not (a and b);
    layer2_outputs(1750) <= b and not a;
    layer2_outputs(1751) <= '0';
    layer2_outputs(1752) <= not b;
    layer2_outputs(1753) <= not (a and b);
    layer2_outputs(1754) <= a and b;
    layer2_outputs(1755) <= not (a or b);
    layer2_outputs(1756) <= not (a and b);
    layer2_outputs(1757) <= not b or a;
    layer2_outputs(1758) <= '1';
    layer2_outputs(1759) <= a and b;
    layer2_outputs(1760) <= not (a and b);
    layer2_outputs(1761) <= b and not a;
    layer2_outputs(1762) <= a or b;
    layer2_outputs(1763) <= not (a or b);
    layer2_outputs(1764) <= not a or b;
    layer2_outputs(1765) <= '0';
    layer2_outputs(1766) <= a and b;
    layer2_outputs(1767) <= a and not b;
    layer2_outputs(1768) <= a;
    layer2_outputs(1769) <= a and not b;
    layer2_outputs(1770) <= a;
    layer2_outputs(1771) <= '1';
    layer2_outputs(1772) <= a xor b;
    layer2_outputs(1773) <= b;
    layer2_outputs(1774) <= not (a or b);
    layer2_outputs(1775) <= a or b;
    layer2_outputs(1776) <= not (a and b);
    layer2_outputs(1777) <= not a;
    layer2_outputs(1778) <= a;
    layer2_outputs(1779) <= b;
    layer2_outputs(1780) <= '1';
    layer2_outputs(1781) <= b and not a;
    layer2_outputs(1782) <= a;
    layer2_outputs(1783) <= '0';
    layer2_outputs(1784) <= not (a and b);
    layer2_outputs(1785) <= b and not a;
    layer2_outputs(1786) <= '1';
    layer2_outputs(1787) <= '1';
    layer2_outputs(1788) <= not a;
    layer2_outputs(1789) <= not b;
    layer2_outputs(1790) <= a and b;
    layer2_outputs(1791) <= not a;
    layer2_outputs(1792) <= a;
    layer2_outputs(1793) <= b;
    layer2_outputs(1794) <= not b or a;
    layer2_outputs(1795) <= b;
    layer2_outputs(1796) <= b;
    layer2_outputs(1797) <= a and not b;
    layer2_outputs(1798) <= not (a or b);
    layer2_outputs(1799) <= a and b;
    layer2_outputs(1800) <= a and not b;
    layer2_outputs(1801) <= not a;
    layer2_outputs(1802) <= not a or b;
    layer2_outputs(1803) <= '0';
    layer2_outputs(1804) <= not a or b;
    layer2_outputs(1805) <= a;
    layer2_outputs(1806) <= a;
    layer2_outputs(1807) <= a or b;
    layer2_outputs(1808) <= not b or a;
    layer2_outputs(1809) <= a xor b;
    layer2_outputs(1810) <= not (a and b);
    layer2_outputs(1811) <= not b or a;
    layer2_outputs(1812) <= a and b;
    layer2_outputs(1813) <= '1';
    layer2_outputs(1814) <= b;
    layer2_outputs(1815) <= a or b;
    layer2_outputs(1816) <= a and b;
    layer2_outputs(1817) <= a or b;
    layer2_outputs(1818) <= '0';
    layer2_outputs(1819) <= not (a and b);
    layer2_outputs(1820) <= not (a or b);
    layer2_outputs(1821) <= not (a xor b);
    layer2_outputs(1822) <= a;
    layer2_outputs(1823) <= not b;
    layer2_outputs(1824) <= '0';
    layer2_outputs(1825) <= a or b;
    layer2_outputs(1826) <= not a;
    layer2_outputs(1827) <= a;
    layer2_outputs(1828) <= '1';
    layer2_outputs(1829) <= '1';
    layer2_outputs(1830) <= a or b;
    layer2_outputs(1831) <= b and not a;
    layer2_outputs(1832) <= a and b;
    layer2_outputs(1833) <= '0';
    layer2_outputs(1834) <= '1';
    layer2_outputs(1835) <= a xor b;
    layer2_outputs(1836) <= '1';
    layer2_outputs(1837) <= a and b;
    layer2_outputs(1838) <= a and b;
    layer2_outputs(1839) <= a and b;
    layer2_outputs(1840) <= b;
    layer2_outputs(1841) <= b;
    layer2_outputs(1842) <= b and not a;
    layer2_outputs(1843) <= not (a and b);
    layer2_outputs(1844) <= '1';
    layer2_outputs(1845) <= not a;
    layer2_outputs(1846) <= not b or a;
    layer2_outputs(1847) <= not (a and b);
    layer2_outputs(1848) <= not a;
    layer2_outputs(1849) <= b;
    layer2_outputs(1850) <= not (a and b);
    layer2_outputs(1851) <= '0';
    layer2_outputs(1852) <= '0';
    layer2_outputs(1853) <= '1';
    layer2_outputs(1854) <= '1';
    layer2_outputs(1855) <= not a;
    layer2_outputs(1856) <= a and b;
    layer2_outputs(1857) <= '0';
    layer2_outputs(1858) <= a and not b;
    layer2_outputs(1859) <= not b;
    layer2_outputs(1860) <= a;
    layer2_outputs(1861) <= b and not a;
    layer2_outputs(1862) <= a;
    layer2_outputs(1863) <= b;
    layer2_outputs(1864) <= b and not a;
    layer2_outputs(1865) <= a;
    layer2_outputs(1866) <= a;
    layer2_outputs(1867) <= '1';
    layer2_outputs(1868) <= not b;
    layer2_outputs(1869) <= b;
    layer2_outputs(1870) <= not a;
    layer2_outputs(1871) <= a;
    layer2_outputs(1872) <= a and not b;
    layer2_outputs(1873) <= not a or b;
    layer2_outputs(1874) <= not a or b;
    layer2_outputs(1875) <= a and b;
    layer2_outputs(1876) <= not a;
    layer2_outputs(1877) <= a or b;
    layer2_outputs(1878) <= '1';
    layer2_outputs(1879) <= not (a and b);
    layer2_outputs(1880) <= '0';
    layer2_outputs(1881) <= not a;
    layer2_outputs(1882) <= '0';
    layer2_outputs(1883) <= '1';
    layer2_outputs(1884) <= a and not b;
    layer2_outputs(1885) <= not b;
    layer2_outputs(1886) <= a and not b;
    layer2_outputs(1887) <= not (a and b);
    layer2_outputs(1888) <= '1';
    layer2_outputs(1889) <= b and not a;
    layer2_outputs(1890) <= a or b;
    layer2_outputs(1891) <= a and b;
    layer2_outputs(1892) <= not a or b;
    layer2_outputs(1893) <= not (a and b);
    layer2_outputs(1894) <= not (a and b);
    layer2_outputs(1895) <= b and not a;
    layer2_outputs(1896) <= not a or b;
    layer2_outputs(1897) <= not (a and b);
    layer2_outputs(1898) <= not a;
    layer2_outputs(1899) <= not b or a;
    layer2_outputs(1900) <= not a or b;
    layer2_outputs(1901) <= a or b;
    layer2_outputs(1902) <= '0';
    layer2_outputs(1903) <= a or b;
    layer2_outputs(1904) <= '0';
    layer2_outputs(1905) <= '1';
    layer2_outputs(1906) <= a and not b;
    layer2_outputs(1907) <= not a;
    layer2_outputs(1908) <= not a;
    layer2_outputs(1909) <= a;
    layer2_outputs(1910) <= not a or b;
    layer2_outputs(1911) <= b and not a;
    layer2_outputs(1912) <= b;
    layer2_outputs(1913) <= not (a and b);
    layer2_outputs(1914) <= not b or a;
    layer2_outputs(1915) <= not b or a;
    layer2_outputs(1916) <= a and b;
    layer2_outputs(1917) <= not (a and b);
    layer2_outputs(1918) <= not (a and b);
    layer2_outputs(1919) <= not (a and b);
    layer2_outputs(1920) <= not (a xor b);
    layer2_outputs(1921) <= '0';
    layer2_outputs(1922) <= a xor b;
    layer2_outputs(1923) <= not a or b;
    layer2_outputs(1924) <= '0';
    layer2_outputs(1925) <= not b or a;
    layer2_outputs(1926) <= b and not a;
    layer2_outputs(1927) <= b;
    layer2_outputs(1928) <= '0';
    layer2_outputs(1929) <= not (a or b);
    layer2_outputs(1930) <= not a;
    layer2_outputs(1931) <= '0';
    layer2_outputs(1932) <= b and not a;
    layer2_outputs(1933) <= not a or b;
    layer2_outputs(1934) <= a or b;
    layer2_outputs(1935) <= not b or a;
    layer2_outputs(1936) <= not (a and b);
    layer2_outputs(1937) <= a and not b;
    layer2_outputs(1938) <= '1';
    layer2_outputs(1939) <= not b or a;
    layer2_outputs(1940) <= b and not a;
    layer2_outputs(1941) <= not b or a;
    layer2_outputs(1942) <= a xor b;
    layer2_outputs(1943) <= not b or a;
    layer2_outputs(1944) <= a and b;
    layer2_outputs(1945) <= not b;
    layer2_outputs(1946) <= a and not b;
    layer2_outputs(1947) <= b and not a;
    layer2_outputs(1948) <= not (a and b);
    layer2_outputs(1949) <= b;
    layer2_outputs(1950) <= a and not b;
    layer2_outputs(1951) <= a;
    layer2_outputs(1952) <= '0';
    layer2_outputs(1953) <= not b;
    layer2_outputs(1954) <= b and not a;
    layer2_outputs(1955) <= '0';
    layer2_outputs(1956) <= not (a and b);
    layer2_outputs(1957) <= a or b;
    layer2_outputs(1958) <= not (a or b);
    layer2_outputs(1959) <= not a;
    layer2_outputs(1960) <= not b or a;
    layer2_outputs(1961) <= b and not a;
    layer2_outputs(1962) <= not (a or b);
    layer2_outputs(1963) <= not (a or b);
    layer2_outputs(1964) <= a and b;
    layer2_outputs(1965) <= not (a or b);
    layer2_outputs(1966) <= b;
    layer2_outputs(1967) <= b;
    layer2_outputs(1968) <= '0';
    layer2_outputs(1969) <= '1';
    layer2_outputs(1970) <= not b;
    layer2_outputs(1971) <= b and not a;
    layer2_outputs(1972) <= a and b;
    layer2_outputs(1973) <= a or b;
    layer2_outputs(1974) <= not b;
    layer2_outputs(1975) <= not a or b;
    layer2_outputs(1976) <= '1';
    layer2_outputs(1977) <= not a;
    layer2_outputs(1978) <= a;
    layer2_outputs(1979) <= not a;
    layer2_outputs(1980) <= b and not a;
    layer2_outputs(1981) <= not (a and b);
    layer2_outputs(1982) <= a;
    layer2_outputs(1983) <= a;
    layer2_outputs(1984) <= not b or a;
    layer2_outputs(1985) <= b;
    layer2_outputs(1986) <= '1';
    layer2_outputs(1987) <= b;
    layer2_outputs(1988) <= a;
    layer2_outputs(1989) <= a or b;
    layer2_outputs(1990) <= not (a and b);
    layer2_outputs(1991) <= '1';
    layer2_outputs(1992) <= not a;
    layer2_outputs(1993) <= not b;
    layer2_outputs(1994) <= '0';
    layer2_outputs(1995) <= not b;
    layer2_outputs(1996) <= b and not a;
    layer2_outputs(1997) <= not a or b;
    layer2_outputs(1998) <= a and not b;
    layer2_outputs(1999) <= not a;
    layer2_outputs(2000) <= a and not b;
    layer2_outputs(2001) <= not a or b;
    layer2_outputs(2002) <= '0';
    layer2_outputs(2003) <= not (a and b);
    layer2_outputs(2004) <= not (a or b);
    layer2_outputs(2005) <= not (a or b);
    layer2_outputs(2006) <= not a or b;
    layer2_outputs(2007) <= a or b;
    layer2_outputs(2008) <= not (a and b);
    layer2_outputs(2009) <= b and not a;
    layer2_outputs(2010) <= not (a and b);
    layer2_outputs(2011) <= not b;
    layer2_outputs(2012) <= not (a and b);
    layer2_outputs(2013) <= '0';
    layer2_outputs(2014) <= not a or b;
    layer2_outputs(2015) <= not a or b;
    layer2_outputs(2016) <= not a;
    layer2_outputs(2017) <= a and not b;
    layer2_outputs(2018) <= not (a and b);
    layer2_outputs(2019) <= a and b;
    layer2_outputs(2020) <= '0';
    layer2_outputs(2021) <= '0';
    layer2_outputs(2022) <= '1';
    layer2_outputs(2023) <= not (a xor b);
    layer2_outputs(2024) <= not a or b;
    layer2_outputs(2025) <= a and b;
    layer2_outputs(2026) <= not a;
    layer2_outputs(2027) <= not a or b;
    layer2_outputs(2028) <= a or b;
    layer2_outputs(2029) <= not (a and b);
    layer2_outputs(2030) <= a and not b;
    layer2_outputs(2031) <= b;
    layer2_outputs(2032) <= '1';
    layer2_outputs(2033) <= '0';
    layer2_outputs(2034) <= a or b;
    layer2_outputs(2035) <= not a or b;
    layer2_outputs(2036) <= not a or b;
    layer2_outputs(2037) <= not (a or b);
    layer2_outputs(2038) <= not b or a;
    layer2_outputs(2039) <= b and not a;
    layer2_outputs(2040) <= a;
    layer2_outputs(2041) <= a;
    layer2_outputs(2042) <= a and b;
    layer2_outputs(2043) <= '0';
    layer2_outputs(2044) <= b;
    layer2_outputs(2045) <= a or b;
    layer2_outputs(2046) <= not a;
    layer2_outputs(2047) <= not (a or b);
    layer2_outputs(2048) <= '1';
    layer2_outputs(2049) <= not (a and b);
    layer2_outputs(2050) <= '0';
    layer2_outputs(2051) <= b;
    layer2_outputs(2052) <= '1';
    layer2_outputs(2053) <= b;
    layer2_outputs(2054) <= b;
    layer2_outputs(2055) <= not b;
    layer2_outputs(2056) <= not a;
    layer2_outputs(2057) <= b;
    layer2_outputs(2058) <= b;
    layer2_outputs(2059) <= '1';
    layer2_outputs(2060) <= not a;
    layer2_outputs(2061) <= not a or b;
    layer2_outputs(2062) <= b and not a;
    layer2_outputs(2063) <= a and b;
    layer2_outputs(2064) <= not (a and b);
    layer2_outputs(2065) <= a or b;
    layer2_outputs(2066) <= '0';
    layer2_outputs(2067) <= not b;
    layer2_outputs(2068) <= a or b;
    layer2_outputs(2069) <= '0';
    layer2_outputs(2070) <= a or b;
    layer2_outputs(2071) <= b;
    layer2_outputs(2072) <= '0';
    layer2_outputs(2073) <= not a;
    layer2_outputs(2074) <= not a;
    layer2_outputs(2075) <= a;
    layer2_outputs(2076) <= a or b;
    layer2_outputs(2077) <= '0';
    layer2_outputs(2078) <= b and not a;
    layer2_outputs(2079) <= '0';
    layer2_outputs(2080) <= '1';
    layer2_outputs(2081) <= b;
    layer2_outputs(2082) <= '0';
    layer2_outputs(2083) <= '0';
    layer2_outputs(2084) <= a and not b;
    layer2_outputs(2085) <= not a or b;
    layer2_outputs(2086) <= a;
    layer2_outputs(2087) <= not b or a;
    layer2_outputs(2088) <= not b or a;
    layer2_outputs(2089) <= a or b;
    layer2_outputs(2090) <= not (a and b);
    layer2_outputs(2091) <= b;
    layer2_outputs(2092) <= a or b;
    layer2_outputs(2093) <= not b or a;
    layer2_outputs(2094) <= a or b;
    layer2_outputs(2095) <= a;
    layer2_outputs(2096) <= a;
    layer2_outputs(2097) <= b and not a;
    layer2_outputs(2098) <= not a or b;
    layer2_outputs(2099) <= a or b;
    layer2_outputs(2100) <= not a;
    layer2_outputs(2101) <= a and b;
    layer2_outputs(2102) <= a and not b;
    layer2_outputs(2103) <= b and not a;
    layer2_outputs(2104) <= b;
    layer2_outputs(2105) <= b and not a;
    layer2_outputs(2106) <= not (a or b);
    layer2_outputs(2107) <= a or b;
    layer2_outputs(2108) <= '1';
    layer2_outputs(2109) <= not (a and b);
    layer2_outputs(2110) <= '1';
    layer2_outputs(2111) <= not (a and b);
    layer2_outputs(2112) <= not b;
    layer2_outputs(2113) <= '1';
    layer2_outputs(2114) <= not a or b;
    layer2_outputs(2115) <= not b;
    layer2_outputs(2116) <= not b;
    layer2_outputs(2117) <= a and not b;
    layer2_outputs(2118) <= a or b;
    layer2_outputs(2119) <= '1';
    layer2_outputs(2120) <= '1';
    layer2_outputs(2121) <= a and not b;
    layer2_outputs(2122) <= a;
    layer2_outputs(2123) <= '0';
    layer2_outputs(2124) <= not (a and b);
    layer2_outputs(2125) <= b;
    layer2_outputs(2126) <= a xor b;
    layer2_outputs(2127) <= not b;
    layer2_outputs(2128) <= b and not a;
    layer2_outputs(2129) <= b and not a;
    layer2_outputs(2130) <= '1';
    layer2_outputs(2131) <= b;
    layer2_outputs(2132) <= not (a and b);
    layer2_outputs(2133) <= b;
    layer2_outputs(2134) <= '1';
    layer2_outputs(2135) <= not b or a;
    layer2_outputs(2136) <= not (a and b);
    layer2_outputs(2137) <= a;
    layer2_outputs(2138) <= b;
    layer2_outputs(2139) <= '0';
    layer2_outputs(2140) <= not a;
    layer2_outputs(2141) <= a;
    layer2_outputs(2142) <= not (a or b);
    layer2_outputs(2143) <= b;
    layer2_outputs(2144) <= not (a or b);
    layer2_outputs(2145) <= b and not a;
    layer2_outputs(2146) <= '1';
    layer2_outputs(2147) <= '0';
    layer2_outputs(2148) <= a or b;
    layer2_outputs(2149) <= a or b;
    layer2_outputs(2150) <= not a or b;
    layer2_outputs(2151) <= not b or a;
    layer2_outputs(2152) <= a or b;
    layer2_outputs(2153) <= not a or b;
    layer2_outputs(2154) <= a or b;
    layer2_outputs(2155) <= '1';
    layer2_outputs(2156) <= not b;
    layer2_outputs(2157) <= a and not b;
    layer2_outputs(2158) <= a;
    layer2_outputs(2159) <= not a or b;
    layer2_outputs(2160) <= not (a or b);
    layer2_outputs(2161) <= a and not b;
    layer2_outputs(2162) <= not b;
    layer2_outputs(2163) <= not b;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= '0';
    layer2_outputs(2166) <= a and not b;
    layer2_outputs(2167) <= b;
    layer2_outputs(2168) <= a xor b;
    layer2_outputs(2169) <= '1';
    layer2_outputs(2170) <= not b;
    layer2_outputs(2171) <= a or b;
    layer2_outputs(2172) <= not a or b;
    layer2_outputs(2173) <= b;
    layer2_outputs(2174) <= b and not a;
    layer2_outputs(2175) <= not (a or b);
    layer2_outputs(2176) <= a and not b;
    layer2_outputs(2177) <= not (a or b);
    layer2_outputs(2178) <= not a or b;
    layer2_outputs(2179) <= a;
    layer2_outputs(2180) <= not b or a;
    layer2_outputs(2181) <= not a;
    layer2_outputs(2182) <= a or b;
    layer2_outputs(2183) <= '0';
    layer2_outputs(2184) <= a;
    layer2_outputs(2185) <= not (a or b);
    layer2_outputs(2186) <= a and b;
    layer2_outputs(2187) <= not a;
    layer2_outputs(2188) <= b;
    layer2_outputs(2189) <= '1';
    layer2_outputs(2190) <= b and not a;
    layer2_outputs(2191) <= a and not b;
    layer2_outputs(2192) <= a and b;
    layer2_outputs(2193) <= '0';
    layer2_outputs(2194) <= b and not a;
    layer2_outputs(2195) <= '1';
    layer2_outputs(2196) <= not (a or b);
    layer2_outputs(2197) <= '1';
    layer2_outputs(2198) <= not (a and b);
    layer2_outputs(2199) <= b;
    layer2_outputs(2200) <= not (a and b);
    layer2_outputs(2201) <= not a or b;
    layer2_outputs(2202) <= not a or b;
    layer2_outputs(2203) <= b;
    layer2_outputs(2204) <= not (a and b);
    layer2_outputs(2205) <= '0';
    layer2_outputs(2206) <= b;
    layer2_outputs(2207) <= not b;
    layer2_outputs(2208) <= not (a and b);
    layer2_outputs(2209) <= '0';
    layer2_outputs(2210) <= b;
    layer2_outputs(2211) <= '1';
    layer2_outputs(2212) <= not a;
    layer2_outputs(2213) <= not a or b;
    layer2_outputs(2214) <= not a;
    layer2_outputs(2215) <= not a or b;
    layer2_outputs(2216) <= not a or b;
    layer2_outputs(2217) <= not b or a;
    layer2_outputs(2218) <= not b or a;
    layer2_outputs(2219) <= '0';
    layer2_outputs(2220) <= a;
    layer2_outputs(2221) <= a;
    layer2_outputs(2222) <= '1';
    layer2_outputs(2223) <= not a or b;
    layer2_outputs(2224) <= a;
    layer2_outputs(2225) <= a or b;
    layer2_outputs(2226) <= '0';
    layer2_outputs(2227) <= '0';
    layer2_outputs(2228) <= a and b;
    layer2_outputs(2229) <= a or b;
    layer2_outputs(2230) <= not b;
    layer2_outputs(2231) <= '0';
    layer2_outputs(2232) <= a or b;
    layer2_outputs(2233) <= not b or a;
    layer2_outputs(2234) <= not b or a;
    layer2_outputs(2235) <= b;
    layer2_outputs(2236) <= a or b;
    layer2_outputs(2237) <= a and not b;
    layer2_outputs(2238) <= a or b;
    layer2_outputs(2239) <= '1';
    layer2_outputs(2240) <= not b or a;
    layer2_outputs(2241) <= a and b;
    layer2_outputs(2242) <= not a;
    layer2_outputs(2243) <= '1';
    layer2_outputs(2244) <= a;
    layer2_outputs(2245) <= a or b;
    layer2_outputs(2246) <= a;
    layer2_outputs(2247) <= not b or a;
    layer2_outputs(2248) <= b and not a;
    layer2_outputs(2249) <= not b or a;
    layer2_outputs(2250) <= '1';
    layer2_outputs(2251) <= '0';
    layer2_outputs(2252) <= a and b;
    layer2_outputs(2253) <= a and b;
    layer2_outputs(2254) <= not (a or b);
    layer2_outputs(2255) <= not b or a;
    layer2_outputs(2256) <= not a or b;
    layer2_outputs(2257) <= '1';
    layer2_outputs(2258) <= a and not b;
    layer2_outputs(2259) <= not a;
    layer2_outputs(2260) <= a xor b;
    layer2_outputs(2261) <= b and not a;
    layer2_outputs(2262) <= '1';
    layer2_outputs(2263) <= not b;
    layer2_outputs(2264) <= not (a or b);
    layer2_outputs(2265) <= not a;
    layer2_outputs(2266) <= '0';
    layer2_outputs(2267) <= not (a xor b);
    layer2_outputs(2268) <= a or b;
    layer2_outputs(2269) <= not b or a;
    layer2_outputs(2270) <= '0';
    layer2_outputs(2271) <= a and not b;
    layer2_outputs(2272) <= not b;
    layer2_outputs(2273) <= not (a or b);
    layer2_outputs(2274) <= not a or b;
    layer2_outputs(2275) <= not b;
    layer2_outputs(2276) <= '1';
    layer2_outputs(2277) <= a or b;
    layer2_outputs(2278) <= '0';
    layer2_outputs(2279) <= a and not b;
    layer2_outputs(2280) <= a or b;
    layer2_outputs(2281) <= a or b;
    layer2_outputs(2282) <= not b;
    layer2_outputs(2283) <= not b;
    layer2_outputs(2284) <= a;
    layer2_outputs(2285) <= not (a or b);
    layer2_outputs(2286) <= '1';
    layer2_outputs(2287) <= b;
    layer2_outputs(2288) <= '1';
    layer2_outputs(2289) <= not (a and b);
    layer2_outputs(2290) <= b and not a;
    layer2_outputs(2291) <= not b;
    layer2_outputs(2292) <= not (a or b);
    layer2_outputs(2293) <= not b;
    layer2_outputs(2294) <= not b;
    layer2_outputs(2295) <= a or b;
    layer2_outputs(2296) <= a or b;
    layer2_outputs(2297) <= '0';
    layer2_outputs(2298) <= b and not a;
    layer2_outputs(2299) <= not (a and b);
    layer2_outputs(2300) <= a or b;
    layer2_outputs(2301) <= '0';
    layer2_outputs(2302) <= '0';
    layer2_outputs(2303) <= not a or b;
    layer2_outputs(2304) <= not b or a;
    layer2_outputs(2305) <= '0';
    layer2_outputs(2306) <= a;
    layer2_outputs(2307) <= a and b;
    layer2_outputs(2308) <= a or b;
    layer2_outputs(2309) <= not (a or b);
    layer2_outputs(2310) <= not a or b;
    layer2_outputs(2311) <= a and not b;
    layer2_outputs(2312) <= a;
    layer2_outputs(2313) <= a and b;
    layer2_outputs(2314) <= not a;
    layer2_outputs(2315) <= a or b;
    layer2_outputs(2316) <= a;
    layer2_outputs(2317) <= b;
    layer2_outputs(2318) <= '0';
    layer2_outputs(2319) <= not (a or b);
    layer2_outputs(2320) <= not (a or b);
    layer2_outputs(2321) <= not (a or b);
    layer2_outputs(2322) <= a;
    layer2_outputs(2323) <= b;
    layer2_outputs(2324) <= b;
    layer2_outputs(2325) <= not a or b;
    layer2_outputs(2326) <= '1';
    layer2_outputs(2327) <= not b;
    layer2_outputs(2328) <= not (a xor b);
    layer2_outputs(2329) <= a or b;
    layer2_outputs(2330) <= not (a and b);
    layer2_outputs(2331) <= '1';
    layer2_outputs(2332) <= '0';
    layer2_outputs(2333) <= not b;
    layer2_outputs(2334) <= a and b;
    layer2_outputs(2335) <= b;
    layer2_outputs(2336) <= not b;
    layer2_outputs(2337) <= a and not b;
    layer2_outputs(2338) <= a and not b;
    layer2_outputs(2339) <= '0';
    layer2_outputs(2340) <= a or b;
    layer2_outputs(2341) <= not (a or b);
    layer2_outputs(2342) <= not b or a;
    layer2_outputs(2343) <= b and not a;
    layer2_outputs(2344) <= not (a or b);
    layer2_outputs(2345) <= a and b;
    layer2_outputs(2346) <= b;
    layer2_outputs(2347) <= a;
    layer2_outputs(2348) <= not (a or b);
    layer2_outputs(2349) <= not (a or b);
    layer2_outputs(2350) <= not (a xor b);
    layer2_outputs(2351) <= b and not a;
    layer2_outputs(2352) <= b and not a;
    layer2_outputs(2353) <= '1';
    layer2_outputs(2354) <= b;
    layer2_outputs(2355) <= not (a or b);
    layer2_outputs(2356) <= b;
    layer2_outputs(2357) <= not a;
    layer2_outputs(2358) <= not a or b;
    layer2_outputs(2359) <= not b or a;
    layer2_outputs(2360) <= b;
    layer2_outputs(2361) <= not b or a;
    layer2_outputs(2362) <= a and not b;
    layer2_outputs(2363) <= not b;
    layer2_outputs(2364) <= a or b;
    layer2_outputs(2365) <= not b or a;
    layer2_outputs(2366) <= '1';
    layer2_outputs(2367) <= a or b;
    layer2_outputs(2368) <= not (a or b);
    layer2_outputs(2369) <= not (a xor b);
    layer2_outputs(2370) <= '0';
    layer2_outputs(2371) <= a or b;
    layer2_outputs(2372) <= not b;
    layer2_outputs(2373) <= not a;
    layer2_outputs(2374) <= a and not b;
    layer2_outputs(2375) <= b;
    layer2_outputs(2376) <= not (a xor b);
    layer2_outputs(2377) <= '0';
    layer2_outputs(2378) <= a and not b;
    layer2_outputs(2379) <= a and b;
    layer2_outputs(2380) <= not (a xor b);
    layer2_outputs(2381) <= a or b;
    layer2_outputs(2382) <= not b or a;
    layer2_outputs(2383) <= not (a and b);
    layer2_outputs(2384) <= not (a or b);
    layer2_outputs(2385) <= not (a or b);
    layer2_outputs(2386) <= a;
    layer2_outputs(2387) <= not b or a;
    layer2_outputs(2388) <= not (a and b);
    layer2_outputs(2389) <= not b or a;
    layer2_outputs(2390) <= '0';
    layer2_outputs(2391) <= '0';
    layer2_outputs(2392) <= a and not b;
    layer2_outputs(2393) <= '0';
    layer2_outputs(2394) <= not (a and b);
    layer2_outputs(2395) <= '1';
    layer2_outputs(2396) <= a and not b;
    layer2_outputs(2397) <= not (a and b);
    layer2_outputs(2398) <= '1';
    layer2_outputs(2399) <= not a or b;
    layer2_outputs(2400) <= '1';
    layer2_outputs(2401) <= not (a xor b);
    layer2_outputs(2402) <= '0';
    layer2_outputs(2403) <= not b or a;
    layer2_outputs(2404) <= not a;
    layer2_outputs(2405) <= a and b;
    layer2_outputs(2406) <= not b or a;
    layer2_outputs(2407) <= a or b;
    layer2_outputs(2408) <= not (a and b);
    layer2_outputs(2409) <= not a or b;
    layer2_outputs(2410) <= not a;
    layer2_outputs(2411) <= b;
    layer2_outputs(2412) <= '0';
    layer2_outputs(2413) <= '1';
    layer2_outputs(2414) <= a or b;
    layer2_outputs(2415) <= a or b;
    layer2_outputs(2416) <= '0';
    layer2_outputs(2417) <= a or b;
    layer2_outputs(2418) <= not a;
    layer2_outputs(2419) <= not b;
    layer2_outputs(2420) <= '1';
    layer2_outputs(2421) <= not (a xor b);
    layer2_outputs(2422) <= b;
    layer2_outputs(2423) <= not b;
    layer2_outputs(2424) <= not (a or b);
    layer2_outputs(2425) <= a or b;
    layer2_outputs(2426) <= a;
    layer2_outputs(2427) <= '0';
    layer2_outputs(2428) <= not (a and b);
    layer2_outputs(2429) <= not (a and b);
    layer2_outputs(2430) <= '1';
    layer2_outputs(2431) <= '1';
    layer2_outputs(2432) <= a and not b;
    layer2_outputs(2433) <= '0';
    layer2_outputs(2434) <= not b or a;
    layer2_outputs(2435) <= not (a and b);
    layer2_outputs(2436) <= a or b;
    layer2_outputs(2437) <= a and not b;
    layer2_outputs(2438) <= not a;
    layer2_outputs(2439) <= not b or a;
    layer2_outputs(2440) <= not a or b;
    layer2_outputs(2441) <= not (a and b);
    layer2_outputs(2442) <= a and b;
    layer2_outputs(2443) <= '1';
    layer2_outputs(2444) <= not b;
    layer2_outputs(2445) <= not b or a;
    layer2_outputs(2446) <= a and b;
    layer2_outputs(2447) <= a and not b;
    layer2_outputs(2448) <= b and not a;
    layer2_outputs(2449) <= b and not a;
    layer2_outputs(2450) <= not b;
    layer2_outputs(2451) <= a and b;
    layer2_outputs(2452) <= '0';
    layer2_outputs(2453) <= not b or a;
    layer2_outputs(2454) <= b and not a;
    layer2_outputs(2455) <= b and not a;
    layer2_outputs(2456) <= a and not b;
    layer2_outputs(2457) <= b;
    layer2_outputs(2458) <= a and b;
    layer2_outputs(2459) <= '0';
    layer2_outputs(2460) <= not (a and b);
    layer2_outputs(2461) <= a and b;
    layer2_outputs(2462) <= not (a or b);
    layer2_outputs(2463) <= not a or b;
    layer2_outputs(2464) <= not (a and b);
    layer2_outputs(2465) <= a or b;
    layer2_outputs(2466) <= not a or b;
    layer2_outputs(2467) <= b and not a;
    layer2_outputs(2468) <= a and not b;
    layer2_outputs(2469) <= not b;
    layer2_outputs(2470) <= not a or b;
    layer2_outputs(2471) <= not (a or b);
    layer2_outputs(2472) <= a;
    layer2_outputs(2473) <= not (a or b);
    layer2_outputs(2474) <= b;
    layer2_outputs(2475) <= not b;
    layer2_outputs(2476) <= '1';
    layer2_outputs(2477) <= a and not b;
    layer2_outputs(2478) <= '1';
    layer2_outputs(2479) <= a and b;
    layer2_outputs(2480) <= b;
    layer2_outputs(2481) <= '0';
    layer2_outputs(2482) <= '0';
    layer2_outputs(2483) <= a and b;
    layer2_outputs(2484) <= '1';
    layer2_outputs(2485) <= a or b;
    layer2_outputs(2486) <= a or b;
    layer2_outputs(2487) <= not a;
    layer2_outputs(2488) <= not (a and b);
    layer2_outputs(2489) <= '0';
    layer2_outputs(2490) <= not a or b;
    layer2_outputs(2491) <= not b;
    layer2_outputs(2492) <= a and b;
    layer2_outputs(2493) <= a and not b;
    layer2_outputs(2494) <= '0';
    layer2_outputs(2495) <= a or b;
    layer2_outputs(2496) <= '1';
    layer2_outputs(2497) <= '1';
    layer2_outputs(2498) <= '0';
    layer2_outputs(2499) <= not (a and b);
    layer2_outputs(2500) <= not a;
    layer2_outputs(2501) <= '0';
    layer2_outputs(2502) <= a or b;
    layer2_outputs(2503) <= not a or b;
    layer2_outputs(2504) <= a xor b;
    layer2_outputs(2505) <= not b or a;
    layer2_outputs(2506) <= b;
    layer2_outputs(2507) <= not b or a;
    layer2_outputs(2508) <= a;
    layer2_outputs(2509) <= a and b;
    layer2_outputs(2510) <= not a or b;
    layer2_outputs(2511) <= not (a and b);
    layer2_outputs(2512) <= '0';
    layer2_outputs(2513) <= not a or b;
    layer2_outputs(2514) <= not a;
    layer2_outputs(2515) <= not b;
    layer2_outputs(2516) <= not a or b;
    layer2_outputs(2517) <= not a or b;
    layer2_outputs(2518) <= b;
    layer2_outputs(2519) <= b;
    layer2_outputs(2520) <= not b or a;
    layer2_outputs(2521) <= b;
    layer2_outputs(2522) <= a;
    layer2_outputs(2523) <= '0';
    layer2_outputs(2524) <= not (a or b);
    layer2_outputs(2525) <= a and not b;
    layer2_outputs(2526) <= b and not a;
    layer2_outputs(2527) <= not b;
    layer2_outputs(2528) <= not a or b;
    layer2_outputs(2529) <= b;
    layer2_outputs(2530) <= '0';
    layer2_outputs(2531) <= '0';
    layer2_outputs(2532) <= not (a xor b);
    layer2_outputs(2533) <= not b or a;
    layer2_outputs(2534) <= not (a or b);
    layer2_outputs(2535) <= not b;
    layer2_outputs(2536) <= not (a or b);
    layer2_outputs(2537) <= b and not a;
    layer2_outputs(2538) <= a and b;
    layer2_outputs(2539) <= a or b;
    layer2_outputs(2540) <= not (a and b);
    layer2_outputs(2541) <= a and not b;
    layer2_outputs(2542) <= not b or a;
    layer2_outputs(2543) <= not b or a;
    layer2_outputs(2544) <= a and b;
    layer2_outputs(2545) <= b and not a;
    layer2_outputs(2546) <= a and not b;
    layer2_outputs(2547) <= '1';
    layer2_outputs(2548) <= not a;
    layer2_outputs(2549) <= not a;
    layer2_outputs(2550) <= '1';
    layer2_outputs(2551) <= not (a and b);
    layer2_outputs(2552) <= not b;
    layer2_outputs(2553) <= not (a or b);
    layer2_outputs(2554) <= a and b;
    layer2_outputs(2555) <= not (a and b);
    layer2_outputs(2556) <= '1';
    layer2_outputs(2557) <= not (a and b);
    layer2_outputs(2558) <= a and b;
    layer2_outputs(2559) <= '1';
    layer2_outputs(2560) <= a xor b;
    layer2_outputs(2561) <= not b or a;
    layer2_outputs(2562) <= b;
    layer2_outputs(2563) <= '1';
    layer2_outputs(2564) <= b and not a;
    layer2_outputs(2565) <= a and b;
    layer2_outputs(2566) <= not b;
    layer2_outputs(2567) <= '1';
    layer2_outputs(2568) <= not (a or b);
    layer2_outputs(2569) <= not b;
    layer2_outputs(2570) <= not b or a;
    layer2_outputs(2571) <= a and b;
    layer2_outputs(2572) <= '0';
    layer2_outputs(2573) <= not a;
    layer2_outputs(2574) <= a;
    layer2_outputs(2575) <= not a;
    layer2_outputs(2576) <= not a;
    layer2_outputs(2577) <= b;
    layer2_outputs(2578) <= '0';
    layer2_outputs(2579) <= a and b;
    layer2_outputs(2580) <= b and not a;
    layer2_outputs(2581) <= a or b;
    layer2_outputs(2582) <= not b or a;
    layer2_outputs(2583) <= a and not b;
    layer2_outputs(2584) <= not b;
    layer2_outputs(2585) <= not (a xor b);
    layer2_outputs(2586) <= b;
    layer2_outputs(2587) <= not b or a;
    layer2_outputs(2588) <= not (a and b);
    layer2_outputs(2589) <= a xor b;
    layer2_outputs(2590) <= '0';
    layer2_outputs(2591) <= not (a xor b);
    layer2_outputs(2592) <= a and not b;
    layer2_outputs(2593) <= not (a xor b);
    layer2_outputs(2594) <= '1';
    layer2_outputs(2595) <= not b or a;
    layer2_outputs(2596) <= a and b;
    layer2_outputs(2597) <= not (a or b);
    layer2_outputs(2598) <= b and not a;
    layer2_outputs(2599) <= not (a or b);
    layer2_outputs(2600) <= '0';
    layer2_outputs(2601) <= a or b;
    layer2_outputs(2602) <= a or b;
    layer2_outputs(2603) <= not (a xor b);
    layer2_outputs(2604) <= not a or b;
    layer2_outputs(2605) <= '1';
    layer2_outputs(2606) <= not (a and b);
    layer2_outputs(2607) <= not (a and b);
    layer2_outputs(2608) <= a and not b;
    layer2_outputs(2609) <= a;
    layer2_outputs(2610) <= a;
    layer2_outputs(2611) <= b;
    layer2_outputs(2612) <= not b or a;
    layer2_outputs(2613) <= '1';
    layer2_outputs(2614) <= a;
    layer2_outputs(2615) <= a and b;
    layer2_outputs(2616) <= not b;
    layer2_outputs(2617) <= a or b;
    layer2_outputs(2618) <= not (a and b);
    layer2_outputs(2619) <= not b or a;
    layer2_outputs(2620) <= not (a or b);
    layer2_outputs(2621) <= '0';
    layer2_outputs(2622) <= not a or b;
    layer2_outputs(2623) <= b;
    layer2_outputs(2624) <= '0';
    layer2_outputs(2625) <= not a;
    layer2_outputs(2626) <= not b;
    layer2_outputs(2627) <= '1';
    layer2_outputs(2628) <= not a or b;
    layer2_outputs(2629) <= not b or a;
    layer2_outputs(2630) <= not (a or b);
    layer2_outputs(2631) <= not b or a;
    layer2_outputs(2632) <= not b;
    layer2_outputs(2633) <= '1';
    layer2_outputs(2634) <= not a;
    layer2_outputs(2635) <= not a or b;
    layer2_outputs(2636) <= not a;
    layer2_outputs(2637) <= not b;
    layer2_outputs(2638) <= a;
    layer2_outputs(2639) <= not a;
    layer2_outputs(2640) <= a or b;
    layer2_outputs(2641) <= a;
    layer2_outputs(2642) <= not (a and b);
    layer2_outputs(2643) <= '1';
    layer2_outputs(2644) <= not b;
    layer2_outputs(2645) <= a;
    layer2_outputs(2646) <= '1';
    layer2_outputs(2647) <= not (a or b);
    layer2_outputs(2648) <= a;
    layer2_outputs(2649) <= not (a or b);
    layer2_outputs(2650) <= '0';
    layer2_outputs(2651) <= b;
    layer2_outputs(2652) <= a;
    layer2_outputs(2653) <= not a;
    layer2_outputs(2654) <= a and b;
    layer2_outputs(2655) <= b;
    layer2_outputs(2656) <= not b or a;
    layer2_outputs(2657) <= not b;
    layer2_outputs(2658) <= not (a xor b);
    layer2_outputs(2659) <= '1';
    layer2_outputs(2660) <= '0';
    layer2_outputs(2661) <= not a;
    layer2_outputs(2662) <= not (a or b);
    layer2_outputs(2663) <= not a or b;
    layer2_outputs(2664) <= '1';
    layer2_outputs(2665) <= a xor b;
    layer2_outputs(2666) <= not (a and b);
    layer2_outputs(2667) <= not b or a;
    layer2_outputs(2668) <= '1';
    layer2_outputs(2669) <= not (a or b);
    layer2_outputs(2670) <= not a or b;
    layer2_outputs(2671) <= b;
    layer2_outputs(2672) <= not a;
    layer2_outputs(2673) <= a;
    layer2_outputs(2674) <= not b or a;
    layer2_outputs(2675) <= not a;
    layer2_outputs(2676) <= a;
    layer2_outputs(2677) <= a;
    layer2_outputs(2678) <= a;
    layer2_outputs(2679) <= not (a or b);
    layer2_outputs(2680) <= a;
    layer2_outputs(2681) <= b and not a;
    layer2_outputs(2682) <= b;
    layer2_outputs(2683) <= not a;
    layer2_outputs(2684) <= a or b;
    layer2_outputs(2685) <= not b or a;
    layer2_outputs(2686) <= a;
    layer2_outputs(2687) <= '1';
    layer2_outputs(2688) <= not a;
    layer2_outputs(2689) <= not b;
    layer2_outputs(2690) <= a and not b;
    layer2_outputs(2691) <= a and b;
    layer2_outputs(2692) <= a xor b;
    layer2_outputs(2693) <= not a;
    layer2_outputs(2694) <= a or b;
    layer2_outputs(2695) <= not a;
    layer2_outputs(2696) <= a;
    layer2_outputs(2697) <= a or b;
    layer2_outputs(2698) <= not b or a;
    layer2_outputs(2699) <= not (a and b);
    layer2_outputs(2700) <= not (a xor b);
    layer2_outputs(2701) <= '0';
    layer2_outputs(2702) <= b and not a;
    layer2_outputs(2703) <= a and b;
    layer2_outputs(2704) <= not a;
    layer2_outputs(2705) <= b and not a;
    layer2_outputs(2706) <= a or b;
    layer2_outputs(2707) <= not b or a;
    layer2_outputs(2708) <= b and not a;
    layer2_outputs(2709) <= a and not b;
    layer2_outputs(2710) <= '0';
    layer2_outputs(2711) <= a and b;
    layer2_outputs(2712) <= not (a and b);
    layer2_outputs(2713) <= b and not a;
    layer2_outputs(2714) <= not (a or b);
    layer2_outputs(2715) <= not b;
    layer2_outputs(2716) <= not b;
    layer2_outputs(2717) <= not (a and b);
    layer2_outputs(2718) <= not b or a;
    layer2_outputs(2719) <= not (a or b);
    layer2_outputs(2720) <= '1';
    layer2_outputs(2721) <= a;
    layer2_outputs(2722) <= not a;
    layer2_outputs(2723) <= not a;
    layer2_outputs(2724) <= a or b;
    layer2_outputs(2725) <= a and not b;
    layer2_outputs(2726) <= a or b;
    layer2_outputs(2727) <= '0';
    layer2_outputs(2728) <= a;
    layer2_outputs(2729) <= a and not b;
    layer2_outputs(2730) <= b;
    layer2_outputs(2731) <= a or b;
    layer2_outputs(2732) <= a or b;
    layer2_outputs(2733) <= '0';
    layer2_outputs(2734) <= a or b;
    layer2_outputs(2735) <= '1';
    layer2_outputs(2736) <= not b or a;
    layer2_outputs(2737) <= a;
    layer2_outputs(2738) <= '1';
    layer2_outputs(2739) <= not a or b;
    layer2_outputs(2740) <= a;
    layer2_outputs(2741) <= not a;
    layer2_outputs(2742) <= '1';
    layer2_outputs(2743) <= a;
    layer2_outputs(2744) <= b and not a;
    layer2_outputs(2745) <= a and not b;
    layer2_outputs(2746) <= not a;
    layer2_outputs(2747) <= a and not b;
    layer2_outputs(2748) <= not (a and b);
    layer2_outputs(2749) <= not b;
    layer2_outputs(2750) <= not a;
    layer2_outputs(2751) <= a or b;
    layer2_outputs(2752) <= not (a or b);
    layer2_outputs(2753) <= a and b;
    layer2_outputs(2754) <= '1';
    layer2_outputs(2755) <= '1';
    layer2_outputs(2756) <= not (a xor b);
    layer2_outputs(2757) <= not (a and b);
    layer2_outputs(2758) <= a or b;
    layer2_outputs(2759) <= a;
    layer2_outputs(2760) <= a and not b;
    layer2_outputs(2761) <= not (a or b);
    layer2_outputs(2762) <= not b or a;
    layer2_outputs(2763) <= a and not b;
    layer2_outputs(2764) <= a;
    layer2_outputs(2765) <= not (a and b);
    layer2_outputs(2766) <= a and not b;
    layer2_outputs(2767) <= '1';
    layer2_outputs(2768) <= a and not b;
    layer2_outputs(2769) <= a and b;
    layer2_outputs(2770) <= b and not a;
    layer2_outputs(2771) <= a or b;
    layer2_outputs(2772) <= '0';
    layer2_outputs(2773) <= not a or b;
    layer2_outputs(2774) <= not (a or b);
    layer2_outputs(2775) <= a and not b;
    layer2_outputs(2776) <= not (a xor b);
    layer2_outputs(2777) <= a and not b;
    layer2_outputs(2778) <= a;
    layer2_outputs(2779) <= not a or b;
    layer2_outputs(2780) <= '0';
    layer2_outputs(2781) <= not (a xor b);
    layer2_outputs(2782) <= '1';
    layer2_outputs(2783) <= '1';
    layer2_outputs(2784) <= not a or b;
    layer2_outputs(2785) <= b and not a;
    layer2_outputs(2786) <= not (a or b);
    layer2_outputs(2787) <= a and b;
    layer2_outputs(2788) <= not b;
    layer2_outputs(2789) <= not b or a;
    layer2_outputs(2790) <= b and not a;
    layer2_outputs(2791) <= not (a or b);
    layer2_outputs(2792) <= not a;
    layer2_outputs(2793) <= a;
    layer2_outputs(2794) <= not b or a;
    layer2_outputs(2795) <= not a;
    layer2_outputs(2796) <= not b;
    layer2_outputs(2797) <= '0';
    layer2_outputs(2798) <= b and not a;
    layer2_outputs(2799) <= a and not b;
    layer2_outputs(2800) <= not b or a;
    layer2_outputs(2801) <= a;
    layer2_outputs(2802) <= not b or a;
    layer2_outputs(2803) <= b;
    layer2_outputs(2804) <= a and b;
    layer2_outputs(2805) <= '0';
    layer2_outputs(2806) <= b and not a;
    layer2_outputs(2807) <= '0';
    layer2_outputs(2808) <= not (a xor b);
    layer2_outputs(2809) <= not b;
    layer2_outputs(2810) <= not a;
    layer2_outputs(2811) <= not a;
    layer2_outputs(2812) <= a and not b;
    layer2_outputs(2813) <= not b or a;
    layer2_outputs(2814) <= not b;
    layer2_outputs(2815) <= a xor b;
    layer2_outputs(2816) <= '1';
    layer2_outputs(2817) <= a and not b;
    layer2_outputs(2818) <= a and b;
    layer2_outputs(2819) <= not (a or b);
    layer2_outputs(2820) <= not a;
    layer2_outputs(2821) <= '0';
    layer2_outputs(2822) <= a;
    layer2_outputs(2823) <= '0';
    layer2_outputs(2824) <= '0';
    layer2_outputs(2825) <= '1';
    layer2_outputs(2826) <= not (a and b);
    layer2_outputs(2827) <= not b;
    layer2_outputs(2828) <= '0';
    layer2_outputs(2829) <= a or b;
    layer2_outputs(2830) <= a or b;
    layer2_outputs(2831) <= '0';
    layer2_outputs(2832) <= not a or b;
    layer2_outputs(2833) <= '0';
    layer2_outputs(2834) <= a or b;
    layer2_outputs(2835) <= b;
    layer2_outputs(2836) <= not a;
    layer2_outputs(2837) <= '1';
    layer2_outputs(2838) <= not b;
    layer2_outputs(2839) <= not (a or b);
    layer2_outputs(2840) <= b;
    layer2_outputs(2841) <= b;
    layer2_outputs(2842) <= '0';
    layer2_outputs(2843) <= a and b;
    layer2_outputs(2844) <= not b or a;
    layer2_outputs(2845) <= a;
    layer2_outputs(2846) <= '1';
    layer2_outputs(2847) <= b and not a;
    layer2_outputs(2848) <= not (a or b);
    layer2_outputs(2849) <= not (a and b);
    layer2_outputs(2850) <= not a or b;
    layer2_outputs(2851) <= not a;
    layer2_outputs(2852) <= '1';
    layer2_outputs(2853) <= a;
    layer2_outputs(2854) <= not a or b;
    layer2_outputs(2855) <= b and not a;
    layer2_outputs(2856) <= a or b;
    layer2_outputs(2857) <= '0';
    layer2_outputs(2858) <= a and not b;
    layer2_outputs(2859) <= not b or a;
    layer2_outputs(2860) <= b;
    layer2_outputs(2861) <= a;
    layer2_outputs(2862) <= '1';
    layer2_outputs(2863) <= '0';
    layer2_outputs(2864) <= '0';
    layer2_outputs(2865) <= b and not a;
    layer2_outputs(2866) <= a and b;
    layer2_outputs(2867) <= b;
    layer2_outputs(2868) <= a and b;
    layer2_outputs(2869) <= not (a xor b);
    layer2_outputs(2870) <= a;
    layer2_outputs(2871) <= a;
    layer2_outputs(2872) <= not b;
    layer2_outputs(2873) <= not a;
    layer2_outputs(2874) <= not a or b;
    layer2_outputs(2875) <= b;
    layer2_outputs(2876) <= not b;
    layer2_outputs(2877) <= '1';
    layer2_outputs(2878) <= not a;
    layer2_outputs(2879) <= not (a or b);
    layer2_outputs(2880) <= '0';
    layer2_outputs(2881) <= a and not b;
    layer2_outputs(2882) <= a and not b;
    layer2_outputs(2883) <= a and not b;
    layer2_outputs(2884) <= not a or b;
    layer2_outputs(2885) <= a or b;
    layer2_outputs(2886) <= not a or b;
    layer2_outputs(2887) <= '0';
    layer2_outputs(2888) <= not (a or b);
    layer2_outputs(2889) <= a or b;
    layer2_outputs(2890) <= not a;
    layer2_outputs(2891) <= not b;
    layer2_outputs(2892) <= not (a xor b);
    layer2_outputs(2893) <= not (a or b);
    layer2_outputs(2894) <= a and not b;
    layer2_outputs(2895) <= not a;
    layer2_outputs(2896) <= b and not a;
    layer2_outputs(2897) <= not a;
    layer2_outputs(2898) <= not a or b;
    layer2_outputs(2899) <= b;
    layer2_outputs(2900) <= '1';
    layer2_outputs(2901) <= not b;
    layer2_outputs(2902) <= a and not b;
    layer2_outputs(2903) <= a and b;
    layer2_outputs(2904) <= not b;
    layer2_outputs(2905) <= not a;
    layer2_outputs(2906) <= not (a and b);
    layer2_outputs(2907) <= '1';
    layer2_outputs(2908) <= not a;
    layer2_outputs(2909) <= b and not a;
    layer2_outputs(2910) <= not b or a;
    layer2_outputs(2911) <= a or b;
    layer2_outputs(2912) <= '1';
    layer2_outputs(2913) <= '1';
    layer2_outputs(2914) <= b;
    layer2_outputs(2915) <= b;
    layer2_outputs(2916) <= not (a or b);
    layer2_outputs(2917) <= a;
    layer2_outputs(2918) <= not b;
    layer2_outputs(2919) <= a xor b;
    layer2_outputs(2920) <= a;
    layer2_outputs(2921) <= not b;
    layer2_outputs(2922) <= not (a or b);
    layer2_outputs(2923) <= not (a or b);
    layer2_outputs(2924) <= '0';
    layer2_outputs(2925) <= a and not b;
    layer2_outputs(2926) <= not a or b;
    layer2_outputs(2927) <= a or b;
    layer2_outputs(2928) <= '0';
    layer2_outputs(2929) <= not a;
    layer2_outputs(2930) <= b;
    layer2_outputs(2931) <= '1';
    layer2_outputs(2932) <= not (a and b);
    layer2_outputs(2933) <= a and b;
    layer2_outputs(2934) <= a or b;
    layer2_outputs(2935) <= not b;
    layer2_outputs(2936) <= '1';
    layer2_outputs(2937) <= not (a or b);
    layer2_outputs(2938) <= a xor b;
    layer2_outputs(2939) <= not (a or b);
    layer2_outputs(2940) <= '0';
    layer2_outputs(2941) <= not a or b;
    layer2_outputs(2942) <= a or b;
    layer2_outputs(2943) <= a or b;
    layer2_outputs(2944) <= a and not b;
    layer2_outputs(2945) <= '0';
    layer2_outputs(2946) <= not (a or b);
    layer2_outputs(2947) <= not a;
    layer2_outputs(2948) <= a;
    layer2_outputs(2949) <= a;
    layer2_outputs(2950) <= a and not b;
    layer2_outputs(2951) <= a or b;
    layer2_outputs(2952) <= not (a and b);
    layer2_outputs(2953) <= not a or b;
    layer2_outputs(2954) <= not b or a;
    layer2_outputs(2955) <= b;
    layer2_outputs(2956) <= '1';
    layer2_outputs(2957) <= not (a and b);
    layer2_outputs(2958) <= not (a or b);
    layer2_outputs(2959) <= b and not a;
    layer2_outputs(2960) <= a or b;
    layer2_outputs(2961) <= '1';
    layer2_outputs(2962) <= not b;
    layer2_outputs(2963) <= b and not a;
    layer2_outputs(2964) <= not b or a;
    layer2_outputs(2965) <= '0';
    layer2_outputs(2966) <= a and not b;
    layer2_outputs(2967) <= not a or b;
    layer2_outputs(2968) <= a and not b;
    layer2_outputs(2969) <= not a or b;
    layer2_outputs(2970) <= '0';
    layer2_outputs(2971) <= not b or a;
    layer2_outputs(2972) <= b;
    layer2_outputs(2973) <= '0';
    layer2_outputs(2974) <= not a or b;
    layer2_outputs(2975) <= '0';
    layer2_outputs(2976) <= a;
    layer2_outputs(2977) <= a or b;
    layer2_outputs(2978) <= b and not a;
    layer2_outputs(2979) <= not (a or b);
    layer2_outputs(2980) <= a;
    layer2_outputs(2981) <= a or b;
    layer2_outputs(2982) <= not b;
    layer2_outputs(2983) <= '0';
    layer2_outputs(2984) <= not a or b;
    layer2_outputs(2985) <= not b or a;
    layer2_outputs(2986) <= a and not b;
    layer2_outputs(2987) <= b;
    layer2_outputs(2988) <= a or b;
    layer2_outputs(2989) <= b;
    layer2_outputs(2990) <= b and not a;
    layer2_outputs(2991) <= '0';
    layer2_outputs(2992) <= '1';
    layer2_outputs(2993) <= a xor b;
    layer2_outputs(2994) <= '0';
    layer2_outputs(2995) <= '0';
    layer2_outputs(2996) <= '1';
    layer2_outputs(2997) <= not a or b;
    layer2_outputs(2998) <= b and not a;
    layer2_outputs(2999) <= not (a and b);
    layer2_outputs(3000) <= not b;
    layer2_outputs(3001) <= '1';
    layer2_outputs(3002) <= not (a xor b);
    layer2_outputs(3003) <= '1';
    layer2_outputs(3004) <= not a or b;
    layer2_outputs(3005) <= not b;
    layer2_outputs(3006) <= '1';
    layer2_outputs(3007) <= '0';
    layer2_outputs(3008) <= a;
    layer2_outputs(3009) <= a;
    layer2_outputs(3010) <= not (a and b);
    layer2_outputs(3011) <= a xor b;
    layer2_outputs(3012) <= b and not a;
    layer2_outputs(3013) <= not b;
    layer2_outputs(3014) <= not b or a;
    layer2_outputs(3015) <= '0';
    layer2_outputs(3016) <= a or b;
    layer2_outputs(3017) <= b;
    layer2_outputs(3018) <= not (a and b);
    layer2_outputs(3019) <= not b;
    layer2_outputs(3020) <= '0';
    layer2_outputs(3021) <= '0';
    layer2_outputs(3022) <= '1';
    layer2_outputs(3023) <= a and not b;
    layer2_outputs(3024) <= not (a and b);
    layer2_outputs(3025) <= b;
    layer2_outputs(3026) <= a xor b;
    layer2_outputs(3027) <= not (a or b);
    layer2_outputs(3028) <= '1';
    layer2_outputs(3029) <= not a;
    layer2_outputs(3030) <= not (a and b);
    layer2_outputs(3031) <= not (a and b);
    layer2_outputs(3032) <= a or b;
    layer2_outputs(3033) <= a;
    layer2_outputs(3034) <= not (a and b);
    layer2_outputs(3035) <= '1';
    layer2_outputs(3036) <= not b;
    layer2_outputs(3037) <= not (a and b);
    layer2_outputs(3038) <= not (a and b);
    layer2_outputs(3039) <= a xor b;
    layer2_outputs(3040) <= not (a and b);
    layer2_outputs(3041) <= b;
    layer2_outputs(3042) <= not b;
    layer2_outputs(3043) <= not a;
    layer2_outputs(3044) <= not b;
    layer2_outputs(3045) <= not a;
    layer2_outputs(3046) <= not (a or b);
    layer2_outputs(3047) <= a or b;
    layer2_outputs(3048) <= not a or b;
    layer2_outputs(3049) <= not a or b;
    layer2_outputs(3050) <= '0';
    layer2_outputs(3051) <= not a;
    layer2_outputs(3052) <= b;
    layer2_outputs(3053) <= a and b;
    layer2_outputs(3054) <= a and b;
    layer2_outputs(3055) <= a and b;
    layer2_outputs(3056) <= not a or b;
    layer2_outputs(3057) <= not a or b;
    layer2_outputs(3058) <= not (a or b);
    layer2_outputs(3059) <= '1';
    layer2_outputs(3060) <= not b;
    layer2_outputs(3061) <= not (a and b);
    layer2_outputs(3062) <= not (a or b);
    layer2_outputs(3063) <= '0';
    layer2_outputs(3064) <= '0';
    layer2_outputs(3065) <= not a or b;
    layer2_outputs(3066) <= not (a and b);
    layer2_outputs(3067) <= a and b;
    layer2_outputs(3068) <= not b or a;
    layer2_outputs(3069) <= a and b;
    layer2_outputs(3070) <= b and not a;
    layer2_outputs(3071) <= '0';
    layer2_outputs(3072) <= a or b;
    layer2_outputs(3073) <= b and not a;
    layer2_outputs(3074) <= not (a or b);
    layer2_outputs(3075) <= b and not a;
    layer2_outputs(3076) <= b;
    layer2_outputs(3077) <= not b;
    layer2_outputs(3078) <= not b;
    layer2_outputs(3079) <= b and not a;
    layer2_outputs(3080) <= '1';
    layer2_outputs(3081) <= a or b;
    layer2_outputs(3082) <= not a;
    layer2_outputs(3083) <= b;
    layer2_outputs(3084) <= not b or a;
    layer2_outputs(3085) <= b;
    layer2_outputs(3086) <= not a;
    layer2_outputs(3087) <= b;
    layer2_outputs(3088) <= '1';
    layer2_outputs(3089) <= not b or a;
    layer2_outputs(3090) <= not b;
    layer2_outputs(3091) <= a and not b;
    layer2_outputs(3092) <= not b;
    layer2_outputs(3093) <= '0';
    layer2_outputs(3094) <= not a or b;
    layer2_outputs(3095) <= '0';
    layer2_outputs(3096) <= '0';
    layer2_outputs(3097) <= b;
    layer2_outputs(3098) <= not b or a;
    layer2_outputs(3099) <= b;
    layer2_outputs(3100) <= not a;
    layer2_outputs(3101) <= a and not b;
    layer2_outputs(3102) <= not b or a;
    layer2_outputs(3103) <= b;
    layer2_outputs(3104) <= '0';
    layer2_outputs(3105) <= not (a or b);
    layer2_outputs(3106) <= not (a xor b);
    layer2_outputs(3107) <= '1';
    layer2_outputs(3108) <= not a;
    layer2_outputs(3109) <= a;
    layer2_outputs(3110) <= not b;
    layer2_outputs(3111) <= b;
    layer2_outputs(3112) <= b;
    layer2_outputs(3113) <= a;
    layer2_outputs(3114) <= not b;
    layer2_outputs(3115) <= not a;
    layer2_outputs(3116) <= a and not b;
    layer2_outputs(3117) <= not (a and b);
    layer2_outputs(3118) <= not (a xor b);
    layer2_outputs(3119) <= not a or b;
    layer2_outputs(3120) <= a and not b;
    layer2_outputs(3121) <= not (a xor b);
    layer2_outputs(3122) <= '0';
    layer2_outputs(3123) <= not (a or b);
    layer2_outputs(3124) <= a and not b;
    layer2_outputs(3125) <= b and not a;
    layer2_outputs(3126) <= not (a or b);
    layer2_outputs(3127) <= a and not b;
    layer2_outputs(3128) <= not b or a;
    layer2_outputs(3129) <= a and b;
    layer2_outputs(3130) <= a or b;
    layer2_outputs(3131) <= a or b;
    layer2_outputs(3132) <= not a or b;
    layer2_outputs(3133) <= b;
    layer2_outputs(3134) <= a;
    layer2_outputs(3135) <= a or b;
    layer2_outputs(3136) <= not b or a;
    layer2_outputs(3137) <= not b;
    layer2_outputs(3138) <= b;
    layer2_outputs(3139) <= not (a and b);
    layer2_outputs(3140) <= '1';
    layer2_outputs(3141) <= '1';
    layer2_outputs(3142) <= b and not a;
    layer2_outputs(3143) <= a and b;
    layer2_outputs(3144) <= not (a and b);
    layer2_outputs(3145) <= b and not a;
    layer2_outputs(3146) <= '0';
    layer2_outputs(3147) <= '1';
    layer2_outputs(3148) <= not a or b;
    layer2_outputs(3149) <= not (a and b);
    layer2_outputs(3150) <= not (a and b);
    layer2_outputs(3151) <= a or b;
    layer2_outputs(3152) <= not a;
    layer2_outputs(3153) <= '1';
    layer2_outputs(3154) <= not b or a;
    layer2_outputs(3155) <= a or b;
    layer2_outputs(3156) <= not (a and b);
    layer2_outputs(3157) <= a;
    layer2_outputs(3158) <= not a;
    layer2_outputs(3159) <= not (a or b);
    layer2_outputs(3160) <= '1';
    layer2_outputs(3161) <= b;
    layer2_outputs(3162) <= not (a and b);
    layer2_outputs(3163) <= a;
    layer2_outputs(3164) <= a and b;
    layer2_outputs(3165) <= not a;
    layer2_outputs(3166) <= not b or a;
    layer2_outputs(3167) <= not a;
    layer2_outputs(3168) <= a or b;
    layer2_outputs(3169) <= '1';
    layer2_outputs(3170) <= b;
    layer2_outputs(3171) <= not b;
    layer2_outputs(3172) <= a and b;
    layer2_outputs(3173) <= not a;
    layer2_outputs(3174) <= not b or a;
    layer2_outputs(3175) <= a or b;
    layer2_outputs(3176) <= b;
    layer2_outputs(3177) <= a or b;
    layer2_outputs(3178) <= a or b;
    layer2_outputs(3179) <= not (a or b);
    layer2_outputs(3180) <= b and not a;
    layer2_outputs(3181) <= a xor b;
    layer2_outputs(3182) <= not (a or b);
    layer2_outputs(3183) <= a and not b;
    layer2_outputs(3184) <= '1';
    layer2_outputs(3185) <= a and not b;
    layer2_outputs(3186) <= not (a and b);
    layer2_outputs(3187) <= a or b;
    layer2_outputs(3188) <= not (a xor b);
    layer2_outputs(3189) <= not a or b;
    layer2_outputs(3190) <= '1';
    layer2_outputs(3191) <= a and not b;
    layer2_outputs(3192) <= '0';
    layer2_outputs(3193) <= b and not a;
    layer2_outputs(3194) <= not a;
    layer2_outputs(3195) <= '0';
    layer2_outputs(3196) <= not a;
    layer2_outputs(3197) <= not b;
    layer2_outputs(3198) <= a xor b;
    layer2_outputs(3199) <= b and not a;
    layer2_outputs(3200) <= '0';
    layer2_outputs(3201) <= not b or a;
    layer2_outputs(3202) <= a and b;
    layer2_outputs(3203) <= a and not b;
    layer2_outputs(3204) <= not (a and b);
    layer2_outputs(3205) <= a and b;
    layer2_outputs(3206) <= a;
    layer2_outputs(3207) <= b;
    layer2_outputs(3208) <= '1';
    layer2_outputs(3209) <= '0';
    layer2_outputs(3210) <= a xor b;
    layer2_outputs(3211) <= not (a and b);
    layer2_outputs(3212) <= not a or b;
    layer2_outputs(3213) <= not (a and b);
    layer2_outputs(3214) <= a or b;
    layer2_outputs(3215) <= a or b;
    layer2_outputs(3216) <= a xor b;
    layer2_outputs(3217) <= a and b;
    layer2_outputs(3218) <= not b;
    layer2_outputs(3219) <= not (a and b);
    layer2_outputs(3220) <= a and not b;
    layer2_outputs(3221) <= a or b;
    layer2_outputs(3222) <= a and b;
    layer2_outputs(3223) <= a;
    layer2_outputs(3224) <= a;
    layer2_outputs(3225) <= not (a or b);
    layer2_outputs(3226) <= a xor b;
    layer2_outputs(3227) <= not b;
    layer2_outputs(3228) <= a and b;
    layer2_outputs(3229) <= b;
    layer2_outputs(3230) <= '0';
    layer2_outputs(3231) <= b and not a;
    layer2_outputs(3232) <= a xor b;
    layer2_outputs(3233) <= b;
    layer2_outputs(3234) <= not a;
    layer2_outputs(3235) <= not (a and b);
    layer2_outputs(3236) <= a and b;
    layer2_outputs(3237) <= not (a and b);
    layer2_outputs(3238) <= not (a or b);
    layer2_outputs(3239) <= not a or b;
    layer2_outputs(3240) <= b and not a;
    layer2_outputs(3241) <= not a;
    layer2_outputs(3242) <= not a;
    layer2_outputs(3243) <= not b;
    layer2_outputs(3244) <= not b or a;
    layer2_outputs(3245) <= a;
    layer2_outputs(3246) <= '0';
    layer2_outputs(3247) <= a or b;
    layer2_outputs(3248) <= not b or a;
    layer2_outputs(3249) <= b and not a;
    layer2_outputs(3250) <= not b or a;
    layer2_outputs(3251) <= not b;
    layer2_outputs(3252) <= a;
    layer2_outputs(3253) <= a;
    layer2_outputs(3254) <= a xor b;
    layer2_outputs(3255) <= '1';
    layer2_outputs(3256) <= a xor b;
    layer2_outputs(3257) <= '0';
    layer2_outputs(3258) <= '1';
    layer2_outputs(3259) <= '0';
    layer2_outputs(3260) <= b;
    layer2_outputs(3261) <= '0';
    layer2_outputs(3262) <= '0';
    layer2_outputs(3263) <= not b or a;
    layer2_outputs(3264) <= not (a xor b);
    layer2_outputs(3265) <= a or b;
    layer2_outputs(3266) <= a;
    layer2_outputs(3267) <= '0';
    layer2_outputs(3268) <= '1';
    layer2_outputs(3269) <= '1';
    layer2_outputs(3270) <= a or b;
    layer2_outputs(3271) <= not a or b;
    layer2_outputs(3272) <= not a;
    layer2_outputs(3273) <= a and not b;
    layer2_outputs(3274) <= a and b;
    layer2_outputs(3275) <= a and not b;
    layer2_outputs(3276) <= not b or a;
    layer2_outputs(3277) <= a;
    layer2_outputs(3278) <= '1';
    layer2_outputs(3279) <= '0';
    layer2_outputs(3280) <= not (a or b);
    layer2_outputs(3281) <= a or b;
    layer2_outputs(3282) <= not a or b;
    layer2_outputs(3283) <= a xor b;
    layer2_outputs(3284) <= not (a and b);
    layer2_outputs(3285) <= a and b;
    layer2_outputs(3286) <= a or b;
    layer2_outputs(3287) <= '1';
    layer2_outputs(3288) <= not a or b;
    layer2_outputs(3289) <= not b or a;
    layer2_outputs(3290) <= not b or a;
    layer2_outputs(3291) <= b and not a;
    layer2_outputs(3292) <= not (a and b);
    layer2_outputs(3293) <= not (a or b);
    layer2_outputs(3294) <= a;
    layer2_outputs(3295) <= a and b;
    layer2_outputs(3296) <= a and not b;
    layer2_outputs(3297) <= a or b;
    layer2_outputs(3298) <= a and b;
    layer2_outputs(3299) <= not (a and b);
    layer2_outputs(3300) <= b;
    layer2_outputs(3301) <= b and not a;
    layer2_outputs(3302) <= a or b;
    layer2_outputs(3303) <= a or b;
    layer2_outputs(3304) <= not (a and b);
    layer2_outputs(3305) <= a and b;
    layer2_outputs(3306) <= a or b;
    layer2_outputs(3307) <= not a;
    layer2_outputs(3308) <= b and not a;
    layer2_outputs(3309) <= not a;
    layer2_outputs(3310) <= '0';
    layer2_outputs(3311) <= not b or a;
    layer2_outputs(3312) <= not a;
    layer2_outputs(3313) <= a;
    layer2_outputs(3314) <= a or b;
    layer2_outputs(3315) <= '0';
    layer2_outputs(3316) <= b and not a;
    layer2_outputs(3317) <= not a or b;
    layer2_outputs(3318) <= a xor b;
    layer2_outputs(3319) <= not (a or b);
    layer2_outputs(3320) <= not (a or b);
    layer2_outputs(3321) <= not b;
    layer2_outputs(3322) <= not a or b;
    layer2_outputs(3323) <= not a or b;
    layer2_outputs(3324) <= '1';
    layer2_outputs(3325) <= b;
    layer2_outputs(3326) <= not (a and b);
    layer2_outputs(3327) <= not (a or b);
    layer2_outputs(3328) <= a xor b;
    layer2_outputs(3329) <= b and not a;
    layer2_outputs(3330) <= a and not b;
    layer2_outputs(3331) <= a and not b;
    layer2_outputs(3332) <= not a;
    layer2_outputs(3333) <= not a or b;
    layer2_outputs(3334) <= not a or b;
    layer2_outputs(3335) <= not (a xor b);
    layer2_outputs(3336) <= b and not a;
    layer2_outputs(3337) <= a and not b;
    layer2_outputs(3338) <= '1';
    layer2_outputs(3339) <= '0';
    layer2_outputs(3340) <= not (a or b);
    layer2_outputs(3341) <= '0';
    layer2_outputs(3342) <= a or b;
    layer2_outputs(3343) <= not (a xor b);
    layer2_outputs(3344) <= '1';
    layer2_outputs(3345) <= not a or b;
    layer2_outputs(3346) <= not a or b;
    layer2_outputs(3347) <= a and not b;
    layer2_outputs(3348) <= b;
    layer2_outputs(3349) <= not b;
    layer2_outputs(3350) <= a xor b;
    layer2_outputs(3351) <= '1';
    layer2_outputs(3352) <= a and not b;
    layer2_outputs(3353) <= b and not a;
    layer2_outputs(3354) <= a or b;
    layer2_outputs(3355) <= a;
    layer2_outputs(3356) <= not b or a;
    layer2_outputs(3357) <= not b;
    layer2_outputs(3358) <= not a;
    layer2_outputs(3359) <= not b or a;
    layer2_outputs(3360) <= b and not a;
    layer2_outputs(3361) <= a and not b;
    layer2_outputs(3362) <= not (a or b);
    layer2_outputs(3363) <= a and b;
    layer2_outputs(3364) <= a;
    layer2_outputs(3365) <= a and not b;
    layer2_outputs(3366) <= a or b;
    layer2_outputs(3367) <= not a or b;
    layer2_outputs(3368) <= a;
    layer2_outputs(3369) <= not (a or b);
    layer2_outputs(3370) <= '0';
    layer2_outputs(3371) <= '1';
    layer2_outputs(3372) <= b;
    layer2_outputs(3373) <= '0';
    layer2_outputs(3374) <= not (a xor b);
    layer2_outputs(3375) <= b;
    layer2_outputs(3376) <= '0';
    layer2_outputs(3377) <= not a or b;
    layer2_outputs(3378) <= a and b;
    layer2_outputs(3379) <= a and not b;
    layer2_outputs(3380) <= not (a or b);
    layer2_outputs(3381) <= b;
    layer2_outputs(3382) <= not a or b;
    layer2_outputs(3383) <= '0';
    layer2_outputs(3384) <= a and not b;
    layer2_outputs(3385) <= a and b;
    layer2_outputs(3386) <= not (a or b);
    layer2_outputs(3387) <= '0';
    layer2_outputs(3388) <= not a or b;
    layer2_outputs(3389) <= '1';
    layer2_outputs(3390) <= not a or b;
    layer2_outputs(3391) <= a;
    layer2_outputs(3392) <= not b or a;
    layer2_outputs(3393) <= not (a or b);
    layer2_outputs(3394) <= not (a or b);
    layer2_outputs(3395) <= a and b;
    layer2_outputs(3396) <= not a or b;
    layer2_outputs(3397) <= not b or a;
    layer2_outputs(3398) <= a and not b;
    layer2_outputs(3399) <= b;
    layer2_outputs(3400) <= not a;
    layer2_outputs(3401) <= b and not a;
    layer2_outputs(3402) <= b;
    layer2_outputs(3403) <= not b or a;
    layer2_outputs(3404) <= not b;
    layer2_outputs(3405) <= b;
    layer2_outputs(3406) <= not (a or b);
    layer2_outputs(3407) <= '0';
    layer2_outputs(3408) <= a and b;
    layer2_outputs(3409) <= '1';
    layer2_outputs(3410) <= a and b;
    layer2_outputs(3411) <= not (a and b);
    layer2_outputs(3412) <= not (a xor b);
    layer2_outputs(3413) <= a and b;
    layer2_outputs(3414) <= '1';
    layer2_outputs(3415) <= not (a xor b);
    layer2_outputs(3416) <= a and not b;
    layer2_outputs(3417) <= '1';
    layer2_outputs(3418) <= a and not b;
    layer2_outputs(3419) <= '1';
    layer2_outputs(3420) <= not (a or b);
    layer2_outputs(3421) <= a and not b;
    layer2_outputs(3422) <= not b;
    layer2_outputs(3423) <= '0';
    layer2_outputs(3424) <= not a or b;
    layer2_outputs(3425) <= not b;
    layer2_outputs(3426) <= not a;
    layer2_outputs(3427) <= not (a or b);
    layer2_outputs(3428) <= b;
    layer2_outputs(3429) <= '1';
    layer2_outputs(3430) <= not (a or b);
    layer2_outputs(3431) <= not (a and b);
    layer2_outputs(3432) <= a or b;
    layer2_outputs(3433) <= not a or b;
    layer2_outputs(3434) <= not (a and b);
    layer2_outputs(3435) <= a xor b;
    layer2_outputs(3436) <= a;
    layer2_outputs(3437) <= '0';
    layer2_outputs(3438) <= b and not a;
    layer2_outputs(3439) <= not (a or b);
    layer2_outputs(3440) <= not b or a;
    layer2_outputs(3441) <= not (a and b);
    layer2_outputs(3442) <= not b;
    layer2_outputs(3443) <= b and not a;
    layer2_outputs(3444) <= a and b;
    layer2_outputs(3445) <= b and not a;
    layer2_outputs(3446) <= not (a and b);
    layer2_outputs(3447) <= not b;
    layer2_outputs(3448) <= b;
    layer2_outputs(3449) <= a;
    layer2_outputs(3450) <= a and b;
    layer2_outputs(3451) <= '1';
    layer2_outputs(3452) <= not b;
    layer2_outputs(3453) <= a and not b;
    layer2_outputs(3454) <= not b;
    layer2_outputs(3455) <= not (a or b);
    layer2_outputs(3456) <= b;
    layer2_outputs(3457) <= a or b;
    layer2_outputs(3458) <= b and not a;
    layer2_outputs(3459) <= a and b;
    layer2_outputs(3460) <= a;
    layer2_outputs(3461) <= a or b;
    layer2_outputs(3462) <= not (a or b);
    layer2_outputs(3463) <= a and b;
    layer2_outputs(3464) <= not (a and b);
    layer2_outputs(3465) <= a and b;
    layer2_outputs(3466) <= not (a xor b);
    layer2_outputs(3467) <= not (a and b);
    layer2_outputs(3468) <= a and b;
    layer2_outputs(3469) <= a and not b;
    layer2_outputs(3470) <= b;
    layer2_outputs(3471) <= b and not a;
    layer2_outputs(3472) <= b and not a;
    layer2_outputs(3473) <= a and b;
    layer2_outputs(3474) <= a or b;
    layer2_outputs(3475) <= a and b;
    layer2_outputs(3476) <= a or b;
    layer2_outputs(3477) <= not (a and b);
    layer2_outputs(3478) <= '1';
    layer2_outputs(3479) <= not (a and b);
    layer2_outputs(3480) <= b;
    layer2_outputs(3481) <= a and not b;
    layer2_outputs(3482) <= not b;
    layer2_outputs(3483) <= b and not a;
    layer2_outputs(3484) <= a or b;
    layer2_outputs(3485) <= a and not b;
    layer2_outputs(3486) <= a and not b;
    layer2_outputs(3487) <= not b;
    layer2_outputs(3488) <= not (a and b);
    layer2_outputs(3489) <= '0';
    layer2_outputs(3490) <= b and not a;
    layer2_outputs(3491) <= not a;
    layer2_outputs(3492) <= b and not a;
    layer2_outputs(3493) <= b;
    layer2_outputs(3494) <= '0';
    layer2_outputs(3495) <= not a;
    layer2_outputs(3496) <= not a or b;
    layer2_outputs(3497) <= not (a or b);
    layer2_outputs(3498) <= not (a or b);
    layer2_outputs(3499) <= not (a and b);
    layer2_outputs(3500) <= not a or b;
    layer2_outputs(3501) <= not (a or b);
    layer2_outputs(3502) <= not (a and b);
    layer2_outputs(3503) <= a;
    layer2_outputs(3504) <= a and b;
    layer2_outputs(3505) <= '0';
    layer2_outputs(3506) <= a;
    layer2_outputs(3507) <= b and not a;
    layer2_outputs(3508) <= a xor b;
    layer2_outputs(3509) <= b and not a;
    layer2_outputs(3510) <= '1';
    layer2_outputs(3511) <= '0';
    layer2_outputs(3512) <= '1';
    layer2_outputs(3513) <= not (a or b);
    layer2_outputs(3514) <= not (a xor b);
    layer2_outputs(3515) <= a and not b;
    layer2_outputs(3516) <= a and not b;
    layer2_outputs(3517) <= not (a and b);
    layer2_outputs(3518) <= not (a or b);
    layer2_outputs(3519) <= not (a xor b);
    layer2_outputs(3520) <= a and not b;
    layer2_outputs(3521) <= '0';
    layer2_outputs(3522) <= b and not a;
    layer2_outputs(3523) <= a;
    layer2_outputs(3524) <= a or b;
    layer2_outputs(3525) <= not a or b;
    layer2_outputs(3526) <= '1';
    layer2_outputs(3527) <= not (a and b);
    layer2_outputs(3528) <= a;
    layer2_outputs(3529) <= a or b;
    layer2_outputs(3530) <= not a or b;
    layer2_outputs(3531) <= not b or a;
    layer2_outputs(3532) <= a and not b;
    layer2_outputs(3533) <= '1';
    layer2_outputs(3534) <= a or b;
    layer2_outputs(3535) <= '0';
    layer2_outputs(3536) <= '1';
    layer2_outputs(3537) <= not b or a;
    layer2_outputs(3538) <= not b or a;
    layer2_outputs(3539) <= a and not b;
    layer2_outputs(3540) <= not (a or b);
    layer2_outputs(3541) <= a xor b;
    layer2_outputs(3542) <= '1';
    layer2_outputs(3543) <= not a or b;
    layer2_outputs(3544) <= '1';
    layer2_outputs(3545) <= not b;
    layer2_outputs(3546) <= not a;
    layer2_outputs(3547) <= b;
    layer2_outputs(3548) <= a and b;
    layer2_outputs(3549) <= not (a or b);
    layer2_outputs(3550) <= a and b;
    layer2_outputs(3551) <= not a;
    layer2_outputs(3552) <= a or b;
    layer2_outputs(3553) <= not b;
    layer2_outputs(3554) <= not b or a;
    layer2_outputs(3555) <= a and b;
    layer2_outputs(3556) <= '1';
    layer2_outputs(3557) <= not (a or b);
    layer2_outputs(3558) <= not a;
    layer2_outputs(3559) <= not a;
    layer2_outputs(3560) <= '0';
    layer2_outputs(3561) <= b and not a;
    layer2_outputs(3562) <= not a or b;
    layer2_outputs(3563) <= not (a or b);
    layer2_outputs(3564) <= a and not b;
    layer2_outputs(3565) <= '0';
    layer2_outputs(3566) <= a;
    layer2_outputs(3567) <= b;
    layer2_outputs(3568) <= a and not b;
    layer2_outputs(3569) <= not a;
    layer2_outputs(3570) <= not a or b;
    layer2_outputs(3571) <= '0';
    layer2_outputs(3572) <= not b or a;
    layer2_outputs(3573) <= b;
    layer2_outputs(3574) <= a or b;
    layer2_outputs(3575) <= '1';
    layer2_outputs(3576) <= a;
    layer2_outputs(3577) <= not b or a;
    layer2_outputs(3578) <= not (a or b);
    layer2_outputs(3579) <= '0';
    layer2_outputs(3580) <= '1';
    layer2_outputs(3581) <= not (a or b);
    layer2_outputs(3582) <= '1';
    layer2_outputs(3583) <= not b;
    layer2_outputs(3584) <= a and not b;
    layer2_outputs(3585) <= not (a or b);
    layer2_outputs(3586) <= a;
    layer2_outputs(3587) <= not b or a;
    layer2_outputs(3588) <= not a or b;
    layer2_outputs(3589) <= a;
    layer2_outputs(3590) <= '1';
    layer2_outputs(3591) <= not b or a;
    layer2_outputs(3592) <= a;
    layer2_outputs(3593) <= '0';
    layer2_outputs(3594) <= not (a or b);
    layer2_outputs(3595) <= a or b;
    layer2_outputs(3596) <= '1';
    layer2_outputs(3597) <= not a or b;
    layer2_outputs(3598) <= a and b;
    layer2_outputs(3599) <= a;
    layer2_outputs(3600) <= not (a or b);
    layer2_outputs(3601) <= not (a and b);
    layer2_outputs(3602) <= a and b;
    layer2_outputs(3603) <= not (a and b);
    layer2_outputs(3604) <= not (a or b);
    layer2_outputs(3605) <= '1';
    layer2_outputs(3606) <= a;
    layer2_outputs(3607) <= a;
    layer2_outputs(3608) <= b and not a;
    layer2_outputs(3609) <= not a;
    layer2_outputs(3610) <= b;
    layer2_outputs(3611) <= a and b;
    layer2_outputs(3612) <= not (a or b);
    layer2_outputs(3613) <= not a;
    layer2_outputs(3614) <= not (a or b);
    layer2_outputs(3615) <= not a;
    layer2_outputs(3616) <= not b;
    layer2_outputs(3617) <= '0';
    layer2_outputs(3618) <= a and not b;
    layer2_outputs(3619) <= a and b;
    layer2_outputs(3620) <= not a or b;
    layer2_outputs(3621) <= '1';
    layer2_outputs(3622) <= not a or b;
    layer2_outputs(3623) <= b and not a;
    layer2_outputs(3624) <= b and not a;
    layer2_outputs(3625) <= not a or b;
    layer2_outputs(3626) <= '0';
    layer2_outputs(3627) <= not b;
    layer2_outputs(3628) <= not b;
    layer2_outputs(3629) <= not a or b;
    layer2_outputs(3630) <= '0';
    layer2_outputs(3631) <= not a or b;
    layer2_outputs(3632) <= '0';
    layer2_outputs(3633) <= not b or a;
    layer2_outputs(3634) <= b and not a;
    layer2_outputs(3635) <= not a or b;
    layer2_outputs(3636) <= not b or a;
    layer2_outputs(3637) <= b and not a;
    layer2_outputs(3638) <= a xor b;
    layer2_outputs(3639) <= a and b;
    layer2_outputs(3640) <= not b;
    layer2_outputs(3641) <= '0';
    layer2_outputs(3642) <= not a or b;
    layer2_outputs(3643) <= a and b;
    layer2_outputs(3644) <= a and not b;
    layer2_outputs(3645) <= b and not a;
    layer2_outputs(3646) <= '0';
    layer2_outputs(3647) <= b;
    layer2_outputs(3648) <= not a or b;
    layer2_outputs(3649) <= not a;
    layer2_outputs(3650) <= '1';
    layer2_outputs(3651) <= not (a or b);
    layer2_outputs(3652) <= a and not b;
    layer2_outputs(3653) <= b;
    layer2_outputs(3654) <= not (a or b);
    layer2_outputs(3655) <= a xor b;
    layer2_outputs(3656) <= b;
    layer2_outputs(3657) <= b and not a;
    layer2_outputs(3658) <= not b or a;
    layer2_outputs(3659) <= '1';
    layer2_outputs(3660) <= not b or a;
    layer2_outputs(3661) <= a or b;
    layer2_outputs(3662) <= b;
    layer2_outputs(3663) <= a or b;
    layer2_outputs(3664) <= not (a and b);
    layer2_outputs(3665) <= not a;
    layer2_outputs(3666) <= not (a and b);
    layer2_outputs(3667) <= not b;
    layer2_outputs(3668) <= not b;
    layer2_outputs(3669) <= not (a or b);
    layer2_outputs(3670) <= a or b;
    layer2_outputs(3671) <= not (a xor b);
    layer2_outputs(3672) <= a;
    layer2_outputs(3673) <= not (a or b);
    layer2_outputs(3674) <= '0';
    layer2_outputs(3675) <= not (a or b);
    layer2_outputs(3676) <= not a;
    layer2_outputs(3677) <= '0';
    layer2_outputs(3678) <= not a or b;
    layer2_outputs(3679) <= '1';
    layer2_outputs(3680) <= not (a xor b);
    layer2_outputs(3681) <= a or b;
    layer2_outputs(3682) <= '1';
    layer2_outputs(3683) <= not b or a;
    layer2_outputs(3684) <= a and not b;
    layer2_outputs(3685) <= b and not a;
    layer2_outputs(3686) <= not a;
    layer2_outputs(3687) <= a or b;
    layer2_outputs(3688) <= not b;
    layer2_outputs(3689) <= '0';
    layer2_outputs(3690) <= '1';
    layer2_outputs(3691) <= not a or b;
    layer2_outputs(3692) <= b;
    layer2_outputs(3693) <= not (a or b);
    layer2_outputs(3694) <= not b;
    layer2_outputs(3695) <= '1';
    layer2_outputs(3696) <= '0';
    layer2_outputs(3697) <= '1';
    layer2_outputs(3698) <= not (a and b);
    layer2_outputs(3699) <= a and b;
    layer2_outputs(3700) <= '1';
    layer2_outputs(3701) <= '1';
    layer2_outputs(3702) <= a xor b;
    layer2_outputs(3703) <= not (a xor b);
    layer2_outputs(3704) <= '0';
    layer2_outputs(3705) <= a;
    layer2_outputs(3706) <= '0';
    layer2_outputs(3707) <= '1';
    layer2_outputs(3708) <= a;
    layer2_outputs(3709) <= not a or b;
    layer2_outputs(3710) <= a;
    layer2_outputs(3711) <= '1';
    layer2_outputs(3712) <= not (a xor b);
    layer2_outputs(3713) <= not b or a;
    layer2_outputs(3714) <= not (a or b);
    layer2_outputs(3715) <= '0';
    layer2_outputs(3716) <= a and b;
    layer2_outputs(3717) <= not (a or b);
    layer2_outputs(3718) <= a;
    layer2_outputs(3719) <= not (a and b);
    layer2_outputs(3720) <= not b or a;
    layer2_outputs(3721) <= b and not a;
    layer2_outputs(3722) <= not (a and b);
    layer2_outputs(3723) <= '1';
    layer2_outputs(3724) <= not b;
    layer2_outputs(3725) <= not a;
    layer2_outputs(3726) <= not a;
    layer2_outputs(3727) <= not (a xor b);
    layer2_outputs(3728) <= a and not b;
    layer2_outputs(3729) <= '1';
    layer2_outputs(3730) <= '1';
    layer2_outputs(3731) <= '0';
    layer2_outputs(3732) <= b and not a;
    layer2_outputs(3733) <= not b;
    layer2_outputs(3734) <= not (a or b);
    layer2_outputs(3735) <= '1';
    layer2_outputs(3736) <= '1';
    layer2_outputs(3737) <= not b;
    layer2_outputs(3738) <= a and not b;
    layer2_outputs(3739) <= '0';
    layer2_outputs(3740) <= b and not a;
    layer2_outputs(3741) <= not (a and b);
    layer2_outputs(3742) <= a;
    layer2_outputs(3743) <= not a or b;
    layer2_outputs(3744) <= a or b;
    layer2_outputs(3745) <= a or b;
    layer2_outputs(3746) <= a and b;
    layer2_outputs(3747) <= b and not a;
    layer2_outputs(3748) <= '1';
    layer2_outputs(3749) <= a and b;
    layer2_outputs(3750) <= '1';
    layer2_outputs(3751) <= '0';
    layer2_outputs(3752) <= '1';
    layer2_outputs(3753) <= not a;
    layer2_outputs(3754) <= not a;
    layer2_outputs(3755) <= not b;
    layer2_outputs(3756) <= not a;
    layer2_outputs(3757) <= not b or a;
    layer2_outputs(3758) <= '0';
    layer2_outputs(3759) <= b and not a;
    layer2_outputs(3760) <= '1';
    layer2_outputs(3761) <= not a or b;
    layer2_outputs(3762) <= b and not a;
    layer2_outputs(3763) <= not (a and b);
    layer2_outputs(3764) <= a and not b;
    layer2_outputs(3765) <= a xor b;
    layer2_outputs(3766) <= not b;
    layer2_outputs(3767) <= not b;
    layer2_outputs(3768) <= not (a or b);
    layer2_outputs(3769) <= a and not b;
    layer2_outputs(3770) <= a or b;
    layer2_outputs(3771) <= a and b;
    layer2_outputs(3772) <= b;
    layer2_outputs(3773) <= not a or b;
    layer2_outputs(3774) <= a or b;
    layer2_outputs(3775) <= not (a and b);
    layer2_outputs(3776) <= a xor b;
    layer2_outputs(3777) <= a and not b;
    layer2_outputs(3778) <= not b;
    layer2_outputs(3779) <= '1';
    layer2_outputs(3780) <= a or b;
    layer2_outputs(3781) <= not b;
    layer2_outputs(3782) <= b and not a;
    layer2_outputs(3783) <= b;
    layer2_outputs(3784) <= b;
    layer2_outputs(3785) <= not b;
    layer2_outputs(3786) <= not b;
    layer2_outputs(3787) <= '0';
    layer2_outputs(3788) <= b;
    layer2_outputs(3789) <= not b or a;
    layer2_outputs(3790) <= not b;
    layer2_outputs(3791) <= not (a or b);
    layer2_outputs(3792) <= '1';
    layer2_outputs(3793) <= b and not a;
    layer2_outputs(3794) <= a or b;
    layer2_outputs(3795) <= a and not b;
    layer2_outputs(3796) <= not (a or b);
    layer2_outputs(3797) <= not b;
    layer2_outputs(3798) <= a or b;
    layer2_outputs(3799) <= not (a and b);
    layer2_outputs(3800) <= '0';
    layer2_outputs(3801) <= b and not a;
    layer2_outputs(3802) <= not (a and b);
    layer2_outputs(3803) <= not a;
    layer2_outputs(3804) <= not (a and b);
    layer2_outputs(3805) <= not a or b;
    layer2_outputs(3806) <= '0';
    layer2_outputs(3807) <= not (a and b);
    layer2_outputs(3808) <= not a;
    layer2_outputs(3809) <= a;
    layer2_outputs(3810) <= a or b;
    layer2_outputs(3811) <= '0';
    layer2_outputs(3812) <= not b;
    layer2_outputs(3813) <= not a or b;
    layer2_outputs(3814) <= not (a or b);
    layer2_outputs(3815) <= '1';
    layer2_outputs(3816) <= '1';
    layer2_outputs(3817) <= '1';
    layer2_outputs(3818) <= not b or a;
    layer2_outputs(3819) <= not (a or b);
    layer2_outputs(3820) <= not (a and b);
    layer2_outputs(3821) <= a or b;
    layer2_outputs(3822) <= b;
    layer2_outputs(3823) <= '0';
    layer2_outputs(3824) <= not (a and b);
    layer2_outputs(3825) <= not (a and b);
    layer2_outputs(3826) <= a and not b;
    layer2_outputs(3827) <= not (a and b);
    layer2_outputs(3828) <= a;
    layer2_outputs(3829) <= not b or a;
    layer2_outputs(3830) <= b and not a;
    layer2_outputs(3831) <= not a or b;
    layer2_outputs(3832) <= a xor b;
    layer2_outputs(3833) <= not a;
    layer2_outputs(3834) <= a;
    layer2_outputs(3835) <= not b or a;
    layer2_outputs(3836) <= not (a and b);
    layer2_outputs(3837) <= not (a xor b);
    layer2_outputs(3838) <= not a or b;
    layer2_outputs(3839) <= b;
    layer2_outputs(3840) <= '1';
    layer2_outputs(3841) <= not b;
    layer2_outputs(3842) <= a and not b;
    layer2_outputs(3843) <= '0';
    layer2_outputs(3844) <= '0';
    layer2_outputs(3845) <= a or b;
    layer2_outputs(3846) <= not b;
    layer2_outputs(3847) <= '1';
    layer2_outputs(3848) <= not b;
    layer2_outputs(3849) <= '1';
    layer2_outputs(3850) <= a and not b;
    layer2_outputs(3851) <= '1';
    layer2_outputs(3852) <= not (a xor b);
    layer2_outputs(3853) <= '1';
    layer2_outputs(3854) <= not a;
    layer2_outputs(3855) <= not b;
    layer2_outputs(3856) <= '0';
    layer2_outputs(3857) <= '1';
    layer2_outputs(3858) <= not b or a;
    layer2_outputs(3859) <= a and not b;
    layer2_outputs(3860) <= '1';
    layer2_outputs(3861) <= not a or b;
    layer2_outputs(3862) <= a and not b;
    layer2_outputs(3863) <= not a;
    layer2_outputs(3864) <= a;
    layer2_outputs(3865) <= not (a and b);
    layer2_outputs(3866) <= '1';
    layer2_outputs(3867) <= '1';
    layer2_outputs(3868) <= b and not a;
    layer2_outputs(3869) <= a and not b;
    layer2_outputs(3870) <= a;
    layer2_outputs(3871) <= not (a and b);
    layer2_outputs(3872) <= b;
    layer2_outputs(3873) <= a and not b;
    layer2_outputs(3874) <= a;
    layer2_outputs(3875) <= not (a or b);
    layer2_outputs(3876) <= not (a or b);
    layer2_outputs(3877) <= not a or b;
    layer2_outputs(3878) <= not (a and b);
    layer2_outputs(3879) <= a or b;
    layer2_outputs(3880) <= a and b;
    layer2_outputs(3881) <= not (a and b);
    layer2_outputs(3882) <= a;
    layer2_outputs(3883) <= '0';
    layer2_outputs(3884) <= not (a or b);
    layer2_outputs(3885) <= b;
    layer2_outputs(3886) <= not (a and b);
    layer2_outputs(3887) <= a and b;
    layer2_outputs(3888) <= b and not a;
    layer2_outputs(3889) <= '1';
    layer2_outputs(3890) <= '0';
    layer2_outputs(3891) <= a and not b;
    layer2_outputs(3892) <= '1';
    layer2_outputs(3893) <= not (a xor b);
    layer2_outputs(3894) <= not (a and b);
    layer2_outputs(3895) <= not a or b;
    layer2_outputs(3896) <= a;
    layer2_outputs(3897) <= b;
    layer2_outputs(3898) <= not (a or b);
    layer2_outputs(3899) <= b;
    layer2_outputs(3900) <= not (a and b);
    layer2_outputs(3901) <= b and not a;
    layer2_outputs(3902) <= b and not a;
    layer2_outputs(3903) <= b;
    layer2_outputs(3904) <= not b;
    layer2_outputs(3905) <= not a or b;
    layer2_outputs(3906) <= not (a or b);
    layer2_outputs(3907) <= not a;
    layer2_outputs(3908) <= b and not a;
    layer2_outputs(3909) <= a or b;
    layer2_outputs(3910) <= a xor b;
    layer2_outputs(3911) <= not a;
    layer2_outputs(3912) <= a and not b;
    layer2_outputs(3913) <= a or b;
    layer2_outputs(3914) <= b and not a;
    layer2_outputs(3915) <= '0';
    layer2_outputs(3916) <= not (a and b);
    layer2_outputs(3917) <= not b or a;
    layer2_outputs(3918) <= b and not a;
    layer2_outputs(3919) <= a or b;
    layer2_outputs(3920) <= not a;
    layer2_outputs(3921) <= '1';
    layer2_outputs(3922) <= not a;
    layer2_outputs(3923) <= a and b;
    layer2_outputs(3924) <= not (a xor b);
    layer2_outputs(3925) <= a and b;
    layer2_outputs(3926) <= not a;
    layer2_outputs(3927) <= not a or b;
    layer2_outputs(3928) <= a and not b;
    layer2_outputs(3929) <= not b;
    layer2_outputs(3930) <= '1';
    layer2_outputs(3931) <= not b;
    layer2_outputs(3932) <= a and b;
    layer2_outputs(3933) <= not (a or b);
    layer2_outputs(3934) <= '0';
    layer2_outputs(3935) <= '1';
    layer2_outputs(3936) <= a or b;
    layer2_outputs(3937) <= not (a xor b);
    layer2_outputs(3938) <= b;
    layer2_outputs(3939) <= a and b;
    layer2_outputs(3940) <= not (a and b);
    layer2_outputs(3941) <= not (a or b);
    layer2_outputs(3942) <= not b or a;
    layer2_outputs(3943) <= '0';
    layer2_outputs(3944) <= a and b;
    layer2_outputs(3945) <= a and b;
    layer2_outputs(3946) <= not b;
    layer2_outputs(3947) <= b;
    layer2_outputs(3948) <= a xor b;
    layer2_outputs(3949) <= not (a or b);
    layer2_outputs(3950) <= '1';
    layer2_outputs(3951) <= a and b;
    layer2_outputs(3952) <= a or b;
    layer2_outputs(3953) <= '1';
    layer2_outputs(3954) <= a and not b;
    layer2_outputs(3955) <= not (a or b);
    layer2_outputs(3956) <= not b;
    layer2_outputs(3957) <= not b or a;
    layer2_outputs(3958) <= '0';
    layer2_outputs(3959) <= b;
    layer2_outputs(3960) <= '0';
    layer2_outputs(3961) <= a and b;
    layer2_outputs(3962) <= a or b;
    layer2_outputs(3963) <= b and not a;
    layer2_outputs(3964) <= not (a xor b);
    layer2_outputs(3965) <= not (a and b);
    layer2_outputs(3966) <= not b or a;
    layer2_outputs(3967) <= '0';
    layer2_outputs(3968) <= a;
    layer2_outputs(3969) <= not b or a;
    layer2_outputs(3970) <= b and not a;
    layer2_outputs(3971) <= a;
    layer2_outputs(3972) <= not (a and b);
    layer2_outputs(3973) <= not a;
    layer2_outputs(3974) <= b and not a;
    layer2_outputs(3975) <= not b or a;
    layer2_outputs(3976) <= a or b;
    layer2_outputs(3977) <= a and not b;
    layer2_outputs(3978) <= '0';
    layer2_outputs(3979) <= a and not b;
    layer2_outputs(3980) <= not b;
    layer2_outputs(3981) <= b and not a;
    layer2_outputs(3982) <= not a;
    layer2_outputs(3983) <= not a or b;
    layer2_outputs(3984) <= a or b;
    layer2_outputs(3985) <= b;
    layer2_outputs(3986) <= '0';
    layer2_outputs(3987) <= a or b;
    layer2_outputs(3988) <= b and not a;
    layer2_outputs(3989) <= '0';
    layer2_outputs(3990) <= a and not b;
    layer2_outputs(3991) <= a;
    layer2_outputs(3992) <= not a or b;
    layer2_outputs(3993) <= not a;
    layer2_outputs(3994) <= a;
    layer2_outputs(3995) <= b and not a;
    layer2_outputs(3996) <= '0';
    layer2_outputs(3997) <= not (a or b);
    layer2_outputs(3998) <= a and b;
    layer2_outputs(3999) <= not b;
    layer2_outputs(4000) <= '1';
    layer2_outputs(4001) <= not a or b;
    layer2_outputs(4002) <= not (a or b);
    layer2_outputs(4003) <= not (a and b);
    layer2_outputs(4004) <= b;
    layer2_outputs(4005) <= not (a or b);
    layer2_outputs(4006) <= b;
    layer2_outputs(4007) <= not b or a;
    layer2_outputs(4008) <= not (a xor b);
    layer2_outputs(4009) <= not a;
    layer2_outputs(4010) <= not b or a;
    layer2_outputs(4011) <= a and not b;
    layer2_outputs(4012) <= a xor b;
    layer2_outputs(4013) <= a;
    layer2_outputs(4014) <= a and not b;
    layer2_outputs(4015) <= a or b;
    layer2_outputs(4016) <= not a or b;
    layer2_outputs(4017) <= a and not b;
    layer2_outputs(4018) <= a or b;
    layer2_outputs(4019) <= not a or b;
    layer2_outputs(4020) <= a;
    layer2_outputs(4021) <= a or b;
    layer2_outputs(4022) <= '0';
    layer2_outputs(4023) <= a xor b;
    layer2_outputs(4024) <= not a;
    layer2_outputs(4025) <= a;
    layer2_outputs(4026) <= a and b;
    layer2_outputs(4027) <= not a;
    layer2_outputs(4028) <= b;
    layer2_outputs(4029) <= a and not b;
    layer2_outputs(4030) <= not a;
    layer2_outputs(4031) <= not (a or b);
    layer2_outputs(4032) <= not a;
    layer2_outputs(4033) <= a and not b;
    layer2_outputs(4034) <= not a or b;
    layer2_outputs(4035) <= a and b;
    layer2_outputs(4036) <= '1';
    layer2_outputs(4037) <= b and not a;
    layer2_outputs(4038) <= not (a and b);
    layer2_outputs(4039) <= not b;
    layer2_outputs(4040) <= a and not b;
    layer2_outputs(4041) <= '1';
    layer2_outputs(4042) <= a or b;
    layer2_outputs(4043) <= '1';
    layer2_outputs(4044) <= not (a or b);
    layer2_outputs(4045) <= a;
    layer2_outputs(4046) <= b;
    layer2_outputs(4047) <= a or b;
    layer2_outputs(4048) <= not (a and b);
    layer2_outputs(4049) <= b;
    layer2_outputs(4050) <= a or b;
    layer2_outputs(4051) <= not b or a;
    layer2_outputs(4052) <= not a or b;
    layer2_outputs(4053) <= not a;
    layer2_outputs(4054) <= a and not b;
    layer2_outputs(4055) <= not (a or b);
    layer2_outputs(4056) <= not a;
    layer2_outputs(4057) <= a or b;
    layer2_outputs(4058) <= not b;
    layer2_outputs(4059) <= a and b;
    layer2_outputs(4060) <= a and not b;
    layer2_outputs(4061) <= not a or b;
    layer2_outputs(4062) <= not (a or b);
    layer2_outputs(4063) <= not (a and b);
    layer2_outputs(4064) <= a and b;
    layer2_outputs(4065) <= not (a and b);
    layer2_outputs(4066) <= b and not a;
    layer2_outputs(4067) <= '1';
    layer2_outputs(4068) <= a and not b;
    layer2_outputs(4069) <= a;
    layer2_outputs(4070) <= '1';
    layer2_outputs(4071) <= not (a or b);
    layer2_outputs(4072) <= a and not b;
    layer2_outputs(4073) <= a or b;
    layer2_outputs(4074) <= not (a or b);
    layer2_outputs(4075) <= not (a and b);
    layer2_outputs(4076) <= not b or a;
    layer2_outputs(4077) <= b;
    layer2_outputs(4078) <= '0';
    layer2_outputs(4079) <= not b;
    layer2_outputs(4080) <= a and b;
    layer2_outputs(4081) <= a;
    layer2_outputs(4082) <= '0';
    layer2_outputs(4083) <= not b;
    layer2_outputs(4084) <= a and not b;
    layer2_outputs(4085) <= b and not a;
    layer2_outputs(4086) <= not b;
    layer2_outputs(4087) <= a and b;
    layer2_outputs(4088) <= not b;
    layer2_outputs(4089) <= not a;
    layer2_outputs(4090) <= not (a and b);
    layer2_outputs(4091) <= '1';
    layer2_outputs(4092) <= not b or a;
    layer2_outputs(4093) <= not b or a;
    layer2_outputs(4094) <= a or b;
    layer2_outputs(4095) <= not (a and b);
    layer2_outputs(4096) <= not (a and b);
    layer2_outputs(4097) <= a and not b;
    layer2_outputs(4098) <= b;
    layer2_outputs(4099) <= not b or a;
    layer2_outputs(4100) <= a or b;
    layer2_outputs(4101) <= not b or a;
    layer2_outputs(4102) <= a or b;
    layer2_outputs(4103) <= not b;
    layer2_outputs(4104) <= not b;
    layer2_outputs(4105) <= not a or b;
    layer2_outputs(4106) <= not (a xor b);
    layer2_outputs(4107) <= not (a or b);
    layer2_outputs(4108) <= a;
    layer2_outputs(4109) <= not b;
    layer2_outputs(4110) <= a and b;
    layer2_outputs(4111) <= '0';
    layer2_outputs(4112) <= not (a and b);
    layer2_outputs(4113) <= not (a or b);
    layer2_outputs(4114) <= '0';
    layer2_outputs(4115) <= not a;
    layer2_outputs(4116) <= not (a or b);
    layer2_outputs(4117) <= a and b;
    layer2_outputs(4118) <= not (a xor b);
    layer2_outputs(4119) <= '1';
    layer2_outputs(4120) <= b;
    layer2_outputs(4121) <= not a or b;
    layer2_outputs(4122) <= b and not a;
    layer2_outputs(4123) <= '0';
    layer2_outputs(4124) <= '0';
    layer2_outputs(4125) <= a and not b;
    layer2_outputs(4126) <= '1';
    layer2_outputs(4127) <= b and not a;
    layer2_outputs(4128) <= a and b;
    layer2_outputs(4129) <= b;
    layer2_outputs(4130) <= not a;
    layer2_outputs(4131) <= not (a or b);
    layer2_outputs(4132) <= not b or a;
    layer2_outputs(4133) <= not a or b;
    layer2_outputs(4134) <= b;
    layer2_outputs(4135) <= '1';
    layer2_outputs(4136) <= not b;
    layer2_outputs(4137) <= '0';
    layer2_outputs(4138) <= b and not a;
    layer2_outputs(4139) <= a and b;
    layer2_outputs(4140) <= not (a or b);
    layer2_outputs(4141) <= not (a and b);
    layer2_outputs(4142) <= '1';
    layer2_outputs(4143) <= not a;
    layer2_outputs(4144) <= '0';
    layer2_outputs(4145) <= a and not b;
    layer2_outputs(4146) <= a;
    layer2_outputs(4147) <= not b;
    layer2_outputs(4148) <= '1';
    layer2_outputs(4149) <= b;
    layer2_outputs(4150) <= not b;
    layer2_outputs(4151) <= not (a and b);
    layer2_outputs(4152) <= b;
    layer2_outputs(4153) <= not (a or b);
    layer2_outputs(4154) <= '0';
    layer2_outputs(4155) <= b;
    layer2_outputs(4156) <= '1';
    layer2_outputs(4157) <= a xor b;
    layer2_outputs(4158) <= b;
    layer2_outputs(4159) <= a and not b;
    layer2_outputs(4160) <= b;
    layer2_outputs(4161) <= '0';
    layer2_outputs(4162) <= not (a and b);
    layer2_outputs(4163) <= not b or a;
    layer2_outputs(4164) <= '0';
    layer2_outputs(4165) <= a;
    layer2_outputs(4166) <= a or b;
    layer2_outputs(4167) <= not (a or b);
    layer2_outputs(4168) <= not (a or b);
    layer2_outputs(4169) <= not b;
    layer2_outputs(4170) <= not (a xor b);
    layer2_outputs(4171) <= not a or b;
    layer2_outputs(4172) <= not b or a;
    layer2_outputs(4173) <= not (a and b);
    layer2_outputs(4174) <= a and b;
    layer2_outputs(4175) <= not b or a;
    layer2_outputs(4176) <= '0';
    layer2_outputs(4177) <= not b;
    layer2_outputs(4178) <= b;
    layer2_outputs(4179) <= a and not b;
    layer2_outputs(4180) <= not (a or b);
    layer2_outputs(4181) <= a and not b;
    layer2_outputs(4182) <= '1';
    layer2_outputs(4183) <= a and not b;
    layer2_outputs(4184) <= not (a xor b);
    layer2_outputs(4185) <= '1';
    layer2_outputs(4186) <= not b or a;
    layer2_outputs(4187) <= not (a or b);
    layer2_outputs(4188) <= not b;
    layer2_outputs(4189) <= not a;
    layer2_outputs(4190) <= a;
    layer2_outputs(4191) <= '0';
    layer2_outputs(4192) <= a and not b;
    layer2_outputs(4193) <= a and b;
    layer2_outputs(4194) <= '0';
    layer2_outputs(4195) <= not b;
    layer2_outputs(4196) <= '1';
    layer2_outputs(4197) <= a;
    layer2_outputs(4198) <= '0';
    layer2_outputs(4199) <= not a;
    layer2_outputs(4200) <= a or b;
    layer2_outputs(4201) <= not (a or b);
    layer2_outputs(4202) <= not b;
    layer2_outputs(4203) <= '1';
    layer2_outputs(4204) <= not (a or b);
    layer2_outputs(4205) <= not a or b;
    layer2_outputs(4206) <= not (a or b);
    layer2_outputs(4207) <= not b or a;
    layer2_outputs(4208) <= not a or b;
    layer2_outputs(4209) <= a or b;
    layer2_outputs(4210) <= a and not b;
    layer2_outputs(4211) <= not (a or b);
    layer2_outputs(4212) <= not b or a;
    layer2_outputs(4213) <= a;
    layer2_outputs(4214) <= not (a or b);
    layer2_outputs(4215) <= not (a or b);
    layer2_outputs(4216) <= a and not b;
    layer2_outputs(4217) <= '0';
    layer2_outputs(4218) <= a or b;
    layer2_outputs(4219) <= a and b;
    layer2_outputs(4220) <= a or b;
    layer2_outputs(4221) <= not (a and b);
    layer2_outputs(4222) <= b;
    layer2_outputs(4223) <= '0';
    layer2_outputs(4224) <= a;
    layer2_outputs(4225) <= not (a and b);
    layer2_outputs(4226) <= '0';
    layer2_outputs(4227) <= a xor b;
    layer2_outputs(4228) <= '0';
    layer2_outputs(4229) <= not a or b;
    layer2_outputs(4230) <= not (a and b);
    layer2_outputs(4231) <= not (a and b);
    layer2_outputs(4232) <= b and not a;
    layer2_outputs(4233) <= not b;
    layer2_outputs(4234) <= not b;
    layer2_outputs(4235) <= not (a and b);
    layer2_outputs(4236) <= not b or a;
    layer2_outputs(4237) <= '0';
    layer2_outputs(4238) <= '1';
    layer2_outputs(4239) <= not a or b;
    layer2_outputs(4240) <= '0';
    layer2_outputs(4241) <= b;
    layer2_outputs(4242) <= a and b;
    layer2_outputs(4243) <= b;
    layer2_outputs(4244) <= not a or b;
    layer2_outputs(4245) <= not b;
    layer2_outputs(4246) <= not (a or b);
    layer2_outputs(4247) <= '1';
    layer2_outputs(4248) <= not b or a;
    layer2_outputs(4249) <= '0';
    layer2_outputs(4250) <= not b;
    layer2_outputs(4251) <= not (a or b);
    layer2_outputs(4252) <= not (a or b);
    layer2_outputs(4253) <= not (a or b);
    layer2_outputs(4254) <= not (a and b);
    layer2_outputs(4255) <= not (a and b);
    layer2_outputs(4256) <= not (a and b);
    layer2_outputs(4257) <= not b;
    layer2_outputs(4258) <= a;
    layer2_outputs(4259) <= '0';
    layer2_outputs(4260) <= b and not a;
    layer2_outputs(4261) <= a or b;
    layer2_outputs(4262) <= '0';
    layer2_outputs(4263) <= a and not b;
    layer2_outputs(4264) <= not (a and b);
    layer2_outputs(4265) <= '1';
    layer2_outputs(4266) <= a and not b;
    layer2_outputs(4267) <= '1';
    layer2_outputs(4268) <= a and not b;
    layer2_outputs(4269) <= not (a and b);
    layer2_outputs(4270) <= not a;
    layer2_outputs(4271) <= a or b;
    layer2_outputs(4272) <= a and b;
    layer2_outputs(4273) <= not a or b;
    layer2_outputs(4274) <= '1';
    layer2_outputs(4275) <= not a or b;
    layer2_outputs(4276) <= '0';
    layer2_outputs(4277) <= not a or b;
    layer2_outputs(4278) <= not a;
    layer2_outputs(4279) <= a or b;
    layer2_outputs(4280) <= a and b;
    layer2_outputs(4281) <= '1';
    layer2_outputs(4282) <= a xor b;
    layer2_outputs(4283) <= a or b;
    layer2_outputs(4284) <= a or b;
    layer2_outputs(4285) <= b;
    layer2_outputs(4286) <= '0';
    layer2_outputs(4287) <= '1';
    layer2_outputs(4288) <= not b;
    layer2_outputs(4289) <= not b or a;
    layer2_outputs(4290) <= '1';
    layer2_outputs(4291) <= not (a and b);
    layer2_outputs(4292) <= not (a or b);
    layer2_outputs(4293) <= not b;
    layer2_outputs(4294) <= a and not b;
    layer2_outputs(4295) <= not a;
    layer2_outputs(4296) <= '1';
    layer2_outputs(4297) <= a;
    layer2_outputs(4298) <= not b;
    layer2_outputs(4299) <= not (a and b);
    layer2_outputs(4300) <= not (a and b);
    layer2_outputs(4301) <= not (a or b);
    layer2_outputs(4302) <= not a;
    layer2_outputs(4303) <= not b or a;
    layer2_outputs(4304) <= not (a or b);
    layer2_outputs(4305) <= not (a or b);
    layer2_outputs(4306) <= not b or a;
    layer2_outputs(4307) <= not a or b;
    layer2_outputs(4308) <= a or b;
    layer2_outputs(4309) <= '1';
    layer2_outputs(4310) <= b and not a;
    layer2_outputs(4311) <= not (a and b);
    layer2_outputs(4312) <= not (a and b);
    layer2_outputs(4313) <= not a;
    layer2_outputs(4314) <= a or b;
    layer2_outputs(4315) <= not b or a;
    layer2_outputs(4316) <= a and b;
    layer2_outputs(4317) <= not b or a;
    layer2_outputs(4318) <= a or b;
    layer2_outputs(4319) <= a and b;
    layer2_outputs(4320) <= a or b;
    layer2_outputs(4321) <= not (a and b);
    layer2_outputs(4322) <= b;
    layer2_outputs(4323) <= '0';
    layer2_outputs(4324) <= not b;
    layer2_outputs(4325) <= '1';
    layer2_outputs(4326) <= a and not b;
    layer2_outputs(4327) <= not a;
    layer2_outputs(4328) <= not a;
    layer2_outputs(4329) <= not (a or b);
    layer2_outputs(4330) <= not b;
    layer2_outputs(4331) <= a or b;
    layer2_outputs(4332) <= b;
    layer2_outputs(4333) <= b and not a;
    layer2_outputs(4334) <= a;
    layer2_outputs(4335) <= a and not b;
    layer2_outputs(4336) <= a or b;
    layer2_outputs(4337) <= not b;
    layer2_outputs(4338) <= a or b;
    layer2_outputs(4339) <= not (a or b);
    layer2_outputs(4340) <= '0';
    layer2_outputs(4341) <= not (a or b);
    layer2_outputs(4342) <= not b or a;
    layer2_outputs(4343) <= not a or b;
    layer2_outputs(4344) <= '0';
    layer2_outputs(4345) <= not (a and b);
    layer2_outputs(4346) <= '0';
    layer2_outputs(4347) <= b;
    layer2_outputs(4348) <= '1';
    layer2_outputs(4349) <= a;
    layer2_outputs(4350) <= '0';
    layer2_outputs(4351) <= a;
    layer2_outputs(4352) <= b and not a;
    layer2_outputs(4353) <= '0';
    layer2_outputs(4354) <= not a or b;
    layer2_outputs(4355) <= a and b;
    layer2_outputs(4356) <= b;
    layer2_outputs(4357) <= not b;
    layer2_outputs(4358) <= b and not a;
    layer2_outputs(4359) <= '0';
    layer2_outputs(4360) <= not (a and b);
    layer2_outputs(4361) <= not a or b;
    layer2_outputs(4362) <= a;
    layer2_outputs(4363) <= '1';
    layer2_outputs(4364) <= a;
    layer2_outputs(4365) <= '0';
    layer2_outputs(4366) <= '1';
    layer2_outputs(4367) <= not (a and b);
    layer2_outputs(4368) <= not (a and b);
    layer2_outputs(4369) <= a;
    layer2_outputs(4370) <= a;
    layer2_outputs(4371) <= not (a and b);
    layer2_outputs(4372) <= not a;
    layer2_outputs(4373) <= not a;
    layer2_outputs(4374) <= b;
    layer2_outputs(4375) <= not (a and b);
    layer2_outputs(4376) <= not (a or b);
    layer2_outputs(4377) <= not a;
    layer2_outputs(4378) <= '0';
    layer2_outputs(4379) <= a and b;
    layer2_outputs(4380) <= not a;
    layer2_outputs(4381) <= a and b;
    layer2_outputs(4382) <= b and not a;
    layer2_outputs(4383) <= '1';
    layer2_outputs(4384) <= not b;
    layer2_outputs(4385) <= '1';
    layer2_outputs(4386) <= '0';
    layer2_outputs(4387) <= b and not a;
    layer2_outputs(4388) <= '1';
    layer2_outputs(4389) <= not (a or b);
    layer2_outputs(4390) <= a and b;
    layer2_outputs(4391) <= '1';
    layer2_outputs(4392) <= not (a and b);
    layer2_outputs(4393) <= not (a or b);
    layer2_outputs(4394) <= b and not a;
    layer2_outputs(4395) <= not b;
    layer2_outputs(4396) <= not (a or b);
    layer2_outputs(4397) <= '0';
    layer2_outputs(4398) <= a and not b;
    layer2_outputs(4399) <= '1';
    layer2_outputs(4400) <= not a;
    layer2_outputs(4401) <= '0';
    layer2_outputs(4402) <= a or b;
    layer2_outputs(4403) <= a or b;
    layer2_outputs(4404) <= not b;
    layer2_outputs(4405) <= not b;
    layer2_outputs(4406) <= '1';
    layer2_outputs(4407) <= a xor b;
    layer2_outputs(4408) <= not (a or b);
    layer2_outputs(4409) <= not b;
    layer2_outputs(4410) <= '1';
    layer2_outputs(4411) <= not (a or b);
    layer2_outputs(4412) <= b and not a;
    layer2_outputs(4413) <= not a;
    layer2_outputs(4414) <= not b or a;
    layer2_outputs(4415) <= b and not a;
    layer2_outputs(4416) <= not b;
    layer2_outputs(4417) <= not b or a;
    layer2_outputs(4418) <= a xor b;
    layer2_outputs(4419) <= '0';
    layer2_outputs(4420) <= not b;
    layer2_outputs(4421) <= a xor b;
    layer2_outputs(4422) <= b;
    layer2_outputs(4423) <= a or b;
    layer2_outputs(4424) <= '1';
    layer2_outputs(4425) <= '1';
    layer2_outputs(4426) <= a;
    layer2_outputs(4427) <= '1';
    layer2_outputs(4428) <= not b or a;
    layer2_outputs(4429) <= not (a and b);
    layer2_outputs(4430) <= not (a or b);
    layer2_outputs(4431) <= not a;
    layer2_outputs(4432) <= not a;
    layer2_outputs(4433) <= a;
    layer2_outputs(4434) <= '0';
    layer2_outputs(4435) <= a;
    layer2_outputs(4436) <= not a or b;
    layer2_outputs(4437) <= not (a or b);
    layer2_outputs(4438) <= not b or a;
    layer2_outputs(4439) <= a and b;
    layer2_outputs(4440) <= not (a or b);
    layer2_outputs(4441) <= not (a or b);
    layer2_outputs(4442) <= not a or b;
    layer2_outputs(4443) <= a and not b;
    layer2_outputs(4444) <= '1';
    layer2_outputs(4445) <= not (a or b);
    layer2_outputs(4446) <= b and not a;
    layer2_outputs(4447) <= b and not a;
    layer2_outputs(4448) <= a and b;
    layer2_outputs(4449) <= not b;
    layer2_outputs(4450) <= not a;
    layer2_outputs(4451) <= not b or a;
    layer2_outputs(4452) <= a or b;
    layer2_outputs(4453) <= '1';
    layer2_outputs(4454) <= not a or b;
    layer2_outputs(4455) <= a or b;
    layer2_outputs(4456) <= a;
    layer2_outputs(4457) <= a and not b;
    layer2_outputs(4458) <= a or b;
    layer2_outputs(4459) <= not a or b;
    layer2_outputs(4460) <= not (a and b);
    layer2_outputs(4461) <= b;
    layer2_outputs(4462) <= '1';
    layer2_outputs(4463) <= b and not a;
    layer2_outputs(4464) <= not b;
    layer2_outputs(4465) <= not b;
    layer2_outputs(4466) <= a;
    layer2_outputs(4467) <= not a;
    layer2_outputs(4468) <= not a;
    layer2_outputs(4469) <= a and not b;
    layer2_outputs(4470) <= not b;
    layer2_outputs(4471) <= a or b;
    layer2_outputs(4472) <= a and not b;
    layer2_outputs(4473) <= b and not a;
    layer2_outputs(4474) <= '0';
    layer2_outputs(4475) <= not (a or b);
    layer2_outputs(4476) <= a or b;
    layer2_outputs(4477) <= not (a and b);
    layer2_outputs(4478) <= a;
    layer2_outputs(4479) <= b;
    layer2_outputs(4480) <= '0';
    layer2_outputs(4481) <= not (a and b);
    layer2_outputs(4482) <= not b or a;
    layer2_outputs(4483) <= not (a or b);
    layer2_outputs(4484) <= b and not a;
    layer2_outputs(4485) <= not b;
    layer2_outputs(4486) <= b and not a;
    layer2_outputs(4487) <= not b or a;
    layer2_outputs(4488) <= b and not a;
    layer2_outputs(4489) <= '1';
    layer2_outputs(4490) <= a and b;
    layer2_outputs(4491) <= not a;
    layer2_outputs(4492) <= '1';
    layer2_outputs(4493) <= '0';
    layer2_outputs(4494) <= '0';
    layer2_outputs(4495) <= not (a and b);
    layer2_outputs(4496) <= a or b;
    layer2_outputs(4497) <= not a or b;
    layer2_outputs(4498) <= not (a or b);
    layer2_outputs(4499) <= a xor b;
    layer2_outputs(4500) <= a;
    layer2_outputs(4501) <= a;
    layer2_outputs(4502) <= not a;
    layer2_outputs(4503) <= a and b;
    layer2_outputs(4504) <= not a or b;
    layer2_outputs(4505) <= b and not a;
    layer2_outputs(4506) <= not (a and b);
    layer2_outputs(4507) <= '1';
    layer2_outputs(4508) <= a;
    layer2_outputs(4509) <= a and not b;
    layer2_outputs(4510) <= a xor b;
    layer2_outputs(4511) <= '1';
    layer2_outputs(4512) <= '1';
    layer2_outputs(4513) <= not a or b;
    layer2_outputs(4514) <= not b or a;
    layer2_outputs(4515) <= not (a and b);
    layer2_outputs(4516) <= not (a or b);
    layer2_outputs(4517) <= a;
    layer2_outputs(4518) <= not a or b;
    layer2_outputs(4519) <= not (a or b);
    layer2_outputs(4520) <= not (a and b);
    layer2_outputs(4521) <= not (a or b);
    layer2_outputs(4522) <= a;
    layer2_outputs(4523) <= a and b;
    layer2_outputs(4524) <= not (a or b);
    layer2_outputs(4525) <= not a or b;
    layer2_outputs(4526) <= not b;
    layer2_outputs(4527) <= not (a and b);
    layer2_outputs(4528) <= not (a xor b);
    layer2_outputs(4529) <= not (a or b);
    layer2_outputs(4530) <= not b;
    layer2_outputs(4531) <= not a;
    layer2_outputs(4532) <= '1';
    layer2_outputs(4533) <= not (a or b);
    layer2_outputs(4534) <= '0';
    layer2_outputs(4535) <= b;
    layer2_outputs(4536) <= a;
    layer2_outputs(4537) <= a or b;
    layer2_outputs(4538) <= a xor b;
    layer2_outputs(4539) <= '0';
    layer2_outputs(4540) <= not (a or b);
    layer2_outputs(4541) <= a;
    layer2_outputs(4542) <= not b or a;
    layer2_outputs(4543) <= not a or b;
    layer2_outputs(4544) <= not b or a;
    layer2_outputs(4545) <= '1';
    layer2_outputs(4546) <= a and b;
    layer2_outputs(4547) <= b;
    layer2_outputs(4548) <= not a;
    layer2_outputs(4549) <= not a or b;
    layer2_outputs(4550) <= '0';
    layer2_outputs(4551) <= not a or b;
    layer2_outputs(4552) <= not a or b;
    layer2_outputs(4553) <= a and not b;
    layer2_outputs(4554) <= not a or b;
    layer2_outputs(4555) <= not a;
    layer2_outputs(4556) <= a or b;
    layer2_outputs(4557) <= not b or a;
    layer2_outputs(4558) <= not a or b;
    layer2_outputs(4559) <= not a;
    layer2_outputs(4560) <= '1';
    layer2_outputs(4561) <= a or b;
    layer2_outputs(4562) <= not (a xor b);
    layer2_outputs(4563) <= not (a and b);
    layer2_outputs(4564) <= not b;
    layer2_outputs(4565) <= not b or a;
    layer2_outputs(4566) <= a;
    layer2_outputs(4567) <= not (a and b);
    layer2_outputs(4568) <= a or b;
    layer2_outputs(4569) <= a;
    layer2_outputs(4570) <= a and not b;
    layer2_outputs(4571) <= not (a xor b);
    layer2_outputs(4572) <= '1';
    layer2_outputs(4573) <= not b;
    layer2_outputs(4574) <= '0';
    layer2_outputs(4575) <= not (a or b);
    layer2_outputs(4576) <= '1';
    layer2_outputs(4577) <= b;
    layer2_outputs(4578) <= not a or b;
    layer2_outputs(4579) <= '1';
    layer2_outputs(4580) <= not a or b;
    layer2_outputs(4581) <= a or b;
    layer2_outputs(4582) <= '1';
    layer2_outputs(4583) <= b;
    layer2_outputs(4584) <= a;
    layer2_outputs(4585) <= not a or b;
    layer2_outputs(4586) <= not (a and b);
    layer2_outputs(4587) <= b;
    layer2_outputs(4588) <= a or b;
    layer2_outputs(4589) <= b and not a;
    layer2_outputs(4590) <= b;
    layer2_outputs(4591) <= '0';
    layer2_outputs(4592) <= not b or a;
    layer2_outputs(4593) <= a or b;
    layer2_outputs(4594) <= '0';
    layer2_outputs(4595) <= not b or a;
    layer2_outputs(4596) <= b and not a;
    layer2_outputs(4597) <= a and b;
    layer2_outputs(4598) <= not (a and b);
    layer2_outputs(4599) <= '0';
    layer2_outputs(4600) <= not (a or b);
    layer2_outputs(4601) <= not b or a;
    layer2_outputs(4602) <= not b or a;
    layer2_outputs(4603) <= '1';
    layer2_outputs(4604) <= '0';
    layer2_outputs(4605) <= a xor b;
    layer2_outputs(4606) <= '1';
    layer2_outputs(4607) <= a and b;
    layer2_outputs(4608) <= not a or b;
    layer2_outputs(4609) <= not a;
    layer2_outputs(4610) <= '1';
    layer2_outputs(4611) <= a or b;
    layer2_outputs(4612) <= '0';
    layer2_outputs(4613) <= not (a xor b);
    layer2_outputs(4614) <= a and not b;
    layer2_outputs(4615) <= a and not b;
    layer2_outputs(4616) <= '0';
    layer2_outputs(4617) <= '0';
    layer2_outputs(4618) <= not b or a;
    layer2_outputs(4619) <= not (a or b);
    layer2_outputs(4620) <= b and not a;
    layer2_outputs(4621) <= '1';
    layer2_outputs(4622) <= not a or b;
    layer2_outputs(4623) <= not (a or b);
    layer2_outputs(4624) <= '1';
    layer2_outputs(4625) <= not (a and b);
    layer2_outputs(4626) <= a or b;
    layer2_outputs(4627) <= a xor b;
    layer2_outputs(4628) <= a or b;
    layer2_outputs(4629) <= not a;
    layer2_outputs(4630) <= '0';
    layer2_outputs(4631) <= not a or b;
    layer2_outputs(4632) <= b;
    layer2_outputs(4633) <= not a or b;
    layer2_outputs(4634) <= not a or b;
    layer2_outputs(4635) <= not a or b;
    layer2_outputs(4636) <= a;
    layer2_outputs(4637) <= a and b;
    layer2_outputs(4638) <= '1';
    layer2_outputs(4639) <= b;
    layer2_outputs(4640) <= a;
    layer2_outputs(4641) <= not (a and b);
    layer2_outputs(4642) <= b and not a;
    layer2_outputs(4643) <= not a;
    layer2_outputs(4644) <= '1';
    layer2_outputs(4645) <= a;
    layer2_outputs(4646) <= a or b;
    layer2_outputs(4647) <= not (a and b);
    layer2_outputs(4648) <= b and not a;
    layer2_outputs(4649) <= '1';
    layer2_outputs(4650) <= b and not a;
    layer2_outputs(4651) <= a xor b;
    layer2_outputs(4652) <= a and not b;
    layer2_outputs(4653) <= b and not a;
    layer2_outputs(4654) <= not (a or b);
    layer2_outputs(4655) <= b;
    layer2_outputs(4656) <= a and b;
    layer2_outputs(4657) <= not b;
    layer2_outputs(4658) <= b and not a;
    layer2_outputs(4659) <= not a;
    layer2_outputs(4660) <= b;
    layer2_outputs(4661) <= '1';
    layer2_outputs(4662) <= '1';
    layer2_outputs(4663) <= not b or a;
    layer2_outputs(4664) <= a xor b;
    layer2_outputs(4665) <= not (a or b);
    layer2_outputs(4666) <= a or b;
    layer2_outputs(4667) <= '1';
    layer2_outputs(4668) <= not a;
    layer2_outputs(4669) <= b;
    layer2_outputs(4670) <= not a;
    layer2_outputs(4671) <= b;
    layer2_outputs(4672) <= not (a or b);
    layer2_outputs(4673) <= not (a or b);
    layer2_outputs(4674) <= not (a and b);
    layer2_outputs(4675) <= '0';
    layer2_outputs(4676) <= a and b;
    layer2_outputs(4677) <= not b or a;
    layer2_outputs(4678) <= not (a and b);
    layer2_outputs(4679) <= '1';
    layer2_outputs(4680) <= '1';
    layer2_outputs(4681) <= not a or b;
    layer2_outputs(4682) <= '0';
    layer2_outputs(4683) <= b and not a;
    layer2_outputs(4684) <= b and not a;
    layer2_outputs(4685) <= not a or b;
    layer2_outputs(4686) <= not b;
    layer2_outputs(4687) <= '1';
    layer2_outputs(4688) <= not b;
    layer2_outputs(4689) <= b;
    layer2_outputs(4690) <= a and not b;
    layer2_outputs(4691) <= not a or b;
    layer2_outputs(4692) <= not a or b;
    layer2_outputs(4693) <= not (a and b);
    layer2_outputs(4694) <= '1';
    layer2_outputs(4695) <= a and b;
    layer2_outputs(4696) <= not (a and b);
    layer2_outputs(4697) <= not b;
    layer2_outputs(4698) <= b and not a;
    layer2_outputs(4699) <= not a or b;
    layer2_outputs(4700) <= not b or a;
    layer2_outputs(4701) <= not b or a;
    layer2_outputs(4702) <= a and b;
    layer2_outputs(4703) <= a;
    layer2_outputs(4704) <= not b;
    layer2_outputs(4705) <= not (a or b);
    layer2_outputs(4706) <= not (a or b);
    layer2_outputs(4707) <= '0';
    layer2_outputs(4708) <= b and not a;
    layer2_outputs(4709) <= '0';
    layer2_outputs(4710) <= not a;
    layer2_outputs(4711) <= a or b;
    layer2_outputs(4712) <= not (a or b);
    layer2_outputs(4713) <= a and b;
    layer2_outputs(4714) <= a or b;
    layer2_outputs(4715) <= not (a xor b);
    layer2_outputs(4716) <= not a or b;
    layer2_outputs(4717) <= b and not a;
    layer2_outputs(4718) <= a or b;
    layer2_outputs(4719) <= not b or a;
    layer2_outputs(4720) <= not b or a;
    layer2_outputs(4721) <= a and b;
    layer2_outputs(4722) <= not a or b;
    layer2_outputs(4723) <= b and not a;
    layer2_outputs(4724) <= '0';
    layer2_outputs(4725) <= not a;
    layer2_outputs(4726) <= a;
    layer2_outputs(4727) <= not (a or b);
    layer2_outputs(4728) <= not a;
    layer2_outputs(4729) <= not (a and b);
    layer2_outputs(4730) <= a or b;
    layer2_outputs(4731) <= not (a xor b);
    layer2_outputs(4732) <= b;
    layer2_outputs(4733) <= not (a or b);
    layer2_outputs(4734) <= a;
    layer2_outputs(4735) <= a and not b;
    layer2_outputs(4736) <= a and b;
    layer2_outputs(4737) <= a;
    layer2_outputs(4738) <= '1';
    layer2_outputs(4739) <= not (a or b);
    layer2_outputs(4740) <= not b or a;
    layer2_outputs(4741) <= b and not a;
    layer2_outputs(4742) <= a and b;
    layer2_outputs(4743) <= '0';
    layer2_outputs(4744) <= b and not a;
    layer2_outputs(4745) <= '0';
    layer2_outputs(4746) <= not (a and b);
    layer2_outputs(4747) <= not a;
    layer2_outputs(4748) <= b and not a;
    layer2_outputs(4749) <= a and not b;
    layer2_outputs(4750) <= '1';
    layer2_outputs(4751) <= '1';
    layer2_outputs(4752) <= a;
    layer2_outputs(4753) <= a and b;
    layer2_outputs(4754) <= a and b;
    layer2_outputs(4755) <= b;
    layer2_outputs(4756) <= a and b;
    layer2_outputs(4757) <= a xor b;
    layer2_outputs(4758) <= not b or a;
    layer2_outputs(4759) <= not a or b;
    layer2_outputs(4760) <= '1';
    layer2_outputs(4761) <= not b;
    layer2_outputs(4762) <= not a;
    layer2_outputs(4763) <= not (a xor b);
    layer2_outputs(4764) <= b;
    layer2_outputs(4765) <= b and not a;
    layer2_outputs(4766) <= a;
    layer2_outputs(4767) <= a;
    layer2_outputs(4768) <= a or b;
    layer2_outputs(4769) <= not b;
    layer2_outputs(4770) <= b;
    layer2_outputs(4771) <= not (a and b);
    layer2_outputs(4772) <= a and b;
    layer2_outputs(4773) <= not (a or b);
    layer2_outputs(4774) <= not b or a;
    layer2_outputs(4775) <= '1';
    layer2_outputs(4776) <= not b or a;
    layer2_outputs(4777) <= not a or b;
    layer2_outputs(4778) <= a;
    layer2_outputs(4779) <= not a or b;
    layer2_outputs(4780) <= '0';
    layer2_outputs(4781) <= '1';
    layer2_outputs(4782) <= not (a and b);
    layer2_outputs(4783) <= '0';
    layer2_outputs(4784) <= a and not b;
    layer2_outputs(4785) <= b;
    layer2_outputs(4786) <= a xor b;
    layer2_outputs(4787) <= b;
    layer2_outputs(4788) <= b;
    layer2_outputs(4789) <= not b or a;
    layer2_outputs(4790) <= a or b;
    layer2_outputs(4791) <= '0';
    layer2_outputs(4792) <= not (a or b);
    layer2_outputs(4793) <= a or b;
    layer2_outputs(4794) <= b;
    layer2_outputs(4795) <= not (a xor b);
    layer2_outputs(4796) <= b;
    layer2_outputs(4797) <= a or b;
    layer2_outputs(4798) <= not a or b;
    layer2_outputs(4799) <= a and b;
    layer2_outputs(4800) <= b and not a;
    layer2_outputs(4801) <= a and b;
    layer2_outputs(4802) <= a or b;
    layer2_outputs(4803) <= not a;
    layer2_outputs(4804) <= a;
    layer2_outputs(4805) <= not (a and b);
    layer2_outputs(4806) <= not (a or b);
    layer2_outputs(4807) <= not b or a;
    layer2_outputs(4808) <= '0';
    layer2_outputs(4809) <= a and b;
    layer2_outputs(4810) <= a and b;
    layer2_outputs(4811) <= not a;
    layer2_outputs(4812) <= a and not b;
    layer2_outputs(4813) <= b and not a;
    layer2_outputs(4814) <= not (a and b);
    layer2_outputs(4815) <= not a or b;
    layer2_outputs(4816) <= not b or a;
    layer2_outputs(4817) <= b and not a;
    layer2_outputs(4818) <= not (a or b);
    layer2_outputs(4819) <= not (a xor b);
    layer2_outputs(4820) <= a xor b;
    layer2_outputs(4821) <= b;
    layer2_outputs(4822) <= b and not a;
    layer2_outputs(4823) <= a and not b;
    layer2_outputs(4824) <= not (a xor b);
    layer2_outputs(4825) <= not (a or b);
    layer2_outputs(4826) <= not (a and b);
    layer2_outputs(4827) <= not (a and b);
    layer2_outputs(4828) <= not b or a;
    layer2_outputs(4829) <= b and not a;
    layer2_outputs(4830) <= a or b;
    layer2_outputs(4831) <= a and not b;
    layer2_outputs(4832) <= '1';
    layer2_outputs(4833) <= '1';
    layer2_outputs(4834) <= not (a and b);
    layer2_outputs(4835) <= b;
    layer2_outputs(4836) <= a xor b;
    layer2_outputs(4837) <= a or b;
    layer2_outputs(4838) <= not (a xor b);
    layer2_outputs(4839) <= not (a or b);
    layer2_outputs(4840) <= a and not b;
    layer2_outputs(4841) <= not a;
    layer2_outputs(4842) <= b and not a;
    layer2_outputs(4843) <= '1';
    layer2_outputs(4844) <= not a;
    layer2_outputs(4845) <= not (a or b);
    layer2_outputs(4846) <= not (a and b);
    layer2_outputs(4847) <= a;
    layer2_outputs(4848) <= a and not b;
    layer2_outputs(4849) <= not a;
    layer2_outputs(4850) <= not b;
    layer2_outputs(4851) <= a and not b;
    layer2_outputs(4852) <= b;
    layer2_outputs(4853) <= not (a or b);
    layer2_outputs(4854) <= '1';
    layer2_outputs(4855) <= not a or b;
    layer2_outputs(4856) <= a and not b;
    layer2_outputs(4857) <= not b or a;
    layer2_outputs(4858) <= not (a and b);
    layer2_outputs(4859) <= not a;
    layer2_outputs(4860) <= a and b;
    layer2_outputs(4861) <= '1';
    layer2_outputs(4862) <= '0';
    layer2_outputs(4863) <= not (a or b);
    layer2_outputs(4864) <= b and not a;
    layer2_outputs(4865) <= '1';
    layer2_outputs(4866) <= not b;
    layer2_outputs(4867) <= not a or b;
    layer2_outputs(4868) <= not a or b;
    layer2_outputs(4869) <= a and not b;
    layer2_outputs(4870) <= not a or b;
    layer2_outputs(4871) <= not (a or b);
    layer2_outputs(4872) <= a and b;
    layer2_outputs(4873) <= a or b;
    layer2_outputs(4874) <= not a;
    layer2_outputs(4875) <= a and not b;
    layer2_outputs(4876) <= a;
    layer2_outputs(4877) <= not a or b;
    layer2_outputs(4878) <= not a or b;
    layer2_outputs(4879) <= not (a and b);
    layer2_outputs(4880) <= not (a or b);
    layer2_outputs(4881) <= '1';
    layer2_outputs(4882) <= a or b;
    layer2_outputs(4883) <= a;
    layer2_outputs(4884) <= '0';
    layer2_outputs(4885) <= '1';
    layer2_outputs(4886) <= a and not b;
    layer2_outputs(4887) <= b;
    layer2_outputs(4888) <= a and b;
    layer2_outputs(4889) <= not (a xor b);
    layer2_outputs(4890) <= b and not a;
    layer2_outputs(4891) <= a;
    layer2_outputs(4892) <= a and not b;
    layer2_outputs(4893) <= not b or a;
    layer2_outputs(4894) <= not b or a;
    layer2_outputs(4895) <= not a;
    layer2_outputs(4896) <= not (a or b);
    layer2_outputs(4897) <= not a;
    layer2_outputs(4898) <= a;
    layer2_outputs(4899) <= not b;
    layer2_outputs(4900) <= '1';
    layer2_outputs(4901) <= not b;
    layer2_outputs(4902) <= a or b;
    layer2_outputs(4903) <= a or b;
    layer2_outputs(4904) <= not (a and b);
    layer2_outputs(4905) <= not a or b;
    layer2_outputs(4906) <= not (a xor b);
    layer2_outputs(4907) <= a or b;
    layer2_outputs(4908) <= '0';
    layer2_outputs(4909) <= '0';
    layer2_outputs(4910) <= a and b;
    layer2_outputs(4911) <= a or b;
    layer2_outputs(4912) <= b;
    layer2_outputs(4913) <= not a or b;
    layer2_outputs(4914) <= not (a or b);
    layer2_outputs(4915) <= b;
    layer2_outputs(4916) <= b and not a;
    layer2_outputs(4917) <= '0';
    layer2_outputs(4918) <= b;
    layer2_outputs(4919) <= a or b;
    layer2_outputs(4920) <= not b or a;
    layer2_outputs(4921) <= not b;
    layer2_outputs(4922) <= b and not a;
    layer2_outputs(4923) <= not (a and b);
    layer2_outputs(4924) <= not a or b;
    layer2_outputs(4925) <= b;
    layer2_outputs(4926) <= '1';
    layer2_outputs(4927) <= not b or a;
    layer2_outputs(4928) <= not b;
    layer2_outputs(4929) <= not (a and b);
    layer2_outputs(4930) <= not b or a;
    layer2_outputs(4931) <= not (a and b);
    layer2_outputs(4932) <= '1';
    layer2_outputs(4933) <= not b;
    layer2_outputs(4934) <= '0';
    layer2_outputs(4935) <= not a or b;
    layer2_outputs(4936) <= a and not b;
    layer2_outputs(4937) <= not a;
    layer2_outputs(4938) <= not a;
    layer2_outputs(4939) <= not (a and b);
    layer2_outputs(4940) <= not b;
    layer2_outputs(4941) <= not b or a;
    layer2_outputs(4942) <= a and not b;
    layer2_outputs(4943) <= not a;
    layer2_outputs(4944) <= not b;
    layer2_outputs(4945) <= not (a or b);
    layer2_outputs(4946) <= a and b;
    layer2_outputs(4947) <= not a or b;
    layer2_outputs(4948) <= a or b;
    layer2_outputs(4949) <= not b or a;
    layer2_outputs(4950) <= '0';
    layer2_outputs(4951) <= not b or a;
    layer2_outputs(4952) <= not (a and b);
    layer2_outputs(4953) <= a;
    layer2_outputs(4954) <= not b;
    layer2_outputs(4955) <= a and not b;
    layer2_outputs(4956) <= not (a xor b);
    layer2_outputs(4957) <= a and b;
    layer2_outputs(4958) <= a;
    layer2_outputs(4959) <= not b or a;
    layer2_outputs(4960) <= b and not a;
    layer2_outputs(4961) <= not (a and b);
    layer2_outputs(4962) <= '0';
    layer2_outputs(4963) <= a;
    layer2_outputs(4964) <= a and b;
    layer2_outputs(4965) <= a and not b;
    layer2_outputs(4966) <= b and not a;
    layer2_outputs(4967) <= '0';
    layer2_outputs(4968) <= a and not b;
    layer2_outputs(4969) <= not a or b;
    layer2_outputs(4970) <= not b;
    layer2_outputs(4971) <= not a;
    layer2_outputs(4972) <= b and not a;
    layer2_outputs(4973) <= not (a or b);
    layer2_outputs(4974) <= not b;
    layer2_outputs(4975) <= not b;
    layer2_outputs(4976) <= b and not a;
    layer2_outputs(4977) <= a;
    layer2_outputs(4978) <= not b;
    layer2_outputs(4979) <= not (a xor b);
    layer2_outputs(4980) <= not b or a;
    layer2_outputs(4981) <= '0';
    layer2_outputs(4982) <= a and not b;
    layer2_outputs(4983) <= not (a and b);
    layer2_outputs(4984) <= '0';
    layer2_outputs(4985) <= '1';
    layer2_outputs(4986) <= not a or b;
    layer2_outputs(4987) <= '0';
    layer2_outputs(4988) <= '0';
    layer2_outputs(4989) <= not a or b;
    layer2_outputs(4990) <= not (a and b);
    layer2_outputs(4991) <= a or b;
    layer2_outputs(4992) <= not b or a;
    layer2_outputs(4993) <= a and not b;
    layer2_outputs(4994) <= not b or a;
    layer2_outputs(4995) <= b and not a;
    layer2_outputs(4996) <= not (a or b);
    layer2_outputs(4997) <= a or b;
    layer2_outputs(4998) <= not b or a;
    layer2_outputs(4999) <= '0';
    layer2_outputs(5000) <= '1';
    layer2_outputs(5001) <= '1';
    layer2_outputs(5002) <= not (a or b);
    layer2_outputs(5003) <= '0';
    layer2_outputs(5004) <= b;
    layer2_outputs(5005) <= not a or b;
    layer2_outputs(5006) <= a or b;
    layer2_outputs(5007) <= a or b;
    layer2_outputs(5008) <= not b or a;
    layer2_outputs(5009) <= not a;
    layer2_outputs(5010) <= not (a or b);
    layer2_outputs(5011) <= b and not a;
    layer2_outputs(5012) <= a or b;
    layer2_outputs(5013) <= a and not b;
    layer2_outputs(5014) <= a or b;
    layer2_outputs(5015) <= '1';
    layer2_outputs(5016) <= b;
    layer2_outputs(5017) <= not a;
    layer2_outputs(5018) <= not a;
    layer2_outputs(5019) <= b and not a;
    layer2_outputs(5020) <= '0';
    layer2_outputs(5021) <= b and not a;
    layer2_outputs(5022) <= not (a xor b);
    layer2_outputs(5023) <= a and not b;
    layer2_outputs(5024) <= not b;
    layer2_outputs(5025) <= not (a or b);
    layer2_outputs(5026) <= not (a and b);
    layer2_outputs(5027) <= a and not b;
    layer2_outputs(5028) <= '0';
    layer2_outputs(5029) <= a and not b;
    layer2_outputs(5030) <= '0';
    layer2_outputs(5031) <= a and not b;
    layer2_outputs(5032) <= b and not a;
    layer2_outputs(5033) <= not b or a;
    layer2_outputs(5034) <= not b or a;
    layer2_outputs(5035) <= a and not b;
    layer2_outputs(5036) <= '1';
    layer2_outputs(5037) <= not b or a;
    layer2_outputs(5038) <= '1';
    layer2_outputs(5039) <= b and not a;
    layer2_outputs(5040) <= not b;
    layer2_outputs(5041) <= a and not b;
    layer2_outputs(5042) <= '0';
    layer2_outputs(5043) <= a and b;
    layer2_outputs(5044) <= a;
    layer2_outputs(5045) <= b;
    layer2_outputs(5046) <= a;
    layer2_outputs(5047) <= a and not b;
    layer2_outputs(5048) <= not a or b;
    layer2_outputs(5049) <= a or b;
    layer2_outputs(5050) <= b;
    layer2_outputs(5051) <= b and not a;
    layer2_outputs(5052) <= b;
    layer2_outputs(5053) <= '1';
    layer2_outputs(5054) <= a;
    layer2_outputs(5055) <= a;
    layer2_outputs(5056) <= not a or b;
    layer2_outputs(5057) <= '0';
    layer2_outputs(5058) <= not a;
    layer2_outputs(5059) <= not (a xor b);
    layer2_outputs(5060) <= a and not b;
    layer2_outputs(5061) <= a and b;
    layer2_outputs(5062) <= not b or a;
    layer2_outputs(5063) <= b;
    layer2_outputs(5064) <= not (a and b);
    layer2_outputs(5065) <= '0';
    layer2_outputs(5066) <= a;
    layer2_outputs(5067) <= a or b;
    layer2_outputs(5068) <= b and not a;
    layer2_outputs(5069) <= not a;
    layer2_outputs(5070) <= a xor b;
    layer2_outputs(5071) <= a or b;
    layer2_outputs(5072) <= a or b;
    layer2_outputs(5073) <= b and not a;
    layer2_outputs(5074) <= '0';
    layer2_outputs(5075) <= a xor b;
    layer2_outputs(5076) <= a or b;
    layer2_outputs(5077) <= not (a or b);
    layer2_outputs(5078) <= b;
    layer2_outputs(5079) <= not (a and b);
    layer2_outputs(5080) <= a or b;
    layer2_outputs(5081) <= not (a and b);
    layer2_outputs(5082) <= a and not b;
    layer2_outputs(5083) <= not b or a;
    layer2_outputs(5084) <= '0';
    layer2_outputs(5085) <= not (a xor b);
    layer2_outputs(5086) <= a or b;
    layer2_outputs(5087) <= a and b;
    layer2_outputs(5088) <= a or b;
    layer2_outputs(5089) <= a xor b;
    layer2_outputs(5090) <= a and not b;
    layer2_outputs(5091) <= a or b;
    layer2_outputs(5092) <= '0';
    layer2_outputs(5093) <= not (a xor b);
    layer2_outputs(5094) <= '1';
    layer2_outputs(5095) <= '0';
    layer2_outputs(5096) <= '1';
    layer2_outputs(5097) <= not b;
    layer2_outputs(5098) <= a or b;
    layer2_outputs(5099) <= a and not b;
    layer2_outputs(5100) <= '1';
    layer2_outputs(5101) <= a and not b;
    layer2_outputs(5102) <= a and b;
    layer2_outputs(5103) <= not (a and b);
    layer2_outputs(5104) <= a;
    layer2_outputs(5105) <= a;
    layer2_outputs(5106) <= '1';
    layer2_outputs(5107) <= a xor b;
    layer2_outputs(5108) <= a and b;
    layer2_outputs(5109) <= not b or a;
    layer2_outputs(5110) <= a;
    layer2_outputs(5111) <= a and b;
    layer2_outputs(5112) <= '1';
    layer2_outputs(5113) <= not a or b;
    layer2_outputs(5114) <= not (a or b);
    layer2_outputs(5115) <= '0';
    layer2_outputs(5116) <= b;
    layer2_outputs(5117) <= not a or b;
    layer2_outputs(5118) <= not (a and b);
    layer2_outputs(5119) <= a xor b;
    layer2_outputs(5120) <= a;
    layer2_outputs(5121) <= not (a and b);
    layer2_outputs(5122) <= a and b;
    layer2_outputs(5123) <= '0';
    layer2_outputs(5124) <= not (a and b);
    layer2_outputs(5125) <= not (a and b);
    layer2_outputs(5126) <= a and not b;
    layer2_outputs(5127) <= a and b;
    layer2_outputs(5128) <= not (a and b);
    layer2_outputs(5129) <= '1';
    layer2_outputs(5130) <= '0';
    layer2_outputs(5131) <= '0';
    layer2_outputs(5132) <= not (a or b);
    layer2_outputs(5133) <= not (a or b);
    layer2_outputs(5134) <= '1';
    layer2_outputs(5135) <= '0';
    layer2_outputs(5136) <= not b;
    layer2_outputs(5137) <= '0';
    layer2_outputs(5138) <= a;
    layer2_outputs(5139) <= a;
    layer2_outputs(5140) <= b;
    layer2_outputs(5141) <= a and b;
    layer2_outputs(5142) <= b;
    layer2_outputs(5143) <= '1';
    layer2_outputs(5144) <= a and not b;
    layer2_outputs(5145) <= not (a or b);
    layer2_outputs(5146) <= not b;
    layer2_outputs(5147) <= '1';
    layer2_outputs(5148) <= a;
    layer2_outputs(5149) <= '0';
    layer2_outputs(5150) <= a and not b;
    layer2_outputs(5151) <= b;
    layer2_outputs(5152) <= not a;
    layer2_outputs(5153) <= not (a and b);
    layer2_outputs(5154) <= not a or b;
    layer2_outputs(5155) <= not b;
    layer2_outputs(5156) <= '0';
    layer2_outputs(5157) <= not (a or b);
    layer2_outputs(5158) <= not a;
    layer2_outputs(5159) <= b;
    layer2_outputs(5160) <= not b or a;
    layer2_outputs(5161) <= not (a and b);
    layer2_outputs(5162) <= not a or b;
    layer2_outputs(5163) <= not b or a;
    layer2_outputs(5164) <= b and not a;
    layer2_outputs(5165) <= '1';
    layer2_outputs(5166) <= not (a and b);
    layer2_outputs(5167) <= a and not b;
    layer2_outputs(5168) <= not b;
    layer2_outputs(5169) <= not b;
    layer2_outputs(5170) <= a or b;
    layer2_outputs(5171) <= a and not b;
    layer2_outputs(5172) <= b;
    layer2_outputs(5173) <= b and not a;
    layer2_outputs(5174) <= not a;
    layer2_outputs(5175) <= a xor b;
    layer2_outputs(5176) <= b;
    layer2_outputs(5177) <= a or b;
    layer2_outputs(5178) <= b and not a;
    layer2_outputs(5179) <= not (a and b);
    layer2_outputs(5180) <= a and not b;
    layer2_outputs(5181) <= not (a and b);
    layer2_outputs(5182) <= not b or a;
    layer2_outputs(5183) <= not b;
    layer2_outputs(5184) <= '1';
    layer2_outputs(5185) <= a and not b;
    layer2_outputs(5186) <= a and b;
    layer2_outputs(5187) <= a and b;
    layer2_outputs(5188) <= a and not b;
    layer2_outputs(5189) <= a or b;
    layer2_outputs(5190) <= not a;
    layer2_outputs(5191) <= a and not b;
    layer2_outputs(5192) <= '0';
    layer2_outputs(5193) <= '0';
    layer2_outputs(5194) <= not b;
    layer2_outputs(5195) <= not b or a;
    layer2_outputs(5196) <= '1';
    layer2_outputs(5197) <= not (a xor b);
    layer2_outputs(5198) <= b and not a;
    layer2_outputs(5199) <= not (a xor b);
    layer2_outputs(5200) <= not (a and b);
    layer2_outputs(5201) <= a and not b;
    layer2_outputs(5202) <= a or b;
    layer2_outputs(5203) <= not (a and b);
    layer2_outputs(5204) <= b;
    layer2_outputs(5205) <= not a or b;
    layer2_outputs(5206) <= a;
    layer2_outputs(5207) <= b and not a;
    layer2_outputs(5208) <= not a or b;
    layer2_outputs(5209) <= not (a or b);
    layer2_outputs(5210) <= not a;
    layer2_outputs(5211) <= not b;
    layer2_outputs(5212) <= '0';
    layer2_outputs(5213) <= not (a or b);
    layer2_outputs(5214) <= b and not a;
    layer2_outputs(5215) <= a and b;
    layer2_outputs(5216) <= not (a and b);
    layer2_outputs(5217) <= not a;
    layer2_outputs(5218) <= '0';
    layer2_outputs(5219) <= b and not a;
    layer2_outputs(5220) <= not (a and b);
    layer2_outputs(5221) <= a and b;
    layer2_outputs(5222) <= '0';
    layer2_outputs(5223) <= '1';
    layer2_outputs(5224) <= b;
    layer2_outputs(5225) <= not a or b;
    layer2_outputs(5226) <= not b;
    layer2_outputs(5227) <= a;
    layer2_outputs(5228) <= '1';
    layer2_outputs(5229) <= a and not b;
    layer2_outputs(5230) <= a;
    layer2_outputs(5231) <= not a or b;
    layer2_outputs(5232) <= a;
    layer2_outputs(5233) <= b;
    layer2_outputs(5234) <= '0';
    layer2_outputs(5235) <= not b;
    layer2_outputs(5236) <= not a;
    layer2_outputs(5237) <= '0';
    layer2_outputs(5238) <= a;
    layer2_outputs(5239) <= not a or b;
    layer2_outputs(5240) <= b and not a;
    layer2_outputs(5241) <= a;
    layer2_outputs(5242) <= not (a and b);
    layer2_outputs(5243) <= '0';
    layer2_outputs(5244) <= not (a and b);
    layer2_outputs(5245) <= not (a or b);
    layer2_outputs(5246) <= not b or a;
    layer2_outputs(5247) <= a;
    layer2_outputs(5248) <= not a;
    layer2_outputs(5249) <= not b or a;
    layer2_outputs(5250) <= not a;
    layer2_outputs(5251) <= '0';
    layer2_outputs(5252) <= not (a and b);
    layer2_outputs(5253) <= '1';
    layer2_outputs(5254) <= a and not b;
    layer2_outputs(5255) <= a or b;
    layer2_outputs(5256) <= not a;
    layer2_outputs(5257) <= a xor b;
    layer2_outputs(5258) <= not (a xor b);
    layer2_outputs(5259) <= b;
    layer2_outputs(5260) <= not a or b;
    layer2_outputs(5261) <= a or b;
    layer2_outputs(5262) <= a and b;
    layer2_outputs(5263) <= '1';
    layer2_outputs(5264) <= b;
    layer2_outputs(5265) <= '0';
    layer2_outputs(5266) <= not b or a;
    layer2_outputs(5267) <= a and not b;
    layer2_outputs(5268) <= a;
    layer2_outputs(5269) <= '0';
    layer2_outputs(5270) <= not b;
    layer2_outputs(5271) <= a and b;
    layer2_outputs(5272) <= a and not b;
    layer2_outputs(5273) <= not (a and b);
    layer2_outputs(5274) <= a or b;
    layer2_outputs(5275) <= a and b;
    layer2_outputs(5276) <= b and not a;
    layer2_outputs(5277) <= a or b;
    layer2_outputs(5278) <= not (a or b);
    layer2_outputs(5279) <= a and b;
    layer2_outputs(5280) <= not b;
    layer2_outputs(5281) <= a and b;
    layer2_outputs(5282) <= not b;
    layer2_outputs(5283) <= '0';
    layer2_outputs(5284) <= '0';
    layer2_outputs(5285) <= '1';
    layer2_outputs(5286) <= '0';
    layer2_outputs(5287) <= not a;
    layer2_outputs(5288) <= not (a or b);
    layer2_outputs(5289) <= not b or a;
    layer2_outputs(5290) <= not (a and b);
    layer2_outputs(5291) <= not (a and b);
    layer2_outputs(5292) <= a and b;
    layer2_outputs(5293) <= a;
    layer2_outputs(5294) <= not a;
    layer2_outputs(5295) <= not b or a;
    layer2_outputs(5296) <= a and not b;
    layer2_outputs(5297) <= a and b;
    layer2_outputs(5298) <= '0';
    layer2_outputs(5299) <= not b or a;
    layer2_outputs(5300) <= a and not b;
    layer2_outputs(5301) <= not (a or b);
    layer2_outputs(5302) <= a;
    layer2_outputs(5303) <= '1';
    layer2_outputs(5304) <= not (a and b);
    layer2_outputs(5305) <= not b or a;
    layer2_outputs(5306) <= not a or b;
    layer2_outputs(5307) <= not a or b;
    layer2_outputs(5308) <= not b;
    layer2_outputs(5309) <= a and b;
    layer2_outputs(5310) <= not b or a;
    layer2_outputs(5311) <= a and not b;
    layer2_outputs(5312) <= a or b;
    layer2_outputs(5313) <= a or b;
    layer2_outputs(5314) <= not a or b;
    layer2_outputs(5315) <= not a;
    layer2_outputs(5316) <= not b or a;
    layer2_outputs(5317) <= a;
    layer2_outputs(5318) <= a and not b;
    layer2_outputs(5319) <= b and not a;
    layer2_outputs(5320) <= not a;
    layer2_outputs(5321) <= '0';
    layer2_outputs(5322) <= not a;
    layer2_outputs(5323) <= not b;
    layer2_outputs(5324) <= a and not b;
    layer2_outputs(5325) <= not a;
    layer2_outputs(5326) <= not b;
    layer2_outputs(5327) <= not a;
    layer2_outputs(5328) <= a and b;
    layer2_outputs(5329) <= '1';
    layer2_outputs(5330) <= not a;
    layer2_outputs(5331) <= not b or a;
    layer2_outputs(5332) <= a;
    layer2_outputs(5333) <= '0';
    layer2_outputs(5334) <= a;
    layer2_outputs(5335) <= b and not a;
    layer2_outputs(5336) <= b;
    layer2_outputs(5337) <= not a or b;
    layer2_outputs(5338) <= not (a and b);
    layer2_outputs(5339) <= a;
    layer2_outputs(5340) <= a and not b;
    layer2_outputs(5341) <= a and not b;
    layer2_outputs(5342) <= not (a and b);
    layer2_outputs(5343) <= not (a and b);
    layer2_outputs(5344) <= b;
    layer2_outputs(5345) <= a and not b;
    layer2_outputs(5346) <= not a or b;
    layer2_outputs(5347) <= not (a or b);
    layer2_outputs(5348) <= not b or a;
    layer2_outputs(5349) <= b and not a;
    layer2_outputs(5350) <= b and not a;
    layer2_outputs(5351) <= b and not a;
    layer2_outputs(5352) <= not b;
    layer2_outputs(5353) <= b;
    layer2_outputs(5354) <= '1';
    layer2_outputs(5355) <= b and not a;
    layer2_outputs(5356) <= b and not a;
    layer2_outputs(5357) <= b and not a;
    layer2_outputs(5358) <= not b or a;
    layer2_outputs(5359) <= not b or a;
    layer2_outputs(5360) <= '1';
    layer2_outputs(5361) <= '1';
    layer2_outputs(5362) <= not a;
    layer2_outputs(5363) <= b and not a;
    layer2_outputs(5364) <= a and not b;
    layer2_outputs(5365) <= '0';
    layer2_outputs(5366) <= a;
    layer2_outputs(5367) <= not b;
    layer2_outputs(5368) <= not a;
    layer2_outputs(5369) <= '1';
    layer2_outputs(5370) <= not b;
    layer2_outputs(5371) <= '0';
    layer2_outputs(5372) <= b and not a;
    layer2_outputs(5373) <= b;
    layer2_outputs(5374) <= not a or b;
    layer2_outputs(5375) <= b;
    layer2_outputs(5376) <= not b or a;
    layer2_outputs(5377) <= '1';
    layer2_outputs(5378) <= a and b;
    layer2_outputs(5379) <= not (a and b);
    layer2_outputs(5380) <= a and not b;
    layer2_outputs(5381) <= '0';
    layer2_outputs(5382) <= a xor b;
    layer2_outputs(5383) <= '1';
    layer2_outputs(5384) <= not a or b;
    layer2_outputs(5385) <= not a;
    layer2_outputs(5386) <= a and not b;
    layer2_outputs(5387) <= a xor b;
    layer2_outputs(5388) <= '0';
    layer2_outputs(5389) <= a;
    layer2_outputs(5390) <= '1';
    layer2_outputs(5391) <= a and b;
    layer2_outputs(5392) <= a and not b;
    layer2_outputs(5393) <= a or b;
    layer2_outputs(5394) <= b;
    layer2_outputs(5395) <= b and not a;
    layer2_outputs(5396) <= not a or b;
    layer2_outputs(5397) <= not a;
    layer2_outputs(5398) <= a or b;
    layer2_outputs(5399) <= '1';
    layer2_outputs(5400) <= '1';
    layer2_outputs(5401) <= not (a or b);
    layer2_outputs(5402) <= not (a or b);
    layer2_outputs(5403) <= not (a or b);
    layer2_outputs(5404) <= not (a and b);
    layer2_outputs(5405) <= not (a and b);
    layer2_outputs(5406) <= a and not b;
    layer2_outputs(5407) <= '0';
    layer2_outputs(5408) <= not a or b;
    layer2_outputs(5409) <= a xor b;
    layer2_outputs(5410) <= not (a or b);
    layer2_outputs(5411) <= '1';
    layer2_outputs(5412) <= '1';
    layer2_outputs(5413) <= a or b;
    layer2_outputs(5414) <= not b or a;
    layer2_outputs(5415) <= a;
    layer2_outputs(5416) <= a or b;
    layer2_outputs(5417) <= '0';
    layer2_outputs(5418) <= a and not b;
    layer2_outputs(5419) <= '1';
    layer2_outputs(5420) <= b and not a;
    layer2_outputs(5421) <= not (a or b);
    layer2_outputs(5422) <= a;
    layer2_outputs(5423) <= '1';
    layer2_outputs(5424) <= a;
    layer2_outputs(5425) <= b;
    layer2_outputs(5426) <= not (a or b);
    layer2_outputs(5427) <= a or b;
    layer2_outputs(5428) <= a and not b;
    layer2_outputs(5429) <= b;
    layer2_outputs(5430) <= a and b;
    layer2_outputs(5431) <= a;
    layer2_outputs(5432) <= '1';
    layer2_outputs(5433) <= not b or a;
    layer2_outputs(5434) <= b and not a;
    layer2_outputs(5435) <= b and not a;
    layer2_outputs(5436) <= not a or b;
    layer2_outputs(5437) <= not a or b;
    layer2_outputs(5438) <= not a or b;
    layer2_outputs(5439) <= a and b;
    layer2_outputs(5440) <= not a;
    layer2_outputs(5441) <= not a;
    layer2_outputs(5442) <= '0';
    layer2_outputs(5443) <= not a or b;
    layer2_outputs(5444) <= a;
    layer2_outputs(5445) <= b and not a;
    layer2_outputs(5446) <= '1';
    layer2_outputs(5447) <= '0';
    layer2_outputs(5448) <= a or b;
    layer2_outputs(5449) <= not (a and b);
    layer2_outputs(5450) <= not (a or b);
    layer2_outputs(5451) <= not a or b;
    layer2_outputs(5452) <= '0';
    layer2_outputs(5453) <= not b or a;
    layer2_outputs(5454) <= not a;
    layer2_outputs(5455) <= '1';
    layer2_outputs(5456) <= not a or b;
    layer2_outputs(5457) <= '0';
    layer2_outputs(5458) <= not (a and b);
    layer2_outputs(5459) <= a xor b;
    layer2_outputs(5460) <= a;
    layer2_outputs(5461) <= not b or a;
    layer2_outputs(5462) <= '1';
    layer2_outputs(5463) <= not b;
    layer2_outputs(5464) <= a and b;
    layer2_outputs(5465) <= '1';
    layer2_outputs(5466) <= not (a or b);
    layer2_outputs(5467) <= b and not a;
    layer2_outputs(5468) <= not a;
    layer2_outputs(5469) <= not (a and b);
    layer2_outputs(5470) <= b;
    layer2_outputs(5471) <= a;
    layer2_outputs(5472) <= not (a and b);
    layer2_outputs(5473) <= not a;
    layer2_outputs(5474) <= a or b;
    layer2_outputs(5475) <= not (a and b);
    layer2_outputs(5476) <= '0';
    layer2_outputs(5477) <= not (a xor b);
    layer2_outputs(5478) <= a;
    layer2_outputs(5479) <= a and not b;
    layer2_outputs(5480) <= not b or a;
    layer2_outputs(5481) <= not a or b;
    layer2_outputs(5482) <= a and not b;
    layer2_outputs(5483) <= b and not a;
    layer2_outputs(5484) <= not (a and b);
    layer2_outputs(5485) <= not (a and b);
    layer2_outputs(5486) <= not (a or b);
    layer2_outputs(5487) <= a and b;
    layer2_outputs(5488) <= not (a or b);
    layer2_outputs(5489) <= not b;
    layer2_outputs(5490) <= a and not b;
    layer2_outputs(5491) <= a or b;
    layer2_outputs(5492) <= '0';
    layer2_outputs(5493) <= a or b;
    layer2_outputs(5494) <= '1';
    layer2_outputs(5495) <= '1';
    layer2_outputs(5496) <= not a;
    layer2_outputs(5497) <= a or b;
    layer2_outputs(5498) <= '0';
    layer2_outputs(5499) <= '1';
    layer2_outputs(5500) <= '0';
    layer2_outputs(5501) <= '0';
    layer2_outputs(5502) <= a and b;
    layer2_outputs(5503) <= not b;
    layer2_outputs(5504) <= b;
    layer2_outputs(5505) <= not a;
    layer2_outputs(5506) <= b;
    layer2_outputs(5507) <= not (a or b);
    layer2_outputs(5508) <= a or b;
    layer2_outputs(5509) <= '0';
    layer2_outputs(5510) <= not b;
    layer2_outputs(5511) <= b and not a;
    layer2_outputs(5512) <= a and b;
    layer2_outputs(5513) <= '1';
    layer2_outputs(5514) <= not (a and b);
    layer2_outputs(5515) <= '0';
    layer2_outputs(5516) <= '0';
    layer2_outputs(5517) <= b;
    layer2_outputs(5518) <= b and not a;
    layer2_outputs(5519) <= not a or b;
    layer2_outputs(5520) <= not a or b;
    layer2_outputs(5521) <= a or b;
    layer2_outputs(5522) <= '0';
    layer2_outputs(5523) <= a xor b;
    layer2_outputs(5524) <= not b;
    layer2_outputs(5525) <= '1';
    layer2_outputs(5526) <= '0';
    layer2_outputs(5527) <= a and b;
    layer2_outputs(5528) <= a and not b;
    layer2_outputs(5529) <= a;
    layer2_outputs(5530) <= not (a and b);
    layer2_outputs(5531) <= '0';
    layer2_outputs(5532) <= not a;
    layer2_outputs(5533) <= b;
    layer2_outputs(5534) <= a xor b;
    layer2_outputs(5535) <= not (a and b);
    layer2_outputs(5536) <= not b or a;
    layer2_outputs(5537) <= not b;
    layer2_outputs(5538) <= '0';
    layer2_outputs(5539) <= not (a xor b);
    layer2_outputs(5540) <= not (a or b);
    layer2_outputs(5541) <= a;
    layer2_outputs(5542) <= not b;
    layer2_outputs(5543) <= '1';
    layer2_outputs(5544) <= not b or a;
    layer2_outputs(5545) <= b;
    layer2_outputs(5546) <= '0';
    layer2_outputs(5547) <= not (a and b);
    layer2_outputs(5548) <= '0';
    layer2_outputs(5549) <= a and not b;
    layer2_outputs(5550) <= not b;
    layer2_outputs(5551) <= b;
    layer2_outputs(5552) <= '1';
    layer2_outputs(5553) <= not (a and b);
    layer2_outputs(5554) <= '1';
    layer2_outputs(5555) <= '1';
    layer2_outputs(5556) <= not a;
    layer2_outputs(5557) <= not a or b;
    layer2_outputs(5558) <= not (a and b);
    layer2_outputs(5559) <= not a or b;
    layer2_outputs(5560) <= b and not a;
    layer2_outputs(5561) <= a and not b;
    layer2_outputs(5562) <= not (a and b);
    layer2_outputs(5563) <= not (a or b);
    layer2_outputs(5564) <= '0';
    layer2_outputs(5565) <= a and b;
    layer2_outputs(5566) <= not (a and b);
    layer2_outputs(5567) <= b;
    layer2_outputs(5568) <= '1';
    layer2_outputs(5569) <= a;
    layer2_outputs(5570) <= '0';
    layer2_outputs(5571) <= b;
    layer2_outputs(5572) <= not a or b;
    layer2_outputs(5573) <= not (a and b);
    layer2_outputs(5574) <= not a;
    layer2_outputs(5575) <= not b;
    layer2_outputs(5576) <= '0';
    layer2_outputs(5577) <= a or b;
    layer2_outputs(5578) <= a and b;
    layer2_outputs(5579) <= b;
    layer2_outputs(5580) <= not a;
    layer2_outputs(5581) <= a or b;
    layer2_outputs(5582) <= '0';
    layer2_outputs(5583) <= not b or a;
    layer2_outputs(5584) <= not a;
    layer2_outputs(5585) <= not (a and b);
    layer2_outputs(5586) <= not a or b;
    layer2_outputs(5587) <= a;
    layer2_outputs(5588) <= '1';
    layer2_outputs(5589) <= '1';
    layer2_outputs(5590) <= not a;
    layer2_outputs(5591) <= a and not b;
    layer2_outputs(5592) <= a xor b;
    layer2_outputs(5593) <= a and not b;
    layer2_outputs(5594) <= a or b;
    layer2_outputs(5595) <= not (a and b);
    layer2_outputs(5596) <= b;
    layer2_outputs(5597) <= '0';
    layer2_outputs(5598) <= b;
    layer2_outputs(5599) <= not a or b;
    layer2_outputs(5600) <= not b or a;
    layer2_outputs(5601) <= not a;
    layer2_outputs(5602) <= a or b;
    layer2_outputs(5603) <= not (a or b);
    layer2_outputs(5604) <= not (a and b);
    layer2_outputs(5605) <= a;
    layer2_outputs(5606) <= a or b;
    layer2_outputs(5607) <= not b or a;
    layer2_outputs(5608) <= a and not b;
    layer2_outputs(5609) <= a;
    layer2_outputs(5610) <= a or b;
    layer2_outputs(5611) <= '0';
    layer2_outputs(5612) <= b;
    layer2_outputs(5613) <= a and not b;
    layer2_outputs(5614) <= a and b;
    layer2_outputs(5615) <= a or b;
    layer2_outputs(5616) <= a and b;
    layer2_outputs(5617) <= not b;
    layer2_outputs(5618) <= b;
    layer2_outputs(5619) <= b and not a;
    layer2_outputs(5620) <= a and b;
    layer2_outputs(5621) <= '1';
    layer2_outputs(5622) <= not b or a;
    layer2_outputs(5623) <= not (a or b);
    layer2_outputs(5624) <= b and not a;
    layer2_outputs(5625) <= not (a or b);
    layer2_outputs(5626) <= a and not b;
    layer2_outputs(5627) <= a;
    layer2_outputs(5628) <= a xor b;
    layer2_outputs(5629) <= a xor b;
    layer2_outputs(5630) <= '0';
    layer2_outputs(5631) <= '1';
    layer2_outputs(5632) <= '0';
    layer2_outputs(5633) <= a and b;
    layer2_outputs(5634) <= not b;
    layer2_outputs(5635) <= a and not b;
    layer2_outputs(5636) <= a or b;
    layer2_outputs(5637) <= a;
    layer2_outputs(5638) <= b and not a;
    layer2_outputs(5639) <= b and not a;
    layer2_outputs(5640) <= a and not b;
    layer2_outputs(5641) <= a xor b;
    layer2_outputs(5642) <= '1';
    layer2_outputs(5643) <= a or b;
    layer2_outputs(5644) <= '0';
    layer2_outputs(5645) <= not b;
    layer2_outputs(5646) <= a and b;
    layer2_outputs(5647) <= b;
    layer2_outputs(5648) <= a and not b;
    layer2_outputs(5649) <= not b;
    layer2_outputs(5650) <= not (a and b);
    layer2_outputs(5651) <= not a;
    layer2_outputs(5652) <= '0';
    layer2_outputs(5653) <= '1';
    layer2_outputs(5654) <= a and not b;
    layer2_outputs(5655) <= not b;
    layer2_outputs(5656) <= b and not a;
    layer2_outputs(5657) <= not (a and b);
    layer2_outputs(5658) <= a or b;
    layer2_outputs(5659) <= '1';
    layer2_outputs(5660) <= a or b;
    layer2_outputs(5661) <= '1';
    layer2_outputs(5662) <= '0';
    layer2_outputs(5663) <= b and not a;
    layer2_outputs(5664) <= not b;
    layer2_outputs(5665) <= not b or a;
    layer2_outputs(5666) <= a or b;
    layer2_outputs(5667) <= not (a xor b);
    layer2_outputs(5668) <= '0';
    layer2_outputs(5669) <= a;
    layer2_outputs(5670) <= '0';
    layer2_outputs(5671) <= a and not b;
    layer2_outputs(5672) <= a and b;
    layer2_outputs(5673) <= '1';
    layer2_outputs(5674) <= b;
    layer2_outputs(5675) <= a;
    layer2_outputs(5676) <= not b or a;
    layer2_outputs(5677) <= not a or b;
    layer2_outputs(5678) <= not b;
    layer2_outputs(5679) <= b and not a;
    layer2_outputs(5680) <= a and not b;
    layer2_outputs(5681) <= a or b;
    layer2_outputs(5682) <= not (a or b);
    layer2_outputs(5683) <= not b;
    layer2_outputs(5684) <= not b or a;
    layer2_outputs(5685) <= a and not b;
    layer2_outputs(5686) <= '0';
    layer2_outputs(5687) <= not a;
    layer2_outputs(5688) <= a and not b;
    layer2_outputs(5689) <= not a or b;
    layer2_outputs(5690) <= b and not a;
    layer2_outputs(5691) <= a and b;
    layer2_outputs(5692) <= a and not b;
    layer2_outputs(5693) <= not (a or b);
    layer2_outputs(5694) <= not (a or b);
    layer2_outputs(5695) <= a and b;
    layer2_outputs(5696) <= not a or b;
    layer2_outputs(5697) <= a;
    layer2_outputs(5698) <= not (a or b);
    layer2_outputs(5699) <= a and b;
    layer2_outputs(5700) <= a and not b;
    layer2_outputs(5701) <= not a;
    layer2_outputs(5702) <= a and not b;
    layer2_outputs(5703) <= not (a or b);
    layer2_outputs(5704) <= '0';
    layer2_outputs(5705) <= not b or a;
    layer2_outputs(5706) <= '1';
    layer2_outputs(5707) <= a;
    layer2_outputs(5708) <= a xor b;
    layer2_outputs(5709) <= not (a and b);
    layer2_outputs(5710) <= not a or b;
    layer2_outputs(5711) <= not (a xor b);
    layer2_outputs(5712) <= not a or b;
    layer2_outputs(5713) <= b;
    layer2_outputs(5714) <= not (a and b);
    layer2_outputs(5715) <= a and not b;
    layer2_outputs(5716) <= b and not a;
    layer2_outputs(5717) <= a and not b;
    layer2_outputs(5718) <= '0';
    layer2_outputs(5719) <= not a;
    layer2_outputs(5720) <= a or b;
    layer2_outputs(5721) <= not (a or b);
    layer2_outputs(5722) <= b and not a;
    layer2_outputs(5723) <= b;
    layer2_outputs(5724) <= a;
    layer2_outputs(5725) <= a or b;
    layer2_outputs(5726) <= not a;
    layer2_outputs(5727) <= b and not a;
    layer2_outputs(5728) <= not (a or b);
    layer2_outputs(5729) <= not b;
    layer2_outputs(5730) <= b;
    layer2_outputs(5731) <= not b or a;
    layer2_outputs(5732) <= a and not b;
    layer2_outputs(5733) <= not a;
    layer2_outputs(5734) <= a or b;
    layer2_outputs(5735) <= '0';
    layer2_outputs(5736) <= b and not a;
    layer2_outputs(5737) <= '0';
    layer2_outputs(5738) <= not a;
    layer2_outputs(5739) <= a and b;
    layer2_outputs(5740) <= not (a or b);
    layer2_outputs(5741) <= '1';
    layer2_outputs(5742) <= not (a or b);
    layer2_outputs(5743) <= b and not a;
    layer2_outputs(5744) <= a and not b;
    layer2_outputs(5745) <= not a or b;
    layer2_outputs(5746) <= b and not a;
    layer2_outputs(5747) <= not b or a;
    layer2_outputs(5748) <= a;
    layer2_outputs(5749) <= a and not b;
    layer2_outputs(5750) <= '0';
    layer2_outputs(5751) <= not (a or b);
    layer2_outputs(5752) <= not b;
    layer2_outputs(5753) <= not (a and b);
    layer2_outputs(5754) <= a or b;
    layer2_outputs(5755) <= b and not a;
    layer2_outputs(5756) <= '0';
    layer2_outputs(5757) <= a and not b;
    layer2_outputs(5758) <= '1';
    layer2_outputs(5759) <= not a;
    layer2_outputs(5760) <= a or b;
    layer2_outputs(5761) <= not a or b;
    layer2_outputs(5762) <= '1';
    layer2_outputs(5763) <= '1';
    layer2_outputs(5764) <= '1';
    layer2_outputs(5765) <= a and not b;
    layer2_outputs(5766) <= '1';
    layer2_outputs(5767) <= b and not a;
    layer2_outputs(5768) <= '0';
    layer2_outputs(5769) <= '1';
    layer2_outputs(5770) <= a and not b;
    layer2_outputs(5771) <= '1';
    layer2_outputs(5772) <= '0';
    layer2_outputs(5773) <= not (a and b);
    layer2_outputs(5774) <= not (a or b);
    layer2_outputs(5775) <= not a;
    layer2_outputs(5776) <= not a or b;
    layer2_outputs(5777) <= not a or b;
    layer2_outputs(5778) <= not (a or b);
    layer2_outputs(5779) <= b;
    layer2_outputs(5780) <= not a;
    layer2_outputs(5781) <= not b or a;
    layer2_outputs(5782) <= a and b;
    layer2_outputs(5783) <= not b;
    layer2_outputs(5784) <= '0';
    layer2_outputs(5785) <= a xor b;
    layer2_outputs(5786) <= not b or a;
    layer2_outputs(5787) <= '0';
    layer2_outputs(5788) <= a and not b;
    layer2_outputs(5789) <= a;
    layer2_outputs(5790) <= not (a or b);
    layer2_outputs(5791) <= not b;
    layer2_outputs(5792) <= a and b;
    layer2_outputs(5793) <= a or b;
    layer2_outputs(5794) <= a or b;
    layer2_outputs(5795) <= not a;
    layer2_outputs(5796) <= b and not a;
    layer2_outputs(5797) <= not a or b;
    layer2_outputs(5798) <= not (a and b);
    layer2_outputs(5799) <= b;
    layer2_outputs(5800) <= '1';
    layer2_outputs(5801) <= '0';
    layer2_outputs(5802) <= not b or a;
    layer2_outputs(5803) <= not a;
    layer2_outputs(5804) <= not (a and b);
    layer2_outputs(5805) <= '0';
    layer2_outputs(5806) <= b;
    layer2_outputs(5807) <= not (a or b);
    layer2_outputs(5808) <= '1';
    layer2_outputs(5809) <= '0';
    layer2_outputs(5810) <= not b or a;
    layer2_outputs(5811) <= '1';
    layer2_outputs(5812) <= a or b;
    layer2_outputs(5813) <= a and not b;
    layer2_outputs(5814) <= '0';
    layer2_outputs(5815) <= not (a xor b);
    layer2_outputs(5816) <= not b;
    layer2_outputs(5817) <= a or b;
    layer2_outputs(5818) <= a;
    layer2_outputs(5819) <= not b;
    layer2_outputs(5820) <= not (a and b);
    layer2_outputs(5821) <= not a or b;
    layer2_outputs(5822) <= a xor b;
    layer2_outputs(5823) <= a or b;
    layer2_outputs(5824) <= a;
    layer2_outputs(5825) <= not a or b;
    layer2_outputs(5826) <= not (a and b);
    layer2_outputs(5827) <= not a or b;
    layer2_outputs(5828) <= b and not a;
    layer2_outputs(5829) <= not (a and b);
    layer2_outputs(5830) <= '0';
    layer2_outputs(5831) <= a or b;
    layer2_outputs(5832) <= a and not b;
    layer2_outputs(5833) <= not a or b;
    layer2_outputs(5834) <= not (a or b);
    layer2_outputs(5835) <= '0';
    layer2_outputs(5836) <= b and not a;
    layer2_outputs(5837) <= '1';
    layer2_outputs(5838) <= b;
    layer2_outputs(5839) <= b;
    layer2_outputs(5840) <= a and not b;
    layer2_outputs(5841) <= b;
    layer2_outputs(5842) <= not b or a;
    layer2_outputs(5843) <= '1';
    layer2_outputs(5844) <= a and not b;
    layer2_outputs(5845) <= not (a or b);
    layer2_outputs(5846) <= b;
    layer2_outputs(5847) <= not (a or b);
    layer2_outputs(5848) <= not (a and b);
    layer2_outputs(5849) <= a and not b;
    layer2_outputs(5850) <= not b or a;
    layer2_outputs(5851) <= '1';
    layer2_outputs(5852) <= '0';
    layer2_outputs(5853) <= b and not a;
    layer2_outputs(5854) <= '0';
    layer2_outputs(5855) <= a;
    layer2_outputs(5856) <= a;
    layer2_outputs(5857) <= a and b;
    layer2_outputs(5858) <= a and not b;
    layer2_outputs(5859) <= b;
    layer2_outputs(5860) <= a and not b;
    layer2_outputs(5861) <= b and not a;
    layer2_outputs(5862) <= a and b;
    layer2_outputs(5863) <= b and not a;
    layer2_outputs(5864) <= a;
    layer2_outputs(5865) <= '0';
    layer2_outputs(5866) <= '0';
    layer2_outputs(5867) <= a;
    layer2_outputs(5868) <= not (a or b);
    layer2_outputs(5869) <= not a or b;
    layer2_outputs(5870) <= '0';
    layer2_outputs(5871) <= not (a and b);
    layer2_outputs(5872) <= a or b;
    layer2_outputs(5873) <= not b or a;
    layer2_outputs(5874) <= not b or a;
    layer2_outputs(5875) <= not b;
    layer2_outputs(5876) <= a;
    layer2_outputs(5877) <= not a or b;
    layer2_outputs(5878) <= not (a and b);
    layer2_outputs(5879) <= '0';
    layer2_outputs(5880) <= a;
    layer2_outputs(5881) <= b;
    layer2_outputs(5882) <= not a;
    layer2_outputs(5883) <= a and not b;
    layer2_outputs(5884) <= not b;
    layer2_outputs(5885) <= not b;
    layer2_outputs(5886) <= a or b;
    layer2_outputs(5887) <= b;
    layer2_outputs(5888) <= not (a or b);
    layer2_outputs(5889) <= a;
    layer2_outputs(5890) <= a and b;
    layer2_outputs(5891) <= not b or a;
    layer2_outputs(5892) <= a and not b;
    layer2_outputs(5893) <= a and b;
    layer2_outputs(5894) <= '1';
    layer2_outputs(5895) <= b and not a;
    layer2_outputs(5896) <= not (a and b);
    layer2_outputs(5897) <= not a;
    layer2_outputs(5898) <= a;
    layer2_outputs(5899) <= a and not b;
    layer2_outputs(5900) <= b and not a;
    layer2_outputs(5901) <= a or b;
    layer2_outputs(5902) <= a and b;
    layer2_outputs(5903) <= not a or b;
    layer2_outputs(5904) <= '0';
    layer2_outputs(5905) <= not a or b;
    layer2_outputs(5906) <= a or b;
    layer2_outputs(5907) <= b and not a;
    layer2_outputs(5908) <= not b or a;
    layer2_outputs(5909) <= a;
    layer2_outputs(5910) <= '1';
    layer2_outputs(5911) <= a;
    layer2_outputs(5912) <= '0';
    layer2_outputs(5913) <= not b or a;
    layer2_outputs(5914) <= b and not a;
    layer2_outputs(5915) <= not a or b;
    layer2_outputs(5916) <= a;
    layer2_outputs(5917) <= not b;
    layer2_outputs(5918) <= not b;
    layer2_outputs(5919) <= not a;
    layer2_outputs(5920) <= '0';
    layer2_outputs(5921) <= '0';
    layer2_outputs(5922) <= a and b;
    layer2_outputs(5923) <= not b;
    layer2_outputs(5924) <= a and b;
    layer2_outputs(5925) <= not b;
    layer2_outputs(5926) <= '0';
    layer2_outputs(5927) <= '0';
    layer2_outputs(5928) <= b and not a;
    layer2_outputs(5929) <= not b or a;
    layer2_outputs(5930) <= b;
    layer2_outputs(5931) <= a;
    layer2_outputs(5932) <= not (a xor b);
    layer2_outputs(5933) <= '0';
    layer2_outputs(5934) <= a and b;
    layer2_outputs(5935) <= not a;
    layer2_outputs(5936) <= '0';
    layer2_outputs(5937) <= a and not b;
    layer2_outputs(5938) <= a and not b;
    layer2_outputs(5939) <= b;
    layer2_outputs(5940) <= not a or b;
    layer2_outputs(5941) <= a and not b;
    layer2_outputs(5942) <= '0';
    layer2_outputs(5943) <= b;
    layer2_outputs(5944) <= a and not b;
    layer2_outputs(5945) <= '0';
    layer2_outputs(5946) <= a and not b;
    layer2_outputs(5947) <= a;
    layer2_outputs(5948) <= '0';
    layer2_outputs(5949) <= b and not a;
    layer2_outputs(5950) <= not a or b;
    layer2_outputs(5951) <= a and b;
    layer2_outputs(5952) <= b and not a;
    layer2_outputs(5953) <= not a;
    layer2_outputs(5954) <= a;
    layer2_outputs(5955) <= '1';
    layer2_outputs(5956) <= b;
    layer2_outputs(5957) <= b;
    layer2_outputs(5958) <= a or b;
    layer2_outputs(5959) <= not b or a;
    layer2_outputs(5960) <= not a or b;
    layer2_outputs(5961) <= a;
    layer2_outputs(5962) <= not (a and b);
    layer2_outputs(5963) <= '1';
    layer2_outputs(5964) <= not (a and b);
    layer2_outputs(5965) <= a xor b;
    layer2_outputs(5966) <= not b;
    layer2_outputs(5967) <= not b;
    layer2_outputs(5968) <= not (a and b);
    layer2_outputs(5969) <= a and b;
    layer2_outputs(5970) <= '1';
    layer2_outputs(5971) <= not a;
    layer2_outputs(5972) <= not (a and b);
    layer2_outputs(5973) <= a and b;
    layer2_outputs(5974) <= '1';
    layer2_outputs(5975) <= not b or a;
    layer2_outputs(5976) <= a xor b;
    layer2_outputs(5977) <= a and b;
    layer2_outputs(5978) <= '1';
    layer2_outputs(5979) <= a;
    layer2_outputs(5980) <= b;
    layer2_outputs(5981) <= '1';
    layer2_outputs(5982) <= not (a or b);
    layer2_outputs(5983) <= a or b;
    layer2_outputs(5984) <= not (a or b);
    layer2_outputs(5985) <= not (a and b);
    layer2_outputs(5986) <= a or b;
    layer2_outputs(5987) <= '0';
    layer2_outputs(5988) <= '0';
    layer2_outputs(5989) <= not (a or b);
    layer2_outputs(5990) <= not a;
    layer2_outputs(5991) <= not a or b;
    layer2_outputs(5992) <= not (a and b);
    layer2_outputs(5993) <= a or b;
    layer2_outputs(5994) <= not a;
    layer2_outputs(5995) <= not b;
    layer2_outputs(5996) <= not (a xor b);
    layer2_outputs(5997) <= not (a and b);
    layer2_outputs(5998) <= a or b;
    layer2_outputs(5999) <= not (a and b);
    layer2_outputs(6000) <= not b or a;
    layer2_outputs(6001) <= '0';
    layer2_outputs(6002) <= not (a or b);
    layer2_outputs(6003) <= not (a xor b);
    layer2_outputs(6004) <= a xor b;
    layer2_outputs(6005) <= b;
    layer2_outputs(6006) <= not b;
    layer2_outputs(6007) <= b;
    layer2_outputs(6008) <= a and not b;
    layer2_outputs(6009) <= not a;
    layer2_outputs(6010) <= not (a and b);
    layer2_outputs(6011) <= not (a and b);
    layer2_outputs(6012) <= '1';
    layer2_outputs(6013) <= not a or b;
    layer2_outputs(6014) <= not b or a;
    layer2_outputs(6015) <= not (a and b);
    layer2_outputs(6016) <= b and not a;
    layer2_outputs(6017) <= '1';
    layer2_outputs(6018) <= a xor b;
    layer2_outputs(6019) <= a and not b;
    layer2_outputs(6020) <= '1';
    layer2_outputs(6021) <= b;
    layer2_outputs(6022) <= not (a and b);
    layer2_outputs(6023) <= b and not a;
    layer2_outputs(6024) <= b;
    layer2_outputs(6025) <= b and not a;
    layer2_outputs(6026) <= a and b;
    layer2_outputs(6027) <= not a;
    layer2_outputs(6028) <= a or b;
    layer2_outputs(6029) <= not b or a;
    layer2_outputs(6030) <= a or b;
    layer2_outputs(6031) <= a;
    layer2_outputs(6032) <= b and not a;
    layer2_outputs(6033) <= not a or b;
    layer2_outputs(6034) <= '0';
    layer2_outputs(6035) <= '1';
    layer2_outputs(6036) <= a and b;
    layer2_outputs(6037) <= a xor b;
    layer2_outputs(6038) <= not a or b;
    layer2_outputs(6039) <= not a;
    layer2_outputs(6040) <= not b;
    layer2_outputs(6041) <= a;
    layer2_outputs(6042) <= not b or a;
    layer2_outputs(6043) <= not b;
    layer2_outputs(6044) <= a or b;
    layer2_outputs(6045) <= not (a or b);
    layer2_outputs(6046) <= not a or b;
    layer2_outputs(6047) <= b and not a;
    layer2_outputs(6048) <= not (a or b);
    layer2_outputs(6049) <= b and not a;
    layer2_outputs(6050) <= b and not a;
    layer2_outputs(6051) <= a;
    layer2_outputs(6052) <= a and b;
    layer2_outputs(6053) <= not (a and b);
    layer2_outputs(6054) <= a and not b;
    layer2_outputs(6055) <= a and not b;
    layer2_outputs(6056) <= a;
    layer2_outputs(6057) <= not (a and b);
    layer2_outputs(6058) <= not b or a;
    layer2_outputs(6059) <= '1';
    layer2_outputs(6060) <= '1';
    layer2_outputs(6061) <= not a;
    layer2_outputs(6062) <= not b;
    layer2_outputs(6063) <= not a or b;
    layer2_outputs(6064) <= not a;
    layer2_outputs(6065) <= not (a or b);
    layer2_outputs(6066) <= not (a and b);
    layer2_outputs(6067) <= '1';
    layer2_outputs(6068) <= not a;
    layer2_outputs(6069) <= '1';
    layer2_outputs(6070) <= a and b;
    layer2_outputs(6071) <= a;
    layer2_outputs(6072) <= '0';
    layer2_outputs(6073) <= not a or b;
    layer2_outputs(6074) <= a or b;
    layer2_outputs(6075) <= b and not a;
    layer2_outputs(6076) <= not b;
    layer2_outputs(6077) <= a or b;
    layer2_outputs(6078) <= b and not a;
    layer2_outputs(6079) <= not (a and b);
    layer2_outputs(6080) <= not (a and b);
    layer2_outputs(6081) <= b;
    layer2_outputs(6082) <= '0';
    layer2_outputs(6083) <= not (a xor b);
    layer2_outputs(6084) <= a;
    layer2_outputs(6085) <= a and not b;
    layer2_outputs(6086) <= '1';
    layer2_outputs(6087) <= a and b;
    layer2_outputs(6088) <= a and b;
    layer2_outputs(6089) <= b and not a;
    layer2_outputs(6090) <= a and b;
    layer2_outputs(6091) <= not b or a;
    layer2_outputs(6092) <= '0';
    layer2_outputs(6093) <= a and not b;
    layer2_outputs(6094) <= a and b;
    layer2_outputs(6095) <= '1';
    layer2_outputs(6096) <= b and not a;
    layer2_outputs(6097) <= a;
    layer2_outputs(6098) <= not (a or b);
    layer2_outputs(6099) <= '0';
    layer2_outputs(6100) <= a and b;
    layer2_outputs(6101) <= not (a or b);
    layer2_outputs(6102) <= not (a and b);
    layer2_outputs(6103) <= '1';
    layer2_outputs(6104) <= not a;
    layer2_outputs(6105) <= not b;
    layer2_outputs(6106) <= not b;
    layer2_outputs(6107) <= not b;
    layer2_outputs(6108) <= a and not b;
    layer2_outputs(6109) <= a and not b;
    layer2_outputs(6110) <= '1';
    layer2_outputs(6111) <= a and b;
    layer2_outputs(6112) <= a;
    layer2_outputs(6113) <= a;
    layer2_outputs(6114) <= not a or b;
    layer2_outputs(6115) <= not (a and b);
    layer2_outputs(6116) <= not a or b;
    layer2_outputs(6117) <= b;
    layer2_outputs(6118) <= a and b;
    layer2_outputs(6119) <= '0';
    layer2_outputs(6120) <= not a;
    layer2_outputs(6121) <= not b or a;
    layer2_outputs(6122) <= not (a or b);
    layer2_outputs(6123) <= not (a and b);
    layer2_outputs(6124) <= a;
    layer2_outputs(6125) <= not b or a;
    layer2_outputs(6126) <= not (a or b);
    layer2_outputs(6127) <= not (a and b);
    layer2_outputs(6128) <= not (a and b);
    layer2_outputs(6129) <= not a;
    layer2_outputs(6130) <= '0';
    layer2_outputs(6131) <= not b or a;
    layer2_outputs(6132) <= b and not a;
    layer2_outputs(6133) <= not (a and b);
    layer2_outputs(6134) <= not (a and b);
    layer2_outputs(6135) <= b;
    layer2_outputs(6136) <= not a;
    layer2_outputs(6137) <= not (a or b);
    layer2_outputs(6138) <= not (a or b);
    layer2_outputs(6139) <= a;
    layer2_outputs(6140) <= not a;
    layer2_outputs(6141) <= '1';
    layer2_outputs(6142) <= a and b;
    layer2_outputs(6143) <= not b or a;
    layer2_outputs(6144) <= not (a and b);
    layer2_outputs(6145) <= not (a or b);
    layer2_outputs(6146) <= a or b;
    layer2_outputs(6147) <= '1';
    layer2_outputs(6148) <= a and not b;
    layer2_outputs(6149) <= b;
    layer2_outputs(6150) <= a or b;
    layer2_outputs(6151) <= not b or a;
    layer2_outputs(6152) <= b and not a;
    layer2_outputs(6153) <= a xor b;
    layer2_outputs(6154) <= b;
    layer2_outputs(6155) <= a and not b;
    layer2_outputs(6156) <= not b or a;
    layer2_outputs(6157) <= '1';
    layer2_outputs(6158) <= not (a or b);
    layer2_outputs(6159) <= not b;
    layer2_outputs(6160) <= not b or a;
    layer2_outputs(6161) <= not b or a;
    layer2_outputs(6162) <= '0';
    layer2_outputs(6163) <= a and b;
    layer2_outputs(6164) <= not (a or b);
    layer2_outputs(6165) <= a and b;
    layer2_outputs(6166) <= a and b;
    layer2_outputs(6167) <= not (a or b);
    layer2_outputs(6168) <= a or b;
    layer2_outputs(6169) <= a;
    layer2_outputs(6170) <= a and not b;
    layer2_outputs(6171) <= b;
    layer2_outputs(6172) <= a or b;
    layer2_outputs(6173) <= not (a or b);
    layer2_outputs(6174) <= '0';
    layer2_outputs(6175) <= b and not a;
    layer2_outputs(6176) <= not b or a;
    layer2_outputs(6177) <= a and b;
    layer2_outputs(6178) <= b and not a;
    layer2_outputs(6179) <= b and not a;
    layer2_outputs(6180) <= b;
    layer2_outputs(6181) <= '1';
    layer2_outputs(6182) <= not (a or b);
    layer2_outputs(6183) <= not b;
    layer2_outputs(6184) <= not (a or b);
    layer2_outputs(6185) <= '1';
    layer2_outputs(6186) <= a;
    layer2_outputs(6187) <= b;
    layer2_outputs(6188) <= a;
    layer2_outputs(6189) <= not (a xor b);
    layer2_outputs(6190) <= '0';
    layer2_outputs(6191) <= b;
    layer2_outputs(6192) <= not (a and b);
    layer2_outputs(6193) <= a;
    layer2_outputs(6194) <= a or b;
    layer2_outputs(6195) <= not (a or b);
    layer2_outputs(6196) <= a and b;
    layer2_outputs(6197) <= b and not a;
    layer2_outputs(6198) <= '0';
    layer2_outputs(6199) <= not a;
    layer2_outputs(6200) <= a and b;
    layer2_outputs(6201) <= a xor b;
    layer2_outputs(6202) <= b and not a;
    layer2_outputs(6203) <= a or b;
    layer2_outputs(6204) <= a and not b;
    layer2_outputs(6205) <= '1';
    layer2_outputs(6206) <= a and not b;
    layer2_outputs(6207) <= a;
    layer2_outputs(6208) <= '0';
    layer2_outputs(6209) <= not (a xor b);
    layer2_outputs(6210) <= b and not a;
    layer2_outputs(6211) <= not b;
    layer2_outputs(6212) <= not (a or b);
    layer2_outputs(6213) <= a or b;
    layer2_outputs(6214) <= b and not a;
    layer2_outputs(6215) <= not (a and b);
    layer2_outputs(6216) <= not b;
    layer2_outputs(6217) <= '1';
    layer2_outputs(6218) <= '1';
    layer2_outputs(6219) <= a and not b;
    layer2_outputs(6220) <= b;
    layer2_outputs(6221) <= a;
    layer2_outputs(6222) <= not (a or b);
    layer2_outputs(6223) <= not (a xor b);
    layer2_outputs(6224) <= b and not a;
    layer2_outputs(6225) <= a or b;
    layer2_outputs(6226) <= not a;
    layer2_outputs(6227) <= '1';
    layer2_outputs(6228) <= not b;
    layer2_outputs(6229) <= '1';
    layer2_outputs(6230) <= b and not a;
    layer2_outputs(6231) <= not b or a;
    layer2_outputs(6232) <= not a;
    layer2_outputs(6233) <= b and not a;
    layer2_outputs(6234) <= b;
    layer2_outputs(6235) <= not (a and b);
    layer2_outputs(6236) <= '1';
    layer2_outputs(6237) <= '1';
    layer2_outputs(6238) <= '0';
    layer2_outputs(6239) <= not b;
    layer2_outputs(6240) <= a and b;
    layer2_outputs(6241) <= not b;
    layer2_outputs(6242) <= not a;
    layer2_outputs(6243) <= a and not b;
    layer2_outputs(6244) <= a and not b;
    layer2_outputs(6245) <= '0';
    layer2_outputs(6246) <= not b;
    layer2_outputs(6247) <= not a or b;
    layer2_outputs(6248) <= not (a or b);
    layer2_outputs(6249) <= '1';
    layer2_outputs(6250) <= '0';
    layer2_outputs(6251) <= a xor b;
    layer2_outputs(6252) <= b and not a;
    layer2_outputs(6253) <= a and not b;
    layer2_outputs(6254) <= b;
    layer2_outputs(6255) <= '0';
    layer2_outputs(6256) <= '0';
    layer2_outputs(6257) <= not a;
    layer2_outputs(6258) <= a or b;
    layer2_outputs(6259) <= a;
    layer2_outputs(6260) <= b and not a;
    layer2_outputs(6261) <= a;
    layer2_outputs(6262) <= not a;
    layer2_outputs(6263) <= a or b;
    layer2_outputs(6264) <= not (a and b);
    layer2_outputs(6265) <= not b;
    layer2_outputs(6266) <= a and not b;
    layer2_outputs(6267) <= a and not b;
    layer2_outputs(6268) <= not b;
    layer2_outputs(6269) <= '0';
    layer2_outputs(6270) <= a and not b;
    layer2_outputs(6271) <= a and not b;
    layer2_outputs(6272) <= not a;
    layer2_outputs(6273) <= a or b;
    layer2_outputs(6274) <= b;
    layer2_outputs(6275) <= a or b;
    layer2_outputs(6276) <= not b;
    layer2_outputs(6277) <= not b or a;
    layer2_outputs(6278) <= not b or a;
    layer2_outputs(6279) <= '0';
    layer2_outputs(6280) <= not b or a;
    layer2_outputs(6281) <= not (a or b);
    layer2_outputs(6282) <= '1';
    layer2_outputs(6283) <= a and not b;
    layer2_outputs(6284) <= not b;
    layer2_outputs(6285) <= not b;
    layer2_outputs(6286) <= a;
    layer2_outputs(6287) <= not (a or b);
    layer2_outputs(6288) <= not b;
    layer2_outputs(6289) <= not a or b;
    layer2_outputs(6290) <= b and not a;
    layer2_outputs(6291) <= a and not b;
    layer2_outputs(6292) <= a or b;
    layer2_outputs(6293) <= a and not b;
    layer2_outputs(6294) <= not b or a;
    layer2_outputs(6295) <= '0';
    layer2_outputs(6296) <= b;
    layer2_outputs(6297) <= a and b;
    layer2_outputs(6298) <= not a;
    layer2_outputs(6299) <= not a or b;
    layer2_outputs(6300) <= a and not b;
    layer2_outputs(6301) <= a xor b;
    layer2_outputs(6302) <= '0';
    layer2_outputs(6303) <= '1';
    layer2_outputs(6304) <= a or b;
    layer2_outputs(6305) <= not b or a;
    layer2_outputs(6306) <= b and not a;
    layer2_outputs(6307) <= not (a and b);
    layer2_outputs(6308) <= a and not b;
    layer2_outputs(6309) <= '1';
    layer2_outputs(6310) <= b and not a;
    layer2_outputs(6311) <= not b or a;
    layer2_outputs(6312) <= '1';
    layer2_outputs(6313) <= not b or a;
    layer2_outputs(6314) <= not a or b;
    layer2_outputs(6315) <= '1';
    layer2_outputs(6316) <= '1';
    layer2_outputs(6317) <= b;
    layer2_outputs(6318) <= not b;
    layer2_outputs(6319) <= '1';
    layer2_outputs(6320) <= a or b;
    layer2_outputs(6321) <= not b;
    layer2_outputs(6322) <= not (a and b);
    layer2_outputs(6323) <= '1';
    layer2_outputs(6324) <= not (a and b);
    layer2_outputs(6325) <= '0';
    layer2_outputs(6326) <= not a or b;
    layer2_outputs(6327) <= a or b;
    layer2_outputs(6328) <= a;
    layer2_outputs(6329) <= a;
    layer2_outputs(6330) <= not (a and b);
    layer2_outputs(6331) <= not (a and b);
    layer2_outputs(6332) <= '0';
    layer2_outputs(6333) <= not (a and b);
    layer2_outputs(6334) <= not (a xor b);
    layer2_outputs(6335) <= a;
    layer2_outputs(6336) <= a or b;
    layer2_outputs(6337) <= not (a or b);
    layer2_outputs(6338) <= b;
    layer2_outputs(6339) <= b and not a;
    layer2_outputs(6340) <= not b;
    layer2_outputs(6341) <= not (a or b);
    layer2_outputs(6342) <= a;
    layer2_outputs(6343) <= '1';
    layer2_outputs(6344) <= not b or a;
    layer2_outputs(6345) <= a and not b;
    layer2_outputs(6346) <= '1';
    layer2_outputs(6347) <= not (a and b);
    layer2_outputs(6348) <= not (a xor b);
    layer2_outputs(6349) <= not a or b;
    layer2_outputs(6350) <= a and not b;
    layer2_outputs(6351) <= a and not b;
    layer2_outputs(6352) <= not a;
    layer2_outputs(6353) <= b;
    layer2_outputs(6354) <= a and b;
    layer2_outputs(6355) <= a and b;
    layer2_outputs(6356) <= a and not b;
    layer2_outputs(6357) <= not b or a;
    layer2_outputs(6358) <= not b;
    layer2_outputs(6359) <= not (a and b);
    layer2_outputs(6360) <= not a;
    layer2_outputs(6361) <= a and not b;
    layer2_outputs(6362) <= a and b;
    layer2_outputs(6363) <= not (a or b);
    layer2_outputs(6364) <= not a;
    layer2_outputs(6365) <= a;
    layer2_outputs(6366) <= '0';
    layer2_outputs(6367) <= '1';
    layer2_outputs(6368) <= '1';
    layer2_outputs(6369) <= not a;
    layer2_outputs(6370) <= b;
    layer2_outputs(6371) <= not a or b;
    layer2_outputs(6372) <= '0';
    layer2_outputs(6373) <= a and b;
    layer2_outputs(6374) <= a or b;
    layer2_outputs(6375) <= not b;
    layer2_outputs(6376) <= a and not b;
    layer2_outputs(6377) <= a and b;
    layer2_outputs(6378) <= not b or a;
    layer2_outputs(6379) <= a or b;
    layer2_outputs(6380) <= not a or b;
    layer2_outputs(6381) <= '0';
    layer2_outputs(6382) <= not (a or b);
    layer2_outputs(6383) <= not a or b;
    layer2_outputs(6384) <= b and not a;
    layer2_outputs(6385) <= '1';
    layer2_outputs(6386) <= not a or b;
    layer2_outputs(6387) <= not b or a;
    layer2_outputs(6388) <= not (a or b);
    layer2_outputs(6389) <= '1';
    layer2_outputs(6390) <= a or b;
    layer2_outputs(6391) <= not a;
    layer2_outputs(6392) <= b;
    layer2_outputs(6393) <= b and not a;
    layer2_outputs(6394) <= '1';
    layer2_outputs(6395) <= a and not b;
    layer2_outputs(6396) <= not a;
    layer2_outputs(6397) <= a and b;
    layer2_outputs(6398) <= not b or a;
    layer2_outputs(6399) <= not b or a;
    layer2_outputs(6400) <= b and not a;
    layer2_outputs(6401) <= not (a and b);
    layer2_outputs(6402) <= b and not a;
    layer2_outputs(6403) <= a and not b;
    layer2_outputs(6404) <= not a or b;
    layer2_outputs(6405) <= not b or a;
    layer2_outputs(6406) <= not (a or b);
    layer2_outputs(6407) <= not a;
    layer2_outputs(6408) <= '1';
    layer2_outputs(6409) <= b and not a;
    layer2_outputs(6410) <= not (a or b);
    layer2_outputs(6411) <= a or b;
    layer2_outputs(6412) <= a and not b;
    layer2_outputs(6413) <= not (a and b);
    layer2_outputs(6414) <= not (a and b);
    layer2_outputs(6415) <= not b;
    layer2_outputs(6416) <= not (a and b);
    layer2_outputs(6417) <= a and not b;
    layer2_outputs(6418) <= a and not b;
    layer2_outputs(6419) <= '1';
    layer2_outputs(6420) <= not (a or b);
    layer2_outputs(6421) <= b;
    layer2_outputs(6422) <= not a or b;
    layer2_outputs(6423) <= not (a or b);
    layer2_outputs(6424) <= not b or a;
    layer2_outputs(6425) <= not (a or b);
    layer2_outputs(6426) <= not b or a;
    layer2_outputs(6427) <= '1';
    layer2_outputs(6428) <= a and not b;
    layer2_outputs(6429) <= a and b;
    layer2_outputs(6430) <= a and not b;
    layer2_outputs(6431) <= '1';
    layer2_outputs(6432) <= not (a and b);
    layer2_outputs(6433) <= '1';
    layer2_outputs(6434) <= not (a or b);
    layer2_outputs(6435) <= not (a xor b);
    layer2_outputs(6436) <= a and b;
    layer2_outputs(6437) <= a or b;
    layer2_outputs(6438) <= '1';
    layer2_outputs(6439) <= '0';
    layer2_outputs(6440) <= a;
    layer2_outputs(6441) <= not (a and b);
    layer2_outputs(6442) <= b;
    layer2_outputs(6443) <= not (a or b);
    layer2_outputs(6444) <= not (a and b);
    layer2_outputs(6445) <= a and not b;
    layer2_outputs(6446) <= not b or a;
    layer2_outputs(6447) <= b;
    layer2_outputs(6448) <= not a;
    layer2_outputs(6449) <= a and not b;
    layer2_outputs(6450) <= '0';
    layer2_outputs(6451) <= not b or a;
    layer2_outputs(6452) <= '1';
    layer2_outputs(6453) <= a and not b;
    layer2_outputs(6454) <= '1';
    layer2_outputs(6455) <= '0';
    layer2_outputs(6456) <= a;
    layer2_outputs(6457) <= not b or a;
    layer2_outputs(6458) <= '1';
    layer2_outputs(6459) <= not a or b;
    layer2_outputs(6460) <= not (a and b);
    layer2_outputs(6461) <= a;
    layer2_outputs(6462) <= not (a and b);
    layer2_outputs(6463) <= '1';
    layer2_outputs(6464) <= a;
    layer2_outputs(6465) <= not a;
    layer2_outputs(6466) <= not b or a;
    layer2_outputs(6467) <= a;
    layer2_outputs(6468) <= not a or b;
    layer2_outputs(6469) <= a and b;
    layer2_outputs(6470) <= '1';
    layer2_outputs(6471) <= not (a or b);
    layer2_outputs(6472) <= b;
    layer2_outputs(6473) <= b;
    layer2_outputs(6474) <= not (a or b);
    layer2_outputs(6475) <= a;
    layer2_outputs(6476) <= not b or a;
    layer2_outputs(6477) <= a and b;
    layer2_outputs(6478) <= a and b;
    layer2_outputs(6479) <= b;
    layer2_outputs(6480) <= not a;
    layer2_outputs(6481) <= not (a and b);
    layer2_outputs(6482) <= a and b;
    layer2_outputs(6483) <= not b or a;
    layer2_outputs(6484) <= a or b;
    layer2_outputs(6485) <= not b;
    layer2_outputs(6486) <= not b;
    layer2_outputs(6487) <= not a;
    layer2_outputs(6488) <= not a or b;
    layer2_outputs(6489) <= a xor b;
    layer2_outputs(6490) <= '0';
    layer2_outputs(6491) <= a and not b;
    layer2_outputs(6492) <= b and not a;
    layer2_outputs(6493) <= not a;
    layer2_outputs(6494) <= a;
    layer2_outputs(6495) <= '0';
    layer2_outputs(6496) <= b and not a;
    layer2_outputs(6497) <= not (a and b);
    layer2_outputs(6498) <= not b or a;
    layer2_outputs(6499) <= b and not a;
    layer2_outputs(6500) <= not b or a;
    layer2_outputs(6501) <= a;
    layer2_outputs(6502) <= not a or b;
    layer2_outputs(6503) <= a or b;
    layer2_outputs(6504) <= not a or b;
    layer2_outputs(6505) <= a;
    layer2_outputs(6506) <= not b or a;
    layer2_outputs(6507) <= not (a and b);
    layer2_outputs(6508) <= a or b;
    layer2_outputs(6509) <= '1';
    layer2_outputs(6510) <= a;
    layer2_outputs(6511) <= a and not b;
    layer2_outputs(6512) <= '0';
    layer2_outputs(6513) <= b;
    layer2_outputs(6514) <= not (a or b);
    layer2_outputs(6515) <= not (a or b);
    layer2_outputs(6516) <= b;
    layer2_outputs(6517) <= a or b;
    layer2_outputs(6518) <= a or b;
    layer2_outputs(6519) <= not a;
    layer2_outputs(6520) <= not (a and b);
    layer2_outputs(6521) <= b and not a;
    layer2_outputs(6522) <= '0';
    layer2_outputs(6523) <= a and b;
    layer2_outputs(6524) <= not b;
    layer2_outputs(6525) <= a and not b;
    layer2_outputs(6526) <= not b;
    layer2_outputs(6527) <= a;
    layer2_outputs(6528) <= a and not b;
    layer2_outputs(6529) <= b;
    layer2_outputs(6530) <= a xor b;
    layer2_outputs(6531) <= '1';
    layer2_outputs(6532) <= a and b;
    layer2_outputs(6533) <= not b;
    layer2_outputs(6534) <= not a or b;
    layer2_outputs(6535) <= a;
    layer2_outputs(6536) <= a;
    layer2_outputs(6537) <= not a or b;
    layer2_outputs(6538) <= a or b;
    layer2_outputs(6539) <= a and b;
    layer2_outputs(6540) <= '0';
    layer2_outputs(6541) <= a;
    layer2_outputs(6542) <= b and not a;
    layer2_outputs(6543) <= a;
    layer2_outputs(6544) <= a and not b;
    layer2_outputs(6545) <= not (a or b);
    layer2_outputs(6546) <= a;
    layer2_outputs(6547) <= not (a and b);
    layer2_outputs(6548) <= b and not a;
    layer2_outputs(6549) <= not b;
    layer2_outputs(6550) <= not b or a;
    layer2_outputs(6551) <= not (a or b);
    layer2_outputs(6552) <= a and b;
    layer2_outputs(6553) <= not b;
    layer2_outputs(6554) <= not (a and b);
    layer2_outputs(6555) <= b;
    layer2_outputs(6556) <= a xor b;
    layer2_outputs(6557) <= not (a or b);
    layer2_outputs(6558) <= not (a or b);
    layer2_outputs(6559) <= '0';
    layer2_outputs(6560) <= b;
    layer2_outputs(6561) <= b;
    layer2_outputs(6562) <= b and not a;
    layer2_outputs(6563) <= not a or b;
    layer2_outputs(6564) <= a;
    layer2_outputs(6565) <= not a;
    layer2_outputs(6566) <= b and not a;
    layer2_outputs(6567) <= not (a or b);
    layer2_outputs(6568) <= b and not a;
    layer2_outputs(6569) <= not b or a;
    layer2_outputs(6570) <= a;
    layer2_outputs(6571) <= not a;
    layer2_outputs(6572) <= a or b;
    layer2_outputs(6573) <= a or b;
    layer2_outputs(6574) <= not b;
    layer2_outputs(6575) <= b and not a;
    layer2_outputs(6576) <= '1';
    layer2_outputs(6577) <= a;
    layer2_outputs(6578) <= a and b;
    layer2_outputs(6579) <= '1';
    layer2_outputs(6580) <= b;
    layer2_outputs(6581) <= not a or b;
    layer2_outputs(6582) <= not a;
    layer2_outputs(6583) <= a;
    layer2_outputs(6584) <= b;
    layer2_outputs(6585) <= not (a and b);
    layer2_outputs(6586) <= a or b;
    layer2_outputs(6587) <= a and b;
    layer2_outputs(6588) <= a or b;
    layer2_outputs(6589) <= a and b;
    layer2_outputs(6590) <= not b;
    layer2_outputs(6591) <= '0';
    layer2_outputs(6592) <= not (a and b);
    layer2_outputs(6593) <= not a;
    layer2_outputs(6594) <= a or b;
    layer2_outputs(6595) <= '1';
    layer2_outputs(6596) <= not a;
    layer2_outputs(6597) <= not b;
    layer2_outputs(6598) <= not a;
    layer2_outputs(6599) <= b;
    layer2_outputs(6600) <= not (a and b);
    layer2_outputs(6601) <= b;
    layer2_outputs(6602) <= b;
    layer2_outputs(6603) <= b and not a;
    layer2_outputs(6604) <= b;
    layer2_outputs(6605) <= a or b;
    layer2_outputs(6606) <= a and not b;
    layer2_outputs(6607) <= not b or a;
    layer2_outputs(6608) <= b and not a;
    layer2_outputs(6609) <= not b or a;
    layer2_outputs(6610) <= not (a or b);
    layer2_outputs(6611) <= a and not b;
    layer2_outputs(6612) <= not a or b;
    layer2_outputs(6613) <= not (a and b);
    layer2_outputs(6614) <= not a;
    layer2_outputs(6615) <= '1';
    layer2_outputs(6616) <= not b or a;
    layer2_outputs(6617) <= not b or a;
    layer2_outputs(6618) <= a or b;
    layer2_outputs(6619) <= '1';
    layer2_outputs(6620) <= a;
    layer2_outputs(6621) <= not a;
    layer2_outputs(6622) <= '1';
    layer2_outputs(6623) <= '0';
    layer2_outputs(6624) <= not (a and b);
    layer2_outputs(6625) <= a xor b;
    layer2_outputs(6626) <= '0';
    layer2_outputs(6627) <= a or b;
    layer2_outputs(6628) <= b and not a;
    layer2_outputs(6629) <= not a;
    layer2_outputs(6630) <= a and not b;
    layer2_outputs(6631) <= not (a and b);
    layer2_outputs(6632) <= b;
    layer2_outputs(6633) <= not (a or b);
    layer2_outputs(6634) <= a and not b;
    layer2_outputs(6635) <= b and not a;
    layer2_outputs(6636) <= not (a or b);
    layer2_outputs(6637) <= a and b;
    layer2_outputs(6638) <= a or b;
    layer2_outputs(6639) <= a or b;
    layer2_outputs(6640) <= a;
    layer2_outputs(6641) <= a or b;
    layer2_outputs(6642) <= '0';
    layer2_outputs(6643) <= b;
    layer2_outputs(6644) <= not (a or b);
    layer2_outputs(6645) <= a or b;
    layer2_outputs(6646) <= b;
    layer2_outputs(6647) <= not (a or b);
    layer2_outputs(6648) <= a and b;
    layer2_outputs(6649) <= not a or b;
    layer2_outputs(6650) <= not a or b;
    layer2_outputs(6651) <= not (a or b);
    layer2_outputs(6652) <= b and not a;
    layer2_outputs(6653) <= a;
    layer2_outputs(6654) <= not a or b;
    layer2_outputs(6655) <= b;
    layer2_outputs(6656) <= not a or b;
    layer2_outputs(6657) <= not a;
    layer2_outputs(6658) <= a and not b;
    layer2_outputs(6659) <= a;
    layer2_outputs(6660) <= a and b;
    layer2_outputs(6661) <= b;
    layer2_outputs(6662) <= '1';
    layer2_outputs(6663) <= not a or b;
    layer2_outputs(6664) <= not b or a;
    layer2_outputs(6665) <= not (a and b);
    layer2_outputs(6666) <= a;
    layer2_outputs(6667) <= '0';
    layer2_outputs(6668) <= a;
    layer2_outputs(6669) <= a or b;
    layer2_outputs(6670) <= a;
    layer2_outputs(6671) <= not a;
    layer2_outputs(6672) <= b and not a;
    layer2_outputs(6673) <= not b or a;
    layer2_outputs(6674) <= not b;
    layer2_outputs(6675) <= not (a and b);
    layer2_outputs(6676) <= not (a and b);
    layer2_outputs(6677) <= a or b;
    layer2_outputs(6678) <= a or b;
    layer2_outputs(6679) <= not (a and b);
    layer2_outputs(6680) <= '1';
    layer2_outputs(6681) <= b;
    layer2_outputs(6682) <= a and b;
    layer2_outputs(6683) <= not b;
    layer2_outputs(6684) <= not a or b;
    layer2_outputs(6685) <= '0';
    layer2_outputs(6686) <= not a or b;
    layer2_outputs(6687) <= not (a or b);
    layer2_outputs(6688) <= '0';
    layer2_outputs(6689) <= b;
    layer2_outputs(6690) <= not (a or b);
    layer2_outputs(6691) <= a and b;
    layer2_outputs(6692) <= a and not b;
    layer2_outputs(6693) <= a and b;
    layer2_outputs(6694) <= a and b;
    layer2_outputs(6695) <= a and not b;
    layer2_outputs(6696) <= b;
    layer2_outputs(6697) <= '0';
    layer2_outputs(6698) <= a xor b;
    layer2_outputs(6699) <= not (a and b);
    layer2_outputs(6700) <= '1';
    layer2_outputs(6701) <= not a or b;
    layer2_outputs(6702) <= not (a or b);
    layer2_outputs(6703) <= not (a and b);
    layer2_outputs(6704) <= a or b;
    layer2_outputs(6705) <= not b or a;
    layer2_outputs(6706) <= a or b;
    layer2_outputs(6707) <= not b;
    layer2_outputs(6708) <= a xor b;
    layer2_outputs(6709) <= not a;
    layer2_outputs(6710) <= not b or a;
    layer2_outputs(6711) <= not (a or b);
    layer2_outputs(6712) <= a and b;
    layer2_outputs(6713) <= not (a xor b);
    layer2_outputs(6714) <= a or b;
    layer2_outputs(6715) <= not a or b;
    layer2_outputs(6716) <= not (a or b);
    layer2_outputs(6717) <= a and not b;
    layer2_outputs(6718) <= not b or a;
    layer2_outputs(6719) <= not b or a;
    layer2_outputs(6720) <= not (a xor b);
    layer2_outputs(6721) <= '0';
    layer2_outputs(6722) <= not b;
    layer2_outputs(6723) <= not (a or b);
    layer2_outputs(6724) <= b;
    layer2_outputs(6725) <= b;
    layer2_outputs(6726) <= a and not b;
    layer2_outputs(6727) <= '1';
    layer2_outputs(6728) <= a and b;
    layer2_outputs(6729) <= not b;
    layer2_outputs(6730) <= b;
    layer2_outputs(6731) <= a or b;
    layer2_outputs(6732) <= b;
    layer2_outputs(6733) <= not b;
    layer2_outputs(6734) <= '0';
    layer2_outputs(6735) <= '1';
    layer2_outputs(6736) <= not b or a;
    layer2_outputs(6737) <= a and b;
    layer2_outputs(6738) <= a and not b;
    layer2_outputs(6739) <= a or b;
    layer2_outputs(6740) <= not a or b;
    layer2_outputs(6741) <= '1';
    layer2_outputs(6742) <= not a or b;
    layer2_outputs(6743) <= '0';
    layer2_outputs(6744) <= not b;
    layer2_outputs(6745) <= a or b;
    layer2_outputs(6746) <= not a;
    layer2_outputs(6747) <= not (a or b);
    layer2_outputs(6748) <= '0';
    layer2_outputs(6749) <= not b;
    layer2_outputs(6750) <= not a;
    layer2_outputs(6751) <= a xor b;
    layer2_outputs(6752) <= a xor b;
    layer2_outputs(6753) <= b;
    layer2_outputs(6754) <= not a;
    layer2_outputs(6755) <= '1';
    layer2_outputs(6756) <= a and not b;
    layer2_outputs(6757) <= b;
    layer2_outputs(6758) <= '0';
    layer2_outputs(6759) <= '0';
    layer2_outputs(6760) <= not b;
    layer2_outputs(6761) <= '0';
    layer2_outputs(6762) <= b and not a;
    layer2_outputs(6763) <= b;
    layer2_outputs(6764) <= not (a or b);
    layer2_outputs(6765) <= not b;
    layer2_outputs(6766) <= not (a and b);
    layer2_outputs(6767) <= not (a and b);
    layer2_outputs(6768) <= a or b;
    layer2_outputs(6769) <= b;
    layer2_outputs(6770) <= b;
    layer2_outputs(6771) <= not (a xor b);
    layer2_outputs(6772) <= not (a and b);
    layer2_outputs(6773) <= b and not a;
    layer2_outputs(6774) <= not b;
    layer2_outputs(6775) <= not (a xor b);
    layer2_outputs(6776) <= not a;
    layer2_outputs(6777) <= not b;
    layer2_outputs(6778) <= not (a and b);
    layer2_outputs(6779) <= a;
    layer2_outputs(6780) <= '1';
    layer2_outputs(6781) <= not (a and b);
    layer2_outputs(6782) <= not (a and b);
    layer2_outputs(6783) <= not (a or b);
    layer2_outputs(6784) <= not b;
    layer2_outputs(6785) <= not a;
    layer2_outputs(6786) <= a xor b;
    layer2_outputs(6787) <= not (a or b);
    layer2_outputs(6788) <= b and not a;
    layer2_outputs(6789) <= a and not b;
    layer2_outputs(6790) <= not a or b;
    layer2_outputs(6791) <= '0';
    layer2_outputs(6792) <= not b;
    layer2_outputs(6793) <= a and b;
    layer2_outputs(6794) <= '0';
    layer2_outputs(6795) <= '1';
    layer2_outputs(6796) <= a or b;
    layer2_outputs(6797) <= a xor b;
    layer2_outputs(6798) <= '1';
    layer2_outputs(6799) <= not (a xor b);
    layer2_outputs(6800) <= b and not a;
    layer2_outputs(6801) <= not (a and b);
    layer2_outputs(6802) <= b;
    layer2_outputs(6803) <= a and not b;
    layer2_outputs(6804) <= '0';
    layer2_outputs(6805) <= '1';
    layer2_outputs(6806) <= '1';
    layer2_outputs(6807) <= b;
    layer2_outputs(6808) <= not (a and b);
    layer2_outputs(6809) <= a and b;
    layer2_outputs(6810) <= a and b;
    layer2_outputs(6811) <= b and not a;
    layer2_outputs(6812) <= not (a or b);
    layer2_outputs(6813) <= not a or b;
    layer2_outputs(6814) <= not (a and b);
    layer2_outputs(6815) <= a;
    layer2_outputs(6816) <= a or b;
    layer2_outputs(6817) <= a and b;
    layer2_outputs(6818) <= a and b;
    layer2_outputs(6819) <= not b or a;
    layer2_outputs(6820) <= not a or b;
    layer2_outputs(6821) <= not (a or b);
    layer2_outputs(6822) <= not (a or b);
    layer2_outputs(6823) <= not b or a;
    layer2_outputs(6824) <= b;
    layer2_outputs(6825) <= a and not b;
    layer2_outputs(6826) <= a;
    layer2_outputs(6827) <= '0';
    layer2_outputs(6828) <= a and b;
    layer2_outputs(6829) <= a and b;
    layer2_outputs(6830) <= not a;
    layer2_outputs(6831) <= not a or b;
    layer2_outputs(6832) <= b and not a;
    layer2_outputs(6833) <= not a;
    layer2_outputs(6834) <= b;
    layer2_outputs(6835) <= '1';
    layer2_outputs(6836) <= not b;
    layer2_outputs(6837) <= a;
    layer2_outputs(6838) <= not b or a;
    layer2_outputs(6839) <= not b;
    layer2_outputs(6840) <= not a or b;
    layer2_outputs(6841) <= not b or a;
    layer2_outputs(6842) <= '0';
    layer2_outputs(6843) <= not b or a;
    layer2_outputs(6844) <= not (a or b);
    layer2_outputs(6845) <= a and not b;
    layer2_outputs(6846) <= not (a xor b);
    layer2_outputs(6847) <= not b or a;
    layer2_outputs(6848) <= a xor b;
    layer2_outputs(6849) <= a and b;
    layer2_outputs(6850) <= not b;
    layer2_outputs(6851) <= '0';
    layer2_outputs(6852) <= a;
    layer2_outputs(6853) <= '1';
    layer2_outputs(6854) <= a or b;
    layer2_outputs(6855) <= not b or a;
    layer2_outputs(6856) <= not (a xor b);
    layer2_outputs(6857) <= not b or a;
    layer2_outputs(6858) <= not b or a;
    layer2_outputs(6859) <= not (a and b);
    layer2_outputs(6860) <= '0';
    layer2_outputs(6861) <= not (a or b);
    layer2_outputs(6862) <= a and b;
    layer2_outputs(6863) <= a;
    layer2_outputs(6864) <= a or b;
    layer2_outputs(6865) <= not (a and b);
    layer2_outputs(6866) <= b and not a;
    layer2_outputs(6867) <= a and not b;
    layer2_outputs(6868) <= '1';
    layer2_outputs(6869) <= a and not b;
    layer2_outputs(6870) <= not (a and b);
    layer2_outputs(6871) <= not (a and b);
    layer2_outputs(6872) <= a and b;
    layer2_outputs(6873) <= not (a and b);
    layer2_outputs(6874) <= not b;
    layer2_outputs(6875) <= not a;
    layer2_outputs(6876) <= a and b;
    layer2_outputs(6877) <= b;
    layer2_outputs(6878) <= '0';
    layer2_outputs(6879) <= not (a or b);
    layer2_outputs(6880) <= '1';
    layer2_outputs(6881) <= not a;
    layer2_outputs(6882) <= a or b;
    layer2_outputs(6883) <= b and not a;
    layer2_outputs(6884) <= a xor b;
    layer2_outputs(6885) <= '1';
    layer2_outputs(6886) <= not a;
    layer2_outputs(6887) <= b;
    layer2_outputs(6888) <= a or b;
    layer2_outputs(6889) <= not a;
    layer2_outputs(6890) <= not (a and b);
    layer2_outputs(6891) <= not a;
    layer2_outputs(6892) <= not b;
    layer2_outputs(6893) <= not (a and b);
    layer2_outputs(6894) <= not (a or b);
    layer2_outputs(6895) <= a xor b;
    layer2_outputs(6896) <= not b;
    layer2_outputs(6897) <= b and not a;
    layer2_outputs(6898) <= not (a or b);
    layer2_outputs(6899) <= a and not b;
    layer2_outputs(6900) <= a;
    layer2_outputs(6901) <= not (a or b);
    layer2_outputs(6902) <= a or b;
    layer2_outputs(6903) <= a or b;
    layer2_outputs(6904) <= b and not a;
    layer2_outputs(6905) <= a;
    layer2_outputs(6906) <= '0';
    layer2_outputs(6907) <= '1';
    layer2_outputs(6908) <= not a or b;
    layer2_outputs(6909) <= a and b;
    layer2_outputs(6910) <= a and not b;
    layer2_outputs(6911) <= not (a or b);
    layer2_outputs(6912) <= '0';
    layer2_outputs(6913) <= '0';
    layer2_outputs(6914) <= a and b;
    layer2_outputs(6915) <= not a or b;
    layer2_outputs(6916) <= b;
    layer2_outputs(6917) <= b;
    layer2_outputs(6918) <= not b or a;
    layer2_outputs(6919) <= not a or b;
    layer2_outputs(6920) <= not (a and b);
    layer2_outputs(6921) <= not a;
    layer2_outputs(6922) <= a and not b;
    layer2_outputs(6923) <= b and not a;
    layer2_outputs(6924) <= b and not a;
    layer2_outputs(6925) <= not a or b;
    layer2_outputs(6926) <= a or b;
    layer2_outputs(6927) <= not (a or b);
    layer2_outputs(6928) <= '0';
    layer2_outputs(6929) <= '1';
    layer2_outputs(6930) <= a or b;
    layer2_outputs(6931) <= a and not b;
    layer2_outputs(6932) <= not b;
    layer2_outputs(6933) <= not (a or b);
    layer2_outputs(6934) <= not (a or b);
    layer2_outputs(6935) <= a and not b;
    layer2_outputs(6936) <= not b or a;
    layer2_outputs(6937) <= b and not a;
    layer2_outputs(6938) <= not b or a;
    layer2_outputs(6939) <= '0';
    layer2_outputs(6940) <= not b;
    layer2_outputs(6941) <= '0';
    layer2_outputs(6942) <= not a;
    layer2_outputs(6943) <= '0';
    layer2_outputs(6944) <= not (a xor b);
    layer2_outputs(6945) <= a or b;
    layer2_outputs(6946) <= a;
    layer2_outputs(6947) <= not (a or b);
    layer2_outputs(6948) <= b and not a;
    layer2_outputs(6949) <= a and not b;
    layer2_outputs(6950) <= not a or b;
    layer2_outputs(6951) <= not (a or b);
    layer2_outputs(6952) <= a and b;
    layer2_outputs(6953) <= not a;
    layer2_outputs(6954) <= b and not a;
    layer2_outputs(6955) <= not a;
    layer2_outputs(6956) <= a;
    layer2_outputs(6957) <= a;
    layer2_outputs(6958) <= a and b;
    layer2_outputs(6959) <= not a or b;
    layer2_outputs(6960) <= b;
    layer2_outputs(6961) <= b and not a;
    layer2_outputs(6962) <= b;
    layer2_outputs(6963) <= not (a and b);
    layer2_outputs(6964) <= not (a or b);
    layer2_outputs(6965) <= not b;
    layer2_outputs(6966) <= not a;
    layer2_outputs(6967) <= '0';
    layer2_outputs(6968) <= not b or a;
    layer2_outputs(6969) <= a and b;
    layer2_outputs(6970) <= b and not a;
    layer2_outputs(6971) <= a or b;
    layer2_outputs(6972) <= not b or a;
    layer2_outputs(6973) <= a or b;
    layer2_outputs(6974) <= b;
    layer2_outputs(6975) <= '1';
    layer2_outputs(6976) <= not b;
    layer2_outputs(6977) <= not a or b;
    layer2_outputs(6978) <= not (a or b);
    layer2_outputs(6979) <= not a or b;
    layer2_outputs(6980) <= '1';
    layer2_outputs(6981) <= b;
    layer2_outputs(6982) <= not a or b;
    layer2_outputs(6983) <= '0';
    layer2_outputs(6984) <= '1';
    layer2_outputs(6985) <= a and not b;
    layer2_outputs(6986) <= a and b;
    layer2_outputs(6987) <= not a or b;
    layer2_outputs(6988) <= a or b;
    layer2_outputs(6989) <= not b;
    layer2_outputs(6990) <= not (a or b);
    layer2_outputs(6991) <= '1';
    layer2_outputs(6992) <= '0';
    layer2_outputs(6993) <= b;
    layer2_outputs(6994) <= '0';
    layer2_outputs(6995) <= '1';
    layer2_outputs(6996) <= b;
    layer2_outputs(6997) <= not a;
    layer2_outputs(6998) <= not a or b;
    layer2_outputs(6999) <= '1';
    layer2_outputs(7000) <= not (a and b);
    layer2_outputs(7001) <= b;
    layer2_outputs(7002) <= a and b;
    layer2_outputs(7003) <= not a;
    layer2_outputs(7004) <= a and not b;
    layer2_outputs(7005) <= '1';
    layer2_outputs(7006) <= '1';
    layer2_outputs(7007) <= not b or a;
    layer2_outputs(7008) <= not (a or b);
    layer2_outputs(7009) <= not b;
    layer2_outputs(7010) <= '1';
    layer2_outputs(7011) <= not a or b;
    layer2_outputs(7012) <= not (a or b);
    layer2_outputs(7013) <= b and not a;
    layer2_outputs(7014) <= a xor b;
    layer2_outputs(7015) <= a;
    layer2_outputs(7016) <= '1';
    layer2_outputs(7017) <= b and not a;
    layer2_outputs(7018) <= a or b;
    layer2_outputs(7019) <= a and not b;
    layer2_outputs(7020) <= a and b;
    layer2_outputs(7021) <= not b or a;
    layer2_outputs(7022) <= a and b;
    layer2_outputs(7023) <= '1';
    layer2_outputs(7024) <= not b or a;
    layer2_outputs(7025) <= not (a xor b);
    layer2_outputs(7026) <= '1';
    layer2_outputs(7027) <= a and b;
    layer2_outputs(7028) <= not a;
    layer2_outputs(7029) <= not a;
    layer2_outputs(7030) <= '1';
    layer2_outputs(7031) <= '0';
    layer2_outputs(7032) <= not b or a;
    layer2_outputs(7033) <= not b;
    layer2_outputs(7034) <= not (a or b);
    layer2_outputs(7035) <= '0';
    layer2_outputs(7036) <= '1';
    layer2_outputs(7037) <= not (a and b);
    layer2_outputs(7038) <= not b;
    layer2_outputs(7039) <= a and not b;
    layer2_outputs(7040) <= not (a and b);
    layer2_outputs(7041) <= a or b;
    layer2_outputs(7042) <= a or b;
    layer2_outputs(7043) <= not a;
    layer2_outputs(7044) <= b;
    layer2_outputs(7045) <= b and not a;
    layer2_outputs(7046) <= not a;
    layer2_outputs(7047) <= b;
    layer2_outputs(7048) <= not (a or b);
    layer2_outputs(7049) <= b and not a;
    layer2_outputs(7050) <= not a;
    layer2_outputs(7051) <= a;
    layer2_outputs(7052) <= '0';
    layer2_outputs(7053) <= not b or a;
    layer2_outputs(7054) <= not b or a;
    layer2_outputs(7055) <= not (a and b);
    layer2_outputs(7056) <= '1';
    layer2_outputs(7057) <= not (a or b);
    layer2_outputs(7058) <= a and not b;
    layer2_outputs(7059) <= '0';
    layer2_outputs(7060) <= '1';
    layer2_outputs(7061) <= '1';
    layer2_outputs(7062) <= '0';
    layer2_outputs(7063) <= not (a xor b);
    layer2_outputs(7064) <= not (a and b);
    layer2_outputs(7065) <= not b;
    layer2_outputs(7066) <= not (a xor b);
    layer2_outputs(7067) <= '1';
    layer2_outputs(7068) <= b and not a;
    layer2_outputs(7069) <= b;
    layer2_outputs(7070) <= '1';
    layer2_outputs(7071) <= a xor b;
    layer2_outputs(7072) <= '0';
    layer2_outputs(7073) <= a or b;
    layer2_outputs(7074) <= a xor b;
    layer2_outputs(7075) <= a;
    layer2_outputs(7076) <= not (a or b);
    layer2_outputs(7077) <= not (a xor b);
    layer2_outputs(7078) <= '1';
    layer2_outputs(7079) <= a;
    layer2_outputs(7080) <= not (a or b);
    layer2_outputs(7081) <= b and not a;
    layer2_outputs(7082) <= a or b;
    layer2_outputs(7083) <= '0';
    layer2_outputs(7084) <= a;
    layer2_outputs(7085) <= b and not a;
    layer2_outputs(7086) <= not b or a;
    layer2_outputs(7087) <= not b;
    layer2_outputs(7088) <= not b;
    layer2_outputs(7089) <= '1';
    layer2_outputs(7090) <= not b or a;
    layer2_outputs(7091) <= not (a and b);
    layer2_outputs(7092) <= a;
    layer2_outputs(7093) <= '1';
    layer2_outputs(7094) <= not a or b;
    layer2_outputs(7095) <= not a;
    layer2_outputs(7096) <= not (a or b);
    layer2_outputs(7097) <= a;
    layer2_outputs(7098) <= not (a xor b);
    layer2_outputs(7099) <= a;
    layer2_outputs(7100) <= not a;
    layer2_outputs(7101) <= '1';
    layer2_outputs(7102) <= a;
    layer2_outputs(7103) <= '1';
    layer2_outputs(7104) <= not a or b;
    layer2_outputs(7105) <= not b;
    layer2_outputs(7106) <= '1';
    layer2_outputs(7107) <= not b;
    layer2_outputs(7108) <= '0';
    layer2_outputs(7109) <= a;
    layer2_outputs(7110) <= b;
    layer2_outputs(7111) <= b and not a;
    layer2_outputs(7112) <= b;
    layer2_outputs(7113) <= not a or b;
    layer2_outputs(7114) <= not b;
    layer2_outputs(7115) <= a and not b;
    layer2_outputs(7116) <= not a or b;
    layer2_outputs(7117) <= a;
    layer2_outputs(7118) <= not a or b;
    layer2_outputs(7119) <= '1';
    layer2_outputs(7120) <= '0';
    layer2_outputs(7121) <= '1';
    layer2_outputs(7122) <= b;
    layer2_outputs(7123) <= '0';
    layer2_outputs(7124) <= a or b;
    layer2_outputs(7125) <= not a;
    layer2_outputs(7126) <= a or b;
    layer2_outputs(7127) <= not b or a;
    layer2_outputs(7128) <= a;
    layer2_outputs(7129) <= not (a or b);
    layer2_outputs(7130) <= not (a or b);
    layer2_outputs(7131) <= '1';
    layer2_outputs(7132) <= not (a and b);
    layer2_outputs(7133) <= b;
    layer2_outputs(7134) <= a or b;
    layer2_outputs(7135) <= a;
    layer2_outputs(7136) <= '1';
    layer2_outputs(7137) <= not (a and b);
    layer2_outputs(7138) <= '0';
    layer2_outputs(7139) <= '1';
    layer2_outputs(7140) <= not b;
    layer2_outputs(7141) <= not b or a;
    layer2_outputs(7142) <= b;
    layer2_outputs(7143) <= '0';
    layer2_outputs(7144) <= a;
    layer2_outputs(7145) <= not a or b;
    layer2_outputs(7146) <= not a;
    layer2_outputs(7147) <= a and b;
    layer2_outputs(7148) <= not (a and b);
    layer2_outputs(7149) <= '0';
    layer2_outputs(7150) <= a and b;
    layer2_outputs(7151) <= a or b;
    layer2_outputs(7152) <= '0';
    layer2_outputs(7153) <= a and not b;
    layer2_outputs(7154) <= a and b;
    layer2_outputs(7155) <= a;
    layer2_outputs(7156) <= a;
    layer2_outputs(7157) <= '1';
    layer2_outputs(7158) <= a;
    layer2_outputs(7159) <= not a or b;
    layer2_outputs(7160) <= not b or a;
    layer2_outputs(7161) <= a or b;
    layer2_outputs(7162) <= '0';
    layer2_outputs(7163) <= a and not b;
    layer2_outputs(7164) <= not b or a;
    layer2_outputs(7165) <= not a;
    layer2_outputs(7166) <= a or b;
    layer2_outputs(7167) <= not (a or b);
    layer2_outputs(7168) <= a and b;
    layer2_outputs(7169) <= a and b;
    layer2_outputs(7170) <= not (a or b);
    layer2_outputs(7171) <= b;
    layer2_outputs(7172) <= not (a and b);
    layer2_outputs(7173) <= not (a and b);
    layer2_outputs(7174) <= not a;
    layer2_outputs(7175) <= a and not b;
    layer2_outputs(7176) <= not (a and b);
    layer2_outputs(7177) <= '1';
    layer2_outputs(7178) <= not (a or b);
    layer2_outputs(7179) <= a or b;
    layer2_outputs(7180) <= not (a and b);
    layer2_outputs(7181) <= not b;
    layer2_outputs(7182) <= not b or a;
    layer2_outputs(7183) <= not b;
    layer2_outputs(7184) <= '1';
    layer2_outputs(7185) <= not b;
    layer2_outputs(7186) <= a or b;
    layer2_outputs(7187) <= not a or b;
    layer2_outputs(7188) <= a or b;
    layer2_outputs(7189) <= a and not b;
    layer2_outputs(7190) <= not (a or b);
    layer2_outputs(7191) <= not (a or b);
    layer2_outputs(7192) <= '1';
    layer2_outputs(7193) <= a xor b;
    layer2_outputs(7194) <= '1';
    layer2_outputs(7195) <= not (a or b);
    layer2_outputs(7196) <= a;
    layer2_outputs(7197) <= a and b;
    layer2_outputs(7198) <= not (a and b);
    layer2_outputs(7199) <= a or b;
    layer2_outputs(7200) <= a or b;
    layer2_outputs(7201) <= b and not a;
    layer2_outputs(7202) <= '1';
    layer2_outputs(7203) <= a and not b;
    layer2_outputs(7204) <= not (a and b);
    layer2_outputs(7205) <= b;
    layer2_outputs(7206) <= '1';
    layer2_outputs(7207) <= a xor b;
    layer2_outputs(7208) <= b;
    layer2_outputs(7209) <= not a;
    layer2_outputs(7210) <= a and not b;
    layer2_outputs(7211) <= a and not b;
    layer2_outputs(7212) <= '1';
    layer2_outputs(7213) <= b and not a;
    layer2_outputs(7214) <= '1';
    layer2_outputs(7215) <= a;
    layer2_outputs(7216) <= not a or b;
    layer2_outputs(7217) <= not a;
    layer2_outputs(7218) <= not (a or b);
    layer2_outputs(7219) <= not (a or b);
    layer2_outputs(7220) <= not (a xor b);
    layer2_outputs(7221) <= b;
    layer2_outputs(7222) <= not a or b;
    layer2_outputs(7223) <= a;
    layer2_outputs(7224) <= '1';
    layer2_outputs(7225) <= a and b;
    layer2_outputs(7226) <= '0';
    layer2_outputs(7227) <= not (a xor b);
    layer2_outputs(7228) <= b;
    layer2_outputs(7229) <= not b;
    layer2_outputs(7230) <= not b;
    layer2_outputs(7231) <= not (a and b);
    layer2_outputs(7232) <= not b;
    layer2_outputs(7233) <= not a;
    layer2_outputs(7234) <= not b;
    layer2_outputs(7235) <= not a or b;
    layer2_outputs(7236) <= b;
    layer2_outputs(7237) <= not a;
    layer2_outputs(7238) <= not b;
    layer2_outputs(7239) <= a and b;
    layer2_outputs(7240) <= not (a and b);
    layer2_outputs(7241) <= a or b;
    layer2_outputs(7242) <= '0';
    layer2_outputs(7243) <= b and not a;
    layer2_outputs(7244) <= a or b;
    layer2_outputs(7245) <= b and not a;
    layer2_outputs(7246) <= not b;
    layer2_outputs(7247) <= not a;
    layer2_outputs(7248) <= not (a xor b);
    layer2_outputs(7249) <= not b;
    layer2_outputs(7250) <= not (a and b);
    layer2_outputs(7251) <= not (a or b);
    layer2_outputs(7252) <= not (a or b);
    layer2_outputs(7253) <= not a or b;
    layer2_outputs(7254) <= '1';
    layer2_outputs(7255) <= b and not a;
    layer2_outputs(7256) <= a and not b;
    layer2_outputs(7257) <= not b or a;
    layer2_outputs(7258) <= not a;
    layer2_outputs(7259) <= not a;
    layer2_outputs(7260) <= not (a xor b);
    layer2_outputs(7261) <= not a or b;
    layer2_outputs(7262) <= '0';
    layer2_outputs(7263) <= '1';
    layer2_outputs(7264) <= not a;
    layer2_outputs(7265) <= a;
    layer2_outputs(7266) <= not b;
    layer2_outputs(7267) <= a xor b;
    layer2_outputs(7268) <= not a or b;
    layer2_outputs(7269) <= not (a and b);
    layer2_outputs(7270) <= b;
    layer2_outputs(7271) <= not a;
    layer2_outputs(7272) <= a or b;
    layer2_outputs(7273) <= not b or a;
    layer2_outputs(7274) <= a or b;
    layer2_outputs(7275) <= '0';
    layer2_outputs(7276) <= a;
    layer2_outputs(7277) <= b and not a;
    layer2_outputs(7278) <= not b or a;
    layer2_outputs(7279) <= not b;
    layer2_outputs(7280) <= not (a and b);
    layer2_outputs(7281) <= b and not a;
    layer2_outputs(7282) <= not (a and b);
    layer2_outputs(7283) <= a or b;
    layer2_outputs(7284) <= not (a or b);
    layer2_outputs(7285) <= b and not a;
    layer2_outputs(7286) <= not a;
    layer2_outputs(7287) <= '0';
    layer2_outputs(7288) <= a or b;
    layer2_outputs(7289) <= b and not a;
    layer2_outputs(7290) <= a;
    layer2_outputs(7291) <= '1';
    layer2_outputs(7292) <= a and not b;
    layer2_outputs(7293) <= a;
    layer2_outputs(7294) <= a or b;
    layer2_outputs(7295) <= not (a xor b);
    layer2_outputs(7296) <= not b;
    layer2_outputs(7297) <= not b;
    layer2_outputs(7298) <= not b or a;
    layer2_outputs(7299) <= not (a xor b);
    layer2_outputs(7300) <= a;
    layer2_outputs(7301) <= not a;
    layer2_outputs(7302) <= not b;
    layer2_outputs(7303) <= not a or b;
    layer2_outputs(7304) <= not a;
    layer2_outputs(7305) <= b and not a;
    layer2_outputs(7306) <= a;
    layer2_outputs(7307) <= '0';
    layer2_outputs(7308) <= '1';
    layer2_outputs(7309) <= not a;
    layer2_outputs(7310) <= a or b;
    layer2_outputs(7311) <= not a or b;
    layer2_outputs(7312) <= '1';
    layer2_outputs(7313) <= '1';
    layer2_outputs(7314) <= a and b;
    layer2_outputs(7315) <= a and b;
    layer2_outputs(7316) <= a and b;
    layer2_outputs(7317) <= b;
    layer2_outputs(7318) <= not b;
    layer2_outputs(7319) <= '1';
    layer2_outputs(7320) <= a;
    layer2_outputs(7321) <= not a;
    layer2_outputs(7322) <= '0';
    layer2_outputs(7323) <= not b;
    layer2_outputs(7324) <= not a or b;
    layer2_outputs(7325) <= a and b;
    layer2_outputs(7326) <= a or b;
    layer2_outputs(7327) <= a xor b;
    layer2_outputs(7328) <= '0';
    layer2_outputs(7329) <= not a;
    layer2_outputs(7330) <= not b or a;
    layer2_outputs(7331) <= a and b;
    layer2_outputs(7332) <= a;
    layer2_outputs(7333) <= '0';
    layer2_outputs(7334) <= not a or b;
    layer2_outputs(7335) <= not b or a;
    layer2_outputs(7336) <= b;
    layer2_outputs(7337) <= not b or a;
    layer2_outputs(7338) <= not a;
    layer2_outputs(7339) <= a and not b;
    layer2_outputs(7340) <= not b;
    layer2_outputs(7341) <= b and not a;
    layer2_outputs(7342) <= not b or a;
    layer2_outputs(7343) <= b;
    layer2_outputs(7344) <= b and not a;
    layer2_outputs(7345) <= not b or a;
    layer2_outputs(7346) <= b and not a;
    layer2_outputs(7347) <= a and not b;
    layer2_outputs(7348) <= not a;
    layer2_outputs(7349) <= a or b;
    layer2_outputs(7350) <= not a or b;
    layer2_outputs(7351) <= b;
    layer2_outputs(7352) <= not a or b;
    layer2_outputs(7353) <= '0';
    layer2_outputs(7354) <= a;
    layer2_outputs(7355) <= a;
    layer2_outputs(7356) <= not b;
    layer2_outputs(7357) <= a or b;
    layer2_outputs(7358) <= not b or a;
    layer2_outputs(7359) <= '1';
    layer2_outputs(7360) <= b and not a;
    layer2_outputs(7361) <= '0';
    layer2_outputs(7362) <= not b or a;
    layer2_outputs(7363) <= not a or b;
    layer2_outputs(7364) <= '1';
    layer2_outputs(7365) <= '1';
    layer2_outputs(7366) <= a and not b;
    layer2_outputs(7367) <= '0';
    layer2_outputs(7368) <= not b or a;
    layer2_outputs(7369) <= a or b;
    layer2_outputs(7370) <= a and not b;
    layer2_outputs(7371) <= not (a or b);
    layer2_outputs(7372) <= a or b;
    layer2_outputs(7373) <= '1';
    layer2_outputs(7374) <= b;
    layer2_outputs(7375) <= a;
    layer2_outputs(7376) <= not b or a;
    layer2_outputs(7377) <= not (a or b);
    layer2_outputs(7378) <= a;
    layer2_outputs(7379) <= not (a and b);
    layer2_outputs(7380) <= a xor b;
    layer2_outputs(7381) <= not b or a;
    layer2_outputs(7382) <= b and not a;
    layer2_outputs(7383) <= not (a or b);
    layer2_outputs(7384) <= not b or a;
    layer2_outputs(7385) <= not a or b;
    layer2_outputs(7386) <= not a or b;
    layer2_outputs(7387) <= a;
    layer2_outputs(7388) <= not b;
    layer2_outputs(7389) <= '0';
    layer2_outputs(7390) <= '0';
    layer2_outputs(7391) <= '0';
    layer2_outputs(7392) <= not b or a;
    layer2_outputs(7393) <= '0';
    layer2_outputs(7394) <= '0';
    layer2_outputs(7395) <= not a or b;
    layer2_outputs(7396) <= not (a or b);
    layer2_outputs(7397) <= a and not b;
    layer2_outputs(7398) <= a xor b;
    layer2_outputs(7399) <= not a or b;
    layer2_outputs(7400) <= not a;
    layer2_outputs(7401) <= '1';
    layer2_outputs(7402) <= not (a and b);
    layer2_outputs(7403) <= not a or b;
    layer2_outputs(7404) <= a and not b;
    layer2_outputs(7405) <= b;
    layer2_outputs(7406) <= '0';
    layer2_outputs(7407) <= b;
    layer2_outputs(7408) <= not b;
    layer2_outputs(7409) <= a;
    layer2_outputs(7410) <= not (a and b);
    layer2_outputs(7411) <= b and not a;
    layer2_outputs(7412) <= not a;
    layer2_outputs(7413) <= not a or b;
    layer2_outputs(7414) <= a;
    layer2_outputs(7415) <= not a or b;
    layer2_outputs(7416) <= not a or b;
    layer2_outputs(7417) <= a;
    layer2_outputs(7418) <= '1';
    layer2_outputs(7419) <= b and not a;
    layer2_outputs(7420) <= '0';
    layer2_outputs(7421) <= a or b;
    layer2_outputs(7422) <= a or b;
    layer2_outputs(7423) <= '1';
    layer2_outputs(7424) <= a and b;
    layer2_outputs(7425) <= not b or a;
    layer2_outputs(7426) <= not (a and b);
    layer2_outputs(7427) <= not a;
    layer2_outputs(7428) <= not a;
    layer2_outputs(7429) <= '0';
    layer2_outputs(7430) <= a and not b;
    layer2_outputs(7431) <= '1';
    layer2_outputs(7432) <= a and not b;
    layer2_outputs(7433) <= not (a or b);
    layer2_outputs(7434) <= not a;
    layer2_outputs(7435) <= b;
    layer2_outputs(7436) <= '0';
    layer2_outputs(7437) <= not (a or b);
    layer2_outputs(7438) <= not a;
    layer2_outputs(7439) <= '1';
    layer2_outputs(7440) <= b;
    layer2_outputs(7441) <= not (a and b);
    layer2_outputs(7442) <= '1';
    layer2_outputs(7443) <= not (a or b);
    layer2_outputs(7444) <= not (a and b);
    layer2_outputs(7445) <= not a;
    layer2_outputs(7446) <= '0';
    layer2_outputs(7447) <= a xor b;
    layer2_outputs(7448) <= not (a or b);
    layer2_outputs(7449) <= not (a and b);
    layer2_outputs(7450) <= b and not a;
    layer2_outputs(7451) <= a;
    layer2_outputs(7452) <= not b or a;
    layer2_outputs(7453) <= not b;
    layer2_outputs(7454) <= a and b;
    layer2_outputs(7455) <= not b or a;
    layer2_outputs(7456) <= not a;
    layer2_outputs(7457) <= not (a or b);
    layer2_outputs(7458) <= not a or b;
    layer2_outputs(7459) <= b and not a;
    layer2_outputs(7460) <= a and not b;
    layer2_outputs(7461) <= b and not a;
    layer2_outputs(7462) <= not (a xor b);
    layer2_outputs(7463) <= not b;
    layer2_outputs(7464) <= a and not b;
    layer2_outputs(7465) <= a;
    layer2_outputs(7466) <= not (a or b);
    layer2_outputs(7467) <= '0';
    layer2_outputs(7468) <= b and not a;
    layer2_outputs(7469) <= a and b;
    layer2_outputs(7470) <= not a;
    layer2_outputs(7471) <= b;
    layer2_outputs(7472) <= not b;
    layer2_outputs(7473) <= not (a and b);
    layer2_outputs(7474) <= b;
    layer2_outputs(7475) <= a and b;
    layer2_outputs(7476) <= a or b;
    layer2_outputs(7477) <= a and not b;
    layer2_outputs(7478) <= a xor b;
    layer2_outputs(7479) <= not (a or b);
    layer2_outputs(7480) <= a or b;
    layer2_outputs(7481) <= a or b;
    layer2_outputs(7482) <= not b;
    layer2_outputs(7483) <= a xor b;
    layer2_outputs(7484) <= a and b;
    layer2_outputs(7485) <= '1';
    layer2_outputs(7486) <= '0';
    layer2_outputs(7487) <= '0';
    layer2_outputs(7488) <= a and not b;
    layer2_outputs(7489) <= a or b;
    layer2_outputs(7490) <= a;
    layer2_outputs(7491) <= a and b;
    layer2_outputs(7492) <= not b;
    layer2_outputs(7493) <= not (a xor b);
    layer2_outputs(7494) <= not b or a;
    layer2_outputs(7495) <= not (a and b);
    layer2_outputs(7496) <= not (a or b);
    layer2_outputs(7497) <= a and b;
    layer2_outputs(7498) <= b and not a;
    layer2_outputs(7499) <= b;
    layer2_outputs(7500) <= a or b;
    layer2_outputs(7501) <= not (a xor b);
    layer2_outputs(7502) <= not a or b;
    layer2_outputs(7503) <= not (a and b);
    layer2_outputs(7504) <= not a;
    layer2_outputs(7505) <= a and b;
    layer2_outputs(7506) <= '0';
    layer2_outputs(7507) <= a xor b;
    layer2_outputs(7508) <= a or b;
    layer2_outputs(7509) <= a and b;
    layer2_outputs(7510) <= not b or a;
    layer2_outputs(7511) <= '0';
    layer2_outputs(7512) <= a;
    layer2_outputs(7513) <= not (a or b);
    layer2_outputs(7514) <= not a;
    layer2_outputs(7515) <= not (a or b);
    layer2_outputs(7516) <= a and b;
    layer2_outputs(7517) <= b and not a;
    layer2_outputs(7518) <= a and b;
    layer2_outputs(7519) <= not a or b;
    layer2_outputs(7520) <= a or b;
    layer2_outputs(7521) <= a and b;
    layer2_outputs(7522) <= not a;
    layer2_outputs(7523) <= '1';
    layer2_outputs(7524) <= not b or a;
    layer2_outputs(7525) <= not b;
    layer2_outputs(7526) <= b and not a;
    layer2_outputs(7527) <= a and b;
    layer2_outputs(7528) <= a;
    layer2_outputs(7529) <= a;
    layer2_outputs(7530) <= a;
    layer2_outputs(7531) <= not b;
    layer2_outputs(7532) <= not b or a;
    layer2_outputs(7533) <= '1';
    layer2_outputs(7534) <= not (a or b);
    layer2_outputs(7535) <= not a or b;
    layer2_outputs(7536) <= '1';
    layer2_outputs(7537) <= a or b;
    layer2_outputs(7538) <= not (a and b);
    layer2_outputs(7539) <= '0';
    layer2_outputs(7540) <= not a or b;
    layer2_outputs(7541) <= not b;
    layer2_outputs(7542) <= not b or a;
    layer2_outputs(7543) <= b and not a;
    layer2_outputs(7544) <= a xor b;
    layer2_outputs(7545) <= a and not b;
    layer2_outputs(7546) <= not (a or b);
    layer2_outputs(7547) <= a and b;
    layer2_outputs(7548) <= '0';
    layer2_outputs(7549) <= '0';
    layer2_outputs(7550) <= not a;
    layer2_outputs(7551) <= a and b;
    layer2_outputs(7552) <= not (a xor b);
    layer2_outputs(7553) <= not a or b;
    layer2_outputs(7554) <= a;
    layer2_outputs(7555) <= not a;
    layer2_outputs(7556) <= a and not b;
    layer2_outputs(7557) <= a and b;
    layer2_outputs(7558) <= not (a and b);
    layer2_outputs(7559) <= a and b;
    layer2_outputs(7560) <= not (a and b);
    layer2_outputs(7561) <= b and not a;
    layer2_outputs(7562) <= '0';
    layer2_outputs(7563) <= not (a and b);
    layer2_outputs(7564) <= b;
    layer2_outputs(7565) <= b;
    layer2_outputs(7566) <= not (a or b);
    layer2_outputs(7567) <= a and not b;
    layer2_outputs(7568) <= '0';
    layer2_outputs(7569) <= '1';
    layer2_outputs(7570) <= a or b;
    layer2_outputs(7571) <= b and not a;
    layer2_outputs(7572) <= not (a and b);
    layer2_outputs(7573) <= '1';
    layer2_outputs(7574) <= not b or a;
    layer2_outputs(7575) <= not a;
    layer2_outputs(7576) <= not (a and b);
    layer2_outputs(7577) <= not (a xor b);
    layer2_outputs(7578) <= not b;
    layer2_outputs(7579) <= not (a or b);
    layer2_outputs(7580) <= a or b;
    layer2_outputs(7581) <= not (a or b);
    layer2_outputs(7582) <= a;
    layer2_outputs(7583) <= '1';
    layer2_outputs(7584) <= a;
    layer2_outputs(7585) <= not b or a;
    layer2_outputs(7586) <= '0';
    layer2_outputs(7587) <= not (a or b);
    layer2_outputs(7588) <= a;
    layer2_outputs(7589) <= b and not a;
    layer2_outputs(7590) <= a and b;
    layer2_outputs(7591) <= b;
    layer2_outputs(7592) <= not a or b;
    layer2_outputs(7593) <= '1';
    layer2_outputs(7594) <= a or b;
    layer2_outputs(7595) <= '1';
    layer2_outputs(7596) <= '1';
    layer2_outputs(7597) <= a and b;
    layer2_outputs(7598) <= not (a and b);
    layer2_outputs(7599) <= not (a and b);
    layer2_outputs(7600) <= b and not a;
    layer2_outputs(7601) <= not (a or b);
    layer2_outputs(7602) <= a;
    layer2_outputs(7603) <= not (a or b);
    layer2_outputs(7604) <= '0';
    layer2_outputs(7605) <= not b or a;
    layer2_outputs(7606) <= b and not a;
    layer2_outputs(7607) <= a;
    layer2_outputs(7608) <= a and not b;
    layer2_outputs(7609) <= a or b;
    layer2_outputs(7610) <= a or b;
    layer2_outputs(7611) <= not a;
    layer2_outputs(7612) <= '0';
    layer2_outputs(7613) <= a and not b;
    layer2_outputs(7614) <= not a;
    layer2_outputs(7615) <= b;
    layer2_outputs(7616) <= '1';
    layer2_outputs(7617) <= not (a and b);
    layer2_outputs(7618) <= not (a or b);
    layer2_outputs(7619) <= not (a or b);
    layer2_outputs(7620) <= a and not b;
    layer2_outputs(7621) <= '1';
    layer2_outputs(7622) <= '1';
    layer2_outputs(7623) <= '0';
    layer2_outputs(7624) <= '0';
    layer2_outputs(7625) <= '0';
    layer2_outputs(7626) <= a or b;
    layer2_outputs(7627) <= '1';
    layer2_outputs(7628) <= not a or b;
    layer2_outputs(7629) <= not a;
    layer2_outputs(7630) <= not (a or b);
    layer2_outputs(7631) <= b;
    layer2_outputs(7632) <= b and not a;
    layer2_outputs(7633) <= '0';
    layer2_outputs(7634) <= '1';
    layer2_outputs(7635) <= b;
    layer2_outputs(7636) <= a and not b;
    layer2_outputs(7637) <= b and not a;
    layer2_outputs(7638) <= not a or b;
    layer2_outputs(7639) <= not (a and b);
    layer2_outputs(7640) <= not (a and b);
    layer2_outputs(7641) <= '1';
    layer2_outputs(7642) <= a or b;
    layer2_outputs(7643) <= not a;
    layer2_outputs(7644) <= not (a or b);
    layer2_outputs(7645) <= '1';
    layer2_outputs(7646) <= not b or a;
    layer2_outputs(7647) <= not a;
    layer2_outputs(7648) <= '0';
    layer2_outputs(7649) <= a and b;
    layer2_outputs(7650) <= '1';
    layer2_outputs(7651) <= not (a and b);
    layer2_outputs(7652) <= not (a and b);
    layer2_outputs(7653) <= a and b;
    layer2_outputs(7654) <= not a;
    layer2_outputs(7655) <= not b;
    layer2_outputs(7656) <= a;
    layer2_outputs(7657) <= not (a and b);
    layer2_outputs(7658) <= not (a and b);
    layer2_outputs(7659) <= not (a and b);
    layer2_outputs(7660) <= not b or a;
    layer2_outputs(7661) <= b;
    layer2_outputs(7662) <= not a;
    layer2_outputs(7663) <= '0';
    layer2_outputs(7664) <= not b or a;
    layer2_outputs(7665) <= '0';
    layer2_outputs(7666) <= a and b;
    layer2_outputs(7667) <= '0';
    layer2_outputs(7668) <= not (a or b);
    layer2_outputs(7669) <= '1';
    layer2_outputs(7670) <= '1';
    layer2_outputs(7671) <= '1';
    layer2_outputs(7672) <= b;
    layer2_outputs(7673) <= a and not b;
    layer2_outputs(7674) <= a and not b;
    layer2_outputs(7675) <= not (a or b);
    layer2_outputs(7676) <= a and not b;
    layer2_outputs(7677) <= a xor b;
    layer2_outputs(7678) <= '1';
    layer2_outputs(7679) <= not a;
    layer3_outputs(0) <= a and not b;
    layer3_outputs(1) <= not (a xor b);
    layer3_outputs(2) <= not b;
    layer3_outputs(3) <= a or b;
    layer3_outputs(4) <= a and not b;
    layer3_outputs(5) <= a and b;
    layer3_outputs(6) <= not a;
    layer3_outputs(7) <= a and not b;
    layer3_outputs(8) <= '1';
    layer3_outputs(9) <= not b;
    layer3_outputs(10) <= not a;
    layer3_outputs(11) <= a and b;
    layer3_outputs(12) <= '1';
    layer3_outputs(13) <= not b or a;
    layer3_outputs(14) <= b and not a;
    layer3_outputs(15) <= '1';
    layer3_outputs(16) <= not a;
    layer3_outputs(17) <= a;
    layer3_outputs(18) <= not b;
    layer3_outputs(19) <= a;
    layer3_outputs(20) <= not (a and b);
    layer3_outputs(21) <= not (a or b);
    layer3_outputs(22) <= not b;
    layer3_outputs(23) <= not a;
    layer3_outputs(24) <= '0';
    layer3_outputs(25) <= not (a or b);
    layer3_outputs(26) <= a xor b;
    layer3_outputs(27) <= a xor b;
    layer3_outputs(28) <= a;
    layer3_outputs(29) <= not b or a;
    layer3_outputs(30) <= not a;
    layer3_outputs(31) <= not (a or b);
    layer3_outputs(32) <= not b or a;
    layer3_outputs(33) <= '0';
    layer3_outputs(34) <= not a or b;
    layer3_outputs(35) <= a and not b;
    layer3_outputs(36) <= b;
    layer3_outputs(37) <= not b;
    layer3_outputs(38) <= a xor b;
    layer3_outputs(39) <= not b or a;
    layer3_outputs(40) <= a and b;
    layer3_outputs(41) <= b;
    layer3_outputs(42) <= not (a and b);
    layer3_outputs(43) <= not b;
    layer3_outputs(44) <= a or b;
    layer3_outputs(45) <= not b or a;
    layer3_outputs(46) <= not a or b;
    layer3_outputs(47) <= not a or b;
    layer3_outputs(48) <= a and b;
    layer3_outputs(49) <= a and not b;
    layer3_outputs(50) <= not b or a;
    layer3_outputs(51) <= a and not b;
    layer3_outputs(52) <= '0';
    layer3_outputs(53) <= a and b;
    layer3_outputs(54) <= not (a xor b);
    layer3_outputs(55) <= a and b;
    layer3_outputs(56) <= a and not b;
    layer3_outputs(57) <= not (a xor b);
    layer3_outputs(58) <= a;
    layer3_outputs(59) <= not a or b;
    layer3_outputs(60) <= not (a or b);
    layer3_outputs(61) <= a and not b;
    layer3_outputs(62) <= not b or a;
    layer3_outputs(63) <= not a;
    layer3_outputs(64) <= b and not a;
    layer3_outputs(65) <= not (a xor b);
    layer3_outputs(66) <= b;
    layer3_outputs(67) <= not b or a;
    layer3_outputs(68) <= not a;
    layer3_outputs(69) <= not a;
    layer3_outputs(70) <= not (a or b);
    layer3_outputs(71) <= not a;
    layer3_outputs(72) <= b and not a;
    layer3_outputs(73) <= a and b;
    layer3_outputs(74) <= not b;
    layer3_outputs(75) <= '1';
    layer3_outputs(76) <= b and not a;
    layer3_outputs(77) <= a and b;
    layer3_outputs(78) <= b;
    layer3_outputs(79) <= not a;
    layer3_outputs(80) <= not a or b;
    layer3_outputs(81) <= a and not b;
    layer3_outputs(82) <= not (a or b);
    layer3_outputs(83) <= '0';
    layer3_outputs(84) <= not b;
    layer3_outputs(85) <= b;
    layer3_outputs(86) <= b and not a;
    layer3_outputs(87) <= b;
    layer3_outputs(88) <= a;
    layer3_outputs(89) <= '1';
    layer3_outputs(90) <= not (a or b);
    layer3_outputs(91) <= not a or b;
    layer3_outputs(92) <= not b;
    layer3_outputs(93) <= not a or b;
    layer3_outputs(94) <= not a or b;
    layer3_outputs(95) <= not (a and b);
    layer3_outputs(96) <= not a;
    layer3_outputs(97) <= not a;
    layer3_outputs(98) <= b;
    layer3_outputs(99) <= '0';
    layer3_outputs(100) <= b and not a;
    layer3_outputs(101) <= a and b;
    layer3_outputs(102) <= a and not b;
    layer3_outputs(103) <= not a;
    layer3_outputs(104) <= not (a xor b);
    layer3_outputs(105) <= not a or b;
    layer3_outputs(106) <= not (a or b);
    layer3_outputs(107) <= not (a or b);
    layer3_outputs(108) <= a;
    layer3_outputs(109) <= a and not b;
    layer3_outputs(110) <= not (a xor b);
    layer3_outputs(111) <= not a or b;
    layer3_outputs(112) <= '1';
    layer3_outputs(113) <= not (a xor b);
    layer3_outputs(114) <= a xor b;
    layer3_outputs(115) <= a xor b;
    layer3_outputs(116) <= a and b;
    layer3_outputs(117) <= not a or b;
    layer3_outputs(118) <= not b or a;
    layer3_outputs(119) <= not b;
    layer3_outputs(120) <= a and not b;
    layer3_outputs(121) <= not (a and b);
    layer3_outputs(122) <= not b;
    layer3_outputs(123) <= '1';
    layer3_outputs(124) <= not b;
    layer3_outputs(125) <= a and not b;
    layer3_outputs(126) <= a xor b;
    layer3_outputs(127) <= a;
    layer3_outputs(128) <= not (a and b);
    layer3_outputs(129) <= a and not b;
    layer3_outputs(130) <= a or b;
    layer3_outputs(131) <= not b or a;
    layer3_outputs(132) <= not (a xor b);
    layer3_outputs(133) <= not (a and b);
    layer3_outputs(134) <= not b or a;
    layer3_outputs(135) <= not a;
    layer3_outputs(136) <= '0';
    layer3_outputs(137) <= b;
    layer3_outputs(138) <= not a;
    layer3_outputs(139) <= b and not a;
    layer3_outputs(140) <= b and not a;
    layer3_outputs(141) <= '1';
    layer3_outputs(142) <= b and not a;
    layer3_outputs(143) <= not a or b;
    layer3_outputs(144) <= b;
    layer3_outputs(145) <= b;
    layer3_outputs(146) <= not (a or b);
    layer3_outputs(147) <= not (a and b);
    layer3_outputs(148) <= a and b;
    layer3_outputs(149) <= a xor b;
    layer3_outputs(150) <= not (a and b);
    layer3_outputs(151) <= not a or b;
    layer3_outputs(152) <= a;
    layer3_outputs(153) <= not a;
    layer3_outputs(154) <= b;
    layer3_outputs(155) <= '0';
    layer3_outputs(156) <= not b;
    layer3_outputs(157) <= a;
    layer3_outputs(158) <= a;
    layer3_outputs(159) <= b and not a;
    layer3_outputs(160) <= not b or a;
    layer3_outputs(161) <= a;
    layer3_outputs(162) <= '0';
    layer3_outputs(163) <= a;
    layer3_outputs(164) <= '0';
    layer3_outputs(165) <= a and b;
    layer3_outputs(166) <= '1';
    layer3_outputs(167) <= not a;
    layer3_outputs(168) <= a and not b;
    layer3_outputs(169) <= not a or b;
    layer3_outputs(170) <= not a;
    layer3_outputs(171) <= not a;
    layer3_outputs(172) <= a or b;
    layer3_outputs(173) <= a or b;
    layer3_outputs(174) <= a and b;
    layer3_outputs(175) <= b;
    layer3_outputs(176) <= '1';
    layer3_outputs(177) <= '0';
    layer3_outputs(178) <= b;
    layer3_outputs(179) <= not b or a;
    layer3_outputs(180) <= not (a or b);
    layer3_outputs(181) <= not a;
    layer3_outputs(182) <= not (a and b);
    layer3_outputs(183) <= '0';
    layer3_outputs(184) <= not (a or b);
    layer3_outputs(185) <= b;
    layer3_outputs(186) <= a;
    layer3_outputs(187) <= not a or b;
    layer3_outputs(188) <= not (a and b);
    layer3_outputs(189) <= not a;
    layer3_outputs(190) <= b;
    layer3_outputs(191) <= b and not a;
    layer3_outputs(192) <= not a;
    layer3_outputs(193) <= b and not a;
    layer3_outputs(194) <= a and not b;
    layer3_outputs(195) <= not b or a;
    layer3_outputs(196) <= b and not a;
    layer3_outputs(197) <= '0';
    layer3_outputs(198) <= not a;
    layer3_outputs(199) <= a or b;
    layer3_outputs(200) <= a and b;
    layer3_outputs(201) <= b and not a;
    layer3_outputs(202) <= not a;
    layer3_outputs(203) <= a and not b;
    layer3_outputs(204) <= '1';
    layer3_outputs(205) <= not a or b;
    layer3_outputs(206) <= b;
    layer3_outputs(207) <= not a;
    layer3_outputs(208) <= '0';
    layer3_outputs(209) <= '0';
    layer3_outputs(210) <= a and not b;
    layer3_outputs(211) <= not a;
    layer3_outputs(212) <= not (a or b);
    layer3_outputs(213) <= not a;
    layer3_outputs(214) <= '1';
    layer3_outputs(215) <= not a;
    layer3_outputs(216) <= not (a or b);
    layer3_outputs(217) <= '0';
    layer3_outputs(218) <= not a or b;
    layer3_outputs(219) <= not b;
    layer3_outputs(220) <= a or b;
    layer3_outputs(221) <= not a;
    layer3_outputs(222) <= not (a xor b);
    layer3_outputs(223) <= a and b;
    layer3_outputs(224) <= a and not b;
    layer3_outputs(225) <= '1';
    layer3_outputs(226) <= not b or a;
    layer3_outputs(227) <= b and not a;
    layer3_outputs(228) <= not (a or b);
    layer3_outputs(229) <= not a or b;
    layer3_outputs(230) <= b and not a;
    layer3_outputs(231) <= not (a xor b);
    layer3_outputs(232) <= not (a and b);
    layer3_outputs(233) <= a and b;
    layer3_outputs(234) <= not (a and b);
    layer3_outputs(235) <= not a;
    layer3_outputs(236) <= b and not a;
    layer3_outputs(237) <= b and not a;
    layer3_outputs(238) <= b;
    layer3_outputs(239) <= a and not b;
    layer3_outputs(240) <= b and not a;
    layer3_outputs(241) <= b and not a;
    layer3_outputs(242) <= not b;
    layer3_outputs(243) <= b and not a;
    layer3_outputs(244) <= a and b;
    layer3_outputs(245) <= a and b;
    layer3_outputs(246) <= not a;
    layer3_outputs(247) <= not b or a;
    layer3_outputs(248) <= not (a xor b);
    layer3_outputs(249) <= a and not b;
    layer3_outputs(250) <= not b or a;
    layer3_outputs(251) <= not b;
    layer3_outputs(252) <= not (a and b);
    layer3_outputs(253) <= a and not b;
    layer3_outputs(254) <= not a;
    layer3_outputs(255) <= '0';
    layer3_outputs(256) <= not b;
    layer3_outputs(257) <= not a or b;
    layer3_outputs(258) <= a and b;
    layer3_outputs(259) <= not b or a;
    layer3_outputs(260) <= a and b;
    layer3_outputs(261) <= a and not b;
    layer3_outputs(262) <= '0';
    layer3_outputs(263) <= '1';
    layer3_outputs(264) <= not b or a;
    layer3_outputs(265) <= not b or a;
    layer3_outputs(266) <= not a;
    layer3_outputs(267) <= not a;
    layer3_outputs(268) <= a or b;
    layer3_outputs(269) <= b and not a;
    layer3_outputs(270) <= not b or a;
    layer3_outputs(271) <= not a;
    layer3_outputs(272) <= a or b;
    layer3_outputs(273) <= a;
    layer3_outputs(274) <= a and not b;
    layer3_outputs(275) <= not (a and b);
    layer3_outputs(276) <= not b or a;
    layer3_outputs(277) <= not (a and b);
    layer3_outputs(278) <= not (a and b);
    layer3_outputs(279) <= a;
    layer3_outputs(280) <= a and not b;
    layer3_outputs(281) <= '0';
    layer3_outputs(282) <= b;
    layer3_outputs(283) <= a xor b;
    layer3_outputs(284) <= b and not a;
    layer3_outputs(285) <= not (a and b);
    layer3_outputs(286) <= a and not b;
    layer3_outputs(287) <= a or b;
    layer3_outputs(288) <= b;
    layer3_outputs(289) <= not (a or b);
    layer3_outputs(290) <= not a;
    layer3_outputs(291) <= not (a or b);
    layer3_outputs(292) <= b and not a;
    layer3_outputs(293) <= a and b;
    layer3_outputs(294) <= not b;
    layer3_outputs(295) <= a;
    layer3_outputs(296) <= not b or a;
    layer3_outputs(297) <= '1';
    layer3_outputs(298) <= not (a and b);
    layer3_outputs(299) <= not b;
    layer3_outputs(300) <= not (a or b);
    layer3_outputs(301) <= '0';
    layer3_outputs(302) <= '0';
    layer3_outputs(303) <= not a;
    layer3_outputs(304) <= '1';
    layer3_outputs(305) <= not a;
    layer3_outputs(306) <= not b or a;
    layer3_outputs(307) <= not (a or b);
    layer3_outputs(308) <= not a or b;
    layer3_outputs(309) <= '0';
    layer3_outputs(310) <= not (a and b);
    layer3_outputs(311) <= b;
    layer3_outputs(312) <= a and b;
    layer3_outputs(313) <= b and not a;
    layer3_outputs(314) <= not b;
    layer3_outputs(315) <= not b or a;
    layer3_outputs(316) <= not b;
    layer3_outputs(317) <= a and b;
    layer3_outputs(318) <= a;
    layer3_outputs(319) <= not b or a;
    layer3_outputs(320) <= not (a or b);
    layer3_outputs(321) <= not a or b;
    layer3_outputs(322) <= not a;
    layer3_outputs(323) <= not (a and b);
    layer3_outputs(324) <= a xor b;
    layer3_outputs(325) <= not (a or b);
    layer3_outputs(326) <= not a or b;
    layer3_outputs(327) <= a or b;
    layer3_outputs(328) <= a;
    layer3_outputs(329) <= b;
    layer3_outputs(330) <= a;
    layer3_outputs(331) <= not a or b;
    layer3_outputs(332) <= a;
    layer3_outputs(333) <= not a or b;
    layer3_outputs(334) <= not a;
    layer3_outputs(335) <= a and b;
    layer3_outputs(336) <= a and b;
    layer3_outputs(337) <= not (a or b);
    layer3_outputs(338) <= not b;
    layer3_outputs(339) <= '1';
    layer3_outputs(340) <= b and not a;
    layer3_outputs(341) <= '1';
    layer3_outputs(342) <= not b;
    layer3_outputs(343) <= a or b;
    layer3_outputs(344) <= not a or b;
    layer3_outputs(345) <= a and b;
    layer3_outputs(346) <= a;
    layer3_outputs(347) <= not (a or b);
    layer3_outputs(348) <= a or b;
    layer3_outputs(349) <= a and b;
    layer3_outputs(350) <= not a or b;
    layer3_outputs(351) <= a or b;
    layer3_outputs(352) <= not a or b;
    layer3_outputs(353) <= a and b;
    layer3_outputs(354) <= b and not a;
    layer3_outputs(355) <= not (a or b);
    layer3_outputs(356) <= b and not a;
    layer3_outputs(357) <= not b or a;
    layer3_outputs(358) <= a;
    layer3_outputs(359) <= not a;
    layer3_outputs(360) <= not b or a;
    layer3_outputs(361) <= not b;
    layer3_outputs(362) <= not (a or b);
    layer3_outputs(363) <= a;
    layer3_outputs(364) <= not b or a;
    layer3_outputs(365) <= a xor b;
    layer3_outputs(366) <= '1';
    layer3_outputs(367) <= not (a or b);
    layer3_outputs(368) <= not b;
    layer3_outputs(369) <= not a or b;
    layer3_outputs(370) <= a and not b;
    layer3_outputs(371) <= b;
    layer3_outputs(372) <= a;
    layer3_outputs(373) <= a xor b;
    layer3_outputs(374) <= '0';
    layer3_outputs(375) <= a xor b;
    layer3_outputs(376) <= b and not a;
    layer3_outputs(377) <= not b;
    layer3_outputs(378) <= a and not b;
    layer3_outputs(379) <= not b or a;
    layer3_outputs(380) <= a;
    layer3_outputs(381) <= not b;
    layer3_outputs(382) <= a and b;
    layer3_outputs(383) <= a and not b;
    layer3_outputs(384) <= a or b;
    layer3_outputs(385) <= a and b;
    layer3_outputs(386) <= b and not a;
    layer3_outputs(387) <= '0';
    layer3_outputs(388) <= b;
    layer3_outputs(389) <= a and not b;
    layer3_outputs(390) <= '0';
    layer3_outputs(391) <= a or b;
    layer3_outputs(392) <= '1';
    layer3_outputs(393) <= b and not a;
    layer3_outputs(394) <= a or b;
    layer3_outputs(395) <= b;
    layer3_outputs(396) <= a xor b;
    layer3_outputs(397) <= not (a and b);
    layer3_outputs(398) <= a and b;
    layer3_outputs(399) <= not b;
    layer3_outputs(400) <= not b;
    layer3_outputs(401) <= a;
    layer3_outputs(402) <= a and b;
    layer3_outputs(403) <= not a;
    layer3_outputs(404) <= b;
    layer3_outputs(405) <= a or b;
    layer3_outputs(406) <= a or b;
    layer3_outputs(407) <= b;
    layer3_outputs(408) <= not a;
    layer3_outputs(409) <= a and b;
    layer3_outputs(410) <= b;
    layer3_outputs(411) <= a or b;
    layer3_outputs(412) <= not (a or b);
    layer3_outputs(413) <= '0';
    layer3_outputs(414) <= a;
    layer3_outputs(415) <= not b or a;
    layer3_outputs(416) <= '0';
    layer3_outputs(417) <= not (a or b);
    layer3_outputs(418) <= not (a and b);
    layer3_outputs(419) <= not a;
    layer3_outputs(420) <= not (a and b);
    layer3_outputs(421) <= '0';
    layer3_outputs(422) <= not b or a;
    layer3_outputs(423) <= b and not a;
    layer3_outputs(424) <= not a;
    layer3_outputs(425) <= not (a or b);
    layer3_outputs(426) <= not (a or b);
    layer3_outputs(427) <= b;
    layer3_outputs(428) <= not a or b;
    layer3_outputs(429) <= a;
    layer3_outputs(430) <= b and not a;
    layer3_outputs(431) <= a and not b;
    layer3_outputs(432) <= not (a and b);
    layer3_outputs(433) <= a and b;
    layer3_outputs(434) <= a and not b;
    layer3_outputs(435) <= not b or a;
    layer3_outputs(436) <= b and not a;
    layer3_outputs(437) <= not a or b;
    layer3_outputs(438) <= b;
    layer3_outputs(439) <= a and not b;
    layer3_outputs(440) <= '0';
    layer3_outputs(441) <= not (a or b);
    layer3_outputs(442) <= not (a and b);
    layer3_outputs(443) <= a and not b;
    layer3_outputs(444) <= b;
    layer3_outputs(445) <= a;
    layer3_outputs(446) <= a;
    layer3_outputs(447) <= b;
    layer3_outputs(448) <= not (a xor b);
    layer3_outputs(449) <= a and b;
    layer3_outputs(450) <= not b or a;
    layer3_outputs(451) <= a or b;
    layer3_outputs(452) <= not a or b;
    layer3_outputs(453) <= '1';
    layer3_outputs(454) <= '0';
    layer3_outputs(455) <= not b or a;
    layer3_outputs(456) <= b and not a;
    layer3_outputs(457) <= a or b;
    layer3_outputs(458) <= b;
    layer3_outputs(459) <= '1';
    layer3_outputs(460) <= not (a or b);
    layer3_outputs(461) <= not a or b;
    layer3_outputs(462) <= not (a xor b);
    layer3_outputs(463) <= a and not b;
    layer3_outputs(464) <= not (a or b);
    layer3_outputs(465) <= not a or b;
    layer3_outputs(466) <= b;
    layer3_outputs(467) <= not b;
    layer3_outputs(468) <= not a;
    layer3_outputs(469) <= not (a or b);
    layer3_outputs(470) <= '1';
    layer3_outputs(471) <= a or b;
    layer3_outputs(472) <= a and b;
    layer3_outputs(473) <= b;
    layer3_outputs(474) <= not a;
    layer3_outputs(475) <= '0';
    layer3_outputs(476) <= a and b;
    layer3_outputs(477) <= b and not a;
    layer3_outputs(478) <= a;
    layer3_outputs(479) <= a or b;
    layer3_outputs(480) <= '0';
    layer3_outputs(481) <= not a;
    layer3_outputs(482) <= a xor b;
    layer3_outputs(483) <= not a or b;
    layer3_outputs(484) <= not (a or b);
    layer3_outputs(485) <= not b or a;
    layer3_outputs(486) <= not b or a;
    layer3_outputs(487) <= b and not a;
    layer3_outputs(488) <= b;
    layer3_outputs(489) <= a and not b;
    layer3_outputs(490) <= a and b;
    layer3_outputs(491) <= '1';
    layer3_outputs(492) <= not b or a;
    layer3_outputs(493) <= not b;
    layer3_outputs(494) <= not (a or b);
    layer3_outputs(495) <= not b or a;
    layer3_outputs(496) <= not b or a;
    layer3_outputs(497) <= not b or a;
    layer3_outputs(498) <= b and not a;
    layer3_outputs(499) <= not b;
    layer3_outputs(500) <= '1';
    layer3_outputs(501) <= a and b;
    layer3_outputs(502) <= a and b;
    layer3_outputs(503) <= '0';
    layer3_outputs(504) <= not a;
    layer3_outputs(505) <= not b or a;
    layer3_outputs(506) <= '0';
    layer3_outputs(507) <= '1';
    layer3_outputs(508) <= a and b;
    layer3_outputs(509) <= not a;
    layer3_outputs(510) <= not (a or b);
    layer3_outputs(511) <= b;
    layer3_outputs(512) <= b;
    layer3_outputs(513) <= a;
    layer3_outputs(514) <= not b or a;
    layer3_outputs(515) <= a or b;
    layer3_outputs(516) <= '1';
    layer3_outputs(517) <= '1';
    layer3_outputs(518) <= a;
    layer3_outputs(519) <= not (a and b);
    layer3_outputs(520) <= '0';
    layer3_outputs(521) <= a;
    layer3_outputs(522) <= not b;
    layer3_outputs(523) <= '0';
    layer3_outputs(524) <= not a;
    layer3_outputs(525) <= a;
    layer3_outputs(526) <= not a;
    layer3_outputs(527) <= '1';
    layer3_outputs(528) <= b;
    layer3_outputs(529) <= not a or b;
    layer3_outputs(530) <= a and not b;
    layer3_outputs(531) <= '1';
    layer3_outputs(532) <= not (a or b);
    layer3_outputs(533) <= a or b;
    layer3_outputs(534) <= not b;
    layer3_outputs(535) <= not (a and b);
    layer3_outputs(536) <= a and b;
    layer3_outputs(537) <= b and not a;
    layer3_outputs(538) <= '0';
    layer3_outputs(539) <= a;
    layer3_outputs(540) <= not (a or b);
    layer3_outputs(541) <= '0';
    layer3_outputs(542) <= a or b;
    layer3_outputs(543) <= not (a or b);
    layer3_outputs(544) <= not (a xor b);
    layer3_outputs(545) <= not b;
    layer3_outputs(546) <= not b;
    layer3_outputs(547) <= '1';
    layer3_outputs(548) <= b and not a;
    layer3_outputs(549) <= '1';
    layer3_outputs(550) <= not b;
    layer3_outputs(551) <= not b;
    layer3_outputs(552) <= b;
    layer3_outputs(553) <= not a or b;
    layer3_outputs(554) <= not a;
    layer3_outputs(555) <= not b or a;
    layer3_outputs(556) <= b;
    layer3_outputs(557) <= '1';
    layer3_outputs(558) <= not a or b;
    layer3_outputs(559) <= a or b;
    layer3_outputs(560) <= not a or b;
    layer3_outputs(561) <= '1';
    layer3_outputs(562) <= a and not b;
    layer3_outputs(563) <= not b or a;
    layer3_outputs(564) <= a;
    layer3_outputs(565) <= a xor b;
    layer3_outputs(566) <= b;
    layer3_outputs(567) <= '1';
    layer3_outputs(568) <= not a;
    layer3_outputs(569) <= b;
    layer3_outputs(570) <= a and b;
    layer3_outputs(571) <= '1';
    layer3_outputs(572) <= '1';
    layer3_outputs(573) <= '0';
    layer3_outputs(574) <= not b or a;
    layer3_outputs(575) <= a and not b;
    layer3_outputs(576) <= b;
    layer3_outputs(577) <= a and not b;
    layer3_outputs(578) <= not b;
    layer3_outputs(579) <= '1';
    layer3_outputs(580) <= not b or a;
    layer3_outputs(581) <= not a or b;
    layer3_outputs(582) <= not a;
    layer3_outputs(583) <= a or b;
    layer3_outputs(584) <= not a or b;
    layer3_outputs(585) <= not (a or b);
    layer3_outputs(586) <= a or b;
    layer3_outputs(587) <= a xor b;
    layer3_outputs(588) <= b;
    layer3_outputs(589) <= not (a and b);
    layer3_outputs(590) <= not b;
    layer3_outputs(591) <= a and b;
    layer3_outputs(592) <= a or b;
    layer3_outputs(593) <= '0';
    layer3_outputs(594) <= b;
    layer3_outputs(595) <= b;
    layer3_outputs(596) <= not b;
    layer3_outputs(597) <= a or b;
    layer3_outputs(598) <= not a;
    layer3_outputs(599) <= not a or b;
    layer3_outputs(600) <= not b or a;
    layer3_outputs(601) <= b;
    layer3_outputs(602) <= a and not b;
    layer3_outputs(603) <= a and not b;
    layer3_outputs(604) <= a and b;
    layer3_outputs(605) <= not a;
    layer3_outputs(606) <= a;
    layer3_outputs(607) <= '0';
    layer3_outputs(608) <= a and b;
    layer3_outputs(609) <= not a or b;
    layer3_outputs(610) <= not a;
    layer3_outputs(611) <= b and not a;
    layer3_outputs(612) <= '1';
    layer3_outputs(613) <= a;
    layer3_outputs(614) <= not (a and b);
    layer3_outputs(615) <= not (a or b);
    layer3_outputs(616) <= not (a and b);
    layer3_outputs(617) <= not a or b;
    layer3_outputs(618) <= not (a xor b);
    layer3_outputs(619) <= not (a and b);
    layer3_outputs(620) <= not a or b;
    layer3_outputs(621) <= '1';
    layer3_outputs(622) <= '0';
    layer3_outputs(623) <= a or b;
    layer3_outputs(624) <= a and not b;
    layer3_outputs(625) <= a or b;
    layer3_outputs(626) <= not b or a;
    layer3_outputs(627) <= b;
    layer3_outputs(628) <= not b or a;
    layer3_outputs(629) <= not (a or b);
    layer3_outputs(630) <= not (a and b);
    layer3_outputs(631) <= a;
    layer3_outputs(632) <= not b;
    layer3_outputs(633) <= not a;
    layer3_outputs(634) <= not b or a;
    layer3_outputs(635) <= not (a or b);
    layer3_outputs(636) <= a or b;
    layer3_outputs(637) <= a and b;
    layer3_outputs(638) <= a;
    layer3_outputs(639) <= '1';
    layer3_outputs(640) <= not (a and b);
    layer3_outputs(641) <= not a or b;
    layer3_outputs(642) <= a;
    layer3_outputs(643) <= not b or a;
    layer3_outputs(644) <= a and not b;
    layer3_outputs(645) <= b and not a;
    layer3_outputs(646) <= not b or a;
    layer3_outputs(647) <= not b or a;
    layer3_outputs(648) <= not a;
    layer3_outputs(649) <= not b;
    layer3_outputs(650) <= a;
    layer3_outputs(651) <= a and b;
    layer3_outputs(652) <= not (a xor b);
    layer3_outputs(653) <= not (a and b);
    layer3_outputs(654) <= a;
    layer3_outputs(655) <= '0';
    layer3_outputs(656) <= a and not b;
    layer3_outputs(657) <= a or b;
    layer3_outputs(658) <= a xor b;
    layer3_outputs(659) <= not b;
    layer3_outputs(660) <= a;
    layer3_outputs(661) <= a and not b;
    layer3_outputs(662) <= a or b;
    layer3_outputs(663) <= not (a and b);
    layer3_outputs(664) <= not (a or b);
    layer3_outputs(665) <= not b;
    layer3_outputs(666) <= not a;
    layer3_outputs(667) <= not a;
    layer3_outputs(668) <= not (a or b);
    layer3_outputs(669) <= not a;
    layer3_outputs(670) <= '1';
    layer3_outputs(671) <= a or b;
    layer3_outputs(672) <= '1';
    layer3_outputs(673) <= a;
    layer3_outputs(674) <= b;
    layer3_outputs(675) <= '1';
    layer3_outputs(676) <= not (a xor b);
    layer3_outputs(677) <= '0';
    layer3_outputs(678) <= b;
    layer3_outputs(679) <= not (a and b);
    layer3_outputs(680) <= not b;
    layer3_outputs(681) <= not a or b;
    layer3_outputs(682) <= not b;
    layer3_outputs(683) <= not a or b;
    layer3_outputs(684) <= not b or a;
    layer3_outputs(685) <= not (a xor b);
    layer3_outputs(686) <= not a;
    layer3_outputs(687) <= not a or b;
    layer3_outputs(688) <= not (a and b);
    layer3_outputs(689) <= b and not a;
    layer3_outputs(690) <= not b;
    layer3_outputs(691) <= a and b;
    layer3_outputs(692) <= a or b;
    layer3_outputs(693) <= '1';
    layer3_outputs(694) <= b and not a;
    layer3_outputs(695) <= not b;
    layer3_outputs(696) <= '0';
    layer3_outputs(697) <= b;
    layer3_outputs(698) <= not b or a;
    layer3_outputs(699) <= b;
    layer3_outputs(700) <= '1';
    layer3_outputs(701) <= not (a and b);
    layer3_outputs(702) <= not a or b;
    layer3_outputs(703) <= not b or a;
    layer3_outputs(704) <= not a;
    layer3_outputs(705) <= a;
    layer3_outputs(706) <= not a;
    layer3_outputs(707) <= a;
    layer3_outputs(708) <= not (a or b);
    layer3_outputs(709) <= not a or b;
    layer3_outputs(710) <= a and b;
    layer3_outputs(711) <= not (a and b);
    layer3_outputs(712) <= b;
    layer3_outputs(713) <= b and not a;
    layer3_outputs(714) <= not (a and b);
    layer3_outputs(715) <= b and not a;
    layer3_outputs(716) <= b;
    layer3_outputs(717) <= b;
    layer3_outputs(718) <= a and not b;
    layer3_outputs(719) <= not (a and b);
    layer3_outputs(720) <= b and not a;
    layer3_outputs(721) <= not a;
    layer3_outputs(722) <= '1';
    layer3_outputs(723) <= '1';
    layer3_outputs(724) <= b and not a;
    layer3_outputs(725) <= a and b;
    layer3_outputs(726) <= a;
    layer3_outputs(727) <= not a;
    layer3_outputs(728) <= not a or b;
    layer3_outputs(729) <= a and b;
    layer3_outputs(730) <= '1';
    layer3_outputs(731) <= a and b;
    layer3_outputs(732) <= a;
    layer3_outputs(733) <= not a or b;
    layer3_outputs(734) <= a;
    layer3_outputs(735) <= not b or a;
    layer3_outputs(736) <= b;
    layer3_outputs(737) <= not a;
    layer3_outputs(738) <= not b or a;
    layer3_outputs(739) <= not (a and b);
    layer3_outputs(740) <= '1';
    layer3_outputs(741) <= not a or b;
    layer3_outputs(742) <= b;
    layer3_outputs(743) <= b and not a;
    layer3_outputs(744) <= '1';
    layer3_outputs(745) <= b;
    layer3_outputs(746) <= not a;
    layer3_outputs(747) <= a and not b;
    layer3_outputs(748) <= a and b;
    layer3_outputs(749) <= not a;
    layer3_outputs(750) <= a and b;
    layer3_outputs(751) <= not (a or b);
    layer3_outputs(752) <= b;
    layer3_outputs(753) <= a xor b;
    layer3_outputs(754) <= not a;
    layer3_outputs(755) <= '1';
    layer3_outputs(756) <= not b;
    layer3_outputs(757) <= a or b;
    layer3_outputs(758) <= not (a and b);
    layer3_outputs(759) <= not (a and b);
    layer3_outputs(760) <= not b or a;
    layer3_outputs(761) <= a and not b;
    layer3_outputs(762) <= not a;
    layer3_outputs(763) <= not (a and b);
    layer3_outputs(764) <= not (a or b);
    layer3_outputs(765) <= a and not b;
    layer3_outputs(766) <= '0';
    layer3_outputs(767) <= not b;
    layer3_outputs(768) <= a and b;
    layer3_outputs(769) <= a or b;
    layer3_outputs(770) <= not (a or b);
    layer3_outputs(771) <= a xor b;
    layer3_outputs(772) <= a or b;
    layer3_outputs(773) <= '1';
    layer3_outputs(774) <= b and not a;
    layer3_outputs(775) <= b;
    layer3_outputs(776) <= not a or b;
    layer3_outputs(777) <= a;
    layer3_outputs(778) <= not b or a;
    layer3_outputs(779) <= b;
    layer3_outputs(780) <= a;
    layer3_outputs(781) <= a;
    layer3_outputs(782) <= not a;
    layer3_outputs(783) <= a and not b;
    layer3_outputs(784) <= a or b;
    layer3_outputs(785) <= not b or a;
    layer3_outputs(786) <= not (a or b);
    layer3_outputs(787) <= '0';
    layer3_outputs(788) <= not (a or b);
    layer3_outputs(789) <= not a;
    layer3_outputs(790) <= '0';
    layer3_outputs(791) <= a and b;
    layer3_outputs(792) <= not b or a;
    layer3_outputs(793) <= a;
    layer3_outputs(794) <= not a;
    layer3_outputs(795) <= '0';
    layer3_outputs(796) <= b and not a;
    layer3_outputs(797) <= not a or b;
    layer3_outputs(798) <= not (a or b);
    layer3_outputs(799) <= not (a and b);
    layer3_outputs(800) <= not b or a;
    layer3_outputs(801) <= a and not b;
    layer3_outputs(802) <= not a or b;
    layer3_outputs(803) <= b and not a;
    layer3_outputs(804) <= '0';
    layer3_outputs(805) <= not a;
    layer3_outputs(806) <= a or b;
    layer3_outputs(807) <= a or b;
    layer3_outputs(808) <= '0';
    layer3_outputs(809) <= a;
    layer3_outputs(810) <= b;
    layer3_outputs(811) <= not a;
    layer3_outputs(812) <= not (a or b);
    layer3_outputs(813) <= a or b;
    layer3_outputs(814) <= '0';
    layer3_outputs(815) <= not a;
    layer3_outputs(816) <= a and not b;
    layer3_outputs(817) <= '0';
    layer3_outputs(818) <= a xor b;
    layer3_outputs(819) <= not (a xor b);
    layer3_outputs(820) <= '0';
    layer3_outputs(821) <= a and not b;
    layer3_outputs(822) <= not (a and b);
    layer3_outputs(823) <= '1';
    layer3_outputs(824) <= not a;
    layer3_outputs(825) <= not a;
    layer3_outputs(826) <= a and b;
    layer3_outputs(827) <= b and not a;
    layer3_outputs(828) <= a or b;
    layer3_outputs(829) <= a and not b;
    layer3_outputs(830) <= not (a xor b);
    layer3_outputs(831) <= b and not a;
    layer3_outputs(832) <= b and not a;
    layer3_outputs(833) <= '1';
    layer3_outputs(834) <= a and b;
    layer3_outputs(835) <= a xor b;
    layer3_outputs(836) <= b and not a;
    layer3_outputs(837) <= a and not b;
    layer3_outputs(838) <= not a;
    layer3_outputs(839) <= '1';
    layer3_outputs(840) <= a or b;
    layer3_outputs(841) <= not a;
    layer3_outputs(842) <= '0';
    layer3_outputs(843) <= not a or b;
    layer3_outputs(844) <= not b or a;
    layer3_outputs(845) <= b and not a;
    layer3_outputs(846) <= a or b;
    layer3_outputs(847) <= a and b;
    layer3_outputs(848) <= not b;
    layer3_outputs(849) <= not b;
    layer3_outputs(850) <= a and not b;
    layer3_outputs(851) <= a or b;
    layer3_outputs(852) <= not b;
    layer3_outputs(853) <= b and not a;
    layer3_outputs(854) <= a xor b;
    layer3_outputs(855) <= '0';
    layer3_outputs(856) <= not (a and b);
    layer3_outputs(857) <= not (a and b);
    layer3_outputs(858) <= not b or a;
    layer3_outputs(859) <= a;
    layer3_outputs(860) <= a xor b;
    layer3_outputs(861) <= '0';
    layer3_outputs(862) <= a or b;
    layer3_outputs(863) <= a and b;
    layer3_outputs(864) <= a xor b;
    layer3_outputs(865) <= a or b;
    layer3_outputs(866) <= not a or b;
    layer3_outputs(867) <= not b;
    layer3_outputs(868) <= a;
    layer3_outputs(869) <= not a or b;
    layer3_outputs(870) <= a;
    layer3_outputs(871) <= a or b;
    layer3_outputs(872) <= not (a xor b);
    layer3_outputs(873) <= not a or b;
    layer3_outputs(874) <= b;
    layer3_outputs(875) <= a and b;
    layer3_outputs(876) <= not (a and b);
    layer3_outputs(877) <= a and b;
    layer3_outputs(878) <= b and not a;
    layer3_outputs(879) <= b and not a;
    layer3_outputs(880) <= b;
    layer3_outputs(881) <= b;
    layer3_outputs(882) <= not (a and b);
    layer3_outputs(883) <= '0';
    layer3_outputs(884) <= a and b;
    layer3_outputs(885) <= a or b;
    layer3_outputs(886) <= a and b;
    layer3_outputs(887) <= a;
    layer3_outputs(888) <= not a or b;
    layer3_outputs(889) <= '0';
    layer3_outputs(890) <= a and not b;
    layer3_outputs(891) <= '0';
    layer3_outputs(892) <= not b;
    layer3_outputs(893) <= b and not a;
    layer3_outputs(894) <= a xor b;
    layer3_outputs(895) <= not a or b;
    layer3_outputs(896) <= not b or a;
    layer3_outputs(897) <= '0';
    layer3_outputs(898) <= not a;
    layer3_outputs(899) <= a and not b;
    layer3_outputs(900) <= not b or a;
    layer3_outputs(901) <= a or b;
    layer3_outputs(902) <= not a or b;
    layer3_outputs(903) <= a and not b;
    layer3_outputs(904) <= not (a and b);
    layer3_outputs(905) <= a and not b;
    layer3_outputs(906) <= a and b;
    layer3_outputs(907) <= a;
    layer3_outputs(908) <= '0';
    layer3_outputs(909) <= a xor b;
    layer3_outputs(910) <= not (a xor b);
    layer3_outputs(911) <= not (a or b);
    layer3_outputs(912) <= not (a and b);
    layer3_outputs(913) <= not b;
    layer3_outputs(914) <= b;
    layer3_outputs(915) <= '0';
    layer3_outputs(916) <= not a or b;
    layer3_outputs(917) <= not (a or b);
    layer3_outputs(918) <= a xor b;
    layer3_outputs(919) <= not a or b;
    layer3_outputs(920) <= '0';
    layer3_outputs(921) <= not b;
    layer3_outputs(922) <= a;
    layer3_outputs(923) <= a and not b;
    layer3_outputs(924) <= not (a or b);
    layer3_outputs(925) <= a and not b;
    layer3_outputs(926) <= not b;
    layer3_outputs(927) <= not (a and b);
    layer3_outputs(928) <= a or b;
    layer3_outputs(929) <= not (a and b);
    layer3_outputs(930) <= b;
    layer3_outputs(931) <= not (a or b);
    layer3_outputs(932) <= not a;
    layer3_outputs(933) <= not b;
    layer3_outputs(934) <= not b;
    layer3_outputs(935) <= not (a or b);
    layer3_outputs(936) <= a or b;
    layer3_outputs(937) <= not b or a;
    layer3_outputs(938) <= a and not b;
    layer3_outputs(939) <= not b or a;
    layer3_outputs(940) <= not b;
    layer3_outputs(941) <= '0';
    layer3_outputs(942) <= a;
    layer3_outputs(943) <= not b or a;
    layer3_outputs(944) <= a or b;
    layer3_outputs(945) <= not (a or b);
    layer3_outputs(946) <= not (a and b);
    layer3_outputs(947) <= not b or a;
    layer3_outputs(948) <= b;
    layer3_outputs(949) <= a and not b;
    layer3_outputs(950) <= '1';
    layer3_outputs(951) <= a and b;
    layer3_outputs(952) <= a;
    layer3_outputs(953) <= a and b;
    layer3_outputs(954) <= a and b;
    layer3_outputs(955) <= b;
    layer3_outputs(956) <= not (a or b);
    layer3_outputs(957) <= a and not b;
    layer3_outputs(958) <= not a;
    layer3_outputs(959) <= '1';
    layer3_outputs(960) <= not (a or b);
    layer3_outputs(961) <= b and not a;
    layer3_outputs(962) <= a or b;
    layer3_outputs(963) <= not b;
    layer3_outputs(964) <= b;
    layer3_outputs(965) <= not b;
    layer3_outputs(966) <= not b;
    layer3_outputs(967) <= b;
    layer3_outputs(968) <= '0';
    layer3_outputs(969) <= not a;
    layer3_outputs(970) <= b;
    layer3_outputs(971) <= b and not a;
    layer3_outputs(972) <= not a or b;
    layer3_outputs(973) <= b;
    layer3_outputs(974) <= not b;
    layer3_outputs(975) <= not (a or b);
    layer3_outputs(976) <= not b;
    layer3_outputs(977) <= '0';
    layer3_outputs(978) <= not a;
    layer3_outputs(979) <= '1';
    layer3_outputs(980) <= not b;
    layer3_outputs(981) <= a and b;
    layer3_outputs(982) <= not (a and b);
    layer3_outputs(983) <= a or b;
    layer3_outputs(984) <= a xor b;
    layer3_outputs(985) <= a or b;
    layer3_outputs(986) <= '1';
    layer3_outputs(987) <= '0';
    layer3_outputs(988) <= not b or a;
    layer3_outputs(989) <= b and not a;
    layer3_outputs(990) <= '0';
    layer3_outputs(991) <= not (a and b);
    layer3_outputs(992) <= a;
    layer3_outputs(993) <= not a or b;
    layer3_outputs(994) <= a xor b;
    layer3_outputs(995) <= not a or b;
    layer3_outputs(996) <= '1';
    layer3_outputs(997) <= '1';
    layer3_outputs(998) <= a and b;
    layer3_outputs(999) <= not b or a;
    layer3_outputs(1000) <= not b;
    layer3_outputs(1001) <= not (a and b);
    layer3_outputs(1002) <= a xor b;
    layer3_outputs(1003) <= '0';
    layer3_outputs(1004) <= not (a and b);
    layer3_outputs(1005) <= '1';
    layer3_outputs(1006) <= '1';
    layer3_outputs(1007) <= not (a or b);
    layer3_outputs(1008) <= not a or b;
    layer3_outputs(1009) <= not b;
    layer3_outputs(1010) <= a or b;
    layer3_outputs(1011) <= a and b;
    layer3_outputs(1012) <= a or b;
    layer3_outputs(1013) <= a and b;
    layer3_outputs(1014) <= a and b;
    layer3_outputs(1015) <= a and b;
    layer3_outputs(1016) <= a;
    layer3_outputs(1017) <= b;
    layer3_outputs(1018) <= a;
    layer3_outputs(1019) <= not a or b;
    layer3_outputs(1020) <= b;
    layer3_outputs(1021) <= b;
    layer3_outputs(1022) <= not (a or b);
    layer3_outputs(1023) <= a;
    layer3_outputs(1024) <= '1';
    layer3_outputs(1025) <= not (a or b);
    layer3_outputs(1026) <= a or b;
    layer3_outputs(1027) <= a;
    layer3_outputs(1028) <= not (a or b);
    layer3_outputs(1029) <= not (a or b);
    layer3_outputs(1030) <= not b;
    layer3_outputs(1031) <= a and not b;
    layer3_outputs(1032) <= b and not a;
    layer3_outputs(1033) <= b;
    layer3_outputs(1034) <= not (a and b);
    layer3_outputs(1035) <= not b or a;
    layer3_outputs(1036) <= not (a xor b);
    layer3_outputs(1037) <= not (a or b);
    layer3_outputs(1038) <= '1';
    layer3_outputs(1039) <= a and b;
    layer3_outputs(1040) <= not (a or b);
    layer3_outputs(1041) <= not b;
    layer3_outputs(1042) <= not (a and b);
    layer3_outputs(1043) <= a;
    layer3_outputs(1044) <= '0';
    layer3_outputs(1045) <= not (a or b);
    layer3_outputs(1046) <= not (a and b);
    layer3_outputs(1047) <= a or b;
    layer3_outputs(1048) <= a or b;
    layer3_outputs(1049) <= '0';
    layer3_outputs(1050) <= '1';
    layer3_outputs(1051) <= a and not b;
    layer3_outputs(1052) <= a;
    layer3_outputs(1053) <= not b or a;
    layer3_outputs(1054) <= not b or a;
    layer3_outputs(1055) <= a and b;
    layer3_outputs(1056) <= not a;
    layer3_outputs(1057) <= not a;
    layer3_outputs(1058) <= a;
    layer3_outputs(1059) <= not b;
    layer3_outputs(1060) <= a or b;
    layer3_outputs(1061) <= not b;
    layer3_outputs(1062) <= not a or b;
    layer3_outputs(1063) <= b and not a;
    layer3_outputs(1064) <= not a;
    layer3_outputs(1065) <= '1';
    layer3_outputs(1066) <= a;
    layer3_outputs(1067) <= '1';
    layer3_outputs(1068) <= not a or b;
    layer3_outputs(1069) <= not a;
    layer3_outputs(1070) <= not (a xor b);
    layer3_outputs(1071) <= b and not a;
    layer3_outputs(1072) <= '1';
    layer3_outputs(1073) <= b;
    layer3_outputs(1074) <= not a;
    layer3_outputs(1075) <= not b;
    layer3_outputs(1076) <= not (a or b);
    layer3_outputs(1077) <= a and b;
    layer3_outputs(1078) <= a or b;
    layer3_outputs(1079) <= a;
    layer3_outputs(1080) <= not b;
    layer3_outputs(1081) <= a;
    layer3_outputs(1082) <= not a or b;
    layer3_outputs(1083) <= a and b;
    layer3_outputs(1084) <= not a;
    layer3_outputs(1085) <= '1';
    layer3_outputs(1086) <= '0';
    layer3_outputs(1087) <= a and not b;
    layer3_outputs(1088) <= not a;
    layer3_outputs(1089) <= not (a or b);
    layer3_outputs(1090) <= not (a and b);
    layer3_outputs(1091) <= '0';
    layer3_outputs(1092) <= a or b;
    layer3_outputs(1093) <= not a or b;
    layer3_outputs(1094) <= not b;
    layer3_outputs(1095) <= '1';
    layer3_outputs(1096) <= a and not b;
    layer3_outputs(1097) <= not a;
    layer3_outputs(1098) <= not b or a;
    layer3_outputs(1099) <= not b or a;
    layer3_outputs(1100) <= b and not a;
    layer3_outputs(1101) <= a and not b;
    layer3_outputs(1102) <= '0';
    layer3_outputs(1103) <= not b;
    layer3_outputs(1104) <= b;
    layer3_outputs(1105) <= not a or b;
    layer3_outputs(1106) <= b and not a;
    layer3_outputs(1107) <= not b;
    layer3_outputs(1108) <= a;
    layer3_outputs(1109) <= b and not a;
    layer3_outputs(1110) <= not b or a;
    layer3_outputs(1111) <= not (a and b);
    layer3_outputs(1112) <= not (a or b);
    layer3_outputs(1113) <= b;
    layer3_outputs(1114) <= a;
    layer3_outputs(1115) <= not a;
    layer3_outputs(1116) <= not a or b;
    layer3_outputs(1117) <= not a;
    layer3_outputs(1118) <= a;
    layer3_outputs(1119) <= not b or a;
    layer3_outputs(1120) <= '0';
    layer3_outputs(1121) <= b and not a;
    layer3_outputs(1122) <= '0';
    layer3_outputs(1123) <= a;
    layer3_outputs(1124) <= a;
    layer3_outputs(1125) <= '1';
    layer3_outputs(1126) <= not (a or b);
    layer3_outputs(1127) <= not (a and b);
    layer3_outputs(1128) <= a and not b;
    layer3_outputs(1129) <= '1';
    layer3_outputs(1130) <= not a or b;
    layer3_outputs(1131) <= a and b;
    layer3_outputs(1132) <= '1';
    layer3_outputs(1133) <= b and not a;
    layer3_outputs(1134) <= a and b;
    layer3_outputs(1135) <= a and not b;
    layer3_outputs(1136) <= a and not b;
    layer3_outputs(1137) <= not a;
    layer3_outputs(1138) <= a or b;
    layer3_outputs(1139) <= '0';
    layer3_outputs(1140) <= not (a and b);
    layer3_outputs(1141) <= not a;
    layer3_outputs(1142) <= a or b;
    layer3_outputs(1143) <= not b or a;
    layer3_outputs(1144) <= '1';
    layer3_outputs(1145) <= not a;
    layer3_outputs(1146) <= b and not a;
    layer3_outputs(1147) <= a and not b;
    layer3_outputs(1148) <= not b;
    layer3_outputs(1149) <= not b;
    layer3_outputs(1150) <= b and not a;
    layer3_outputs(1151) <= not b or a;
    layer3_outputs(1152) <= a and b;
    layer3_outputs(1153) <= '0';
    layer3_outputs(1154) <= not a;
    layer3_outputs(1155) <= '1';
    layer3_outputs(1156) <= not a;
    layer3_outputs(1157) <= not (a or b);
    layer3_outputs(1158) <= b and not a;
    layer3_outputs(1159) <= not a or b;
    layer3_outputs(1160) <= not b;
    layer3_outputs(1161) <= '0';
    layer3_outputs(1162) <= not (a and b);
    layer3_outputs(1163) <= b;
    layer3_outputs(1164) <= a and not b;
    layer3_outputs(1165) <= not (a or b);
    layer3_outputs(1166) <= not (a and b);
    layer3_outputs(1167) <= a and not b;
    layer3_outputs(1168) <= not (a or b);
    layer3_outputs(1169) <= not b or a;
    layer3_outputs(1170) <= b;
    layer3_outputs(1171) <= not (a xor b);
    layer3_outputs(1172) <= not (a or b);
    layer3_outputs(1173) <= a;
    layer3_outputs(1174) <= not (a or b);
    layer3_outputs(1175) <= a and b;
    layer3_outputs(1176) <= '1';
    layer3_outputs(1177) <= b;
    layer3_outputs(1178) <= not a or b;
    layer3_outputs(1179) <= not a or b;
    layer3_outputs(1180) <= b and not a;
    layer3_outputs(1181) <= a and not b;
    layer3_outputs(1182) <= a;
    layer3_outputs(1183) <= '0';
    layer3_outputs(1184) <= '0';
    layer3_outputs(1185) <= not b;
    layer3_outputs(1186) <= not a;
    layer3_outputs(1187) <= a and b;
    layer3_outputs(1188) <= b and not a;
    layer3_outputs(1189) <= not b;
    layer3_outputs(1190) <= a or b;
    layer3_outputs(1191) <= not (a and b);
    layer3_outputs(1192) <= not b;
    layer3_outputs(1193) <= not (a and b);
    layer3_outputs(1194) <= a and not b;
    layer3_outputs(1195) <= a and b;
    layer3_outputs(1196) <= not a;
    layer3_outputs(1197) <= not b;
    layer3_outputs(1198) <= not b or a;
    layer3_outputs(1199) <= b;
    layer3_outputs(1200) <= not (a or b);
    layer3_outputs(1201) <= not (a and b);
    layer3_outputs(1202) <= not b;
    layer3_outputs(1203) <= not b;
    layer3_outputs(1204) <= b and not a;
    layer3_outputs(1205) <= not (a and b);
    layer3_outputs(1206) <= '1';
    layer3_outputs(1207) <= not (a and b);
    layer3_outputs(1208) <= not (a or b);
    layer3_outputs(1209) <= a and not b;
    layer3_outputs(1210) <= not a or b;
    layer3_outputs(1211) <= not b or a;
    layer3_outputs(1212) <= not b or a;
    layer3_outputs(1213) <= b;
    layer3_outputs(1214) <= not b or a;
    layer3_outputs(1215) <= a and not b;
    layer3_outputs(1216) <= not (a and b);
    layer3_outputs(1217) <= '0';
    layer3_outputs(1218) <= b and not a;
    layer3_outputs(1219) <= a and b;
    layer3_outputs(1220) <= not b;
    layer3_outputs(1221) <= '1';
    layer3_outputs(1222) <= not (a and b);
    layer3_outputs(1223) <= not a;
    layer3_outputs(1224) <= a or b;
    layer3_outputs(1225) <= not (a and b);
    layer3_outputs(1226) <= '0';
    layer3_outputs(1227) <= b and not a;
    layer3_outputs(1228) <= a;
    layer3_outputs(1229) <= a and not b;
    layer3_outputs(1230) <= '1';
    layer3_outputs(1231) <= a or b;
    layer3_outputs(1232) <= not (a or b);
    layer3_outputs(1233) <= a and b;
    layer3_outputs(1234) <= '0';
    layer3_outputs(1235) <= '1';
    layer3_outputs(1236) <= a and b;
    layer3_outputs(1237) <= not a or b;
    layer3_outputs(1238) <= not (a or b);
    layer3_outputs(1239) <= b and not a;
    layer3_outputs(1240) <= not b;
    layer3_outputs(1241) <= not (a or b);
    layer3_outputs(1242) <= a xor b;
    layer3_outputs(1243) <= not b or a;
    layer3_outputs(1244) <= '1';
    layer3_outputs(1245) <= '0';
    layer3_outputs(1246) <= not (a or b);
    layer3_outputs(1247) <= not (a and b);
    layer3_outputs(1248) <= b and not a;
    layer3_outputs(1249) <= b;
    layer3_outputs(1250) <= '0';
    layer3_outputs(1251) <= '0';
    layer3_outputs(1252) <= a and not b;
    layer3_outputs(1253) <= a and b;
    layer3_outputs(1254) <= not (a and b);
    layer3_outputs(1255) <= not b or a;
    layer3_outputs(1256) <= a and b;
    layer3_outputs(1257) <= a or b;
    layer3_outputs(1258) <= not (a xor b);
    layer3_outputs(1259) <= a or b;
    layer3_outputs(1260) <= not b or a;
    layer3_outputs(1261) <= a;
    layer3_outputs(1262) <= b;
    layer3_outputs(1263) <= not (a or b);
    layer3_outputs(1264) <= b and not a;
    layer3_outputs(1265) <= not a or b;
    layer3_outputs(1266) <= not a or b;
    layer3_outputs(1267) <= b;
    layer3_outputs(1268) <= not a;
    layer3_outputs(1269) <= '1';
    layer3_outputs(1270) <= not (a or b);
    layer3_outputs(1271) <= a or b;
    layer3_outputs(1272) <= a and not b;
    layer3_outputs(1273) <= not a or b;
    layer3_outputs(1274) <= not b;
    layer3_outputs(1275) <= a or b;
    layer3_outputs(1276) <= a and b;
    layer3_outputs(1277) <= a and not b;
    layer3_outputs(1278) <= a and b;
    layer3_outputs(1279) <= a;
    layer3_outputs(1280) <= not a or b;
    layer3_outputs(1281) <= not a or b;
    layer3_outputs(1282) <= not b or a;
    layer3_outputs(1283) <= not b;
    layer3_outputs(1284) <= '0';
    layer3_outputs(1285) <= not (a or b);
    layer3_outputs(1286) <= not a or b;
    layer3_outputs(1287) <= b and not a;
    layer3_outputs(1288) <= a and b;
    layer3_outputs(1289) <= not b;
    layer3_outputs(1290) <= a;
    layer3_outputs(1291) <= not b;
    layer3_outputs(1292) <= a;
    layer3_outputs(1293) <= '0';
    layer3_outputs(1294) <= b;
    layer3_outputs(1295) <= b and not a;
    layer3_outputs(1296) <= '0';
    layer3_outputs(1297) <= not a or b;
    layer3_outputs(1298) <= a or b;
    layer3_outputs(1299) <= not (a and b);
    layer3_outputs(1300) <= not (a or b);
    layer3_outputs(1301) <= b and not a;
    layer3_outputs(1302) <= '1';
    layer3_outputs(1303) <= b and not a;
    layer3_outputs(1304) <= a or b;
    layer3_outputs(1305) <= not a;
    layer3_outputs(1306) <= '1';
    layer3_outputs(1307) <= not (a or b);
    layer3_outputs(1308) <= '0';
    layer3_outputs(1309) <= not a or b;
    layer3_outputs(1310) <= not (a or b);
    layer3_outputs(1311) <= b and not a;
    layer3_outputs(1312) <= a and not b;
    layer3_outputs(1313) <= not b;
    layer3_outputs(1314) <= not b or a;
    layer3_outputs(1315) <= '1';
    layer3_outputs(1316) <= b;
    layer3_outputs(1317) <= a or b;
    layer3_outputs(1318) <= not a;
    layer3_outputs(1319) <= a or b;
    layer3_outputs(1320) <= not (a and b);
    layer3_outputs(1321) <= a or b;
    layer3_outputs(1322) <= not b or a;
    layer3_outputs(1323) <= b and not a;
    layer3_outputs(1324) <= a and not b;
    layer3_outputs(1325) <= a and b;
    layer3_outputs(1326) <= not (a or b);
    layer3_outputs(1327) <= not b or a;
    layer3_outputs(1328) <= not (a or b);
    layer3_outputs(1329) <= not a or b;
    layer3_outputs(1330) <= not b;
    layer3_outputs(1331) <= not (a and b);
    layer3_outputs(1332) <= not (a and b);
    layer3_outputs(1333) <= b and not a;
    layer3_outputs(1334) <= a xor b;
    layer3_outputs(1335) <= not (a or b);
    layer3_outputs(1336) <= a or b;
    layer3_outputs(1337) <= not b;
    layer3_outputs(1338) <= not (a and b);
    layer3_outputs(1339) <= b;
    layer3_outputs(1340) <= not b or a;
    layer3_outputs(1341) <= not a;
    layer3_outputs(1342) <= b and not a;
    layer3_outputs(1343) <= b and not a;
    layer3_outputs(1344) <= a xor b;
    layer3_outputs(1345) <= b;
    layer3_outputs(1346) <= not a or b;
    layer3_outputs(1347) <= b and not a;
    layer3_outputs(1348) <= not b;
    layer3_outputs(1349) <= b and not a;
    layer3_outputs(1350) <= not (a xor b);
    layer3_outputs(1351) <= a or b;
    layer3_outputs(1352) <= not (a xor b);
    layer3_outputs(1353) <= a and b;
    layer3_outputs(1354) <= a;
    layer3_outputs(1355) <= not a or b;
    layer3_outputs(1356) <= not b or a;
    layer3_outputs(1357) <= not b;
    layer3_outputs(1358) <= b and not a;
    layer3_outputs(1359) <= not (a or b);
    layer3_outputs(1360) <= '0';
    layer3_outputs(1361) <= a and b;
    layer3_outputs(1362) <= not (a or b);
    layer3_outputs(1363) <= '1';
    layer3_outputs(1364) <= a;
    layer3_outputs(1365) <= b;
    layer3_outputs(1366) <= not (a and b);
    layer3_outputs(1367) <= a and not b;
    layer3_outputs(1368) <= not a;
    layer3_outputs(1369) <= a or b;
    layer3_outputs(1370) <= not b or a;
    layer3_outputs(1371) <= b and not a;
    layer3_outputs(1372) <= not b;
    layer3_outputs(1373) <= a and b;
    layer3_outputs(1374) <= not a or b;
    layer3_outputs(1375) <= a and b;
    layer3_outputs(1376) <= a and b;
    layer3_outputs(1377) <= b;
    layer3_outputs(1378) <= not (a and b);
    layer3_outputs(1379) <= a and b;
    layer3_outputs(1380) <= a;
    layer3_outputs(1381) <= '1';
    layer3_outputs(1382) <= a;
    layer3_outputs(1383) <= not b;
    layer3_outputs(1384) <= not (a or b);
    layer3_outputs(1385) <= not (a or b);
    layer3_outputs(1386) <= b and not a;
    layer3_outputs(1387) <= not (a or b);
    layer3_outputs(1388) <= not a;
    layer3_outputs(1389) <= '0';
    layer3_outputs(1390) <= not (a and b);
    layer3_outputs(1391) <= a and not b;
    layer3_outputs(1392) <= not (a or b);
    layer3_outputs(1393) <= a and not b;
    layer3_outputs(1394) <= not (a and b);
    layer3_outputs(1395) <= not a;
    layer3_outputs(1396) <= '1';
    layer3_outputs(1397) <= b and not a;
    layer3_outputs(1398) <= not b or a;
    layer3_outputs(1399) <= a;
    layer3_outputs(1400) <= not (a or b);
    layer3_outputs(1401) <= not a;
    layer3_outputs(1402) <= not b or a;
    layer3_outputs(1403) <= not b or a;
    layer3_outputs(1404) <= not (a or b);
    layer3_outputs(1405) <= not a or b;
    layer3_outputs(1406) <= '1';
    layer3_outputs(1407) <= not a;
    layer3_outputs(1408) <= not (a and b);
    layer3_outputs(1409) <= a and not b;
    layer3_outputs(1410) <= not a;
    layer3_outputs(1411) <= a or b;
    layer3_outputs(1412) <= not b or a;
    layer3_outputs(1413) <= b;
    layer3_outputs(1414) <= not (a and b);
    layer3_outputs(1415) <= b;
    layer3_outputs(1416) <= a and b;
    layer3_outputs(1417) <= not b or a;
    layer3_outputs(1418) <= not (a and b);
    layer3_outputs(1419) <= a or b;
    layer3_outputs(1420) <= not (a and b);
    layer3_outputs(1421) <= a and not b;
    layer3_outputs(1422) <= '0';
    layer3_outputs(1423) <= not a;
    layer3_outputs(1424) <= '1';
    layer3_outputs(1425) <= b and not a;
    layer3_outputs(1426) <= not (a or b);
    layer3_outputs(1427) <= not a or b;
    layer3_outputs(1428) <= a and not b;
    layer3_outputs(1429) <= b and not a;
    layer3_outputs(1430) <= a or b;
    layer3_outputs(1431) <= not b or a;
    layer3_outputs(1432) <= not b;
    layer3_outputs(1433) <= '0';
    layer3_outputs(1434) <= not a;
    layer3_outputs(1435) <= a;
    layer3_outputs(1436) <= a and b;
    layer3_outputs(1437) <= b and not a;
    layer3_outputs(1438) <= '0';
    layer3_outputs(1439) <= '0';
    layer3_outputs(1440) <= not b or a;
    layer3_outputs(1441) <= b and not a;
    layer3_outputs(1442) <= a and not b;
    layer3_outputs(1443) <= b and not a;
    layer3_outputs(1444) <= b;
    layer3_outputs(1445) <= '0';
    layer3_outputs(1446) <= '0';
    layer3_outputs(1447) <= not (a or b);
    layer3_outputs(1448) <= not a or b;
    layer3_outputs(1449) <= a and not b;
    layer3_outputs(1450) <= '1';
    layer3_outputs(1451) <= a;
    layer3_outputs(1452) <= a and b;
    layer3_outputs(1453) <= not b or a;
    layer3_outputs(1454) <= '0';
    layer3_outputs(1455) <= a;
    layer3_outputs(1456) <= '1';
    layer3_outputs(1457) <= a or b;
    layer3_outputs(1458) <= a and b;
    layer3_outputs(1459) <= not b or a;
    layer3_outputs(1460) <= b and not a;
    layer3_outputs(1461) <= not a or b;
    layer3_outputs(1462) <= not (a or b);
    layer3_outputs(1463) <= not (a and b);
    layer3_outputs(1464) <= a or b;
    layer3_outputs(1465) <= not (a and b);
    layer3_outputs(1466) <= not (a or b);
    layer3_outputs(1467) <= a and b;
    layer3_outputs(1468) <= '0';
    layer3_outputs(1469) <= a and not b;
    layer3_outputs(1470) <= '1';
    layer3_outputs(1471) <= b and not a;
    layer3_outputs(1472) <= not a;
    layer3_outputs(1473) <= b;
    layer3_outputs(1474) <= not b;
    layer3_outputs(1475) <= b;
    layer3_outputs(1476) <= not a or b;
    layer3_outputs(1477) <= not a;
    layer3_outputs(1478) <= not a;
    layer3_outputs(1479) <= not a or b;
    layer3_outputs(1480) <= not a;
    layer3_outputs(1481) <= '0';
    layer3_outputs(1482) <= not (a or b);
    layer3_outputs(1483) <= not a;
    layer3_outputs(1484) <= a;
    layer3_outputs(1485) <= a;
    layer3_outputs(1486) <= not b or a;
    layer3_outputs(1487) <= b;
    layer3_outputs(1488) <= not b;
    layer3_outputs(1489) <= '0';
    layer3_outputs(1490) <= a or b;
    layer3_outputs(1491) <= a;
    layer3_outputs(1492) <= '1';
    layer3_outputs(1493) <= b and not a;
    layer3_outputs(1494) <= a or b;
    layer3_outputs(1495) <= a and b;
    layer3_outputs(1496) <= a and not b;
    layer3_outputs(1497) <= a and not b;
    layer3_outputs(1498) <= not (a or b);
    layer3_outputs(1499) <= not b;
    layer3_outputs(1500) <= a or b;
    layer3_outputs(1501) <= not (a xor b);
    layer3_outputs(1502) <= b;
    layer3_outputs(1503) <= not (a and b);
    layer3_outputs(1504) <= b and not a;
    layer3_outputs(1505) <= not (a or b);
    layer3_outputs(1506) <= a or b;
    layer3_outputs(1507) <= a and b;
    layer3_outputs(1508) <= b and not a;
    layer3_outputs(1509) <= a;
    layer3_outputs(1510) <= a or b;
    layer3_outputs(1511) <= b;
    layer3_outputs(1512) <= not (a or b);
    layer3_outputs(1513) <= not (a or b);
    layer3_outputs(1514) <= not (a xor b);
    layer3_outputs(1515) <= b;
    layer3_outputs(1516) <= b and not a;
    layer3_outputs(1517) <= not (a and b);
    layer3_outputs(1518) <= not b or a;
    layer3_outputs(1519) <= a;
    layer3_outputs(1520) <= not b or a;
    layer3_outputs(1521) <= b;
    layer3_outputs(1522) <= a;
    layer3_outputs(1523) <= not b or a;
    layer3_outputs(1524) <= not b or a;
    layer3_outputs(1525) <= not (a or b);
    layer3_outputs(1526) <= b and not a;
    layer3_outputs(1527) <= not b;
    layer3_outputs(1528) <= a;
    layer3_outputs(1529) <= not a;
    layer3_outputs(1530) <= '0';
    layer3_outputs(1531) <= a xor b;
    layer3_outputs(1532) <= not a;
    layer3_outputs(1533) <= '1';
    layer3_outputs(1534) <= not (a and b);
    layer3_outputs(1535) <= not a or b;
    layer3_outputs(1536) <= a and not b;
    layer3_outputs(1537) <= not b;
    layer3_outputs(1538) <= not (a or b);
    layer3_outputs(1539) <= not b;
    layer3_outputs(1540) <= b and not a;
    layer3_outputs(1541) <= a or b;
    layer3_outputs(1542) <= not (a and b);
    layer3_outputs(1543) <= not b;
    layer3_outputs(1544) <= not a or b;
    layer3_outputs(1545) <= not b or a;
    layer3_outputs(1546) <= not (a or b);
    layer3_outputs(1547) <= a and b;
    layer3_outputs(1548) <= '1';
    layer3_outputs(1549) <= a and not b;
    layer3_outputs(1550) <= a and b;
    layer3_outputs(1551) <= not (a xor b);
    layer3_outputs(1552) <= a and not b;
    layer3_outputs(1553) <= a and b;
    layer3_outputs(1554) <= b;
    layer3_outputs(1555) <= not (a and b);
    layer3_outputs(1556) <= not b;
    layer3_outputs(1557) <= '0';
    layer3_outputs(1558) <= not a or b;
    layer3_outputs(1559) <= not a;
    layer3_outputs(1560) <= not a;
    layer3_outputs(1561) <= not (a xor b);
    layer3_outputs(1562) <= a xor b;
    layer3_outputs(1563) <= not (a or b);
    layer3_outputs(1564) <= b and not a;
    layer3_outputs(1565) <= a or b;
    layer3_outputs(1566) <= '0';
    layer3_outputs(1567) <= a and b;
    layer3_outputs(1568) <= not (a or b);
    layer3_outputs(1569) <= a and not b;
    layer3_outputs(1570) <= a;
    layer3_outputs(1571) <= not (a or b);
    layer3_outputs(1572) <= not (a or b);
    layer3_outputs(1573) <= not (a or b);
    layer3_outputs(1574) <= a and b;
    layer3_outputs(1575) <= a and not b;
    layer3_outputs(1576) <= not b;
    layer3_outputs(1577) <= '1';
    layer3_outputs(1578) <= not (a and b);
    layer3_outputs(1579) <= a or b;
    layer3_outputs(1580) <= '1';
    layer3_outputs(1581) <= a xor b;
    layer3_outputs(1582) <= b and not a;
    layer3_outputs(1583) <= '1';
    layer3_outputs(1584) <= b and not a;
    layer3_outputs(1585) <= b;
    layer3_outputs(1586) <= a;
    layer3_outputs(1587) <= '0';
    layer3_outputs(1588) <= not (a and b);
    layer3_outputs(1589) <= not (a and b);
    layer3_outputs(1590) <= not (a and b);
    layer3_outputs(1591) <= a and b;
    layer3_outputs(1592) <= not a or b;
    layer3_outputs(1593) <= not (a or b);
    layer3_outputs(1594) <= b and not a;
    layer3_outputs(1595) <= a;
    layer3_outputs(1596) <= not b or a;
    layer3_outputs(1597) <= a;
    layer3_outputs(1598) <= '0';
    layer3_outputs(1599) <= '1';
    layer3_outputs(1600) <= '1';
    layer3_outputs(1601) <= b and not a;
    layer3_outputs(1602) <= b and not a;
    layer3_outputs(1603) <= a or b;
    layer3_outputs(1604) <= a and b;
    layer3_outputs(1605) <= b;
    layer3_outputs(1606) <= not b;
    layer3_outputs(1607) <= '0';
    layer3_outputs(1608) <= '0';
    layer3_outputs(1609) <= a and not b;
    layer3_outputs(1610) <= not a or b;
    layer3_outputs(1611) <= not b or a;
    layer3_outputs(1612) <= b;
    layer3_outputs(1613) <= a or b;
    layer3_outputs(1614) <= b and not a;
    layer3_outputs(1615) <= not (a or b);
    layer3_outputs(1616) <= not a or b;
    layer3_outputs(1617) <= b;
    layer3_outputs(1618) <= not a;
    layer3_outputs(1619) <= a xor b;
    layer3_outputs(1620) <= not a;
    layer3_outputs(1621) <= a and b;
    layer3_outputs(1622) <= b and not a;
    layer3_outputs(1623) <= not b;
    layer3_outputs(1624) <= a and not b;
    layer3_outputs(1625) <= not a;
    layer3_outputs(1626) <= '0';
    layer3_outputs(1627) <= not b or a;
    layer3_outputs(1628) <= a;
    layer3_outputs(1629) <= not (a and b);
    layer3_outputs(1630) <= b and not a;
    layer3_outputs(1631) <= a and not b;
    layer3_outputs(1632) <= a and b;
    layer3_outputs(1633) <= b;
    layer3_outputs(1634) <= b;
    layer3_outputs(1635) <= a;
    layer3_outputs(1636) <= b and not a;
    layer3_outputs(1637) <= not a or b;
    layer3_outputs(1638) <= a and b;
    layer3_outputs(1639) <= b and not a;
    layer3_outputs(1640) <= a and not b;
    layer3_outputs(1641) <= not (a and b);
    layer3_outputs(1642) <= a and not b;
    layer3_outputs(1643) <= a and b;
    layer3_outputs(1644) <= b and not a;
    layer3_outputs(1645) <= b;
    layer3_outputs(1646) <= '1';
    layer3_outputs(1647) <= a;
    layer3_outputs(1648) <= b and not a;
    layer3_outputs(1649) <= a xor b;
    layer3_outputs(1650) <= not (a or b);
    layer3_outputs(1651) <= not (a or b);
    layer3_outputs(1652) <= not b;
    layer3_outputs(1653) <= '0';
    layer3_outputs(1654) <= a xor b;
    layer3_outputs(1655) <= not (a or b);
    layer3_outputs(1656) <= b and not a;
    layer3_outputs(1657) <= a and b;
    layer3_outputs(1658) <= '1';
    layer3_outputs(1659) <= '1';
    layer3_outputs(1660) <= a and not b;
    layer3_outputs(1661) <= not b or a;
    layer3_outputs(1662) <= b and not a;
    layer3_outputs(1663) <= '1';
    layer3_outputs(1664) <= not (a or b);
    layer3_outputs(1665) <= b;
    layer3_outputs(1666) <= b and not a;
    layer3_outputs(1667) <= a and not b;
    layer3_outputs(1668) <= not b or a;
    layer3_outputs(1669) <= a or b;
    layer3_outputs(1670) <= '1';
    layer3_outputs(1671) <= not (a and b);
    layer3_outputs(1672) <= a and b;
    layer3_outputs(1673) <= not b;
    layer3_outputs(1674) <= a and b;
    layer3_outputs(1675) <= a and not b;
    layer3_outputs(1676) <= a and not b;
    layer3_outputs(1677) <= a and not b;
    layer3_outputs(1678) <= not (a and b);
    layer3_outputs(1679) <= not b or a;
    layer3_outputs(1680) <= not b or a;
    layer3_outputs(1681) <= a or b;
    layer3_outputs(1682) <= a xor b;
    layer3_outputs(1683) <= b;
    layer3_outputs(1684) <= not b or a;
    layer3_outputs(1685) <= not (a xor b);
    layer3_outputs(1686) <= not a;
    layer3_outputs(1687) <= not a or b;
    layer3_outputs(1688) <= not (a or b);
    layer3_outputs(1689) <= a xor b;
    layer3_outputs(1690) <= a and b;
    layer3_outputs(1691) <= b and not a;
    layer3_outputs(1692) <= '1';
    layer3_outputs(1693) <= not a or b;
    layer3_outputs(1694) <= not b;
    layer3_outputs(1695) <= a and b;
    layer3_outputs(1696) <= not b or a;
    layer3_outputs(1697) <= not (a and b);
    layer3_outputs(1698) <= b;
    layer3_outputs(1699) <= not b or a;
    layer3_outputs(1700) <= b;
    layer3_outputs(1701) <= a and not b;
    layer3_outputs(1702) <= '1';
    layer3_outputs(1703) <= a or b;
    layer3_outputs(1704) <= a xor b;
    layer3_outputs(1705) <= a and b;
    layer3_outputs(1706) <= not (a or b);
    layer3_outputs(1707) <= b and not a;
    layer3_outputs(1708) <= not b;
    layer3_outputs(1709) <= b;
    layer3_outputs(1710) <= b and not a;
    layer3_outputs(1711) <= a and b;
    layer3_outputs(1712) <= not b;
    layer3_outputs(1713) <= a and not b;
    layer3_outputs(1714) <= '0';
    layer3_outputs(1715) <= not b;
    layer3_outputs(1716) <= a;
    layer3_outputs(1717) <= a and b;
    layer3_outputs(1718) <= not b or a;
    layer3_outputs(1719) <= b and not a;
    layer3_outputs(1720) <= b and not a;
    layer3_outputs(1721) <= not b or a;
    layer3_outputs(1722) <= not (a or b);
    layer3_outputs(1723) <= a and b;
    layer3_outputs(1724) <= a and b;
    layer3_outputs(1725) <= '0';
    layer3_outputs(1726) <= not a or b;
    layer3_outputs(1727) <= b and not a;
    layer3_outputs(1728) <= not b;
    layer3_outputs(1729) <= '1';
    layer3_outputs(1730) <= a and not b;
    layer3_outputs(1731) <= a;
    layer3_outputs(1732) <= '1';
    layer3_outputs(1733) <= not b or a;
    layer3_outputs(1734) <= not a or b;
    layer3_outputs(1735) <= a and b;
    layer3_outputs(1736) <= not a;
    layer3_outputs(1737) <= not b;
    layer3_outputs(1738) <= not a or b;
    layer3_outputs(1739) <= b and not a;
    layer3_outputs(1740) <= b;
    layer3_outputs(1741) <= not (a or b);
    layer3_outputs(1742) <= not b or a;
    layer3_outputs(1743) <= not a or b;
    layer3_outputs(1744) <= not a;
    layer3_outputs(1745) <= not (a xor b);
    layer3_outputs(1746) <= a and not b;
    layer3_outputs(1747) <= '1';
    layer3_outputs(1748) <= b;
    layer3_outputs(1749) <= not (a and b);
    layer3_outputs(1750) <= b and not a;
    layer3_outputs(1751) <= '0';
    layer3_outputs(1752) <= not a;
    layer3_outputs(1753) <= a and not b;
    layer3_outputs(1754) <= '0';
    layer3_outputs(1755) <= a and b;
    layer3_outputs(1756) <= a and not b;
    layer3_outputs(1757) <= '1';
    layer3_outputs(1758) <= a;
    layer3_outputs(1759) <= not (a and b);
    layer3_outputs(1760) <= a or b;
    layer3_outputs(1761) <= not b;
    layer3_outputs(1762) <= not a or b;
    layer3_outputs(1763) <= not (a and b);
    layer3_outputs(1764) <= a;
    layer3_outputs(1765) <= a or b;
    layer3_outputs(1766) <= '0';
    layer3_outputs(1767) <= not (a and b);
    layer3_outputs(1768) <= not b or a;
    layer3_outputs(1769) <= not (a and b);
    layer3_outputs(1770) <= '1';
    layer3_outputs(1771) <= not (a or b);
    layer3_outputs(1772) <= '0';
    layer3_outputs(1773) <= a xor b;
    layer3_outputs(1774) <= a and b;
    layer3_outputs(1775) <= a and b;
    layer3_outputs(1776) <= a and b;
    layer3_outputs(1777) <= not (a or b);
    layer3_outputs(1778) <= not b;
    layer3_outputs(1779) <= a xor b;
    layer3_outputs(1780) <= a and not b;
    layer3_outputs(1781) <= '1';
    layer3_outputs(1782) <= a and b;
    layer3_outputs(1783) <= '0';
    layer3_outputs(1784) <= not (a or b);
    layer3_outputs(1785) <= not b;
    layer3_outputs(1786) <= '0';
    layer3_outputs(1787) <= a and not b;
    layer3_outputs(1788) <= not a or b;
    layer3_outputs(1789) <= a xor b;
    layer3_outputs(1790) <= not a;
    layer3_outputs(1791) <= '0';
    layer3_outputs(1792) <= b;
    layer3_outputs(1793) <= not a;
    layer3_outputs(1794) <= not a or b;
    layer3_outputs(1795) <= a and b;
    layer3_outputs(1796) <= b;
    layer3_outputs(1797) <= a and not b;
    layer3_outputs(1798) <= '1';
    layer3_outputs(1799) <= not a;
    layer3_outputs(1800) <= not a;
    layer3_outputs(1801) <= not a or b;
    layer3_outputs(1802) <= a;
    layer3_outputs(1803) <= a;
    layer3_outputs(1804) <= a and b;
    layer3_outputs(1805) <= not b;
    layer3_outputs(1806) <= not b or a;
    layer3_outputs(1807) <= a and not b;
    layer3_outputs(1808) <= not a or b;
    layer3_outputs(1809) <= not b;
    layer3_outputs(1810) <= a;
    layer3_outputs(1811) <= not (a and b);
    layer3_outputs(1812) <= '1';
    layer3_outputs(1813) <= not a;
    layer3_outputs(1814) <= a or b;
    layer3_outputs(1815) <= '1';
    layer3_outputs(1816) <= a and b;
    layer3_outputs(1817) <= b and not a;
    layer3_outputs(1818) <= not (a or b);
    layer3_outputs(1819) <= '1';
    layer3_outputs(1820) <= '1';
    layer3_outputs(1821) <= not (a or b);
    layer3_outputs(1822) <= a xor b;
    layer3_outputs(1823) <= not a;
    layer3_outputs(1824) <= a and not b;
    layer3_outputs(1825) <= not (a and b);
    layer3_outputs(1826) <= not a;
    layer3_outputs(1827) <= b and not a;
    layer3_outputs(1828) <= '1';
    layer3_outputs(1829) <= '1';
    layer3_outputs(1830) <= not b or a;
    layer3_outputs(1831) <= '1';
    layer3_outputs(1832) <= '0';
    layer3_outputs(1833) <= not b;
    layer3_outputs(1834) <= not a;
    layer3_outputs(1835) <= not a;
    layer3_outputs(1836) <= not a or b;
    layer3_outputs(1837) <= b;
    layer3_outputs(1838) <= '1';
    layer3_outputs(1839) <= not a;
    layer3_outputs(1840) <= a or b;
    layer3_outputs(1841) <= not b;
    layer3_outputs(1842) <= b;
    layer3_outputs(1843) <= not b or a;
    layer3_outputs(1844) <= '1';
    layer3_outputs(1845) <= not b;
    layer3_outputs(1846) <= a and b;
    layer3_outputs(1847) <= not (a and b);
    layer3_outputs(1848) <= '1';
    layer3_outputs(1849) <= a and b;
    layer3_outputs(1850) <= a and b;
    layer3_outputs(1851) <= a;
    layer3_outputs(1852) <= not a;
    layer3_outputs(1853) <= not (a and b);
    layer3_outputs(1854) <= not a;
    layer3_outputs(1855) <= a or b;
    layer3_outputs(1856) <= '0';
    layer3_outputs(1857) <= a or b;
    layer3_outputs(1858) <= a and not b;
    layer3_outputs(1859) <= not b;
    layer3_outputs(1860) <= b and not a;
    layer3_outputs(1861) <= a;
    layer3_outputs(1862) <= not a or b;
    layer3_outputs(1863) <= a;
    layer3_outputs(1864) <= '0';
    layer3_outputs(1865) <= a and not b;
    layer3_outputs(1866) <= '1';
    layer3_outputs(1867) <= not a;
    layer3_outputs(1868) <= a xor b;
    layer3_outputs(1869) <= not a;
    layer3_outputs(1870) <= not b;
    layer3_outputs(1871) <= a and b;
    layer3_outputs(1872) <= not a;
    layer3_outputs(1873) <= not b;
    layer3_outputs(1874) <= not b;
    layer3_outputs(1875) <= a and b;
    layer3_outputs(1876) <= not (a and b);
    layer3_outputs(1877) <= '0';
    layer3_outputs(1878) <= not a;
    layer3_outputs(1879) <= a;
    layer3_outputs(1880) <= a;
    layer3_outputs(1881) <= a and not b;
    layer3_outputs(1882) <= '0';
    layer3_outputs(1883) <= not (a xor b);
    layer3_outputs(1884) <= not (a or b);
    layer3_outputs(1885) <= b and not a;
    layer3_outputs(1886) <= b and not a;
    layer3_outputs(1887) <= a and b;
    layer3_outputs(1888) <= not (a or b);
    layer3_outputs(1889) <= '0';
    layer3_outputs(1890) <= '0';
    layer3_outputs(1891) <= a and not b;
    layer3_outputs(1892) <= '0';
    layer3_outputs(1893) <= b and not a;
    layer3_outputs(1894) <= b and not a;
    layer3_outputs(1895) <= b and not a;
    layer3_outputs(1896) <= not b or a;
    layer3_outputs(1897) <= a and b;
    layer3_outputs(1898) <= not (a xor b);
    layer3_outputs(1899) <= not a or b;
    layer3_outputs(1900) <= a;
    layer3_outputs(1901) <= b;
    layer3_outputs(1902) <= '1';
    layer3_outputs(1903) <= not b;
    layer3_outputs(1904) <= not a;
    layer3_outputs(1905) <= not b or a;
    layer3_outputs(1906) <= b;
    layer3_outputs(1907) <= b;
    layer3_outputs(1908) <= a and not b;
    layer3_outputs(1909) <= '0';
    layer3_outputs(1910) <= a;
    layer3_outputs(1911) <= '0';
    layer3_outputs(1912) <= not (a or b);
    layer3_outputs(1913) <= not a;
    layer3_outputs(1914) <= not (a or b);
    layer3_outputs(1915) <= a and not b;
    layer3_outputs(1916) <= not (a xor b);
    layer3_outputs(1917) <= '1';
    layer3_outputs(1918) <= not (a or b);
    layer3_outputs(1919) <= not b or a;
    layer3_outputs(1920) <= a;
    layer3_outputs(1921) <= a and b;
    layer3_outputs(1922) <= a or b;
    layer3_outputs(1923) <= a xor b;
    layer3_outputs(1924) <= not b;
    layer3_outputs(1925) <= a or b;
    layer3_outputs(1926) <= '0';
    layer3_outputs(1927) <= not (a and b);
    layer3_outputs(1928) <= b;
    layer3_outputs(1929) <= a;
    layer3_outputs(1930) <= a or b;
    layer3_outputs(1931) <= not b;
    layer3_outputs(1932) <= '1';
    layer3_outputs(1933) <= '1';
    layer3_outputs(1934) <= not (a and b);
    layer3_outputs(1935) <= a and b;
    layer3_outputs(1936) <= a and not b;
    layer3_outputs(1937) <= '1';
    layer3_outputs(1938) <= '0';
    layer3_outputs(1939) <= '0';
    layer3_outputs(1940) <= '1';
    layer3_outputs(1941) <= not a or b;
    layer3_outputs(1942) <= not b or a;
    layer3_outputs(1943) <= not b or a;
    layer3_outputs(1944) <= b and not a;
    layer3_outputs(1945) <= not a or b;
    layer3_outputs(1946) <= b;
    layer3_outputs(1947) <= not a or b;
    layer3_outputs(1948) <= not (a or b);
    layer3_outputs(1949) <= not b;
    layer3_outputs(1950) <= '1';
    layer3_outputs(1951) <= a xor b;
    layer3_outputs(1952) <= b;
    layer3_outputs(1953) <= '0';
    layer3_outputs(1954) <= not b;
    layer3_outputs(1955) <= '0';
    layer3_outputs(1956) <= not (a and b);
    layer3_outputs(1957) <= '0';
    layer3_outputs(1958) <= a and b;
    layer3_outputs(1959) <= not a;
    layer3_outputs(1960) <= not b or a;
    layer3_outputs(1961) <= a;
    layer3_outputs(1962) <= not b or a;
    layer3_outputs(1963) <= '1';
    layer3_outputs(1964) <= '0';
    layer3_outputs(1965) <= not (a xor b);
    layer3_outputs(1966) <= not (a xor b);
    layer3_outputs(1967) <= b;
    layer3_outputs(1968) <= a and not b;
    layer3_outputs(1969) <= b;
    layer3_outputs(1970) <= '1';
    layer3_outputs(1971) <= not (a or b);
    layer3_outputs(1972) <= '1';
    layer3_outputs(1973) <= a and not b;
    layer3_outputs(1974) <= a and not b;
    layer3_outputs(1975) <= a xor b;
    layer3_outputs(1976) <= not (a and b);
    layer3_outputs(1977) <= '0';
    layer3_outputs(1978) <= not (a and b);
    layer3_outputs(1979) <= not b or a;
    layer3_outputs(1980) <= not b or a;
    layer3_outputs(1981) <= not (a xor b);
    layer3_outputs(1982) <= a;
    layer3_outputs(1983) <= a;
    layer3_outputs(1984) <= a and b;
    layer3_outputs(1985) <= a xor b;
    layer3_outputs(1986) <= '0';
    layer3_outputs(1987) <= not b;
    layer3_outputs(1988) <= not b;
    layer3_outputs(1989) <= not (a and b);
    layer3_outputs(1990) <= not a or b;
    layer3_outputs(1991) <= not a;
    layer3_outputs(1992) <= b and not a;
    layer3_outputs(1993) <= a or b;
    layer3_outputs(1994) <= a and not b;
    layer3_outputs(1995) <= not b or a;
    layer3_outputs(1996) <= '0';
    layer3_outputs(1997) <= b;
    layer3_outputs(1998) <= a and b;
    layer3_outputs(1999) <= not (a or b);
    layer3_outputs(2000) <= not (a and b);
    layer3_outputs(2001) <= '0';
    layer3_outputs(2002) <= '0';
    layer3_outputs(2003) <= a or b;
    layer3_outputs(2004) <= b and not a;
    layer3_outputs(2005) <= a and not b;
    layer3_outputs(2006) <= not b;
    layer3_outputs(2007) <= a and b;
    layer3_outputs(2008) <= not b;
    layer3_outputs(2009) <= '1';
    layer3_outputs(2010) <= '0';
    layer3_outputs(2011) <= b;
    layer3_outputs(2012) <= b and not a;
    layer3_outputs(2013) <= b;
    layer3_outputs(2014) <= a or b;
    layer3_outputs(2015) <= not b;
    layer3_outputs(2016) <= b;
    layer3_outputs(2017) <= not (a and b);
    layer3_outputs(2018) <= not a or b;
    layer3_outputs(2019) <= not (a and b);
    layer3_outputs(2020) <= not (a xor b);
    layer3_outputs(2021) <= a and not b;
    layer3_outputs(2022) <= b and not a;
    layer3_outputs(2023) <= not a or b;
    layer3_outputs(2024) <= '1';
    layer3_outputs(2025) <= not a or b;
    layer3_outputs(2026) <= a and b;
    layer3_outputs(2027) <= not b or a;
    layer3_outputs(2028) <= not a or b;
    layer3_outputs(2029) <= a;
    layer3_outputs(2030) <= '0';
    layer3_outputs(2031) <= '1';
    layer3_outputs(2032) <= a or b;
    layer3_outputs(2033) <= a;
    layer3_outputs(2034) <= b;
    layer3_outputs(2035) <= '1';
    layer3_outputs(2036) <= '0';
    layer3_outputs(2037) <= not a;
    layer3_outputs(2038) <= '1';
    layer3_outputs(2039) <= a;
    layer3_outputs(2040) <= '1';
    layer3_outputs(2041) <= b;
    layer3_outputs(2042) <= not a;
    layer3_outputs(2043) <= not (a or b);
    layer3_outputs(2044) <= '1';
    layer3_outputs(2045) <= a;
    layer3_outputs(2046) <= '1';
    layer3_outputs(2047) <= b and not a;
    layer3_outputs(2048) <= b and not a;
    layer3_outputs(2049) <= a and b;
    layer3_outputs(2050) <= a and not b;
    layer3_outputs(2051) <= a or b;
    layer3_outputs(2052) <= not (a or b);
    layer3_outputs(2053) <= '0';
    layer3_outputs(2054) <= not b;
    layer3_outputs(2055) <= '1';
    layer3_outputs(2056) <= '0';
    layer3_outputs(2057) <= not (a and b);
    layer3_outputs(2058) <= '0';
    layer3_outputs(2059) <= b;
    layer3_outputs(2060) <= b and not a;
    layer3_outputs(2061) <= a or b;
    layer3_outputs(2062) <= not a or b;
    layer3_outputs(2063) <= not a;
    layer3_outputs(2064) <= '1';
    layer3_outputs(2065) <= not a;
    layer3_outputs(2066) <= '1';
    layer3_outputs(2067) <= not b;
    layer3_outputs(2068) <= '0';
    layer3_outputs(2069) <= '0';
    layer3_outputs(2070) <= '1';
    layer3_outputs(2071) <= a and not b;
    layer3_outputs(2072) <= b and not a;
    layer3_outputs(2073) <= a;
    layer3_outputs(2074) <= '1';
    layer3_outputs(2075) <= not (a or b);
    layer3_outputs(2076) <= '0';
    layer3_outputs(2077) <= not b or a;
    layer3_outputs(2078) <= a or b;
    layer3_outputs(2079) <= not a;
    layer3_outputs(2080) <= a and b;
    layer3_outputs(2081) <= b and not a;
    layer3_outputs(2082) <= b;
    layer3_outputs(2083) <= not b;
    layer3_outputs(2084) <= not a or b;
    layer3_outputs(2085) <= b and not a;
    layer3_outputs(2086) <= not (a xor b);
    layer3_outputs(2087) <= a and not b;
    layer3_outputs(2088) <= '0';
    layer3_outputs(2089) <= not (a and b);
    layer3_outputs(2090) <= not (a or b);
    layer3_outputs(2091) <= not (a or b);
    layer3_outputs(2092) <= not a;
    layer3_outputs(2093) <= '1';
    layer3_outputs(2094) <= '0';
    layer3_outputs(2095) <= not b;
    layer3_outputs(2096) <= not a or b;
    layer3_outputs(2097) <= a or b;
    layer3_outputs(2098) <= '1';
    layer3_outputs(2099) <= not (a xor b);
    layer3_outputs(2100) <= '0';
    layer3_outputs(2101) <= not (a and b);
    layer3_outputs(2102) <= not (a and b);
    layer3_outputs(2103) <= a or b;
    layer3_outputs(2104) <= not (a and b);
    layer3_outputs(2105) <= a or b;
    layer3_outputs(2106) <= a or b;
    layer3_outputs(2107) <= b;
    layer3_outputs(2108) <= '1';
    layer3_outputs(2109) <= not (a xor b);
    layer3_outputs(2110) <= '1';
    layer3_outputs(2111) <= a or b;
    layer3_outputs(2112) <= '0';
    layer3_outputs(2113) <= b;
    layer3_outputs(2114) <= not (a or b);
    layer3_outputs(2115) <= not (a and b);
    layer3_outputs(2116) <= '1';
    layer3_outputs(2117) <= not b or a;
    layer3_outputs(2118) <= a or b;
    layer3_outputs(2119) <= not (a or b);
    layer3_outputs(2120) <= b;
    layer3_outputs(2121) <= not (a xor b);
    layer3_outputs(2122) <= '1';
    layer3_outputs(2123) <= not a;
    layer3_outputs(2124) <= not (a or b);
    layer3_outputs(2125) <= not (a xor b);
    layer3_outputs(2126) <= a or b;
    layer3_outputs(2127) <= '0';
    layer3_outputs(2128) <= a;
    layer3_outputs(2129) <= '0';
    layer3_outputs(2130) <= a and not b;
    layer3_outputs(2131) <= a and not b;
    layer3_outputs(2132) <= a and b;
    layer3_outputs(2133) <= not a;
    layer3_outputs(2134) <= not a;
    layer3_outputs(2135) <= a and not b;
    layer3_outputs(2136) <= b and not a;
    layer3_outputs(2137) <= a or b;
    layer3_outputs(2138) <= not (a and b);
    layer3_outputs(2139) <= '0';
    layer3_outputs(2140) <= a or b;
    layer3_outputs(2141) <= '0';
    layer3_outputs(2142) <= not (a and b);
    layer3_outputs(2143) <= b and not a;
    layer3_outputs(2144) <= a;
    layer3_outputs(2145) <= a and not b;
    layer3_outputs(2146) <= not a or b;
    layer3_outputs(2147) <= not (a and b);
    layer3_outputs(2148) <= not b;
    layer3_outputs(2149) <= a;
    layer3_outputs(2150) <= '0';
    layer3_outputs(2151) <= '1';
    layer3_outputs(2152) <= b and not a;
    layer3_outputs(2153) <= not (a xor b);
    layer3_outputs(2154) <= not a;
    layer3_outputs(2155) <= not (a or b);
    layer3_outputs(2156) <= not a or b;
    layer3_outputs(2157) <= not b;
    layer3_outputs(2158) <= '1';
    layer3_outputs(2159) <= '1';
    layer3_outputs(2160) <= a or b;
    layer3_outputs(2161) <= b and not a;
    layer3_outputs(2162) <= a or b;
    layer3_outputs(2163) <= not b or a;
    layer3_outputs(2164) <= '0';
    layer3_outputs(2165) <= b;
    layer3_outputs(2166) <= not a;
    layer3_outputs(2167) <= b;
    layer3_outputs(2168) <= a;
    layer3_outputs(2169) <= b and not a;
    layer3_outputs(2170) <= a and not b;
    layer3_outputs(2171) <= not b or a;
    layer3_outputs(2172) <= not (a and b);
    layer3_outputs(2173) <= a and b;
    layer3_outputs(2174) <= a;
    layer3_outputs(2175) <= b;
    layer3_outputs(2176) <= not (a and b);
    layer3_outputs(2177) <= '1';
    layer3_outputs(2178) <= not (a or b);
    layer3_outputs(2179) <= not (a or b);
    layer3_outputs(2180) <= '0';
    layer3_outputs(2181) <= not (a xor b);
    layer3_outputs(2182) <= '1';
    layer3_outputs(2183) <= not (a and b);
    layer3_outputs(2184) <= b;
    layer3_outputs(2185) <= not b;
    layer3_outputs(2186) <= '0';
    layer3_outputs(2187) <= b and not a;
    layer3_outputs(2188) <= not b;
    layer3_outputs(2189) <= b;
    layer3_outputs(2190) <= not b or a;
    layer3_outputs(2191) <= not (a or b);
    layer3_outputs(2192) <= a and not b;
    layer3_outputs(2193) <= a and not b;
    layer3_outputs(2194) <= a and not b;
    layer3_outputs(2195) <= a or b;
    layer3_outputs(2196) <= not a;
    layer3_outputs(2197) <= not (a and b);
    layer3_outputs(2198) <= '1';
    layer3_outputs(2199) <= not (a or b);
    layer3_outputs(2200) <= b and not a;
    layer3_outputs(2201) <= not (a or b);
    layer3_outputs(2202) <= not (a and b);
    layer3_outputs(2203) <= not (a or b);
    layer3_outputs(2204) <= not (a and b);
    layer3_outputs(2205) <= not (a and b);
    layer3_outputs(2206) <= not b or a;
    layer3_outputs(2207) <= not b or a;
    layer3_outputs(2208) <= a or b;
    layer3_outputs(2209) <= '1';
    layer3_outputs(2210) <= b;
    layer3_outputs(2211) <= a and not b;
    layer3_outputs(2212) <= not (a and b);
    layer3_outputs(2213) <= '0';
    layer3_outputs(2214) <= a and b;
    layer3_outputs(2215) <= '0';
    layer3_outputs(2216) <= a and b;
    layer3_outputs(2217) <= not b or a;
    layer3_outputs(2218) <= not (a and b);
    layer3_outputs(2219) <= a or b;
    layer3_outputs(2220) <= not b or a;
    layer3_outputs(2221) <= '1';
    layer3_outputs(2222) <= a or b;
    layer3_outputs(2223) <= not b;
    layer3_outputs(2224) <= a and not b;
    layer3_outputs(2225) <= b and not a;
    layer3_outputs(2226) <= not (a and b);
    layer3_outputs(2227) <= '0';
    layer3_outputs(2228) <= '1';
    layer3_outputs(2229) <= not b;
    layer3_outputs(2230) <= not b;
    layer3_outputs(2231) <= not (a or b);
    layer3_outputs(2232) <= a;
    layer3_outputs(2233) <= '1';
    layer3_outputs(2234) <= not a;
    layer3_outputs(2235) <= a or b;
    layer3_outputs(2236) <= not (a and b);
    layer3_outputs(2237) <= a and b;
    layer3_outputs(2238) <= not (a xor b);
    layer3_outputs(2239) <= not (a or b);
    layer3_outputs(2240) <= a and not b;
    layer3_outputs(2241) <= not b;
    layer3_outputs(2242) <= a or b;
    layer3_outputs(2243) <= not (a and b);
    layer3_outputs(2244) <= not (a and b);
    layer3_outputs(2245) <= not b or a;
    layer3_outputs(2246) <= a;
    layer3_outputs(2247) <= b;
    layer3_outputs(2248) <= a and b;
    layer3_outputs(2249) <= b and not a;
    layer3_outputs(2250) <= not b;
    layer3_outputs(2251) <= a and b;
    layer3_outputs(2252) <= '1';
    layer3_outputs(2253) <= '0';
    layer3_outputs(2254) <= not (a or b);
    layer3_outputs(2255) <= '0';
    layer3_outputs(2256) <= not b or a;
    layer3_outputs(2257) <= not b;
    layer3_outputs(2258) <= b and not a;
    layer3_outputs(2259) <= a or b;
    layer3_outputs(2260) <= a or b;
    layer3_outputs(2261) <= not (a or b);
    layer3_outputs(2262) <= not a;
    layer3_outputs(2263) <= not (a and b);
    layer3_outputs(2264) <= '0';
    layer3_outputs(2265) <= a xor b;
    layer3_outputs(2266) <= a and b;
    layer3_outputs(2267) <= not (a or b);
    layer3_outputs(2268) <= not a or b;
    layer3_outputs(2269) <= not (a xor b);
    layer3_outputs(2270) <= not b;
    layer3_outputs(2271) <= not (a xor b);
    layer3_outputs(2272) <= not (a and b);
    layer3_outputs(2273) <= not a or b;
    layer3_outputs(2274) <= '1';
    layer3_outputs(2275) <= b and not a;
    layer3_outputs(2276) <= not (a or b);
    layer3_outputs(2277) <= not (a and b);
    layer3_outputs(2278) <= not (a or b);
    layer3_outputs(2279) <= b;
    layer3_outputs(2280) <= a and not b;
    layer3_outputs(2281) <= b and not a;
    layer3_outputs(2282) <= not a or b;
    layer3_outputs(2283) <= not (a and b);
    layer3_outputs(2284) <= b and not a;
    layer3_outputs(2285) <= not b or a;
    layer3_outputs(2286) <= '1';
    layer3_outputs(2287) <= a and b;
    layer3_outputs(2288) <= a and not b;
    layer3_outputs(2289) <= a and b;
    layer3_outputs(2290) <= a and not b;
    layer3_outputs(2291) <= not a;
    layer3_outputs(2292) <= not b;
    layer3_outputs(2293) <= a or b;
    layer3_outputs(2294) <= not (a and b);
    layer3_outputs(2295) <= a;
    layer3_outputs(2296) <= not b or a;
    layer3_outputs(2297) <= not (a xor b);
    layer3_outputs(2298) <= a and b;
    layer3_outputs(2299) <= '1';
    layer3_outputs(2300) <= not (a or b);
    layer3_outputs(2301) <= a and not b;
    layer3_outputs(2302) <= b and not a;
    layer3_outputs(2303) <= b and not a;
    layer3_outputs(2304) <= a or b;
    layer3_outputs(2305) <= not a or b;
    layer3_outputs(2306) <= not a or b;
    layer3_outputs(2307) <= not b;
    layer3_outputs(2308) <= b and not a;
    layer3_outputs(2309) <= not b;
    layer3_outputs(2310) <= not (a and b);
    layer3_outputs(2311) <= a and not b;
    layer3_outputs(2312) <= b and not a;
    layer3_outputs(2313) <= a;
    layer3_outputs(2314) <= not b or a;
    layer3_outputs(2315) <= '1';
    layer3_outputs(2316) <= a and b;
    layer3_outputs(2317) <= '0';
    layer3_outputs(2318) <= not b;
    layer3_outputs(2319) <= not a or b;
    layer3_outputs(2320) <= '1';
    layer3_outputs(2321) <= a and b;
    layer3_outputs(2322) <= not b or a;
    layer3_outputs(2323) <= '1';
    layer3_outputs(2324) <= not a;
    layer3_outputs(2325) <= a or b;
    layer3_outputs(2326) <= not b;
    layer3_outputs(2327) <= a and b;
    layer3_outputs(2328) <= not a or b;
    layer3_outputs(2329) <= a and b;
    layer3_outputs(2330) <= not (a or b);
    layer3_outputs(2331) <= not (a or b);
    layer3_outputs(2332) <= a and not b;
    layer3_outputs(2333) <= '1';
    layer3_outputs(2334) <= '0';
    layer3_outputs(2335) <= '1';
    layer3_outputs(2336) <= not b or a;
    layer3_outputs(2337) <= not a;
    layer3_outputs(2338) <= not (a and b);
    layer3_outputs(2339) <= not b;
    layer3_outputs(2340) <= not a or b;
    layer3_outputs(2341) <= a xor b;
    layer3_outputs(2342) <= '0';
    layer3_outputs(2343) <= '1';
    layer3_outputs(2344) <= b;
    layer3_outputs(2345) <= a;
    layer3_outputs(2346) <= a or b;
    layer3_outputs(2347) <= not b or a;
    layer3_outputs(2348) <= b;
    layer3_outputs(2349) <= not b;
    layer3_outputs(2350) <= a;
    layer3_outputs(2351) <= not (a and b);
    layer3_outputs(2352) <= not (a or b);
    layer3_outputs(2353) <= not a;
    layer3_outputs(2354) <= not b;
    layer3_outputs(2355) <= a and b;
    layer3_outputs(2356) <= a;
    layer3_outputs(2357) <= '1';
    layer3_outputs(2358) <= not (a and b);
    layer3_outputs(2359) <= b;
    layer3_outputs(2360) <= a or b;
    layer3_outputs(2361) <= not (a and b);
    layer3_outputs(2362) <= not b;
    layer3_outputs(2363) <= b;
    layer3_outputs(2364) <= not (a or b);
    layer3_outputs(2365) <= not (a and b);
    layer3_outputs(2366) <= a xor b;
    layer3_outputs(2367) <= not a;
    layer3_outputs(2368) <= not b;
    layer3_outputs(2369) <= a and not b;
    layer3_outputs(2370) <= a and b;
    layer3_outputs(2371) <= '1';
    layer3_outputs(2372) <= a and b;
    layer3_outputs(2373) <= not (a and b);
    layer3_outputs(2374) <= '0';
    layer3_outputs(2375) <= a or b;
    layer3_outputs(2376) <= not (a or b);
    layer3_outputs(2377) <= not b or a;
    layer3_outputs(2378) <= a or b;
    layer3_outputs(2379) <= not (a and b);
    layer3_outputs(2380) <= not a;
    layer3_outputs(2381) <= b and not a;
    layer3_outputs(2382) <= not b or a;
    layer3_outputs(2383) <= not a or b;
    layer3_outputs(2384) <= '1';
    layer3_outputs(2385) <= a and b;
    layer3_outputs(2386) <= a or b;
    layer3_outputs(2387) <= not b;
    layer3_outputs(2388) <= not b;
    layer3_outputs(2389) <= not (a or b);
    layer3_outputs(2390) <= not b;
    layer3_outputs(2391) <= a and b;
    layer3_outputs(2392) <= a or b;
    layer3_outputs(2393) <= '0';
    layer3_outputs(2394) <= not (a and b);
    layer3_outputs(2395) <= '1';
    layer3_outputs(2396) <= not a or b;
    layer3_outputs(2397) <= not (a and b);
    layer3_outputs(2398) <= b and not a;
    layer3_outputs(2399) <= a or b;
    layer3_outputs(2400) <= not a;
    layer3_outputs(2401) <= a;
    layer3_outputs(2402) <= not (a or b);
    layer3_outputs(2403) <= not a or b;
    layer3_outputs(2404) <= b;
    layer3_outputs(2405) <= b;
    layer3_outputs(2406) <= b and not a;
    layer3_outputs(2407) <= a and b;
    layer3_outputs(2408) <= not (a and b);
    layer3_outputs(2409) <= b;
    layer3_outputs(2410) <= a or b;
    layer3_outputs(2411) <= not (a and b);
    layer3_outputs(2412) <= not a;
    layer3_outputs(2413) <= a xor b;
    layer3_outputs(2414) <= a and b;
    layer3_outputs(2415) <= not a or b;
    layer3_outputs(2416) <= not b or a;
    layer3_outputs(2417) <= not a or b;
    layer3_outputs(2418) <= not b or a;
    layer3_outputs(2419) <= b and not a;
    layer3_outputs(2420) <= b and not a;
    layer3_outputs(2421) <= a;
    layer3_outputs(2422) <= '1';
    layer3_outputs(2423) <= b and not a;
    layer3_outputs(2424) <= not a;
    layer3_outputs(2425) <= '0';
    layer3_outputs(2426) <= a and not b;
    layer3_outputs(2427) <= b;
    layer3_outputs(2428) <= a and b;
    layer3_outputs(2429) <= a and b;
    layer3_outputs(2430) <= b and not a;
    layer3_outputs(2431) <= a and b;
    layer3_outputs(2432) <= '0';
    layer3_outputs(2433) <= not b;
    layer3_outputs(2434) <= '1';
    layer3_outputs(2435) <= not a;
    layer3_outputs(2436) <= a;
    layer3_outputs(2437) <= not b;
    layer3_outputs(2438) <= not (a or b);
    layer3_outputs(2439) <= not a;
    layer3_outputs(2440) <= '0';
    layer3_outputs(2441) <= a or b;
    layer3_outputs(2442) <= not b or a;
    layer3_outputs(2443) <= not a or b;
    layer3_outputs(2444) <= not b or a;
    layer3_outputs(2445) <= not b or a;
    layer3_outputs(2446) <= not a or b;
    layer3_outputs(2447) <= not a or b;
    layer3_outputs(2448) <= not b or a;
    layer3_outputs(2449) <= not b;
    layer3_outputs(2450) <= not b or a;
    layer3_outputs(2451) <= '0';
    layer3_outputs(2452) <= not (a and b);
    layer3_outputs(2453) <= b;
    layer3_outputs(2454) <= not (a and b);
    layer3_outputs(2455) <= not a or b;
    layer3_outputs(2456) <= b and not a;
    layer3_outputs(2457) <= a and b;
    layer3_outputs(2458) <= b and not a;
    layer3_outputs(2459) <= a or b;
    layer3_outputs(2460) <= '1';
    layer3_outputs(2461) <= a;
    layer3_outputs(2462) <= not (a or b);
    layer3_outputs(2463) <= b and not a;
    layer3_outputs(2464) <= '1';
    layer3_outputs(2465) <= '1';
    layer3_outputs(2466) <= b and not a;
    layer3_outputs(2467) <= '0';
    layer3_outputs(2468) <= not (a or b);
    layer3_outputs(2469) <= not b;
    layer3_outputs(2470) <= a and b;
    layer3_outputs(2471) <= a and b;
    layer3_outputs(2472) <= not a;
    layer3_outputs(2473) <= not b or a;
    layer3_outputs(2474) <= a;
    layer3_outputs(2475) <= not a or b;
    layer3_outputs(2476) <= not a or b;
    layer3_outputs(2477) <= not (a or b);
    layer3_outputs(2478) <= a;
    layer3_outputs(2479) <= not b or a;
    layer3_outputs(2480) <= not a;
    layer3_outputs(2481) <= '0';
    layer3_outputs(2482) <= not (a or b);
    layer3_outputs(2483) <= not a or b;
    layer3_outputs(2484) <= a;
    layer3_outputs(2485) <= a and not b;
    layer3_outputs(2486) <= '1';
    layer3_outputs(2487) <= not a;
    layer3_outputs(2488) <= not b or a;
    layer3_outputs(2489) <= not (a and b);
    layer3_outputs(2490) <= not (a xor b);
    layer3_outputs(2491) <= b;
    layer3_outputs(2492) <= not (a or b);
    layer3_outputs(2493) <= a and not b;
    layer3_outputs(2494) <= a;
    layer3_outputs(2495) <= '1';
    layer3_outputs(2496) <= not (a and b);
    layer3_outputs(2497) <= not b;
    layer3_outputs(2498) <= not (a xor b);
    layer3_outputs(2499) <= b and not a;
    layer3_outputs(2500) <= '1';
    layer3_outputs(2501) <= a xor b;
    layer3_outputs(2502) <= b and not a;
    layer3_outputs(2503) <= '0';
    layer3_outputs(2504) <= a;
    layer3_outputs(2505) <= not (a and b);
    layer3_outputs(2506) <= '0';
    layer3_outputs(2507) <= '0';
    layer3_outputs(2508) <= a and b;
    layer3_outputs(2509) <= not b or a;
    layer3_outputs(2510) <= '0';
    layer3_outputs(2511) <= not a or b;
    layer3_outputs(2512) <= b;
    layer3_outputs(2513) <= not b or a;
    layer3_outputs(2514) <= not b or a;
    layer3_outputs(2515) <= a or b;
    layer3_outputs(2516) <= b and not a;
    layer3_outputs(2517) <= not a or b;
    layer3_outputs(2518) <= not (a and b);
    layer3_outputs(2519) <= b and not a;
    layer3_outputs(2520) <= not (a and b);
    layer3_outputs(2521) <= '0';
    layer3_outputs(2522) <= b;
    layer3_outputs(2523) <= not b or a;
    layer3_outputs(2524) <= not a;
    layer3_outputs(2525) <= '1';
    layer3_outputs(2526) <= not b;
    layer3_outputs(2527) <= a;
    layer3_outputs(2528) <= '0';
    layer3_outputs(2529) <= not (a or b);
    layer3_outputs(2530) <= not b;
    layer3_outputs(2531) <= '0';
    layer3_outputs(2532) <= '1';
    layer3_outputs(2533) <= not b or a;
    layer3_outputs(2534) <= a or b;
    layer3_outputs(2535) <= '0';
    layer3_outputs(2536) <= not (a and b);
    layer3_outputs(2537) <= not a or b;
    layer3_outputs(2538) <= a;
    layer3_outputs(2539) <= a;
    layer3_outputs(2540) <= a and not b;
    layer3_outputs(2541) <= a and not b;
    layer3_outputs(2542) <= a and b;
    layer3_outputs(2543) <= not (a xor b);
    layer3_outputs(2544) <= b;
    layer3_outputs(2545) <= a and b;
    layer3_outputs(2546) <= b and not a;
    layer3_outputs(2547) <= a or b;
    layer3_outputs(2548) <= not (a or b);
    layer3_outputs(2549) <= a or b;
    layer3_outputs(2550) <= '0';
    layer3_outputs(2551) <= a;
    layer3_outputs(2552) <= not a or b;
    layer3_outputs(2553) <= b;
    layer3_outputs(2554) <= b and not a;
    layer3_outputs(2555) <= a;
    layer3_outputs(2556) <= '0';
    layer3_outputs(2557) <= not a;
    layer3_outputs(2558) <= not (a or b);
    layer3_outputs(2559) <= not b or a;
    layer3_outputs(2560) <= not (a and b);
    layer3_outputs(2561) <= '0';
    layer3_outputs(2562) <= '1';
    layer3_outputs(2563) <= a or b;
    layer3_outputs(2564) <= not (a or b);
    layer3_outputs(2565) <= b;
    layer3_outputs(2566) <= not b;
    layer3_outputs(2567) <= not (a and b);
    layer3_outputs(2568) <= b and not a;
    layer3_outputs(2569) <= a and b;
    layer3_outputs(2570) <= '0';
    layer3_outputs(2571) <= b and not a;
    layer3_outputs(2572) <= '1';
    layer3_outputs(2573) <= not a;
    layer3_outputs(2574) <= not a;
    layer3_outputs(2575) <= b and not a;
    layer3_outputs(2576) <= a or b;
    layer3_outputs(2577) <= b;
    layer3_outputs(2578) <= not b or a;
    layer3_outputs(2579) <= not b;
    layer3_outputs(2580) <= not a or b;
    layer3_outputs(2581) <= not (a or b);
    layer3_outputs(2582) <= a;
    layer3_outputs(2583) <= not b;
    layer3_outputs(2584) <= '1';
    layer3_outputs(2585) <= a or b;
    layer3_outputs(2586) <= not (a and b);
    layer3_outputs(2587) <= a and not b;
    layer3_outputs(2588) <= a and not b;
    layer3_outputs(2589) <= '1';
    layer3_outputs(2590) <= not (a and b);
    layer3_outputs(2591) <= not a or b;
    layer3_outputs(2592) <= a;
    layer3_outputs(2593) <= not b or a;
    layer3_outputs(2594) <= '0';
    layer3_outputs(2595) <= b;
    layer3_outputs(2596) <= not b;
    layer3_outputs(2597) <= a;
    layer3_outputs(2598) <= b;
    layer3_outputs(2599) <= a or b;
    layer3_outputs(2600) <= '1';
    layer3_outputs(2601) <= b and not a;
    layer3_outputs(2602) <= '1';
    layer3_outputs(2603) <= '0';
    layer3_outputs(2604) <= not (a or b);
    layer3_outputs(2605) <= a and b;
    layer3_outputs(2606) <= not (a and b);
    layer3_outputs(2607) <= not (a xor b);
    layer3_outputs(2608) <= a;
    layer3_outputs(2609) <= '0';
    layer3_outputs(2610) <= not b;
    layer3_outputs(2611) <= b and not a;
    layer3_outputs(2612) <= not b;
    layer3_outputs(2613) <= not a or b;
    layer3_outputs(2614) <= b and not a;
    layer3_outputs(2615) <= not b;
    layer3_outputs(2616) <= b and not a;
    layer3_outputs(2617) <= a;
    layer3_outputs(2618) <= not b;
    layer3_outputs(2619) <= '1';
    layer3_outputs(2620) <= not b or a;
    layer3_outputs(2621) <= not a or b;
    layer3_outputs(2622) <= b;
    layer3_outputs(2623) <= not (a or b);
    layer3_outputs(2624) <= a and not b;
    layer3_outputs(2625) <= not a;
    layer3_outputs(2626) <= b and not a;
    layer3_outputs(2627) <= not (a xor b);
    layer3_outputs(2628) <= a and not b;
    layer3_outputs(2629) <= not a;
    layer3_outputs(2630) <= a or b;
    layer3_outputs(2631) <= a;
    layer3_outputs(2632) <= not b;
    layer3_outputs(2633) <= b and not a;
    layer3_outputs(2634) <= not (a or b);
    layer3_outputs(2635) <= a or b;
    layer3_outputs(2636) <= not b or a;
    layer3_outputs(2637) <= a and b;
    layer3_outputs(2638) <= a or b;
    layer3_outputs(2639) <= not a or b;
    layer3_outputs(2640) <= '0';
    layer3_outputs(2641) <= a or b;
    layer3_outputs(2642) <= '1';
    layer3_outputs(2643) <= a;
    layer3_outputs(2644) <= a;
    layer3_outputs(2645) <= not (a or b);
    layer3_outputs(2646) <= b;
    layer3_outputs(2647) <= b and not a;
    layer3_outputs(2648) <= a and b;
    layer3_outputs(2649) <= '0';
    layer3_outputs(2650) <= b and not a;
    layer3_outputs(2651) <= '0';
    layer3_outputs(2652) <= a and not b;
    layer3_outputs(2653) <= b and not a;
    layer3_outputs(2654) <= not a or b;
    layer3_outputs(2655) <= not (a or b);
    layer3_outputs(2656) <= b;
    layer3_outputs(2657) <= not (a or b);
    layer3_outputs(2658) <= not (a and b);
    layer3_outputs(2659) <= '1';
    layer3_outputs(2660) <= not (a or b);
    layer3_outputs(2661) <= a and b;
    layer3_outputs(2662) <= a and not b;
    layer3_outputs(2663) <= b and not a;
    layer3_outputs(2664) <= '1';
    layer3_outputs(2665) <= not a or b;
    layer3_outputs(2666) <= '1';
    layer3_outputs(2667) <= a or b;
    layer3_outputs(2668) <= b;
    layer3_outputs(2669) <= not b;
    layer3_outputs(2670) <= not (a and b);
    layer3_outputs(2671) <= not b or a;
    layer3_outputs(2672) <= not a;
    layer3_outputs(2673) <= a;
    layer3_outputs(2674) <= a and b;
    layer3_outputs(2675) <= not a or b;
    layer3_outputs(2676) <= '1';
    layer3_outputs(2677) <= not a;
    layer3_outputs(2678) <= not b or a;
    layer3_outputs(2679) <= not a or b;
    layer3_outputs(2680) <= not (a and b);
    layer3_outputs(2681) <= a;
    layer3_outputs(2682) <= '1';
    layer3_outputs(2683) <= a and not b;
    layer3_outputs(2684) <= not (a and b);
    layer3_outputs(2685) <= a and not b;
    layer3_outputs(2686) <= not b or a;
    layer3_outputs(2687) <= a or b;
    layer3_outputs(2688) <= b;
    layer3_outputs(2689) <= a xor b;
    layer3_outputs(2690) <= '1';
    layer3_outputs(2691) <= not a;
    layer3_outputs(2692) <= not (a or b);
    layer3_outputs(2693) <= not b;
    layer3_outputs(2694) <= a;
    layer3_outputs(2695) <= not (a or b);
    layer3_outputs(2696) <= not a;
    layer3_outputs(2697) <= not (a or b);
    layer3_outputs(2698) <= b;
    layer3_outputs(2699) <= a;
    layer3_outputs(2700) <= a or b;
    layer3_outputs(2701) <= a xor b;
    layer3_outputs(2702) <= not b or a;
    layer3_outputs(2703) <= not (a or b);
    layer3_outputs(2704) <= not b;
    layer3_outputs(2705) <= a and not b;
    layer3_outputs(2706) <= not (a and b);
    layer3_outputs(2707) <= '1';
    layer3_outputs(2708) <= '1';
    layer3_outputs(2709) <= a and not b;
    layer3_outputs(2710) <= b and not a;
    layer3_outputs(2711) <= a;
    layer3_outputs(2712) <= '0';
    layer3_outputs(2713) <= a or b;
    layer3_outputs(2714) <= a and not b;
    layer3_outputs(2715) <= not a;
    layer3_outputs(2716) <= not (a and b);
    layer3_outputs(2717) <= a and not b;
    layer3_outputs(2718) <= a and not b;
    layer3_outputs(2719) <= not b;
    layer3_outputs(2720) <= not (a and b);
    layer3_outputs(2721) <= b;
    layer3_outputs(2722) <= a and not b;
    layer3_outputs(2723) <= not a or b;
    layer3_outputs(2724) <= a and not b;
    layer3_outputs(2725) <= b and not a;
    layer3_outputs(2726) <= a and not b;
    layer3_outputs(2727) <= a or b;
    layer3_outputs(2728) <= a and not b;
    layer3_outputs(2729) <= not a;
    layer3_outputs(2730) <= '0';
    layer3_outputs(2731) <= b;
    layer3_outputs(2732) <= not b;
    layer3_outputs(2733) <= '0';
    layer3_outputs(2734) <= b and not a;
    layer3_outputs(2735) <= not a or b;
    layer3_outputs(2736) <= '0';
    layer3_outputs(2737) <= not (a or b);
    layer3_outputs(2738) <= a or b;
    layer3_outputs(2739) <= a and b;
    layer3_outputs(2740) <= a and not b;
    layer3_outputs(2741) <= not b or a;
    layer3_outputs(2742) <= a xor b;
    layer3_outputs(2743) <= not (a xor b);
    layer3_outputs(2744) <= not (a or b);
    layer3_outputs(2745) <= a and b;
    layer3_outputs(2746) <= not a or b;
    layer3_outputs(2747) <= a and not b;
    layer3_outputs(2748) <= '1';
    layer3_outputs(2749) <= a and b;
    layer3_outputs(2750) <= not (a or b);
    layer3_outputs(2751) <= not (a or b);
    layer3_outputs(2752) <= not (a and b);
    layer3_outputs(2753) <= a;
    layer3_outputs(2754) <= not b or a;
    layer3_outputs(2755) <= not b or a;
    layer3_outputs(2756) <= '1';
    layer3_outputs(2757) <= b and not a;
    layer3_outputs(2758) <= '1';
    layer3_outputs(2759) <= a;
    layer3_outputs(2760) <= not b;
    layer3_outputs(2761) <= not (a or b);
    layer3_outputs(2762) <= not (a or b);
    layer3_outputs(2763) <= a;
    layer3_outputs(2764) <= a or b;
    layer3_outputs(2765) <= a;
    layer3_outputs(2766) <= b and not a;
    layer3_outputs(2767) <= b and not a;
    layer3_outputs(2768) <= b and not a;
    layer3_outputs(2769) <= a and b;
    layer3_outputs(2770) <= not (a or b);
    layer3_outputs(2771) <= a xor b;
    layer3_outputs(2772) <= not b;
    layer3_outputs(2773) <= b and not a;
    layer3_outputs(2774) <= '0';
    layer3_outputs(2775) <= a and b;
    layer3_outputs(2776) <= a and not b;
    layer3_outputs(2777) <= not (a and b);
    layer3_outputs(2778) <= not b;
    layer3_outputs(2779) <= '1';
    layer3_outputs(2780) <= '0';
    layer3_outputs(2781) <= not b;
    layer3_outputs(2782) <= a and b;
    layer3_outputs(2783) <= '1';
    layer3_outputs(2784) <= a and b;
    layer3_outputs(2785) <= not (a xor b);
    layer3_outputs(2786) <= not a or b;
    layer3_outputs(2787) <= not (a xor b);
    layer3_outputs(2788) <= a;
    layer3_outputs(2789) <= not (a or b);
    layer3_outputs(2790) <= '0';
    layer3_outputs(2791) <= not b or a;
    layer3_outputs(2792) <= a and not b;
    layer3_outputs(2793) <= a and not b;
    layer3_outputs(2794) <= '0';
    layer3_outputs(2795) <= not a;
    layer3_outputs(2796) <= a;
    layer3_outputs(2797) <= '0';
    layer3_outputs(2798) <= b;
    layer3_outputs(2799) <= not (a or b);
    layer3_outputs(2800) <= a;
    layer3_outputs(2801) <= a;
    layer3_outputs(2802) <= a and not b;
    layer3_outputs(2803) <= not (a and b);
    layer3_outputs(2804) <= a and not b;
    layer3_outputs(2805) <= a and b;
    layer3_outputs(2806) <= a or b;
    layer3_outputs(2807) <= not b or a;
    layer3_outputs(2808) <= a and not b;
    layer3_outputs(2809) <= a;
    layer3_outputs(2810) <= not a;
    layer3_outputs(2811) <= a and not b;
    layer3_outputs(2812) <= '1';
    layer3_outputs(2813) <= not (a xor b);
    layer3_outputs(2814) <= a and not b;
    layer3_outputs(2815) <= not b;
    layer3_outputs(2816) <= a and b;
    layer3_outputs(2817) <= '0';
    layer3_outputs(2818) <= not a or b;
    layer3_outputs(2819) <= a;
    layer3_outputs(2820) <= '0';
    layer3_outputs(2821) <= not (a and b);
    layer3_outputs(2822) <= b;
    layer3_outputs(2823) <= a and b;
    layer3_outputs(2824) <= a or b;
    layer3_outputs(2825) <= '1';
    layer3_outputs(2826) <= a xor b;
    layer3_outputs(2827) <= not b or a;
    layer3_outputs(2828) <= a and not b;
    layer3_outputs(2829) <= '0';
    layer3_outputs(2830) <= a or b;
    layer3_outputs(2831) <= not b;
    layer3_outputs(2832) <= a and b;
    layer3_outputs(2833) <= not a or b;
    layer3_outputs(2834) <= not b;
    layer3_outputs(2835) <= not a or b;
    layer3_outputs(2836) <= '0';
    layer3_outputs(2837) <= b and not a;
    layer3_outputs(2838) <= a;
    layer3_outputs(2839) <= not (a xor b);
    layer3_outputs(2840) <= b;
    layer3_outputs(2841) <= b and not a;
    layer3_outputs(2842) <= b;
    layer3_outputs(2843) <= a or b;
    layer3_outputs(2844) <= not b;
    layer3_outputs(2845) <= a and b;
    layer3_outputs(2846) <= b and not a;
    layer3_outputs(2847) <= not (a or b);
    layer3_outputs(2848) <= '0';
    layer3_outputs(2849) <= b and not a;
    layer3_outputs(2850) <= not b;
    layer3_outputs(2851) <= a and not b;
    layer3_outputs(2852) <= not a;
    layer3_outputs(2853) <= not a;
    layer3_outputs(2854) <= '0';
    layer3_outputs(2855) <= '1';
    layer3_outputs(2856) <= a or b;
    layer3_outputs(2857) <= not b or a;
    layer3_outputs(2858) <= '0';
    layer3_outputs(2859) <= '1';
    layer3_outputs(2860) <= a and b;
    layer3_outputs(2861) <= '0';
    layer3_outputs(2862) <= b and not a;
    layer3_outputs(2863) <= a and not b;
    layer3_outputs(2864) <= a;
    layer3_outputs(2865) <= a or b;
    layer3_outputs(2866) <= a and not b;
    layer3_outputs(2867) <= not a or b;
    layer3_outputs(2868) <= not (a or b);
    layer3_outputs(2869) <= not (a or b);
    layer3_outputs(2870) <= '1';
    layer3_outputs(2871) <= '1';
    layer3_outputs(2872) <= not b;
    layer3_outputs(2873) <= not (a and b);
    layer3_outputs(2874) <= a and not b;
    layer3_outputs(2875) <= a or b;
    layer3_outputs(2876) <= b and not a;
    layer3_outputs(2877) <= a and b;
    layer3_outputs(2878) <= not b;
    layer3_outputs(2879) <= '0';
    layer3_outputs(2880) <= not (a or b);
    layer3_outputs(2881) <= a or b;
    layer3_outputs(2882) <= a and b;
    layer3_outputs(2883) <= '0';
    layer3_outputs(2884) <= a or b;
    layer3_outputs(2885) <= not (a or b);
    layer3_outputs(2886) <= not (a and b);
    layer3_outputs(2887) <= '0';
    layer3_outputs(2888) <= '0';
    layer3_outputs(2889) <= a and b;
    layer3_outputs(2890) <= not (a and b);
    layer3_outputs(2891) <= not (a and b);
    layer3_outputs(2892) <= a and b;
    layer3_outputs(2893) <= not (a and b);
    layer3_outputs(2894) <= '1';
    layer3_outputs(2895) <= a or b;
    layer3_outputs(2896) <= '0';
    layer3_outputs(2897) <= b and not a;
    layer3_outputs(2898) <= not b;
    layer3_outputs(2899) <= a;
    layer3_outputs(2900) <= b;
    layer3_outputs(2901) <= not a;
    layer3_outputs(2902) <= a and not b;
    layer3_outputs(2903) <= not (a and b);
    layer3_outputs(2904) <= '1';
    layer3_outputs(2905) <= a xor b;
    layer3_outputs(2906) <= not (a or b);
    layer3_outputs(2907) <= '0';
    layer3_outputs(2908) <= a xor b;
    layer3_outputs(2909) <= '0';
    layer3_outputs(2910) <= not a;
    layer3_outputs(2911) <= '1';
    layer3_outputs(2912) <= a and b;
    layer3_outputs(2913) <= a;
    layer3_outputs(2914) <= '1';
    layer3_outputs(2915) <= '0';
    layer3_outputs(2916) <= not b or a;
    layer3_outputs(2917) <= '0';
    layer3_outputs(2918) <= not a;
    layer3_outputs(2919) <= '0';
    layer3_outputs(2920) <= a and b;
    layer3_outputs(2921) <= a or b;
    layer3_outputs(2922) <= '1';
    layer3_outputs(2923) <= a and not b;
    layer3_outputs(2924) <= not a;
    layer3_outputs(2925) <= a or b;
    layer3_outputs(2926) <= not (a or b);
    layer3_outputs(2927) <= not (a or b);
    layer3_outputs(2928) <= not a;
    layer3_outputs(2929) <= not (a and b);
    layer3_outputs(2930) <= not a or b;
    layer3_outputs(2931) <= a;
    layer3_outputs(2932) <= a and b;
    layer3_outputs(2933) <= not a or b;
    layer3_outputs(2934) <= not (a and b);
    layer3_outputs(2935) <= not b;
    layer3_outputs(2936) <= a and not b;
    layer3_outputs(2937) <= a or b;
    layer3_outputs(2938) <= a and b;
    layer3_outputs(2939) <= not a or b;
    layer3_outputs(2940) <= b;
    layer3_outputs(2941) <= not a or b;
    layer3_outputs(2942) <= '0';
    layer3_outputs(2943) <= a or b;
    layer3_outputs(2944) <= '1';
    layer3_outputs(2945) <= not (a or b);
    layer3_outputs(2946) <= a and b;
    layer3_outputs(2947) <= a or b;
    layer3_outputs(2948) <= not b or a;
    layer3_outputs(2949) <= not b or a;
    layer3_outputs(2950) <= a and b;
    layer3_outputs(2951) <= '0';
    layer3_outputs(2952) <= a or b;
    layer3_outputs(2953) <= not a;
    layer3_outputs(2954) <= not b;
    layer3_outputs(2955) <= not (a and b);
    layer3_outputs(2956) <= not a or b;
    layer3_outputs(2957) <= a and b;
    layer3_outputs(2958) <= not a;
    layer3_outputs(2959) <= a and b;
    layer3_outputs(2960) <= a or b;
    layer3_outputs(2961) <= a or b;
    layer3_outputs(2962) <= not a;
    layer3_outputs(2963) <= not (a and b);
    layer3_outputs(2964) <= not a or b;
    layer3_outputs(2965) <= a xor b;
    layer3_outputs(2966) <= not (a or b);
    layer3_outputs(2967) <= not b or a;
    layer3_outputs(2968) <= a and b;
    layer3_outputs(2969) <= not (a and b);
    layer3_outputs(2970) <= not (a and b);
    layer3_outputs(2971) <= a or b;
    layer3_outputs(2972) <= a;
    layer3_outputs(2973) <= not (a and b);
    layer3_outputs(2974) <= '1';
    layer3_outputs(2975) <= a or b;
    layer3_outputs(2976) <= a and b;
    layer3_outputs(2977) <= not b or a;
    layer3_outputs(2978) <= a;
    layer3_outputs(2979) <= b;
    layer3_outputs(2980) <= b;
    layer3_outputs(2981) <= not (a xor b);
    layer3_outputs(2982) <= not a or b;
    layer3_outputs(2983) <= '0';
    layer3_outputs(2984) <= b and not a;
    layer3_outputs(2985) <= not (a or b);
    layer3_outputs(2986) <= b;
    layer3_outputs(2987) <= not a or b;
    layer3_outputs(2988) <= not (a xor b);
    layer3_outputs(2989) <= not b;
    layer3_outputs(2990) <= not (a xor b);
    layer3_outputs(2991) <= not a;
    layer3_outputs(2992) <= not a;
    layer3_outputs(2993) <= not (a and b);
    layer3_outputs(2994) <= a;
    layer3_outputs(2995) <= not (a and b);
    layer3_outputs(2996) <= not (a and b);
    layer3_outputs(2997) <= '1';
    layer3_outputs(2998) <= a and not b;
    layer3_outputs(2999) <= not a;
    layer3_outputs(3000) <= not a or b;
    layer3_outputs(3001) <= a or b;
    layer3_outputs(3002) <= '0';
    layer3_outputs(3003) <= b and not a;
    layer3_outputs(3004) <= not a;
    layer3_outputs(3005) <= a xor b;
    layer3_outputs(3006) <= a;
    layer3_outputs(3007) <= '0';
    layer3_outputs(3008) <= not (a xor b);
    layer3_outputs(3009) <= not (a or b);
    layer3_outputs(3010) <= not a or b;
    layer3_outputs(3011) <= not (a or b);
    layer3_outputs(3012) <= a xor b;
    layer3_outputs(3013) <= a;
    layer3_outputs(3014) <= not b;
    layer3_outputs(3015) <= not a;
    layer3_outputs(3016) <= a;
    layer3_outputs(3017) <= a;
    layer3_outputs(3018) <= not (a and b);
    layer3_outputs(3019) <= not b;
    layer3_outputs(3020) <= not b or a;
    layer3_outputs(3021) <= not (a or b);
    layer3_outputs(3022) <= not b or a;
    layer3_outputs(3023) <= not a or b;
    layer3_outputs(3024) <= '1';
    layer3_outputs(3025) <= not b or a;
    layer3_outputs(3026) <= a and b;
    layer3_outputs(3027) <= not (a or b);
    layer3_outputs(3028) <= not a or b;
    layer3_outputs(3029) <= not (a or b);
    layer3_outputs(3030) <= not (a or b);
    layer3_outputs(3031) <= not b or a;
    layer3_outputs(3032) <= not b;
    layer3_outputs(3033) <= not a or b;
    layer3_outputs(3034) <= b;
    layer3_outputs(3035) <= not a;
    layer3_outputs(3036) <= not a;
    layer3_outputs(3037) <= a and not b;
    layer3_outputs(3038) <= a and b;
    layer3_outputs(3039) <= b;
    layer3_outputs(3040) <= '1';
    layer3_outputs(3041) <= a and not b;
    layer3_outputs(3042) <= not (a or b);
    layer3_outputs(3043) <= a and b;
    layer3_outputs(3044) <= '0';
    layer3_outputs(3045) <= b;
    layer3_outputs(3046) <= not (a and b);
    layer3_outputs(3047) <= b and not a;
    layer3_outputs(3048) <= a and b;
    layer3_outputs(3049) <= a and not b;
    layer3_outputs(3050) <= b;
    layer3_outputs(3051) <= b and not a;
    layer3_outputs(3052) <= not a;
    layer3_outputs(3053) <= not b or a;
    layer3_outputs(3054) <= b;
    layer3_outputs(3055) <= not b or a;
    layer3_outputs(3056) <= not (a and b);
    layer3_outputs(3057) <= a or b;
    layer3_outputs(3058) <= not a;
    layer3_outputs(3059) <= not (a and b);
    layer3_outputs(3060) <= not (a or b);
    layer3_outputs(3061) <= '0';
    layer3_outputs(3062) <= '0';
    layer3_outputs(3063) <= '1';
    layer3_outputs(3064) <= '0';
    layer3_outputs(3065) <= not a;
    layer3_outputs(3066) <= a or b;
    layer3_outputs(3067) <= not a;
    layer3_outputs(3068) <= a and not b;
    layer3_outputs(3069) <= a or b;
    layer3_outputs(3070) <= a;
    layer3_outputs(3071) <= not (a and b);
    layer3_outputs(3072) <= a;
    layer3_outputs(3073) <= b;
    layer3_outputs(3074) <= '1';
    layer3_outputs(3075) <= a;
    layer3_outputs(3076) <= a or b;
    layer3_outputs(3077) <= not (a or b);
    layer3_outputs(3078) <= b;
    layer3_outputs(3079) <= not b or a;
    layer3_outputs(3080) <= b and not a;
    layer3_outputs(3081) <= '0';
    layer3_outputs(3082) <= not a;
    layer3_outputs(3083) <= a and not b;
    layer3_outputs(3084) <= '0';
    layer3_outputs(3085) <= not (a xor b);
    layer3_outputs(3086) <= not a or b;
    layer3_outputs(3087) <= not (a or b);
    layer3_outputs(3088) <= not b;
    layer3_outputs(3089) <= a and not b;
    layer3_outputs(3090) <= a or b;
    layer3_outputs(3091) <= b and not a;
    layer3_outputs(3092) <= b and not a;
    layer3_outputs(3093) <= a or b;
    layer3_outputs(3094) <= a xor b;
    layer3_outputs(3095) <= not (a and b);
    layer3_outputs(3096) <= a and not b;
    layer3_outputs(3097) <= '0';
    layer3_outputs(3098) <= a;
    layer3_outputs(3099) <= a;
    layer3_outputs(3100) <= '1';
    layer3_outputs(3101) <= not a or b;
    layer3_outputs(3102) <= not a;
    layer3_outputs(3103) <= a or b;
    layer3_outputs(3104) <= not a;
    layer3_outputs(3105) <= not a;
    layer3_outputs(3106) <= not (a and b);
    layer3_outputs(3107) <= not a or b;
    layer3_outputs(3108) <= a and b;
    layer3_outputs(3109) <= '1';
    layer3_outputs(3110) <= b;
    layer3_outputs(3111) <= not (a and b);
    layer3_outputs(3112) <= a xor b;
    layer3_outputs(3113) <= a or b;
    layer3_outputs(3114) <= '1';
    layer3_outputs(3115) <= b;
    layer3_outputs(3116) <= not a;
    layer3_outputs(3117) <= not a;
    layer3_outputs(3118) <= a or b;
    layer3_outputs(3119) <= not a;
    layer3_outputs(3120) <= '1';
    layer3_outputs(3121) <= a or b;
    layer3_outputs(3122) <= a and b;
    layer3_outputs(3123) <= b;
    layer3_outputs(3124) <= a;
    layer3_outputs(3125) <= a or b;
    layer3_outputs(3126) <= not (a and b);
    layer3_outputs(3127) <= not a or b;
    layer3_outputs(3128) <= not a;
    layer3_outputs(3129) <= a;
    layer3_outputs(3130) <= a;
    layer3_outputs(3131) <= not b or a;
    layer3_outputs(3132) <= not b;
    layer3_outputs(3133) <= b and not a;
    layer3_outputs(3134) <= b and not a;
    layer3_outputs(3135) <= a and b;
    layer3_outputs(3136) <= a and b;
    layer3_outputs(3137) <= not (a and b);
    layer3_outputs(3138) <= '0';
    layer3_outputs(3139) <= not a or b;
    layer3_outputs(3140) <= not b or a;
    layer3_outputs(3141) <= '1';
    layer3_outputs(3142) <= not b;
    layer3_outputs(3143) <= '0';
    layer3_outputs(3144) <= not a;
    layer3_outputs(3145) <= a and not b;
    layer3_outputs(3146) <= not (a and b);
    layer3_outputs(3147) <= '1';
    layer3_outputs(3148) <= not a or b;
    layer3_outputs(3149) <= a or b;
    layer3_outputs(3150) <= '1';
    layer3_outputs(3151) <= b;
    layer3_outputs(3152) <= not (a and b);
    layer3_outputs(3153) <= '0';
    layer3_outputs(3154) <= a and not b;
    layer3_outputs(3155) <= a;
    layer3_outputs(3156) <= not b or a;
    layer3_outputs(3157) <= b;
    layer3_outputs(3158) <= a and b;
    layer3_outputs(3159) <= a xor b;
    layer3_outputs(3160) <= '1';
    layer3_outputs(3161) <= a and not b;
    layer3_outputs(3162) <= a;
    layer3_outputs(3163) <= a xor b;
    layer3_outputs(3164) <= b;
    layer3_outputs(3165) <= not (a or b);
    layer3_outputs(3166) <= b and not a;
    layer3_outputs(3167) <= not b or a;
    layer3_outputs(3168) <= not (a and b);
    layer3_outputs(3169) <= not a;
    layer3_outputs(3170) <= not (a and b);
    layer3_outputs(3171) <= a and b;
    layer3_outputs(3172) <= '1';
    layer3_outputs(3173) <= a and not b;
    layer3_outputs(3174) <= not b;
    layer3_outputs(3175) <= a xor b;
    layer3_outputs(3176) <= a;
    layer3_outputs(3177) <= not b;
    layer3_outputs(3178) <= a;
    layer3_outputs(3179) <= not (a and b);
    layer3_outputs(3180) <= a;
    layer3_outputs(3181) <= b and not a;
    layer3_outputs(3182) <= b;
    layer3_outputs(3183) <= a or b;
    layer3_outputs(3184) <= not (a or b);
    layer3_outputs(3185) <= a and not b;
    layer3_outputs(3186) <= not b or a;
    layer3_outputs(3187) <= not b;
    layer3_outputs(3188) <= not b;
    layer3_outputs(3189) <= not b;
    layer3_outputs(3190) <= not (a or b);
    layer3_outputs(3191) <= not b;
    layer3_outputs(3192) <= not a or b;
    layer3_outputs(3193) <= a;
    layer3_outputs(3194) <= '1';
    layer3_outputs(3195) <= a and b;
    layer3_outputs(3196) <= a;
    layer3_outputs(3197) <= a;
    layer3_outputs(3198) <= not b;
    layer3_outputs(3199) <= not (a and b);
    layer3_outputs(3200) <= a and b;
    layer3_outputs(3201) <= '1';
    layer3_outputs(3202) <= not b or a;
    layer3_outputs(3203) <= b;
    layer3_outputs(3204) <= a and not b;
    layer3_outputs(3205) <= b;
    layer3_outputs(3206) <= not (a or b);
    layer3_outputs(3207) <= '1';
    layer3_outputs(3208) <= b and not a;
    layer3_outputs(3209) <= a;
    layer3_outputs(3210) <= not b or a;
    layer3_outputs(3211) <= '0';
    layer3_outputs(3212) <= a and not b;
    layer3_outputs(3213) <= not b or a;
    layer3_outputs(3214) <= not a;
    layer3_outputs(3215) <= a and not b;
    layer3_outputs(3216) <= not (a or b);
    layer3_outputs(3217) <= not b;
    layer3_outputs(3218) <= not a;
    layer3_outputs(3219) <= not (a or b);
    layer3_outputs(3220) <= '0';
    layer3_outputs(3221) <= b;
    layer3_outputs(3222) <= not a;
    layer3_outputs(3223) <= a or b;
    layer3_outputs(3224) <= b;
    layer3_outputs(3225) <= not (a and b);
    layer3_outputs(3226) <= b and not a;
    layer3_outputs(3227) <= a and not b;
    layer3_outputs(3228) <= not (a or b);
    layer3_outputs(3229) <= b and not a;
    layer3_outputs(3230) <= '0';
    layer3_outputs(3231) <= not a;
    layer3_outputs(3232) <= not (a or b);
    layer3_outputs(3233) <= '1';
    layer3_outputs(3234) <= b and not a;
    layer3_outputs(3235) <= not b;
    layer3_outputs(3236) <= not (a or b);
    layer3_outputs(3237) <= not b;
    layer3_outputs(3238) <= b and not a;
    layer3_outputs(3239) <= not b;
    layer3_outputs(3240) <= a or b;
    layer3_outputs(3241) <= a;
    layer3_outputs(3242) <= not (a or b);
    layer3_outputs(3243) <= b and not a;
    layer3_outputs(3244) <= not b or a;
    layer3_outputs(3245) <= not b or a;
    layer3_outputs(3246) <= not b or a;
    layer3_outputs(3247) <= b and not a;
    layer3_outputs(3248) <= a and not b;
    layer3_outputs(3249) <= a and b;
    layer3_outputs(3250) <= a;
    layer3_outputs(3251) <= not (a or b);
    layer3_outputs(3252) <= a and not b;
    layer3_outputs(3253) <= not a;
    layer3_outputs(3254) <= not (a and b);
    layer3_outputs(3255) <= a xor b;
    layer3_outputs(3256) <= not (a or b);
    layer3_outputs(3257) <= not (a or b);
    layer3_outputs(3258) <= not a or b;
    layer3_outputs(3259) <= b;
    layer3_outputs(3260) <= '1';
    layer3_outputs(3261) <= '0';
    layer3_outputs(3262) <= b and not a;
    layer3_outputs(3263) <= a or b;
    layer3_outputs(3264) <= '1';
    layer3_outputs(3265) <= not a;
    layer3_outputs(3266) <= '1';
    layer3_outputs(3267) <= not (a and b);
    layer3_outputs(3268) <= '1';
    layer3_outputs(3269) <= not a or b;
    layer3_outputs(3270) <= '1';
    layer3_outputs(3271) <= a and b;
    layer3_outputs(3272) <= not a;
    layer3_outputs(3273) <= a and not b;
    layer3_outputs(3274) <= '0';
    layer3_outputs(3275) <= '1';
    layer3_outputs(3276) <= not b;
    layer3_outputs(3277) <= '1';
    layer3_outputs(3278) <= a or b;
    layer3_outputs(3279) <= not b;
    layer3_outputs(3280) <= '0';
    layer3_outputs(3281) <= a and not b;
    layer3_outputs(3282) <= not b or a;
    layer3_outputs(3283) <= b;
    layer3_outputs(3284) <= not a;
    layer3_outputs(3285) <= not b or a;
    layer3_outputs(3286) <= not b;
    layer3_outputs(3287) <= not b;
    layer3_outputs(3288) <= a and b;
    layer3_outputs(3289) <= a and not b;
    layer3_outputs(3290) <= not b;
    layer3_outputs(3291) <= a and not b;
    layer3_outputs(3292) <= '0';
    layer3_outputs(3293) <= not b;
    layer3_outputs(3294) <= '1';
    layer3_outputs(3295) <= '0';
    layer3_outputs(3296) <= not b or a;
    layer3_outputs(3297) <= a;
    layer3_outputs(3298) <= not a or b;
    layer3_outputs(3299) <= a or b;
    layer3_outputs(3300) <= not b or a;
    layer3_outputs(3301) <= a;
    layer3_outputs(3302) <= a or b;
    layer3_outputs(3303) <= not b;
    layer3_outputs(3304) <= a;
    layer3_outputs(3305) <= not a;
    layer3_outputs(3306) <= '0';
    layer3_outputs(3307) <= a;
    layer3_outputs(3308) <= a and not b;
    layer3_outputs(3309) <= a;
    layer3_outputs(3310) <= not a or b;
    layer3_outputs(3311) <= not (a or b);
    layer3_outputs(3312) <= b;
    layer3_outputs(3313) <= not (a or b);
    layer3_outputs(3314) <= '0';
    layer3_outputs(3315) <= a and b;
    layer3_outputs(3316) <= not (a or b);
    layer3_outputs(3317) <= not (a and b);
    layer3_outputs(3318) <= a and b;
    layer3_outputs(3319) <= '0';
    layer3_outputs(3320) <= a and b;
    layer3_outputs(3321) <= not a or b;
    layer3_outputs(3322) <= not a;
    layer3_outputs(3323) <= not b;
    layer3_outputs(3324) <= not b;
    layer3_outputs(3325) <= a and not b;
    layer3_outputs(3326) <= not a;
    layer3_outputs(3327) <= not b;
    layer3_outputs(3328) <= not a;
    layer3_outputs(3329) <= b;
    layer3_outputs(3330) <= a or b;
    layer3_outputs(3331) <= a and b;
    layer3_outputs(3332) <= a and b;
    layer3_outputs(3333) <= '0';
    layer3_outputs(3334) <= '0';
    layer3_outputs(3335) <= not (a and b);
    layer3_outputs(3336) <= a;
    layer3_outputs(3337) <= '1';
    layer3_outputs(3338) <= a and b;
    layer3_outputs(3339) <= b and not a;
    layer3_outputs(3340) <= not a or b;
    layer3_outputs(3341) <= '0';
    layer3_outputs(3342) <= '1';
    layer3_outputs(3343) <= not (a or b);
    layer3_outputs(3344) <= not a or b;
    layer3_outputs(3345) <= a xor b;
    layer3_outputs(3346) <= not a;
    layer3_outputs(3347) <= not b or a;
    layer3_outputs(3348) <= '0';
    layer3_outputs(3349) <= not b or a;
    layer3_outputs(3350) <= b and not a;
    layer3_outputs(3351) <= '0';
    layer3_outputs(3352) <= not b;
    layer3_outputs(3353) <= not b;
    layer3_outputs(3354) <= not a;
    layer3_outputs(3355) <= not a or b;
    layer3_outputs(3356) <= not a or b;
    layer3_outputs(3357) <= a or b;
    layer3_outputs(3358) <= not b;
    layer3_outputs(3359) <= a xor b;
    layer3_outputs(3360) <= a and b;
    layer3_outputs(3361) <= not a or b;
    layer3_outputs(3362) <= not a;
    layer3_outputs(3363) <= b and not a;
    layer3_outputs(3364) <= not (a and b);
    layer3_outputs(3365) <= a and not b;
    layer3_outputs(3366) <= '0';
    layer3_outputs(3367) <= not b or a;
    layer3_outputs(3368) <= not b;
    layer3_outputs(3369) <= not b or a;
    layer3_outputs(3370) <= not a;
    layer3_outputs(3371) <= b and not a;
    layer3_outputs(3372) <= a and b;
    layer3_outputs(3373) <= a;
    layer3_outputs(3374) <= '0';
    layer3_outputs(3375) <= a and b;
    layer3_outputs(3376) <= not a;
    layer3_outputs(3377) <= not a;
    layer3_outputs(3378) <= a;
    layer3_outputs(3379) <= not (a or b);
    layer3_outputs(3380) <= not a;
    layer3_outputs(3381) <= b;
    layer3_outputs(3382) <= b and not a;
    layer3_outputs(3383) <= a;
    layer3_outputs(3384) <= b;
    layer3_outputs(3385) <= not a or b;
    layer3_outputs(3386) <= b and not a;
    layer3_outputs(3387) <= a or b;
    layer3_outputs(3388) <= a and not b;
    layer3_outputs(3389) <= not b;
    layer3_outputs(3390) <= a and b;
    layer3_outputs(3391) <= not (a xor b);
    layer3_outputs(3392) <= '1';
    layer3_outputs(3393) <= not b or a;
    layer3_outputs(3394) <= not (a and b);
    layer3_outputs(3395) <= a and b;
    layer3_outputs(3396) <= '1';
    layer3_outputs(3397) <= not a or b;
    layer3_outputs(3398) <= b;
    layer3_outputs(3399) <= not (a or b);
    layer3_outputs(3400) <= not b;
    layer3_outputs(3401) <= '0';
    layer3_outputs(3402) <= b and not a;
    layer3_outputs(3403) <= not a or b;
    layer3_outputs(3404) <= not (a and b);
    layer3_outputs(3405) <= not (a and b);
    layer3_outputs(3406) <= not b;
    layer3_outputs(3407) <= a and b;
    layer3_outputs(3408) <= '0';
    layer3_outputs(3409) <= not a or b;
    layer3_outputs(3410) <= a and b;
    layer3_outputs(3411) <= not b or a;
    layer3_outputs(3412) <= '1';
    layer3_outputs(3413) <= not (a and b);
    layer3_outputs(3414) <= not a or b;
    layer3_outputs(3415) <= not a;
    layer3_outputs(3416) <= a;
    layer3_outputs(3417) <= '1';
    layer3_outputs(3418) <= a and not b;
    layer3_outputs(3419) <= '0';
    layer3_outputs(3420) <= '1';
    layer3_outputs(3421) <= not b or a;
    layer3_outputs(3422) <= a or b;
    layer3_outputs(3423) <= not a or b;
    layer3_outputs(3424) <= '0';
    layer3_outputs(3425) <= b and not a;
    layer3_outputs(3426) <= a;
    layer3_outputs(3427) <= a and b;
    layer3_outputs(3428) <= a and not b;
    layer3_outputs(3429) <= a and b;
    layer3_outputs(3430) <= a and b;
    layer3_outputs(3431) <= a or b;
    layer3_outputs(3432) <= not b;
    layer3_outputs(3433) <= not b or a;
    layer3_outputs(3434) <= a or b;
    layer3_outputs(3435) <= a;
    layer3_outputs(3436) <= not a or b;
    layer3_outputs(3437) <= not a or b;
    layer3_outputs(3438) <= '0';
    layer3_outputs(3439) <= not a or b;
    layer3_outputs(3440) <= a;
    layer3_outputs(3441) <= not (a and b);
    layer3_outputs(3442) <= a and not b;
    layer3_outputs(3443) <= '1';
    layer3_outputs(3444) <= a and not b;
    layer3_outputs(3445) <= '1';
    layer3_outputs(3446) <= not a or b;
    layer3_outputs(3447) <= '1';
    layer3_outputs(3448) <= '0';
    layer3_outputs(3449) <= not b or a;
    layer3_outputs(3450) <= not b or a;
    layer3_outputs(3451) <= not a;
    layer3_outputs(3452) <= b;
    layer3_outputs(3453) <= not (a or b);
    layer3_outputs(3454) <= b and not a;
    layer3_outputs(3455) <= not (a or b);
    layer3_outputs(3456) <= a and b;
    layer3_outputs(3457) <= b;
    layer3_outputs(3458) <= b;
    layer3_outputs(3459) <= not (a or b);
    layer3_outputs(3460) <= b and not a;
    layer3_outputs(3461) <= a;
    layer3_outputs(3462) <= not a or b;
    layer3_outputs(3463) <= '1';
    layer3_outputs(3464) <= b;
    layer3_outputs(3465) <= '0';
    layer3_outputs(3466) <= '0';
    layer3_outputs(3467) <= b;
    layer3_outputs(3468) <= not (a or b);
    layer3_outputs(3469) <= not b;
    layer3_outputs(3470) <= '0';
    layer3_outputs(3471) <= not b;
    layer3_outputs(3472) <= a and b;
    layer3_outputs(3473) <= a;
    layer3_outputs(3474) <= a and b;
    layer3_outputs(3475) <= '1';
    layer3_outputs(3476) <= not b;
    layer3_outputs(3477) <= '1';
    layer3_outputs(3478) <= not a;
    layer3_outputs(3479) <= not (a or b);
    layer3_outputs(3480) <= a or b;
    layer3_outputs(3481) <= a or b;
    layer3_outputs(3482) <= b and not a;
    layer3_outputs(3483) <= a and not b;
    layer3_outputs(3484) <= not b or a;
    layer3_outputs(3485) <= b;
    layer3_outputs(3486) <= b;
    layer3_outputs(3487) <= b and not a;
    layer3_outputs(3488) <= a xor b;
    layer3_outputs(3489) <= not b or a;
    layer3_outputs(3490) <= not (a xor b);
    layer3_outputs(3491) <= not b or a;
    layer3_outputs(3492) <= b and not a;
    layer3_outputs(3493) <= a;
    layer3_outputs(3494) <= a or b;
    layer3_outputs(3495) <= not a or b;
    layer3_outputs(3496) <= not (a or b);
    layer3_outputs(3497) <= not b;
    layer3_outputs(3498) <= b;
    layer3_outputs(3499) <= a or b;
    layer3_outputs(3500) <= '1';
    layer3_outputs(3501) <= not a or b;
    layer3_outputs(3502) <= not (a and b);
    layer3_outputs(3503) <= b and not a;
    layer3_outputs(3504) <= b and not a;
    layer3_outputs(3505) <= a and not b;
    layer3_outputs(3506) <= a and b;
    layer3_outputs(3507) <= a and not b;
    layer3_outputs(3508) <= a and not b;
    layer3_outputs(3509) <= '1';
    layer3_outputs(3510) <= not b or a;
    layer3_outputs(3511) <= not (a or b);
    layer3_outputs(3512) <= a;
    layer3_outputs(3513) <= not b;
    layer3_outputs(3514) <= a;
    layer3_outputs(3515) <= not a or b;
    layer3_outputs(3516) <= '1';
    layer3_outputs(3517) <= a and b;
    layer3_outputs(3518) <= a and b;
    layer3_outputs(3519) <= a and b;
    layer3_outputs(3520) <= not a or b;
    layer3_outputs(3521) <= not (a and b);
    layer3_outputs(3522) <= a;
    layer3_outputs(3523) <= '1';
    layer3_outputs(3524) <= a xor b;
    layer3_outputs(3525) <= '1';
    layer3_outputs(3526) <= not b or a;
    layer3_outputs(3527) <= not (a or b);
    layer3_outputs(3528) <= b;
    layer3_outputs(3529) <= '0';
    layer3_outputs(3530) <= not a;
    layer3_outputs(3531) <= not (a and b);
    layer3_outputs(3532) <= a;
    layer3_outputs(3533) <= b;
    layer3_outputs(3534) <= not (a or b);
    layer3_outputs(3535) <= b;
    layer3_outputs(3536) <= a or b;
    layer3_outputs(3537) <= '1';
    layer3_outputs(3538) <= a;
    layer3_outputs(3539) <= a;
    layer3_outputs(3540) <= not b;
    layer3_outputs(3541) <= a or b;
    layer3_outputs(3542) <= not (a or b);
    layer3_outputs(3543) <= '1';
    layer3_outputs(3544) <= b;
    layer3_outputs(3545) <= '0';
    layer3_outputs(3546) <= '0';
    layer3_outputs(3547) <= not (a xor b);
    layer3_outputs(3548) <= not b or a;
    layer3_outputs(3549) <= b;
    layer3_outputs(3550) <= b and not a;
    layer3_outputs(3551) <= not b;
    layer3_outputs(3552) <= a or b;
    layer3_outputs(3553) <= '1';
    layer3_outputs(3554) <= a;
    layer3_outputs(3555) <= a or b;
    layer3_outputs(3556) <= not a or b;
    layer3_outputs(3557) <= b and not a;
    layer3_outputs(3558) <= '1';
    layer3_outputs(3559) <= not (a or b);
    layer3_outputs(3560) <= a;
    layer3_outputs(3561) <= not a or b;
    layer3_outputs(3562) <= not b;
    layer3_outputs(3563) <= not b;
    layer3_outputs(3564) <= a or b;
    layer3_outputs(3565) <= b and not a;
    layer3_outputs(3566) <= a and b;
    layer3_outputs(3567) <= not (a xor b);
    layer3_outputs(3568) <= a and b;
    layer3_outputs(3569) <= not a;
    layer3_outputs(3570) <= not a or b;
    layer3_outputs(3571) <= '0';
    layer3_outputs(3572) <= a and not b;
    layer3_outputs(3573) <= not (a or b);
    layer3_outputs(3574) <= b;
    layer3_outputs(3575) <= not (a or b);
    layer3_outputs(3576) <= a and b;
    layer3_outputs(3577) <= '1';
    layer3_outputs(3578) <= a or b;
    layer3_outputs(3579) <= not (a or b);
    layer3_outputs(3580) <= b;
    layer3_outputs(3581) <= a and b;
    layer3_outputs(3582) <= not (a and b);
    layer3_outputs(3583) <= '0';
    layer3_outputs(3584) <= not a;
    layer3_outputs(3585) <= b and not a;
    layer3_outputs(3586) <= a;
    layer3_outputs(3587) <= '0';
    layer3_outputs(3588) <= a or b;
    layer3_outputs(3589) <= b;
    layer3_outputs(3590) <= b and not a;
    layer3_outputs(3591) <= a and b;
    layer3_outputs(3592) <= '1';
    layer3_outputs(3593) <= a or b;
    layer3_outputs(3594) <= not (a and b);
    layer3_outputs(3595) <= a and not b;
    layer3_outputs(3596) <= not a or b;
    layer3_outputs(3597) <= not a;
    layer3_outputs(3598) <= not (a or b);
    layer3_outputs(3599) <= '0';
    layer3_outputs(3600) <= b;
    layer3_outputs(3601) <= not a or b;
    layer3_outputs(3602) <= not a;
    layer3_outputs(3603) <= not a;
    layer3_outputs(3604) <= not (a or b);
    layer3_outputs(3605) <= a;
    layer3_outputs(3606) <= '1';
    layer3_outputs(3607) <= a;
    layer3_outputs(3608) <= not (a and b);
    layer3_outputs(3609) <= a;
    layer3_outputs(3610) <= not a;
    layer3_outputs(3611) <= b;
    layer3_outputs(3612) <= not (a or b);
    layer3_outputs(3613) <= not b or a;
    layer3_outputs(3614) <= a and not b;
    layer3_outputs(3615) <= not a;
    layer3_outputs(3616) <= not a or b;
    layer3_outputs(3617) <= a;
    layer3_outputs(3618) <= b and not a;
    layer3_outputs(3619) <= not b;
    layer3_outputs(3620) <= a xor b;
    layer3_outputs(3621) <= '0';
    layer3_outputs(3622) <= b;
    layer3_outputs(3623) <= not a;
    layer3_outputs(3624) <= '0';
    layer3_outputs(3625) <= b and not a;
    layer3_outputs(3626) <= not (a and b);
    layer3_outputs(3627) <= a and b;
    layer3_outputs(3628) <= not a;
    layer3_outputs(3629) <= not a;
    layer3_outputs(3630) <= '1';
    layer3_outputs(3631) <= a and not b;
    layer3_outputs(3632) <= '0';
    layer3_outputs(3633) <= '0';
    layer3_outputs(3634) <= a or b;
    layer3_outputs(3635) <= not b;
    layer3_outputs(3636) <= not b;
    layer3_outputs(3637) <= not (a or b);
    layer3_outputs(3638) <= not (a or b);
    layer3_outputs(3639) <= b and not a;
    layer3_outputs(3640) <= b and not a;
    layer3_outputs(3641) <= not b or a;
    layer3_outputs(3642) <= a and b;
    layer3_outputs(3643) <= a and not b;
    layer3_outputs(3644) <= not (a or b);
    layer3_outputs(3645) <= '0';
    layer3_outputs(3646) <= '1';
    layer3_outputs(3647) <= a and not b;
    layer3_outputs(3648) <= '0';
    layer3_outputs(3649) <= not (a and b);
    layer3_outputs(3650) <= b and not a;
    layer3_outputs(3651) <= not b;
    layer3_outputs(3652) <= not b or a;
    layer3_outputs(3653) <= not (a or b);
    layer3_outputs(3654) <= '1';
    layer3_outputs(3655) <= b and not a;
    layer3_outputs(3656) <= a;
    layer3_outputs(3657) <= not b;
    layer3_outputs(3658) <= a and not b;
    layer3_outputs(3659) <= not (a and b);
    layer3_outputs(3660) <= not b;
    layer3_outputs(3661) <= not b or a;
    layer3_outputs(3662) <= not (a or b);
    layer3_outputs(3663) <= '0';
    layer3_outputs(3664) <= not (a or b);
    layer3_outputs(3665) <= a;
    layer3_outputs(3666) <= b;
    layer3_outputs(3667) <= '0';
    layer3_outputs(3668) <= not a;
    layer3_outputs(3669) <= a and b;
    layer3_outputs(3670) <= not b or a;
    layer3_outputs(3671) <= not a or b;
    layer3_outputs(3672) <= not a;
    layer3_outputs(3673) <= '1';
    layer3_outputs(3674) <= not b or a;
    layer3_outputs(3675) <= b and not a;
    layer3_outputs(3676) <= not a;
    layer3_outputs(3677) <= not a or b;
    layer3_outputs(3678) <= not b or a;
    layer3_outputs(3679) <= not b or a;
    layer3_outputs(3680) <= a and not b;
    layer3_outputs(3681) <= not b or a;
    layer3_outputs(3682) <= not a or b;
    layer3_outputs(3683) <= a and b;
    layer3_outputs(3684) <= a and b;
    layer3_outputs(3685) <= a;
    layer3_outputs(3686) <= b;
    layer3_outputs(3687) <= a and not b;
    layer3_outputs(3688) <= '0';
    layer3_outputs(3689) <= not a;
    layer3_outputs(3690) <= not (a xor b);
    layer3_outputs(3691) <= not b;
    layer3_outputs(3692) <= not a;
    layer3_outputs(3693) <= not b;
    layer3_outputs(3694) <= not (a xor b);
    layer3_outputs(3695) <= b;
    layer3_outputs(3696) <= not (a and b);
    layer3_outputs(3697) <= a and b;
    layer3_outputs(3698) <= not b or a;
    layer3_outputs(3699) <= a and not b;
    layer3_outputs(3700) <= '0';
    layer3_outputs(3701) <= not b;
    layer3_outputs(3702) <= a and not b;
    layer3_outputs(3703) <= not b;
    layer3_outputs(3704) <= a and not b;
    layer3_outputs(3705) <= not (a xor b);
    layer3_outputs(3706) <= '0';
    layer3_outputs(3707) <= not a or b;
    layer3_outputs(3708) <= '0';
    layer3_outputs(3709) <= b and not a;
    layer3_outputs(3710) <= a;
    layer3_outputs(3711) <= not a or b;
    layer3_outputs(3712) <= a;
    layer3_outputs(3713) <= a or b;
    layer3_outputs(3714) <= '0';
    layer3_outputs(3715) <= b and not a;
    layer3_outputs(3716) <= not a;
    layer3_outputs(3717) <= a and not b;
    layer3_outputs(3718) <= b and not a;
    layer3_outputs(3719) <= not a or b;
    layer3_outputs(3720) <= a or b;
    layer3_outputs(3721) <= not a or b;
    layer3_outputs(3722) <= b;
    layer3_outputs(3723) <= '0';
    layer3_outputs(3724) <= b and not a;
    layer3_outputs(3725) <= a and b;
    layer3_outputs(3726) <= '1';
    layer3_outputs(3727) <= '0';
    layer3_outputs(3728) <= a and not b;
    layer3_outputs(3729) <= '0';
    layer3_outputs(3730) <= '1';
    layer3_outputs(3731) <= not (a or b);
    layer3_outputs(3732) <= not a;
    layer3_outputs(3733) <= a or b;
    layer3_outputs(3734) <= not a;
    layer3_outputs(3735) <= not a;
    layer3_outputs(3736) <= not a or b;
    layer3_outputs(3737) <= not b;
    layer3_outputs(3738) <= a and not b;
    layer3_outputs(3739) <= a and b;
    layer3_outputs(3740) <= a or b;
    layer3_outputs(3741) <= '0';
    layer3_outputs(3742) <= b;
    layer3_outputs(3743) <= '0';
    layer3_outputs(3744) <= not (a xor b);
    layer3_outputs(3745) <= a and not b;
    layer3_outputs(3746) <= a;
    layer3_outputs(3747) <= '0';
    layer3_outputs(3748) <= '1';
    layer3_outputs(3749) <= '0';
    layer3_outputs(3750) <= a or b;
    layer3_outputs(3751) <= b;
    layer3_outputs(3752) <= a and not b;
    layer3_outputs(3753) <= '0';
    layer3_outputs(3754) <= not b or a;
    layer3_outputs(3755) <= a;
    layer3_outputs(3756) <= not (a and b);
    layer3_outputs(3757) <= a xor b;
    layer3_outputs(3758) <= b;
    layer3_outputs(3759) <= not a;
    layer3_outputs(3760) <= b;
    layer3_outputs(3761) <= a and b;
    layer3_outputs(3762) <= '0';
    layer3_outputs(3763) <= not b or a;
    layer3_outputs(3764) <= a or b;
    layer3_outputs(3765) <= a and not b;
    layer3_outputs(3766) <= a and b;
    layer3_outputs(3767) <= not a;
    layer3_outputs(3768) <= not a or b;
    layer3_outputs(3769) <= a or b;
    layer3_outputs(3770) <= not (a or b);
    layer3_outputs(3771) <= '0';
    layer3_outputs(3772) <= a;
    layer3_outputs(3773) <= a or b;
    layer3_outputs(3774) <= not (a and b);
    layer3_outputs(3775) <= not a or b;
    layer3_outputs(3776) <= '0';
    layer3_outputs(3777) <= a xor b;
    layer3_outputs(3778) <= b;
    layer3_outputs(3779) <= a or b;
    layer3_outputs(3780) <= not (a and b);
    layer3_outputs(3781) <= not a;
    layer3_outputs(3782) <= not (a or b);
    layer3_outputs(3783) <= '1';
    layer3_outputs(3784) <= b and not a;
    layer3_outputs(3785) <= not (a or b);
    layer3_outputs(3786) <= a;
    layer3_outputs(3787) <= b and not a;
    layer3_outputs(3788) <= b;
    layer3_outputs(3789) <= b;
    layer3_outputs(3790) <= a and b;
    layer3_outputs(3791) <= not (a and b);
    layer3_outputs(3792) <= a or b;
    layer3_outputs(3793) <= b;
    layer3_outputs(3794) <= not a or b;
    layer3_outputs(3795) <= a and not b;
    layer3_outputs(3796) <= a or b;
    layer3_outputs(3797) <= not (a and b);
    layer3_outputs(3798) <= not a or b;
    layer3_outputs(3799) <= a and b;
    layer3_outputs(3800) <= '1';
    layer3_outputs(3801) <= '1';
    layer3_outputs(3802) <= a and not b;
    layer3_outputs(3803) <= a and b;
    layer3_outputs(3804) <= not (a and b);
    layer3_outputs(3805) <= a and b;
    layer3_outputs(3806) <= not (a or b);
    layer3_outputs(3807) <= '0';
    layer3_outputs(3808) <= a and not b;
    layer3_outputs(3809) <= a xor b;
    layer3_outputs(3810) <= not (a and b);
    layer3_outputs(3811) <= not b;
    layer3_outputs(3812) <= a xor b;
    layer3_outputs(3813) <= b and not a;
    layer3_outputs(3814) <= not (a and b);
    layer3_outputs(3815) <= '1';
    layer3_outputs(3816) <= not (a and b);
    layer3_outputs(3817) <= not a;
    layer3_outputs(3818) <= b;
    layer3_outputs(3819) <= not (a and b);
    layer3_outputs(3820) <= not b;
    layer3_outputs(3821) <= a;
    layer3_outputs(3822) <= not b;
    layer3_outputs(3823) <= not b;
    layer3_outputs(3824) <= a and not b;
    layer3_outputs(3825) <= not a or b;
    layer3_outputs(3826) <= not a;
    layer3_outputs(3827) <= not (a or b);
    layer3_outputs(3828) <= b;
    layer3_outputs(3829) <= '0';
    layer3_outputs(3830) <= not a;
    layer3_outputs(3831) <= not a or b;
    layer3_outputs(3832) <= not a or b;
    layer3_outputs(3833) <= a and b;
    layer3_outputs(3834) <= '1';
    layer3_outputs(3835) <= a and not b;
    layer3_outputs(3836) <= b;
    layer3_outputs(3837) <= a;
    layer3_outputs(3838) <= not b;
    layer3_outputs(3839) <= b;
    layer3_outputs(3840) <= a and not b;
    layer3_outputs(3841) <= '0';
    layer3_outputs(3842) <= not a or b;
    layer3_outputs(3843) <= not (a and b);
    layer3_outputs(3844) <= b and not a;
    layer3_outputs(3845) <= a;
    layer3_outputs(3846) <= not a or b;
    layer3_outputs(3847) <= b and not a;
    layer3_outputs(3848) <= not b or a;
    layer3_outputs(3849) <= '1';
    layer3_outputs(3850) <= not a or b;
    layer3_outputs(3851) <= b and not a;
    layer3_outputs(3852) <= '1';
    layer3_outputs(3853) <= b;
    layer3_outputs(3854) <= a and not b;
    layer3_outputs(3855) <= b;
    layer3_outputs(3856) <= not b or a;
    layer3_outputs(3857) <= not b or a;
    layer3_outputs(3858) <= b and not a;
    layer3_outputs(3859) <= a and not b;
    layer3_outputs(3860) <= not (a xor b);
    layer3_outputs(3861) <= not (a or b);
    layer3_outputs(3862) <= not a or b;
    layer3_outputs(3863) <= '1';
    layer3_outputs(3864) <= not (a and b);
    layer3_outputs(3865) <= not (a xor b);
    layer3_outputs(3866) <= not b;
    layer3_outputs(3867) <= not a or b;
    layer3_outputs(3868) <= a or b;
    layer3_outputs(3869) <= b and not a;
    layer3_outputs(3870) <= not (a or b);
    layer3_outputs(3871) <= not (a and b);
    layer3_outputs(3872) <= not b;
    layer3_outputs(3873) <= not a or b;
    layer3_outputs(3874) <= a and not b;
    layer3_outputs(3875) <= a or b;
    layer3_outputs(3876) <= '1';
    layer3_outputs(3877) <= a or b;
    layer3_outputs(3878) <= a;
    layer3_outputs(3879) <= '1';
    layer3_outputs(3880) <= b;
    layer3_outputs(3881) <= not (a and b);
    layer3_outputs(3882) <= not b or a;
    layer3_outputs(3883) <= not b or a;
    layer3_outputs(3884) <= b and not a;
    layer3_outputs(3885) <= '0';
    layer3_outputs(3886) <= b;
    layer3_outputs(3887) <= a or b;
    layer3_outputs(3888) <= not (a or b);
    layer3_outputs(3889) <= not (a or b);
    layer3_outputs(3890) <= not (a and b);
    layer3_outputs(3891) <= '1';
    layer3_outputs(3892) <= not (a or b);
    layer3_outputs(3893) <= not a or b;
    layer3_outputs(3894) <= not (a and b);
    layer3_outputs(3895) <= not a or b;
    layer3_outputs(3896) <= a and b;
    layer3_outputs(3897) <= a xor b;
    layer3_outputs(3898) <= not b;
    layer3_outputs(3899) <= b;
    layer3_outputs(3900) <= a and not b;
    layer3_outputs(3901) <= not b or a;
    layer3_outputs(3902) <= '1';
    layer3_outputs(3903) <= a or b;
    layer3_outputs(3904) <= not a or b;
    layer3_outputs(3905) <= not a or b;
    layer3_outputs(3906) <= b and not a;
    layer3_outputs(3907) <= a xor b;
    layer3_outputs(3908) <= a and b;
    layer3_outputs(3909) <= '1';
    layer3_outputs(3910) <= not b;
    layer3_outputs(3911) <= not (a and b);
    layer3_outputs(3912) <= not a or b;
    layer3_outputs(3913) <= a;
    layer3_outputs(3914) <= not (a and b);
    layer3_outputs(3915) <= not (a and b);
    layer3_outputs(3916) <= '0';
    layer3_outputs(3917) <= not a or b;
    layer3_outputs(3918) <= a;
    layer3_outputs(3919) <= not a;
    layer3_outputs(3920) <= a;
    layer3_outputs(3921) <= '1';
    layer3_outputs(3922) <= a or b;
    layer3_outputs(3923) <= not a or b;
    layer3_outputs(3924) <= b;
    layer3_outputs(3925) <= '1';
    layer3_outputs(3926) <= '1';
    layer3_outputs(3927) <= a and not b;
    layer3_outputs(3928) <= not (a and b);
    layer3_outputs(3929) <= not (a and b);
    layer3_outputs(3930) <= not (a xor b);
    layer3_outputs(3931) <= '0';
    layer3_outputs(3932) <= not b or a;
    layer3_outputs(3933) <= a and not b;
    layer3_outputs(3934) <= a or b;
    layer3_outputs(3935) <= '1';
    layer3_outputs(3936) <= not (a xor b);
    layer3_outputs(3937) <= a and not b;
    layer3_outputs(3938) <= a or b;
    layer3_outputs(3939) <= not (a xor b);
    layer3_outputs(3940) <= a;
    layer3_outputs(3941) <= a and b;
    layer3_outputs(3942) <= not a or b;
    layer3_outputs(3943) <= '1';
    layer3_outputs(3944) <= b;
    layer3_outputs(3945) <= b and not a;
    layer3_outputs(3946) <= not b;
    layer3_outputs(3947) <= not (a xor b);
    layer3_outputs(3948) <= b;
    layer3_outputs(3949) <= a and not b;
    layer3_outputs(3950) <= a or b;
    layer3_outputs(3951) <= b and not a;
    layer3_outputs(3952) <= not a or b;
    layer3_outputs(3953) <= not a;
    layer3_outputs(3954) <= not (a or b);
    layer3_outputs(3955) <= a or b;
    layer3_outputs(3956) <= '0';
    layer3_outputs(3957) <= not b or a;
    layer3_outputs(3958) <= a or b;
    layer3_outputs(3959) <= not a;
    layer3_outputs(3960) <= b;
    layer3_outputs(3961) <= not b or a;
    layer3_outputs(3962) <= a;
    layer3_outputs(3963) <= b;
    layer3_outputs(3964) <= b;
    layer3_outputs(3965) <= a and not b;
    layer3_outputs(3966) <= a or b;
    layer3_outputs(3967) <= not b;
    layer3_outputs(3968) <= '0';
    layer3_outputs(3969) <= b;
    layer3_outputs(3970) <= a or b;
    layer3_outputs(3971) <= not b;
    layer3_outputs(3972) <= '0';
    layer3_outputs(3973) <= not (a and b);
    layer3_outputs(3974) <= a or b;
    layer3_outputs(3975) <= a and not b;
    layer3_outputs(3976) <= not b;
    layer3_outputs(3977) <= not b;
    layer3_outputs(3978) <= not b or a;
    layer3_outputs(3979) <= a;
    layer3_outputs(3980) <= b;
    layer3_outputs(3981) <= not a;
    layer3_outputs(3982) <= a or b;
    layer3_outputs(3983) <= not (a and b);
    layer3_outputs(3984) <= not b or a;
    layer3_outputs(3985) <= a;
    layer3_outputs(3986) <= not a;
    layer3_outputs(3987) <= not (a xor b);
    layer3_outputs(3988) <= '0';
    layer3_outputs(3989) <= b and not a;
    layer3_outputs(3990) <= not a;
    layer3_outputs(3991) <= '0';
    layer3_outputs(3992) <= '1';
    layer3_outputs(3993) <= a xor b;
    layer3_outputs(3994) <= a or b;
    layer3_outputs(3995) <= '0';
    layer3_outputs(3996) <= b;
    layer3_outputs(3997) <= b and not a;
    layer3_outputs(3998) <= not b;
    layer3_outputs(3999) <= not a or b;
    layer3_outputs(4000) <= a or b;
    layer3_outputs(4001) <= not b or a;
    layer3_outputs(4002) <= a;
    layer3_outputs(4003) <= not (a and b);
    layer3_outputs(4004) <= b and not a;
    layer3_outputs(4005) <= not (a or b);
    layer3_outputs(4006) <= b;
    layer3_outputs(4007) <= not b;
    layer3_outputs(4008) <= a and b;
    layer3_outputs(4009) <= not (a or b);
    layer3_outputs(4010) <= not a;
    layer3_outputs(4011) <= b;
    layer3_outputs(4012) <= not b;
    layer3_outputs(4013) <= not b;
    layer3_outputs(4014) <= not a or b;
    layer3_outputs(4015) <= not b;
    layer3_outputs(4016) <= b;
    layer3_outputs(4017) <= not a;
    layer3_outputs(4018) <= a and not b;
    layer3_outputs(4019) <= a xor b;
    layer3_outputs(4020) <= not (a or b);
    layer3_outputs(4021) <= a;
    layer3_outputs(4022) <= not (a xor b);
    layer3_outputs(4023) <= '1';
    layer3_outputs(4024) <= b and not a;
    layer3_outputs(4025) <= not (a xor b);
    layer3_outputs(4026) <= a and b;
    layer3_outputs(4027) <= '1';
    layer3_outputs(4028) <= a or b;
    layer3_outputs(4029) <= b;
    layer3_outputs(4030) <= a and not b;
    layer3_outputs(4031) <= b and not a;
    layer3_outputs(4032) <= a and not b;
    layer3_outputs(4033) <= '0';
    layer3_outputs(4034) <= a and b;
    layer3_outputs(4035) <= a and b;
    layer3_outputs(4036) <= not (a and b);
    layer3_outputs(4037) <= not b or a;
    layer3_outputs(4038) <= not a or b;
    layer3_outputs(4039) <= a xor b;
    layer3_outputs(4040) <= b;
    layer3_outputs(4041) <= a;
    layer3_outputs(4042) <= not (a and b);
    layer3_outputs(4043) <= b;
    layer3_outputs(4044) <= a;
    layer3_outputs(4045) <= a and b;
    layer3_outputs(4046) <= not (a or b);
    layer3_outputs(4047) <= not a or b;
    layer3_outputs(4048) <= not (a xor b);
    layer3_outputs(4049) <= not b;
    layer3_outputs(4050) <= not b or a;
    layer3_outputs(4051) <= a;
    layer3_outputs(4052) <= not (a and b);
    layer3_outputs(4053) <= not a or b;
    layer3_outputs(4054) <= a and b;
    layer3_outputs(4055) <= b;
    layer3_outputs(4056) <= not a or b;
    layer3_outputs(4057) <= '1';
    layer3_outputs(4058) <= not a or b;
    layer3_outputs(4059) <= not (a or b);
    layer3_outputs(4060) <= a and not b;
    layer3_outputs(4061) <= a and b;
    layer3_outputs(4062) <= a;
    layer3_outputs(4063) <= a and not b;
    layer3_outputs(4064) <= '0';
    layer3_outputs(4065) <= b;
    layer3_outputs(4066) <= a and b;
    layer3_outputs(4067) <= not b or a;
    layer3_outputs(4068) <= b;
    layer3_outputs(4069) <= not a or b;
    layer3_outputs(4070) <= not b;
    layer3_outputs(4071) <= '0';
    layer3_outputs(4072) <= not b or a;
    layer3_outputs(4073) <= '0';
    layer3_outputs(4074) <= a;
    layer3_outputs(4075) <= not b or a;
    layer3_outputs(4076) <= not b;
    layer3_outputs(4077) <= not (a or b);
    layer3_outputs(4078) <= not a;
    layer3_outputs(4079) <= not b;
    layer3_outputs(4080) <= not (a and b);
    layer3_outputs(4081) <= not b;
    layer3_outputs(4082) <= '1';
    layer3_outputs(4083) <= '1';
    layer3_outputs(4084) <= not b;
    layer3_outputs(4085) <= not b;
    layer3_outputs(4086) <= not (a and b);
    layer3_outputs(4087) <= not a or b;
    layer3_outputs(4088) <= a and not b;
    layer3_outputs(4089) <= b;
    layer3_outputs(4090) <= a and b;
    layer3_outputs(4091) <= '0';
    layer3_outputs(4092) <= a xor b;
    layer3_outputs(4093) <= a or b;
    layer3_outputs(4094) <= not (a or b);
    layer3_outputs(4095) <= b;
    layer3_outputs(4096) <= '1';
    layer3_outputs(4097) <= b;
    layer3_outputs(4098) <= not (a and b);
    layer3_outputs(4099) <= b;
    layer3_outputs(4100) <= a and b;
    layer3_outputs(4101) <= not b or a;
    layer3_outputs(4102) <= not b or a;
    layer3_outputs(4103) <= not a;
    layer3_outputs(4104) <= b and not a;
    layer3_outputs(4105) <= a and not b;
    layer3_outputs(4106) <= a or b;
    layer3_outputs(4107) <= not (a and b);
    layer3_outputs(4108) <= not (a and b);
    layer3_outputs(4109) <= not (a and b);
    layer3_outputs(4110) <= not a or b;
    layer3_outputs(4111) <= b and not a;
    layer3_outputs(4112) <= a xor b;
    layer3_outputs(4113) <= b;
    layer3_outputs(4114) <= a;
    layer3_outputs(4115) <= not (a or b);
    layer3_outputs(4116) <= not (a or b);
    layer3_outputs(4117) <= '0';
    layer3_outputs(4118) <= not a or b;
    layer3_outputs(4119) <= not (a or b);
    layer3_outputs(4120) <= a and not b;
    layer3_outputs(4121) <= b;
    layer3_outputs(4122) <= not (a and b);
    layer3_outputs(4123) <= not b or a;
    layer3_outputs(4124) <= not (a and b);
    layer3_outputs(4125) <= not (a and b);
    layer3_outputs(4126) <= not b or a;
    layer3_outputs(4127) <= not b;
    layer3_outputs(4128) <= a and b;
    layer3_outputs(4129) <= not b;
    layer3_outputs(4130) <= '0';
    layer3_outputs(4131) <= a or b;
    layer3_outputs(4132) <= not b or a;
    layer3_outputs(4133) <= not (a and b);
    layer3_outputs(4134) <= not b;
    layer3_outputs(4135) <= not (a and b);
    layer3_outputs(4136) <= '0';
    layer3_outputs(4137) <= a and not b;
    layer3_outputs(4138) <= a;
    layer3_outputs(4139) <= b;
    layer3_outputs(4140) <= not (a or b);
    layer3_outputs(4141) <= a;
    layer3_outputs(4142) <= a and not b;
    layer3_outputs(4143) <= '1';
    layer3_outputs(4144) <= '0';
    layer3_outputs(4145) <= a and not b;
    layer3_outputs(4146) <= not (a xor b);
    layer3_outputs(4147) <= a and b;
    layer3_outputs(4148) <= a and not b;
    layer3_outputs(4149) <= a and not b;
    layer3_outputs(4150) <= not b or a;
    layer3_outputs(4151) <= a and not b;
    layer3_outputs(4152) <= a and not b;
    layer3_outputs(4153) <= not (a xor b);
    layer3_outputs(4154) <= '1';
    layer3_outputs(4155) <= not b or a;
    layer3_outputs(4156) <= b and not a;
    layer3_outputs(4157) <= a or b;
    layer3_outputs(4158) <= b and not a;
    layer3_outputs(4159) <= not a;
    layer3_outputs(4160) <= a and not b;
    layer3_outputs(4161) <= not b;
    layer3_outputs(4162) <= not (a or b);
    layer3_outputs(4163) <= not a or b;
    layer3_outputs(4164) <= not (a or b);
    layer3_outputs(4165) <= b;
    layer3_outputs(4166) <= b and not a;
    layer3_outputs(4167) <= a or b;
    layer3_outputs(4168) <= a;
    layer3_outputs(4169) <= not a;
    layer3_outputs(4170) <= '1';
    layer3_outputs(4171) <= a and b;
    layer3_outputs(4172) <= '1';
    layer3_outputs(4173) <= not a or b;
    layer3_outputs(4174) <= not b;
    layer3_outputs(4175) <= b;
    layer3_outputs(4176) <= not b or a;
    layer3_outputs(4177) <= not b or a;
    layer3_outputs(4178) <= '1';
    layer3_outputs(4179) <= not b or a;
    layer3_outputs(4180) <= not a or b;
    layer3_outputs(4181) <= a and b;
    layer3_outputs(4182) <= b and not a;
    layer3_outputs(4183) <= b;
    layer3_outputs(4184) <= not (a and b);
    layer3_outputs(4185) <= not (a or b);
    layer3_outputs(4186) <= not a or b;
    layer3_outputs(4187) <= a and b;
    layer3_outputs(4188) <= a or b;
    layer3_outputs(4189) <= a and not b;
    layer3_outputs(4190) <= '0';
    layer3_outputs(4191) <= a;
    layer3_outputs(4192) <= not a;
    layer3_outputs(4193) <= not (a or b);
    layer3_outputs(4194) <= '1';
    layer3_outputs(4195) <= b;
    layer3_outputs(4196) <= not a;
    layer3_outputs(4197) <= '1';
    layer3_outputs(4198) <= not a or b;
    layer3_outputs(4199) <= a or b;
    layer3_outputs(4200) <= a;
    layer3_outputs(4201) <= not (a and b);
    layer3_outputs(4202) <= '1';
    layer3_outputs(4203) <= '0';
    layer3_outputs(4204) <= a and not b;
    layer3_outputs(4205) <= not b;
    layer3_outputs(4206) <= a;
    layer3_outputs(4207) <= a and not b;
    layer3_outputs(4208) <= '1';
    layer3_outputs(4209) <= b and not a;
    layer3_outputs(4210) <= a and not b;
    layer3_outputs(4211) <= not b;
    layer3_outputs(4212) <= b and not a;
    layer3_outputs(4213) <= a;
    layer3_outputs(4214) <= not b;
    layer3_outputs(4215) <= a xor b;
    layer3_outputs(4216) <= a xor b;
    layer3_outputs(4217) <= not a or b;
    layer3_outputs(4218) <= a;
    layer3_outputs(4219) <= a;
    layer3_outputs(4220) <= a;
    layer3_outputs(4221) <= not b;
    layer3_outputs(4222) <= a or b;
    layer3_outputs(4223) <= not b;
    layer3_outputs(4224) <= not a;
    layer3_outputs(4225) <= a xor b;
    layer3_outputs(4226) <= a and b;
    layer3_outputs(4227) <= '1';
    layer3_outputs(4228) <= not a;
    layer3_outputs(4229) <= '0';
    layer3_outputs(4230) <= '0';
    layer3_outputs(4231) <= not (a and b);
    layer3_outputs(4232) <= '0';
    layer3_outputs(4233) <= b;
    layer3_outputs(4234) <= b and not a;
    layer3_outputs(4235) <= a;
    layer3_outputs(4236) <= not (a and b);
    layer3_outputs(4237) <= not a;
    layer3_outputs(4238) <= not (a and b);
    layer3_outputs(4239) <= b and not a;
    layer3_outputs(4240) <= a or b;
    layer3_outputs(4241) <= not a or b;
    layer3_outputs(4242) <= not a;
    layer3_outputs(4243) <= not b or a;
    layer3_outputs(4244) <= a and b;
    layer3_outputs(4245) <= not b;
    layer3_outputs(4246) <= not b or a;
    layer3_outputs(4247) <= not b or a;
    layer3_outputs(4248) <= not b or a;
    layer3_outputs(4249) <= a and b;
    layer3_outputs(4250) <= not a or b;
    layer3_outputs(4251) <= a;
    layer3_outputs(4252) <= not (a and b);
    layer3_outputs(4253) <= not b;
    layer3_outputs(4254) <= not b or a;
    layer3_outputs(4255) <= a xor b;
    layer3_outputs(4256) <= not a;
    layer3_outputs(4257) <= not b or a;
    layer3_outputs(4258) <= not a;
    layer3_outputs(4259) <= '0';
    layer3_outputs(4260) <= a and b;
    layer3_outputs(4261) <= not a;
    layer3_outputs(4262) <= not a or b;
    layer3_outputs(4263) <= b and not a;
    layer3_outputs(4264) <= '0';
    layer3_outputs(4265) <= not b or a;
    layer3_outputs(4266) <= b;
    layer3_outputs(4267) <= b;
    layer3_outputs(4268) <= a or b;
    layer3_outputs(4269) <= a xor b;
    layer3_outputs(4270) <= a and b;
    layer3_outputs(4271) <= '0';
    layer3_outputs(4272) <= b and not a;
    layer3_outputs(4273) <= b and not a;
    layer3_outputs(4274) <= a xor b;
    layer3_outputs(4275) <= not (a and b);
    layer3_outputs(4276) <= not (a xor b);
    layer3_outputs(4277) <= b and not a;
    layer3_outputs(4278) <= not (a and b);
    layer3_outputs(4279) <= not (a xor b);
    layer3_outputs(4280) <= not (a xor b);
    layer3_outputs(4281) <= '0';
    layer3_outputs(4282) <= a or b;
    layer3_outputs(4283) <= b;
    layer3_outputs(4284) <= a;
    layer3_outputs(4285) <= a xor b;
    layer3_outputs(4286) <= a;
    layer3_outputs(4287) <= b and not a;
    layer3_outputs(4288) <= a xor b;
    layer3_outputs(4289) <= a or b;
    layer3_outputs(4290) <= b and not a;
    layer3_outputs(4291) <= a and b;
    layer3_outputs(4292) <= not b;
    layer3_outputs(4293) <= not (a or b);
    layer3_outputs(4294) <= a and not b;
    layer3_outputs(4295) <= a and not b;
    layer3_outputs(4296) <= not (a and b);
    layer3_outputs(4297) <= a or b;
    layer3_outputs(4298) <= a and not b;
    layer3_outputs(4299) <= a and b;
    layer3_outputs(4300) <= not a or b;
    layer3_outputs(4301) <= '0';
    layer3_outputs(4302) <= not b or a;
    layer3_outputs(4303) <= b;
    layer3_outputs(4304) <= a and not b;
    layer3_outputs(4305) <= a or b;
    layer3_outputs(4306) <= a and b;
    layer3_outputs(4307) <= not a or b;
    layer3_outputs(4308) <= '1';
    layer3_outputs(4309) <= not (a or b);
    layer3_outputs(4310) <= not a;
    layer3_outputs(4311) <= b;
    layer3_outputs(4312) <= '0';
    layer3_outputs(4313) <= not (a or b);
    layer3_outputs(4314) <= '0';
    layer3_outputs(4315) <= not (a xor b);
    layer3_outputs(4316) <= not b or a;
    layer3_outputs(4317) <= not (a or b);
    layer3_outputs(4318) <= a and b;
    layer3_outputs(4319) <= not a;
    layer3_outputs(4320) <= a or b;
    layer3_outputs(4321) <= not (a or b);
    layer3_outputs(4322) <= not b;
    layer3_outputs(4323) <= not b;
    layer3_outputs(4324) <= not b;
    layer3_outputs(4325) <= not (a or b);
    layer3_outputs(4326) <= not a;
    layer3_outputs(4327) <= '0';
    layer3_outputs(4328) <= a;
    layer3_outputs(4329) <= a and not b;
    layer3_outputs(4330) <= not b or a;
    layer3_outputs(4331) <= not b or a;
    layer3_outputs(4332) <= not a;
    layer3_outputs(4333) <= not a or b;
    layer3_outputs(4334) <= a xor b;
    layer3_outputs(4335) <= not a;
    layer3_outputs(4336) <= not b;
    layer3_outputs(4337) <= not a;
    layer3_outputs(4338) <= '1';
    layer3_outputs(4339) <= not b;
    layer3_outputs(4340) <= a or b;
    layer3_outputs(4341) <= not (a or b);
    layer3_outputs(4342) <= b and not a;
    layer3_outputs(4343) <= a and not b;
    layer3_outputs(4344) <= a;
    layer3_outputs(4345) <= not b;
    layer3_outputs(4346) <= a;
    layer3_outputs(4347) <= a and not b;
    layer3_outputs(4348) <= a or b;
    layer3_outputs(4349) <= not b or a;
    layer3_outputs(4350) <= not a or b;
    layer3_outputs(4351) <= '1';
    layer3_outputs(4352) <= not (a and b);
    layer3_outputs(4353) <= a and b;
    layer3_outputs(4354) <= not a or b;
    layer3_outputs(4355) <= b;
    layer3_outputs(4356) <= not a or b;
    layer3_outputs(4357) <= a;
    layer3_outputs(4358) <= '1';
    layer3_outputs(4359) <= '0';
    layer3_outputs(4360) <= b;
    layer3_outputs(4361) <= a and b;
    layer3_outputs(4362) <= not (a or b);
    layer3_outputs(4363) <= a and not b;
    layer3_outputs(4364) <= '0';
    layer3_outputs(4365) <= not b;
    layer3_outputs(4366) <= not (a and b);
    layer3_outputs(4367) <= '0';
    layer3_outputs(4368) <= not a or b;
    layer3_outputs(4369) <= '1';
    layer3_outputs(4370) <= not a;
    layer3_outputs(4371) <= not a or b;
    layer3_outputs(4372) <= a;
    layer3_outputs(4373) <= not (a or b);
    layer3_outputs(4374) <= not a or b;
    layer3_outputs(4375) <= not a or b;
    layer3_outputs(4376) <= '0';
    layer3_outputs(4377) <= a and not b;
    layer3_outputs(4378) <= not b or a;
    layer3_outputs(4379) <= a or b;
    layer3_outputs(4380) <= b;
    layer3_outputs(4381) <= '0';
    layer3_outputs(4382) <= a or b;
    layer3_outputs(4383) <= a and not b;
    layer3_outputs(4384) <= '1';
    layer3_outputs(4385) <= not (a xor b);
    layer3_outputs(4386) <= a or b;
    layer3_outputs(4387) <= a;
    layer3_outputs(4388) <= not (a and b);
    layer3_outputs(4389) <= a and not b;
    layer3_outputs(4390) <= a and b;
    layer3_outputs(4391) <= not (a and b);
    layer3_outputs(4392) <= not b or a;
    layer3_outputs(4393) <= a and not b;
    layer3_outputs(4394) <= a;
    layer3_outputs(4395) <= not a;
    layer3_outputs(4396) <= a;
    layer3_outputs(4397) <= not a;
    layer3_outputs(4398) <= not (a or b);
    layer3_outputs(4399) <= a and b;
    layer3_outputs(4400) <= not a;
    layer3_outputs(4401) <= b;
    layer3_outputs(4402) <= '0';
    layer3_outputs(4403) <= not (a xor b);
    layer3_outputs(4404) <= not (a and b);
    layer3_outputs(4405) <= a xor b;
    layer3_outputs(4406) <= not b or a;
    layer3_outputs(4407) <= not a or b;
    layer3_outputs(4408) <= '1';
    layer3_outputs(4409) <= a and b;
    layer3_outputs(4410) <= a;
    layer3_outputs(4411) <= not (a and b);
    layer3_outputs(4412) <= not b;
    layer3_outputs(4413) <= a and b;
    layer3_outputs(4414) <= b;
    layer3_outputs(4415) <= a and not b;
    layer3_outputs(4416) <= a and not b;
    layer3_outputs(4417) <= '0';
    layer3_outputs(4418) <= not b;
    layer3_outputs(4419) <= a or b;
    layer3_outputs(4420) <= '1';
    layer3_outputs(4421) <= not (a xor b);
    layer3_outputs(4422) <= not b or a;
    layer3_outputs(4423) <= not a or b;
    layer3_outputs(4424) <= not a or b;
    layer3_outputs(4425) <= a;
    layer3_outputs(4426) <= not b or a;
    layer3_outputs(4427) <= '0';
    layer3_outputs(4428) <= not (a or b);
    layer3_outputs(4429) <= not a;
    layer3_outputs(4430) <= a and not b;
    layer3_outputs(4431) <= not (a or b);
    layer3_outputs(4432) <= '1';
    layer3_outputs(4433) <= '0';
    layer3_outputs(4434) <= not (a xor b);
    layer3_outputs(4435) <= a or b;
    layer3_outputs(4436) <= not (a and b);
    layer3_outputs(4437) <= not (a or b);
    layer3_outputs(4438) <= not a;
    layer3_outputs(4439) <= b;
    layer3_outputs(4440) <= a and b;
    layer3_outputs(4441) <= b and not a;
    layer3_outputs(4442) <= not a or b;
    layer3_outputs(4443) <= b;
    layer3_outputs(4444) <= a and not b;
    layer3_outputs(4445) <= '0';
    layer3_outputs(4446) <= not b or a;
    layer3_outputs(4447) <= a;
    layer3_outputs(4448) <= a and b;
    layer3_outputs(4449) <= not (a or b);
    layer3_outputs(4450) <= b and not a;
    layer3_outputs(4451) <= b;
    layer3_outputs(4452) <= not b or a;
    layer3_outputs(4453) <= a and not b;
    layer3_outputs(4454) <= a;
    layer3_outputs(4455) <= not b;
    layer3_outputs(4456) <= '0';
    layer3_outputs(4457) <= not a or b;
    layer3_outputs(4458) <= not b or a;
    layer3_outputs(4459) <= a;
    layer3_outputs(4460) <= a and not b;
    layer3_outputs(4461) <= '1';
    layer3_outputs(4462) <= b and not a;
    layer3_outputs(4463) <= not b or a;
    layer3_outputs(4464) <= b and not a;
    layer3_outputs(4465) <= not (a and b);
    layer3_outputs(4466) <= not (a or b);
    layer3_outputs(4467) <= b and not a;
    layer3_outputs(4468) <= '1';
    layer3_outputs(4469) <= not (a and b);
    layer3_outputs(4470) <= b and not a;
    layer3_outputs(4471) <= not a;
    layer3_outputs(4472) <= '0';
    layer3_outputs(4473) <= not (a and b);
    layer3_outputs(4474) <= not b;
    layer3_outputs(4475) <= not b;
    layer3_outputs(4476) <= not (a and b);
    layer3_outputs(4477) <= '1';
    layer3_outputs(4478) <= not a or b;
    layer3_outputs(4479) <= not b or a;
    layer3_outputs(4480) <= a and b;
    layer3_outputs(4481) <= not b;
    layer3_outputs(4482) <= not a or b;
    layer3_outputs(4483) <= not (a and b);
    layer3_outputs(4484) <= not b;
    layer3_outputs(4485) <= not a or b;
    layer3_outputs(4486) <= not (a or b);
    layer3_outputs(4487) <= b;
    layer3_outputs(4488) <= not a;
    layer3_outputs(4489) <= not a;
    layer3_outputs(4490) <= '0';
    layer3_outputs(4491) <= not (a and b);
    layer3_outputs(4492) <= '1';
    layer3_outputs(4493) <= not a;
    layer3_outputs(4494) <= not b or a;
    layer3_outputs(4495) <= b;
    layer3_outputs(4496) <= a and b;
    layer3_outputs(4497) <= a and b;
    layer3_outputs(4498) <= '0';
    layer3_outputs(4499) <= a and not b;
    layer3_outputs(4500) <= not (a xor b);
    layer3_outputs(4501) <= not (a or b);
    layer3_outputs(4502) <= not (a and b);
    layer3_outputs(4503) <= a;
    layer3_outputs(4504) <= not (a and b);
    layer3_outputs(4505) <= a and b;
    layer3_outputs(4506) <= not a or b;
    layer3_outputs(4507) <= not a;
    layer3_outputs(4508) <= not b;
    layer3_outputs(4509) <= not a or b;
    layer3_outputs(4510) <= not (a and b);
    layer3_outputs(4511) <= a;
    layer3_outputs(4512) <= not (a and b);
    layer3_outputs(4513) <= a or b;
    layer3_outputs(4514) <= not a;
    layer3_outputs(4515) <= '1';
    layer3_outputs(4516) <= not a;
    layer3_outputs(4517) <= not b;
    layer3_outputs(4518) <= a xor b;
    layer3_outputs(4519) <= not (a or b);
    layer3_outputs(4520) <= not b;
    layer3_outputs(4521) <= not (a or b);
    layer3_outputs(4522) <= a and b;
    layer3_outputs(4523) <= not a;
    layer3_outputs(4524) <= not (a and b);
    layer3_outputs(4525) <= not a or b;
    layer3_outputs(4526) <= b;
    layer3_outputs(4527) <= not b;
    layer3_outputs(4528) <= not b;
    layer3_outputs(4529) <= '1';
    layer3_outputs(4530) <= not a;
    layer3_outputs(4531) <= not (a or b);
    layer3_outputs(4532) <= not a or b;
    layer3_outputs(4533) <= a or b;
    layer3_outputs(4534) <= not (a and b);
    layer3_outputs(4535) <= not a;
    layer3_outputs(4536) <= not (a or b);
    layer3_outputs(4537) <= not (a or b);
    layer3_outputs(4538) <= b and not a;
    layer3_outputs(4539) <= b and not a;
    layer3_outputs(4540) <= b;
    layer3_outputs(4541) <= not b or a;
    layer3_outputs(4542) <= a xor b;
    layer3_outputs(4543) <= b;
    layer3_outputs(4544) <= a and b;
    layer3_outputs(4545) <= not b;
    layer3_outputs(4546) <= not a;
    layer3_outputs(4547) <= a and b;
    layer3_outputs(4548) <= '1';
    layer3_outputs(4549) <= b;
    layer3_outputs(4550) <= not b or a;
    layer3_outputs(4551) <= '0';
    layer3_outputs(4552) <= not b;
    layer3_outputs(4553) <= '0';
    layer3_outputs(4554) <= '1';
    layer3_outputs(4555) <= b;
    layer3_outputs(4556) <= '1';
    layer3_outputs(4557) <= a;
    layer3_outputs(4558) <= not (a and b);
    layer3_outputs(4559) <= b;
    layer3_outputs(4560) <= not a;
    layer3_outputs(4561) <= not a or b;
    layer3_outputs(4562) <= '0';
    layer3_outputs(4563) <= '1';
    layer3_outputs(4564) <= a and b;
    layer3_outputs(4565) <= a and b;
    layer3_outputs(4566) <= a and b;
    layer3_outputs(4567) <= '0';
    layer3_outputs(4568) <= a or b;
    layer3_outputs(4569) <= '0';
    layer3_outputs(4570) <= a;
    layer3_outputs(4571) <= a and not b;
    layer3_outputs(4572) <= a or b;
    layer3_outputs(4573) <= not a;
    layer3_outputs(4574) <= b and not a;
    layer3_outputs(4575) <= not (a or b);
    layer3_outputs(4576) <= not (a and b);
    layer3_outputs(4577) <= a xor b;
    layer3_outputs(4578) <= b;
    layer3_outputs(4579) <= a;
    layer3_outputs(4580) <= a and b;
    layer3_outputs(4581) <= a and b;
    layer3_outputs(4582) <= a and not b;
    layer3_outputs(4583) <= not b or a;
    layer3_outputs(4584) <= not a or b;
    layer3_outputs(4585) <= not (a and b);
    layer3_outputs(4586) <= a and b;
    layer3_outputs(4587) <= '0';
    layer3_outputs(4588) <= not b;
    layer3_outputs(4589) <= '1';
    layer3_outputs(4590) <= not a;
    layer3_outputs(4591) <= not a or b;
    layer3_outputs(4592) <= not a or b;
    layer3_outputs(4593) <= b;
    layer3_outputs(4594) <= b and not a;
    layer3_outputs(4595) <= a and not b;
    layer3_outputs(4596) <= a or b;
    layer3_outputs(4597) <= a and not b;
    layer3_outputs(4598) <= not (a or b);
    layer3_outputs(4599) <= a and not b;
    layer3_outputs(4600) <= '1';
    layer3_outputs(4601) <= not (a and b);
    layer3_outputs(4602) <= not a;
    layer3_outputs(4603) <= not b;
    layer3_outputs(4604) <= a and b;
    layer3_outputs(4605) <= b;
    layer3_outputs(4606) <= a or b;
    layer3_outputs(4607) <= not b or a;
    layer3_outputs(4608) <= not b or a;
    layer3_outputs(4609) <= not (a xor b);
    layer3_outputs(4610) <= b;
    layer3_outputs(4611) <= not b or a;
    layer3_outputs(4612) <= not (a or b);
    layer3_outputs(4613) <= not (a or b);
    layer3_outputs(4614) <= not a;
    layer3_outputs(4615) <= a and b;
    layer3_outputs(4616) <= b;
    layer3_outputs(4617) <= not a or b;
    layer3_outputs(4618) <= a or b;
    layer3_outputs(4619) <= not (a or b);
    layer3_outputs(4620) <= a and not b;
    layer3_outputs(4621) <= not (a or b);
    layer3_outputs(4622) <= b;
    layer3_outputs(4623) <= a xor b;
    layer3_outputs(4624) <= a or b;
    layer3_outputs(4625) <= '0';
    layer3_outputs(4626) <= a or b;
    layer3_outputs(4627) <= b and not a;
    layer3_outputs(4628) <= not b or a;
    layer3_outputs(4629) <= a and not b;
    layer3_outputs(4630) <= not b or a;
    layer3_outputs(4631) <= not (a or b);
    layer3_outputs(4632) <= not a;
    layer3_outputs(4633) <= not a or b;
    layer3_outputs(4634) <= not (a and b);
    layer3_outputs(4635) <= not b or a;
    layer3_outputs(4636) <= a or b;
    layer3_outputs(4637) <= not (a or b);
    layer3_outputs(4638) <= '0';
    layer3_outputs(4639) <= a and b;
    layer3_outputs(4640) <= not (a and b);
    layer3_outputs(4641) <= a;
    layer3_outputs(4642) <= not (a or b);
    layer3_outputs(4643) <= not a;
    layer3_outputs(4644) <= not a;
    layer3_outputs(4645) <= '1';
    layer3_outputs(4646) <= '1';
    layer3_outputs(4647) <= b and not a;
    layer3_outputs(4648) <= not (a and b);
    layer3_outputs(4649) <= a or b;
    layer3_outputs(4650) <= a and b;
    layer3_outputs(4651) <= a xor b;
    layer3_outputs(4652) <= b;
    layer3_outputs(4653) <= not b;
    layer3_outputs(4654) <= not b or a;
    layer3_outputs(4655) <= not b;
    layer3_outputs(4656) <= '1';
    layer3_outputs(4657) <= not b or a;
    layer3_outputs(4658) <= a and b;
    layer3_outputs(4659) <= a or b;
    layer3_outputs(4660) <= a xor b;
    layer3_outputs(4661) <= a;
    layer3_outputs(4662) <= not a;
    layer3_outputs(4663) <= '1';
    layer3_outputs(4664) <= '1';
    layer3_outputs(4665) <= a and b;
    layer3_outputs(4666) <= not (a or b);
    layer3_outputs(4667) <= '1';
    layer3_outputs(4668) <= b and not a;
    layer3_outputs(4669) <= a and not b;
    layer3_outputs(4670) <= not a or b;
    layer3_outputs(4671) <= not (a and b);
    layer3_outputs(4672) <= not (a and b);
    layer3_outputs(4673) <= '1';
    layer3_outputs(4674) <= a and b;
    layer3_outputs(4675) <= b and not a;
    layer3_outputs(4676) <= a or b;
    layer3_outputs(4677) <= not (a or b);
    layer3_outputs(4678) <= not (a xor b);
    layer3_outputs(4679) <= not a;
    layer3_outputs(4680) <= a and not b;
    layer3_outputs(4681) <= a and b;
    layer3_outputs(4682) <= not a or b;
    layer3_outputs(4683) <= not a or b;
    layer3_outputs(4684) <= not b or a;
    layer3_outputs(4685) <= not b;
    layer3_outputs(4686) <= a or b;
    layer3_outputs(4687) <= b;
    layer3_outputs(4688) <= not b or a;
    layer3_outputs(4689) <= '1';
    layer3_outputs(4690) <= a;
    layer3_outputs(4691) <= '0';
    layer3_outputs(4692) <= not (a or b);
    layer3_outputs(4693) <= b;
    layer3_outputs(4694) <= a;
    layer3_outputs(4695) <= a and not b;
    layer3_outputs(4696) <= not (a and b);
    layer3_outputs(4697) <= not b or a;
    layer3_outputs(4698) <= b and not a;
    layer3_outputs(4699) <= a and b;
    layer3_outputs(4700) <= not (a xor b);
    layer3_outputs(4701) <= a and b;
    layer3_outputs(4702) <= a and not b;
    layer3_outputs(4703) <= not a;
    layer3_outputs(4704) <= not b;
    layer3_outputs(4705) <= not b;
    layer3_outputs(4706) <= not (a and b);
    layer3_outputs(4707) <= '1';
    layer3_outputs(4708) <= not (a xor b);
    layer3_outputs(4709) <= '0';
    layer3_outputs(4710) <= '1';
    layer3_outputs(4711) <= a xor b;
    layer3_outputs(4712) <= not a or b;
    layer3_outputs(4713) <= not b;
    layer3_outputs(4714) <= '1';
    layer3_outputs(4715) <= not (a and b);
    layer3_outputs(4716) <= not b or a;
    layer3_outputs(4717) <= not a or b;
    layer3_outputs(4718) <= a or b;
    layer3_outputs(4719) <= a and b;
    layer3_outputs(4720) <= a and not b;
    layer3_outputs(4721) <= not b;
    layer3_outputs(4722) <= a or b;
    layer3_outputs(4723) <= not (a and b);
    layer3_outputs(4724) <= not b;
    layer3_outputs(4725) <= b;
    layer3_outputs(4726) <= not (a or b);
    layer3_outputs(4727) <= a and not b;
    layer3_outputs(4728) <= b and not a;
    layer3_outputs(4729) <= a and not b;
    layer3_outputs(4730) <= not (a and b);
    layer3_outputs(4731) <= a or b;
    layer3_outputs(4732) <= b;
    layer3_outputs(4733) <= '0';
    layer3_outputs(4734) <= a or b;
    layer3_outputs(4735) <= '1';
    layer3_outputs(4736) <= a;
    layer3_outputs(4737) <= a or b;
    layer3_outputs(4738) <= not (a and b);
    layer3_outputs(4739) <= a;
    layer3_outputs(4740) <= not a;
    layer3_outputs(4741) <= a and not b;
    layer3_outputs(4742) <= b and not a;
    layer3_outputs(4743) <= b;
    layer3_outputs(4744) <= '1';
    layer3_outputs(4745) <= a and b;
    layer3_outputs(4746) <= '1';
    layer3_outputs(4747) <= not (a and b);
    layer3_outputs(4748) <= not b or a;
    layer3_outputs(4749) <= '0';
    layer3_outputs(4750) <= a and b;
    layer3_outputs(4751) <= a;
    layer3_outputs(4752) <= b;
    layer3_outputs(4753) <= a and b;
    layer3_outputs(4754) <= not a or b;
    layer3_outputs(4755) <= not b or a;
    layer3_outputs(4756) <= a;
    layer3_outputs(4757) <= b and not a;
    layer3_outputs(4758) <= '1';
    layer3_outputs(4759) <= not b or a;
    layer3_outputs(4760) <= a and not b;
    layer3_outputs(4761) <= not b;
    layer3_outputs(4762) <= a;
    layer3_outputs(4763) <= not (a or b);
    layer3_outputs(4764) <= b and not a;
    layer3_outputs(4765) <= not (a or b);
    layer3_outputs(4766) <= '0';
    layer3_outputs(4767) <= a or b;
    layer3_outputs(4768) <= b;
    layer3_outputs(4769) <= a;
    layer3_outputs(4770) <= '1';
    layer3_outputs(4771) <= not b or a;
    layer3_outputs(4772) <= not b or a;
    layer3_outputs(4773) <= not b;
    layer3_outputs(4774) <= not (a or b);
    layer3_outputs(4775) <= a;
    layer3_outputs(4776) <= not b;
    layer3_outputs(4777) <= not (a and b);
    layer3_outputs(4778) <= a and not b;
    layer3_outputs(4779) <= not a or b;
    layer3_outputs(4780) <= not (a or b);
    layer3_outputs(4781) <= '0';
    layer3_outputs(4782) <= not a;
    layer3_outputs(4783) <= a and b;
    layer3_outputs(4784) <= not a;
    layer3_outputs(4785) <= a or b;
    layer3_outputs(4786) <= not a or b;
    layer3_outputs(4787) <= not (a or b);
    layer3_outputs(4788) <= not (a and b);
    layer3_outputs(4789) <= not (a and b);
    layer3_outputs(4790) <= not b or a;
    layer3_outputs(4791) <= not (a and b);
    layer3_outputs(4792) <= not b or a;
    layer3_outputs(4793) <= not b;
    layer3_outputs(4794) <= not b;
    layer3_outputs(4795) <= not b;
    layer3_outputs(4796) <= not a;
    layer3_outputs(4797) <= not a;
    layer3_outputs(4798) <= '0';
    layer3_outputs(4799) <= '1';
    layer3_outputs(4800) <= not a or b;
    layer3_outputs(4801) <= not (a and b);
    layer3_outputs(4802) <= not a;
    layer3_outputs(4803) <= '0';
    layer3_outputs(4804) <= '0';
    layer3_outputs(4805) <= '1';
    layer3_outputs(4806) <= not a;
    layer3_outputs(4807) <= '0';
    layer3_outputs(4808) <= '1';
    layer3_outputs(4809) <= not (a or b);
    layer3_outputs(4810) <= '1';
    layer3_outputs(4811) <= not b;
    layer3_outputs(4812) <= a and b;
    layer3_outputs(4813) <= not a or b;
    layer3_outputs(4814) <= not (a and b);
    layer3_outputs(4815) <= not (a or b);
    layer3_outputs(4816) <= a;
    layer3_outputs(4817) <= a and not b;
    layer3_outputs(4818) <= a xor b;
    layer3_outputs(4819) <= not a;
    layer3_outputs(4820) <= a or b;
    layer3_outputs(4821) <= '1';
    layer3_outputs(4822) <= not (a and b);
    layer3_outputs(4823) <= not b;
    layer3_outputs(4824) <= a and b;
    layer3_outputs(4825) <= not a or b;
    layer3_outputs(4826) <= not (a and b);
    layer3_outputs(4827) <= not (a and b);
    layer3_outputs(4828) <= not a;
    layer3_outputs(4829) <= '1';
    layer3_outputs(4830) <= b;
    layer3_outputs(4831) <= not (a and b);
    layer3_outputs(4832) <= b and not a;
    layer3_outputs(4833) <= not a;
    layer3_outputs(4834) <= b and not a;
    layer3_outputs(4835) <= '0';
    layer3_outputs(4836) <= '0';
    layer3_outputs(4837) <= a and b;
    layer3_outputs(4838) <= not (a or b);
    layer3_outputs(4839) <= not (a or b);
    layer3_outputs(4840) <= not a;
    layer3_outputs(4841) <= b and not a;
    layer3_outputs(4842) <= not (a xor b);
    layer3_outputs(4843) <= not (a or b);
    layer3_outputs(4844) <= not b or a;
    layer3_outputs(4845) <= a;
    layer3_outputs(4846) <= not (a or b);
    layer3_outputs(4847) <= a and not b;
    layer3_outputs(4848) <= a xor b;
    layer3_outputs(4849) <= not b;
    layer3_outputs(4850) <= not (a xor b);
    layer3_outputs(4851) <= not b;
    layer3_outputs(4852) <= b and not a;
    layer3_outputs(4853) <= a and not b;
    layer3_outputs(4854) <= b;
    layer3_outputs(4855) <= not (a or b);
    layer3_outputs(4856) <= a and not b;
    layer3_outputs(4857) <= not (a and b);
    layer3_outputs(4858) <= not (a and b);
    layer3_outputs(4859) <= b and not a;
    layer3_outputs(4860) <= b;
    layer3_outputs(4861) <= not a or b;
    layer3_outputs(4862) <= '0';
    layer3_outputs(4863) <= a or b;
    layer3_outputs(4864) <= a and not b;
    layer3_outputs(4865) <= not a or b;
    layer3_outputs(4866) <= a;
    layer3_outputs(4867) <= not b or a;
    layer3_outputs(4868) <= '0';
    layer3_outputs(4869) <= a and b;
    layer3_outputs(4870) <= not (a and b);
    layer3_outputs(4871) <= a or b;
    layer3_outputs(4872) <= a or b;
    layer3_outputs(4873) <= not a;
    layer3_outputs(4874) <= not b;
    layer3_outputs(4875) <= not b or a;
    layer3_outputs(4876) <= a xor b;
    layer3_outputs(4877) <= '0';
    layer3_outputs(4878) <= a or b;
    layer3_outputs(4879) <= not a or b;
    layer3_outputs(4880) <= not a;
    layer3_outputs(4881) <= not a;
    layer3_outputs(4882) <= not b or a;
    layer3_outputs(4883) <= a and b;
    layer3_outputs(4884) <= not (a xor b);
    layer3_outputs(4885) <= not a or b;
    layer3_outputs(4886) <= not (a or b);
    layer3_outputs(4887) <= '1';
    layer3_outputs(4888) <= a and not b;
    layer3_outputs(4889) <= a;
    layer3_outputs(4890) <= not (a or b);
    layer3_outputs(4891) <= '0';
    layer3_outputs(4892) <= not (a or b);
    layer3_outputs(4893) <= not b;
    layer3_outputs(4894) <= a and b;
    layer3_outputs(4895) <= not a or b;
    layer3_outputs(4896) <= not a or b;
    layer3_outputs(4897) <= b and not a;
    layer3_outputs(4898) <= a and b;
    layer3_outputs(4899) <= a and b;
    layer3_outputs(4900) <= not (a or b);
    layer3_outputs(4901) <= not (a and b);
    layer3_outputs(4902) <= not b or a;
    layer3_outputs(4903) <= not b or a;
    layer3_outputs(4904) <= not a or b;
    layer3_outputs(4905) <= a and not b;
    layer3_outputs(4906) <= not a;
    layer3_outputs(4907) <= not (a or b);
    layer3_outputs(4908) <= a and not b;
    layer3_outputs(4909) <= not b or a;
    layer3_outputs(4910) <= not a;
    layer3_outputs(4911) <= b and not a;
    layer3_outputs(4912) <= not (a or b);
    layer3_outputs(4913) <= a;
    layer3_outputs(4914) <= not a or b;
    layer3_outputs(4915) <= a;
    layer3_outputs(4916) <= not b;
    layer3_outputs(4917) <= b and not a;
    layer3_outputs(4918) <= b;
    layer3_outputs(4919) <= b;
    layer3_outputs(4920) <= not b;
    layer3_outputs(4921) <= not (a xor b);
    layer3_outputs(4922) <= not a or b;
    layer3_outputs(4923) <= not b;
    layer3_outputs(4924) <= b and not a;
    layer3_outputs(4925) <= not a or b;
    layer3_outputs(4926) <= a;
    layer3_outputs(4927) <= not b;
    layer3_outputs(4928) <= '0';
    layer3_outputs(4929) <= not (a and b);
    layer3_outputs(4930) <= '1';
    layer3_outputs(4931) <= '1';
    layer3_outputs(4932) <= not a;
    layer3_outputs(4933) <= not (a or b);
    layer3_outputs(4934) <= a or b;
    layer3_outputs(4935) <= a and not b;
    layer3_outputs(4936) <= b and not a;
    layer3_outputs(4937) <= b and not a;
    layer3_outputs(4938) <= not a or b;
    layer3_outputs(4939) <= '1';
    layer3_outputs(4940) <= not (a or b);
    layer3_outputs(4941) <= a and not b;
    layer3_outputs(4942) <= a xor b;
    layer3_outputs(4943) <= not a or b;
    layer3_outputs(4944) <= not b;
    layer3_outputs(4945) <= not b;
    layer3_outputs(4946) <= b;
    layer3_outputs(4947) <= a or b;
    layer3_outputs(4948) <= not b;
    layer3_outputs(4949) <= '0';
    layer3_outputs(4950) <= not (a or b);
    layer3_outputs(4951) <= a;
    layer3_outputs(4952) <= not b;
    layer3_outputs(4953) <= '1';
    layer3_outputs(4954) <= not (a or b);
    layer3_outputs(4955) <= a and b;
    layer3_outputs(4956) <= a;
    layer3_outputs(4957) <= a and b;
    layer3_outputs(4958) <= b;
    layer3_outputs(4959) <= not a or b;
    layer3_outputs(4960) <= a;
    layer3_outputs(4961) <= a or b;
    layer3_outputs(4962) <= a and not b;
    layer3_outputs(4963) <= a or b;
    layer3_outputs(4964) <= not (a and b);
    layer3_outputs(4965) <= not a or b;
    layer3_outputs(4966) <= not (a and b);
    layer3_outputs(4967) <= b and not a;
    layer3_outputs(4968) <= a and not b;
    layer3_outputs(4969) <= not (a and b);
    layer3_outputs(4970) <= a and b;
    layer3_outputs(4971) <= '0';
    layer3_outputs(4972) <= a xor b;
    layer3_outputs(4973) <= a and b;
    layer3_outputs(4974) <= not (a and b);
    layer3_outputs(4975) <= '1';
    layer3_outputs(4976) <= a and not b;
    layer3_outputs(4977) <= '1';
    layer3_outputs(4978) <= not b or a;
    layer3_outputs(4979) <= '0';
    layer3_outputs(4980) <= '1';
    layer3_outputs(4981) <= not a;
    layer3_outputs(4982) <= not a or b;
    layer3_outputs(4983) <= a and not b;
    layer3_outputs(4984) <= b;
    layer3_outputs(4985) <= not a;
    layer3_outputs(4986) <= '1';
    layer3_outputs(4987) <= not (a or b);
    layer3_outputs(4988) <= a and b;
    layer3_outputs(4989) <= a and b;
    layer3_outputs(4990) <= a xor b;
    layer3_outputs(4991) <= a and not b;
    layer3_outputs(4992) <= not b or a;
    layer3_outputs(4993) <= a or b;
    layer3_outputs(4994) <= not b or a;
    layer3_outputs(4995) <= not b;
    layer3_outputs(4996) <= a and not b;
    layer3_outputs(4997) <= not b or a;
    layer3_outputs(4998) <= not (a and b);
    layer3_outputs(4999) <= a or b;
    layer3_outputs(5000) <= a and b;
    layer3_outputs(5001) <= '0';
    layer3_outputs(5002) <= not b;
    layer3_outputs(5003) <= not (a xor b);
    layer3_outputs(5004) <= '0';
    layer3_outputs(5005) <= not b;
    layer3_outputs(5006) <= a and b;
    layer3_outputs(5007) <= not (a or b);
    layer3_outputs(5008) <= not a or b;
    layer3_outputs(5009) <= not (a and b);
    layer3_outputs(5010) <= b;
    layer3_outputs(5011) <= a and b;
    layer3_outputs(5012) <= '1';
    layer3_outputs(5013) <= a and not b;
    layer3_outputs(5014) <= not a or b;
    layer3_outputs(5015) <= a;
    layer3_outputs(5016) <= not a or b;
    layer3_outputs(5017) <= not b;
    layer3_outputs(5018) <= not a;
    layer3_outputs(5019) <= b;
    layer3_outputs(5020) <= a or b;
    layer3_outputs(5021) <= not a;
    layer3_outputs(5022) <= not a or b;
    layer3_outputs(5023) <= not a or b;
    layer3_outputs(5024) <= '0';
    layer3_outputs(5025) <= not b;
    layer3_outputs(5026) <= not b or a;
    layer3_outputs(5027) <= b and not a;
    layer3_outputs(5028) <= not (a or b);
    layer3_outputs(5029) <= not a;
    layer3_outputs(5030) <= b;
    layer3_outputs(5031) <= '0';
    layer3_outputs(5032) <= a;
    layer3_outputs(5033) <= b;
    layer3_outputs(5034) <= '1';
    layer3_outputs(5035) <= not (a xor b);
    layer3_outputs(5036) <= not (a or b);
    layer3_outputs(5037) <= '0';
    layer3_outputs(5038) <= a or b;
    layer3_outputs(5039) <= '0';
    layer3_outputs(5040) <= a and b;
    layer3_outputs(5041) <= a and not b;
    layer3_outputs(5042) <= a and b;
    layer3_outputs(5043) <= b and not a;
    layer3_outputs(5044) <= a or b;
    layer3_outputs(5045) <= b;
    layer3_outputs(5046) <= not a or b;
    layer3_outputs(5047) <= '0';
    layer3_outputs(5048) <= not a or b;
    layer3_outputs(5049) <= '0';
    layer3_outputs(5050) <= '0';
    layer3_outputs(5051) <= not b or a;
    layer3_outputs(5052) <= not (a or b);
    layer3_outputs(5053) <= not b or a;
    layer3_outputs(5054) <= not b or a;
    layer3_outputs(5055) <= a;
    layer3_outputs(5056) <= a and not b;
    layer3_outputs(5057) <= b and not a;
    layer3_outputs(5058) <= a or b;
    layer3_outputs(5059) <= not b or a;
    layer3_outputs(5060) <= a and b;
    layer3_outputs(5061) <= not a or b;
    layer3_outputs(5062) <= not a;
    layer3_outputs(5063) <= not b;
    layer3_outputs(5064) <= not b;
    layer3_outputs(5065) <= b;
    layer3_outputs(5066) <= '0';
    layer3_outputs(5067) <= not (a or b);
    layer3_outputs(5068) <= b;
    layer3_outputs(5069) <= a and not b;
    layer3_outputs(5070) <= a and not b;
    layer3_outputs(5071) <= not (a xor b);
    layer3_outputs(5072) <= not a or b;
    layer3_outputs(5073) <= not a;
    layer3_outputs(5074) <= not a or b;
    layer3_outputs(5075) <= not (a or b);
    layer3_outputs(5076) <= '1';
    layer3_outputs(5077) <= b;
    layer3_outputs(5078) <= b and not a;
    layer3_outputs(5079) <= '0';
    layer3_outputs(5080) <= b and not a;
    layer3_outputs(5081) <= not a or b;
    layer3_outputs(5082) <= '0';
    layer3_outputs(5083) <= not b or a;
    layer3_outputs(5084) <= not (a and b);
    layer3_outputs(5085) <= '1';
    layer3_outputs(5086) <= a;
    layer3_outputs(5087) <= '0';
    layer3_outputs(5088) <= a;
    layer3_outputs(5089) <= not (a and b);
    layer3_outputs(5090) <= '0';
    layer3_outputs(5091) <= not a or b;
    layer3_outputs(5092) <= b and not a;
    layer3_outputs(5093) <= not (a and b);
    layer3_outputs(5094) <= not a;
    layer3_outputs(5095) <= a;
    layer3_outputs(5096) <= '1';
    layer3_outputs(5097) <= a or b;
    layer3_outputs(5098) <= a or b;
    layer3_outputs(5099) <= b;
    layer3_outputs(5100) <= a and not b;
    layer3_outputs(5101) <= not (a xor b);
    layer3_outputs(5102) <= a and b;
    layer3_outputs(5103) <= not (a or b);
    layer3_outputs(5104) <= b and not a;
    layer3_outputs(5105) <= a or b;
    layer3_outputs(5106) <= a or b;
    layer3_outputs(5107) <= a and not b;
    layer3_outputs(5108) <= not b or a;
    layer3_outputs(5109) <= b and not a;
    layer3_outputs(5110) <= b and not a;
    layer3_outputs(5111) <= not (a or b);
    layer3_outputs(5112) <= b;
    layer3_outputs(5113) <= a;
    layer3_outputs(5114) <= '0';
    layer3_outputs(5115) <= not b or a;
    layer3_outputs(5116) <= b;
    layer3_outputs(5117) <= '0';
    layer3_outputs(5118) <= a and not b;
    layer3_outputs(5119) <= '0';
    layer3_outputs(5120) <= not a or b;
    layer3_outputs(5121) <= a and not b;
    layer3_outputs(5122) <= not b;
    layer3_outputs(5123) <= a and not b;
    layer3_outputs(5124) <= not a;
    layer3_outputs(5125) <= not (a or b);
    layer3_outputs(5126) <= a and b;
    layer3_outputs(5127) <= a;
    layer3_outputs(5128) <= b;
    layer3_outputs(5129) <= a xor b;
    layer3_outputs(5130) <= not (a and b);
    layer3_outputs(5131) <= b and not a;
    layer3_outputs(5132) <= a and b;
    layer3_outputs(5133) <= b;
    layer3_outputs(5134) <= a;
    layer3_outputs(5135) <= not a;
    layer3_outputs(5136) <= b and not a;
    layer3_outputs(5137) <= '0';
    layer3_outputs(5138) <= not b;
    layer3_outputs(5139) <= a and not b;
    layer3_outputs(5140) <= not a;
    layer3_outputs(5141) <= not a or b;
    layer3_outputs(5142) <= a and not b;
    layer3_outputs(5143) <= not b or a;
    layer3_outputs(5144) <= not a;
    layer3_outputs(5145) <= not (a or b);
    layer3_outputs(5146) <= not (a and b);
    layer3_outputs(5147) <= a;
    layer3_outputs(5148) <= not b;
    layer3_outputs(5149) <= '0';
    layer3_outputs(5150) <= not a;
    layer3_outputs(5151) <= a;
    layer3_outputs(5152) <= a and b;
    layer3_outputs(5153) <= a and b;
    layer3_outputs(5154) <= '1';
    layer3_outputs(5155) <= b;
    layer3_outputs(5156) <= a;
    layer3_outputs(5157) <= not (a or b);
    layer3_outputs(5158) <= a or b;
    layer3_outputs(5159) <= '1';
    layer3_outputs(5160) <= not b or a;
    layer3_outputs(5161) <= b;
    layer3_outputs(5162) <= '1';
    layer3_outputs(5163) <= not a or b;
    layer3_outputs(5164) <= not (a or b);
    layer3_outputs(5165) <= a and not b;
    layer3_outputs(5166) <= not (a or b);
    layer3_outputs(5167) <= b and not a;
    layer3_outputs(5168) <= not a or b;
    layer3_outputs(5169) <= not b;
    layer3_outputs(5170) <= '1';
    layer3_outputs(5171) <= a;
    layer3_outputs(5172) <= '0';
    layer3_outputs(5173) <= not b;
    layer3_outputs(5174) <= a and b;
    layer3_outputs(5175) <= '0';
    layer3_outputs(5176) <= not a or b;
    layer3_outputs(5177) <= a or b;
    layer3_outputs(5178) <= not (a or b);
    layer3_outputs(5179) <= not b or a;
    layer3_outputs(5180) <= not (a or b);
    layer3_outputs(5181) <= not b;
    layer3_outputs(5182) <= not (a and b);
    layer3_outputs(5183) <= not (a or b);
    layer3_outputs(5184) <= not a;
    layer3_outputs(5185) <= '1';
    layer3_outputs(5186) <= '0';
    layer3_outputs(5187) <= not b;
    layer3_outputs(5188) <= not a;
    layer3_outputs(5189) <= not b;
    layer3_outputs(5190) <= not (a or b);
    layer3_outputs(5191) <= not (a xor b);
    layer3_outputs(5192) <= '1';
    layer3_outputs(5193) <= a or b;
    layer3_outputs(5194) <= b;
    layer3_outputs(5195) <= a;
    layer3_outputs(5196) <= a;
    layer3_outputs(5197) <= not (a and b);
    layer3_outputs(5198) <= '1';
    layer3_outputs(5199) <= b and not a;
    layer3_outputs(5200) <= b and not a;
    layer3_outputs(5201) <= a and b;
    layer3_outputs(5202) <= not (a and b);
    layer3_outputs(5203) <= '1';
    layer3_outputs(5204) <= a;
    layer3_outputs(5205) <= b and not a;
    layer3_outputs(5206) <= a and b;
    layer3_outputs(5207) <= '1';
    layer3_outputs(5208) <= a and not b;
    layer3_outputs(5209) <= b and not a;
    layer3_outputs(5210) <= not a or b;
    layer3_outputs(5211) <= a and not b;
    layer3_outputs(5212) <= a;
    layer3_outputs(5213) <= a and not b;
    layer3_outputs(5214) <= not a or b;
    layer3_outputs(5215) <= a and not b;
    layer3_outputs(5216) <= a or b;
    layer3_outputs(5217) <= not a;
    layer3_outputs(5218) <= a or b;
    layer3_outputs(5219) <= '0';
    layer3_outputs(5220) <= not b or a;
    layer3_outputs(5221) <= not (a and b);
    layer3_outputs(5222) <= not (a and b);
    layer3_outputs(5223) <= b and not a;
    layer3_outputs(5224) <= '1';
    layer3_outputs(5225) <= a and not b;
    layer3_outputs(5226) <= not a or b;
    layer3_outputs(5227) <= '1';
    layer3_outputs(5228) <= not a or b;
    layer3_outputs(5229) <= a or b;
    layer3_outputs(5230) <= not a;
    layer3_outputs(5231) <= not (a or b);
    layer3_outputs(5232) <= '1';
    layer3_outputs(5233) <= '0';
    layer3_outputs(5234) <= a and b;
    layer3_outputs(5235) <= b;
    layer3_outputs(5236) <= not b or a;
    layer3_outputs(5237) <= '0';
    layer3_outputs(5238) <= a and b;
    layer3_outputs(5239) <= '1';
    layer3_outputs(5240) <= '0';
    layer3_outputs(5241) <= not b;
    layer3_outputs(5242) <= b;
    layer3_outputs(5243) <= not (a and b);
    layer3_outputs(5244) <= a and b;
    layer3_outputs(5245) <= b and not a;
    layer3_outputs(5246) <= a or b;
    layer3_outputs(5247) <= a and b;
    layer3_outputs(5248) <= '0';
    layer3_outputs(5249) <= not (a and b);
    layer3_outputs(5250) <= a and b;
    layer3_outputs(5251) <= not a;
    layer3_outputs(5252) <= '1';
    layer3_outputs(5253) <= not a or b;
    layer3_outputs(5254) <= a and b;
    layer3_outputs(5255) <= a or b;
    layer3_outputs(5256) <= '1';
    layer3_outputs(5257) <= not (a or b);
    layer3_outputs(5258) <= not b;
    layer3_outputs(5259) <= a or b;
    layer3_outputs(5260) <= not a or b;
    layer3_outputs(5261) <= not (a or b);
    layer3_outputs(5262) <= not a;
    layer3_outputs(5263) <= b and not a;
    layer3_outputs(5264) <= not b;
    layer3_outputs(5265) <= '0';
    layer3_outputs(5266) <= '1';
    layer3_outputs(5267) <= b;
    layer3_outputs(5268) <= a or b;
    layer3_outputs(5269) <= not b;
    layer3_outputs(5270) <= a and not b;
    layer3_outputs(5271) <= a or b;
    layer3_outputs(5272) <= b;
    layer3_outputs(5273) <= not (a and b);
    layer3_outputs(5274) <= a;
    layer3_outputs(5275) <= b;
    layer3_outputs(5276) <= b;
    layer3_outputs(5277) <= a;
    layer3_outputs(5278) <= not a or b;
    layer3_outputs(5279) <= a;
    layer3_outputs(5280) <= a;
    layer3_outputs(5281) <= '1';
    layer3_outputs(5282) <= not b or a;
    layer3_outputs(5283) <= b and not a;
    layer3_outputs(5284) <= not (a xor b);
    layer3_outputs(5285) <= a;
    layer3_outputs(5286) <= b;
    layer3_outputs(5287) <= not (a xor b);
    layer3_outputs(5288) <= not (a xor b);
    layer3_outputs(5289) <= not (a or b);
    layer3_outputs(5290) <= a and b;
    layer3_outputs(5291) <= '1';
    layer3_outputs(5292) <= a and b;
    layer3_outputs(5293) <= b;
    layer3_outputs(5294) <= '1';
    layer3_outputs(5295) <= not (a and b);
    layer3_outputs(5296) <= '0';
    layer3_outputs(5297) <= b;
    layer3_outputs(5298) <= a and not b;
    layer3_outputs(5299) <= b;
    layer3_outputs(5300) <= not a or b;
    layer3_outputs(5301) <= a and not b;
    layer3_outputs(5302) <= '0';
    layer3_outputs(5303) <= '0';
    layer3_outputs(5304) <= b;
    layer3_outputs(5305) <= not (a or b);
    layer3_outputs(5306) <= '0';
    layer3_outputs(5307) <= b;
    layer3_outputs(5308) <= a or b;
    layer3_outputs(5309) <= b and not a;
    layer3_outputs(5310) <= a and b;
    layer3_outputs(5311) <= a or b;
    layer3_outputs(5312) <= a;
    layer3_outputs(5313) <= not b;
    layer3_outputs(5314) <= '0';
    layer3_outputs(5315) <= not a;
    layer3_outputs(5316) <= not (a and b);
    layer3_outputs(5317) <= a and b;
    layer3_outputs(5318) <= '0';
    layer3_outputs(5319) <= not b or a;
    layer3_outputs(5320) <= a and b;
    layer3_outputs(5321) <= not a or b;
    layer3_outputs(5322) <= '0';
    layer3_outputs(5323) <= not (a xor b);
    layer3_outputs(5324) <= not (a and b);
    layer3_outputs(5325) <= a and b;
    layer3_outputs(5326) <= '0';
    layer3_outputs(5327) <= '1';
    layer3_outputs(5328) <= '0';
    layer3_outputs(5329) <= b and not a;
    layer3_outputs(5330) <= not (a xor b);
    layer3_outputs(5331) <= not b;
    layer3_outputs(5332) <= a;
    layer3_outputs(5333) <= a and not b;
    layer3_outputs(5334) <= not b or a;
    layer3_outputs(5335) <= not a;
    layer3_outputs(5336) <= b and not a;
    layer3_outputs(5337) <= not (a and b);
    layer3_outputs(5338) <= '1';
    layer3_outputs(5339) <= a or b;
    layer3_outputs(5340) <= a and b;
    layer3_outputs(5341) <= not (a and b);
    layer3_outputs(5342) <= b and not a;
    layer3_outputs(5343) <= '0';
    layer3_outputs(5344) <= not b or a;
    layer3_outputs(5345) <= '0';
    layer3_outputs(5346) <= not a or b;
    layer3_outputs(5347) <= not (a or b);
    layer3_outputs(5348) <= '0';
    layer3_outputs(5349) <= b;
    layer3_outputs(5350) <= not b or a;
    layer3_outputs(5351) <= not (a or b);
    layer3_outputs(5352) <= b and not a;
    layer3_outputs(5353) <= a and b;
    layer3_outputs(5354) <= '1';
    layer3_outputs(5355) <= a and not b;
    layer3_outputs(5356) <= a;
    layer3_outputs(5357) <= not a;
    layer3_outputs(5358) <= b;
    layer3_outputs(5359) <= '0';
    layer3_outputs(5360) <= not a;
    layer3_outputs(5361) <= b;
    layer3_outputs(5362) <= a;
    layer3_outputs(5363) <= not a;
    layer3_outputs(5364) <= not (a or b);
    layer3_outputs(5365) <= not b;
    layer3_outputs(5366) <= a;
    layer3_outputs(5367) <= '1';
    layer3_outputs(5368) <= b and not a;
    layer3_outputs(5369) <= not (a or b);
    layer3_outputs(5370) <= not a;
    layer3_outputs(5371) <= not a or b;
    layer3_outputs(5372) <= '1';
    layer3_outputs(5373) <= a and b;
    layer3_outputs(5374) <= a;
    layer3_outputs(5375) <= b and not a;
    layer3_outputs(5376) <= not (a or b);
    layer3_outputs(5377) <= '1';
    layer3_outputs(5378) <= not a;
    layer3_outputs(5379) <= not b or a;
    layer3_outputs(5380) <= a and not b;
    layer3_outputs(5381) <= a;
    layer3_outputs(5382) <= a or b;
    layer3_outputs(5383) <= not (a xor b);
    layer3_outputs(5384) <= not (a or b);
    layer3_outputs(5385) <= a and not b;
    layer3_outputs(5386) <= b;
    layer3_outputs(5387) <= not b or a;
    layer3_outputs(5388) <= '1';
    layer3_outputs(5389) <= b and not a;
    layer3_outputs(5390) <= a and b;
    layer3_outputs(5391) <= not a or b;
    layer3_outputs(5392) <= a;
    layer3_outputs(5393) <= a and not b;
    layer3_outputs(5394) <= a;
    layer3_outputs(5395) <= a and b;
    layer3_outputs(5396) <= a and not b;
    layer3_outputs(5397) <= a;
    layer3_outputs(5398) <= a and not b;
    layer3_outputs(5399) <= a and not b;
    layer3_outputs(5400) <= b and not a;
    layer3_outputs(5401) <= not (a and b);
    layer3_outputs(5402) <= not b;
    layer3_outputs(5403) <= a and b;
    layer3_outputs(5404) <= a xor b;
    layer3_outputs(5405) <= not b;
    layer3_outputs(5406) <= not (a xor b);
    layer3_outputs(5407) <= a;
    layer3_outputs(5408) <= a and b;
    layer3_outputs(5409) <= a or b;
    layer3_outputs(5410) <= not (a or b);
    layer3_outputs(5411) <= b and not a;
    layer3_outputs(5412) <= a;
    layer3_outputs(5413) <= b and not a;
    layer3_outputs(5414) <= b;
    layer3_outputs(5415) <= a;
    layer3_outputs(5416) <= b and not a;
    layer3_outputs(5417) <= a;
    layer3_outputs(5418) <= a and b;
    layer3_outputs(5419) <= not (a or b);
    layer3_outputs(5420) <= not b or a;
    layer3_outputs(5421) <= a and b;
    layer3_outputs(5422) <= b and not a;
    layer3_outputs(5423) <= b and not a;
    layer3_outputs(5424) <= a and not b;
    layer3_outputs(5425) <= b;
    layer3_outputs(5426) <= b;
    layer3_outputs(5427) <= not a or b;
    layer3_outputs(5428) <= a and b;
    layer3_outputs(5429) <= not (a and b);
    layer3_outputs(5430) <= not a or b;
    layer3_outputs(5431) <= not (a and b);
    layer3_outputs(5432) <= a or b;
    layer3_outputs(5433) <= not a;
    layer3_outputs(5434) <= not b or a;
    layer3_outputs(5435) <= b and not a;
    layer3_outputs(5436) <= '1';
    layer3_outputs(5437) <= not b;
    layer3_outputs(5438) <= not b;
    layer3_outputs(5439) <= a or b;
    layer3_outputs(5440) <= a or b;
    layer3_outputs(5441) <= '1';
    layer3_outputs(5442) <= b;
    layer3_outputs(5443) <= b;
    layer3_outputs(5444) <= not b;
    layer3_outputs(5445) <= a;
    layer3_outputs(5446) <= not (a and b);
    layer3_outputs(5447) <= a and not b;
    layer3_outputs(5448) <= not (a or b);
    layer3_outputs(5449) <= not a or b;
    layer3_outputs(5450) <= not a;
    layer3_outputs(5451) <= a;
    layer3_outputs(5452) <= not b or a;
    layer3_outputs(5453) <= not (a and b);
    layer3_outputs(5454) <= a;
    layer3_outputs(5455) <= a and not b;
    layer3_outputs(5456) <= not (a or b);
    layer3_outputs(5457) <= not (a and b);
    layer3_outputs(5458) <= not a;
    layer3_outputs(5459) <= a;
    layer3_outputs(5460) <= not b or a;
    layer3_outputs(5461) <= a and not b;
    layer3_outputs(5462) <= not b or a;
    layer3_outputs(5463) <= not b or a;
    layer3_outputs(5464) <= b and not a;
    layer3_outputs(5465) <= '0';
    layer3_outputs(5466) <= b and not a;
    layer3_outputs(5467) <= not a or b;
    layer3_outputs(5468) <= not (a and b);
    layer3_outputs(5469) <= a and b;
    layer3_outputs(5470) <= not a or b;
    layer3_outputs(5471) <= '0';
    layer3_outputs(5472) <= b and not a;
    layer3_outputs(5473) <= a xor b;
    layer3_outputs(5474) <= b and not a;
    layer3_outputs(5475) <= b and not a;
    layer3_outputs(5476) <= not b or a;
    layer3_outputs(5477) <= b;
    layer3_outputs(5478) <= '1';
    layer3_outputs(5479) <= '1';
    layer3_outputs(5480) <= not a;
    layer3_outputs(5481) <= a;
    layer3_outputs(5482) <= a xor b;
    layer3_outputs(5483) <= not b or a;
    layer3_outputs(5484) <= a and b;
    layer3_outputs(5485) <= not (a and b);
    layer3_outputs(5486) <= a;
    layer3_outputs(5487) <= not (a or b);
    layer3_outputs(5488) <= a and b;
    layer3_outputs(5489) <= not a;
    layer3_outputs(5490) <= a or b;
    layer3_outputs(5491) <= '0';
    layer3_outputs(5492) <= b and not a;
    layer3_outputs(5493) <= a and not b;
    layer3_outputs(5494) <= not a;
    layer3_outputs(5495) <= a and b;
    layer3_outputs(5496) <= not a or b;
    layer3_outputs(5497) <= '0';
    layer3_outputs(5498) <= '0';
    layer3_outputs(5499) <= '1';
    layer3_outputs(5500) <= b;
    layer3_outputs(5501) <= '0';
    layer3_outputs(5502) <= b;
    layer3_outputs(5503) <= b and not a;
    layer3_outputs(5504) <= b and not a;
    layer3_outputs(5505) <= a and b;
    layer3_outputs(5506) <= '0';
    layer3_outputs(5507) <= not b;
    layer3_outputs(5508) <= not b;
    layer3_outputs(5509) <= b and not a;
    layer3_outputs(5510) <= '1';
    layer3_outputs(5511) <= a and b;
    layer3_outputs(5512) <= not b;
    layer3_outputs(5513) <= a and not b;
    layer3_outputs(5514) <= a or b;
    layer3_outputs(5515) <= b and not a;
    layer3_outputs(5516) <= '0';
    layer3_outputs(5517) <= not (a and b);
    layer3_outputs(5518) <= not b;
    layer3_outputs(5519) <= a and not b;
    layer3_outputs(5520) <= '1';
    layer3_outputs(5521) <= not a or b;
    layer3_outputs(5522) <= not b;
    layer3_outputs(5523) <= a or b;
    layer3_outputs(5524) <= '0';
    layer3_outputs(5525) <= b;
    layer3_outputs(5526) <= a and b;
    layer3_outputs(5527) <= not b;
    layer3_outputs(5528) <= a or b;
    layer3_outputs(5529) <= a and not b;
    layer3_outputs(5530) <= not b;
    layer3_outputs(5531) <= not a;
    layer3_outputs(5532) <= b;
    layer3_outputs(5533) <= a and b;
    layer3_outputs(5534) <= not a or b;
    layer3_outputs(5535) <= not (a and b);
    layer3_outputs(5536) <= not (a and b);
    layer3_outputs(5537) <= not a;
    layer3_outputs(5538) <= b;
    layer3_outputs(5539) <= not a;
    layer3_outputs(5540) <= a or b;
    layer3_outputs(5541) <= not b or a;
    layer3_outputs(5542) <= not b or a;
    layer3_outputs(5543) <= not (a or b);
    layer3_outputs(5544) <= a and not b;
    layer3_outputs(5545) <= not a or b;
    layer3_outputs(5546) <= a;
    layer3_outputs(5547) <= b;
    layer3_outputs(5548) <= not b;
    layer3_outputs(5549) <= '0';
    layer3_outputs(5550) <= b and not a;
    layer3_outputs(5551) <= a or b;
    layer3_outputs(5552) <= b;
    layer3_outputs(5553) <= b;
    layer3_outputs(5554) <= '0';
    layer3_outputs(5555) <= not a or b;
    layer3_outputs(5556) <= '1';
    layer3_outputs(5557) <= a;
    layer3_outputs(5558) <= not (a and b);
    layer3_outputs(5559) <= not a;
    layer3_outputs(5560) <= b;
    layer3_outputs(5561) <= a and b;
    layer3_outputs(5562) <= not b or a;
    layer3_outputs(5563) <= not a or b;
    layer3_outputs(5564) <= '0';
    layer3_outputs(5565) <= '0';
    layer3_outputs(5566) <= '1';
    layer3_outputs(5567) <= not (a or b);
    layer3_outputs(5568) <= not a;
    layer3_outputs(5569) <= b and not a;
    layer3_outputs(5570) <= a xor b;
    layer3_outputs(5571) <= a or b;
    layer3_outputs(5572) <= b and not a;
    layer3_outputs(5573) <= b;
    layer3_outputs(5574) <= not a;
    layer3_outputs(5575) <= a;
    layer3_outputs(5576) <= not a or b;
    layer3_outputs(5577) <= not a or b;
    layer3_outputs(5578) <= not b or a;
    layer3_outputs(5579) <= b;
    layer3_outputs(5580) <= b and not a;
    layer3_outputs(5581) <= a and not b;
    layer3_outputs(5582) <= a and b;
    layer3_outputs(5583) <= not (a or b);
    layer3_outputs(5584) <= '1';
    layer3_outputs(5585) <= not b or a;
    layer3_outputs(5586) <= a and b;
    layer3_outputs(5587) <= '0';
    layer3_outputs(5588) <= a and not b;
    layer3_outputs(5589) <= a and b;
    layer3_outputs(5590) <= not (a and b);
    layer3_outputs(5591) <= not b;
    layer3_outputs(5592) <= b;
    layer3_outputs(5593) <= '1';
    layer3_outputs(5594) <= not a or b;
    layer3_outputs(5595) <= a and not b;
    layer3_outputs(5596) <= not a;
    layer3_outputs(5597) <= a xor b;
    layer3_outputs(5598) <= not b or a;
    layer3_outputs(5599) <= a or b;
    layer3_outputs(5600) <= not (a or b);
    layer3_outputs(5601) <= not b;
    layer3_outputs(5602) <= a and not b;
    layer3_outputs(5603) <= a or b;
    layer3_outputs(5604) <= a;
    layer3_outputs(5605) <= a;
    layer3_outputs(5606) <= not b or a;
    layer3_outputs(5607) <= b and not a;
    layer3_outputs(5608) <= a and not b;
    layer3_outputs(5609) <= not b or a;
    layer3_outputs(5610) <= not a;
    layer3_outputs(5611) <= not (a and b);
    layer3_outputs(5612) <= a xor b;
    layer3_outputs(5613) <= a or b;
    layer3_outputs(5614) <= not b;
    layer3_outputs(5615) <= b and not a;
    layer3_outputs(5616) <= '0';
    layer3_outputs(5617) <= a or b;
    layer3_outputs(5618) <= '1';
    layer3_outputs(5619) <= '0';
    layer3_outputs(5620) <= not (a xor b);
    layer3_outputs(5621) <= not (a or b);
    layer3_outputs(5622) <= not b or a;
    layer3_outputs(5623) <= not b;
    layer3_outputs(5624) <= a and b;
    layer3_outputs(5625) <= not (a and b);
    layer3_outputs(5626) <= '1';
    layer3_outputs(5627) <= not (a or b);
    layer3_outputs(5628) <= a and not b;
    layer3_outputs(5629) <= b;
    layer3_outputs(5630) <= not (a and b);
    layer3_outputs(5631) <= not (a and b);
    layer3_outputs(5632) <= not b;
    layer3_outputs(5633) <= not (a and b);
    layer3_outputs(5634) <= b and not a;
    layer3_outputs(5635) <= not b or a;
    layer3_outputs(5636) <= a and b;
    layer3_outputs(5637) <= '1';
    layer3_outputs(5638) <= b and not a;
    layer3_outputs(5639) <= '1';
    layer3_outputs(5640) <= not (a or b);
    layer3_outputs(5641) <= not b or a;
    layer3_outputs(5642) <= not b;
    layer3_outputs(5643) <= '0';
    layer3_outputs(5644) <= a and b;
    layer3_outputs(5645) <= not b or a;
    layer3_outputs(5646) <= a or b;
    layer3_outputs(5647) <= not a;
    layer3_outputs(5648) <= not (a or b);
    layer3_outputs(5649) <= not a;
    layer3_outputs(5650) <= not b or a;
    layer3_outputs(5651) <= not (a and b);
    layer3_outputs(5652) <= b and not a;
    layer3_outputs(5653) <= a;
    layer3_outputs(5654) <= not (a or b);
    layer3_outputs(5655) <= not b or a;
    layer3_outputs(5656) <= a and b;
    layer3_outputs(5657) <= not a or b;
    layer3_outputs(5658) <= not b or a;
    layer3_outputs(5659) <= not (a and b);
    layer3_outputs(5660) <= b and not a;
    layer3_outputs(5661) <= not a or b;
    layer3_outputs(5662) <= a and not b;
    layer3_outputs(5663) <= a and b;
    layer3_outputs(5664) <= not a or b;
    layer3_outputs(5665) <= not (a or b);
    layer3_outputs(5666) <= not b or a;
    layer3_outputs(5667) <= not (a xor b);
    layer3_outputs(5668) <= a or b;
    layer3_outputs(5669) <= a and b;
    layer3_outputs(5670) <= a and not b;
    layer3_outputs(5671) <= '0';
    layer3_outputs(5672) <= '0';
    layer3_outputs(5673) <= a and not b;
    layer3_outputs(5674) <= not (a or b);
    layer3_outputs(5675) <= not b;
    layer3_outputs(5676) <= b;
    layer3_outputs(5677) <= a and not b;
    layer3_outputs(5678) <= b;
    layer3_outputs(5679) <= '0';
    layer3_outputs(5680) <= not (a or b);
    layer3_outputs(5681) <= not b or a;
    layer3_outputs(5682) <= not (a or b);
    layer3_outputs(5683) <= a and not b;
    layer3_outputs(5684) <= a;
    layer3_outputs(5685) <= a xor b;
    layer3_outputs(5686) <= '0';
    layer3_outputs(5687) <= not b or a;
    layer3_outputs(5688) <= a and b;
    layer3_outputs(5689) <= a and b;
    layer3_outputs(5690) <= a and not b;
    layer3_outputs(5691) <= not (a or b);
    layer3_outputs(5692) <= '1';
    layer3_outputs(5693) <= '1';
    layer3_outputs(5694) <= a xor b;
    layer3_outputs(5695) <= not b or a;
    layer3_outputs(5696) <= not b or a;
    layer3_outputs(5697) <= a or b;
    layer3_outputs(5698) <= not b or a;
    layer3_outputs(5699) <= a;
    layer3_outputs(5700) <= '0';
    layer3_outputs(5701) <= not a;
    layer3_outputs(5702) <= a xor b;
    layer3_outputs(5703) <= not (a xor b);
    layer3_outputs(5704) <= not b;
    layer3_outputs(5705) <= b and not a;
    layer3_outputs(5706) <= '1';
    layer3_outputs(5707) <= not (a or b);
    layer3_outputs(5708) <= not b;
    layer3_outputs(5709) <= not a or b;
    layer3_outputs(5710) <= a and not b;
    layer3_outputs(5711) <= '1';
    layer3_outputs(5712) <= not b or a;
    layer3_outputs(5713) <= b and not a;
    layer3_outputs(5714) <= not b;
    layer3_outputs(5715) <= not (a xor b);
    layer3_outputs(5716) <= b;
    layer3_outputs(5717) <= not b or a;
    layer3_outputs(5718) <= not a;
    layer3_outputs(5719) <= a or b;
    layer3_outputs(5720) <= a and b;
    layer3_outputs(5721) <= a and b;
    layer3_outputs(5722) <= a and b;
    layer3_outputs(5723) <= a;
    layer3_outputs(5724) <= a or b;
    layer3_outputs(5725) <= not (a or b);
    layer3_outputs(5726) <= not a or b;
    layer3_outputs(5727) <= not (a and b);
    layer3_outputs(5728) <= not b;
    layer3_outputs(5729) <= not (a and b);
    layer3_outputs(5730) <= b and not a;
    layer3_outputs(5731) <= a and not b;
    layer3_outputs(5732) <= not (a xor b);
    layer3_outputs(5733) <= not a;
    layer3_outputs(5734) <= b and not a;
    layer3_outputs(5735) <= b and not a;
    layer3_outputs(5736) <= a;
    layer3_outputs(5737) <= not (a or b);
    layer3_outputs(5738) <= b and not a;
    layer3_outputs(5739) <= not a;
    layer3_outputs(5740) <= not (a and b);
    layer3_outputs(5741) <= not a or b;
    layer3_outputs(5742) <= b and not a;
    layer3_outputs(5743) <= not (a and b);
    layer3_outputs(5744) <= b and not a;
    layer3_outputs(5745) <= not b;
    layer3_outputs(5746) <= not (a xor b);
    layer3_outputs(5747) <= a and b;
    layer3_outputs(5748) <= not a or b;
    layer3_outputs(5749) <= '1';
    layer3_outputs(5750) <= '0';
    layer3_outputs(5751) <= not (a and b);
    layer3_outputs(5752) <= b and not a;
    layer3_outputs(5753) <= '0';
    layer3_outputs(5754) <= not b;
    layer3_outputs(5755) <= '1';
    layer3_outputs(5756) <= a;
    layer3_outputs(5757) <= not b or a;
    layer3_outputs(5758) <= not a;
    layer3_outputs(5759) <= not (a and b);
    layer3_outputs(5760) <= not b or a;
    layer3_outputs(5761) <= not b;
    layer3_outputs(5762) <= a and b;
    layer3_outputs(5763) <= '1';
    layer3_outputs(5764) <= not a;
    layer3_outputs(5765) <= '1';
    layer3_outputs(5766) <= a;
    layer3_outputs(5767) <= not (a and b);
    layer3_outputs(5768) <= a and not b;
    layer3_outputs(5769) <= not a;
    layer3_outputs(5770) <= a xor b;
    layer3_outputs(5771) <= not b or a;
    layer3_outputs(5772) <= not a;
    layer3_outputs(5773) <= a and not b;
    layer3_outputs(5774) <= a and b;
    layer3_outputs(5775) <= not a or b;
    layer3_outputs(5776) <= a or b;
    layer3_outputs(5777) <= a or b;
    layer3_outputs(5778) <= a and b;
    layer3_outputs(5779) <= b and not a;
    layer3_outputs(5780) <= a and not b;
    layer3_outputs(5781) <= '0';
    layer3_outputs(5782) <= not (a or b);
    layer3_outputs(5783) <= a and not b;
    layer3_outputs(5784) <= not (a xor b);
    layer3_outputs(5785) <= not a or b;
    layer3_outputs(5786) <= b and not a;
    layer3_outputs(5787) <= not b or a;
    layer3_outputs(5788) <= a or b;
    layer3_outputs(5789) <= not (a xor b);
    layer3_outputs(5790) <= not (a and b);
    layer3_outputs(5791) <= not (a and b);
    layer3_outputs(5792) <= '0';
    layer3_outputs(5793) <= not b;
    layer3_outputs(5794) <= not b or a;
    layer3_outputs(5795) <= a and not b;
    layer3_outputs(5796) <= '0';
    layer3_outputs(5797) <= a;
    layer3_outputs(5798) <= not a or b;
    layer3_outputs(5799) <= '1';
    layer3_outputs(5800) <= b;
    layer3_outputs(5801) <= b;
    layer3_outputs(5802) <= not a or b;
    layer3_outputs(5803) <= a and not b;
    layer3_outputs(5804) <= not a;
    layer3_outputs(5805) <= b;
    layer3_outputs(5806) <= a and b;
    layer3_outputs(5807) <= b and not a;
    layer3_outputs(5808) <= a;
    layer3_outputs(5809) <= not a or b;
    layer3_outputs(5810) <= a and not b;
    layer3_outputs(5811) <= not (a and b);
    layer3_outputs(5812) <= a or b;
    layer3_outputs(5813) <= a;
    layer3_outputs(5814) <= not (a or b);
    layer3_outputs(5815) <= a and b;
    layer3_outputs(5816) <= '0';
    layer3_outputs(5817) <= b;
    layer3_outputs(5818) <= not a;
    layer3_outputs(5819) <= not b or a;
    layer3_outputs(5820) <= not a or b;
    layer3_outputs(5821) <= not (a and b);
    layer3_outputs(5822) <= '0';
    layer3_outputs(5823) <= not (a or b);
    layer3_outputs(5824) <= b and not a;
    layer3_outputs(5825) <= a or b;
    layer3_outputs(5826) <= not b;
    layer3_outputs(5827) <= not b;
    layer3_outputs(5828) <= a;
    layer3_outputs(5829) <= a;
    layer3_outputs(5830) <= a and b;
    layer3_outputs(5831) <= not b or a;
    layer3_outputs(5832) <= b;
    layer3_outputs(5833) <= a and not b;
    layer3_outputs(5834) <= '0';
    layer3_outputs(5835) <= a and not b;
    layer3_outputs(5836) <= not a;
    layer3_outputs(5837) <= '1';
    layer3_outputs(5838) <= a or b;
    layer3_outputs(5839) <= a;
    layer3_outputs(5840) <= '0';
    layer3_outputs(5841) <= not (a and b);
    layer3_outputs(5842) <= '0';
    layer3_outputs(5843) <= not a;
    layer3_outputs(5844) <= not a;
    layer3_outputs(5845) <= not b or a;
    layer3_outputs(5846) <= not (a or b);
    layer3_outputs(5847) <= not b or a;
    layer3_outputs(5848) <= not b or a;
    layer3_outputs(5849) <= b;
    layer3_outputs(5850) <= not b;
    layer3_outputs(5851) <= not (a or b);
    layer3_outputs(5852) <= not (a and b);
    layer3_outputs(5853) <= not (a xor b);
    layer3_outputs(5854) <= a and not b;
    layer3_outputs(5855) <= a or b;
    layer3_outputs(5856) <= b;
    layer3_outputs(5857) <= not b or a;
    layer3_outputs(5858) <= not a or b;
    layer3_outputs(5859) <= not a or b;
    layer3_outputs(5860) <= b and not a;
    layer3_outputs(5861) <= '1';
    layer3_outputs(5862) <= a and not b;
    layer3_outputs(5863) <= '0';
    layer3_outputs(5864) <= not b;
    layer3_outputs(5865) <= not (a or b);
    layer3_outputs(5866) <= not b;
    layer3_outputs(5867) <= a xor b;
    layer3_outputs(5868) <= a and b;
    layer3_outputs(5869) <= a or b;
    layer3_outputs(5870) <= a and b;
    layer3_outputs(5871) <= not a or b;
    layer3_outputs(5872) <= not b;
    layer3_outputs(5873) <= '0';
    layer3_outputs(5874) <= b and not a;
    layer3_outputs(5875) <= a and b;
    layer3_outputs(5876) <= not (a xor b);
    layer3_outputs(5877) <= not a;
    layer3_outputs(5878) <= a and not b;
    layer3_outputs(5879) <= not b;
    layer3_outputs(5880) <= b;
    layer3_outputs(5881) <= not (a or b);
    layer3_outputs(5882) <= a;
    layer3_outputs(5883) <= b;
    layer3_outputs(5884) <= not b;
    layer3_outputs(5885) <= b and not a;
    layer3_outputs(5886) <= not (a and b);
    layer3_outputs(5887) <= not (a or b);
    layer3_outputs(5888) <= b and not a;
    layer3_outputs(5889) <= a and not b;
    layer3_outputs(5890) <= a;
    layer3_outputs(5891) <= not (a or b);
    layer3_outputs(5892) <= a;
    layer3_outputs(5893) <= not a or b;
    layer3_outputs(5894) <= a or b;
    layer3_outputs(5895) <= a and b;
    layer3_outputs(5896) <= b;
    layer3_outputs(5897) <= not b or a;
    layer3_outputs(5898) <= not (a and b);
    layer3_outputs(5899) <= '0';
    layer3_outputs(5900) <= a and not b;
    layer3_outputs(5901) <= b;
    layer3_outputs(5902) <= b;
    layer3_outputs(5903) <= not (a or b);
    layer3_outputs(5904) <= b;
    layer3_outputs(5905) <= a and not b;
    layer3_outputs(5906) <= a or b;
    layer3_outputs(5907) <= b;
    layer3_outputs(5908) <= not a or b;
    layer3_outputs(5909) <= not (a or b);
    layer3_outputs(5910) <= a xor b;
    layer3_outputs(5911) <= b and not a;
    layer3_outputs(5912) <= a and not b;
    layer3_outputs(5913) <= a and b;
    layer3_outputs(5914) <= b;
    layer3_outputs(5915) <= a and not b;
    layer3_outputs(5916) <= not b;
    layer3_outputs(5917) <= '1';
    layer3_outputs(5918) <= not b;
    layer3_outputs(5919) <= '1';
    layer3_outputs(5920) <= not a or b;
    layer3_outputs(5921) <= not b;
    layer3_outputs(5922) <= not (a and b);
    layer3_outputs(5923) <= b and not a;
    layer3_outputs(5924) <= '1';
    layer3_outputs(5925) <= a and not b;
    layer3_outputs(5926) <= b;
    layer3_outputs(5927) <= not a;
    layer3_outputs(5928) <= '0';
    layer3_outputs(5929) <= b and not a;
    layer3_outputs(5930) <= not (a xor b);
    layer3_outputs(5931) <= not (a xor b);
    layer3_outputs(5932) <= not a;
    layer3_outputs(5933) <= a;
    layer3_outputs(5934) <= b;
    layer3_outputs(5935) <= not (a or b);
    layer3_outputs(5936) <= not b;
    layer3_outputs(5937) <= b;
    layer3_outputs(5938) <= b and not a;
    layer3_outputs(5939) <= a and not b;
    layer3_outputs(5940) <= a and not b;
    layer3_outputs(5941) <= not (a xor b);
    layer3_outputs(5942) <= not b;
    layer3_outputs(5943) <= not b or a;
    layer3_outputs(5944) <= b;
    layer3_outputs(5945) <= not (a and b);
    layer3_outputs(5946) <= not (a or b);
    layer3_outputs(5947) <= not a or b;
    layer3_outputs(5948) <= a or b;
    layer3_outputs(5949) <= not a or b;
    layer3_outputs(5950) <= not b;
    layer3_outputs(5951) <= not a;
    layer3_outputs(5952) <= a and not b;
    layer3_outputs(5953) <= a and b;
    layer3_outputs(5954) <= a or b;
    layer3_outputs(5955) <= not (a xor b);
    layer3_outputs(5956) <= '1';
    layer3_outputs(5957) <= a and not b;
    layer3_outputs(5958) <= not b;
    layer3_outputs(5959) <= a;
    layer3_outputs(5960) <= '1';
    layer3_outputs(5961) <= not a or b;
    layer3_outputs(5962) <= '1';
    layer3_outputs(5963) <= b and not a;
    layer3_outputs(5964) <= not (a or b);
    layer3_outputs(5965) <= a and not b;
    layer3_outputs(5966) <= a and not b;
    layer3_outputs(5967) <= not (a xor b);
    layer3_outputs(5968) <= a and b;
    layer3_outputs(5969) <= a or b;
    layer3_outputs(5970) <= a and not b;
    layer3_outputs(5971) <= not (a xor b);
    layer3_outputs(5972) <= '1';
    layer3_outputs(5973) <= not b or a;
    layer3_outputs(5974) <= not b;
    layer3_outputs(5975) <= a and b;
    layer3_outputs(5976) <= not a or b;
    layer3_outputs(5977) <= not (a and b);
    layer3_outputs(5978) <= not b;
    layer3_outputs(5979) <= a;
    layer3_outputs(5980) <= b;
    layer3_outputs(5981) <= a;
    layer3_outputs(5982) <= not a or b;
    layer3_outputs(5983) <= not (a or b);
    layer3_outputs(5984) <= a;
    layer3_outputs(5985) <= a or b;
    layer3_outputs(5986) <= not (a and b);
    layer3_outputs(5987) <= '1';
    layer3_outputs(5988) <= not (a xor b);
    layer3_outputs(5989) <= not (a and b);
    layer3_outputs(5990) <= b;
    layer3_outputs(5991) <= not b;
    layer3_outputs(5992) <= not a or b;
    layer3_outputs(5993) <= not (a and b);
    layer3_outputs(5994) <= a or b;
    layer3_outputs(5995) <= not b or a;
    layer3_outputs(5996) <= not a or b;
    layer3_outputs(5997) <= b and not a;
    layer3_outputs(5998) <= not a;
    layer3_outputs(5999) <= not a;
    layer3_outputs(6000) <= not (a and b);
    layer3_outputs(6001) <= not (a and b);
    layer3_outputs(6002) <= not b;
    layer3_outputs(6003) <= not a;
    layer3_outputs(6004) <= '0';
    layer3_outputs(6005) <= b;
    layer3_outputs(6006) <= a and not b;
    layer3_outputs(6007) <= b and not a;
    layer3_outputs(6008) <= not a or b;
    layer3_outputs(6009) <= not a;
    layer3_outputs(6010) <= not b or a;
    layer3_outputs(6011) <= not a or b;
    layer3_outputs(6012) <= '0';
    layer3_outputs(6013) <= a and b;
    layer3_outputs(6014) <= '1';
    layer3_outputs(6015) <= a or b;
    layer3_outputs(6016) <= '1';
    layer3_outputs(6017) <= not b;
    layer3_outputs(6018) <= a and not b;
    layer3_outputs(6019) <= not (a or b);
    layer3_outputs(6020) <= not (a or b);
    layer3_outputs(6021) <= not b or a;
    layer3_outputs(6022) <= a;
    layer3_outputs(6023) <= not (a and b);
    layer3_outputs(6024) <= a or b;
    layer3_outputs(6025) <= not (a and b);
    layer3_outputs(6026) <= '0';
    layer3_outputs(6027) <= a or b;
    layer3_outputs(6028) <= a and b;
    layer3_outputs(6029) <= a;
    layer3_outputs(6030) <= not (a xor b);
    layer3_outputs(6031) <= not a;
    layer3_outputs(6032) <= not (a or b);
    layer3_outputs(6033) <= b and not a;
    layer3_outputs(6034) <= a;
    layer3_outputs(6035) <= not b;
    layer3_outputs(6036) <= not a;
    layer3_outputs(6037) <= a and b;
    layer3_outputs(6038) <= a and not b;
    layer3_outputs(6039) <= a xor b;
    layer3_outputs(6040) <= b and not a;
    layer3_outputs(6041) <= not (a xor b);
    layer3_outputs(6042) <= '1';
    layer3_outputs(6043) <= a xor b;
    layer3_outputs(6044) <= not a or b;
    layer3_outputs(6045) <= not b or a;
    layer3_outputs(6046) <= b;
    layer3_outputs(6047) <= not b or a;
    layer3_outputs(6048) <= not (a and b);
    layer3_outputs(6049) <= not (a and b);
    layer3_outputs(6050) <= not (a or b);
    layer3_outputs(6051) <= b and not a;
    layer3_outputs(6052) <= a or b;
    layer3_outputs(6053) <= not (a or b);
    layer3_outputs(6054) <= not (a or b);
    layer3_outputs(6055) <= not a;
    layer3_outputs(6056) <= b;
    layer3_outputs(6057) <= '0';
    layer3_outputs(6058) <= not (a or b);
    layer3_outputs(6059) <= not b;
    layer3_outputs(6060) <= not a or b;
    layer3_outputs(6061) <= not b or a;
    layer3_outputs(6062) <= b;
    layer3_outputs(6063) <= not (a or b);
    layer3_outputs(6064) <= not (a and b);
    layer3_outputs(6065) <= not a;
    layer3_outputs(6066) <= not b or a;
    layer3_outputs(6067) <= a and not b;
    layer3_outputs(6068) <= '1';
    layer3_outputs(6069) <= a or b;
    layer3_outputs(6070) <= '1';
    layer3_outputs(6071) <= a;
    layer3_outputs(6072) <= a;
    layer3_outputs(6073) <= not (a and b);
    layer3_outputs(6074) <= not (a or b);
    layer3_outputs(6075) <= b and not a;
    layer3_outputs(6076) <= not a or b;
    layer3_outputs(6077) <= a and b;
    layer3_outputs(6078) <= not b;
    layer3_outputs(6079) <= not (a or b);
    layer3_outputs(6080) <= not (a and b);
    layer3_outputs(6081) <= a and b;
    layer3_outputs(6082) <= b and not a;
    layer3_outputs(6083) <= a or b;
    layer3_outputs(6084) <= '1';
    layer3_outputs(6085) <= not (a and b);
    layer3_outputs(6086) <= a and not b;
    layer3_outputs(6087) <= not (a and b);
    layer3_outputs(6088) <= a;
    layer3_outputs(6089) <= not a;
    layer3_outputs(6090) <= a and b;
    layer3_outputs(6091) <= b;
    layer3_outputs(6092) <= not b;
    layer3_outputs(6093) <= not (a and b);
    layer3_outputs(6094) <= not a;
    layer3_outputs(6095) <= a and not b;
    layer3_outputs(6096) <= not (a or b);
    layer3_outputs(6097) <= not a or b;
    layer3_outputs(6098) <= b and not a;
    layer3_outputs(6099) <= '0';
    layer3_outputs(6100) <= '1';
    layer3_outputs(6101) <= not a;
    layer3_outputs(6102) <= a or b;
    layer3_outputs(6103) <= a;
    layer3_outputs(6104) <= '1';
    layer3_outputs(6105) <= a and not b;
    layer3_outputs(6106) <= not (a or b);
    layer3_outputs(6107) <= b;
    layer3_outputs(6108) <= not b or a;
    layer3_outputs(6109) <= '0';
    layer3_outputs(6110) <= not b;
    layer3_outputs(6111) <= a and not b;
    layer3_outputs(6112) <= a xor b;
    layer3_outputs(6113) <= not (a and b);
    layer3_outputs(6114) <= not b or a;
    layer3_outputs(6115) <= '1';
    layer3_outputs(6116) <= not (a or b);
    layer3_outputs(6117) <= not a or b;
    layer3_outputs(6118) <= b;
    layer3_outputs(6119) <= a;
    layer3_outputs(6120) <= b and not a;
    layer3_outputs(6121) <= b and not a;
    layer3_outputs(6122) <= b and not a;
    layer3_outputs(6123) <= not b;
    layer3_outputs(6124) <= a and not b;
    layer3_outputs(6125) <= '1';
    layer3_outputs(6126) <= '0';
    layer3_outputs(6127) <= a and b;
    layer3_outputs(6128) <= not (a and b);
    layer3_outputs(6129) <= '1';
    layer3_outputs(6130) <= '0';
    layer3_outputs(6131) <= '0';
    layer3_outputs(6132) <= b;
    layer3_outputs(6133) <= a;
    layer3_outputs(6134) <= not (a xor b);
    layer3_outputs(6135) <= not b or a;
    layer3_outputs(6136) <= a or b;
    layer3_outputs(6137) <= b and not a;
    layer3_outputs(6138) <= '0';
    layer3_outputs(6139) <= a xor b;
    layer3_outputs(6140) <= b and not a;
    layer3_outputs(6141) <= a and not b;
    layer3_outputs(6142) <= a or b;
    layer3_outputs(6143) <= '0';
    layer3_outputs(6144) <= not (a or b);
    layer3_outputs(6145) <= a or b;
    layer3_outputs(6146) <= not a or b;
    layer3_outputs(6147) <= not (a or b);
    layer3_outputs(6148) <= not a or b;
    layer3_outputs(6149) <= not b;
    layer3_outputs(6150) <= a and not b;
    layer3_outputs(6151) <= a and b;
    layer3_outputs(6152) <= b;
    layer3_outputs(6153) <= not a or b;
    layer3_outputs(6154) <= a and b;
    layer3_outputs(6155) <= b and not a;
    layer3_outputs(6156) <= b and not a;
    layer3_outputs(6157) <= a and b;
    layer3_outputs(6158) <= b and not a;
    layer3_outputs(6159) <= not a;
    layer3_outputs(6160) <= '1';
    layer3_outputs(6161) <= a and b;
    layer3_outputs(6162) <= a and not b;
    layer3_outputs(6163) <= '1';
    layer3_outputs(6164) <= a or b;
    layer3_outputs(6165) <= a and b;
    layer3_outputs(6166) <= not b;
    layer3_outputs(6167) <= not b;
    layer3_outputs(6168) <= a and not b;
    layer3_outputs(6169) <= a xor b;
    layer3_outputs(6170) <= not a;
    layer3_outputs(6171) <= a or b;
    layer3_outputs(6172) <= b;
    layer3_outputs(6173) <= not b or a;
    layer3_outputs(6174) <= not (a and b);
    layer3_outputs(6175) <= a;
    layer3_outputs(6176) <= a or b;
    layer3_outputs(6177) <= '0';
    layer3_outputs(6178) <= a or b;
    layer3_outputs(6179) <= not b;
    layer3_outputs(6180) <= a and not b;
    layer3_outputs(6181) <= not (a or b);
    layer3_outputs(6182) <= a and b;
    layer3_outputs(6183) <= not (a and b);
    layer3_outputs(6184) <= a and b;
    layer3_outputs(6185) <= not a;
    layer3_outputs(6186) <= b;
    layer3_outputs(6187) <= a and not b;
    layer3_outputs(6188) <= a or b;
    layer3_outputs(6189) <= b and not a;
    layer3_outputs(6190) <= not a or b;
    layer3_outputs(6191) <= a;
    layer3_outputs(6192) <= '0';
    layer3_outputs(6193) <= not a;
    layer3_outputs(6194) <= '0';
    layer3_outputs(6195) <= not (a or b);
    layer3_outputs(6196) <= a and not b;
    layer3_outputs(6197) <= not a or b;
    layer3_outputs(6198) <= a;
    layer3_outputs(6199) <= a and not b;
    layer3_outputs(6200) <= '1';
    layer3_outputs(6201) <= a xor b;
    layer3_outputs(6202) <= a and not b;
    layer3_outputs(6203) <= b;
    layer3_outputs(6204) <= '1';
    layer3_outputs(6205) <= a or b;
    layer3_outputs(6206) <= a or b;
    layer3_outputs(6207) <= a;
    layer3_outputs(6208) <= not b;
    layer3_outputs(6209) <= not b or a;
    layer3_outputs(6210) <= a;
    layer3_outputs(6211) <= not (a xor b);
    layer3_outputs(6212) <= a;
    layer3_outputs(6213) <= a and not b;
    layer3_outputs(6214) <= b and not a;
    layer3_outputs(6215) <= not a;
    layer3_outputs(6216) <= a or b;
    layer3_outputs(6217) <= '1';
    layer3_outputs(6218) <= b;
    layer3_outputs(6219) <= not b or a;
    layer3_outputs(6220) <= b and not a;
    layer3_outputs(6221) <= not (a or b);
    layer3_outputs(6222) <= not (a xor b);
    layer3_outputs(6223) <= '1';
    layer3_outputs(6224) <= b and not a;
    layer3_outputs(6225) <= not (a xor b);
    layer3_outputs(6226) <= not a;
    layer3_outputs(6227) <= '1';
    layer3_outputs(6228) <= not a;
    layer3_outputs(6229) <= b and not a;
    layer3_outputs(6230) <= a and b;
    layer3_outputs(6231) <= not b;
    layer3_outputs(6232) <= not (a and b);
    layer3_outputs(6233) <= a or b;
    layer3_outputs(6234) <= a and not b;
    layer3_outputs(6235) <= a or b;
    layer3_outputs(6236) <= not b or a;
    layer3_outputs(6237) <= a or b;
    layer3_outputs(6238) <= not b;
    layer3_outputs(6239) <= not (a xor b);
    layer3_outputs(6240) <= a or b;
    layer3_outputs(6241) <= not (a xor b);
    layer3_outputs(6242) <= a or b;
    layer3_outputs(6243) <= not (a xor b);
    layer3_outputs(6244) <= b;
    layer3_outputs(6245) <= b and not a;
    layer3_outputs(6246) <= not b or a;
    layer3_outputs(6247) <= a or b;
    layer3_outputs(6248) <= a;
    layer3_outputs(6249) <= not a;
    layer3_outputs(6250) <= not b;
    layer3_outputs(6251) <= '1';
    layer3_outputs(6252) <= not a;
    layer3_outputs(6253) <= b;
    layer3_outputs(6254) <= not b or a;
    layer3_outputs(6255) <= '0';
    layer3_outputs(6256) <= b;
    layer3_outputs(6257) <= a;
    layer3_outputs(6258) <= not b or a;
    layer3_outputs(6259) <= a;
    layer3_outputs(6260) <= a or b;
    layer3_outputs(6261) <= b;
    layer3_outputs(6262) <= a xor b;
    layer3_outputs(6263) <= b and not a;
    layer3_outputs(6264) <= not a;
    layer3_outputs(6265) <= not b;
    layer3_outputs(6266) <= not a or b;
    layer3_outputs(6267) <= not (a or b);
    layer3_outputs(6268) <= a or b;
    layer3_outputs(6269) <= not (a or b);
    layer3_outputs(6270) <= a or b;
    layer3_outputs(6271) <= a and not b;
    layer3_outputs(6272) <= not a;
    layer3_outputs(6273) <= not a;
    layer3_outputs(6274) <= not b;
    layer3_outputs(6275) <= a and not b;
    layer3_outputs(6276) <= not (a or b);
    layer3_outputs(6277) <= not a or b;
    layer3_outputs(6278) <= not b or a;
    layer3_outputs(6279) <= not b or a;
    layer3_outputs(6280) <= a and not b;
    layer3_outputs(6281) <= a and not b;
    layer3_outputs(6282) <= b;
    layer3_outputs(6283) <= a and b;
    layer3_outputs(6284) <= not a or b;
    layer3_outputs(6285) <= a;
    layer3_outputs(6286) <= not (a and b);
    layer3_outputs(6287) <= b and not a;
    layer3_outputs(6288) <= a or b;
    layer3_outputs(6289) <= not b or a;
    layer3_outputs(6290) <= b and not a;
    layer3_outputs(6291) <= not (a and b);
    layer3_outputs(6292) <= a and not b;
    layer3_outputs(6293) <= '0';
    layer3_outputs(6294) <= a;
    layer3_outputs(6295) <= a and b;
    layer3_outputs(6296) <= not a;
    layer3_outputs(6297) <= not a;
    layer3_outputs(6298) <= a;
    layer3_outputs(6299) <= not b;
    layer3_outputs(6300) <= not b;
    layer3_outputs(6301) <= not (a and b);
    layer3_outputs(6302) <= not b or a;
    layer3_outputs(6303) <= a and not b;
    layer3_outputs(6304) <= a xor b;
    layer3_outputs(6305) <= a and not b;
    layer3_outputs(6306) <= a and b;
    layer3_outputs(6307) <= a;
    layer3_outputs(6308) <= not (a or b);
    layer3_outputs(6309) <= b;
    layer3_outputs(6310) <= b;
    layer3_outputs(6311) <= a and not b;
    layer3_outputs(6312) <= b;
    layer3_outputs(6313) <= b;
    layer3_outputs(6314) <= a and not b;
    layer3_outputs(6315) <= '1';
    layer3_outputs(6316) <= b and not a;
    layer3_outputs(6317) <= '0';
    layer3_outputs(6318) <= a;
    layer3_outputs(6319) <= b and not a;
    layer3_outputs(6320) <= not (a and b);
    layer3_outputs(6321) <= not (a or b);
    layer3_outputs(6322) <= b;
    layer3_outputs(6323) <= not (a or b);
    layer3_outputs(6324) <= '1';
    layer3_outputs(6325) <= a;
    layer3_outputs(6326) <= not a or b;
    layer3_outputs(6327) <= '1';
    layer3_outputs(6328) <= a xor b;
    layer3_outputs(6329) <= a and not b;
    layer3_outputs(6330) <= not a or b;
    layer3_outputs(6331) <= a or b;
    layer3_outputs(6332) <= a and b;
    layer3_outputs(6333) <= not a or b;
    layer3_outputs(6334) <= not (a or b);
    layer3_outputs(6335) <= not b or a;
    layer3_outputs(6336) <= a or b;
    layer3_outputs(6337) <= not a;
    layer3_outputs(6338) <= a;
    layer3_outputs(6339) <= not b or a;
    layer3_outputs(6340) <= '0';
    layer3_outputs(6341) <= '0';
    layer3_outputs(6342) <= a or b;
    layer3_outputs(6343) <= not b or a;
    layer3_outputs(6344) <= b;
    layer3_outputs(6345) <= '1';
    layer3_outputs(6346) <= b and not a;
    layer3_outputs(6347) <= a and not b;
    layer3_outputs(6348) <= a and not b;
    layer3_outputs(6349) <= a and not b;
    layer3_outputs(6350) <= '1';
    layer3_outputs(6351) <= not a or b;
    layer3_outputs(6352) <= not b or a;
    layer3_outputs(6353) <= a xor b;
    layer3_outputs(6354) <= a;
    layer3_outputs(6355) <= a;
    layer3_outputs(6356) <= b;
    layer3_outputs(6357) <= a;
    layer3_outputs(6358) <= a;
    layer3_outputs(6359) <= not b;
    layer3_outputs(6360) <= b and not a;
    layer3_outputs(6361) <= not b;
    layer3_outputs(6362) <= not b or a;
    layer3_outputs(6363) <= not a;
    layer3_outputs(6364) <= a and b;
    layer3_outputs(6365) <= not a or b;
    layer3_outputs(6366) <= b and not a;
    layer3_outputs(6367) <= '1';
    layer3_outputs(6368) <= not a or b;
    layer3_outputs(6369) <= not b or a;
    layer3_outputs(6370) <= b and not a;
    layer3_outputs(6371) <= a or b;
    layer3_outputs(6372) <= a and b;
    layer3_outputs(6373) <= a or b;
    layer3_outputs(6374) <= '0';
    layer3_outputs(6375) <= not b or a;
    layer3_outputs(6376) <= a or b;
    layer3_outputs(6377) <= '0';
    layer3_outputs(6378) <= a;
    layer3_outputs(6379) <= a or b;
    layer3_outputs(6380) <= a;
    layer3_outputs(6381) <= a or b;
    layer3_outputs(6382) <= b and not a;
    layer3_outputs(6383) <= '1';
    layer3_outputs(6384) <= not (a or b);
    layer3_outputs(6385) <= not b or a;
    layer3_outputs(6386) <= not (a and b);
    layer3_outputs(6387) <= not a or b;
    layer3_outputs(6388) <= a or b;
    layer3_outputs(6389) <= a;
    layer3_outputs(6390) <= not a or b;
    layer3_outputs(6391) <= '0';
    layer3_outputs(6392) <= b and not a;
    layer3_outputs(6393) <= a or b;
    layer3_outputs(6394) <= not b;
    layer3_outputs(6395) <= a and b;
    layer3_outputs(6396) <= not b;
    layer3_outputs(6397) <= not a or b;
    layer3_outputs(6398) <= a xor b;
    layer3_outputs(6399) <= a;
    layer3_outputs(6400) <= not (a and b);
    layer3_outputs(6401) <= '1';
    layer3_outputs(6402) <= '0';
    layer3_outputs(6403) <= '1';
    layer3_outputs(6404) <= '1';
    layer3_outputs(6405) <= a and b;
    layer3_outputs(6406) <= b and not a;
    layer3_outputs(6407) <= a and not b;
    layer3_outputs(6408) <= a;
    layer3_outputs(6409) <= not a;
    layer3_outputs(6410) <= not a;
    layer3_outputs(6411) <= a or b;
    layer3_outputs(6412) <= '0';
    layer3_outputs(6413) <= a and not b;
    layer3_outputs(6414) <= b and not a;
    layer3_outputs(6415) <= a;
    layer3_outputs(6416) <= not a or b;
    layer3_outputs(6417) <= b and not a;
    layer3_outputs(6418) <= a and not b;
    layer3_outputs(6419) <= not a;
    layer3_outputs(6420) <= not a;
    layer3_outputs(6421) <= a and not b;
    layer3_outputs(6422) <= '1';
    layer3_outputs(6423) <= not b;
    layer3_outputs(6424) <= a;
    layer3_outputs(6425) <= not b;
    layer3_outputs(6426) <= a and not b;
    layer3_outputs(6427) <= '0';
    layer3_outputs(6428) <= '1';
    layer3_outputs(6429) <= b and not a;
    layer3_outputs(6430) <= '1';
    layer3_outputs(6431) <= not b;
    layer3_outputs(6432) <= a or b;
    layer3_outputs(6433) <= a and not b;
    layer3_outputs(6434) <= a or b;
    layer3_outputs(6435) <= not a or b;
    layer3_outputs(6436) <= a and not b;
    layer3_outputs(6437) <= a and not b;
    layer3_outputs(6438) <= a;
    layer3_outputs(6439) <= a xor b;
    layer3_outputs(6440) <= not (a xor b);
    layer3_outputs(6441) <= not (a or b);
    layer3_outputs(6442) <= a;
    layer3_outputs(6443) <= b;
    layer3_outputs(6444) <= a and b;
    layer3_outputs(6445) <= b;
    layer3_outputs(6446) <= a and b;
    layer3_outputs(6447) <= '1';
    layer3_outputs(6448) <= b and not a;
    layer3_outputs(6449) <= b;
    layer3_outputs(6450) <= b and not a;
    layer3_outputs(6451) <= a and b;
    layer3_outputs(6452) <= not (a or b);
    layer3_outputs(6453) <= '0';
    layer3_outputs(6454) <= not a or b;
    layer3_outputs(6455) <= a and not b;
    layer3_outputs(6456) <= not b;
    layer3_outputs(6457) <= not b;
    layer3_outputs(6458) <= a or b;
    layer3_outputs(6459) <= b;
    layer3_outputs(6460) <= '0';
    layer3_outputs(6461) <= not (a and b);
    layer3_outputs(6462) <= a and not b;
    layer3_outputs(6463) <= not a or b;
    layer3_outputs(6464) <= not a;
    layer3_outputs(6465) <= not (a and b);
    layer3_outputs(6466) <= a and not b;
    layer3_outputs(6467) <= '1';
    layer3_outputs(6468) <= not b;
    layer3_outputs(6469) <= '0';
    layer3_outputs(6470) <= '1';
    layer3_outputs(6471) <= not (a xor b);
    layer3_outputs(6472) <= '1';
    layer3_outputs(6473) <= b;
    layer3_outputs(6474) <= b and not a;
    layer3_outputs(6475) <= a;
    layer3_outputs(6476) <= not a;
    layer3_outputs(6477) <= not (a or b);
    layer3_outputs(6478) <= '0';
    layer3_outputs(6479) <= not a or b;
    layer3_outputs(6480) <= '0';
    layer3_outputs(6481) <= '1';
    layer3_outputs(6482) <= not (a or b);
    layer3_outputs(6483) <= '0';
    layer3_outputs(6484) <= b and not a;
    layer3_outputs(6485) <= not a;
    layer3_outputs(6486) <= b and not a;
    layer3_outputs(6487) <= b;
    layer3_outputs(6488) <= a and not b;
    layer3_outputs(6489) <= not (a or b);
    layer3_outputs(6490) <= a;
    layer3_outputs(6491) <= a and not b;
    layer3_outputs(6492) <= a and b;
    layer3_outputs(6493) <= '1';
    layer3_outputs(6494) <= not (a or b);
    layer3_outputs(6495) <= b;
    layer3_outputs(6496) <= a and not b;
    layer3_outputs(6497) <= a;
    layer3_outputs(6498) <= a;
    layer3_outputs(6499) <= a and not b;
    layer3_outputs(6500) <= not a or b;
    layer3_outputs(6501) <= b and not a;
    layer3_outputs(6502) <= not b or a;
    layer3_outputs(6503) <= '0';
    layer3_outputs(6504) <= '1';
    layer3_outputs(6505) <= not a or b;
    layer3_outputs(6506) <= not (a or b);
    layer3_outputs(6507) <= a;
    layer3_outputs(6508) <= '0';
    layer3_outputs(6509) <= '1';
    layer3_outputs(6510) <= not a or b;
    layer3_outputs(6511) <= not b;
    layer3_outputs(6512) <= a;
    layer3_outputs(6513) <= b;
    layer3_outputs(6514) <= a and b;
    layer3_outputs(6515) <= b;
    layer3_outputs(6516) <= not (a and b);
    layer3_outputs(6517) <= '1';
    layer3_outputs(6518) <= not (a and b);
    layer3_outputs(6519) <= b;
    layer3_outputs(6520) <= not b or a;
    layer3_outputs(6521) <= not a or b;
    layer3_outputs(6522) <= not b;
    layer3_outputs(6523) <= b;
    layer3_outputs(6524) <= not b or a;
    layer3_outputs(6525) <= not b or a;
    layer3_outputs(6526) <= a;
    layer3_outputs(6527) <= a xor b;
    layer3_outputs(6528) <= b and not a;
    layer3_outputs(6529) <= not a;
    layer3_outputs(6530) <= not a or b;
    layer3_outputs(6531) <= not a;
    layer3_outputs(6532) <= a and b;
    layer3_outputs(6533) <= b and not a;
    layer3_outputs(6534) <= b and not a;
    layer3_outputs(6535) <= b and not a;
    layer3_outputs(6536) <= a;
    layer3_outputs(6537) <= a and not b;
    layer3_outputs(6538) <= '0';
    layer3_outputs(6539) <= not (a xor b);
    layer3_outputs(6540) <= not b or a;
    layer3_outputs(6541) <= not b or a;
    layer3_outputs(6542) <= a;
    layer3_outputs(6543) <= a or b;
    layer3_outputs(6544) <= not (a or b);
    layer3_outputs(6545) <= not (a and b);
    layer3_outputs(6546) <= a and b;
    layer3_outputs(6547) <= not a;
    layer3_outputs(6548) <= a;
    layer3_outputs(6549) <= not b;
    layer3_outputs(6550) <= not b or a;
    layer3_outputs(6551) <= not b;
    layer3_outputs(6552) <= a;
    layer3_outputs(6553) <= a and b;
    layer3_outputs(6554) <= a and b;
    layer3_outputs(6555) <= not a;
    layer3_outputs(6556) <= not b;
    layer3_outputs(6557) <= a and b;
    layer3_outputs(6558) <= not (a and b);
    layer3_outputs(6559) <= not (a or b);
    layer3_outputs(6560) <= '1';
    layer3_outputs(6561) <= not b or a;
    layer3_outputs(6562) <= not a or b;
    layer3_outputs(6563) <= '1';
    layer3_outputs(6564) <= not a or b;
    layer3_outputs(6565) <= not b or a;
    layer3_outputs(6566) <= a or b;
    layer3_outputs(6567) <= not (a or b);
    layer3_outputs(6568) <= a and b;
    layer3_outputs(6569) <= not b;
    layer3_outputs(6570) <= not (a and b);
    layer3_outputs(6571) <= not b;
    layer3_outputs(6572) <= not b;
    layer3_outputs(6573) <= not b;
    layer3_outputs(6574) <= '1';
    layer3_outputs(6575) <= b and not a;
    layer3_outputs(6576) <= b and not a;
    layer3_outputs(6577) <= a xor b;
    layer3_outputs(6578) <= not a;
    layer3_outputs(6579) <= a;
    layer3_outputs(6580) <= a;
    layer3_outputs(6581) <= not b or a;
    layer3_outputs(6582) <= a or b;
    layer3_outputs(6583) <= b and not a;
    layer3_outputs(6584) <= not a;
    layer3_outputs(6585) <= a;
    layer3_outputs(6586) <= not a;
    layer3_outputs(6587) <= not (a and b);
    layer3_outputs(6588) <= a;
    layer3_outputs(6589) <= b;
    layer3_outputs(6590) <= not (a and b);
    layer3_outputs(6591) <= a and b;
    layer3_outputs(6592) <= a;
    layer3_outputs(6593) <= a and not b;
    layer3_outputs(6594) <= not a;
    layer3_outputs(6595) <= not a;
    layer3_outputs(6596) <= '1';
    layer3_outputs(6597) <= not (a or b);
    layer3_outputs(6598) <= not (a and b);
    layer3_outputs(6599) <= not (a or b);
    layer3_outputs(6600) <= not (a and b);
    layer3_outputs(6601) <= b and not a;
    layer3_outputs(6602) <= a and b;
    layer3_outputs(6603) <= a xor b;
    layer3_outputs(6604) <= not b;
    layer3_outputs(6605) <= a and b;
    layer3_outputs(6606) <= '1';
    layer3_outputs(6607) <= not a;
    layer3_outputs(6608) <= '1';
    layer3_outputs(6609) <= not a or b;
    layer3_outputs(6610) <= '0';
    layer3_outputs(6611) <= not (a and b);
    layer3_outputs(6612) <= not (a or b);
    layer3_outputs(6613) <= not b or a;
    layer3_outputs(6614) <= b;
    layer3_outputs(6615) <= a or b;
    layer3_outputs(6616) <= '1';
    layer3_outputs(6617) <= not a;
    layer3_outputs(6618) <= not (a or b);
    layer3_outputs(6619) <= b;
    layer3_outputs(6620) <= not (a and b);
    layer3_outputs(6621) <= a and b;
    layer3_outputs(6622) <= a;
    layer3_outputs(6623) <= not (a and b);
    layer3_outputs(6624) <= not a or b;
    layer3_outputs(6625) <= '1';
    layer3_outputs(6626) <= b and not a;
    layer3_outputs(6627) <= a and b;
    layer3_outputs(6628) <= not a or b;
    layer3_outputs(6629) <= not b;
    layer3_outputs(6630) <= not (a or b);
    layer3_outputs(6631) <= not b;
    layer3_outputs(6632) <= a or b;
    layer3_outputs(6633) <= not a or b;
    layer3_outputs(6634) <= a;
    layer3_outputs(6635) <= not (a and b);
    layer3_outputs(6636) <= b;
    layer3_outputs(6637) <= b;
    layer3_outputs(6638) <= a and b;
    layer3_outputs(6639) <= not a;
    layer3_outputs(6640) <= '1';
    layer3_outputs(6641) <= not a;
    layer3_outputs(6642) <= a or b;
    layer3_outputs(6643) <= not (a xor b);
    layer3_outputs(6644) <= b and not a;
    layer3_outputs(6645) <= a or b;
    layer3_outputs(6646) <= not a;
    layer3_outputs(6647) <= not (a or b);
    layer3_outputs(6648) <= not (a and b);
    layer3_outputs(6649) <= not (a or b);
    layer3_outputs(6650) <= not (a and b);
    layer3_outputs(6651) <= not b;
    layer3_outputs(6652) <= '0';
    layer3_outputs(6653) <= a;
    layer3_outputs(6654) <= not (a and b);
    layer3_outputs(6655) <= b;
    layer3_outputs(6656) <= not b or a;
    layer3_outputs(6657) <= not (a or b);
    layer3_outputs(6658) <= not (a or b);
    layer3_outputs(6659) <= not a;
    layer3_outputs(6660) <= a or b;
    layer3_outputs(6661) <= a or b;
    layer3_outputs(6662) <= '1';
    layer3_outputs(6663) <= '1';
    layer3_outputs(6664) <= a xor b;
    layer3_outputs(6665) <= not (a or b);
    layer3_outputs(6666) <= a or b;
    layer3_outputs(6667) <= not b or a;
    layer3_outputs(6668) <= '0';
    layer3_outputs(6669) <= not (a and b);
    layer3_outputs(6670) <= not a or b;
    layer3_outputs(6671) <= not (a and b);
    layer3_outputs(6672) <= not (a and b);
    layer3_outputs(6673) <= '1';
    layer3_outputs(6674) <= not a;
    layer3_outputs(6675) <= '1';
    layer3_outputs(6676) <= not (a or b);
    layer3_outputs(6677) <= a and b;
    layer3_outputs(6678) <= not b;
    layer3_outputs(6679) <= '1';
    layer3_outputs(6680) <= not b;
    layer3_outputs(6681) <= not (a and b);
    layer3_outputs(6682) <= a and not b;
    layer3_outputs(6683) <= not a or b;
    layer3_outputs(6684) <= a or b;
    layer3_outputs(6685) <= not a;
    layer3_outputs(6686) <= not b or a;
    layer3_outputs(6687) <= not a or b;
    layer3_outputs(6688) <= not b;
    layer3_outputs(6689) <= '0';
    layer3_outputs(6690) <= a or b;
    layer3_outputs(6691) <= not (a and b);
    layer3_outputs(6692) <= not a or b;
    layer3_outputs(6693) <= not a or b;
    layer3_outputs(6694) <= not a;
    layer3_outputs(6695) <= b;
    layer3_outputs(6696) <= a and not b;
    layer3_outputs(6697) <= not (a and b);
    layer3_outputs(6698) <= not b;
    layer3_outputs(6699) <= not (a or b);
    layer3_outputs(6700) <= '0';
    layer3_outputs(6701) <= b;
    layer3_outputs(6702) <= not a;
    layer3_outputs(6703) <= a and not b;
    layer3_outputs(6704) <= '0';
    layer3_outputs(6705) <= a;
    layer3_outputs(6706) <= a and b;
    layer3_outputs(6707) <= a xor b;
    layer3_outputs(6708) <= a xor b;
    layer3_outputs(6709) <= '0';
    layer3_outputs(6710) <= not (a xor b);
    layer3_outputs(6711) <= b and not a;
    layer3_outputs(6712) <= a;
    layer3_outputs(6713) <= b;
    layer3_outputs(6714) <= a;
    layer3_outputs(6715) <= not (a and b);
    layer3_outputs(6716) <= not (a or b);
    layer3_outputs(6717) <= not (a or b);
    layer3_outputs(6718) <= not b;
    layer3_outputs(6719) <= not b;
    layer3_outputs(6720) <= not b or a;
    layer3_outputs(6721) <= not b;
    layer3_outputs(6722) <= a or b;
    layer3_outputs(6723) <= a xor b;
    layer3_outputs(6724) <= not (a and b);
    layer3_outputs(6725) <= a or b;
    layer3_outputs(6726) <= a and b;
    layer3_outputs(6727) <= not (a and b);
    layer3_outputs(6728) <= a;
    layer3_outputs(6729) <= not a or b;
    layer3_outputs(6730) <= b and not a;
    layer3_outputs(6731) <= b and not a;
    layer3_outputs(6732) <= a or b;
    layer3_outputs(6733) <= not (a or b);
    layer3_outputs(6734) <= not (a or b);
    layer3_outputs(6735) <= '1';
    layer3_outputs(6736) <= a;
    layer3_outputs(6737) <= b and not a;
    layer3_outputs(6738) <= not (a or b);
    layer3_outputs(6739) <= a or b;
    layer3_outputs(6740) <= a;
    layer3_outputs(6741) <= a;
    layer3_outputs(6742) <= '1';
    layer3_outputs(6743) <= a xor b;
    layer3_outputs(6744) <= '1';
    layer3_outputs(6745) <= not b or a;
    layer3_outputs(6746) <= not (a or b);
    layer3_outputs(6747) <= a and b;
    layer3_outputs(6748) <= '0';
    layer3_outputs(6749) <= not (a xor b);
    layer3_outputs(6750) <= not a or b;
    layer3_outputs(6751) <= not (a and b);
    layer3_outputs(6752) <= not (a or b);
    layer3_outputs(6753) <= a and not b;
    layer3_outputs(6754) <= not a;
    layer3_outputs(6755) <= not a or b;
    layer3_outputs(6756) <= a and b;
    layer3_outputs(6757) <= not a or b;
    layer3_outputs(6758) <= a and b;
    layer3_outputs(6759) <= '1';
    layer3_outputs(6760) <= a and b;
    layer3_outputs(6761) <= not a;
    layer3_outputs(6762) <= not a;
    layer3_outputs(6763) <= a and not b;
    layer3_outputs(6764) <= not (a and b);
    layer3_outputs(6765) <= a or b;
    layer3_outputs(6766) <= '1';
    layer3_outputs(6767) <= b and not a;
    layer3_outputs(6768) <= a xor b;
    layer3_outputs(6769) <= '1';
    layer3_outputs(6770) <= '1';
    layer3_outputs(6771) <= not (a and b);
    layer3_outputs(6772) <= a and not b;
    layer3_outputs(6773) <= '1';
    layer3_outputs(6774) <= a xor b;
    layer3_outputs(6775) <= a xor b;
    layer3_outputs(6776) <= not (a and b);
    layer3_outputs(6777) <= a or b;
    layer3_outputs(6778) <= not (a and b);
    layer3_outputs(6779) <= not (a or b);
    layer3_outputs(6780) <= a;
    layer3_outputs(6781) <= not a;
    layer3_outputs(6782) <= not (a or b);
    layer3_outputs(6783) <= a;
    layer3_outputs(6784) <= '0';
    layer3_outputs(6785) <= '0';
    layer3_outputs(6786) <= '0';
    layer3_outputs(6787) <= b and not a;
    layer3_outputs(6788) <= a and not b;
    layer3_outputs(6789) <= not b or a;
    layer3_outputs(6790) <= not (a xor b);
    layer3_outputs(6791) <= a or b;
    layer3_outputs(6792) <= a and b;
    layer3_outputs(6793) <= not b or a;
    layer3_outputs(6794) <= '1';
    layer3_outputs(6795) <= a xor b;
    layer3_outputs(6796) <= not (a and b);
    layer3_outputs(6797) <= a and b;
    layer3_outputs(6798) <= a and b;
    layer3_outputs(6799) <= a;
    layer3_outputs(6800) <= a xor b;
    layer3_outputs(6801) <= b and not a;
    layer3_outputs(6802) <= not b or a;
    layer3_outputs(6803) <= a and not b;
    layer3_outputs(6804) <= not a;
    layer3_outputs(6805) <= not (a or b);
    layer3_outputs(6806) <= not a;
    layer3_outputs(6807) <= not (a and b);
    layer3_outputs(6808) <= '1';
    layer3_outputs(6809) <= b and not a;
    layer3_outputs(6810) <= a and b;
    layer3_outputs(6811) <= not b;
    layer3_outputs(6812) <= '0';
    layer3_outputs(6813) <= not a or b;
    layer3_outputs(6814) <= a;
    layer3_outputs(6815) <= not b;
    layer3_outputs(6816) <= a and not b;
    layer3_outputs(6817) <= a and not b;
    layer3_outputs(6818) <= not (a or b);
    layer3_outputs(6819) <= b;
    layer3_outputs(6820) <= a or b;
    layer3_outputs(6821) <= not b;
    layer3_outputs(6822) <= a and not b;
    layer3_outputs(6823) <= '1';
    layer3_outputs(6824) <= not a;
    layer3_outputs(6825) <= not b or a;
    layer3_outputs(6826) <= a or b;
    layer3_outputs(6827) <= a or b;
    layer3_outputs(6828) <= not (a xor b);
    layer3_outputs(6829) <= a or b;
    layer3_outputs(6830) <= not b or a;
    layer3_outputs(6831) <= b and not a;
    layer3_outputs(6832) <= not a;
    layer3_outputs(6833) <= '1';
    layer3_outputs(6834) <= a or b;
    layer3_outputs(6835) <= not (a and b);
    layer3_outputs(6836) <= not b or a;
    layer3_outputs(6837) <= b;
    layer3_outputs(6838) <= not a;
    layer3_outputs(6839) <= not (a and b);
    layer3_outputs(6840) <= not b;
    layer3_outputs(6841) <= a and b;
    layer3_outputs(6842) <= not a or b;
    layer3_outputs(6843) <= not (a or b);
    layer3_outputs(6844) <= a;
    layer3_outputs(6845) <= not a;
    layer3_outputs(6846) <= not b or a;
    layer3_outputs(6847) <= '0';
    layer3_outputs(6848) <= not b or a;
    layer3_outputs(6849) <= not a;
    layer3_outputs(6850) <= b and not a;
    layer3_outputs(6851) <= not (a and b);
    layer3_outputs(6852) <= a and b;
    layer3_outputs(6853) <= b;
    layer3_outputs(6854) <= not b or a;
    layer3_outputs(6855) <= not b or a;
    layer3_outputs(6856) <= not a;
    layer3_outputs(6857) <= not b or a;
    layer3_outputs(6858) <= b;
    layer3_outputs(6859) <= not (a and b);
    layer3_outputs(6860) <= a and not b;
    layer3_outputs(6861) <= not (a and b);
    layer3_outputs(6862) <= not a or b;
    layer3_outputs(6863) <= b;
    layer3_outputs(6864) <= b;
    layer3_outputs(6865) <= a and b;
    layer3_outputs(6866) <= a or b;
    layer3_outputs(6867) <= a or b;
    layer3_outputs(6868) <= a and not b;
    layer3_outputs(6869) <= a or b;
    layer3_outputs(6870) <= not b;
    layer3_outputs(6871) <= not b;
    layer3_outputs(6872) <= '1';
    layer3_outputs(6873) <= not (a or b);
    layer3_outputs(6874) <= '1';
    layer3_outputs(6875) <= '1';
    layer3_outputs(6876) <= not a;
    layer3_outputs(6877) <= not b or a;
    layer3_outputs(6878) <= not b;
    layer3_outputs(6879) <= '1';
    layer3_outputs(6880) <= a xor b;
    layer3_outputs(6881) <= a and b;
    layer3_outputs(6882) <= not (a and b);
    layer3_outputs(6883) <= not (a and b);
    layer3_outputs(6884) <= b;
    layer3_outputs(6885) <= a;
    layer3_outputs(6886) <= not (a and b);
    layer3_outputs(6887) <= not b or a;
    layer3_outputs(6888) <= a or b;
    layer3_outputs(6889) <= a or b;
    layer3_outputs(6890) <= '1';
    layer3_outputs(6891) <= a and b;
    layer3_outputs(6892) <= not b or a;
    layer3_outputs(6893) <= b;
    layer3_outputs(6894) <= not (a or b);
    layer3_outputs(6895) <= not (a xor b);
    layer3_outputs(6896) <= a and not b;
    layer3_outputs(6897) <= not a;
    layer3_outputs(6898) <= b;
    layer3_outputs(6899) <= '0';
    layer3_outputs(6900) <= '0';
    layer3_outputs(6901) <= not a;
    layer3_outputs(6902) <= b and not a;
    layer3_outputs(6903) <= b and not a;
    layer3_outputs(6904) <= a xor b;
    layer3_outputs(6905) <= '0';
    layer3_outputs(6906) <= a or b;
    layer3_outputs(6907) <= not (a or b);
    layer3_outputs(6908) <= a and not b;
    layer3_outputs(6909) <= not a or b;
    layer3_outputs(6910) <= not (a or b);
    layer3_outputs(6911) <= not (a and b);
    layer3_outputs(6912) <= b and not a;
    layer3_outputs(6913) <= '1';
    layer3_outputs(6914) <= a and b;
    layer3_outputs(6915) <= a;
    layer3_outputs(6916) <= not (a or b);
    layer3_outputs(6917) <= b and not a;
    layer3_outputs(6918) <= b;
    layer3_outputs(6919) <= not a or b;
    layer3_outputs(6920) <= '0';
    layer3_outputs(6921) <= not a;
    layer3_outputs(6922) <= a and b;
    layer3_outputs(6923) <= a and not b;
    layer3_outputs(6924) <= not (a and b);
    layer3_outputs(6925) <= not b;
    layer3_outputs(6926) <= b and not a;
    layer3_outputs(6927) <= a and not b;
    layer3_outputs(6928) <= '1';
    layer3_outputs(6929) <= not b or a;
    layer3_outputs(6930) <= a and not b;
    layer3_outputs(6931) <= not (a and b);
    layer3_outputs(6932) <= '0';
    layer3_outputs(6933) <= not b or a;
    layer3_outputs(6934) <= '0';
    layer3_outputs(6935) <= not b;
    layer3_outputs(6936) <= not a;
    layer3_outputs(6937) <= '1';
    layer3_outputs(6938) <= '0';
    layer3_outputs(6939) <= not a;
    layer3_outputs(6940) <= a xor b;
    layer3_outputs(6941) <= b and not a;
    layer3_outputs(6942) <= '0';
    layer3_outputs(6943) <= not b;
    layer3_outputs(6944) <= '1';
    layer3_outputs(6945) <= '0';
    layer3_outputs(6946) <= not (a and b);
    layer3_outputs(6947) <= not a or b;
    layer3_outputs(6948) <= not (a and b);
    layer3_outputs(6949) <= not (a and b);
    layer3_outputs(6950) <= not (a or b);
    layer3_outputs(6951) <= not b or a;
    layer3_outputs(6952) <= b;
    layer3_outputs(6953) <= a and not b;
    layer3_outputs(6954) <= not b;
    layer3_outputs(6955) <= not a;
    layer3_outputs(6956) <= not (a or b);
    layer3_outputs(6957) <= not a or b;
    layer3_outputs(6958) <= not b or a;
    layer3_outputs(6959) <= b and not a;
    layer3_outputs(6960) <= not b;
    layer3_outputs(6961) <= a;
    layer3_outputs(6962) <= b;
    layer3_outputs(6963) <= not b or a;
    layer3_outputs(6964) <= b and not a;
    layer3_outputs(6965) <= a xor b;
    layer3_outputs(6966) <= '0';
    layer3_outputs(6967) <= not (a and b);
    layer3_outputs(6968) <= not (a and b);
    layer3_outputs(6969) <= a and b;
    layer3_outputs(6970) <= b and not a;
    layer3_outputs(6971) <= not a or b;
    layer3_outputs(6972) <= not b or a;
    layer3_outputs(6973) <= a and b;
    layer3_outputs(6974) <= not a or b;
    layer3_outputs(6975) <= '0';
    layer3_outputs(6976) <= b and not a;
    layer3_outputs(6977) <= not b;
    layer3_outputs(6978) <= b;
    layer3_outputs(6979) <= not (a or b);
    layer3_outputs(6980) <= b and not a;
    layer3_outputs(6981) <= a and not b;
    layer3_outputs(6982) <= a and not b;
    layer3_outputs(6983) <= not (a or b);
    layer3_outputs(6984) <= a and not b;
    layer3_outputs(6985) <= a and b;
    layer3_outputs(6986) <= not (a xor b);
    layer3_outputs(6987) <= b;
    layer3_outputs(6988) <= not a;
    layer3_outputs(6989) <= '0';
    layer3_outputs(6990) <= a;
    layer3_outputs(6991) <= a xor b;
    layer3_outputs(6992) <= b and not a;
    layer3_outputs(6993) <= a and not b;
    layer3_outputs(6994) <= not (a xor b);
    layer3_outputs(6995) <= a and not b;
    layer3_outputs(6996) <= b and not a;
    layer3_outputs(6997) <= a;
    layer3_outputs(6998) <= a and b;
    layer3_outputs(6999) <= not b or a;
    layer3_outputs(7000) <= not a;
    layer3_outputs(7001) <= not (a or b);
    layer3_outputs(7002) <= a and not b;
    layer3_outputs(7003) <= a and not b;
    layer3_outputs(7004) <= not (a and b);
    layer3_outputs(7005) <= not b or a;
    layer3_outputs(7006) <= b and not a;
    layer3_outputs(7007) <= '0';
    layer3_outputs(7008) <= a and not b;
    layer3_outputs(7009) <= not (a or b);
    layer3_outputs(7010) <= not b;
    layer3_outputs(7011) <= not a;
    layer3_outputs(7012) <= a;
    layer3_outputs(7013) <= a and not b;
    layer3_outputs(7014) <= b and not a;
    layer3_outputs(7015) <= not a or b;
    layer3_outputs(7016) <= not (a or b);
    layer3_outputs(7017) <= a and b;
    layer3_outputs(7018) <= not b or a;
    layer3_outputs(7019) <= '0';
    layer3_outputs(7020) <= b;
    layer3_outputs(7021) <= a and not b;
    layer3_outputs(7022) <= b;
    layer3_outputs(7023) <= '0';
    layer3_outputs(7024) <= a;
    layer3_outputs(7025) <= a;
    layer3_outputs(7026) <= b;
    layer3_outputs(7027) <= b and not a;
    layer3_outputs(7028) <= a;
    layer3_outputs(7029) <= a and b;
    layer3_outputs(7030) <= a;
    layer3_outputs(7031) <= not (a or b);
    layer3_outputs(7032) <= '0';
    layer3_outputs(7033) <= a and not b;
    layer3_outputs(7034) <= a and not b;
    layer3_outputs(7035) <= b and not a;
    layer3_outputs(7036) <= b and not a;
    layer3_outputs(7037) <= a or b;
    layer3_outputs(7038) <= not (a and b);
    layer3_outputs(7039) <= not (a or b);
    layer3_outputs(7040) <= not a;
    layer3_outputs(7041) <= a or b;
    layer3_outputs(7042) <= not (a or b);
    layer3_outputs(7043) <= not (a or b);
    layer3_outputs(7044) <= not a;
    layer3_outputs(7045) <= b;
    layer3_outputs(7046) <= not a or b;
    layer3_outputs(7047) <= b;
    layer3_outputs(7048) <= not a or b;
    layer3_outputs(7049) <= not (a or b);
    layer3_outputs(7050) <= not a;
    layer3_outputs(7051) <= not (a and b);
    layer3_outputs(7052) <= a;
    layer3_outputs(7053) <= '0';
    layer3_outputs(7054) <= a;
    layer3_outputs(7055) <= a xor b;
    layer3_outputs(7056) <= not (a or b);
    layer3_outputs(7057) <= not a or b;
    layer3_outputs(7058) <= not b or a;
    layer3_outputs(7059) <= not a;
    layer3_outputs(7060) <= not a;
    layer3_outputs(7061) <= a and b;
    layer3_outputs(7062) <= b and not a;
    layer3_outputs(7063) <= not a or b;
    layer3_outputs(7064) <= not a or b;
    layer3_outputs(7065) <= a and b;
    layer3_outputs(7066) <= b and not a;
    layer3_outputs(7067) <= a and b;
    layer3_outputs(7068) <= not (a and b);
    layer3_outputs(7069) <= '0';
    layer3_outputs(7070) <= b;
    layer3_outputs(7071) <= not (a or b);
    layer3_outputs(7072) <= a xor b;
    layer3_outputs(7073) <= b and not a;
    layer3_outputs(7074) <= not b or a;
    layer3_outputs(7075) <= not (a xor b);
    layer3_outputs(7076) <= a;
    layer3_outputs(7077) <= not a;
    layer3_outputs(7078) <= a;
    layer3_outputs(7079) <= b and not a;
    layer3_outputs(7080) <= b and not a;
    layer3_outputs(7081) <= not a or b;
    layer3_outputs(7082) <= not b or a;
    layer3_outputs(7083) <= not b;
    layer3_outputs(7084) <= a or b;
    layer3_outputs(7085) <= '1';
    layer3_outputs(7086) <= not b or a;
    layer3_outputs(7087) <= a or b;
    layer3_outputs(7088) <= a and b;
    layer3_outputs(7089) <= a or b;
    layer3_outputs(7090) <= a and b;
    layer3_outputs(7091) <= a and not b;
    layer3_outputs(7092) <= a or b;
    layer3_outputs(7093) <= '0';
    layer3_outputs(7094) <= not a;
    layer3_outputs(7095) <= not (a xor b);
    layer3_outputs(7096) <= not a or b;
    layer3_outputs(7097) <= not b or a;
    layer3_outputs(7098) <= a or b;
    layer3_outputs(7099) <= not b or a;
    layer3_outputs(7100) <= a;
    layer3_outputs(7101) <= not (a or b);
    layer3_outputs(7102) <= b and not a;
    layer3_outputs(7103) <= '1';
    layer3_outputs(7104) <= not b or a;
    layer3_outputs(7105) <= not a;
    layer3_outputs(7106) <= not b or a;
    layer3_outputs(7107) <= a or b;
    layer3_outputs(7108) <= not a or b;
    layer3_outputs(7109) <= not b;
    layer3_outputs(7110) <= a and b;
    layer3_outputs(7111) <= a;
    layer3_outputs(7112) <= not (a xor b);
    layer3_outputs(7113) <= not (a or b);
    layer3_outputs(7114) <= '1';
    layer3_outputs(7115) <= not b;
    layer3_outputs(7116) <= not b or a;
    layer3_outputs(7117) <= not (a or b);
    layer3_outputs(7118) <= '0';
    layer3_outputs(7119) <= a or b;
    layer3_outputs(7120) <= not a;
    layer3_outputs(7121) <= a xor b;
    layer3_outputs(7122) <= b;
    layer3_outputs(7123) <= a and not b;
    layer3_outputs(7124) <= '0';
    layer3_outputs(7125) <= not (a or b);
    layer3_outputs(7126) <= a or b;
    layer3_outputs(7127) <= not a;
    layer3_outputs(7128) <= a and not b;
    layer3_outputs(7129) <= a xor b;
    layer3_outputs(7130) <= not b or a;
    layer3_outputs(7131) <= not a or b;
    layer3_outputs(7132) <= b and not a;
    layer3_outputs(7133) <= '0';
    layer3_outputs(7134) <= '0';
    layer3_outputs(7135) <= b;
    layer3_outputs(7136) <= '1';
    layer3_outputs(7137) <= a or b;
    layer3_outputs(7138) <= '0';
    layer3_outputs(7139) <= b;
    layer3_outputs(7140) <= not b;
    layer3_outputs(7141) <= not b or a;
    layer3_outputs(7142) <= not a or b;
    layer3_outputs(7143) <= b;
    layer3_outputs(7144) <= not b or a;
    layer3_outputs(7145) <= b and not a;
    layer3_outputs(7146) <= not (a or b);
    layer3_outputs(7147) <= '0';
    layer3_outputs(7148) <= a and not b;
    layer3_outputs(7149) <= a and b;
    layer3_outputs(7150) <= not a or b;
    layer3_outputs(7151) <= a;
    layer3_outputs(7152) <= not (a xor b);
    layer3_outputs(7153) <= a and b;
    layer3_outputs(7154) <= not (a or b);
    layer3_outputs(7155) <= not (a and b);
    layer3_outputs(7156) <= a or b;
    layer3_outputs(7157) <= a;
    layer3_outputs(7158) <= '1';
    layer3_outputs(7159) <= a;
    layer3_outputs(7160) <= a and b;
    layer3_outputs(7161) <= not a or b;
    layer3_outputs(7162) <= not a or b;
    layer3_outputs(7163) <= a or b;
    layer3_outputs(7164) <= a or b;
    layer3_outputs(7165) <= a xor b;
    layer3_outputs(7166) <= not b or a;
    layer3_outputs(7167) <= b;
    layer3_outputs(7168) <= '1';
    layer3_outputs(7169) <= a and not b;
    layer3_outputs(7170) <= a and not b;
    layer3_outputs(7171) <= '0';
    layer3_outputs(7172) <= not (a or b);
    layer3_outputs(7173) <= not a or b;
    layer3_outputs(7174) <= not a;
    layer3_outputs(7175) <= b and not a;
    layer3_outputs(7176) <= not (a and b);
    layer3_outputs(7177) <= not (a or b);
    layer3_outputs(7178) <= not b;
    layer3_outputs(7179) <= '0';
    layer3_outputs(7180) <= not b;
    layer3_outputs(7181) <= '0';
    layer3_outputs(7182) <= not (a xor b);
    layer3_outputs(7183) <= a and not b;
    layer3_outputs(7184) <= '0';
    layer3_outputs(7185) <= a and b;
    layer3_outputs(7186) <= not b;
    layer3_outputs(7187) <= '1';
    layer3_outputs(7188) <= not b or a;
    layer3_outputs(7189) <= b and not a;
    layer3_outputs(7190) <= not a or b;
    layer3_outputs(7191) <= not b;
    layer3_outputs(7192) <= a and b;
    layer3_outputs(7193) <= not b;
    layer3_outputs(7194) <= b;
    layer3_outputs(7195) <= not b;
    layer3_outputs(7196) <= not b;
    layer3_outputs(7197) <= not b or a;
    layer3_outputs(7198) <= a;
    layer3_outputs(7199) <= not b or a;
    layer3_outputs(7200) <= a and b;
    layer3_outputs(7201) <= not (a or b);
    layer3_outputs(7202) <= a or b;
    layer3_outputs(7203) <= not (a or b);
    layer3_outputs(7204) <= not (a and b);
    layer3_outputs(7205) <= '1';
    layer3_outputs(7206) <= b and not a;
    layer3_outputs(7207) <= not b or a;
    layer3_outputs(7208) <= a or b;
    layer3_outputs(7209) <= a xor b;
    layer3_outputs(7210) <= a and not b;
    layer3_outputs(7211) <= a and not b;
    layer3_outputs(7212) <= not a;
    layer3_outputs(7213) <= a;
    layer3_outputs(7214) <= '0';
    layer3_outputs(7215) <= not (a and b);
    layer3_outputs(7216) <= not b or a;
    layer3_outputs(7217) <= a or b;
    layer3_outputs(7218) <= b and not a;
    layer3_outputs(7219) <= a or b;
    layer3_outputs(7220) <= not b;
    layer3_outputs(7221) <= not b;
    layer3_outputs(7222) <= b and not a;
    layer3_outputs(7223) <= not a or b;
    layer3_outputs(7224) <= a and not b;
    layer3_outputs(7225) <= not a;
    layer3_outputs(7226) <= not b or a;
    layer3_outputs(7227) <= not a or b;
    layer3_outputs(7228) <= a or b;
    layer3_outputs(7229) <= not a or b;
    layer3_outputs(7230) <= b;
    layer3_outputs(7231) <= b and not a;
    layer3_outputs(7232) <= '1';
    layer3_outputs(7233) <= not a;
    layer3_outputs(7234) <= not a or b;
    layer3_outputs(7235) <= a;
    layer3_outputs(7236) <= a and b;
    layer3_outputs(7237) <= not a;
    layer3_outputs(7238) <= '1';
    layer3_outputs(7239) <= a;
    layer3_outputs(7240) <= not (a and b);
    layer3_outputs(7241) <= not (a and b);
    layer3_outputs(7242) <= a and b;
    layer3_outputs(7243) <= '0';
    layer3_outputs(7244) <= a;
    layer3_outputs(7245) <= not a;
    layer3_outputs(7246) <= not (a xor b);
    layer3_outputs(7247) <= not b;
    layer3_outputs(7248) <= not (a or b);
    layer3_outputs(7249) <= a;
    layer3_outputs(7250) <= a and b;
    layer3_outputs(7251) <= a and b;
    layer3_outputs(7252) <= not b;
    layer3_outputs(7253) <= a;
    layer3_outputs(7254) <= a;
    layer3_outputs(7255) <= not (a or b);
    layer3_outputs(7256) <= a;
    layer3_outputs(7257) <= a or b;
    layer3_outputs(7258) <= not b;
    layer3_outputs(7259) <= b;
    layer3_outputs(7260) <= a or b;
    layer3_outputs(7261) <= not b;
    layer3_outputs(7262) <= not a;
    layer3_outputs(7263) <= a and not b;
    layer3_outputs(7264) <= b;
    layer3_outputs(7265) <= not b or a;
    layer3_outputs(7266) <= a and not b;
    layer3_outputs(7267) <= a xor b;
    layer3_outputs(7268) <= '1';
    layer3_outputs(7269) <= a and not b;
    layer3_outputs(7270) <= b;
    layer3_outputs(7271) <= a or b;
    layer3_outputs(7272) <= not (a xor b);
    layer3_outputs(7273) <= not a or b;
    layer3_outputs(7274) <= b and not a;
    layer3_outputs(7275) <= b;
    layer3_outputs(7276) <= a or b;
    layer3_outputs(7277) <= b and not a;
    layer3_outputs(7278) <= a or b;
    layer3_outputs(7279) <= a and b;
    layer3_outputs(7280) <= b and not a;
    layer3_outputs(7281) <= not b;
    layer3_outputs(7282) <= not b or a;
    layer3_outputs(7283) <= not a;
    layer3_outputs(7284) <= not b;
    layer3_outputs(7285) <= not a or b;
    layer3_outputs(7286) <= a and b;
    layer3_outputs(7287) <= not a;
    layer3_outputs(7288) <= '0';
    layer3_outputs(7289) <= a and not b;
    layer3_outputs(7290) <= a and b;
    layer3_outputs(7291) <= not (a or b);
    layer3_outputs(7292) <= not b or a;
    layer3_outputs(7293) <= not (a or b);
    layer3_outputs(7294) <= b and not a;
    layer3_outputs(7295) <= not b;
    layer3_outputs(7296) <= a and b;
    layer3_outputs(7297) <= '0';
    layer3_outputs(7298) <= not (a or b);
    layer3_outputs(7299) <= not b or a;
    layer3_outputs(7300) <= b and not a;
    layer3_outputs(7301) <= a and not b;
    layer3_outputs(7302) <= b;
    layer3_outputs(7303) <= '0';
    layer3_outputs(7304) <= b and not a;
    layer3_outputs(7305) <= not a or b;
    layer3_outputs(7306) <= b;
    layer3_outputs(7307) <= a or b;
    layer3_outputs(7308) <= a;
    layer3_outputs(7309) <= b and not a;
    layer3_outputs(7310) <= not a;
    layer3_outputs(7311) <= not (a xor b);
    layer3_outputs(7312) <= '1';
    layer3_outputs(7313) <= a and b;
    layer3_outputs(7314) <= '1';
    layer3_outputs(7315) <= not a;
    layer3_outputs(7316) <= '1';
    layer3_outputs(7317) <= '1';
    layer3_outputs(7318) <= not b;
    layer3_outputs(7319) <= not b or a;
    layer3_outputs(7320) <= a or b;
    layer3_outputs(7321) <= b;
    layer3_outputs(7322) <= '0';
    layer3_outputs(7323) <= b;
    layer3_outputs(7324) <= not (a and b);
    layer3_outputs(7325) <= not (a or b);
    layer3_outputs(7326) <= not (a xor b);
    layer3_outputs(7327) <= '1';
    layer3_outputs(7328) <= b;
    layer3_outputs(7329) <= a and b;
    layer3_outputs(7330) <= '0';
    layer3_outputs(7331) <= not a or b;
    layer3_outputs(7332) <= a and not b;
    layer3_outputs(7333) <= a and not b;
    layer3_outputs(7334) <= not b or a;
    layer3_outputs(7335) <= a;
    layer3_outputs(7336) <= not (a or b);
    layer3_outputs(7337) <= '1';
    layer3_outputs(7338) <= not (a and b);
    layer3_outputs(7339) <= b;
    layer3_outputs(7340) <= a;
    layer3_outputs(7341) <= a or b;
    layer3_outputs(7342) <= '0';
    layer3_outputs(7343) <= not b or a;
    layer3_outputs(7344) <= not (a and b);
    layer3_outputs(7345) <= not b;
    layer3_outputs(7346) <= '1';
    layer3_outputs(7347) <= not a;
    layer3_outputs(7348) <= b and not a;
    layer3_outputs(7349) <= not (a and b);
    layer3_outputs(7350) <= not a;
    layer3_outputs(7351) <= a and b;
    layer3_outputs(7352) <= a and b;
    layer3_outputs(7353) <= '1';
    layer3_outputs(7354) <= not b;
    layer3_outputs(7355) <= a or b;
    layer3_outputs(7356) <= a;
    layer3_outputs(7357) <= not a;
    layer3_outputs(7358) <= '0';
    layer3_outputs(7359) <= a or b;
    layer3_outputs(7360) <= not a or b;
    layer3_outputs(7361) <= '1';
    layer3_outputs(7362) <= b and not a;
    layer3_outputs(7363) <= a;
    layer3_outputs(7364) <= '0';
    layer3_outputs(7365) <= not a or b;
    layer3_outputs(7366) <= b and not a;
    layer3_outputs(7367) <= a;
    layer3_outputs(7368) <= not (a or b);
    layer3_outputs(7369) <= '0';
    layer3_outputs(7370) <= not (a and b);
    layer3_outputs(7371) <= '1';
    layer3_outputs(7372) <= a xor b;
    layer3_outputs(7373) <= not (a and b);
    layer3_outputs(7374) <= b and not a;
    layer3_outputs(7375) <= b;
    layer3_outputs(7376) <= not b or a;
    layer3_outputs(7377) <= b;
    layer3_outputs(7378) <= '1';
    layer3_outputs(7379) <= '0';
    layer3_outputs(7380) <= '1';
    layer3_outputs(7381) <= not (a and b);
    layer3_outputs(7382) <= not (a and b);
    layer3_outputs(7383) <= not b;
    layer3_outputs(7384) <= not (a xor b);
    layer3_outputs(7385) <= b;
    layer3_outputs(7386) <= a or b;
    layer3_outputs(7387) <= a;
    layer3_outputs(7388) <= not a;
    layer3_outputs(7389) <= b;
    layer3_outputs(7390) <= b and not a;
    layer3_outputs(7391) <= a;
    layer3_outputs(7392) <= not (a and b);
    layer3_outputs(7393) <= not b or a;
    layer3_outputs(7394) <= '1';
    layer3_outputs(7395) <= not a;
    layer3_outputs(7396) <= not a or b;
    layer3_outputs(7397) <= not (a and b);
    layer3_outputs(7398) <= a and b;
    layer3_outputs(7399) <= b;
    layer3_outputs(7400) <= a or b;
    layer3_outputs(7401) <= a xor b;
    layer3_outputs(7402) <= a or b;
    layer3_outputs(7403) <= b;
    layer3_outputs(7404) <= b;
    layer3_outputs(7405) <= not (a and b);
    layer3_outputs(7406) <= not (a and b);
    layer3_outputs(7407) <= not a or b;
    layer3_outputs(7408) <= a or b;
    layer3_outputs(7409) <= b and not a;
    layer3_outputs(7410) <= not b;
    layer3_outputs(7411) <= not a;
    layer3_outputs(7412) <= '0';
    layer3_outputs(7413) <= not a;
    layer3_outputs(7414) <= a or b;
    layer3_outputs(7415) <= not a;
    layer3_outputs(7416) <= not a;
    layer3_outputs(7417) <= a and not b;
    layer3_outputs(7418) <= a;
    layer3_outputs(7419) <= b;
    layer3_outputs(7420) <= not b or a;
    layer3_outputs(7421) <= not a;
    layer3_outputs(7422) <= '0';
    layer3_outputs(7423) <= a;
    layer3_outputs(7424) <= b;
    layer3_outputs(7425) <= a;
    layer3_outputs(7426) <= not (a or b);
    layer3_outputs(7427) <= not a or b;
    layer3_outputs(7428) <= not a;
    layer3_outputs(7429) <= not a;
    layer3_outputs(7430) <= a;
    layer3_outputs(7431) <= a xor b;
    layer3_outputs(7432) <= not a;
    layer3_outputs(7433) <= b;
    layer3_outputs(7434) <= not (a xor b);
    layer3_outputs(7435) <= b;
    layer3_outputs(7436) <= a and not b;
    layer3_outputs(7437) <= a or b;
    layer3_outputs(7438) <= a;
    layer3_outputs(7439) <= not b;
    layer3_outputs(7440) <= b;
    layer3_outputs(7441) <= a and not b;
    layer3_outputs(7442) <= not b or a;
    layer3_outputs(7443) <= not a or b;
    layer3_outputs(7444) <= not a;
    layer3_outputs(7445) <= a and not b;
    layer3_outputs(7446) <= not (a or b);
    layer3_outputs(7447) <= a and not b;
    layer3_outputs(7448) <= not b or a;
    layer3_outputs(7449) <= b;
    layer3_outputs(7450) <= b and not a;
    layer3_outputs(7451) <= a and b;
    layer3_outputs(7452) <= not b or a;
    layer3_outputs(7453) <= b;
    layer3_outputs(7454) <= not (a and b);
    layer3_outputs(7455) <= not b or a;
    layer3_outputs(7456) <= not a;
    layer3_outputs(7457) <= a;
    layer3_outputs(7458) <= not a or b;
    layer3_outputs(7459) <= b and not a;
    layer3_outputs(7460) <= not a;
    layer3_outputs(7461) <= not a or b;
    layer3_outputs(7462) <= not (a and b);
    layer3_outputs(7463) <= not a or b;
    layer3_outputs(7464) <= a and not b;
    layer3_outputs(7465) <= not b;
    layer3_outputs(7466) <= a;
    layer3_outputs(7467) <= '0';
    layer3_outputs(7468) <= '0';
    layer3_outputs(7469) <= a and not b;
    layer3_outputs(7470) <= '1';
    layer3_outputs(7471) <= b;
    layer3_outputs(7472) <= '1';
    layer3_outputs(7473) <= '0';
    layer3_outputs(7474) <= '1';
    layer3_outputs(7475) <= not a;
    layer3_outputs(7476) <= '0';
    layer3_outputs(7477) <= a or b;
    layer3_outputs(7478) <= not a or b;
    layer3_outputs(7479) <= not b or a;
    layer3_outputs(7480) <= not a;
    layer3_outputs(7481) <= a and b;
    layer3_outputs(7482) <= a and not b;
    layer3_outputs(7483) <= '0';
    layer3_outputs(7484) <= a xor b;
    layer3_outputs(7485) <= not a;
    layer3_outputs(7486) <= not b or a;
    layer3_outputs(7487) <= b and not a;
    layer3_outputs(7488) <= a and not b;
    layer3_outputs(7489) <= not (a or b);
    layer3_outputs(7490) <= not b;
    layer3_outputs(7491) <= not a;
    layer3_outputs(7492) <= not b or a;
    layer3_outputs(7493) <= a;
    layer3_outputs(7494) <= not a or b;
    layer3_outputs(7495) <= not (a or b);
    layer3_outputs(7496) <= not a;
    layer3_outputs(7497) <= b and not a;
    layer3_outputs(7498) <= a and b;
    layer3_outputs(7499) <= b and not a;
    layer3_outputs(7500) <= b and not a;
    layer3_outputs(7501) <= a xor b;
    layer3_outputs(7502) <= a and not b;
    layer3_outputs(7503) <= not (a and b);
    layer3_outputs(7504) <= not a;
    layer3_outputs(7505) <= not b;
    layer3_outputs(7506) <= a and not b;
    layer3_outputs(7507) <= '1';
    layer3_outputs(7508) <= not b;
    layer3_outputs(7509) <= a xor b;
    layer3_outputs(7510) <= not (a or b);
    layer3_outputs(7511) <= a and b;
    layer3_outputs(7512) <= not (a xor b);
    layer3_outputs(7513) <= not b;
    layer3_outputs(7514) <= not b or a;
    layer3_outputs(7515) <= a;
    layer3_outputs(7516) <= a and not b;
    layer3_outputs(7517) <= not b or a;
    layer3_outputs(7518) <= a and not b;
    layer3_outputs(7519) <= not b;
    layer3_outputs(7520) <= b and not a;
    layer3_outputs(7521) <= not b or a;
    layer3_outputs(7522) <= not (a or b);
    layer3_outputs(7523) <= not (a and b);
    layer3_outputs(7524) <= a and not b;
    layer3_outputs(7525) <= a;
    layer3_outputs(7526) <= not (a and b);
    layer3_outputs(7527) <= not a or b;
    layer3_outputs(7528) <= a and not b;
    layer3_outputs(7529) <= '0';
    layer3_outputs(7530) <= not a or b;
    layer3_outputs(7531) <= not a or b;
    layer3_outputs(7532) <= '1';
    layer3_outputs(7533) <= not b or a;
    layer3_outputs(7534) <= a or b;
    layer3_outputs(7535) <= not a or b;
    layer3_outputs(7536) <= a and b;
    layer3_outputs(7537) <= not a;
    layer3_outputs(7538) <= not a or b;
    layer3_outputs(7539) <= b and not a;
    layer3_outputs(7540) <= b and not a;
    layer3_outputs(7541) <= a or b;
    layer3_outputs(7542) <= not a or b;
    layer3_outputs(7543) <= b and not a;
    layer3_outputs(7544) <= a and not b;
    layer3_outputs(7545) <= a and b;
    layer3_outputs(7546) <= a and not b;
    layer3_outputs(7547) <= not b or a;
    layer3_outputs(7548) <= '1';
    layer3_outputs(7549) <= '0';
    layer3_outputs(7550) <= not b or a;
    layer3_outputs(7551) <= '1';
    layer3_outputs(7552) <= b and not a;
    layer3_outputs(7553) <= not (a xor b);
    layer3_outputs(7554) <= not b;
    layer3_outputs(7555) <= b;
    layer3_outputs(7556) <= not a or b;
    layer3_outputs(7557) <= '1';
    layer3_outputs(7558) <= not a or b;
    layer3_outputs(7559) <= not (a or b);
    layer3_outputs(7560) <= not (a or b);
    layer3_outputs(7561) <= a and b;
    layer3_outputs(7562) <= not (a or b);
    layer3_outputs(7563) <= '1';
    layer3_outputs(7564) <= not a;
    layer3_outputs(7565) <= not b;
    layer3_outputs(7566) <= not (a and b);
    layer3_outputs(7567) <= b and not a;
    layer3_outputs(7568) <= a or b;
    layer3_outputs(7569) <= '0';
    layer3_outputs(7570) <= a;
    layer3_outputs(7571) <= '1';
    layer3_outputs(7572) <= a and b;
    layer3_outputs(7573) <= a and b;
    layer3_outputs(7574) <= a and b;
    layer3_outputs(7575) <= a xor b;
    layer3_outputs(7576) <= not a or b;
    layer3_outputs(7577) <= b;
    layer3_outputs(7578) <= b;
    layer3_outputs(7579) <= not (a or b);
    layer3_outputs(7580) <= not a or b;
    layer3_outputs(7581) <= a;
    layer3_outputs(7582) <= not b;
    layer3_outputs(7583) <= a and not b;
    layer3_outputs(7584) <= '1';
    layer3_outputs(7585) <= b;
    layer3_outputs(7586) <= not b;
    layer3_outputs(7587) <= not (a and b);
    layer3_outputs(7588) <= a and not b;
    layer3_outputs(7589) <= '1';
    layer3_outputs(7590) <= b;
    layer3_outputs(7591) <= not a;
    layer3_outputs(7592) <= a xor b;
    layer3_outputs(7593) <= '0';
    layer3_outputs(7594) <= '0';
    layer3_outputs(7595) <= not (a and b);
    layer3_outputs(7596) <= not a;
    layer3_outputs(7597) <= not b or a;
    layer3_outputs(7598) <= not (a and b);
    layer3_outputs(7599) <= not (a or b);
    layer3_outputs(7600) <= a and not b;
    layer3_outputs(7601) <= '1';
    layer3_outputs(7602) <= a;
    layer3_outputs(7603) <= b and not a;
    layer3_outputs(7604) <= not a or b;
    layer3_outputs(7605) <= '0';
    layer3_outputs(7606) <= not (a and b);
    layer3_outputs(7607) <= not b or a;
    layer3_outputs(7608) <= b and not a;
    layer3_outputs(7609) <= not (a xor b);
    layer3_outputs(7610) <= not a or b;
    layer3_outputs(7611) <= not (a or b);
    layer3_outputs(7612) <= a and b;
    layer3_outputs(7613) <= a;
    layer3_outputs(7614) <= '1';
    layer3_outputs(7615) <= not a;
    layer3_outputs(7616) <= not a or b;
    layer3_outputs(7617) <= a xor b;
    layer3_outputs(7618) <= not b;
    layer3_outputs(7619) <= a and b;
    layer3_outputs(7620) <= b and not a;
    layer3_outputs(7621) <= a and b;
    layer3_outputs(7622) <= a and b;
    layer3_outputs(7623) <= a or b;
    layer3_outputs(7624) <= b;
    layer3_outputs(7625) <= a or b;
    layer3_outputs(7626) <= not (a or b);
    layer3_outputs(7627) <= a and not b;
    layer3_outputs(7628) <= a or b;
    layer3_outputs(7629) <= b and not a;
    layer3_outputs(7630) <= a and not b;
    layer3_outputs(7631) <= not (a xor b);
    layer3_outputs(7632) <= not (a and b);
    layer3_outputs(7633) <= a and b;
    layer3_outputs(7634) <= not b or a;
    layer3_outputs(7635) <= a or b;
    layer3_outputs(7636) <= '0';
    layer3_outputs(7637) <= not b;
    layer3_outputs(7638) <= '1';
    layer3_outputs(7639) <= '1';
    layer3_outputs(7640) <= '1';
    layer3_outputs(7641) <= a and not b;
    layer3_outputs(7642) <= a and not b;
    layer3_outputs(7643) <= a and b;
    layer3_outputs(7644) <= a or b;
    layer3_outputs(7645) <= not (a or b);
    layer3_outputs(7646) <= not (a or b);
    layer3_outputs(7647) <= a and b;
    layer3_outputs(7648) <= not a;
    layer3_outputs(7649) <= not (a or b);
    layer3_outputs(7650) <= not b;
    layer3_outputs(7651) <= not (a or b);
    layer3_outputs(7652) <= '0';
    layer3_outputs(7653) <= not b or a;
    layer3_outputs(7654) <= not (a or b);
    layer3_outputs(7655) <= not b or a;
    layer3_outputs(7656) <= not b;
    layer3_outputs(7657) <= '0';
    layer3_outputs(7658) <= not b or a;
    layer3_outputs(7659) <= not a;
    layer3_outputs(7660) <= a and not b;
    layer3_outputs(7661) <= '1';
    layer3_outputs(7662) <= not a or b;
    layer3_outputs(7663) <= b;
    layer3_outputs(7664) <= a and b;
    layer3_outputs(7665) <= b and not a;
    layer3_outputs(7666) <= not a;
    layer3_outputs(7667) <= not a or b;
    layer3_outputs(7668) <= not b;
    layer3_outputs(7669) <= '1';
    layer3_outputs(7670) <= '0';
    layer3_outputs(7671) <= not b or a;
    layer3_outputs(7672) <= a;
    layer3_outputs(7673) <= not (a and b);
    layer3_outputs(7674) <= a and b;
    layer3_outputs(7675) <= not (a or b);
    layer3_outputs(7676) <= a and not b;
    layer3_outputs(7677) <= b;
    layer3_outputs(7678) <= a or b;
    layer3_outputs(7679) <= not a or b;
    layer4_outputs(0) <= not a;
    layer4_outputs(1) <= not b;
    layer4_outputs(2) <= not (a or b);
    layer4_outputs(3) <= a and b;
    layer4_outputs(4) <= not b or a;
    layer4_outputs(5) <= a or b;
    layer4_outputs(6) <= b and not a;
    layer4_outputs(7) <= '0';
    layer4_outputs(8) <= not (a or b);
    layer4_outputs(9) <= a and not b;
    layer4_outputs(10) <= not b or a;
    layer4_outputs(11) <= a;
    layer4_outputs(12) <= a and not b;
    layer4_outputs(13) <= b;
    layer4_outputs(14) <= a and b;
    layer4_outputs(15) <= not a or b;
    layer4_outputs(16) <= not a or b;
    layer4_outputs(17) <= '1';
    layer4_outputs(18) <= not (a xor b);
    layer4_outputs(19) <= b and not a;
    layer4_outputs(20) <= not (a or b);
    layer4_outputs(21) <= not (a or b);
    layer4_outputs(22) <= not a;
    layer4_outputs(23) <= '1';
    layer4_outputs(24) <= '1';
    layer4_outputs(25) <= not a or b;
    layer4_outputs(26) <= a or b;
    layer4_outputs(27) <= not (a and b);
    layer4_outputs(28) <= not b or a;
    layer4_outputs(29) <= not b;
    layer4_outputs(30) <= a;
    layer4_outputs(31) <= '0';
    layer4_outputs(32) <= not a;
    layer4_outputs(33) <= not (a and b);
    layer4_outputs(34) <= a;
    layer4_outputs(35) <= not b or a;
    layer4_outputs(36) <= a or b;
    layer4_outputs(37) <= a or b;
    layer4_outputs(38) <= a xor b;
    layer4_outputs(39) <= not a;
    layer4_outputs(40) <= not (a xor b);
    layer4_outputs(41) <= not a or b;
    layer4_outputs(42) <= not (a and b);
    layer4_outputs(43) <= not a or b;
    layer4_outputs(44) <= '0';
    layer4_outputs(45) <= a;
    layer4_outputs(46) <= a and b;
    layer4_outputs(47) <= '1';
    layer4_outputs(48) <= '0';
    layer4_outputs(49) <= not b;
    layer4_outputs(50) <= a and not b;
    layer4_outputs(51) <= a and not b;
    layer4_outputs(52) <= not b;
    layer4_outputs(53) <= not b or a;
    layer4_outputs(54) <= b and not a;
    layer4_outputs(55) <= a and b;
    layer4_outputs(56) <= b and not a;
    layer4_outputs(57) <= a and not b;
    layer4_outputs(58) <= not a or b;
    layer4_outputs(59) <= not a;
    layer4_outputs(60) <= not (a or b);
    layer4_outputs(61) <= not (a and b);
    layer4_outputs(62) <= not b or a;
    layer4_outputs(63) <= not a or b;
    layer4_outputs(64) <= b;
    layer4_outputs(65) <= b and not a;
    layer4_outputs(66) <= '1';
    layer4_outputs(67) <= not b or a;
    layer4_outputs(68) <= b;
    layer4_outputs(69) <= not b;
    layer4_outputs(70) <= '1';
    layer4_outputs(71) <= a and not b;
    layer4_outputs(72) <= a;
    layer4_outputs(73) <= not (a or b);
    layer4_outputs(74) <= not (a and b);
    layer4_outputs(75) <= a and not b;
    layer4_outputs(76) <= a or b;
    layer4_outputs(77) <= b and not a;
    layer4_outputs(78) <= not (a or b);
    layer4_outputs(79) <= '0';
    layer4_outputs(80) <= a and b;
    layer4_outputs(81) <= a and b;
    layer4_outputs(82) <= '1';
    layer4_outputs(83) <= '1';
    layer4_outputs(84) <= not a or b;
    layer4_outputs(85) <= b;
    layer4_outputs(86) <= not a or b;
    layer4_outputs(87) <= a;
    layer4_outputs(88) <= a xor b;
    layer4_outputs(89) <= not (a and b);
    layer4_outputs(90) <= not b or a;
    layer4_outputs(91) <= '1';
    layer4_outputs(92) <= not a;
    layer4_outputs(93) <= b;
    layer4_outputs(94) <= a and not b;
    layer4_outputs(95) <= '1';
    layer4_outputs(96) <= not b;
    layer4_outputs(97) <= not a;
    layer4_outputs(98) <= not (a and b);
    layer4_outputs(99) <= not (a xor b);
    layer4_outputs(100) <= not (a and b);
    layer4_outputs(101) <= not a;
    layer4_outputs(102) <= a and b;
    layer4_outputs(103) <= a or b;
    layer4_outputs(104) <= not a;
    layer4_outputs(105) <= '0';
    layer4_outputs(106) <= a and not b;
    layer4_outputs(107) <= b;
    layer4_outputs(108) <= b;
    layer4_outputs(109) <= '0';
    layer4_outputs(110) <= '1';
    layer4_outputs(111) <= '1';
    layer4_outputs(112) <= a and not b;
    layer4_outputs(113) <= not b or a;
    layer4_outputs(114) <= a;
    layer4_outputs(115) <= not b or a;
    layer4_outputs(116) <= not (a and b);
    layer4_outputs(117) <= a;
    layer4_outputs(118) <= a and not b;
    layer4_outputs(119) <= b;
    layer4_outputs(120) <= '0';
    layer4_outputs(121) <= not a;
    layer4_outputs(122) <= not b;
    layer4_outputs(123) <= not (a or b);
    layer4_outputs(124) <= not a or b;
    layer4_outputs(125) <= not (a and b);
    layer4_outputs(126) <= a or b;
    layer4_outputs(127) <= not a;
    layer4_outputs(128) <= a or b;
    layer4_outputs(129) <= not (a or b);
    layer4_outputs(130) <= not (a or b);
    layer4_outputs(131) <= a and b;
    layer4_outputs(132) <= not a;
    layer4_outputs(133) <= '0';
    layer4_outputs(134) <= not a or b;
    layer4_outputs(135) <= b and not a;
    layer4_outputs(136) <= not (a and b);
    layer4_outputs(137) <= a;
    layer4_outputs(138) <= not b or a;
    layer4_outputs(139) <= b and not a;
    layer4_outputs(140) <= not a or b;
    layer4_outputs(141) <= b and not a;
    layer4_outputs(142) <= not (a and b);
    layer4_outputs(143) <= a and b;
    layer4_outputs(144) <= a;
    layer4_outputs(145) <= not a;
    layer4_outputs(146) <= a;
    layer4_outputs(147) <= a;
    layer4_outputs(148) <= a and b;
    layer4_outputs(149) <= a;
    layer4_outputs(150) <= b and not a;
    layer4_outputs(151) <= not a;
    layer4_outputs(152) <= b and not a;
    layer4_outputs(153) <= a;
    layer4_outputs(154) <= b and not a;
    layer4_outputs(155) <= a or b;
    layer4_outputs(156) <= a or b;
    layer4_outputs(157) <= a and not b;
    layer4_outputs(158) <= b;
    layer4_outputs(159) <= not (a and b);
    layer4_outputs(160) <= a or b;
    layer4_outputs(161) <= not b or a;
    layer4_outputs(162) <= '1';
    layer4_outputs(163) <= a;
    layer4_outputs(164) <= b and not a;
    layer4_outputs(165) <= not a;
    layer4_outputs(166) <= a;
    layer4_outputs(167) <= not (a or b);
    layer4_outputs(168) <= not (a xor b);
    layer4_outputs(169) <= a;
    layer4_outputs(170) <= '1';
    layer4_outputs(171) <= not (a or b);
    layer4_outputs(172) <= not a or b;
    layer4_outputs(173) <= b and not a;
    layer4_outputs(174) <= b and not a;
    layer4_outputs(175) <= b;
    layer4_outputs(176) <= not (a and b);
    layer4_outputs(177) <= a and not b;
    layer4_outputs(178) <= not (a or b);
    layer4_outputs(179) <= b and not a;
    layer4_outputs(180) <= b;
    layer4_outputs(181) <= not (a xor b);
    layer4_outputs(182) <= a and b;
    layer4_outputs(183) <= not a or b;
    layer4_outputs(184) <= b;
    layer4_outputs(185) <= '1';
    layer4_outputs(186) <= not (a xor b);
    layer4_outputs(187) <= a or b;
    layer4_outputs(188) <= not a;
    layer4_outputs(189) <= a;
    layer4_outputs(190) <= b and not a;
    layer4_outputs(191) <= not b;
    layer4_outputs(192) <= not b;
    layer4_outputs(193) <= not a or b;
    layer4_outputs(194) <= '0';
    layer4_outputs(195) <= '0';
    layer4_outputs(196) <= a and not b;
    layer4_outputs(197) <= not b or a;
    layer4_outputs(198) <= not a or b;
    layer4_outputs(199) <= '0';
    layer4_outputs(200) <= not b;
    layer4_outputs(201) <= not (a and b);
    layer4_outputs(202) <= '1';
    layer4_outputs(203) <= a or b;
    layer4_outputs(204) <= '1';
    layer4_outputs(205) <= a and b;
    layer4_outputs(206) <= not (a and b);
    layer4_outputs(207) <= not a;
    layer4_outputs(208) <= a and b;
    layer4_outputs(209) <= b;
    layer4_outputs(210) <= a and not b;
    layer4_outputs(211) <= '1';
    layer4_outputs(212) <= not a or b;
    layer4_outputs(213) <= a;
    layer4_outputs(214) <= a and not b;
    layer4_outputs(215) <= b;
    layer4_outputs(216) <= a or b;
    layer4_outputs(217) <= a;
    layer4_outputs(218) <= not a or b;
    layer4_outputs(219) <= a;
    layer4_outputs(220) <= a;
    layer4_outputs(221) <= a and not b;
    layer4_outputs(222) <= a or b;
    layer4_outputs(223) <= '0';
    layer4_outputs(224) <= '0';
    layer4_outputs(225) <= a or b;
    layer4_outputs(226) <= not (a and b);
    layer4_outputs(227) <= '1';
    layer4_outputs(228) <= a xor b;
    layer4_outputs(229) <= not a or b;
    layer4_outputs(230) <= not b or a;
    layer4_outputs(231) <= '1';
    layer4_outputs(232) <= not (a and b);
    layer4_outputs(233) <= a or b;
    layer4_outputs(234) <= a or b;
    layer4_outputs(235) <= a;
    layer4_outputs(236) <= a and b;
    layer4_outputs(237) <= not b;
    layer4_outputs(238) <= b and not a;
    layer4_outputs(239) <= a or b;
    layer4_outputs(240) <= a;
    layer4_outputs(241) <= a or b;
    layer4_outputs(242) <= not (a or b);
    layer4_outputs(243) <= not a or b;
    layer4_outputs(244) <= not a;
    layer4_outputs(245) <= not (a or b);
    layer4_outputs(246) <= '0';
    layer4_outputs(247) <= not (a and b);
    layer4_outputs(248) <= '1';
    layer4_outputs(249) <= a and not b;
    layer4_outputs(250) <= '0';
    layer4_outputs(251) <= not (a or b);
    layer4_outputs(252) <= '1';
    layer4_outputs(253) <= a and b;
    layer4_outputs(254) <= a xor b;
    layer4_outputs(255) <= not (a xor b);
    layer4_outputs(256) <= not b;
    layer4_outputs(257) <= not a;
    layer4_outputs(258) <= a and not b;
    layer4_outputs(259) <= not (a or b);
    layer4_outputs(260) <= a and b;
    layer4_outputs(261) <= not a;
    layer4_outputs(262) <= not a;
    layer4_outputs(263) <= a;
    layer4_outputs(264) <= not a or b;
    layer4_outputs(265) <= b;
    layer4_outputs(266) <= not (a or b);
    layer4_outputs(267) <= a and b;
    layer4_outputs(268) <= not a;
    layer4_outputs(269) <= a and not b;
    layer4_outputs(270) <= '1';
    layer4_outputs(271) <= not a;
    layer4_outputs(272) <= a;
    layer4_outputs(273) <= not b;
    layer4_outputs(274) <= b and not a;
    layer4_outputs(275) <= not (a and b);
    layer4_outputs(276) <= a or b;
    layer4_outputs(277) <= '0';
    layer4_outputs(278) <= not (a and b);
    layer4_outputs(279) <= b;
    layer4_outputs(280) <= b;
    layer4_outputs(281) <= not b or a;
    layer4_outputs(282) <= a and not b;
    layer4_outputs(283) <= not a;
    layer4_outputs(284) <= b and not a;
    layer4_outputs(285) <= a or b;
    layer4_outputs(286) <= a;
    layer4_outputs(287) <= a;
    layer4_outputs(288) <= not a or b;
    layer4_outputs(289) <= a;
    layer4_outputs(290) <= '1';
    layer4_outputs(291) <= not b;
    layer4_outputs(292) <= not a;
    layer4_outputs(293) <= not b or a;
    layer4_outputs(294) <= a and not b;
    layer4_outputs(295) <= a or b;
    layer4_outputs(296) <= not b;
    layer4_outputs(297) <= b and not a;
    layer4_outputs(298) <= a or b;
    layer4_outputs(299) <= '1';
    layer4_outputs(300) <= not (a or b);
    layer4_outputs(301) <= not (a xor b);
    layer4_outputs(302) <= '1';
    layer4_outputs(303) <= b;
    layer4_outputs(304) <= not a;
    layer4_outputs(305) <= not a;
    layer4_outputs(306) <= a and b;
    layer4_outputs(307) <= b and not a;
    layer4_outputs(308) <= a;
    layer4_outputs(309) <= b;
    layer4_outputs(310) <= not b;
    layer4_outputs(311) <= a and not b;
    layer4_outputs(312) <= not b or a;
    layer4_outputs(313) <= '1';
    layer4_outputs(314) <= b;
    layer4_outputs(315) <= '0';
    layer4_outputs(316) <= not a;
    layer4_outputs(317) <= not a or b;
    layer4_outputs(318) <= '1';
    layer4_outputs(319) <= a xor b;
    layer4_outputs(320) <= a or b;
    layer4_outputs(321) <= a or b;
    layer4_outputs(322) <= not (a or b);
    layer4_outputs(323) <= not (a and b);
    layer4_outputs(324) <= a;
    layer4_outputs(325) <= not (a and b);
    layer4_outputs(326) <= not b;
    layer4_outputs(327) <= a and b;
    layer4_outputs(328) <= a and not b;
    layer4_outputs(329) <= b and not a;
    layer4_outputs(330) <= not b;
    layer4_outputs(331) <= a and not b;
    layer4_outputs(332) <= not b;
    layer4_outputs(333) <= a and b;
    layer4_outputs(334) <= b and not a;
    layer4_outputs(335) <= not b or a;
    layer4_outputs(336) <= '1';
    layer4_outputs(337) <= not b;
    layer4_outputs(338) <= not b or a;
    layer4_outputs(339) <= a and not b;
    layer4_outputs(340) <= a or b;
    layer4_outputs(341) <= not b;
    layer4_outputs(342) <= not b;
    layer4_outputs(343) <= not a;
    layer4_outputs(344) <= not b;
    layer4_outputs(345) <= a and b;
    layer4_outputs(346) <= not (a and b);
    layer4_outputs(347) <= not a;
    layer4_outputs(348) <= b;
    layer4_outputs(349) <= not b or a;
    layer4_outputs(350) <= a and b;
    layer4_outputs(351) <= not a;
    layer4_outputs(352) <= a and not b;
    layer4_outputs(353) <= a;
    layer4_outputs(354) <= not a;
    layer4_outputs(355) <= '0';
    layer4_outputs(356) <= not (a xor b);
    layer4_outputs(357) <= b;
    layer4_outputs(358) <= a;
    layer4_outputs(359) <= not a or b;
    layer4_outputs(360) <= not a;
    layer4_outputs(361) <= not (a or b);
    layer4_outputs(362) <= not a or b;
    layer4_outputs(363) <= '0';
    layer4_outputs(364) <= a;
    layer4_outputs(365) <= not a;
    layer4_outputs(366) <= not a or b;
    layer4_outputs(367) <= not b;
    layer4_outputs(368) <= '1';
    layer4_outputs(369) <= b;
    layer4_outputs(370) <= not b or a;
    layer4_outputs(371) <= '0';
    layer4_outputs(372) <= b;
    layer4_outputs(373) <= not b or a;
    layer4_outputs(374) <= not b or a;
    layer4_outputs(375) <= not b;
    layer4_outputs(376) <= not (a or b);
    layer4_outputs(377) <= a and not b;
    layer4_outputs(378) <= a and b;
    layer4_outputs(379) <= '1';
    layer4_outputs(380) <= a and not b;
    layer4_outputs(381) <= not b or a;
    layer4_outputs(382) <= not a;
    layer4_outputs(383) <= a;
    layer4_outputs(384) <= not b;
    layer4_outputs(385) <= not b;
    layer4_outputs(386) <= a and not b;
    layer4_outputs(387) <= b and not a;
    layer4_outputs(388) <= not b or a;
    layer4_outputs(389) <= '0';
    layer4_outputs(390) <= a or b;
    layer4_outputs(391) <= not (a and b);
    layer4_outputs(392) <= not b or a;
    layer4_outputs(393) <= not (a xor b);
    layer4_outputs(394) <= b and not a;
    layer4_outputs(395) <= not b or a;
    layer4_outputs(396) <= not a or b;
    layer4_outputs(397) <= not b;
    layer4_outputs(398) <= not b;
    layer4_outputs(399) <= '0';
    layer4_outputs(400) <= b;
    layer4_outputs(401) <= a;
    layer4_outputs(402) <= a;
    layer4_outputs(403) <= a xor b;
    layer4_outputs(404) <= not b;
    layer4_outputs(405) <= a xor b;
    layer4_outputs(406) <= b;
    layer4_outputs(407) <= a;
    layer4_outputs(408) <= '1';
    layer4_outputs(409) <= a;
    layer4_outputs(410) <= b and not a;
    layer4_outputs(411) <= a and not b;
    layer4_outputs(412) <= not b;
    layer4_outputs(413) <= not b;
    layer4_outputs(414) <= not a or b;
    layer4_outputs(415) <= b;
    layer4_outputs(416) <= not (a and b);
    layer4_outputs(417) <= b;
    layer4_outputs(418) <= a and b;
    layer4_outputs(419) <= b;
    layer4_outputs(420) <= not (a and b);
    layer4_outputs(421) <= not b or a;
    layer4_outputs(422) <= '0';
    layer4_outputs(423) <= not a;
    layer4_outputs(424) <= a;
    layer4_outputs(425) <= a xor b;
    layer4_outputs(426) <= a xor b;
    layer4_outputs(427) <= '0';
    layer4_outputs(428) <= not (a or b);
    layer4_outputs(429) <= a and not b;
    layer4_outputs(430) <= not a or b;
    layer4_outputs(431) <= a and not b;
    layer4_outputs(432) <= not (a and b);
    layer4_outputs(433) <= '1';
    layer4_outputs(434) <= b and not a;
    layer4_outputs(435) <= a or b;
    layer4_outputs(436) <= a;
    layer4_outputs(437) <= not a or b;
    layer4_outputs(438) <= '0';
    layer4_outputs(439) <= '1';
    layer4_outputs(440) <= '0';
    layer4_outputs(441) <= '1';
    layer4_outputs(442) <= not (a and b);
    layer4_outputs(443) <= not b or a;
    layer4_outputs(444) <= not b;
    layer4_outputs(445) <= not (a or b);
    layer4_outputs(446) <= not a;
    layer4_outputs(447) <= not b;
    layer4_outputs(448) <= not a;
    layer4_outputs(449) <= a and b;
    layer4_outputs(450) <= not b or a;
    layer4_outputs(451) <= a;
    layer4_outputs(452) <= not b;
    layer4_outputs(453) <= not a or b;
    layer4_outputs(454) <= '1';
    layer4_outputs(455) <= a or b;
    layer4_outputs(456) <= b;
    layer4_outputs(457) <= not (a and b);
    layer4_outputs(458) <= not (a and b);
    layer4_outputs(459) <= not b or a;
    layer4_outputs(460) <= not b or a;
    layer4_outputs(461) <= '0';
    layer4_outputs(462) <= a;
    layer4_outputs(463) <= not b;
    layer4_outputs(464) <= not (a or b);
    layer4_outputs(465) <= a and not b;
    layer4_outputs(466) <= '0';
    layer4_outputs(467) <= '0';
    layer4_outputs(468) <= '1';
    layer4_outputs(469) <= not a or b;
    layer4_outputs(470) <= a;
    layer4_outputs(471) <= not (a and b);
    layer4_outputs(472) <= not b;
    layer4_outputs(473) <= a;
    layer4_outputs(474) <= not a or b;
    layer4_outputs(475) <= a xor b;
    layer4_outputs(476) <= not (a and b);
    layer4_outputs(477) <= not (a or b);
    layer4_outputs(478) <= not b;
    layer4_outputs(479) <= a;
    layer4_outputs(480) <= a and b;
    layer4_outputs(481) <= not (a or b);
    layer4_outputs(482) <= b and not a;
    layer4_outputs(483) <= not a;
    layer4_outputs(484) <= b and not a;
    layer4_outputs(485) <= a or b;
    layer4_outputs(486) <= not b;
    layer4_outputs(487) <= a or b;
    layer4_outputs(488) <= a and b;
    layer4_outputs(489) <= a and not b;
    layer4_outputs(490) <= b and not a;
    layer4_outputs(491) <= not b or a;
    layer4_outputs(492) <= '1';
    layer4_outputs(493) <= not (a and b);
    layer4_outputs(494) <= not b;
    layer4_outputs(495) <= not a;
    layer4_outputs(496) <= not (a and b);
    layer4_outputs(497) <= not b;
    layer4_outputs(498) <= not a;
    layer4_outputs(499) <= b;
    layer4_outputs(500) <= b;
    layer4_outputs(501) <= a and b;
    layer4_outputs(502) <= a xor b;
    layer4_outputs(503) <= a and not b;
    layer4_outputs(504) <= not a;
    layer4_outputs(505) <= a;
    layer4_outputs(506) <= b and not a;
    layer4_outputs(507) <= a and not b;
    layer4_outputs(508) <= not (a xor b);
    layer4_outputs(509) <= b and not a;
    layer4_outputs(510) <= b;
    layer4_outputs(511) <= a;
    layer4_outputs(512) <= b and not a;
    layer4_outputs(513) <= b;
    layer4_outputs(514) <= not a or b;
    layer4_outputs(515) <= a and b;
    layer4_outputs(516) <= a or b;
    layer4_outputs(517) <= b;
    layer4_outputs(518) <= '0';
    layer4_outputs(519) <= b and not a;
    layer4_outputs(520) <= '0';
    layer4_outputs(521) <= b and not a;
    layer4_outputs(522) <= not (a and b);
    layer4_outputs(523) <= not (a or b);
    layer4_outputs(524) <= a and b;
    layer4_outputs(525) <= not b or a;
    layer4_outputs(526) <= not (a xor b);
    layer4_outputs(527) <= not a;
    layer4_outputs(528) <= a and b;
    layer4_outputs(529) <= not b;
    layer4_outputs(530) <= a and b;
    layer4_outputs(531) <= not b or a;
    layer4_outputs(532) <= a;
    layer4_outputs(533) <= b;
    layer4_outputs(534) <= '0';
    layer4_outputs(535) <= '0';
    layer4_outputs(536) <= '1';
    layer4_outputs(537) <= a and not b;
    layer4_outputs(538) <= not b;
    layer4_outputs(539) <= a xor b;
    layer4_outputs(540) <= a;
    layer4_outputs(541) <= not b or a;
    layer4_outputs(542) <= not (a and b);
    layer4_outputs(543) <= a xor b;
    layer4_outputs(544) <= not b or a;
    layer4_outputs(545) <= not a;
    layer4_outputs(546) <= a xor b;
    layer4_outputs(547) <= b;
    layer4_outputs(548) <= a and b;
    layer4_outputs(549) <= a or b;
    layer4_outputs(550) <= a or b;
    layer4_outputs(551) <= a or b;
    layer4_outputs(552) <= not (a and b);
    layer4_outputs(553) <= not (a or b);
    layer4_outputs(554) <= a or b;
    layer4_outputs(555) <= '0';
    layer4_outputs(556) <= '0';
    layer4_outputs(557) <= not a or b;
    layer4_outputs(558) <= not b;
    layer4_outputs(559) <= a or b;
    layer4_outputs(560) <= a and not b;
    layer4_outputs(561) <= not a;
    layer4_outputs(562) <= a;
    layer4_outputs(563) <= a and b;
    layer4_outputs(564) <= '1';
    layer4_outputs(565) <= a;
    layer4_outputs(566) <= not (a or b);
    layer4_outputs(567) <= a and b;
    layer4_outputs(568) <= a and b;
    layer4_outputs(569) <= a;
    layer4_outputs(570) <= not (a and b);
    layer4_outputs(571) <= '0';
    layer4_outputs(572) <= '0';
    layer4_outputs(573) <= not (a or b);
    layer4_outputs(574) <= a and not b;
    layer4_outputs(575) <= not b;
    layer4_outputs(576) <= not b;
    layer4_outputs(577) <= not a or b;
    layer4_outputs(578) <= a and not b;
    layer4_outputs(579) <= a and not b;
    layer4_outputs(580) <= b and not a;
    layer4_outputs(581) <= not a;
    layer4_outputs(582) <= not (a or b);
    layer4_outputs(583) <= a and not b;
    layer4_outputs(584) <= not a or b;
    layer4_outputs(585) <= '1';
    layer4_outputs(586) <= '0';
    layer4_outputs(587) <= '1';
    layer4_outputs(588) <= a;
    layer4_outputs(589) <= a;
    layer4_outputs(590) <= b;
    layer4_outputs(591) <= '0';
    layer4_outputs(592) <= not b;
    layer4_outputs(593) <= a and b;
    layer4_outputs(594) <= a or b;
    layer4_outputs(595) <= not b;
    layer4_outputs(596) <= not b;
    layer4_outputs(597) <= not a or b;
    layer4_outputs(598) <= a;
    layer4_outputs(599) <= a and not b;
    layer4_outputs(600) <= not a or b;
    layer4_outputs(601) <= a and not b;
    layer4_outputs(602) <= not (a or b);
    layer4_outputs(603) <= a and not b;
    layer4_outputs(604) <= a and not b;
    layer4_outputs(605) <= not (a or b);
    layer4_outputs(606) <= not (a or b);
    layer4_outputs(607) <= '0';
    layer4_outputs(608) <= a and b;
    layer4_outputs(609) <= not b or a;
    layer4_outputs(610) <= b and not a;
    layer4_outputs(611) <= '1';
    layer4_outputs(612) <= not b;
    layer4_outputs(613) <= not b or a;
    layer4_outputs(614) <= a and not b;
    layer4_outputs(615) <= a or b;
    layer4_outputs(616) <= b;
    layer4_outputs(617) <= not a;
    layer4_outputs(618) <= '1';
    layer4_outputs(619) <= '1';
    layer4_outputs(620) <= not a;
    layer4_outputs(621) <= not a or b;
    layer4_outputs(622) <= not (a or b);
    layer4_outputs(623) <= '0';
    layer4_outputs(624) <= not a or b;
    layer4_outputs(625) <= a and b;
    layer4_outputs(626) <= not (a xor b);
    layer4_outputs(627) <= a or b;
    layer4_outputs(628) <= b and not a;
    layer4_outputs(629) <= a and b;
    layer4_outputs(630) <= a and b;
    layer4_outputs(631) <= b;
    layer4_outputs(632) <= '1';
    layer4_outputs(633) <= a;
    layer4_outputs(634) <= not (a and b);
    layer4_outputs(635) <= not (a xor b);
    layer4_outputs(636) <= b and not a;
    layer4_outputs(637) <= not (a or b);
    layer4_outputs(638) <= a and not b;
    layer4_outputs(639) <= b;
    layer4_outputs(640) <= a or b;
    layer4_outputs(641) <= a;
    layer4_outputs(642) <= a and not b;
    layer4_outputs(643) <= not b or a;
    layer4_outputs(644) <= a;
    layer4_outputs(645) <= b;
    layer4_outputs(646) <= '1';
    layer4_outputs(647) <= not a or b;
    layer4_outputs(648) <= '1';
    layer4_outputs(649) <= '1';
    layer4_outputs(650) <= b;
    layer4_outputs(651) <= not a;
    layer4_outputs(652) <= a;
    layer4_outputs(653) <= '0';
    layer4_outputs(654) <= a and b;
    layer4_outputs(655) <= b;
    layer4_outputs(656) <= a;
    layer4_outputs(657) <= b and not a;
    layer4_outputs(658) <= b;
    layer4_outputs(659) <= a and b;
    layer4_outputs(660) <= not (a xor b);
    layer4_outputs(661) <= b and not a;
    layer4_outputs(662) <= '1';
    layer4_outputs(663) <= not a;
    layer4_outputs(664) <= not (a or b);
    layer4_outputs(665) <= not b;
    layer4_outputs(666) <= not (a and b);
    layer4_outputs(667) <= a and b;
    layer4_outputs(668) <= not b or a;
    layer4_outputs(669) <= a and b;
    layer4_outputs(670) <= b and not a;
    layer4_outputs(671) <= a;
    layer4_outputs(672) <= a and b;
    layer4_outputs(673) <= a and b;
    layer4_outputs(674) <= a and not b;
    layer4_outputs(675) <= not b;
    layer4_outputs(676) <= not (a and b);
    layer4_outputs(677) <= not (a or b);
    layer4_outputs(678) <= not b;
    layer4_outputs(679) <= b and not a;
    layer4_outputs(680) <= not a or b;
    layer4_outputs(681) <= a and b;
    layer4_outputs(682) <= '1';
    layer4_outputs(683) <= b and not a;
    layer4_outputs(684) <= b;
    layer4_outputs(685) <= b;
    layer4_outputs(686) <= a and b;
    layer4_outputs(687) <= '1';
    layer4_outputs(688) <= not a;
    layer4_outputs(689) <= a and not b;
    layer4_outputs(690) <= b;
    layer4_outputs(691) <= b and not a;
    layer4_outputs(692) <= not a or b;
    layer4_outputs(693) <= not (a or b);
    layer4_outputs(694) <= a or b;
    layer4_outputs(695) <= not (a or b);
    layer4_outputs(696) <= a and not b;
    layer4_outputs(697) <= b and not a;
    layer4_outputs(698) <= not (a or b);
    layer4_outputs(699) <= a xor b;
    layer4_outputs(700) <= b;
    layer4_outputs(701) <= b and not a;
    layer4_outputs(702) <= '1';
    layer4_outputs(703) <= '1';
    layer4_outputs(704) <= not (a or b);
    layer4_outputs(705) <= a or b;
    layer4_outputs(706) <= not (a or b);
    layer4_outputs(707) <= not a;
    layer4_outputs(708) <= not b or a;
    layer4_outputs(709) <= a or b;
    layer4_outputs(710) <= not (a and b);
    layer4_outputs(711) <= not b;
    layer4_outputs(712) <= a and not b;
    layer4_outputs(713) <= a xor b;
    layer4_outputs(714) <= a and b;
    layer4_outputs(715) <= '0';
    layer4_outputs(716) <= a;
    layer4_outputs(717) <= not b or a;
    layer4_outputs(718) <= a and b;
    layer4_outputs(719) <= not a;
    layer4_outputs(720) <= not (a xor b);
    layer4_outputs(721) <= a xor b;
    layer4_outputs(722) <= not (a and b);
    layer4_outputs(723) <= not a;
    layer4_outputs(724) <= not b or a;
    layer4_outputs(725) <= '0';
    layer4_outputs(726) <= a or b;
    layer4_outputs(727) <= '0';
    layer4_outputs(728) <= not a;
    layer4_outputs(729) <= not (a and b);
    layer4_outputs(730) <= b and not a;
    layer4_outputs(731) <= not (a xor b);
    layer4_outputs(732) <= '0';
    layer4_outputs(733) <= '0';
    layer4_outputs(734) <= not a;
    layer4_outputs(735) <= b and not a;
    layer4_outputs(736) <= not b or a;
    layer4_outputs(737) <= not (a and b);
    layer4_outputs(738) <= not (a or b);
    layer4_outputs(739) <= a;
    layer4_outputs(740) <= b;
    layer4_outputs(741) <= a and not b;
    layer4_outputs(742) <= '0';
    layer4_outputs(743) <= not (a or b);
    layer4_outputs(744) <= a;
    layer4_outputs(745) <= not a;
    layer4_outputs(746) <= not (a and b);
    layer4_outputs(747) <= not (a or b);
    layer4_outputs(748) <= b and not a;
    layer4_outputs(749) <= a;
    layer4_outputs(750) <= b;
    layer4_outputs(751) <= '1';
    layer4_outputs(752) <= a or b;
    layer4_outputs(753) <= not (a and b);
    layer4_outputs(754) <= not b;
    layer4_outputs(755) <= '1';
    layer4_outputs(756) <= b;
    layer4_outputs(757) <= not b or a;
    layer4_outputs(758) <= not (a and b);
    layer4_outputs(759) <= a and not b;
    layer4_outputs(760) <= not (a xor b);
    layer4_outputs(761) <= b and not a;
    layer4_outputs(762) <= not (a and b);
    layer4_outputs(763) <= not (a xor b);
    layer4_outputs(764) <= not a or b;
    layer4_outputs(765) <= not b or a;
    layer4_outputs(766) <= not (a or b);
    layer4_outputs(767) <= a xor b;
    layer4_outputs(768) <= a and b;
    layer4_outputs(769) <= a or b;
    layer4_outputs(770) <= a and b;
    layer4_outputs(771) <= not (a and b);
    layer4_outputs(772) <= b;
    layer4_outputs(773) <= not a;
    layer4_outputs(774) <= '0';
    layer4_outputs(775) <= '0';
    layer4_outputs(776) <= a or b;
    layer4_outputs(777) <= not (a and b);
    layer4_outputs(778) <= a;
    layer4_outputs(779) <= not b;
    layer4_outputs(780) <= not b;
    layer4_outputs(781) <= b;
    layer4_outputs(782) <= not b or a;
    layer4_outputs(783) <= not (a or b);
    layer4_outputs(784) <= not a;
    layer4_outputs(785) <= b and not a;
    layer4_outputs(786) <= a or b;
    layer4_outputs(787) <= b and not a;
    layer4_outputs(788) <= a xor b;
    layer4_outputs(789) <= b;
    layer4_outputs(790) <= not a or b;
    layer4_outputs(791) <= not a;
    layer4_outputs(792) <= not b or a;
    layer4_outputs(793) <= not (a xor b);
    layer4_outputs(794) <= a and b;
    layer4_outputs(795) <= a and b;
    layer4_outputs(796) <= a and not b;
    layer4_outputs(797) <= a or b;
    layer4_outputs(798) <= b;
    layer4_outputs(799) <= not a or b;
    layer4_outputs(800) <= not a;
    layer4_outputs(801) <= b;
    layer4_outputs(802) <= a or b;
    layer4_outputs(803) <= not b or a;
    layer4_outputs(804) <= not b;
    layer4_outputs(805) <= not b;
    layer4_outputs(806) <= a and not b;
    layer4_outputs(807) <= not (a xor b);
    layer4_outputs(808) <= not a;
    layer4_outputs(809) <= not (a and b);
    layer4_outputs(810) <= a and not b;
    layer4_outputs(811) <= not b or a;
    layer4_outputs(812) <= a and b;
    layer4_outputs(813) <= a and b;
    layer4_outputs(814) <= a and not b;
    layer4_outputs(815) <= not b;
    layer4_outputs(816) <= a or b;
    layer4_outputs(817) <= not (a and b);
    layer4_outputs(818) <= not (a or b);
    layer4_outputs(819) <= not a;
    layer4_outputs(820) <= not a;
    layer4_outputs(821) <= not b;
    layer4_outputs(822) <= '1';
    layer4_outputs(823) <= b and not a;
    layer4_outputs(824) <= b;
    layer4_outputs(825) <= a;
    layer4_outputs(826) <= not (a and b);
    layer4_outputs(827) <= a;
    layer4_outputs(828) <= not b;
    layer4_outputs(829) <= '1';
    layer4_outputs(830) <= not b;
    layer4_outputs(831) <= a or b;
    layer4_outputs(832) <= a and not b;
    layer4_outputs(833) <= not b;
    layer4_outputs(834) <= a and not b;
    layer4_outputs(835) <= b and not a;
    layer4_outputs(836) <= b and not a;
    layer4_outputs(837) <= a and not b;
    layer4_outputs(838) <= not b;
    layer4_outputs(839) <= a and b;
    layer4_outputs(840) <= not b or a;
    layer4_outputs(841) <= not b or a;
    layer4_outputs(842) <= a or b;
    layer4_outputs(843) <= not (a or b);
    layer4_outputs(844) <= b and not a;
    layer4_outputs(845) <= a and not b;
    layer4_outputs(846) <= '0';
    layer4_outputs(847) <= not b or a;
    layer4_outputs(848) <= not (a and b);
    layer4_outputs(849) <= a and not b;
    layer4_outputs(850) <= b;
    layer4_outputs(851) <= not (a or b);
    layer4_outputs(852) <= a;
    layer4_outputs(853) <= not (a or b);
    layer4_outputs(854) <= not (a or b);
    layer4_outputs(855) <= '1';
    layer4_outputs(856) <= b;
    layer4_outputs(857) <= '0';
    layer4_outputs(858) <= a;
    layer4_outputs(859) <= '0';
    layer4_outputs(860) <= b and not a;
    layer4_outputs(861) <= a or b;
    layer4_outputs(862) <= a or b;
    layer4_outputs(863) <= a;
    layer4_outputs(864) <= a and not b;
    layer4_outputs(865) <= '1';
    layer4_outputs(866) <= not (a or b);
    layer4_outputs(867) <= a or b;
    layer4_outputs(868) <= b;
    layer4_outputs(869) <= a or b;
    layer4_outputs(870) <= a and b;
    layer4_outputs(871) <= b and not a;
    layer4_outputs(872) <= b and not a;
    layer4_outputs(873) <= b;
    layer4_outputs(874) <= b;
    layer4_outputs(875) <= b;
    layer4_outputs(876) <= a xor b;
    layer4_outputs(877) <= not (a or b);
    layer4_outputs(878) <= '1';
    layer4_outputs(879) <= not a or b;
    layer4_outputs(880) <= '0';
    layer4_outputs(881) <= a and not b;
    layer4_outputs(882) <= not b or a;
    layer4_outputs(883) <= a or b;
    layer4_outputs(884) <= not b;
    layer4_outputs(885) <= a and b;
    layer4_outputs(886) <= '1';
    layer4_outputs(887) <= b;
    layer4_outputs(888) <= a xor b;
    layer4_outputs(889) <= not b or a;
    layer4_outputs(890) <= b;
    layer4_outputs(891) <= not (a and b);
    layer4_outputs(892) <= a or b;
    layer4_outputs(893) <= not b;
    layer4_outputs(894) <= a and not b;
    layer4_outputs(895) <= a and not b;
    layer4_outputs(896) <= a or b;
    layer4_outputs(897) <= b;
    layer4_outputs(898) <= not b or a;
    layer4_outputs(899) <= '0';
    layer4_outputs(900) <= a;
    layer4_outputs(901) <= '0';
    layer4_outputs(902) <= not b;
    layer4_outputs(903) <= a;
    layer4_outputs(904) <= not (a or b);
    layer4_outputs(905) <= '0';
    layer4_outputs(906) <= b;
    layer4_outputs(907) <= not a;
    layer4_outputs(908) <= not b or a;
    layer4_outputs(909) <= a and not b;
    layer4_outputs(910) <= a and b;
    layer4_outputs(911) <= not a;
    layer4_outputs(912) <= not a or b;
    layer4_outputs(913) <= b;
    layer4_outputs(914) <= not (a xor b);
    layer4_outputs(915) <= a or b;
    layer4_outputs(916) <= a and not b;
    layer4_outputs(917) <= '0';
    layer4_outputs(918) <= b and not a;
    layer4_outputs(919) <= not b;
    layer4_outputs(920) <= '1';
    layer4_outputs(921) <= not a or b;
    layer4_outputs(922) <= a and b;
    layer4_outputs(923) <= not a;
    layer4_outputs(924) <= not a;
    layer4_outputs(925) <= not b;
    layer4_outputs(926) <= '1';
    layer4_outputs(927) <= not b;
    layer4_outputs(928) <= '1';
    layer4_outputs(929) <= a;
    layer4_outputs(930) <= not a or b;
    layer4_outputs(931) <= not a;
    layer4_outputs(932) <= a or b;
    layer4_outputs(933) <= not (a and b);
    layer4_outputs(934) <= a and b;
    layer4_outputs(935) <= '1';
    layer4_outputs(936) <= not (a and b);
    layer4_outputs(937) <= b and not a;
    layer4_outputs(938) <= not a;
    layer4_outputs(939) <= not (a or b);
    layer4_outputs(940) <= a;
    layer4_outputs(941) <= a or b;
    layer4_outputs(942) <= not (a xor b);
    layer4_outputs(943) <= not b or a;
    layer4_outputs(944) <= a and b;
    layer4_outputs(945) <= '0';
    layer4_outputs(946) <= not a or b;
    layer4_outputs(947) <= not b;
    layer4_outputs(948) <= not a;
    layer4_outputs(949) <= not b or a;
    layer4_outputs(950) <= a;
    layer4_outputs(951) <= not (a xor b);
    layer4_outputs(952) <= '0';
    layer4_outputs(953) <= b and not a;
    layer4_outputs(954) <= not (a and b);
    layer4_outputs(955) <= a xor b;
    layer4_outputs(956) <= not b or a;
    layer4_outputs(957) <= not (a and b);
    layer4_outputs(958) <= not b;
    layer4_outputs(959) <= a xor b;
    layer4_outputs(960) <= a xor b;
    layer4_outputs(961) <= a or b;
    layer4_outputs(962) <= b and not a;
    layer4_outputs(963) <= a xor b;
    layer4_outputs(964) <= a and not b;
    layer4_outputs(965) <= not a or b;
    layer4_outputs(966) <= b;
    layer4_outputs(967) <= a;
    layer4_outputs(968) <= not (a or b);
    layer4_outputs(969) <= not b or a;
    layer4_outputs(970) <= a xor b;
    layer4_outputs(971) <= not a;
    layer4_outputs(972) <= b;
    layer4_outputs(973) <= '1';
    layer4_outputs(974) <= a and b;
    layer4_outputs(975) <= not a;
    layer4_outputs(976) <= not a or b;
    layer4_outputs(977) <= a or b;
    layer4_outputs(978) <= not (a and b);
    layer4_outputs(979) <= a;
    layer4_outputs(980) <= not (a or b);
    layer4_outputs(981) <= b;
    layer4_outputs(982) <= a;
    layer4_outputs(983) <= a;
    layer4_outputs(984) <= not a or b;
    layer4_outputs(985) <= b and not a;
    layer4_outputs(986) <= not b;
    layer4_outputs(987) <= a;
    layer4_outputs(988) <= not a;
    layer4_outputs(989) <= not b or a;
    layer4_outputs(990) <= not (a or b);
    layer4_outputs(991) <= not a;
    layer4_outputs(992) <= not a or b;
    layer4_outputs(993) <= a and b;
    layer4_outputs(994) <= not a or b;
    layer4_outputs(995) <= a or b;
    layer4_outputs(996) <= b;
    layer4_outputs(997) <= '1';
    layer4_outputs(998) <= a and b;
    layer4_outputs(999) <= not a;
    layer4_outputs(1000) <= a or b;
    layer4_outputs(1001) <= not b;
    layer4_outputs(1002) <= not a;
    layer4_outputs(1003) <= a;
    layer4_outputs(1004) <= b and not a;
    layer4_outputs(1005) <= not (a or b);
    layer4_outputs(1006) <= not (a and b);
    layer4_outputs(1007) <= not a;
    layer4_outputs(1008) <= a or b;
    layer4_outputs(1009) <= not b or a;
    layer4_outputs(1010) <= b;
    layer4_outputs(1011) <= '1';
    layer4_outputs(1012) <= not (a or b);
    layer4_outputs(1013) <= a and not b;
    layer4_outputs(1014) <= not (a xor b);
    layer4_outputs(1015) <= not (a and b);
    layer4_outputs(1016) <= a or b;
    layer4_outputs(1017) <= b;
    layer4_outputs(1018) <= not a;
    layer4_outputs(1019) <= not (a xor b);
    layer4_outputs(1020) <= not (a or b);
    layer4_outputs(1021) <= not a or b;
    layer4_outputs(1022) <= not (a and b);
    layer4_outputs(1023) <= a or b;
    layer4_outputs(1024) <= not b;
    layer4_outputs(1025) <= '1';
    layer4_outputs(1026) <= not (a and b);
    layer4_outputs(1027) <= not b;
    layer4_outputs(1028) <= a;
    layer4_outputs(1029) <= b;
    layer4_outputs(1030) <= b;
    layer4_outputs(1031) <= not b or a;
    layer4_outputs(1032) <= b;
    layer4_outputs(1033) <= a and b;
    layer4_outputs(1034) <= '0';
    layer4_outputs(1035) <= a and not b;
    layer4_outputs(1036) <= not b or a;
    layer4_outputs(1037) <= not a or b;
    layer4_outputs(1038) <= a and b;
    layer4_outputs(1039) <= not b or a;
    layer4_outputs(1040) <= not b or a;
    layer4_outputs(1041) <= not a;
    layer4_outputs(1042) <= a or b;
    layer4_outputs(1043) <= b and not a;
    layer4_outputs(1044) <= not b or a;
    layer4_outputs(1045) <= a;
    layer4_outputs(1046) <= not (a or b);
    layer4_outputs(1047) <= a and not b;
    layer4_outputs(1048) <= a and not b;
    layer4_outputs(1049) <= a;
    layer4_outputs(1050) <= not (a and b);
    layer4_outputs(1051) <= not (a and b);
    layer4_outputs(1052) <= '0';
    layer4_outputs(1053) <= a and not b;
    layer4_outputs(1054) <= a or b;
    layer4_outputs(1055) <= a or b;
    layer4_outputs(1056) <= not b;
    layer4_outputs(1057) <= not b;
    layer4_outputs(1058) <= not a;
    layer4_outputs(1059) <= a and not b;
    layer4_outputs(1060) <= b and not a;
    layer4_outputs(1061) <= b;
    layer4_outputs(1062) <= a and b;
    layer4_outputs(1063) <= not (a and b);
    layer4_outputs(1064) <= a or b;
    layer4_outputs(1065) <= a or b;
    layer4_outputs(1066) <= not (a and b);
    layer4_outputs(1067) <= a or b;
    layer4_outputs(1068) <= b;
    layer4_outputs(1069) <= b;
    layer4_outputs(1070) <= a;
    layer4_outputs(1071) <= not (a or b);
    layer4_outputs(1072) <= not (a and b);
    layer4_outputs(1073) <= not (a and b);
    layer4_outputs(1074) <= not a or b;
    layer4_outputs(1075) <= a and b;
    layer4_outputs(1076) <= not b or a;
    layer4_outputs(1077) <= a or b;
    layer4_outputs(1078) <= '1';
    layer4_outputs(1079) <= not a;
    layer4_outputs(1080) <= a or b;
    layer4_outputs(1081) <= not (a or b);
    layer4_outputs(1082) <= '1';
    layer4_outputs(1083) <= a xor b;
    layer4_outputs(1084) <= not b;
    layer4_outputs(1085) <= a and b;
    layer4_outputs(1086) <= not b or a;
    layer4_outputs(1087) <= a or b;
    layer4_outputs(1088) <= not (a and b);
    layer4_outputs(1089) <= not a;
    layer4_outputs(1090) <= not (a or b);
    layer4_outputs(1091) <= a or b;
    layer4_outputs(1092) <= a and not b;
    layer4_outputs(1093) <= a or b;
    layer4_outputs(1094) <= not a or b;
    layer4_outputs(1095) <= a;
    layer4_outputs(1096) <= a or b;
    layer4_outputs(1097) <= not (a and b);
    layer4_outputs(1098) <= not a;
    layer4_outputs(1099) <= not a or b;
    layer4_outputs(1100) <= not (a and b);
    layer4_outputs(1101) <= '1';
    layer4_outputs(1102) <= '0';
    layer4_outputs(1103) <= a xor b;
    layer4_outputs(1104) <= '0';
    layer4_outputs(1105) <= '0';
    layer4_outputs(1106) <= a;
    layer4_outputs(1107) <= not b or a;
    layer4_outputs(1108) <= b and not a;
    layer4_outputs(1109) <= a;
    layer4_outputs(1110) <= not a or b;
    layer4_outputs(1111) <= not a or b;
    layer4_outputs(1112) <= not (a and b);
    layer4_outputs(1113) <= a and not b;
    layer4_outputs(1114) <= '1';
    layer4_outputs(1115) <= a and not b;
    layer4_outputs(1116) <= a xor b;
    layer4_outputs(1117) <= a or b;
    layer4_outputs(1118) <= not b or a;
    layer4_outputs(1119) <= b;
    layer4_outputs(1120) <= not (a or b);
    layer4_outputs(1121) <= '1';
    layer4_outputs(1122) <= b and not a;
    layer4_outputs(1123) <= a;
    layer4_outputs(1124) <= not a or b;
    layer4_outputs(1125) <= b and not a;
    layer4_outputs(1126) <= not b or a;
    layer4_outputs(1127) <= a and not b;
    layer4_outputs(1128) <= not a or b;
    layer4_outputs(1129) <= b;
    layer4_outputs(1130) <= not b;
    layer4_outputs(1131) <= a and not b;
    layer4_outputs(1132) <= not a;
    layer4_outputs(1133) <= a and b;
    layer4_outputs(1134) <= b and not a;
    layer4_outputs(1135) <= not b or a;
    layer4_outputs(1136) <= '0';
    layer4_outputs(1137) <= a or b;
    layer4_outputs(1138) <= not b or a;
    layer4_outputs(1139) <= not b;
    layer4_outputs(1140) <= '1';
    layer4_outputs(1141) <= a and b;
    layer4_outputs(1142) <= not (a and b);
    layer4_outputs(1143) <= not (a or b);
    layer4_outputs(1144) <= a or b;
    layer4_outputs(1145) <= not a;
    layer4_outputs(1146) <= '0';
    layer4_outputs(1147) <= not (a and b);
    layer4_outputs(1148) <= not a or b;
    layer4_outputs(1149) <= a;
    layer4_outputs(1150) <= b and not a;
    layer4_outputs(1151) <= a;
    layer4_outputs(1152) <= not a;
    layer4_outputs(1153) <= b and not a;
    layer4_outputs(1154) <= b and not a;
    layer4_outputs(1155) <= '1';
    layer4_outputs(1156) <= not a;
    layer4_outputs(1157) <= not (a or b);
    layer4_outputs(1158) <= not b;
    layer4_outputs(1159) <= '1';
    layer4_outputs(1160) <= not b;
    layer4_outputs(1161) <= a and b;
    layer4_outputs(1162) <= b;
    layer4_outputs(1163) <= a or b;
    layer4_outputs(1164) <= not (a and b);
    layer4_outputs(1165) <= b;
    layer4_outputs(1166) <= b and not a;
    layer4_outputs(1167) <= b;
    layer4_outputs(1168) <= not (a and b);
    layer4_outputs(1169) <= a;
    layer4_outputs(1170) <= '0';
    layer4_outputs(1171) <= a;
    layer4_outputs(1172) <= not (a or b);
    layer4_outputs(1173) <= not (a or b);
    layer4_outputs(1174) <= a or b;
    layer4_outputs(1175) <= a and not b;
    layer4_outputs(1176) <= not b;
    layer4_outputs(1177) <= b and not a;
    layer4_outputs(1178) <= b;
    layer4_outputs(1179) <= not (a and b);
    layer4_outputs(1180) <= a or b;
    layer4_outputs(1181) <= a and not b;
    layer4_outputs(1182) <= b;
    layer4_outputs(1183) <= not (a xor b);
    layer4_outputs(1184) <= not (a xor b);
    layer4_outputs(1185) <= a and b;
    layer4_outputs(1186) <= not b or a;
    layer4_outputs(1187) <= not b;
    layer4_outputs(1188) <= b and not a;
    layer4_outputs(1189) <= not b;
    layer4_outputs(1190) <= a and b;
    layer4_outputs(1191) <= a or b;
    layer4_outputs(1192) <= not a;
    layer4_outputs(1193) <= not (a or b);
    layer4_outputs(1194) <= b;
    layer4_outputs(1195) <= a and b;
    layer4_outputs(1196) <= not (a or b);
    layer4_outputs(1197) <= a and b;
    layer4_outputs(1198) <= not a or b;
    layer4_outputs(1199) <= '0';
    layer4_outputs(1200) <= not (a xor b);
    layer4_outputs(1201) <= b and not a;
    layer4_outputs(1202) <= a or b;
    layer4_outputs(1203) <= a;
    layer4_outputs(1204) <= '1';
    layer4_outputs(1205) <= not b;
    layer4_outputs(1206) <= b;
    layer4_outputs(1207) <= b and not a;
    layer4_outputs(1208) <= not a or b;
    layer4_outputs(1209) <= b and not a;
    layer4_outputs(1210) <= not b or a;
    layer4_outputs(1211) <= a and b;
    layer4_outputs(1212) <= not (a and b);
    layer4_outputs(1213) <= a and not b;
    layer4_outputs(1214) <= not (a and b);
    layer4_outputs(1215) <= not a;
    layer4_outputs(1216) <= a and not b;
    layer4_outputs(1217) <= a or b;
    layer4_outputs(1218) <= '1';
    layer4_outputs(1219) <= not b or a;
    layer4_outputs(1220) <= not (a and b);
    layer4_outputs(1221) <= a;
    layer4_outputs(1222) <= a and not b;
    layer4_outputs(1223) <= b and not a;
    layer4_outputs(1224) <= b;
    layer4_outputs(1225) <= not a or b;
    layer4_outputs(1226) <= not a or b;
    layer4_outputs(1227) <= not b or a;
    layer4_outputs(1228) <= not (a xor b);
    layer4_outputs(1229) <= not b;
    layer4_outputs(1230) <= a or b;
    layer4_outputs(1231) <= a xor b;
    layer4_outputs(1232) <= a or b;
    layer4_outputs(1233) <= not a or b;
    layer4_outputs(1234) <= a and b;
    layer4_outputs(1235) <= '1';
    layer4_outputs(1236) <= b;
    layer4_outputs(1237) <= '1';
    layer4_outputs(1238) <= not b;
    layer4_outputs(1239) <= '1';
    layer4_outputs(1240) <= b;
    layer4_outputs(1241) <= a;
    layer4_outputs(1242) <= not a or b;
    layer4_outputs(1243) <= '1';
    layer4_outputs(1244) <= a or b;
    layer4_outputs(1245) <= not b;
    layer4_outputs(1246) <= a or b;
    layer4_outputs(1247) <= b and not a;
    layer4_outputs(1248) <= a;
    layer4_outputs(1249) <= b and not a;
    layer4_outputs(1250) <= a;
    layer4_outputs(1251) <= not (a xor b);
    layer4_outputs(1252) <= not b;
    layer4_outputs(1253) <= a;
    layer4_outputs(1254) <= not a;
    layer4_outputs(1255) <= b;
    layer4_outputs(1256) <= not b;
    layer4_outputs(1257) <= b;
    layer4_outputs(1258) <= b;
    layer4_outputs(1259) <= not (a and b);
    layer4_outputs(1260) <= a;
    layer4_outputs(1261) <= a and b;
    layer4_outputs(1262) <= b;
    layer4_outputs(1263) <= a and not b;
    layer4_outputs(1264) <= a;
    layer4_outputs(1265) <= not a or b;
    layer4_outputs(1266) <= a and b;
    layer4_outputs(1267) <= not a;
    layer4_outputs(1268) <= not a;
    layer4_outputs(1269) <= not a or b;
    layer4_outputs(1270) <= not (a or b);
    layer4_outputs(1271) <= not (a and b);
    layer4_outputs(1272) <= '1';
    layer4_outputs(1273) <= not (a and b);
    layer4_outputs(1274) <= not a or b;
    layer4_outputs(1275) <= '1';
    layer4_outputs(1276) <= not (a and b);
    layer4_outputs(1277) <= not a;
    layer4_outputs(1278) <= a;
    layer4_outputs(1279) <= not b or a;
    layer4_outputs(1280) <= not b or a;
    layer4_outputs(1281) <= not b or a;
    layer4_outputs(1282) <= not (a or b);
    layer4_outputs(1283) <= not (a xor b);
    layer4_outputs(1284) <= not a or b;
    layer4_outputs(1285) <= '0';
    layer4_outputs(1286) <= a;
    layer4_outputs(1287) <= '1';
    layer4_outputs(1288) <= not (a or b);
    layer4_outputs(1289) <= a and not b;
    layer4_outputs(1290) <= not (a and b);
    layer4_outputs(1291) <= a;
    layer4_outputs(1292) <= not (a and b);
    layer4_outputs(1293) <= a or b;
    layer4_outputs(1294) <= not a;
    layer4_outputs(1295) <= not a;
    layer4_outputs(1296) <= a and not b;
    layer4_outputs(1297) <= a;
    layer4_outputs(1298) <= a and b;
    layer4_outputs(1299) <= not (a or b);
    layer4_outputs(1300) <= a or b;
    layer4_outputs(1301) <= not a;
    layer4_outputs(1302) <= a xor b;
    layer4_outputs(1303) <= b and not a;
    layer4_outputs(1304) <= not (a and b);
    layer4_outputs(1305) <= a xor b;
    layer4_outputs(1306) <= a and b;
    layer4_outputs(1307) <= not b or a;
    layer4_outputs(1308) <= a and b;
    layer4_outputs(1309) <= not (a or b);
    layer4_outputs(1310) <= a and not b;
    layer4_outputs(1311) <= not (a and b);
    layer4_outputs(1312) <= '0';
    layer4_outputs(1313) <= a and b;
    layer4_outputs(1314) <= not b or a;
    layer4_outputs(1315) <= not a;
    layer4_outputs(1316) <= not b or a;
    layer4_outputs(1317) <= not (a and b);
    layer4_outputs(1318) <= '1';
    layer4_outputs(1319) <= a and not b;
    layer4_outputs(1320) <= not a;
    layer4_outputs(1321) <= '0';
    layer4_outputs(1322) <= not b or a;
    layer4_outputs(1323) <= '0';
    layer4_outputs(1324) <= b;
    layer4_outputs(1325) <= '1';
    layer4_outputs(1326) <= a or b;
    layer4_outputs(1327) <= a and not b;
    layer4_outputs(1328) <= not (a and b);
    layer4_outputs(1329) <= a;
    layer4_outputs(1330) <= not (a xor b);
    layer4_outputs(1331) <= '1';
    layer4_outputs(1332) <= not b;
    layer4_outputs(1333) <= b;
    layer4_outputs(1334) <= not (a and b);
    layer4_outputs(1335) <= not b;
    layer4_outputs(1336) <= not b or a;
    layer4_outputs(1337) <= not b;
    layer4_outputs(1338) <= b and not a;
    layer4_outputs(1339) <= not a;
    layer4_outputs(1340) <= not a;
    layer4_outputs(1341) <= a or b;
    layer4_outputs(1342) <= a;
    layer4_outputs(1343) <= a;
    layer4_outputs(1344) <= a;
    layer4_outputs(1345) <= not a or b;
    layer4_outputs(1346) <= a;
    layer4_outputs(1347) <= a and not b;
    layer4_outputs(1348) <= not (a and b);
    layer4_outputs(1349) <= a;
    layer4_outputs(1350) <= not (a and b);
    layer4_outputs(1351) <= not b;
    layer4_outputs(1352) <= a;
    layer4_outputs(1353) <= b;
    layer4_outputs(1354) <= b;
    layer4_outputs(1355) <= b;
    layer4_outputs(1356) <= '0';
    layer4_outputs(1357) <= a;
    layer4_outputs(1358) <= not b or a;
    layer4_outputs(1359) <= a or b;
    layer4_outputs(1360) <= a;
    layer4_outputs(1361) <= a and b;
    layer4_outputs(1362) <= not a;
    layer4_outputs(1363) <= not b;
    layer4_outputs(1364) <= not b;
    layer4_outputs(1365) <= not b;
    layer4_outputs(1366) <= a and b;
    layer4_outputs(1367) <= a;
    layer4_outputs(1368) <= '1';
    layer4_outputs(1369) <= a and not b;
    layer4_outputs(1370) <= '0';
    layer4_outputs(1371) <= b;
    layer4_outputs(1372) <= not (a xor b);
    layer4_outputs(1373) <= a or b;
    layer4_outputs(1374) <= not (a or b);
    layer4_outputs(1375) <= '0';
    layer4_outputs(1376) <= a or b;
    layer4_outputs(1377) <= not b or a;
    layer4_outputs(1378) <= not b;
    layer4_outputs(1379) <= not (a or b);
    layer4_outputs(1380) <= b;
    layer4_outputs(1381) <= not a or b;
    layer4_outputs(1382) <= a;
    layer4_outputs(1383) <= not b;
    layer4_outputs(1384) <= b;
    layer4_outputs(1385) <= not b;
    layer4_outputs(1386) <= not (a or b);
    layer4_outputs(1387) <= not b or a;
    layer4_outputs(1388) <= not a or b;
    layer4_outputs(1389) <= a and b;
    layer4_outputs(1390) <= not a;
    layer4_outputs(1391) <= not (a or b);
    layer4_outputs(1392) <= not (a and b);
    layer4_outputs(1393) <= not a or b;
    layer4_outputs(1394) <= not a;
    layer4_outputs(1395) <= a;
    layer4_outputs(1396) <= '1';
    layer4_outputs(1397) <= b and not a;
    layer4_outputs(1398) <= not b;
    layer4_outputs(1399) <= a;
    layer4_outputs(1400) <= a;
    layer4_outputs(1401) <= not b or a;
    layer4_outputs(1402) <= not b;
    layer4_outputs(1403) <= not a;
    layer4_outputs(1404) <= not (a xor b);
    layer4_outputs(1405) <= '1';
    layer4_outputs(1406) <= a and not b;
    layer4_outputs(1407) <= not (a and b);
    layer4_outputs(1408) <= not a or b;
    layer4_outputs(1409) <= a;
    layer4_outputs(1410) <= '1';
    layer4_outputs(1411) <= not (a or b);
    layer4_outputs(1412) <= not (a and b);
    layer4_outputs(1413) <= not (a or b);
    layer4_outputs(1414) <= not b or a;
    layer4_outputs(1415) <= not b;
    layer4_outputs(1416) <= not b or a;
    layer4_outputs(1417) <= a;
    layer4_outputs(1418) <= not b;
    layer4_outputs(1419) <= b;
    layer4_outputs(1420) <= not a or b;
    layer4_outputs(1421) <= a xor b;
    layer4_outputs(1422) <= not (a or b);
    layer4_outputs(1423) <= b;
    layer4_outputs(1424) <= not b or a;
    layer4_outputs(1425) <= not (a or b);
    layer4_outputs(1426) <= a and b;
    layer4_outputs(1427) <= not a or b;
    layer4_outputs(1428) <= not a or b;
    layer4_outputs(1429) <= b and not a;
    layer4_outputs(1430) <= a and not b;
    layer4_outputs(1431) <= a and not b;
    layer4_outputs(1432) <= not a;
    layer4_outputs(1433) <= a and not b;
    layer4_outputs(1434) <= not (a or b);
    layer4_outputs(1435) <= '0';
    layer4_outputs(1436) <= not b;
    layer4_outputs(1437) <= not b;
    layer4_outputs(1438) <= b and not a;
    layer4_outputs(1439) <= not (a and b);
    layer4_outputs(1440) <= not b or a;
    layer4_outputs(1441) <= not a;
    layer4_outputs(1442) <= a or b;
    layer4_outputs(1443) <= not b;
    layer4_outputs(1444) <= b;
    layer4_outputs(1445) <= not a;
    layer4_outputs(1446) <= '0';
    layer4_outputs(1447) <= not b;
    layer4_outputs(1448) <= a;
    layer4_outputs(1449) <= not b or a;
    layer4_outputs(1450) <= '0';
    layer4_outputs(1451) <= a or b;
    layer4_outputs(1452) <= a or b;
    layer4_outputs(1453) <= not a;
    layer4_outputs(1454) <= not a or b;
    layer4_outputs(1455) <= not a;
    layer4_outputs(1456) <= not b;
    layer4_outputs(1457) <= not b;
    layer4_outputs(1458) <= not a or b;
    layer4_outputs(1459) <= not a or b;
    layer4_outputs(1460) <= b;
    layer4_outputs(1461) <= not b;
    layer4_outputs(1462) <= a and not b;
    layer4_outputs(1463) <= not a or b;
    layer4_outputs(1464) <= a or b;
    layer4_outputs(1465) <= not (a or b);
    layer4_outputs(1466) <= not b;
    layer4_outputs(1467) <= b and not a;
    layer4_outputs(1468) <= b;
    layer4_outputs(1469) <= a or b;
    layer4_outputs(1470) <= a and not b;
    layer4_outputs(1471) <= not b;
    layer4_outputs(1472) <= not (a and b);
    layer4_outputs(1473) <= b and not a;
    layer4_outputs(1474) <= a;
    layer4_outputs(1475) <= not b;
    layer4_outputs(1476) <= not (a xor b);
    layer4_outputs(1477) <= a or b;
    layer4_outputs(1478) <= '0';
    layer4_outputs(1479) <= not (a xor b);
    layer4_outputs(1480) <= a;
    layer4_outputs(1481) <= not a;
    layer4_outputs(1482) <= not a or b;
    layer4_outputs(1483) <= b and not a;
    layer4_outputs(1484) <= a and b;
    layer4_outputs(1485) <= a and b;
    layer4_outputs(1486) <= not a;
    layer4_outputs(1487) <= b and not a;
    layer4_outputs(1488) <= b and not a;
    layer4_outputs(1489) <= not (a or b);
    layer4_outputs(1490) <= '1';
    layer4_outputs(1491) <= not (a or b);
    layer4_outputs(1492) <= a xor b;
    layer4_outputs(1493) <= a and b;
    layer4_outputs(1494) <= a;
    layer4_outputs(1495) <= not b;
    layer4_outputs(1496) <= b;
    layer4_outputs(1497) <= '0';
    layer4_outputs(1498) <= not b or a;
    layer4_outputs(1499) <= '0';
    layer4_outputs(1500) <= b;
    layer4_outputs(1501) <= '1';
    layer4_outputs(1502) <= not a;
    layer4_outputs(1503) <= not (a and b);
    layer4_outputs(1504) <= a;
    layer4_outputs(1505) <= not (a or b);
    layer4_outputs(1506) <= '0';
    layer4_outputs(1507) <= '1';
    layer4_outputs(1508) <= a and b;
    layer4_outputs(1509) <= a or b;
    layer4_outputs(1510) <= not (a or b);
    layer4_outputs(1511) <= not a or b;
    layer4_outputs(1512) <= not b or a;
    layer4_outputs(1513) <= not (a or b);
    layer4_outputs(1514) <= b;
    layer4_outputs(1515) <= not b or a;
    layer4_outputs(1516) <= '1';
    layer4_outputs(1517) <= b;
    layer4_outputs(1518) <= not a;
    layer4_outputs(1519) <= a and b;
    layer4_outputs(1520) <= b and not a;
    layer4_outputs(1521) <= not a or b;
    layer4_outputs(1522) <= a xor b;
    layer4_outputs(1523) <= not b or a;
    layer4_outputs(1524) <= b and not a;
    layer4_outputs(1525) <= not a or b;
    layer4_outputs(1526) <= not a;
    layer4_outputs(1527) <= '1';
    layer4_outputs(1528) <= not b or a;
    layer4_outputs(1529) <= not a or b;
    layer4_outputs(1530) <= b;
    layer4_outputs(1531) <= a and b;
    layer4_outputs(1532) <= not (a or b);
    layer4_outputs(1533) <= a and not b;
    layer4_outputs(1534) <= a and b;
    layer4_outputs(1535) <= not b or a;
    layer4_outputs(1536) <= '0';
    layer4_outputs(1537) <= not a;
    layer4_outputs(1538) <= not b;
    layer4_outputs(1539) <= '0';
    layer4_outputs(1540) <= '0';
    layer4_outputs(1541) <= not a or b;
    layer4_outputs(1542) <= a and not b;
    layer4_outputs(1543) <= b;
    layer4_outputs(1544) <= a and b;
    layer4_outputs(1545) <= not (a or b);
    layer4_outputs(1546) <= not a or b;
    layer4_outputs(1547) <= not b or a;
    layer4_outputs(1548) <= not b;
    layer4_outputs(1549) <= a and b;
    layer4_outputs(1550) <= a and not b;
    layer4_outputs(1551) <= not (a and b);
    layer4_outputs(1552) <= not b;
    layer4_outputs(1553) <= '1';
    layer4_outputs(1554) <= '1';
    layer4_outputs(1555) <= not (a xor b);
    layer4_outputs(1556) <= not a;
    layer4_outputs(1557) <= not b;
    layer4_outputs(1558) <= a xor b;
    layer4_outputs(1559) <= a and b;
    layer4_outputs(1560) <= not b or a;
    layer4_outputs(1561) <= a and not b;
    layer4_outputs(1562) <= not b or a;
    layer4_outputs(1563) <= not a;
    layer4_outputs(1564) <= '1';
    layer4_outputs(1565) <= '1';
    layer4_outputs(1566) <= b and not a;
    layer4_outputs(1567) <= not a or b;
    layer4_outputs(1568) <= a and not b;
    layer4_outputs(1569) <= not a;
    layer4_outputs(1570) <= a;
    layer4_outputs(1571) <= '0';
    layer4_outputs(1572) <= a or b;
    layer4_outputs(1573) <= not (a and b);
    layer4_outputs(1574) <= not a;
    layer4_outputs(1575) <= a and b;
    layer4_outputs(1576) <= not b or a;
    layer4_outputs(1577) <= not (a or b);
    layer4_outputs(1578) <= b and not a;
    layer4_outputs(1579) <= b and not a;
    layer4_outputs(1580) <= a and not b;
    layer4_outputs(1581) <= a and b;
    layer4_outputs(1582) <= a;
    layer4_outputs(1583) <= '0';
    layer4_outputs(1584) <= not a or b;
    layer4_outputs(1585) <= not (a and b);
    layer4_outputs(1586) <= a or b;
    layer4_outputs(1587) <= not (a or b);
    layer4_outputs(1588) <= a;
    layer4_outputs(1589) <= a;
    layer4_outputs(1590) <= b;
    layer4_outputs(1591) <= '1';
    layer4_outputs(1592) <= '1';
    layer4_outputs(1593) <= b and not a;
    layer4_outputs(1594) <= not b;
    layer4_outputs(1595) <= not b;
    layer4_outputs(1596) <= '1';
    layer4_outputs(1597) <= '0';
    layer4_outputs(1598) <= a or b;
    layer4_outputs(1599) <= not a or b;
    layer4_outputs(1600) <= not (a and b);
    layer4_outputs(1601) <= a and b;
    layer4_outputs(1602) <= a;
    layer4_outputs(1603) <= a or b;
    layer4_outputs(1604) <= not a or b;
    layer4_outputs(1605) <= '1';
    layer4_outputs(1606) <= not b;
    layer4_outputs(1607) <= a and not b;
    layer4_outputs(1608) <= a;
    layer4_outputs(1609) <= a and b;
    layer4_outputs(1610) <= a and not b;
    layer4_outputs(1611) <= b;
    layer4_outputs(1612) <= not a;
    layer4_outputs(1613) <= a and b;
    layer4_outputs(1614) <= a;
    layer4_outputs(1615) <= a or b;
    layer4_outputs(1616) <= '0';
    layer4_outputs(1617) <= not (a or b);
    layer4_outputs(1618) <= not b or a;
    layer4_outputs(1619) <= not b;
    layer4_outputs(1620) <= not b;
    layer4_outputs(1621) <= '0';
    layer4_outputs(1622) <= not (a and b);
    layer4_outputs(1623) <= not (a or b);
    layer4_outputs(1624) <= not a or b;
    layer4_outputs(1625) <= '0';
    layer4_outputs(1626) <= not b or a;
    layer4_outputs(1627) <= not (a or b);
    layer4_outputs(1628) <= not a;
    layer4_outputs(1629) <= not a or b;
    layer4_outputs(1630) <= not b;
    layer4_outputs(1631) <= a or b;
    layer4_outputs(1632) <= b;
    layer4_outputs(1633) <= b;
    layer4_outputs(1634) <= not (a or b);
    layer4_outputs(1635) <= a;
    layer4_outputs(1636) <= not b or a;
    layer4_outputs(1637) <= not (a xor b);
    layer4_outputs(1638) <= '0';
    layer4_outputs(1639) <= a and b;
    layer4_outputs(1640) <= not (a and b);
    layer4_outputs(1641) <= a xor b;
    layer4_outputs(1642) <= a or b;
    layer4_outputs(1643) <= '1';
    layer4_outputs(1644) <= not (a or b);
    layer4_outputs(1645) <= b;
    layer4_outputs(1646) <= b;
    layer4_outputs(1647) <= b;
    layer4_outputs(1648) <= not (a and b);
    layer4_outputs(1649) <= '1';
    layer4_outputs(1650) <= a and not b;
    layer4_outputs(1651) <= b and not a;
    layer4_outputs(1652) <= not a;
    layer4_outputs(1653) <= a or b;
    layer4_outputs(1654) <= a or b;
    layer4_outputs(1655) <= not b or a;
    layer4_outputs(1656) <= not (a xor b);
    layer4_outputs(1657) <= not a;
    layer4_outputs(1658) <= a and b;
    layer4_outputs(1659) <= not (a or b);
    layer4_outputs(1660) <= a and b;
    layer4_outputs(1661) <= a or b;
    layer4_outputs(1662) <= not a or b;
    layer4_outputs(1663) <= not (a or b);
    layer4_outputs(1664) <= not a;
    layer4_outputs(1665) <= not b or a;
    layer4_outputs(1666) <= a and b;
    layer4_outputs(1667) <= a and b;
    layer4_outputs(1668) <= not b;
    layer4_outputs(1669) <= b and not a;
    layer4_outputs(1670) <= a or b;
    layer4_outputs(1671) <= not a or b;
    layer4_outputs(1672) <= a;
    layer4_outputs(1673) <= '0';
    layer4_outputs(1674) <= b;
    layer4_outputs(1675) <= not a;
    layer4_outputs(1676) <= not b;
    layer4_outputs(1677) <= b and not a;
    layer4_outputs(1678) <= not (a and b);
    layer4_outputs(1679) <= not a or b;
    layer4_outputs(1680) <= not a;
    layer4_outputs(1681) <= a and not b;
    layer4_outputs(1682) <= a;
    layer4_outputs(1683) <= '0';
    layer4_outputs(1684) <= b;
    layer4_outputs(1685) <= a;
    layer4_outputs(1686) <= not (a and b);
    layer4_outputs(1687) <= not b;
    layer4_outputs(1688) <= '0';
    layer4_outputs(1689) <= b and not a;
    layer4_outputs(1690) <= a;
    layer4_outputs(1691) <= not (a and b);
    layer4_outputs(1692) <= not b or a;
    layer4_outputs(1693) <= a;
    layer4_outputs(1694) <= not b;
    layer4_outputs(1695) <= not (a or b);
    layer4_outputs(1696) <= a and b;
    layer4_outputs(1697) <= '1';
    layer4_outputs(1698) <= not (a or b);
    layer4_outputs(1699) <= a and not b;
    layer4_outputs(1700) <= not a or b;
    layer4_outputs(1701) <= a and b;
    layer4_outputs(1702) <= a or b;
    layer4_outputs(1703) <= a;
    layer4_outputs(1704) <= b;
    layer4_outputs(1705) <= a;
    layer4_outputs(1706) <= not b;
    layer4_outputs(1707) <= not (a and b);
    layer4_outputs(1708) <= not (a and b);
    layer4_outputs(1709) <= not (a or b);
    layer4_outputs(1710) <= a and not b;
    layer4_outputs(1711) <= a;
    layer4_outputs(1712) <= a and not b;
    layer4_outputs(1713) <= not (a xor b);
    layer4_outputs(1714) <= not b or a;
    layer4_outputs(1715) <= b;
    layer4_outputs(1716) <= a and b;
    layer4_outputs(1717) <= not a or b;
    layer4_outputs(1718) <= not b or a;
    layer4_outputs(1719) <= not b or a;
    layer4_outputs(1720) <= not b;
    layer4_outputs(1721) <= '1';
    layer4_outputs(1722) <= not a;
    layer4_outputs(1723) <= a;
    layer4_outputs(1724) <= a or b;
    layer4_outputs(1725) <= '0';
    layer4_outputs(1726) <= b;
    layer4_outputs(1727) <= a and not b;
    layer4_outputs(1728) <= not (a or b);
    layer4_outputs(1729) <= a;
    layer4_outputs(1730) <= not (a and b);
    layer4_outputs(1731) <= '0';
    layer4_outputs(1732) <= b and not a;
    layer4_outputs(1733) <= a and not b;
    layer4_outputs(1734) <= a;
    layer4_outputs(1735) <= a or b;
    layer4_outputs(1736) <= not a or b;
    layer4_outputs(1737) <= a or b;
    layer4_outputs(1738) <= a and b;
    layer4_outputs(1739) <= not (a and b);
    layer4_outputs(1740) <= not b;
    layer4_outputs(1741) <= a and b;
    layer4_outputs(1742) <= not (a xor b);
    layer4_outputs(1743) <= a xor b;
    layer4_outputs(1744) <= a and not b;
    layer4_outputs(1745) <= a;
    layer4_outputs(1746) <= a and b;
    layer4_outputs(1747) <= a and not b;
    layer4_outputs(1748) <= not (a xor b);
    layer4_outputs(1749) <= a and not b;
    layer4_outputs(1750) <= b and not a;
    layer4_outputs(1751) <= a;
    layer4_outputs(1752) <= not (a and b);
    layer4_outputs(1753) <= b and not a;
    layer4_outputs(1754) <= '0';
    layer4_outputs(1755) <= a;
    layer4_outputs(1756) <= a or b;
    layer4_outputs(1757) <= a or b;
    layer4_outputs(1758) <= a;
    layer4_outputs(1759) <= not (a or b);
    layer4_outputs(1760) <= a xor b;
    layer4_outputs(1761) <= a and not b;
    layer4_outputs(1762) <= not (a and b);
    layer4_outputs(1763) <= '0';
    layer4_outputs(1764) <= b;
    layer4_outputs(1765) <= a and not b;
    layer4_outputs(1766) <= not a;
    layer4_outputs(1767) <= not a or b;
    layer4_outputs(1768) <= not (a xor b);
    layer4_outputs(1769) <= not b;
    layer4_outputs(1770) <= not a;
    layer4_outputs(1771) <= '0';
    layer4_outputs(1772) <= not a;
    layer4_outputs(1773) <= a xor b;
    layer4_outputs(1774) <= a or b;
    layer4_outputs(1775) <= '1';
    layer4_outputs(1776) <= not (a xor b);
    layer4_outputs(1777) <= a and not b;
    layer4_outputs(1778) <= a or b;
    layer4_outputs(1779) <= b;
    layer4_outputs(1780) <= a or b;
    layer4_outputs(1781) <= not a or b;
    layer4_outputs(1782) <= not a or b;
    layer4_outputs(1783) <= not b;
    layer4_outputs(1784) <= a and not b;
    layer4_outputs(1785) <= not b or a;
    layer4_outputs(1786) <= b;
    layer4_outputs(1787) <= not (a or b);
    layer4_outputs(1788) <= not (a and b);
    layer4_outputs(1789) <= not (a or b);
    layer4_outputs(1790) <= a and b;
    layer4_outputs(1791) <= not b or a;
    layer4_outputs(1792) <= b;
    layer4_outputs(1793) <= a;
    layer4_outputs(1794) <= b and not a;
    layer4_outputs(1795) <= not a or b;
    layer4_outputs(1796) <= not b or a;
    layer4_outputs(1797) <= not b or a;
    layer4_outputs(1798) <= '1';
    layer4_outputs(1799) <= not b;
    layer4_outputs(1800) <= b and not a;
    layer4_outputs(1801) <= a and b;
    layer4_outputs(1802) <= not b;
    layer4_outputs(1803) <= b;
    layer4_outputs(1804) <= not a;
    layer4_outputs(1805) <= b;
    layer4_outputs(1806) <= a;
    layer4_outputs(1807) <= a;
    layer4_outputs(1808) <= a and b;
    layer4_outputs(1809) <= a and not b;
    layer4_outputs(1810) <= '1';
    layer4_outputs(1811) <= b;
    layer4_outputs(1812) <= a or b;
    layer4_outputs(1813) <= b;
    layer4_outputs(1814) <= not a;
    layer4_outputs(1815) <= '1';
    layer4_outputs(1816) <= not b or a;
    layer4_outputs(1817) <= not b;
    layer4_outputs(1818) <= '0';
    layer4_outputs(1819) <= a;
    layer4_outputs(1820) <= a or b;
    layer4_outputs(1821) <= b;
    layer4_outputs(1822) <= a;
    layer4_outputs(1823) <= '0';
    layer4_outputs(1824) <= '1';
    layer4_outputs(1825) <= a or b;
    layer4_outputs(1826) <= a and not b;
    layer4_outputs(1827) <= b;
    layer4_outputs(1828) <= a and not b;
    layer4_outputs(1829) <= not a or b;
    layer4_outputs(1830) <= not b;
    layer4_outputs(1831) <= not (a and b);
    layer4_outputs(1832) <= not b;
    layer4_outputs(1833) <= not b or a;
    layer4_outputs(1834) <= not b;
    layer4_outputs(1835) <= a;
    layer4_outputs(1836) <= '0';
    layer4_outputs(1837) <= '0';
    layer4_outputs(1838) <= '1';
    layer4_outputs(1839) <= '0';
    layer4_outputs(1840) <= not a;
    layer4_outputs(1841) <= not b;
    layer4_outputs(1842) <= a and b;
    layer4_outputs(1843) <= '0';
    layer4_outputs(1844) <= not a or b;
    layer4_outputs(1845) <= b;
    layer4_outputs(1846) <= b and not a;
    layer4_outputs(1847) <= not (a or b);
    layer4_outputs(1848) <= a and not b;
    layer4_outputs(1849) <= a and b;
    layer4_outputs(1850) <= a and b;
    layer4_outputs(1851) <= not b;
    layer4_outputs(1852) <= a and b;
    layer4_outputs(1853) <= not a;
    layer4_outputs(1854) <= a and b;
    layer4_outputs(1855) <= a;
    layer4_outputs(1856) <= '1';
    layer4_outputs(1857) <= not b;
    layer4_outputs(1858) <= b and not a;
    layer4_outputs(1859) <= b;
    layer4_outputs(1860) <= a;
    layer4_outputs(1861) <= not a or b;
    layer4_outputs(1862) <= b and not a;
    layer4_outputs(1863) <= a and b;
    layer4_outputs(1864) <= not b;
    layer4_outputs(1865) <= a and not b;
    layer4_outputs(1866) <= '1';
    layer4_outputs(1867) <= not a;
    layer4_outputs(1868) <= a and not b;
    layer4_outputs(1869) <= not b;
    layer4_outputs(1870) <= not a or b;
    layer4_outputs(1871) <= not (a and b);
    layer4_outputs(1872) <= a or b;
    layer4_outputs(1873) <= not (a xor b);
    layer4_outputs(1874) <= a and b;
    layer4_outputs(1875) <= '1';
    layer4_outputs(1876) <= '1';
    layer4_outputs(1877) <= not a or b;
    layer4_outputs(1878) <= not b;
    layer4_outputs(1879) <= b and not a;
    layer4_outputs(1880) <= not (a or b);
    layer4_outputs(1881) <= not a or b;
    layer4_outputs(1882) <= b and not a;
    layer4_outputs(1883) <= '1';
    layer4_outputs(1884) <= '0';
    layer4_outputs(1885) <= not b or a;
    layer4_outputs(1886) <= '0';
    layer4_outputs(1887) <= a and not b;
    layer4_outputs(1888) <= not b or a;
    layer4_outputs(1889) <= a;
    layer4_outputs(1890) <= a;
    layer4_outputs(1891) <= not b;
    layer4_outputs(1892) <= a and not b;
    layer4_outputs(1893) <= not (a or b);
    layer4_outputs(1894) <= a;
    layer4_outputs(1895) <= a;
    layer4_outputs(1896) <= a and b;
    layer4_outputs(1897) <= a and not b;
    layer4_outputs(1898) <= a and b;
    layer4_outputs(1899) <= '1';
    layer4_outputs(1900) <= a and not b;
    layer4_outputs(1901) <= not (a and b);
    layer4_outputs(1902) <= not b or a;
    layer4_outputs(1903) <= '1';
    layer4_outputs(1904) <= not b;
    layer4_outputs(1905) <= not (a xor b);
    layer4_outputs(1906) <= not b or a;
    layer4_outputs(1907) <= not (a xor b);
    layer4_outputs(1908) <= a and not b;
    layer4_outputs(1909) <= a;
    layer4_outputs(1910) <= '0';
    layer4_outputs(1911) <= b;
    layer4_outputs(1912) <= a xor b;
    layer4_outputs(1913) <= not b;
    layer4_outputs(1914) <= a and not b;
    layer4_outputs(1915) <= not (a and b);
    layer4_outputs(1916) <= a or b;
    layer4_outputs(1917) <= '1';
    layer4_outputs(1918) <= a and not b;
    layer4_outputs(1919) <= a and not b;
    layer4_outputs(1920) <= a and b;
    layer4_outputs(1921) <= a and not b;
    layer4_outputs(1922) <= '0';
    layer4_outputs(1923) <= not (a and b);
    layer4_outputs(1924) <= not b or a;
    layer4_outputs(1925) <= a or b;
    layer4_outputs(1926) <= '1';
    layer4_outputs(1927) <= not b or a;
    layer4_outputs(1928) <= b and not a;
    layer4_outputs(1929) <= not b;
    layer4_outputs(1930) <= '1';
    layer4_outputs(1931) <= '1';
    layer4_outputs(1932) <= b;
    layer4_outputs(1933) <= a and not b;
    layer4_outputs(1934) <= not (a or b);
    layer4_outputs(1935) <= a and b;
    layer4_outputs(1936) <= not a;
    layer4_outputs(1937) <= '0';
    layer4_outputs(1938) <= not (a and b);
    layer4_outputs(1939) <= not a;
    layer4_outputs(1940) <= not (a or b);
    layer4_outputs(1941) <= not a;
    layer4_outputs(1942) <= '1';
    layer4_outputs(1943) <= a and b;
    layer4_outputs(1944) <= not b or a;
    layer4_outputs(1945) <= not b or a;
    layer4_outputs(1946) <= a or b;
    layer4_outputs(1947) <= b and not a;
    layer4_outputs(1948) <= a and not b;
    layer4_outputs(1949) <= not a;
    layer4_outputs(1950) <= a and not b;
    layer4_outputs(1951) <= not a or b;
    layer4_outputs(1952) <= b and not a;
    layer4_outputs(1953) <= a;
    layer4_outputs(1954) <= '0';
    layer4_outputs(1955) <= '1';
    layer4_outputs(1956) <= a or b;
    layer4_outputs(1957) <= not b or a;
    layer4_outputs(1958) <= b and not a;
    layer4_outputs(1959) <= a;
    layer4_outputs(1960) <= not b;
    layer4_outputs(1961) <= not b or a;
    layer4_outputs(1962) <= b;
    layer4_outputs(1963) <= not b;
    layer4_outputs(1964) <= not a;
    layer4_outputs(1965) <= '0';
    layer4_outputs(1966) <= not (a or b);
    layer4_outputs(1967) <= a and not b;
    layer4_outputs(1968) <= not (a and b);
    layer4_outputs(1969) <= a or b;
    layer4_outputs(1970) <= not a or b;
    layer4_outputs(1971) <= not b or a;
    layer4_outputs(1972) <= a and b;
    layer4_outputs(1973) <= '1';
    layer4_outputs(1974) <= not b;
    layer4_outputs(1975) <= not a or b;
    layer4_outputs(1976) <= a;
    layer4_outputs(1977) <= '1';
    layer4_outputs(1978) <= not (a and b);
    layer4_outputs(1979) <= not (a and b);
    layer4_outputs(1980) <= '1';
    layer4_outputs(1981) <= not a;
    layer4_outputs(1982) <= not b or a;
    layer4_outputs(1983) <= b and not a;
    layer4_outputs(1984) <= not b or a;
    layer4_outputs(1985) <= not a or b;
    layer4_outputs(1986) <= '1';
    layer4_outputs(1987) <= a xor b;
    layer4_outputs(1988) <= b;
    layer4_outputs(1989) <= not a;
    layer4_outputs(1990) <= a and not b;
    layer4_outputs(1991) <= '1';
    layer4_outputs(1992) <= a;
    layer4_outputs(1993) <= not a;
    layer4_outputs(1994) <= not b;
    layer4_outputs(1995) <= not b;
    layer4_outputs(1996) <= not b or a;
    layer4_outputs(1997) <= not a;
    layer4_outputs(1998) <= not (a and b);
    layer4_outputs(1999) <= not a or b;
    layer4_outputs(2000) <= not b or a;
    layer4_outputs(2001) <= a or b;
    layer4_outputs(2002) <= b and not a;
    layer4_outputs(2003) <= not a;
    layer4_outputs(2004) <= not b;
    layer4_outputs(2005) <= a and not b;
    layer4_outputs(2006) <= a and not b;
    layer4_outputs(2007) <= not a;
    layer4_outputs(2008) <= '1';
    layer4_outputs(2009) <= not (a and b);
    layer4_outputs(2010) <= b;
    layer4_outputs(2011) <= '0';
    layer4_outputs(2012) <= a and not b;
    layer4_outputs(2013) <= b and not a;
    layer4_outputs(2014) <= a and not b;
    layer4_outputs(2015) <= not (a and b);
    layer4_outputs(2016) <= not a;
    layer4_outputs(2017) <= a or b;
    layer4_outputs(2018) <= not b or a;
    layer4_outputs(2019) <= not a;
    layer4_outputs(2020) <= '0';
    layer4_outputs(2021) <= '1';
    layer4_outputs(2022) <= not (a and b);
    layer4_outputs(2023) <= not a;
    layer4_outputs(2024) <= not b;
    layer4_outputs(2025) <= not (a or b);
    layer4_outputs(2026) <= '1';
    layer4_outputs(2027) <= a;
    layer4_outputs(2028) <= a;
    layer4_outputs(2029) <= not a;
    layer4_outputs(2030) <= a;
    layer4_outputs(2031) <= b;
    layer4_outputs(2032) <= not (a xor b);
    layer4_outputs(2033) <= '1';
    layer4_outputs(2034) <= not (a and b);
    layer4_outputs(2035) <= '1';
    layer4_outputs(2036) <= a and not b;
    layer4_outputs(2037) <= not b;
    layer4_outputs(2038) <= not (a or b);
    layer4_outputs(2039) <= a or b;
    layer4_outputs(2040) <= b;
    layer4_outputs(2041) <= a and b;
    layer4_outputs(2042) <= not b or a;
    layer4_outputs(2043) <= b and not a;
    layer4_outputs(2044) <= not (a and b);
    layer4_outputs(2045) <= a or b;
    layer4_outputs(2046) <= not (a and b);
    layer4_outputs(2047) <= not (a xor b);
    layer4_outputs(2048) <= b;
    layer4_outputs(2049) <= not (a and b);
    layer4_outputs(2050) <= b;
    layer4_outputs(2051) <= a xor b;
    layer4_outputs(2052) <= b and not a;
    layer4_outputs(2053) <= a;
    layer4_outputs(2054) <= b and not a;
    layer4_outputs(2055) <= not b or a;
    layer4_outputs(2056) <= not (a or b);
    layer4_outputs(2057) <= not (a or b);
    layer4_outputs(2058) <= '0';
    layer4_outputs(2059) <= a and b;
    layer4_outputs(2060) <= not a;
    layer4_outputs(2061) <= not a;
    layer4_outputs(2062) <= b;
    layer4_outputs(2063) <= not a;
    layer4_outputs(2064) <= '1';
    layer4_outputs(2065) <= not b;
    layer4_outputs(2066) <= not (a or b);
    layer4_outputs(2067) <= b and not a;
    layer4_outputs(2068) <= not a;
    layer4_outputs(2069) <= not a;
    layer4_outputs(2070) <= not b or a;
    layer4_outputs(2071) <= not (a and b);
    layer4_outputs(2072) <= not a;
    layer4_outputs(2073) <= a or b;
    layer4_outputs(2074) <= b;
    layer4_outputs(2075) <= a or b;
    layer4_outputs(2076) <= not b or a;
    layer4_outputs(2077) <= not (a or b);
    layer4_outputs(2078) <= not a or b;
    layer4_outputs(2079) <= not (a or b);
    layer4_outputs(2080) <= a xor b;
    layer4_outputs(2081) <= a xor b;
    layer4_outputs(2082) <= not (a or b);
    layer4_outputs(2083) <= b and not a;
    layer4_outputs(2084) <= not b or a;
    layer4_outputs(2085) <= b;
    layer4_outputs(2086) <= a xor b;
    layer4_outputs(2087) <= not b or a;
    layer4_outputs(2088) <= b and not a;
    layer4_outputs(2089) <= b;
    layer4_outputs(2090) <= not b;
    layer4_outputs(2091) <= not a or b;
    layer4_outputs(2092) <= a;
    layer4_outputs(2093) <= b and not a;
    layer4_outputs(2094) <= not (a xor b);
    layer4_outputs(2095) <= not (a and b);
    layer4_outputs(2096) <= a;
    layer4_outputs(2097) <= not a;
    layer4_outputs(2098) <= not b;
    layer4_outputs(2099) <= '1';
    layer4_outputs(2100) <= b and not a;
    layer4_outputs(2101) <= a and b;
    layer4_outputs(2102) <= a and b;
    layer4_outputs(2103) <= not (a or b);
    layer4_outputs(2104) <= not a or b;
    layer4_outputs(2105) <= not (a or b);
    layer4_outputs(2106) <= not a or b;
    layer4_outputs(2107) <= '0';
    layer4_outputs(2108) <= a or b;
    layer4_outputs(2109) <= b and not a;
    layer4_outputs(2110) <= b and not a;
    layer4_outputs(2111) <= not a or b;
    layer4_outputs(2112) <= not a;
    layer4_outputs(2113) <= b;
    layer4_outputs(2114) <= not b;
    layer4_outputs(2115) <= '0';
    layer4_outputs(2116) <= b and not a;
    layer4_outputs(2117) <= a and not b;
    layer4_outputs(2118) <= '1';
    layer4_outputs(2119) <= '0';
    layer4_outputs(2120) <= not (a and b);
    layer4_outputs(2121) <= not (a or b);
    layer4_outputs(2122) <= b;
    layer4_outputs(2123) <= a or b;
    layer4_outputs(2124) <= a;
    layer4_outputs(2125) <= '0';
    layer4_outputs(2126) <= not (a or b);
    layer4_outputs(2127) <= not b;
    layer4_outputs(2128) <= not a or b;
    layer4_outputs(2129) <= a or b;
    layer4_outputs(2130) <= b and not a;
    layer4_outputs(2131) <= not (a and b);
    layer4_outputs(2132) <= not (a and b);
    layer4_outputs(2133) <= b and not a;
    layer4_outputs(2134) <= not a or b;
    layer4_outputs(2135) <= '0';
    layer4_outputs(2136) <= b and not a;
    layer4_outputs(2137) <= b;
    layer4_outputs(2138) <= a;
    layer4_outputs(2139) <= not a;
    layer4_outputs(2140) <= b and not a;
    layer4_outputs(2141) <= a xor b;
    layer4_outputs(2142) <= a and b;
    layer4_outputs(2143) <= not (a or b);
    layer4_outputs(2144) <= '1';
    layer4_outputs(2145) <= '0';
    layer4_outputs(2146) <= a and b;
    layer4_outputs(2147) <= a;
    layer4_outputs(2148) <= not a;
    layer4_outputs(2149) <= not a or b;
    layer4_outputs(2150) <= not b;
    layer4_outputs(2151) <= '0';
    layer4_outputs(2152) <= b and not a;
    layer4_outputs(2153) <= not a;
    layer4_outputs(2154) <= b;
    layer4_outputs(2155) <= '0';
    layer4_outputs(2156) <= not (a and b);
    layer4_outputs(2157) <= b;
    layer4_outputs(2158) <= not a;
    layer4_outputs(2159) <= a xor b;
    layer4_outputs(2160) <= not (a xor b);
    layer4_outputs(2161) <= not b or a;
    layer4_outputs(2162) <= '0';
    layer4_outputs(2163) <= not b or a;
    layer4_outputs(2164) <= b and not a;
    layer4_outputs(2165) <= not b or a;
    layer4_outputs(2166) <= a;
    layer4_outputs(2167) <= a and not b;
    layer4_outputs(2168) <= a and b;
    layer4_outputs(2169) <= b and not a;
    layer4_outputs(2170) <= '0';
    layer4_outputs(2171) <= not a;
    layer4_outputs(2172) <= '1';
    layer4_outputs(2173) <= not b or a;
    layer4_outputs(2174) <= not a;
    layer4_outputs(2175) <= a;
    layer4_outputs(2176) <= not (a or b);
    layer4_outputs(2177) <= a or b;
    layer4_outputs(2178) <= not b;
    layer4_outputs(2179) <= a;
    layer4_outputs(2180) <= a and not b;
    layer4_outputs(2181) <= a and not b;
    layer4_outputs(2182) <= not a or b;
    layer4_outputs(2183) <= b;
    layer4_outputs(2184) <= b;
    layer4_outputs(2185) <= a and b;
    layer4_outputs(2186) <= '1';
    layer4_outputs(2187) <= a and b;
    layer4_outputs(2188) <= '1';
    layer4_outputs(2189) <= not b;
    layer4_outputs(2190) <= not a or b;
    layer4_outputs(2191) <= '0';
    layer4_outputs(2192) <= not (a and b);
    layer4_outputs(2193) <= not (a and b);
    layer4_outputs(2194) <= not b;
    layer4_outputs(2195) <= a or b;
    layer4_outputs(2196) <= b and not a;
    layer4_outputs(2197) <= not (a and b);
    layer4_outputs(2198) <= a and not b;
    layer4_outputs(2199) <= not a;
    layer4_outputs(2200) <= '1';
    layer4_outputs(2201) <= a and b;
    layer4_outputs(2202) <= '1';
    layer4_outputs(2203) <= not a or b;
    layer4_outputs(2204) <= b and not a;
    layer4_outputs(2205) <= not (a and b);
    layer4_outputs(2206) <= not b or a;
    layer4_outputs(2207) <= b;
    layer4_outputs(2208) <= a and not b;
    layer4_outputs(2209) <= b;
    layer4_outputs(2210) <= not a;
    layer4_outputs(2211) <= not b or a;
    layer4_outputs(2212) <= a;
    layer4_outputs(2213) <= a and b;
    layer4_outputs(2214) <= b and not a;
    layer4_outputs(2215) <= not a;
    layer4_outputs(2216) <= '1';
    layer4_outputs(2217) <= a and not b;
    layer4_outputs(2218) <= b;
    layer4_outputs(2219) <= b;
    layer4_outputs(2220) <= not (a and b);
    layer4_outputs(2221) <= '0';
    layer4_outputs(2222) <= b;
    layer4_outputs(2223) <= '0';
    layer4_outputs(2224) <= a and not b;
    layer4_outputs(2225) <= a;
    layer4_outputs(2226) <= b and not a;
    layer4_outputs(2227) <= '0';
    layer4_outputs(2228) <= not (a and b);
    layer4_outputs(2229) <= not a;
    layer4_outputs(2230) <= '1';
    layer4_outputs(2231) <= b;
    layer4_outputs(2232) <= not a or b;
    layer4_outputs(2233) <= b;
    layer4_outputs(2234) <= a and b;
    layer4_outputs(2235) <= b;
    layer4_outputs(2236) <= not (a and b);
    layer4_outputs(2237) <= not (a or b);
    layer4_outputs(2238) <= '1';
    layer4_outputs(2239) <= not a;
    layer4_outputs(2240) <= not b or a;
    layer4_outputs(2241) <= a;
    layer4_outputs(2242) <= '0';
    layer4_outputs(2243) <= a or b;
    layer4_outputs(2244) <= not a or b;
    layer4_outputs(2245) <= not b or a;
    layer4_outputs(2246) <= not b or a;
    layer4_outputs(2247) <= not b;
    layer4_outputs(2248) <= not a or b;
    layer4_outputs(2249) <= not a or b;
    layer4_outputs(2250) <= not b or a;
    layer4_outputs(2251) <= not b;
    layer4_outputs(2252) <= '0';
    layer4_outputs(2253) <= not (a or b);
    layer4_outputs(2254) <= a and not b;
    layer4_outputs(2255) <= a or b;
    layer4_outputs(2256) <= not b;
    layer4_outputs(2257) <= not (a xor b);
    layer4_outputs(2258) <= a;
    layer4_outputs(2259) <= not b or a;
    layer4_outputs(2260) <= '0';
    layer4_outputs(2261) <= '1';
    layer4_outputs(2262) <= '1';
    layer4_outputs(2263) <= a xor b;
    layer4_outputs(2264) <= not (a or b);
    layer4_outputs(2265) <= not (a and b);
    layer4_outputs(2266) <= b and not a;
    layer4_outputs(2267) <= not a;
    layer4_outputs(2268) <= '0';
    layer4_outputs(2269) <= not (a or b);
    layer4_outputs(2270) <= not b or a;
    layer4_outputs(2271) <= a and not b;
    layer4_outputs(2272) <= not (a or b);
    layer4_outputs(2273) <= b;
    layer4_outputs(2274) <= not a;
    layer4_outputs(2275) <= not a;
    layer4_outputs(2276) <= b and not a;
    layer4_outputs(2277) <= not a or b;
    layer4_outputs(2278) <= b and not a;
    layer4_outputs(2279) <= b;
    layer4_outputs(2280) <= not a;
    layer4_outputs(2281) <= '1';
    layer4_outputs(2282) <= not b or a;
    layer4_outputs(2283) <= b;
    layer4_outputs(2284) <= '1';
    layer4_outputs(2285) <= not b;
    layer4_outputs(2286) <= a or b;
    layer4_outputs(2287) <= a and not b;
    layer4_outputs(2288) <= '1';
    layer4_outputs(2289) <= not (a and b);
    layer4_outputs(2290) <= not b;
    layer4_outputs(2291) <= not (a xor b);
    layer4_outputs(2292) <= not a;
    layer4_outputs(2293) <= b;
    layer4_outputs(2294) <= b and not a;
    layer4_outputs(2295) <= b;
    layer4_outputs(2296) <= a;
    layer4_outputs(2297) <= a or b;
    layer4_outputs(2298) <= a or b;
    layer4_outputs(2299) <= not b;
    layer4_outputs(2300) <= b;
    layer4_outputs(2301) <= not a;
    layer4_outputs(2302) <= a and b;
    layer4_outputs(2303) <= not a or b;
    layer4_outputs(2304) <= a;
    layer4_outputs(2305) <= a and not b;
    layer4_outputs(2306) <= not (a xor b);
    layer4_outputs(2307) <= b;
    layer4_outputs(2308) <= not (a or b);
    layer4_outputs(2309) <= not a or b;
    layer4_outputs(2310) <= b and not a;
    layer4_outputs(2311) <= a and not b;
    layer4_outputs(2312) <= not b;
    layer4_outputs(2313) <= not (a xor b);
    layer4_outputs(2314) <= not a;
    layer4_outputs(2315) <= b and not a;
    layer4_outputs(2316) <= not a;
    layer4_outputs(2317) <= a and not b;
    layer4_outputs(2318) <= '0';
    layer4_outputs(2319) <= not b;
    layer4_outputs(2320) <= a and not b;
    layer4_outputs(2321) <= not b or a;
    layer4_outputs(2322) <= '1';
    layer4_outputs(2323) <= not (a or b);
    layer4_outputs(2324) <= not b;
    layer4_outputs(2325) <= not (a xor b);
    layer4_outputs(2326) <= a and not b;
    layer4_outputs(2327) <= a xor b;
    layer4_outputs(2328) <= a;
    layer4_outputs(2329) <= not b or a;
    layer4_outputs(2330) <= not (a xor b);
    layer4_outputs(2331) <= b and not a;
    layer4_outputs(2332) <= a and b;
    layer4_outputs(2333) <= '1';
    layer4_outputs(2334) <= not a or b;
    layer4_outputs(2335) <= not (a and b);
    layer4_outputs(2336) <= a and not b;
    layer4_outputs(2337) <= a and b;
    layer4_outputs(2338) <= a or b;
    layer4_outputs(2339) <= not (a and b);
    layer4_outputs(2340) <= a;
    layer4_outputs(2341) <= b and not a;
    layer4_outputs(2342) <= not (a or b);
    layer4_outputs(2343) <= not b or a;
    layer4_outputs(2344) <= not (a or b);
    layer4_outputs(2345) <= a or b;
    layer4_outputs(2346) <= b;
    layer4_outputs(2347) <= not b or a;
    layer4_outputs(2348) <= not b;
    layer4_outputs(2349) <= a;
    layer4_outputs(2350) <= not b;
    layer4_outputs(2351) <= not b or a;
    layer4_outputs(2352) <= a or b;
    layer4_outputs(2353) <= '0';
    layer4_outputs(2354) <= b;
    layer4_outputs(2355) <= not b or a;
    layer4_outputs(2356) <= a and not b;
    layer4_outputs(2357) <= not a or b;
    layer4_outputs(2358) <= a and not b;
    layer4_outputs(2359) <= a or b;
    layer4_outputs(2360) <= a or b;
    layer4_outputs(2361) <= a;
    layer4_outputs(2362) <= not a;
    layer4_outputs(2363) <= not a or b;
    layer4_outputs(2364) <= '1';
    layer4_outputs(2365) <= not (a xor b);
    layer4_outputs(2366) <= b;
    layer4_outputs(2367) <= '0';
    layer4_outputs(2368) <= not (a or b);
    layer4_outputs(2369) <= not (a or b);
    layer4_outputs(2370) <= '1';
    layer4_outputs(2371) <= '1';
    layer4_outputs(2372) <= not (a and b);
    layer4_outputs(2373) <= a;
    layer4_outputs(2374) <= a xor b;
    layer4_outputs(2375) <= not b or a;
    layer4_outputs(2376) <= b;
    layer4_outputs(2377) <= a and b;
    layer4_outputs(2378) <= b and not a;
    layer4_outputs(2379) <= not (a and b);
    layer4_outputs(2380) <= b;
    layer4_outputs(2381) <= a or b;
    layer4_outputs(2382) <= a and b;
    layer4_outputs(2383) <= '1';
    layer4_outputs(2384) <= a and b;
    layer4_outputs(2385) <= not (a or b);
    layer4_outputs(2386) <= '1';
    layer4_outputs(2387) <= not a or b;
    layer4_outputs(2388) <= a;
    layer4_outputs(2389) <= b;
    layer4_outputs(2390) <= a and b;
    layer4_outputs(2391) <= not (a and b);
    layer4_outputs(2392) <= b and not a;
    layer4_outputs(2393) <= not (a or b);
    layer4_outputs(2394) <= b;
    layer4_outputs(2395) <= b;
    layer4_outputs(2396) <= not (a or b);
    layer4_outputs(2397) <= a xor b;
    layer4_outputs(2398) <= not b or a;
    layer4_outputs(2399) <= not (a xor b);
    layer4_outputs(2400) <= not (a or b);
    layer4_outputs(2401) <= a and not b;
    layer4_outputs(2402) <= a and not b;
    layer4_outputs(2403) <= a or b;
    layer4_outputs(2404) <= '1';
    layer4_outputs(2405) <= a and not b;
    layer4_outputs(2406) <= not (a or b);
    layer4_outputs(2407) <= not (a or b);
    layer4_outputs(2408) <= b;
    layer4_outputs(2409) <= not b;
    layer4_outputs(2410) <= a;
    layer4_outputs(2411) <= b and not a;
    layer4_outputs(2412) <= b;
    layer4_outputs(2413) <= a and b;
    layer4_outputs(2414) <= '0';
    layer4_outputs(2415) <= b;
    layer4_outputs(2416) <= b and not a;
    layer4_outputs(2417) <= not (a or b);
    layer4_outputs(2418) <= not (a and b);
    layer4_outputs(2419) <= b and not a;
    layer4_outputs(2420) <= not a;
    layer4_outputs(2421) <= not a or b;
    layer4_outputs(2422) <= a xor b;
    layer4_outputs(2423) <= not a;
    layer4_outputs(2424) <= a and not b;
    layer4_outputs(2425) <= a and b;
    layer4_outputs(2426) <= not a or b;
    layer4_outputs(2427) <= b;
    layer4_outputs(2428) <= not (a or b);
    layer4_outputs(2429) <= not (a or b);
    layer4_outputs(2430) <= not (a and b);
    layer4_outputs(2431) <= not b or a;
    layer4_outputs(2432) <= a;
    layer4_outputs(2433) <= a or b;
    layer4_outputs(2434) <= not a;
    layer4_outputs(2435) <= '1';
    layer4_outputs(2436) <= b and not a;
    layer4_outputs(2437) <= a and b;
    layer4_outputs(2438) <= a;
    layer4_outputs(2439) <= not (a or b);
    layer4_outputs(2440) <= not b;
    layer4_outputs(2441) <= a;
    layer4_outputs(2442) <= a or b;
    layer4_outputs(2443) <= not (a xor b);
    layer4_outputs(2444) <= a and b;
    layer4_outputs(2445) <= a;
    layer4_outputs(2446) <= '1';
    layer4_outputs(2447) <= b and not a;
    layer4_outputs(2448) <= not (a and b);
    layer4_outputs(2449) <= '0';
    layer4_outputs(2450) <= not a;
    layer4_outputs(2451) <= b;
    layer4_outputs(2452) <= b;
    layer4_outputs(2453) <= '0';
    layer4_outputs(2454) <= a;
    layer4_outputs(2455) <= not b or a;
    layer4_outputs(2456) <= a and b;
    layer4_outputs(2457) <= a xor b;
    layer4_outputs(2458) <= '0';
    layer4_outputs(2459) <= b and not a;
    layer4_outputs(2460) <= '0';
    layer4_outputs(2461) <= a;
    layer4_outputs(2462) <= b and not a;
    layer4_outputs(2463) <= a xor b;
    layer4_outputs(2464) <= not (a and b);
    layer4_outputs(2465) <= b;
    layer4_outputs(2466) <= a;
    layer4_outputs(2467) <= a and b;
    layer4_outputs(2468) <= a and b;
    layer4_outputs(2469) <= not a;
    layer4_outputs(2470) <= not b or a;
    layer4_outputs(2471) <= '1';
    layer4_outputs(2472) <= b;
    layer4_outputs(2473) <= b;
    layer4_outputs(2474) <= a and b;
    layer4_outputs(2475) <= b and not a;
    layer4_outputs(2476) <= a;
    layer4_outputs(2477) <= b;
    layer4_outputs(2478) <= '1';
    layer4_outputs(2479) <= not b;
    layer4_outputs(2480) <= not b;
    layer4_outputs(2481) <= a or b;
    layer4_outputs(2482) <= b;
    layer4_outputs(2483) <= not (a and b);
    layer4_outputs(2484) <= b and not a;
    layer4_outputs(2485) <= not (a or b);
    layer4_outputs(2486) <= not b or a;
    layer4_outputs(2487) <= b;
    layer4_outputs(2488) <= b;
    layer4_outputs(2489) <= a or b;
    layer4_outputs(2490) <= not b;
    layer4_outputs(2491) <= not a or b;
    layer4_outputs(2492) <= b and not a;
    layer4_outputs(2493) <= b and not a;
    layer4_outputs(2494) <= not a or b;
    layer4_outputs(2495) <= b;
    layer4_outputs(2496) <= not (a or b);
    layer4_outputs(2497) <= not b;
    layer4_outputs(2498) <= not b;
    layer4_outputs(2499) <= not a;
    layer4_outputs(2500) <= a and not b;
    layer4_outputs(2501) <= a;
    layer4_outputs(2502) <= a;
    layer4_outputs(2503) <= not b or a;
    layer4_outputs(2504) <= not (a and b);
    layer4_outputs(2505) <= a xor b;
    layer4_outputs(2506) <= '0';
    layer4_outputs(2507) <= not (a or b);
    layer4_outputs(2508) <= a and b;
    layer4_outputs(2509) <= not (a and b);
    layer4_outputs(2510) <= a and b;
    layer4_outputs(2511) <= a xor b;
    layer4_outputs(2512) <= a;
    layer4_outputs(2513) <= b and not a;
    layer4_outputs(2514) <= a and not b;
    layer4_outputs(2515) <= not b or a;
    layer4_outputs(2516) <= not b;
    layer4_outputs(2517) <= not (a or b);
    layer4_outputs(2518) <= not b;
    layer4_outputs(2519) <= a and not b;
    layer4_outputs(2520) <= b and not a;
    layer4_outputs(2521) <= a and b;
    layer4_outputs(2522) <= not (a and b);
    layer4_outputs(2523) <= not b or a;
    layer4_outputs(2524) <= a;
    layer4_outputs(2525) <= '1';
    layer4_outputs(2526) <= not a or b;
    layer4_outputs(2527) <= b;
    layer4_outputs(2528) <= a and b;
    layer4_outputs(2529) <= not a or b;
    layer4_outputs(2530) <= a;
    layer4_outputs(2531) <= a;
    layer4_outputs(2532) <= not a or b;
    layer4_outputs(2533) <= b;
    layer4_outputs(2534) <= not b or a;
    layer4_outputs(2535) <= a or b;
    layer4_outputs(2536) <= not a;
    layer4_outputs(2537) <= not b or a;
    layer4_outputs(2538) <= not b or a;
    layer4_outputs(2539) <= not b or a;
    layer4_outputs(2540) <= b;
    layer4_outputs(2541) <= not b;
    layer4_outputs(2542) <= b and not a;
    layer4_outputs(2543) <= a and not b;
    layer4_outputs(2544) <= a and b;
    layer4_outputs(2545) <= a;
    layer4_outputs(2546) <= not b;
    layer4_outputs(2547) <= not b or a;
    layer4_outputs(2548) <= a or b;
    layer4_outputs(2549) <= '1';
    layer4_outputs(2550) <= not a or b;
    layer4_outputs(2551) <= not (a and b);
    layer4_outputs(2552) <= b;
    layer4_outputs(2553) <= a;
    layer4_outputs(2554) <= not a;
    layer4_outputs(2555) <= not (a or b);
    layer4_outputs(2556) <= not b or a;
    layer4_outputs(2557) <= not (a and b);
    layer4_outputs(2558) <= a and not b;
    layer4_outputs(2559) <= not b;
    layer4_outputs(2560) <= not b;
    layer4_outputs(2561) <= a and not b;
    layer4_outputs(2562) <= b and not a;
    layer4_outputs(2563) <= not b;
    layer4_outputs(2564) <= not a or b;
    layer4_outputs(2565) <= not b;
    layer4_outputs(2566) <= a;
    layer4_outputs(2567) <= not (a or b);
    layer4_outputs(2568) <= not b or a;
    layer4_outputs(2569) <= not (a or b);
    layer4_outputs(2570) <= '1';
    layer4_outputs(2571) <= not a;
    layer4_outputs(2572) <= b and not a;
    layer4_outputs(2573) <= '1';
    layer4_outputs(2574) <= not a;
    layer4_outputs(2575) <= not (a or b);
    layer4_outputs(2576) <= a;
    layer4_outputs(2577) <= not a;
    layer4_outputs(2578) <= a;
    layer4_outputs(2579) <= not (a and b);
    layer4_outputs(2580) <= not b or a;
    layer4_outputs(2581) <= not b or a;
    layer4_outputs(2582) <= not (a and b);
    layer4_outputs(2583) <= not a;
    layer4_outputs(2584) <= not b or a;
    layer4_outputs(2585) <= not b or a;
    layer4_outputs(2586) <= not b;
    layer4_outputs(2587) <= b;
    layer4_outputs(2588) <= not (a or b);
    layer4_outputs(2589) <= a and not b;
    layer4_outputs(2590) <= not a;
    layer4_outputs(2591) <= a;
    layer4_outputs(2592) <= not a or b;
    layer4_outputs(2593) <= not a or b;
    layer4_outputs(2594) <= a or b;
    layer4_outputs(2595) <= not (a or b);
    layer4_outputs(2596) <= not (a or b);
    layer4_outputs(2597) <= not (a and b);
    layer4_outputs(2598) <= b and not a;
    layer4_outputs(2599) <= not (a or b);
    layer4_outputs(2600) <= not a;
    layer4_outputs(2601) <= not a;
    layer4_outputs(2602) <= '0';
    layer4_outputs(2603) <= not b;
    layer4_outputs(2604) <= b;
    layer4_outputs(2605) <= a and not b;
    layer4_outputs(2606) <= a and not b;
    layer4_outputs(2607) <= not b;
    layer4_outputs(2608) <= a and b;
    layer4_outputs(2609) <= b;
    layer4_outputs(2610) <= a or b;
    layer4_outputs(2611) <= not (a and b);
    layer4_outputs(2612) <= a and not b;
    layer4_outputs(2613) <= not (a or b);
    layer4_outputs(2614) <= not b;
    layer4_outputs(2615) <= not a;
    layer4_outputs(2616) <= not b or a;
    layer4_outputs(2617) <= a and not b;
    layer4_outputs(2618) <= not b or a;
    layer4_outputs(2619) <= a;
    layer4_outputs(2620) <= a;
    layer4_outputs(2621) <= not a;
    layer4_outputs(2622) <= not b;
    layer4_outputs(2623) <= not (a and b);
    layer4_outputs(2624) <= not a or b;
    layer4_outputs(2625) <= a and b;
    layer4_outputs(2626) <= '1';
    layer4_outputs(2627) <= a;
    layer4_outputs(2628) <= '0';
    layer4_outputs(2629) <= not b;
    layer4_outputs(2630) <= b and not a;
    layer4_outputs(2631) <= b;
    layer4_outputs(2632) <= not (a or b);
    layer4_outputs(2633) <= not b;
    layer4_outputs(2634) <= b and not a;
    layer4_outputs(2635) <= not a;
    layer4_outputs(2636) <= a and not b;
    layer4_outputs(2637) <= '0';
    layer4_outputs(2638) <= not (a and b);
    layer4_outputs(2639) <= '1';
    layer4_outputs(2640) <= not (a or b);
    layer4_outputs(2641) <= not (a and b);
    layer4_outputs(2642) <= a;
    layer4_outputs(2643) <= not (a or b);
    layer4_outputs(2644) <= not (a and b);
    layer4_outputs(2645) <= b and not a;
    layer4_outputs(2646) <= not (a or b);
    layer4_outputs(2647) <= not a;
    layer4_outputs(2648) <= not a or b;
    layer4_outputs(2649) <= a and not b;
    layer4_outputs(2650) <= '0';
    layer4_outputs(2651) <= not (a and b);
    layer4_outputs(2652) <= '0';
    layer4_outputs(2653) <= a or b;
    layer4_outputs(2654) <= a xor b;
    layer4_outputs(2655) <= a and b;
    layer4_outputs(2656) <= a or b;
    layer4_outputs(2657) <= not (a or b);
    layer4_outputs(2658) <= '0';
    layer4_outputs(2659) <= '1';
    layer4_outputs(2660) <= a or b;
    layer4_outputs(2661) <= not b or a;
    layer4_outputs(2662) <= not b;
    layer4_outputs(2663) <= not (a or b);
    layer4_outputs(2664) <= a and not b;
    layer4_outputs(2665) <= not b;
    layer4_outputs(2666) <= not a;
    layer4_outputs(2667) <= not (a or b);
    layer4_outputs(2668) <= not b or a;
    layer4_outputs(2669) <= not a;
    layer4_outputs(2670) <= not a or b;
    layer4_outputs(2671) <= a and not b;
    layer4_outputs(2672) <= '1';
    layer4_outputs(2673) <= a and not b;
    layer4_outputs(2674) <= '1';
    layer4_outputs(2675) <= '0';
    layer4_outputs(2676) <= b and not a;
    layer4_outputs(2677) <= not b or a;
    layer4_outputs(2678) <= not a;
    layer4_outputs(2679) <= not a;
    layer4_outputs(2680) <= not a;
    layer4_outputs(2681) <= b;
    layer4_outputs(2682) <= not (a and b);
    layer4_outputs(2683) <= a and not b;
    layer4_outputs(2684) <= not b or a;
    layer4_outputs(2685) <= not b;
    layer4_outputs(2686) <= a and not b;
    layer4_outputs(2687) <= not (a xor b);
    layer4_outputs(2688) <= not b or a;
    layer4_outputs(2689) <= b;
    layer4_outputs(2690) <= a and b;
    layer4_outputs(2691) <= a;
    layer4_outputs(2692) <= a;
    layer4_outputs(2693) <= a and b;
    layer4_outputs(2694) <= a and not b;
    layer4_outputs(2695) <= not a;
    layer4_outputs(2696) <= not (a xor b);
    layer4_outputs(2697) <= b;
    layer4_outputs(2698) <= b;
    layer4_outputs(2699) <= not (a or b);
    layer4_outputs(2700) <= not a or b;
    layer4_outputs(2701) <= b and not a;
    layer4_outputs(2702) <= not b;
    layer4_outputs(2703) <= not b;
    layer4_outputs(2704) <= b;
    layer4_outputs(2705) <= not a;
    layer4_outputs(2706) <= a and b;
    layer4_outputs(2707) <= not b;
    layer4_outputs(2708) <= a;
    layer4_outputs(2709) <= a and not b;
    layer4_outputs(2710) <= not a or b;
    layer4_outputs(2711) <= b;
    layer4_outputs(2712) <= a and not b;
    layer4_outputs(2713) <= a;
    layer4_outputs(2714) <= not a or b;
    layer4_outputs(2715) <= b;
    layer4_outputs(2716) <= '1';
    layer4_outputs(2717) <= b;
    layer4_outputs(2718) <= not b or a;
    layer4_outputs(2719) <= b;
    layer4_outputs(2720) <= not a;
    layer4_outputs(2721) <= not b;
    layer4_outputs(2722) <= not (a and b);
    layer4_outputs(2723) <= not a or b;
    layer4_outputs(2724) <= not b;
    layer4_outputs(2725) <= a and not b;
    layer4_outputs(2726) <= not a or b;
    layer4_outputs(2727) <= not (a or b);
    layer4_outputs(2728) <= '0';
    layer4_outputs(2729) <= a and not b;
    layer4_outputs(2730) <= not a;
    layer4_outputs(2731) <= '1';
    layer4_outputs(2732) <= '0';
    layer4_outputs(2733) <= not b or a;
    layer4_outputs(2734) <= b;
    layer4_outputs(2735) <= not (a or b);
    layer4_outputs(2736) <= not b or a;
    layer4_outputs(2737) <= not b or a;
    layer4_outputs(2738) <= '1';
    layer4_outputs(2739) <= a or b;
    layer4_outputs(2740) <= b and not a;
    layer4_outputs(2741) <= not b or a;
    layer4_outputs(2742) <= a and b;
    layer4_outputs(2743) <= not a or b;
    layer4_outputs(2744) <= not b or a;
    layer4_outputs(2745) <= not (a and b);
    layer4_outputs(2746) <= b and not a;
    layer4_outputs(2747) <= not b;
    layer4_outputs(2748) <= a xor b;
    layer4_outputs(2749) <= a or b;
    layer4_outputs(2750) <= a;
    layer4_outputs(2751) <= not a;
    layer4_outputs(2752) <= a;
    layer4_outputs(2753) <= '0';
    layer4_outputs(2754) <= '1';
    layer4_outputs(2755) <= a and b;
    layer4_outputs(2756) <= b;
    layer4_outputs(2757) <= a and not b;
    layer4_outputs(2758) <= a;
    layer4_outputs(2759) <= not a;
    layer4_outputs(2760) <= b;
    layer4_outputs(2761) <= not a;
    layer4_outputs(2762) <= not (a or b);
    layer4_outputs(2763) <= not a;
    layer4_outputs(2764) <= '0';
    layer4_outputs(2765) <= not b;
    layer4_outputs(2766) <= not b or a;
    layer4_outputs(2767) <= not b;
    layer4_outputs(2768) <= a or b;
    layer4_outputs(2769) <= a and not b;
    layer4_outputs(2770) <= a xor b;
    layer4_outputs(2771) <= b and not a;
    layer4_outputs(2772) <= a or b;
    layer4_outputs(2773) <= not (a or b);
    layer4_outputs(2774) <= '0';
    layer4_outputs(2775) <= '0';
    layer4_outputs(2776) <= a and not b;
    layer4_outputs(2777) <= not a;
    layer4_outputs(2778) <= not a;
    layer4_outputs(2779) <= not (a or b);
    layer4_outputs(2780) <= not (a or b);
    layer4_outputs(2781) <= b and not a;
    layer4_outputs(2782) <= not b or a;
    layer4_outputs(2783) <= not a;
    layer4_outputs(2784) <= not (a xor b);
    layer4_outputs(2785) <= b;
    layer4_outputs(2786) <= a and not b;
    layer4_outputs(2787) <= b and not a;
    layer4_outputs(2788) <= b;
    layer4_outputs(2789) <= not b or a;
    layer4_outputs(2790) <= a or b;
    layer4_outputs(2791) <= a and b;
    layer4_outputs(2792) <= not b;
    layer4_outputs(2793) <= not (a xor b);
    layer4_outputs(2794) <= a or b;
    layer4_outputs(2795) <= a;
    layer4_outputs(2796) <= not (a and b);
    layer4_outputs(2797) <= b and not a;
    layer4_outputs(2798) <= a;
    layer4_outputs(2799) <= a and b;
    layer4_outputs(2800) <= '0';
    layer4_outputs(2801) <= a or b;
    layer4_outputs(2802) <= a and b;
    layer4_outputs(2803) <= not b;
    layer4_outputs(2804) <= b;
    layer4_outputs(2805) <= b and not a;
    layer4_outputs(2806) <= b and not a;
    layer4_outputs(2807) <= a and b;
    layer4_outputs(2808) <= '1';
    layer4_outputs(2809) <= '1';
    layer4_outputs(2810) <= a or b;
    layer4_outputs(2811) <= a and not b;
    layer4_outputs(2812) <= a or b;
    layer4_outputs(2813) <= not (a and b);
    layer4_outputs(2814) <= not b or a;
    layer4_outputs(2815) <= not b;
    layer4_outputs(2816) <= '0';
    layer4_outputs(2817) <= a;
    layer4_outputs(2818) <= not a or b;
    layer4_outputs(2819) <= b;
    layer4_outputs(2820) <= not a;
    layer4_outputs(2821) <= not b;
    layer4_outputs(2822) <= not (a or b);
    layer4_outputs(2823) <= b;
    layer4_outputs(2824) <= not b or a;
    layer4_outputs(2825) <= '1';
    layer4_outputs(2826) <= '1';
    layer4_outputs(2827) <= not b or a;
    layer4_outputs(2828) <= '1';
    layer4_outputs(2829) <= a and not b;
    layer4_outputs(2830) <= b;
    layer4_outputs(2831) <= a and not b;
    layer4_outputs(2832) <= a or b;
    layer4_outputs(2833) <= a and not b;
    layer4_outputs(2834) <= a or b;
    layer4_outputs(2835) <= not (a or b);
    layer4_outputs(2836) <= b and not a;
    layer4_outputs(2837) <= '0';
    layer4_outputs(2838) <= b and not a;
    layer4_outputs(2839) <= b;
    layer4_outputs(2840) <= not b or a;
    layer4_outputs(2841) <= a;
    layer4_outputs(2842) <= a and b;
    layer4_outputs(2843) <= not (a or b);
    layer4_outputs(2844) <= '0';
    layer4_outputs(2845) <= a and b;
    layer4_outputs(2846) <= not b;
    layer4_outputs(2847) <= not b;
    layer4_outputs(2848) <= not (a or b);
    layer4_outputs(2849) <= not a;
    layer4_outputs(2850) <= not b;
    layer4_outputs(2851) <= not (a or b);
    layer4_outputs(2852) <= not b or a;
    layer4_outputs(2853) <= not a or b;
    layer4_outputs(2854) <= not b;
    layer4_outputs(2855) <= not b or a;
    layer4_outputs(2856) <= not b or a;
    layer4_outputs(2857) <= a or b;
    layer4_outputs(2858) <= a or b;
    layer4_outputs(2859) <= a;
    layer4_outputs(2860) <= '0';
    layer4_outputs(2861) <= a and b;
    layer4_outputs(2862) <= a and b;
    layer4_outputs(2863) <= not a or b;
    layer4_outputs(2864) <= not (a and b);
    layer4_outputs(2865) <= not b;
    layer4_outputs(2866) <= b;
    layer4_outputs(2867) <= not a or b;
    layer4_outputs(2868) <= not b or a;
    layer4_outputs(2869) <= not a or b;
    layer4_outputs(2870) <= '1';
    layer4_outputs(2871) <= not b;
    layer4_outputs(2872) <= '0';
    layer4_outputs(2873) <= a and not b;
    layer4_outputs(2874) <= not a;
    layer4_outputs(2875) <= a and not b;
    layer4_outputs(2876) <= a and b;
    layer4_outputs(2877) <= not (a and b);
    layer4_outputs(2878) <= a;
    layer4_outputs(2879) <= not b;
    layer4_outputs(2880) <= not (a or b);
    layer4_outputs(2881) <= '0';
    layer4_outputs(2882) <= b and not a;
    layer4_outputs(2883) <= a xor b;
    layer4_outputs(2884) <= not (a or b);
    layer4_outputs(2885) <= not (a xor b);
    layer4_outputs(2886) <= not a;
    layer4_outputs(2887) <= not a;
    layer4_outputs(2888) <= not a;
    layer4_outputs(2889) <= a xor b;
    layer4_outputs(2890) <= '1';
    layer4_outputs(2891) <= b and not a;
    layer4_outputs(2892) <= not a or b;
    layer4_outputs(2893) <= a or b;
    layer4_outputs(2894) <= not b or a;
    layer4_outputs(2895) <= a and not b;
    layer4_outputs(2896) <= a and b;
    layer4_outputs(2897) <= a or b;
    layer4_outputs(2898) <= '1';
    layer4_outputs(2899) <= not b or a;
    layer4_outputs(2900) <= b and not a;
    layer4_outputs(2901) <= not (a or b);
    layer4_outputs(2902) <= a;
    layer4_outputs(2903) <= not b;
    layer4_outputs(2904) <= b and not a;
    layer4_outputs(2905) <= not a or b;
    layer4_outputs(2906) <= '1';
    layer4_outputs(2907) <= '1';
    layer4_outputs(2908) <= not b;
    layer4_outputs(2909) <= b;
    layer4_outputs(2910) <= a and not b;
    layer4_outputs(2911) <= '1';
    layer4_outputs(2912) <= a and b;
    layer4_outputs(2913) <= not (a xor b);
    layer4_outputs(2914) <= a;
    layer4_outputs(2915) <= a;
    layer4_outputs(2916) <= a or b;
    layer4_outputs(2917) <= not (a or b);
    layer4_outputs(2918) <= not a;
    layer4_outputs(2919) <= not b;
    layer4_outputs(2920) <= not (a and b);
    layer4_outputs(2921) <= a xor b;
    layer4_outputs(2922) <= '1';
    layer4_outputs(2923) <= a and b;
    layer4_outputs(2924) <= a or b;
    layer4_outputs(2925) <= not b or a;
    layer4_outputs(2926) <= not (a and b);
    layer4_outputs(2927) <= '0';
    layer4_outputs(2928) <= not b or a;
    layer4_outputs(2929) <= a and b;
    layer4_outputs(2930) <= not (a or b);
    layer4_outputs(2931) <= not a or b;
    layer4_outputs(2932) <= a;
    layer4_outputs(2933) <= not a or b;
    layer4_outputs(2934) <= not b;
    layer4_outputs(2935) <= '0';
    layer4_outputs(2936) <= a or b;
    layer4_outputs(2937) <= not (a and b);
    layer4_outputs(2938) <= a or b;
    layer4_outputs(2939) <= '0';
    layer4_outputs(2940) <= a and b;
    layer4_outputs(2941) <= '0';
    layer4_outputs(2942) <= b and not a;
    layer4_outputs(2943) <= a and not b;
    layer4_outputs(2944) <= a and b;
    layer4_outputs(2945) <= b and not a;
    layer4_outputs(2946) <= a or b;
    layer4_outputs(2947) <= not a;
    layer4_outputs(2948) <= a and b;
    layer4_outputs(2949) <= '0';
    layer4_outputs(2950) <= b and not a;
    layer4_outputs(2951) <= not (a or b);
    layer4_outputs(2952) <= b;
    layer4_outputs(2953) <= b and not a;
    layer4_outputs(2954) <= not (a or b);
    layer4_outputs(2955) <= '0';
    layer4_outputs(2956) <= not a or b;
    layer4_outputs(2957) <= a or b;
    layer4_outputs(2958) <= not b;
    layer4_outputs(2959) <= '0';
    layer4_outputs(2960) <= not b;
    layer4_outputs(2961) <= not (a or b);
    layer4_outputs(2962) <= a or b;
    layer4_outputs(2963) <= a;
    layer4_outputs(2964) <= a and not b;
    layer4_outputs(2965) <= not b or a;
    layer4_outputs(2966) <= a and b;
    layer4_outputs(2967) <= b and not a;
    layer4_outputs(2968) <= b and not a;
    layer4_outputs(2969) <= a;
    layer4_outputs(2970) <= not a or b;
    layer4_outputs(2971) <= not b or a;
    layer4_outputs(2972) <= not b;
    layer4_outputs(2973) <= a;
    layer4_outputs(2974) <= not (a and b);
    layer4_outputs(2975) <= not (a or b);
    layer4_outputs(2976) <= not b or a;
    layer4_outputs(2977) <= a xor b;
    layer4_outputs(2978) <= not b;
    layer4_outputs(2979) <= b;
    layer4_outputs(2980) <= b;
    layer4_outputs(2981) <= not (a xor b);
    layer4_outputs(2982) <= not (a or b);
    layer4_outputs(2983) <= not (a xor b);
    layer4_outputs(2984) <= a and not b;
    layer4_outputs(2985) <= a or b;
    layer4_outputs(2986) <= a and not b;
    layer4_outputs(2987) <= not a or b;
    layer4_outputs(2988) <= not (a and b);
    layer4_outputs(2989) <= not (a or b);
    layer4_outputs(2990) <= b;
    layer4_outputs(2991) <= not (a or b);
    layer4_outputs(2992) <= not a;
    layer4_outputs(2993) <= not (a and b);
    layer4_outputs(2994) <= not a;
    layer4_outputs(2995) <= not b or a;
    layer4_outputs(2996) <= not a;
    layer4_outputs(2997) <= a or b;
    layer4_outputs(2998) <= not (a or b);
    layer4_outputs(2999) <= b and not a;
    layer4_outputs(3000) <= not b or a;
    layer4_outputs(3001) <= not a;
    layer4_outputs(3002) <= a and b;
    layer4_outputs(3003) <= b;
    layer4_outputs(3004) <= a;
    layer4_outputs(3005) <= not b;
    layer4_outputs(3006) <= a and not b;
    layer4_outputs(3007) <= not (a xor b);
    layer4_outputs(3008) <= a and b;
    layer4_outputs(3009) <= '1';
    layer4_outputs(3010) <= a and b;
    layer4_outputs(3011) <= not b;
    layer4_outputs(3012) <= not b or a;
    layer4_outputs(3013) <= a;
    layer4_outputs(3014) <= a or b;
    layer4_outputs(3015) <= b and not a;
    layer4_outputs(3016) <= a or b;
    layer4_outputs(3017) <= not (a or b);
    layer4_outputs(3018) <= not (a or b);
    layer4_outputs(3019) <= '0';
    layer4_outputs(3020) <= a;
    layer4_outputs(3021) <= not (a and b);
    layer4_outputs(3022) <= a or b;
    layer4_outputs(3023) <= '1';
    layer4_outputs(3024) <= a or b;
    layer4_outputs(3025) <= not (a and b);
    layer4_outputs(3026) <= a and b;
    layer4_outputs(3027) <= not (a or b);
    layer4_outputs(3028) <= a or b;
    layer4_outputs(3029) <= a xor b;
    layer4_outputs(3030) <= a or b;
    layer4_outputs(3031) <= a or b;
    layer4_outputs(3032) <= not b or a;
    layer4_outputs(3033) <= b and not a;
    layer4_outputs(3034) <= a or b;
    layer4_outputs(3035) <= not b;
    layer4_outputs(3036) <= a or b;
    layer4_outputs(3037) <= a and b;
    layer4_outputs(3038) <= a or b;
    layer4_outputs(3039) <= not b or a;
    layer4_outputs(3040) <= '0';
    layer4_outputs(3041) <= not a or b;
    layer4_outputs(3042) <= b;
    layer4_outputs(3043) <= a and not b;
    layer4_outputs(3044) <= not a or b;
    layer4_outputs(3045) <= not a;
    layer4_outputs(3046) <= not b;
    layer4_outputs(3047) <= not (a xor b);
    layer4_outputs(3048) <= not b;
    layer4_outputs(3049) <= not (a xor b);
    layer4_outputs(3050) <= b;
    layer4_outputs(3051) <= a or b;
    layer4_outputs(3052) <= a and b;
    layer4_outputs(3053) <= not b or a;
    layer4_outputs(3054) <= not a;
    layer4_outputs(3055) <= not b or a;
    layer4_outputs(3056) <= a and not b;
    layer4_outputs(3057) <= not b or a;
    layer4_outputs(3058) <= a and b;
    layer4_outputs(3059) <= not (a and b);
    layer4_outputs(3060) <= '1';
    layer4_outputs(3061) <= a;
    layer4_outputs(3062) <= a;
    layer4_outputs(3063) <= b and not a;
    layer4_outputs(3064) <= not b or a;
    layer4_outputs(3065) <= '0';
    layer4_outputs(3066) <= '1';
    layer4_outputs(3067) <= a and b;
    layer4_outputs(3068) <= b;
    layer4_outputs(3069) <= not a;
    layer4_outputs(3070) <= b;
    layer4_outputs(3071) <= not b;
    layer4_outputs(3072) <= not a;
    layer4_outputs(3073) <= '1';
    layer4_outputs(3074) <= a;
    layer4_outputs(3075) <= '0';
    layer4_outputs(3076) <= '0';
    layer4_outputs(3077) <= a and b;
    layer4_outputs(3078) <= a xor b;
    layer4_outputs(3079) <= not b or a;
    layer4_outputs(3080) <= a and b;
    layer4_outputs(3081) <= not a;
    layer4_outputs(3082) <= not a or b;
    layer4_outputs(3083) <= not b;
    layer4_outputs(3084) <= a or b;
    layer4_outputs(3085) <= not a;
    layer4_outputs(3086) <= a;
    layer4_outputs(3087) <= '0';
    layer4_outputs(3088) <= b and not a;
    layer4_outputs(3089) <= '0';
    layer4_outputs(3090) <= b and not a;
    layer4_outputs(3091) <= a and b;
    layer4_outputs(3092) <= '1';
    layer4_outputs(3093) <= not b;
    layer4_outputs(3094) <= a or b;
    layer4_outputs(3095) <= not a or b;
    layer4_outputs(3096) <= b and not a;
    layer4_outputs(3097) <= not a;
    layer4_outputs(3098) <= a and b;
    layer4_outputs(3099) <= a and not b;
    layer4_outputs(3100) <= not a;
    layer4_outputs(3101) <= not b or a;
    layer4_outputs(3102) <= b;
    layer4_outputs(3103) <= not a;
    layer4_outputs(3104) <= not a;
    layer4_outputs(3105) <= not (a and b);
    layer4_outputs(3106) <= not (a and b);
    layer4_outputs(3107) <= b and not a;
    layer4_outputs(3108) <= not (a or b);
    layer4_outputs(3109) <= not a;
    layer4_outputs(3110) <= a and b;
    layer4_outputs(3111) <= not a;
    layer4_outputs(3112) <= '1';
    layer4_outputs(3113) <= a or b;
    layer4_outputs(3114) <= a and b;
    layer4_outputs(3115) <= a and b;
    layer4_outputs(3116) <= not (a or b);
    layer4_outputs(3117) <= b;
    layer4_outputs(3118) <= not (a and b);
    layer4_outputs(3119) <= b;
    layer4_outputs(3120) <= a and b;
    layer4_outputs(3121) <= not a;
    layer4_outputs(3122) <= not (a and b);
    layer4_outputs(3123) <= not (a xor b);
    layer4_outputs(3124) <= not (a or b);
    layer4_outputs(3125) <= a;
    layer4_outputs(3126) <= a and not b;
    layer4_outputs(3127) <= '0';
    layer4_outputs(3128) <= '0';
    layer4_outputs(3129) <= a;
    layer4_outputs(3130) <= not b or a;
    layer4_outputs(3131) <= not a or b;
    layer4_outputs(3132) <= not a or b;
    layer4_outputs(3133) <= not b;
    layer4_outputs(3134) <= not (a or b);
    layer4_outputs(3135) <= a and b;
    layer4_outputs(3136) <= '0';
    layer4_outputs(3137) <= not a;
    layer4_outputs(3138) <= b and not a;
    layer4_outputs(3139) <= a xor b;
    layer4_outputs(3140) <= not b or a;
    layer4_outputs(3141) <= a or b;
    layer4_outputs(3142) <= not a;
    layer4_outputs(3143) <= a or b;
    layer4_outputs(3144) <= a and not b;
    layer4_outputs(3145) <= not (a or b);
    layer4_outputs(3146) <= not (a or b);
    layer4_outputs(3147) <= a and b;
    layer4_outputs(3148) <= a and not b;
    layer4_outputs(3149) <= '0';
    layer4_outputs(3150) <= b;
    layer4_outputs(3151) <= not (a and b);
    layer4_outputs(3152) <= b;
    layer4_outputs(3153) <= not (a and b);
    layer4_outputs(3154) <= a;
    layer4_outputs(3155) <= not a or b;
    layer4_outputs(3156) <= not (a and b);
    layer4_outputs(3157) <= not a or b;
    layer4_outputs(3158) <= b and not a;
    layer4_outputs(3159) <= not b;
    layer4_outputs(3160) <= not b;
    layer4_outputs(3161) <= b and not a;
    layer4_outputs(3162) <= a or b;
    layer4_outputs(3163) <= b and not a;
    layer4_outputs(3164) <= a and not b;
    layer4_outputs(3165) <= not a;
    layer4_outputs(3166) <= b;
    layer4_outputs(3167) <= not b or a;
    layer4_outputs(3168) <= b and not a;
    layer4_outputs(3169) <= a or b;
    layer4_outputs(3170) <= '1';
    layer4_outputs(3171) <= b;
    layer4_outputs(3172) <= not b;
    layer4_outputs(3173) <= b;
    layer4_outputs(3174) <= a and b;
    layer4_outputs(3175) <= b and not a;
    layer4_outputs(3176) <= not b or a;
    layer4_outputs(3177) <= not a;
    layer4_outputs(3178) <= not b or a;
    layer4_outputs(3179) <= not a or b;
    layer4_outputs(3180) <= a and not b;
    layer4_outputs(3181) <= b and not a;
    layer4_outputs(3182) <= not a or b;
    layer4_outputs(3183) <= a and b;
    layer4_outputs(3184) <= '1';
    layer4_outputs(3185) <= not b or a;
    layer4_outputs(3186) <= not b or a;
    layer4_outputs(3187) <= not b;
    layer4_outputs(3188) <= b and not a;
    layer4_outputs(3189) <= not a or b;
    layer4_outputs(3190) <= a and not b;
    layer4_outputs(3191) <= b and not a;
    layer4_outputs(3192) <= a or b;
    layer4_outputs(3193) <= a or b;
    layer4_outputs(3194) <= not (a or b);
    layer4_outputs(3195) <= b;
    layer4_outputs(3196) <= '1';
    layer4_outputs(3197) <= not b or a;
    layer4_outputs(3198) <= not b;
    layer4_outputs(3199) <= a and not b;
    layer4_outputs(3200) <= not a;
    layer4_outputs(3201) <= a and not b;
    layer4_outputs(3202) <= '1';
    layer4_outputs(3203) <= not b or a;
    layer4_outputs(3204) <= '0';
    layer4_outputs(3205) <= not (a and b);
    layer4_outputs(3206) <= not b or a;
    layer4_outputs(3207) <= a or b;
    layer4_outputs(3208) <= not b;
    layer4_outputs(3209) <= a or b;
    layer4_outputs(3210) <= not (a and b);
    layer4_outputs(3211) <= '1';
    layer4_outputs(3212) <= '0';
    layer4_outputs(3213) <= '0';
    layer4_outputs(3214) <= not b;
    layer4_outputs(3215) <= not b;
    layer4_outputs(3216) <= not a or b;
    layer4_outputs(3217) <= a or b;
    layer4_outputs(3218) <= not a;
    layer4_outputs(3219) <= not a or b;
    layer4_outputs(3220) <= a;
    layer4_outputs(3221) <= '0';
    layer4_outputs(3222) <= not a;
    layer4_outputs(3223) <= a and not b;
    layer4_outputs(3224) <= b;
    layer4_outputs(3225) <= a;
    layer4_outputs(3226) <= '1';
    layer4_outputs(3227) <= '0';
    layer4_outputs(3228) <= not a;
    layer4_outputs(3229) <= a and b;
    layer4_outputs(3230) <= not (a and b);
    layer4_outputs(3231) <= a and not b;
    layer4_outputs(3232) <= '0';
    layer4_outputs(3233) <= b and not a;
    layer4_outputs(3234) <= not (a and b);
    layer4_outputs(3235) <= not (a and b);
    layer4_outputs(3236) <= not (a and b);
    layer4_outputs(3237) <= not (a or b);
    layer4_outputs(3238) <= a and b;
    layer4_outputs(3239) <= not b or a;
    layer4_outputs(3240) <= not (a or b);
    layer4_outputs(3241) <= not a or b;
    layer4_outputs(3242) <= a;
    layer4_outputs(3243) <= a;
    layer4_outputs(3244) <= b and not a;
    layer4_outputs(3245) <= not a or b;
    layer4_outputs(3246) <= '0';
    layer4_outputs(3247) <= a;
    layer4_outputs(3248) <= a;
    layer4_outputs(3249) <= '0';
    layer4_outputs(3250) <= a;
    layer4_outputs(3251) <= a and not b;
    layer4_outputs(3252) <= '1';
    layer4_outputs(3253) <= not (a and b);
    layer4_outputs(3254) <= a;
    layer4_outputs(3255) <= not (a and b);
    layer4_outputs(3256) <= b and not a;
    layer4_outputs(3257) <= not b;
    layer4_outputs(3258) <= a or b;
    layer4_outputs(3259) <= not a;
    layer4_outputs(3260) <= b and not a;
    layer4_outputs(3261) <= '1';
    layer4_outputs(3262) <= not a;
    layer4_outputs(3263) <= a;
    layer4_outputs(3264) <= not a or b;
    layer4_outputs(3265) <= a and not b;
    layer4_outputs(3266) <= '1';
    layer4_outputs(3267) <= '0';
    layer4_outputs(3268) <= a xor b;
    layer4_outputs(3269) <= b;
    layer4_outputs(3270) <= not (a and b);
    layer4_outputs(3271) <= '1';
    layer4_outputs(3272) <= a;
    layer4_outputs(3273) <= b and not a;
    layer4_outputs(3274) <= b and not a;
    layer4_outputs(3275) <= a and b;
    layer4_outputs(3276) <= not b;
    layer4_outputs(3277) <= '1';
    layer4_outputs(3278) <= a or b;
    layer4_outputs(3279) <= not b;
    layer4_outputs(3280) <= not b or a;
    layer4_outputs(3281) <= a or b;
    layer4_outputs(3282) <= '1';
    layer4_outputs(3283) <= b;
    layer4_outputs(3284) <= a;
    layer4_outputs(3285) <= not b or a;
    layer4_outputs(3286) <= not b;
    layer4_outputs(3287) <= a and not b;
    layer4_outputs(3288) <= not b or a;
    layer4_outputs(3289) <= not (a and b);
    layer4_outputs(3290) <= not (a or b);
    layer4_outputs(3291) <= b;
    layer4_outputs(3292) <= a;
    layer4_outputs(3293) <= not b or a;
    layer4_outputs(3294) <= not a;
    layer4_outputs(3295) <= not a;
    layer4_outputs(3296) <= b;
    layer4_outputs(3297) <= a and not b;
    layer4_outputs(3298) <= not b;
    layer4_outputs(3299) <= a and b;
    layer4_outputs(3300) <= a and b;
    layer4_outputs(3301) <= a and b;
    layer4_outputs(3302) <= a and not b;
    layer4_outputs(3303) <= not b;
    layer4_outputs(3304) <= not b;
    layer4_outputs(3305) <= '1';
    layer4_outputs(3306) <= not (a xor b);
    layer4_outputs(3307) <= not b;
    layer4_outputs(3308) <= not (a and b);
    layer4_outputs(3309) <= b and not a;
    layer4_outputs(3310) <= a and not b;
    layer4_outputs(3311) <= a and not b;
    layer4_outputs(3312) <= a and b;
    layer4_outputs(3313) <= b and not a;
    layer4_outputs(3314) <= not a or b;
    layer4_outputs(3315) <= not a;
    layer4_outputs(3316) <= a;
    layer4_outputs(3317) <= not a or b;
    layer4_outputs(3318) <= not b or a;
    layer4_outputs(3319) <= b;
    layer4_outputs(3320) <= a and b;
    layer4_outputs(3321) <= b and not a;
    layer4_outputs(3322) <= not (a xor b);
    layer4_outputs(3323) <= not a or b;
    layer4_outputs(3324) <= not a or b;
    layer4_outputs(3325) <= a or b;
    layer4_outputs(3326) <= not b;
    layer4_outputs(3327) <= a;
    layer4_outputs(3328) <= not b;
    layer4_outputs(3329) <= '1';
    layer4_outputs(3330) <= a xor b;
    layer4_outputs(3331) <= a and b;
    layer4_outputs(3332) <= not b;
    layer4_outputs(3333) <= a or b;
    layer4_outputs(3334) <= a and b;
    layer4_outputs(3335) <= a xor b;
    layer4_outputs(3336) <= '1';
    layer4_outputs(3337) <= not b;
    layer4_outputs(3338) <= not a;
    layer4_outputs(3339) <= '1';
    layer4_outputs(3340) <= b and not a;
    layer4_outputs(3341) <= a or b;
    layer4_outputs(3342) <= not b or a;
    layer4_outputs(3343) <= not a or b;
    layer4_outputs(3344) <= not b;
    layer4_outputs(3345) <= '1';
    layer4_outputs(3346) <= b and not a;
    layer4_outputs(3347) <= b and not a;
    layer4_outputs(3348) <= not (a or b);
    layer4_outputs(3349) <= a xor b;
    layer4_outputs(3350) <= '1';
    layer4_outputs(3351) <= a xor b;
    layer4_outputs(3352) <= b and not a;
    layer4_outputs(3353) <= not (a xor b);
    layer4_outputs(3354) <= not (a xor b);
    layer4_outputs(3355) <= not (a and b);
    layer4_outputs(3356) <= b;
    layer4_outputs(3357) <= '0';
    layer4_outputs(3358) <= a or b;
    layer4_outputs(3359) <= not a;
    layer4_outputs(3360) <= b;
    layer4_outputs(3361) <= not a;
    layer4_outputs(3362) <= not a or b;
    layer4_outputs(3363) <= a and not b;
    layer4_outputs(3364) <= a;
    layer4_outputs(3365) <= not (a or b);
    layer4_outputs(3366) <= b and not a;
    layer4_outputs(3367) <= not a;
    layer4_outputs(3368) <= '0';
    layer4_outputs(3369) <= a and not b;
    layer4_outputs(3370) <= b and not a;
    layer4_outputs(3371) <= a or b;
    layer4_outputs(3372) <= not a or b;
    layer4_outputs(3373) <= not b;
    layer4_outputs(3374) <= a;
    layer4_outputs(3375) <= '1';
    layer4_outputs(3376) <= a and not b;
    layer4_outputs(3377) <= b;
    layer4_outputs(3378) <= not b;
    layer4_outputs(3379) <= not a;
    layer4_outputs(3380) <= not (a or b);
    layer4_outputs(3381) <= not (a and b);
    layer4_outputs(3382) <= not a;
    layer4_outputs(3383) <= a and not b;
    layer4_outputs(3384) <= a;
    layer4_outputs(3385) <= not (a xor b);
    layer4_outputs(3386) <= '1';
    layer4_outputs(3387) <= not a or b;
    layer4_outputs(3388) <= '0';
    layer4_outputs(3389) <= not (a and b);
    layer4_outputs(3390) <= '1';
    layer4_outputs(3391) <= not a;
    layer4_outputs(3392) <= b;
    layer4_outputs(3393) <= a and not b;
    layer4_outputs(3394) <= '1';
    layer4_outputs(3395) <= b and not a;
    layer4_outputs(3396) <= a and b;
    layer4_outputs(3397) <= a and not b;
    layer4_outputs(3398) <= a;
    layer4_outputs(3399) <= a and not b;
    layer4_outputs(3400) <= a and b;
    layer4_outputs(3401) <= not b;
    layer4_outputs(3402) <= not b;
    layer4_outputs(3403) <= a;
    layer4_outputs(3404) <= '0';
    layer4_outputs(3405) <= not (a and b);
    layer4_outputs(3406) <= not b or a;
    layer4_outputs(3407) <= '1';
    layer4_outputs(3408) <= not (a or b);
    layer4_outputs(3409) <= not b or a;
    layer4_outputs(3410) <= a;
    layer4_outputs(3411) <= '1';
    layer4_outputs(3412) <= b and not a;
    layer4_outputs(3413) <= not (a xor b);
    layer4_outputs(3414) <= not a;
    layer4_outputs(3415) <= not (a or b);
    layer4_outputs(3416) <= not b;
    layer4_outputs(3417) <= not b;
    layer4_outputs(3418) <= a and not b;
    layer4_outputs(3419) <= a and not b;
    layer4_outputs(3420) <= '1';
    layer4_outputs(3421) <= b and not a;
    layer4_outputs(3422) <= '0';
    layer4_outputs(3423) <= a and not b;
    layer4_outputs(3424) <= a;
    layer4_outputs(3425) <= not (a xor b);
    layer4_outputs(3426) <= a and b;
    layer4_outputs(3427) <= not b or a;
    layer4_outputs(3428) <= a and not b;
    layer4_outputs(3429) <= not a or b;
    layer4_outputs(3430) <= not a or b;
    layer4_outputs(3431) <= a and not b;
    layer4_outputs(3432) <= a;
    layer4_outputs(3433) <= a and b;
    layer4_outputs(3434) <= b;
    layer4_outputs(3435) <= not a;
    layer4_outputs(3436) <= b;
    layer4_outputs(3437) <= not (a xor b);
    layer4_outputs(3438) <= '0';
    layer4_outputs(3439) <= not a;
    layer4_outputs(3440) <= '1';
    layer4_outputs(3441) <= '1';
    layer4_outputs(3442) <= not b or a;
    layer4_outputs(3443) <= a or b;
    layer4_outputs(3444) <= a or b;
    layer4_outputs(3445) <= b;
    layer4_outputs(3446) <= b and not a;
    layer4_outputs(3447) <= not (a or b);
    layer4_outputs(3448) <= b;
    layer4_outputs(3449) <= a;
    layer4_outputs(3450) <= not (a xor b);
    layer4_outputs(3451) <= a or b;
    layer4_outputs(3452) <= not a;
    layer4_outputs(3453) <= not b;
    layer4_outputs(3454) <= a and b;
    layer4_outputs(3455) <= '1';
    layer4_outputs(3456) <= a and not b;
    layer4_outputs(3457) <= a and not b;
    layer4_outputs(3458) <= a;
    layer4_outputs(3459) <= not a or b;
    layer4_outputs(3460) <= not a;
    layer4_outputs(3461) <= not a;
    layer4_outputs(3462) <= b;
    layer4_outputs(3463) <= a and b;
    layer4_outputs(3464) <= not (a or b);
    layer4_outputs(3465) <= not (a and b);
    layer4_outputs(3466) <= not (a xor b);
    layer4_outputs(3467) <= b;
    layer4_outputs(3468) <= b;
    layer4_outputs(3469) <= not b;
    layer4_outputs(3470) <= not (a xor b);
    layer4_outputs(3471) <= not a;
    layer4_outputs(3472) <= a and b;
    layer4_outputs(3473) <= b and not a;
    layer4_outputs(3474) <= b;
    layer4_outputs(3475) <= a;
    layer4_outputs(3476) <= b and not a;
    layer4_outputs(3477) <= '1';
    layer4_outputs(3478) <= a or b;
    layer4_outputs(3479) <= not (a and b);
    layer4_outputs(3480) <= a;
    layer4_outputs(3481) <= not a or b;
    layer4_outputs(3482) <= not (a or b);
    layer4_outputs(3483) <= not (a or b);
    layer4_outputs(3484) <= not (a and b);
    layer4_outputs(3485) <= not a or b;
    layer4_outputs(3486) <= a;
    layer4_outputs(3487) <= not a or b;
    layer4_outputs(3488) <= not (a or b);
    layer4_outputs(3489) <= not a or b;
    layer4_outputs(3490) <= a;
    layer4_outputs(3491) <= '0';
    layer4_outputs(3492) <= not a or b;
    layer4_outputs(3493) <= a;
    layer4_outputs(3494) <= not b or a;
    layer4_outputs(3495) <= a and b;
    layer4_outputs(3496) <= a and b;
    layer4_outputs(3497) <= '1';
    layer4_outputs(3498) <= '0';
    layer4_outputs(3499) <= not a or b;
    layer4_outputs(3500) <= b and not a;
    layer4_outputs(3501) <= not b or a;
    layer4_outputs(3502) <= '0';
    layer4_outputs(3503) <= b;
    layer4_outputs(3504) <= not a or b;
    layer4_outputs(3505) <= a or b;
    layer4_outputs(3506) <= not a or b;
    layer4_outputs(3507) <= not (a xor b);
    layer4_outputs(3508) <= a xor b;
    layer4_outputs(3509) <= not b;
    layer4_outputs(3510) <= not (a xor b);
    layer4_outputs(3511) <= b;
    layer4_outputs(3512) <= not a;
    layer4_outputs(3513) <= not a or b;
    layer4_outputs(3514) <= not (a or b);
    layer4_outputs(3515) <= not b;
    layer4_outputs(3516) <= a;
    layer4_outputs(3517) <= a or b;
    layer4_outputs(3518) <= not b;
    layer4_outputs(3519) <= not a;
    layer4_outputs(3520) <= not (a and b);
    layer4_outputs(3521) <= not a;
    layer4_outputs(3522) <= not a or b;
    layer4_outputs(3523) <= a and b;
    layer4_outputs(3524) <= not b or a;
    layer4_outputs(3525) <= not b;
    layer4_outputs(3526) <= '0';
    layer4_outputs(3527) <= not (a or b);
    layer4_outputs(3528) <= a and not b;
    layer4_outputs(3529) <= b;
    layer4_outputs(3530) <= not a;
    layer4_outputs(3531) <= not b;
    layer4_outputs(3532) <= not a or b;
    layer4_outputs(3533) <= b;
    layer4_outputs(3534) <= not (a xor b);
    layer4_outputs(3535) <= a or b;
    layer4_outputs(3536) <= a;
    layer4_outputs(3537) <= a and not b;
    layer4_outputs(3538) <= a and not b;
    layer4_outputs(3539) <= not b or a;
    layer4_outputs(3540) <= b;
    layer4_outputs(3541) <= not a;
    layer4_outputs(3542) <= a and b;
    layer4_outputs(3543) <= '1';
    layer4_outputs(3544) <= '0';
    layer4_outputs(3545) <= '1';
    layer4_outputs(3546) <= not (a or b);
    layer4_outputs(3547) <= a and not b;
    layer4_outputs(3548) <= not (a and b);
    layer4_outputs(3549) <= b and not a;
    layer4_outputs(3550) <= a or b;
    layer4_outputs(3551) <= not b or a;
    layer4_outputs(3552) <= a xor b;
    layer4_outputs(3553) <= not a;
    layer4_outputs(3554) <= b;
    layer4_outputs(3555) <= a and not b;
    layer4_outputs(3556) <= a and b;
    layer4_outputs(3557) <= a or b;
    layer4_outputs(3558) <= not a;
    layer4_outputs(3559) <= not (a xor b);
    layer4_outputs(3560) <= not (a xor b);
    layer4_outputs(3561) <= a and b;
    layer4_outputs(3562) <= not a;
    layer4_outputs(3563) <= not a or b;
    layer4_outputs(3564) <= not b or a;
    layer4_outputs(3565) <= not (a or b);
    layer4_outputs(3566) <= not a or b;
    layer4_outputs(3567) <= not a;
    layer4_outputs(3568) <= '0';
    layer4_outputs(3569) <= b and not a;
    layer4_outputs(3570) <= a and b;
    layer4_outputs(3571) <= b and not a;
    layer4_outputs(3572) <= '0';
    layer4_outputs(3573) <= '1';
    layer4_outputs(3574) <= b;
    layer4_outputs(3575) <= not (a and b);
    layer4_outputs(3576) <= not a;
    layer4_outputs(3577) <= a and not b;
    layer4_outputs(3578) <= not (a and b);
    layer4_outputs(3579) <= not b;
    layer4_outputs(3580) <= a and not b;
    layer4_outputs(3581) <= '0';
    layer4_outputs(3582) <= b;
    layer4_outputs(3583) <= b;
    layer4_outputs(3584) <= not a;
    layer4_outputs(3585) <= a;
    layer4_outputs(3586) <= b;
    layer4_outputs(3587) <= not a or b;
    layer4_outputs(3588) <= a or b;
    layer4_outputs(3589) <= a;
    layer4_outputs(3590) <= not b or a;
    layer4_outputs(3591) <= '1';
    layer4_outputs(3592) <= not b or a;
    layer4_outputs(3593) <= not (a or b);
    layer4_outputs(3594) <= a;
    layer4_outputs(3595) <= '1';
    layer4_outputs(3596) <= a and b;
    layer4_outputs(3597) <= not b or a;
    layer4_outputs(3598) <= not b;
    layer4_outputs(3599) <= a;
    layer4_outputs(3600) <= not (a xor b);
    layer4_outputs(3601) <= b;
    layer4_outputs(3602) <= '1';
    layer4_outputs(3603) <= a;
    layer4_outputs(3604) <= a and not b;
    layer4_outputs(3605) <= b;
    layer4_outputs(3606) <= a or b;
    layer4_outputs(3607) <= not a;
    layer4_outputs(3608) <= not (a or b);
    layer4_outputs(3609) <= '0';
    layer4_outputs(3610) <= a;
    layer4_outputs(3611) <= '1';
    layer4_outputs(3612) <= b and not a;
    layer4_outputs(3613) <= not a or b;
    layer4_outputs(3614) <= not b;
    layer4_outputs(3615) <= not b;
    layer4_outputs(3616) <= not a or b;
    layer4_outputs(3617) <= not a;
    layer4_outputs(3618) <= a and not b;
    layer4_outputs(3619) <= a and b;
    layer4_outputs(3620) <= '0';
    layer4_outputs(3621) <= not b or a;
    layer4_outputs(3622) <= not a or b;
    layer4_outputs(3623) <= b and not a;
    layer4_outputs(3624) <= not a;
    layer4_outputs(3625) <= a;
    layer4_outputs(3626) <= not a or b;
    layer4_outputs(3627) <= a;
    layer4_outputs(3628) <= b;
    layer4_outputs(3629) <= not (a or b);
    layer4_outputs(3630) <= not a or b;
    layer4_outputs(3631) <= not (a or b);
    layer4_outputs(3632) <= a and not b;
    layer4_outputs(3633) <= a and b;
    layer4_outputs(3634) <= not b;
    layer4_outputs(3635) <= a and b;
    layer4_outputs(3636) <= not (a or b);
    layer4_outputs(3637) <= not a or b;
    layer4_outputs(3638) <= a and not b;
    layer4_outputs(3639) <= a or b;
    layer4_outputs(3640) <= not b or a;
    layer4_outputs(3641) <= not (a and b);
    layer4_outputs(3642) <= a;
    layer4_outputs(3643) <= b and not a;
    layer4_outputs(3644) <= a;
    layer4_outputs(3645) <= a xor b;
    layer4_outputs(3646) <= not a;
    layer4_outputs(3647) <= '0';
    layer4_outputs(3648) <= a and b;
    layer4_outputs(3649) <= not b or a;
    layer4_outputs(3650) <= a and not b;
    layer4_outputs(3651) <= not a;
    layer4_outputs(3652) <= not a;
    layer4_outputs(3653) <= not (a and b);
    layer4_outputs(3654) <= b and not a;
    layer4_outputs(3655) <= a and not b;
    layer4_outputs(3656) <= not (a and b);
    layer4_outputs(3657) <= '0';
    layer4_outputs(3658) <= b;
    layer4_outputs(3659) <= a;
    layer4_outputs(3660) <= b;
    layer4_outputs(3661) <= a or b;
    layer4_outputs(3662) <= b and not a;
    layer4_outputs(3663) <= '0';
    layer4_outputs(3664) <= not (a or b);
    layer4_outputs(3665) <= '0';
    layer4_outputs(3666) <= not b or a;
    layer4_outputs(3667) <= not (a xor b);
    layer4_outputs(3668) <= not a or b;
    layer4_outputs(3669) <= not (a and b);
    layer4_outputs(3670) <= not b or a;
    layer4_outputs(3671) <= '0';
    layer4_outputs(3672) <= b;
    layer4_outputs(3673) <= not b or a;
    layer4_outputs(3674) <= '1';
    layer4_outputs(3675) <= '1';
    layer4_outputs(3676) <= not b or a;
    layer4_outputs(3677) <= a xor b;
    layer4_outputs(3678) <= '1';
    layer4_outputs(3679) <= b and not a;
    layer4_outputs(3680) <= not (a and b);
    layer4_outputs(3681) <= not a;
    layer4_outputs(3682) <= not b;
    layer4_outputs(3683) <= b and not a;
    layer4_outputs(3684) <= b;
    layer4_outputs(3685) <= not b or a;
    layer4_outputs(3686) <= not b;
    layer4_outputs(3687) <= not b or a;
    layer4_outputs(3688) <= not b;
    layer4_outputs(3689) <= '1';
    layer4_outputs(3690) <= a and b;
    layer4_outputs(3691) <= not (a and b);
    layer4_outputs(3692) <= not a;
    layer4_outputs(3693) <= '1';
    layer4_outputs(3694) <= a;
    layer4_outputs(3695) <= a and b;
    layer4_outputs(3696) <= a and not b;
    layer4_outputs(3697) <= b and not a;
    layer4_outputs(3698) <= not a;
    layer4_outputs(3699) <= b and not a;
    layer4_outputs(3700) <= a xor b;
    layer4_outputs(3701) <= not b;
    layer4_outputs(3702) <= b and not a;
    layer4_outputs(3703) <= not b;
    layer4_outputs(3704) <= not a;
    layer4_outputs(3705) <= not a or b;
    layer4_outputs(3706) <= a and b;
    layer4_outputs(3707) <= a or b;
    layer4_outputs(3708) <= a and b;
    layer4_outputs(3709) <= b and not a;
    layer4_outputs(3710) <= '1';
    layer4_outputs(3711) <= a;
    layer4_outputs(3712) <= not (a xor b);
    layer4_outputs(3713) <= a;
    layer4_outputs(3714) <= not a;
    layer4_outputs(3715) <= '0';
    layer4_outputs(3716) <= a and b;
    layer4_outputs(3717) <= b and not a;
    layer4_outputs(3718) <= a and b;
    layer4_outputs(3719) <= not b;
    layer4_outputs(3720) <= '0';
    layer4_outputs(3721) <= a and b;
    layer4_outputs(3722) <= a and not b;
    layer4_outputs(3723) <= a and b;
    layer4_outputs(3724) <= not (a or b);
    layer4_outputs(3725) <= a or b;
    layer4_outputs(3726) <= '0';
    layer4_outputs(3727) <= not b or a;
    layer4_outputs(3728) <= a;
    layer4_outputs(3729) <= a;
    layer4_outputs(3730) <= not a or b;
    layer4_outputs(3731) <= a and not b;
    layer4_outputs(3732) <= b and not a;
    layer4_outputs(3733) <= a and b;
    layer4_outputs(3734) <= not (a xor b);
    layer4_outputs(3735) <= a or b;
    layer4_outputs(3736) <= b and not a;
    layer4_outputs(3737) <= b;
    layer4_outputs(3738) <= '0';
    layer4_outputs(3739) <= not (a and b);
    layer4_outputs(3740) <= b and not a;
    layer4_outputs(3741) <= '1';
    layer4_outputs(3742) <= not (a and b);
    layer4_outputs(3743) <= not a or b;
    layer4_outputs(3744) <= a;
    layer4_outputs(3745) <= not b or a;
    layer4_outputs(3746) <= a or b;
    layer4_outputs(3747) <= not b;
    layer4_outputs(3748) <= not a;
    layer4_outputs(3749) <= not b;
    layer4_outputs(3750) <= b;
    layer4_outputs(3751) <= b;
    layer4_outputs(3752) <= not (a and b);
    layer4_outputs(3753) <= '0';
    layer4_outputs(3754) <= b and not a;
    layer4_outputs(3755) <= a or b;
    layer4_outputs(3756) <= not a;
    layer4_outputs(3757) <= b and not a;
    layer4_outputs(3758) <= b;
    layer4_outputs(3759) <= not a or b;
    layer4_outputs(3760) <= '0';
    layer4_outputs(3761) <= not b;
    layer4_outputs(3762) <= b;
    layer4_outputs(3763) <= not (a xor b);
    layer4_outputs(3764) <= not (a or b);
    layer4_outputs(3765) <= not b;
    layer4_outputs(3766) <= not a or b;
    layer4_outputs(3767) <= not b or a;
    layer4_outputs(3768) <= a xor b;
    layer4_outputs(3769) <= not a or b;
    layer4_outputs(3770) <= not (a or b);
    layer4_outputs(3771) <= not (a xor b);
    layer4_outputs(3772) <= a and not b;
    layer4_outputs(3773) <= '1';
    layer4_outputs(3774) <= a and not b;
    layer4_outputs(3775) <= a;
    layer4_outputs(3776) <= b;
    layer4_outputs(3777) <= a;
    layer4_outputs(3778) <= not (a xor b);
    layer4_outputs(3779) <= not b or a;
    layer4_outputs(3780) <= not a or b;
    layer4_outputs(3781) <= b;
    layer4_outputs(3782) <= not a or b;
    layer4_outputs(3783) <= not b;
    layer4_outputs(3784) <= not a;
    layer4_outputs(3785) <= not (a or b);
    layer4_outputs(3786) <= not a;
    layer4_outputs(3787) <= not (a and b);
    layer4_outputs(3788) <= a and b;
    layer4_outputs(3789) <= a or b;
    layer4_outputs(3790) <= not b or a;
    layer4_outputs(3791) <= a or b;
    layer4_outputs(3792) <= a and b;
    layer4_outputs(3793) <= a and not b;
    layer4_outputs(3794) <= '1';
    layer4_outputs(3795) <= b and not a;
    layer4_outputs(3796) <= a and not b;
    layer4_outputs(3797) <= not (a and b);
    layer4_outputs(3798) <= b;
    layer4_outputs(3799) <= not (a and b);
    layer4_outputs(3800) <= a;
    layer4_outputs(3801) <= b;
    layer4_outputs(3802) <= not b or a;
    layer4_outputs(3803) <= b;
    layer4_outputs(3804) <= b and not a;
    layer4_outputs(3805) <= '1';
    layer4_outputs(3806) <= b;
    layer4_outputs(3807) <= b;
    layer4_outputs(3808) <= b;
    layer4_outputs(3809) <= not (a or b);
    layer4_outputs(3810) <= not (a and b);
    layer4_outputs(3811) <= not a or b;
    layer4_outputs(3812) <= not b;
    layer4_outputs(3813) <= not (a and b);
    layer4_outputs(3814) <= not (a and b);
    layer4_outputs(3815) <= a and b;
    layer4_outputs(3816) <= not a;
    layer4_outputs(3817) <= not b or a;
    layer4_outputs(3818) <= b and not a;
    layer4_outputs(3819) <= not (a xor b);
    layer4_outputs(3820) <= not a or b;
    layer4_outputs(3821) <= not b or a;
    layer4_outputs(3822) <= not a;
    layer4_outputs(3823) <= not a or b;
    layer4_outputs(3824) <= a and not b;
    layer4_outputs(3825) <= a xor b;
    layer4_outputs(3826) <= a and not b;
    layer4_outputs(3827) <= a;
    layer4_outputs(3828) <= a and b;
    layer4_outputs(3829) <= not (a and b);
    layer4_outputs(3830) <= a;
    layer4_outputs(3831) <= b;
    layer4_outputs(3832) <= not (a or b);
    layer4_outputs(3833) <= not (a or b);
    layer4_outputs(3834) <= b and not a;
    layer4_outputs(3835) <= a;
    layer4_outputs(3836) <= '0';
    layer4_outputs(3837) <= '1';
    layer4_outputs(3838) <= '0';
    layer4_outputs(3839) <= not (a and b);
    layer4_outputs(3840) <= '0';
    layer4_outputs(3841) <= not (a and b);
    layer4_outputs(3842) <= a xor b;
    layer4_outputs(3843) <= b;
    layer4_outputs(3844) <= b and not a;
    layer4_outputs(3845) <= b and not a;
    layer4_outputs(3846) <= a or b;
    layer4_outputs(3847) <= not a or b;
    layer4_outputs(3848) <= not a;
    layer4_outputs(3849) <= a;
    layer4_outputs(3850) <= '1';
    layer4_outputs(3851) <= a;
    layer4_outputs(3852) <= not a or b;
    layer4_outputs(3853) <= b and not a;
    layer4_outputs(3854) <= a and not b;
    layer4_outputs(3855) <= not b;
    layer4_outputs(3856) <= not (a or b);
    layer4_outputs(3857) <= a and not b;
    layer4_outputs(3858) <= not (a and b);
    layer4_outputs(3859) <= not a;
    layer4_outputs(3860) <= b and not a;
    layer4_outputs(3861) <= not b or a;
    layer4_outputs(3862) <= a;
    layer4_outputs(3863) <= not b or a;
    layer4_outputs(3864) <= not (a or b);
    layer4_outputs(3865) <= a;
    layer4_outputs(3866) <= '0';
    layer4_outputs(3867) <= not b or a;
    layer4_outputs(3868) <= a or b;
    layer4_outputs(3869) <= a and b;
    layer4_outputs(3870) <= not b;
    layer4_outputs(3871) <= not (a or b);
    layer4_outputs(3872) <= not (a and b);
    layer4_outputs(3873) <= a and not b;
    layer4_outputs(3874) <= not b or a;
    layer4_outputs(3875) <= a and b;
    layer4_outputs(3876) <= '1';
    layer4_outputs(3877) <= not b;
    layer4_outputs(3878) <= not (a and b);
    layer4_outputs(3879) <= not b or a;
    layer4_outputs(3880) <= a and not b;
    layer4_outputs(3881) <= b;
    layer4_outputs(3882) <= b;
    layer4_outputs(3883) <= a and not b;
    layer4_outputs(3884) <= a or b;
    layer4_outputs(3885) <= a and not b;
    layer4_outputs(3886) <= not (a and b);
    layer4_outputs(3887) <= not a or b;
    layer4_outputs(3888) <= a or b;
    layer4_outputs(3889) <= not (a and b);
    layer4_outputs(3890) <= b and not a;
    layer4_outputs(3891) <= not b or a;
    layer4_outputs(3892) <= b;
    layer4_outputs(3893) <= a and b;
    layer4_outputs(3894) <= '0';
    layer4_outputs(3895) <= not b;
    layer4_outputs(3896) <= '1';
    layer4_outputs(3897) <= '1';
    layer4_outputs(3898) <= not b or a;
    layer4_outputs(3899) <= a or b;
    layer4_outputs(3900) <= b and not a;
    layer4_outputs(3901) <= not (a xor b);
    layer4_outputs(3902) <= '1';
    layer4_outputs(3903) <= a;
    layer4_outputs(3904) <= not b;
    layer4_outputs(3905) <= not (a or b);
    layer4_outputs(3906) <= a;
    layer4_outputs(3907) <= not a;
    layer4_outputs(3908) <= not b;
    layer4_outputs(3909) <= a or b;
    layer4_outputs(3910) <= '1';
    layer4_outputs(3911) <= a and not b;
    layer4_outputs(3912) <= not b;
    layer4_outputs(3913) <= b;
    layer4_outputs(3914) <= not (a or b);
    layer4_outputs(3915) <= not a;
    layer4_outputs(3916) <= b and not a;
    layer4_outputs(3917) <= a;
    layer4_outputs(3918) <= not b or a;
    layer4_outputs(3919) <= not a;
    layer4_outputs(3920) <= a;
    layer4_outputs(3921) <= not b or a;
    layer4_outputs(3922) <= not b or a;
    layer4_outputs(3923) <= not a;
    layer4_outputs(3924) <= not b or a;
    layer4_outputs(3925) <= '1';
    layer4_outputs(3926) <= not b;
    layer4_outputs(3927) <= not b or a;
    layer4_outputs(3928) <= not (a xor b);
    layer4_outputs(3929) <= not b;
    layer4_outputs(3930) <= a xor b;
    layer4_outputs(3931) <= a and not b;
    layer4_outputs(3932) <= a and not b;
    layer4_outputs(3933) <= a and not b;
    layer4_outputs(3934) <= not a or b;
    layer4_outputs(3935) <= a xor b;
    layer4_outputs(3936) <= not a;
    layer4_outputs(3937) <= not b or a;
    layer4_outputs(3938) <= '0';
    layer4_outputs(3939) <= b;
    layer4_outputs(3940) <= a and b;
    layer4_outputs(3941) <= not b;
    layer4_outputs(3942) <= a and b;
    layer4_outputs(3943) <= not b or a;
    layer4_outputs(3944) <= b and not a;
    layer4_outputs(3945) <= a and b;
    layer4_outputs(3946) <= a or b;
    layer4_outputs(3947) <= not a or b;
    layer4_outputs(3948) <= not (a and b);
    layer4_outputs(3949) <= not a;
    layer4_outputs(3950) <= not (a or b);
    layer4_outputs(3951) <= a xor b;
    layer4_outputs(3952) <= b;
    layer4_outputs(3953) <= a and not b;
    layer4_outputs(3954) <= b;
    layer4_outputs(3955) <= not (a and b);
    layer4_outputs(3956) <= a and b;
    layer4_outputs(3957) <= not b;
    layer4_outputs(3958) <= a xor b;
    layer4_outputs(3959) <= not a;
    layer4_outputs(3960) <= not (a and b);
    layer4_outputs(3961) <= '0';
    layer4_outputs(3962) <= not a or b;
    layer4_outputs(3963) <= a xor b;
    layer4_outputs(3964) <= not b;
    layer4_outputs(3965) <= not b;
    layer4_outputs(3966) <= a and not b;
    layer4_outputs(3967) <= b and not a;
    layer4_outputs(3968) <= a and not b;
    layer4_outputs(3969) <= '0';
    layer4_outputs(3970) <= not (a and b);
    layer4_outputs(3971) <= not a;
    layer4_outputs(3972) <= not b or a;
    layer4_outputs(3973) <= '1';
    layer4_outputs(3974) <= a;
    layer4_outputs(3975) <= b;
    layer4_outputs(3976) <= not (a and b);
    layer4_outputs(3977) <= not a;
    layer4_outputs(3978) <= not (a xor b);
    layer4_outputs(3979) <= not (a and b);
    layer4_outputs(3980) <= not a or b;
    layer4_outputs(3981) <= '1';
    layer4_outputs(3982) <= b;
    layer4_outputs(3983) <= not b;
    layer4_outputs(3984) <= a and b;
    layer4_outputs(3985) <= not (a or b);
    layer4_outputs(3986) <= a or b;
    layer4_outputs(3987) <= a and b;
    layer4_outputs(3988) <= not a or b;
    layer4_outputs(3989) <= not a or b;
    layer4_outputs(3990) <= a;
    layer4_outputs(3991) <= a;
    layer4_outputs(3992) <= '1';
    layer4_outputs(3993) <= not b;
    layer4_outputs(3994) <= not b;
    layer4_outputs(3995) <= not b;
    layer4_outputs(3996) <= not a;
    layer4_outputs(3997) <= not b or a;
    layer4_outputs(3998) <= not (a and b);
    layer4_outputs(3999) <= not (a and b);
    layer4_outputs(4000) <= b;
    layer4_outputs(4001) <= a;
    layer4_outputs(4002) <= not a;
    layer4_outputs(4003) <= not (a or b);
    layer4_outputs(4004) <= a and not b;
    layer4_outputs(4005) <= not (a and b);
    layer4_outputs(4006) <= not a;
    layer4_outputs(4007) <= b;
    layer4_outputs(4008) <= b and not a;
    layer4_outputs(4009) <= not a;
    layer4_outputs(4010) <= not a or b;
    layer4_outputs(4011) <= a and b;
    layer4_outputs(4012) <= a;
    layer4_outputs(4013) <= a and not b;
    layer4_outputs(4014) <= b;
    layer4_outputs(4015) <= b and not a;
    layer4_outputs(4016) <= a or b;
    layer4_outputs(4017) <= not b;
    layer4_outputs(4018) <= '1';
    layer4_outputs(4019) <= not b;
    layer4_outputs(4020) <= b;
    layer4_outputs(4021) <= a;
    layer4_outputs(4022) <= not b;
    layer4_outputs(4023) <= b;
    layer4_outputs(4024) <= a or b;
    layer4_outputs(4025) <= not (a and b);
    layer4_outputs(4026) <= not a;
    layer4_outputs(4027) <= '1';
    layer4_outputs(4028) <= not (a and b);
    layer4_outputs(4029) <= b;
    layer4_outputs(4030) <= not b or a;
    layer4_outputs(4031) <= a;
    layer4_outputs(4032) <= not b or a;
    layer4_outputs(4033) <= not a or b;
    layer4_outputs(4034) <= a or b;
    layer4_outputs(4035) <= not a;
    layer4_outputs(4036) <= not a;
    layer4_outputs(4037) <= not b or a;
    layer4_outputs(4038) <= a and not b;
    layer4_outputs(4039) <= a and b;
    layer4_outputs(4040) <= b;
    layer4_outputs(4041) <= b;
    layer4_outputs(4042) <= b and not a;
    layer4_outputs(4043) <= not a;
    layer4_outputs(4044) <= not b;
    layer4_outputs(4045) <= a and not b;
    layer4_outputs(4046) <= a or b;
    layer4_outputs(4047) <= '0';
    layer4_outputs(4048) <= not (a and b);
    layer4_outputs(4049) <= a or b;
    layer4_outputs(4050) <= not b or a;
    layer4_outputs(4051) <= '1';
    layer4_outputs(4052) <= a and not b;
    layer4_outputs(4053) <= a;
    layer4_outputs(4054) <= not a;
    layer4_outputs(4055) <= a and not b;
    layer4_outputs(4056) <= not a;
    layer4_outputs(4057) <= b and not a;
    layer4_outputs(4058) <= not b or a;
    layer4_outputs(4059) <= a and b;
    layer4_outputs(4060) <= a and b;
    layer4_outputs(4061) <= not b;
    layer4_outputs(4062) <= not a or b;
    layer4_outputs(4063) <= not b or a;
    layer4_outputs(4064) <= b;
    layer4_outputs(4065) <= a and not b;
    layer4_outputs(4066) <= a;
    layer4_outputs(4067) <= a or b;
    layer4_outputs(4068) <= not (a xor b);
    layer4_outputs(4069) <= a or b;
    layer4_outputs(4070) <= not (a or b);
    layer4_outputs(4071) <= b;
    layer4_outputs(4072) <= not b or a;
    layer4_outputs(4073) <= not b;
    layer4_outputs(4074) <= not b;
    layer4_outputs(4075) <= a xor b;
    layer4_outputs(4076) <= b and not a;
    layer4_outputs(4077) <= a or b;
    layer4_outputs(4078) <= not b or a;
    layer4_outputs(4079) <= b;
    layer4_outputs(4080) <= not b;
    layer4_outputs(4081) <= b and not a;
    layer4_outputs(4082) <= a or b;
    layer4_outputs(4083) <= a and not b;
    layer4_outputs(4084) <= b and not a;
    layer4_outputs(4085) <= not (a or b);
    layer4_outputs(4086) <= b;
    layer4_outputs(4087) <= '1';
    layer4_outputs(4088) <= '0';
    layer4_outputs(4089) <= '1';
    layer4_outputs(4090) <= a xor b;
    layer4_outputs(4091) <= not b or a;
    layer4_outputs(4092) <= b and not a;
    layer4_outputs(4093) <= '1';
    layer4_outputs(4094) <= not (a xor b);
    layer4_outputs(4095) <= '1';
    layer4_outputs(4096) <= not a or b;
    layer4_outputs(4097) <= not (a and b);
    layer4_outputs(4098) <= not (a or b);
    layer4_outputs(4099) <= a and b;
    layer4_outputs(4100) <= a;
    layer4_outputs(4101) <= a and b;
    layer4_outputs(4102) <= not (a and b);
    layer4_outputs(4103) <= b;
    layer4_outputs(4104) <= b;
    layer4_outputs(4105) <= not (a or b);
    layer4_outputs(4106) <= a or b;
    layer4_outputs(4107) <= '0';
    layer4_outputs(4108) <= b;
    layer4_outputs(4109) <= not b or a;
    layer4_outputs(4110) <= a;
    layer4_outputs(4111) <= not a;
    layer4_outputs(4112) <= not a;
    layer4_outputs(4113) <= not b;
    layer4_outputs(4114) <= not a or b;
    layer4_outputs(4115) <= a and not b;
    layer4_outputs(4116) <= b;
    layer4_outputs(4117) <= a;
    layer4_outputs(4118) <= not a;
    layer4_outputs(4119) <= not (a and b);
    layer4_outputs(4120) <= not a;
    layer4_outputs(4121) <= not (a and b);
    layer4_outputs(4122) <= a;
    layer4_outputs(4123) <= not a;
    layer4_outputs(4124) <= b and not a;
    layer4_outputs(4125) <= b;
    layer4_outputs(4126) <= not b;
    layer4_outputs(4127) <= a and b;
    layer4_outputs(4128) <= a and not b;
    layer4_outputs(4129) <= '1';
    layer4_outputs(4130) <= not b or a;
    layer4_outputs(4131) <= not (a and b);
    layer4_outputs(4132) <= not (a or b);
    layer4_outputs(4133) <= not (a or b);
    layer4_outputs(4134) <= b;
    layer4_outputs(4135) <= a and not b;
    layer4_outputs(4136) <= b and not a;
    layer4_outputs(4137) <= a or b;
    layer4_outputs(4138) <= not a or b;
    layer4_outputs(4139) <= not (a and b);
    layer4_outputs(4140) <= not b;
    layer4_outputs(4141) <= a or b;
    layer4_outputs(4142) <= not (a or b);
    layer4_outputs(4143) <= not a;
    layer4_outputs(4144) <= '0';
    layer4_outputs(4145) <= a and b;
    layer4_outputs(4146) <= not b;
    layer4_outputs(4147) <= a;
    layer4_outputs(4148) <= a or b;
    layer4_outputs(4149) <= '1';
    layer4_outputs(4150) <= '0';
    layer4_outputs(4151) <= a or b;
    layer4_outputs(4152) <= not (a and b);
    layer4_outputs(4153) <= not b;
    layer4_outputs(4154) <= '0';
    layer4_outputs(4155) <= not a;
    layer4_outputs(4156) <= b;
    layer4_outputs(4157) <= not a;
    layer4_outputs(4158) <= a xor b;
    layer4_outputs(4159) <= not (a and b);
    layer4_outputs(4160) <= b and not a;
    layer4_outputs(4161) <= not b;
    layer4_outputs(4162) <= a or b;
    layer4_outputs(4163) <= not a or b;
    layer4_outputs(4164) <= not b or a;
    layer4_outputs(4165) <= b and not a;
    layer4_outputs(4166) <= a or b;
    layer4_outputs(4167) <= b;
    layer4_outputs(4168) <= a;
    layer4_outputs(4169) <= not a;
    layer4_outputs(4170) <= a and not b;
    layer4_outputs(4171) <= not b or a;
    layer4_outputs(4172) <= a or b;
    layer4_outputs(4173) <= a or b;
    layer4_outputs(4174) <= not a;
    layer4_outputs(4175) <= a and not b;
    layer4_outputs(4176) <= a or b;
    layer4_outputs(4177) <= not (a and b);
    layer4_outputs(4178) <= b and not a;
    layer4_outputs(4179) <= not a or b;
    layer4_outputs(4180) <= not b;
    layer4_outputs(4181) <= a and not b;
    layer4_outputs(4182) <= not b or a;
    layer4_outputs(4183) <= b;
    layer4_outputs(4184) <= a and not b;
    layer4_outputs(4185) <= not a or b;
    layer4_outputs(4186) <= b;
    layer4_outputs(4187) <= b;
    layer4_outputs(4188) <= not b or a;
    layer4_outputs(4189) <= a xor b;
    layer4_outputs(4190) <= '1';
    layer4_outputs(4191) <= b and not a;
    layer4_outputs(4192) <= '0';
    layer4_outputs(4193) <= '0';
    layer4_outputs(4194) <= not a or b;
    layer4_outputs(4195) <= '0';
    layer4_outputs(4196) <= not a;
    layer4_outputs(4197) <= not (a xor b);
    layer4_outputs(4198) <= not a;
    layer4_outputs(4199) <= '0';
    layer4_outputs(4200) <= a and b;
    layer4_outputs(4201) <= a;
    layer4_outputs(4202) <= not b or a;
    layer4_outputs(4203) <= a and not b;
    layer4_outputs(4204) <= not (a or b);
    layer4_outputs(4205) <= a xor b;
    layer4_outputs(4206) <= not a or b;
    layer4_outputs(4207) <= a or b;
    layer4_outputs(4208) <= b and not a;
    layer4_outputs(4209) <= not b or a;
    layer4_outputs(4210) <= '1';
    layer4_outputs(4211) <= not b or a;
    layer4_outputs(4212) <= not b or a;
    layer4_outputs(4213) <= not b or a;
    layer4_outputs(4214) <= not a;
    layer4_outputs(4215) <= '1';
    layer4_outputs(4216) <= a and b;
    layer4_outputs(4217) <= not a or b;
    layer4_outputs(4218) <= b and not a;
    layer4_outputs(4219) <= b;
    layer4_outputs(4220) <= not (a or b);
    layer4_outputs(4221) <= not (a xor b);
    layer4_outputs(4222) <= '1';
    layer4_outputs(4223) <= a or b;
    layer4_outputs(4224) <= not b;
    layer4_outputs(4225) <= a;
    layer4_outputs(4226) <= a and b;
    layer4_outputs(4227) <= not a;
    layer4_outputs(4228) <= b;
    layer4_outputs(4229) <= a and not b;
    layer4_outputs(4230) <= a and b;
    layer4_outputs(4231) <= not (a or b);
    layer4_outputs(4232) <= not b;
    layer4_outputs(4233) <= not b;
    layer4_outputs(4234) <= not a or b;
    layer4_outputs(4235) <= a;
    layer4_outputs(4236) <= not (a or b);
    layer4_outputs(4237) <= b and not a;
    layer4_outputs(4238) <= '0';
    layer4_outputs(4239) <= a and not b;
    layer4_outputs(4240) <= a and not b;
    layer4_outputs(4241) <= a and b;
    layer4_outputs(4242) <= not b or a;
    layer4_outputs(4243) <= b;
    layer4_outputs(4244) <= a or b;
    layer4_outputs(4245) <= not a;
    layer4_outputs(4246) <= a xor b;
    layer4_outputs(4247) <= not a;
    layer4_outputs(4248) <= not a;
    layer4_outputs(4249) <= a xor b;
    layer4_outputs(4250) <= a;
    layer4_outputs(4251) <= a;
    layer4_outputs(4252) <= a;
    layer4_outputs(4253) <= not b;
    layer4_outputs(4254) <= not (a xor b);
    layer4_outputs(4255) <= not a;
    layer4_outputs(4256) <= not (a and b);
    layer4_outputs(4257) <= not a;
    layer4_outputs(4258) <= a and b;
    layer4_outputs(4259) <= not (a or b);
    layer4_outputs(4260) <= '0';
    layer4_outputs(4261) <= b and not a;
    layer4_outputs(4262) <= a or b;
    layer4_outputs(4263) <= not (a xor b);
    layer4_outputs(4264) <= a and b;
    layer4_outputs(4265) <= '1';
    layer4_outputs(4266) <= b;
    layer4_outputs(4267) <= not b or a;
    layer4_outputs(4268) <= not b or a;
    layer4_outputs(4269) <= b;
    layer4_outputs(4270) <= '1';
    layer4_outputs(4271) <= a and b;
    layer4_outputs(4272) <= a;
    layer4_outputs(4273) <= not b or a;
    layer4_outputs(4274) <= b;
    layer4_outputs(4275) <= not b or a;
    layer4_outputs(4276) <= not (a xor b);
    layer4_outputs(4277) <= not a;
    layer4_outputs(4278) <= not b;
    layer4_outputs(4279) <= not (a and b);
    layer4_outputs(4280) <= a;
    layer4_outputs(4281) <= not b;
    layer4_outputs(4282) <= '1';
    layer4_outputs(4283) <= not a or b;
    layer4_outputs(4284) <= not a or b;
    layer4_outputs(4285) <= a and b;
    layer4_outputs(4286) <= '1';
    layer4_outputs(4287) <= b and not a;
    layer4_outputs(4288) <= not a or b;
    layer4_outputs(4289) <= a and b;
    layer4_outputs(4290) <= not (a and b);
    layer4_outputs(4291) <= '0';
    layer4_outputs(4292) <= b and not a;
    layer4_outputs(4293) <= a;
    layer4_outputs(4294) <= '0';
    layer4_outputs(4295) <= not a;
    layer4_outputs(4296) <= '0';
    layer4_outputs(4297) <= a;
    layer4_outputs(4298) <= a and b;
    layer4_outputs(4299) <= not a or b;
    layer4_outputs(4300) <= not (a and b);
    layer4_outputs(4301) <= b and not a;
    layer4_outputs(4302) <= b and not a;
    layer4_outputs(4303) <= not (a and b);
    layer4_outputs(4304) <= not b;
    layer4_outputs(4305) <= a and b;
    layer4_outputs(4306) <= b and not a;
    layer4_outputs(4307) <= not (a or b);
    layer4_outputs(4308) <= not a or b;
    layer4_outputs(4309) <= b and not a;
    layer4_outputs(4310) <= not a;
    layer4_outputs(4311) <= b and not a;
    layer4_outputs(4312) <= b;
    layer4_outputs(4313) <= a;
    layer4_outputs(4314) <= a;
    layer4_outputs(4315) <= b;
    layer4_outputs(4316) <= a and not b;
    layer4_outputs(4317) <= '1';
    layer4_outputs(4318) <= not (a and b);
    layer4_outputs(4319) <= b and not a;
    layer4_outputs(4320) <= not b or a;
    layer4_outputs(4321) <= not b;
    layer4_outputs(4322) <= not (a and b);
    layer4_outputs(4323) <= a;
    layer4_outputs(4324) <= not b;
    layer4_outputs(4325) <= not a;
    layer4_outputs(4326) <= not a;
    layer4_outputs(4327) <= not a;
    layer4_outputs(4328) <= not a or b;
    layer4_outputs(4329) <= not (a xor b);
    layer4_outputs(4330) <= not b or a;
    layer4_outputs(4331) <= a and b;
    layer4_outputs(4332) <= a or b;
    layer4_outputs(4333) <= a;
    layer4_outputs(4334) <= a and not b;
    layer4_outputs(4335) <= not (a or b);
    layer4_outputs(4336) <= not (a and b);
    layer4_outputs(4337) <= b;
    layer4_outputs(4338) <= b and not a;
    layer4_outputs(4339) <= a and not b;
    layer4_outputs(4340) <= not (a and b);
    layer4_outputs(4341) <= b and not a;
    layer4_outputs(4342) <= not (a xor b);
    layer4_outputs(4343) <= not (a and b);
    layer4_outputs(4344) <= b;
    layer4_outputs(4345) <= a and not b;
    layer4_outputs(4346) <= not (a and b);
    layer4_outputs(4347) <= not a;
    layer4_outputs(4348) <= not a or b;
    layer4_outputs(4349) <= a or b;
    layer4_outputs(4350) <= a;
    layer4_outputs(4351) <= a and b;
    layer4_outputs(4352) <= not a or b;
    layer4_outputs(4353) <= not (a and b);
    layer4_outputs(4354) <= '1';
    layer4_outputs(4355) <= not (a xor b);
    layer4_outputs(4356) <= not b or a;
    layer4_outputs(4357) <= a;
    layer4_outputs(4358) <= b;
    layer4_outputs(4359) <= a and b;
    layer4_outputs(4360) <= a;
    layer4_outputs(4361) <= not b or a;
    layer4_outputs(4362) <= a or b;
    layer4_outputs(4363) <= a and not b;
    layer4_outputs(4364) <= a or b;
    layer4_outputs(4365) <= b;
    layer4_outputs(4366) <= '1';
    layer4_outputs(4367) <= b;
    layer4_outputs(4368) <= not b or a;
    layer4_outputs(4369) <= a xor b;
    layer4_outputs(4370) <= not (a xor b);
    layer4_outputs(4371) <= a and b;
    layer4_outputs(4372) <= a;
    layer4_outputs(4373) <= not (a or b);
    layer4_outputs(4374) <= a and b;
    layer4_outputs(4375) <= not (a and b);
    layer4_outputs(4376) <= not (a xor b);
    layer4_outputs(4377) <= a and not b;
    layer4_outputs(4378) <= not a or b;
    layer4_outputs(4379) <= not b;
    layer4_outputs(4380) <= not b or a;
    layer4_outputs(4381) <= not a;
    layer4_outputs(4382) <= a and not b;
    layer4_outputs(4383) <= not (a and b);
    layer4_outputs(4384) <= a and not b;
    layer4_outputs(4385) <= b;
    layer4_outputs(4386) <= a and b;
    layer4_outputs(4387) <= not a or b;
    layer4_outputs(4388) <= not a;
    layer4_outputs(4389) <= a;
    layer4_outputs(4390) <= not b or a;
    layer4_outputs(4391) <= not (a xor b);
    layer4_outputs(4392) <= '0';
    layer4_outputs(4393) <= a or b;
    layer4_outputs(4394) <= a and b;
    layer4_outputs(4395) <= not b or a;
    layer4_outputs(4396) <= a and b;
    layer4_outputs(4397) <= not (a or b);
    layer4_outputs(4398) <= '1';
    layer4_outputs(4399) <= a and b;
    layer4_outputs(4400) <= not b or a;
    layer4_outputs(4401) <= a xor b;
    layer4_outputs(4402) <= not a;
    layer4_outputs(4403) <= b;
    layer4_outputs(4404) <= not (a and b);
    layer4_outputs(4405) <= a and not b;
    layer4_outputs(4406) <= b;
    layer4_outputs(4407) <= not (a or b);
    layer4_outputs(4408) <= '1';
    layer4_outputs(4409) <= a and not b;
    layer4_outputs(4410) <= a;
    layer4_outputs(4411) <= a or b;
    layer4_outputs(4412) <= a;
    layer4_outputs(4413) <= not a;
    layer4_outputs(4414) <= a and b;
    layer4_outputs(4415) <= '1';
    layer4_outputs(4416) <= not b or a;
    layer4_outputs(4417) <= not a or b;
    layer4_outputs(4418) <= b and not a;
    layer4_outputs(4419) <= a and not b;
    layer4_outputs(4420) <= a or b;
    layer4_outputs(4421) <= not a or b;
    layer4_outputs(4422) <= b and not a;
    layer4_outputs(4423) <= not (a and b);
    layer4_outputs(4424) <= b;
    layer4_outputs(4425) <= a xor b;
    layer4_outputs(4426) <= a and not b;
    layer4_outputs(4427) <= b;
    layer4_outputs(4428) <= a and b;
    layer4_outputs(4429) <= a;
    layer4_outputs(4430) <= a or b;
    layer4_outputs(4431) <= a and not b;
    layer4_outputs(4432) <= not a;
    layer4_outputs(4433) <= '0';
    layer4_outputs(4434) <= a or b;
    layer4_outputs(4435) <= b;
    layer4_outputs(4436) <= a and b;
    layer4_outputs(4437) <= b;
    layer4_outputs(4438) <= '1';
    layer4_outputs(4439) <= not a;
    layer4_outputs(4440) <= not b or a;
    layer4_outputs(4441) <= not (a or b);
    layer4_outputs(4442) <= a;
    layer4_outputs(4443) <= a;
    layer4_outputs(4444) <= a;
    layer4_outputs(4445) <= not a;
    layer4_outputs(4446) <= '1';
    layer4_outputs(4447) <= not (a and b);
    layer4_outputs(4448) <= not (a or b);
    layer4_outputs(4449) <= not a;
    layer4_outputs(4450) <= '0';
    layer4_outputs(4451) <= not (a and b);
    layer4_outputs(4452) <= not b;
    layer4_outputs(4453) <= not (a or b);
    layer4_outputs(4454) <= not (a and b);
    layer4_outputs(4455) <= not (a xor b);
    layer4_outputs(4456) <= a and not b;
    layer4_outputs(4457) <= '1';
    layer4_outputs(4458) <= b and not a;
    layer4_outputs(4459) <= a and b;
    layer4_outputs(4460) <= not (a or b);
    layer4_outputs(4461) <= not b or a;
    layer4_outputs(4462) <= not (a xor b);
    layer4_outputs(4463) <= a;
    layer4_outputs(4464) <= '0';
    layer4_outputs(4465) <= a and not b;
    layer4_outputs(4466) <= not b;
    layer4_outputs(4467) <= b;
    layer4_outputs(4468) <= '1';
    layer4_outputs(4469) <= b and not a;
    layer4_outputs(4470) <= a or b;
    layer4_outputs(4471) <= not a;
    layer4_outputs(4472) <= not a or b;
    layer4_outputs(4473) <= b;
    layer4_outputs(4474) <= not b;
    layer4_outputs(4475) <= a;
    layer4_outputs(4476) <= not a;
    layer4_outputs(4477) <= not a;
    layer4_outputs(4478) <= b;
    layer4_outputs(4479) <= a or b;
    layer4_outputs(4480) <= b;
    layer4_outputs(4481) <= a;
    layer4_outputs(4482) <= not b or a;
    layer4_outputs(4483) <= '1';
    layer4_outputs(4484) <= not (a or b);
    layer4_outputs(4485) <= not (a or b);
    layer4_outputs(4486) <= not a;
    layer4_outputs(4487) <= a or b;
    layer4_outputs(4488) <= '0';
    layer4_outputs(4489) <= not a;
    layer4_outputs(4490) <= a;
    layer4_outputs(4491) <= b;
    layer4_outputs(4492) <= b;
    layer4_outputs(4493) <= '0';
    layer4_outputs(4494) <= not b or a;
    layer4_outputs(4495) <= not a or b;
    layer4_outputs(4496) <= a;
    layer4_outputs(4497) <= not b or a;
    layer4_outputs(4498) <= not b or a;
    layer4_outputs(4499) <= a;
    layer4_outputs(4500) <= a;
    layer4_outputs(4501) <= not b or a;
    layer4_outputs(4502) <= a and not b;
    layer4_outputs(4503) <= '0';
    layer4_outputs(4504) <= not a;
    layer4_outputs(4505) <= '0';
    layer4_outputs(4506) <= not (a xor b);
    layer4_outputs(4507) <= not (a or b);
    layer4_outputs(4508) <= not b;
    layer4_outputs(4509) <= b;
    layer4_outputs(4510) <= '1';
    layer4_outputs(4511) <= '0';
    layer4_outputs(4512) <= not (a and b);
    layer4_outputs(4513) <= b;
    layer4_outputs(4514) <= b and not a;
    layer4_outputs(4515) <= a and not b;
    layer4_outputs(4516) <= a and not b;
    layer4_outputs(4517) <= not a;
    layer4_outputs(4518) <= not b;
    layer4_outputs(4519) <= a xor b;
    layer4_outputs(4520) <= not (a and b);
    layer4_outputs(4521) <= a;
    layer4_outputs(4522) <= not a or b;
    layer4_outputs(4523) <= a and b;
    layer4_outputs(4524) <= not (a and b);
    layer4_outputs(4525) <= b and not a;
    layer4_outputs(4526) <= not a or b;
    layer4_outputs(4527) <= a xor b;
    layer4_outputs(4528) <= '0';
    layer4_outputs(4529) <= a and b;
    layer4_outputs(4530) <= a;
    layer4_outputs(4531) <= '0';
    layer4_outputs(4532) <= a and not b;
    layer4_outputs(4533) <= not b;
    layer4_outputs(4534) <= a and b;
    layer4_outputs(4535) <= not b or a;
    layer4_outputs(4536) <= not (a and b);
    layer4_outputs(4537) <= not (a or b);
    layer4_outputs(4538) <= b and not a;
    layer4_outputs(4539) <= a or b;
    layer4_outputs(4540) <= b and not a;
    layer4_outputs(4541) <= a;
    layer4_outputs(4542) <= a;
    layer4_outputs(4543) <= not a or b;
    layer4_outputs(4544) <= not (a xor b);
    layer4_outputs(4545) <= not (a or b);
    layer4_outputs(4546) <= b;
    layer4_outputs(4547) <= b and not a;
    layer4_outputs(4548) <= b and not a;
    layer4_outputs(4549) <= not (a xor b);
    layer4_outputs(4550) <= a or b;
    layer4_outputs(4551) <= '0';
    layer4_outputs(4552) <= '1';
    layer4_outputs(4553) <= b;
    layer4_outputs(4554) <= a;
    layer4_outputs(4555) <= not b or a;
    layer4_outputs(4556) <= not a;
    layer4_outputs(4557) <= a and b;
    layer4_outputs(4558) <= not (a and b);
    layer4_outputs(4559) <= not b or a;
    layer4_outputs(4560) <= not a;
    layer4_outputs(4561) <= not (a and b);
    layer4_outputs(4562) <= a or b;
    layer4_outputs(4563) <= not (a and b);
    layer4_outputs(4564) <= b;
    layer4_outputs(4565) <= not b or a;
    layer4_outputs(4566) <= a;
    layer4_outputs(4567) <= a or b;
    layer4_outputs(4568) <= '0';
    layer4_outputs(4569) <= not (a and b);
    layer4_outputs(4570) <= '1';
    layer4_outputs(4571) <= not b;
    layer4_outputs(4572) <= not (a and b);
    layer4_outputs(4573) <= not (a and b);
    layer4_outputs(4574) <= a or b;
    layer4_outputs(4575) <= not a;
    layer4_outputs(4576) <= '0';
    layer4_outputs(4577) <= a;
    layer4_outputs(4578) <= a or b;
    layer4_outputs(4579) <= not a or b;
    layer4_outputs(4580) <= b and not a;
    layer4_outputs(4581) <= not a;
    layer4_outputs(4582) <= a;
    layer4_outputs(4583) <= not a;
    layer4_outputs(4584) <= not (a or b);
    layer4_outputs(4585) <= b;
    layer4_outputs(4586) <= not (a xor b);
    layer4_outputs(4587) <= '0';
    layer4_outputs(4588) <= a;
    layer4_outputs(4589) <= not b or a;
    layer4_outputs(4590) <= not b or a;
    layer4_outputs(4591) <= a xor b;
    layer4_outputs(4592) <= not b;
    layer4_outputs(4593) <= b and not a;
    layer4_outputs(4594) <= a or b;
    layer4_outputs(4595) <= '0';
    layer4_outputs(4596) <= '1';
    layer4_outputs(4597) <= a or b;
    layer4_outputs(4598) <= not a or b;
    layer4_outputs(4599) <= b;
    layer4_outputs(4600) <= a;
    layer4_outputs(4601) <= '1';
    layer4_outputs(4602) <= a;
    layer4_outputs(4603) <= '1';
    layer4_outputs(4604) <= not (a or b);
    layer4_outputs(4605) <= not b;
    layer4_outputs(4606) <= a;
    layer4_outputs(4607) <= a and b;
    layer4_outputs(4608) <= b and not a;
    layer4_outputs(4609) <= not (a and b);
    layer4_outputs(4610) <= a;
    layer4_outputs(4611) <= not a;
    layer4_outputs(4612) <= not b;
    layer4_outputs(4613) <= not a or b;
    layer4_outputs(4614) <= not (a and b);
    layer4_outputs(4615) <= not (a and b);
    layer4_outputs(4616) <= '1';
    layer4_outputs(4617) <= not b;
    layer4_outputs(4618) <= '0';
    layer4_outputs(4619) <= a xor b;
    layer4_outputs(4620) <= a;
    layer4_outputs(4621) <= a or b;
    layer4_outputs(4622) <= not a or b;
    layer4_outputs(4623) <= a;
    layer4_outputs(4624) <= not (a and b);
    layer4_outputs(4625) <= b;
    layer4_outputs(4626) <= not a;
    layer4_outputs(4627) <= not b;
    layer4_outputs(4628) <= a and not b;
    layer4_outputs(4629) <= a and b;
    layer4_outputs(4630) <= a or b;
    layer4_outputs(4631) <= not (a and b);
    layer4_outputs(4632) <= not (a or b);
    layer4_outputs(4633) <= '1';
    layer4_outputs(4634) <= a and b;
    layer4_outputs(4635) <= '1';
    layer4_outputs(4636) <= '0';
    layer4_outputs(4637) <= '1';
    layer4_outputs(4638) <= not (a or b);
    layer4_outputs(4639) <= not b;
    layer4_outputs(4640) <= not (a or b);
    layer4_outputs(4641) <= a;
    layer4_outputs(4642) <= not a;
    layer4_outputs(4643) <= not b or a;
    layer4_outputs(4644) <= a and not b;
    layer4_outputs(4645) <= a and b;
    layer4_outputs(4646) <= a or b;
    layer4_outputs(4647) <= a and b;
    layer4_outputs(4648) <= not (a or b);
    layer4_outputs(4649) <= b and not a;
    layer4_outputs(4650) <= a or b;
    layer4_outputs(4651) <= b;
    layer4_outputs(4652) <= a and not b;
    layer4_outputs(4653) <= not (a and b);
    layer4_outputs(4654) <= a and not b;
    layer4_outputs(4655) <= not (a and b);
    layer4_outputs(4656) <= b;
    layer4_outputs(4657) <= b and not a;
    layer4_outputs(4658) <= not a or b;
    layer4_outputs(4659) <= not b;
    layer4_outputs(4660) <= b;
    layer4_outputs(4661) <= a and b;
    layer4_outputs(4662) <= '0';
    layer4_outputs(4663) <= not (a or b);
    layer4_outputs(4664) <= '1';
    layer4_outputs(4665) <= not b;
    layer4_outputs(4666) <= b;
    layer4_outputs(4667) <= not (a and b);
    layer4_outputs(4668) <= a;
    layer4_outputs(4669) <= not (a or b);
    layer4_outputs(4670) <= a;
    layer4_outputs(4671) <= a or b;
    layer4_outputs(4672) <= a xor b;
    layer4_outputs(4673) <= a;
    layer4_outputs(4674) <= not b or a;
    layer4_outputs(4675) <= not (a or b);
    layer4_outputs(4676) <= a or b;
    layer4_outputs(4677) <= '0';
    layer4_outputs(4678) <= b;
    layer4_outputs(4679) <= '1';
    layer4_outputs(4680) <= a;
    layer4_outputs(4681) <= b and not a;
    layer4_outputs(4682) <= not a;
    layer4_outputs(4683) <= not a;
    layer4_outputs(4684) <= a and b;
    layer4_outputs(4685) <= a and not b;
    layer4_outputs(4686) <= b;
    layer4_outputs(4687) <= not b;
    layer4_outputs(4688) <= '0';
    layer4_outputs(4689) <= '0';
    layer4_outputs(4690) <= b and not a;
    layer4_outputs(4691) <= not b;
    layer4_outputs(4692) <= a and not b;
    layer4_outputs(4693) <= a;
    layer4_outputs(4694) <= not a or b;
    layer4_outputs(4695) <= not a;
    layer4_outputs(4696) <= a;
    layer4_outputs(4697) <= '0';
    layer4_outputs(4698) <= a;
    layer4_outputs(4699) <= not (a xor b);
    layer4_outputs(4700) <= not b;
    layer4_outputs(4701) <= b and not a;
    layer4_outputs(4702) <= not b or a;
    layer4_outputs(4703) <= not b;
    layer4_outputs(4704) <= not a or b;
    layer4_outputs(4705) <= not a;
    layer4_outputs(4706) <= not a;
    layer4_outputs(4707) <= not (a and b);
    layer4_outputs(4708) <= b and not a;
    layer4_outputs(4709) <= a and b;
    layer4_outputs(4710) <= a and not b;
    layer4_outputs(4711) <= a;
    layer4_outputs(4712) <= not (a or b);
    layer4_outputs(4713) <= not b or a;
    layer4_outputs(4714) <= a or b;
    layer4_outputs(4715) <= '1';
    layer4_outputs(4716) <= not a;
    layer4_outputs(4717) <= not (a or b);
    layer4_outputs(4718) <= b and not a;
    layer4_outputs(4719) <= '1';
    layer4_outputs(4720) <= '1';
    layer4_outputs(4721) <= not (a and b);
    layer4_outputs(4722) <= not (a and b);
    layer4_outputs(4723) <= a or b;
    layer4_outputs(4724) <= '1';
    layer4_outputs(4725) <= not (a and b);
    layer4_outputs(4726) <= not b;
    layer4_outputs(4727) <= not b or a;
    layer4_outputs(4728) <= not (a xor b);
    layer4_outputs(4729) <= not a or b;
    layer4_outputs(4730) <= '1';
    layer4_outputs(4731) <= a;
    layer4_outputs(4732) <= b;
    layer4_outputs(4733) <= not a or b;
    layer4_outputs(4734) <= not a or b;
    layer4_outputs(4735) <= not (a and b);
    layer4_outputs(4736) <= b and not a;
    layer4_outputs(4737) <= '1';
    layer4_outputs(4738) <= not b;
    layer4_outputs(4739) <= a xor b;
    layer4_outputs(4740) <= '1';
    layer4_outputs(4741) <= a;
    layer4_outputs(4742) <= a;
    layer4_outputs(4743) <= a and not b;
    layer4_outputs(4744) <= b;
    layer4_outputs(4745) <= not a;
    layer4_outputs(4746) <= not (a or b);
    layer4_outputs(4747) <= not b;
    layer4_outputs(4748) <= not a or b;
    layer4_outputs(4749) <= b and not a;
    layer4_outputs(4750) <= not b;
    layer4_outputs(4751) <= not b;
    layer4_outputs(4752) <= not b;
    layer4_outputs(4753) <= '0';
    layer4_outputs(4754) <= a and not b;
    layer4_outputs(4755) <= not b;
    layer4_outputs(4756) <= not a;
    layer4_outputs(4757) <= not b;
    layer4_outputs(4758) <= b and not a;
    layer4_outputs(4759) <= b;
    layer4_outputs(4760) <= '0';
    layer4_outputs(4761) <= a xor b;
    layer4_outputs(4762) <= a;
    layer4_outputs(4763) <= not (a or b);
    layer4_outputs(4764) <= b and not a;
    layer4_outputs(4765) <= '0';
    layer4_outputs(4766) <= a xor b;
    layer4_outputs(4767) <= not (a and b);
    layer4_outputs(4768) <= not b or a;
    layer4_outputs(4769) <= a or b;
    layer4_outputs(4770) <= a and not b;
    layer4_outputs(4771) <= not a or b;
    layer4_outputs(4772) <= a and not b;
    layer4_outputs(4773) <= b;
    layer4_outputs(4774) <= '1';
    layer4_outputs(4775) <= b and not a;
    layer4_outputs(4776) <= a or b;
    layer4_outputs(4777) <= not a or b;
    layer4_outputs(4778) <= a or b;
    layer4_outputs(4779) <= a and b;
    layer4_outputs(4780) <= not (a or b);
    layer4_outputs(4781) <= not (a or b);
    layer4_outputs(4782) <= not b or a;
    layer4_outputs(4783) <= b and not a;
    layer4_outputs(4784) <= not a;
    layer4_outputs(4785) <= a or b;
    layer4_outputs(4786) <= b;
    layer4_outputs(4787) <= a;
    layer4_outputs(4788) <= '0';
    layer4_outputs(4789) <= a;
    layer4_outputs(4790) <= b and not a;
    layer4_outputs(4791) <= b;
    layer4_outputs(4792) <= a or b;
    layer4_outputs(4793) <= b and not a;
    layer4_outputs(4794) <= not a;
    layer4_outputs(4795) <= not (a or b);
    layer4_outputs(4796) <= a and b;
    layer4_outputs(4797) <= not a or b;
    layer4_outputs(4798) <= '0';
    layer4_outputs(4799) <= not a;
    layer4_outputs(4800) <= a;
    layer4_outputs(4801) <= a or b;
    layer4_outputs(4802) <= not a;
    layer4_outputs(4803) <= a;
    layer4_outputs(4804) <= not (a or b);
    layer4_outputs(4805) <= a and b;
    layer4_outputs(4806) <= a and not b;
    layer4_outputs(4807) <= not a;
    layer4_outputs(4808) <= '0';
    layer4_outputs(4809) <= not a;
    layer4_outputs(4810) <= b;
    layer4_outputs(4811) <= not a;
    layer4_outputs(4812) <= a and b;
    layer4_outputs(4813) <= b;
    layer4_outputs(4814) <= not a;
    layer4_outputs(4815) <= not (a and b);
    layer4_outputs(4816) <= a;
    layer4_outputs(4817) <= not (a xor b);
    layer4_outputs(4818) <= '0';
    layer4_outputs(4819) <= not a;
    layer4_outputs(4820) <= '1';
    layer4_outputs(4821) <= b;
    layer4_outputs(4822) <= a xor b;
    layer4_outputs(4823) <= a and not b;
    layer4_outputs(4824) <= a and b;
    layer4_outputs(4825) <= not b;
    layer4_outputs(4826) <= not (a and b);
    layer4_outputs(4827) <= not a or b;
    layer4_outputs(4828) <= not b or a;
    layer4_outputs(4829) <= not (a or b);
    layer4_outputs(4830) <= b;
    layer4_outputs(4831) <= '0';
    layer4_outputs(4832) <= not a;
    layer4_outputs(4833) <= a and not b;
    layer4_outputs(4834) <= '0';
    layer4_outputs(4835) <= '0';
    layer4_outputs(4836) <= '1';
    layer4_outputs(4837) <= not b;
    layer4_outputs(4838) <= b and not a;
    layer4_outputs(4839) <= not a or b;
    layer4_outputs(4840) <= '1';
    layer4_outputs(4841) <= a and not b;
    layer4_outputs(4842) <= not (a and b);
    layer4_outputs(4843) <= a and b;
    layer4_outputs(4844) <= not (a xor b);
    layer4_outputs(4845) <= a;
    layer4_outputs(4846) <= not (a and b);
    layer4_outputs(4847) <= b;
    layer4_outputs(4848) <= b and not a;
    layer4_outputs(4849) <= not (a and b);
    layer4_outputs(4850) <= '1';
    layer4_outputs(4851) <= b and not a;
    layer4_outputs(4852) <= not (a xor b);
    layer4_outputs(4853) <= not a or b;
    layer4_outputs(4854) <= not a;
    layer4_outputs(4855) <= b;
    layer4_outputs(4856) <= b;
    layer4_outputs(4857) <= not (a or b);
    layer4_outputs(4858) <= a;
    layer4_outputs(4859) <= b and not a;
    layer4_outputs(4860) <= not (a xor b);
    layer4_outputs(4861) <= a or b;
    layer4_outputs(4862) <= a;
    layer4_outputs(4863) <= a and b;
    layer4_outputs(4864) <= a and not b;
    layer4_outputs(4865) <= '1';
    layer4_outputs(4866) <= a and not b;
    layer4_outputs(4867) <= b and not a;
    layer4_outputs(4868) <= not a;
    layer4_outputs(4869) <= a or b;
    layer4_outputs(4870) <= not (a and b);
    layer4_outputs(4871) <= '0';
    layer4_outputs(4872) <= '0';
    layer4_outputs(4873) <= a xor b;
    layer4_outputs(4874) <= '0';
    layer4_outputs(4875) <= not b;
    layer4_outputs(4876) <= not b or a;
    layer4_outputs(4877) <= not b or a;
    layer4_outputs(4878) <= not (a and b);
    layer4_outputs(4879) <= a and b;
    layer4_outputs(4880) <= not b;
    layer4_outputs(4881) <= a or b;
    layer4_outputs(4882) <= '1';
    layer4_outputs(4883) <= not (a and b);
    layer4_outputs(4884) <= not b;
    layer4_outputs(4885) <= b and not a;
    layer4_outputs(4886) <= not b or a;
    layer4_outputs(4887) <= a or b;
    layer4_outputs(4888) <= '1';
    layer4_outputs(4889) <= '1';
    layer4_outputs(4890) <= not b;
    layer4_outputs(4891) <= not a;
    layer4_outputs(4892) <= a or b;
    layer4_outputs(4893) <= b;
    layer4_outputs(4894) <= '1';
    layer4_outputs(4895) <= not a or b;
    layer4_outputs(4896) <= not b;
    layer4_outputs(4897) <= a and b;
    layer4_outputs(4898) <= not a;
    layer4_outputs(4899) <= a or b;
    layer4_outputs(4900) <= b and not a;
    layer4_outputs(4901) <= not b;
    layer4_outputs(4902) <= b;
    layer4_outputs(4903) <= a and not b;
    layer4_outputs(4904) <= a;
    layer4_outputs(4905) <= a;
    layer4_outputs(4906) <= '0';
    layer4_outputs(4907) <= not (a or b);
    layer4_outputs(4908) <= not a or b;
    layer4_outputs(4909) <= '1';
    layer4_outputs(4910) <= not a;
    layer4_outputs(4911) <= not a or b;
    layer4_outputs(4912) <= '0';
    layer4_outputs(4913) <= not (a and b);
    layer4_outputs(4914) <= '1';
    layer4_outputs(4915) <= '0';
    layer4_outputs(4916) <= a or b;
    layer4_outputs(4917) <= not (a and b);
    layer4_outputs(4918) <= a;
    layer4_outputs(4919) <= not (a and b);
    layer4_outputs(4920) <= '0';
    layer4_outputs(4921) <= not (a or b);
    layer4_outputs(4922) <= b;
    layer4_outputs(4923) <= not b;
    layer4_outputs(4924) <= b and not a;
    layer4_outputs(4925) <= b and not a;
    layer4_outputs(4926) <= a or b;
    layer4_outputs(4927) <= not a or b;
    layer4_outputs(4928) <= a and b;
    layer4_outputs(4929) <= a and not b;
    layer4_outputs(4930) <= not b;
    layer4_outputs(4931) <= a and not b;
    layer4_outputs(4932) <= not b or a;
    layer4_outputs(4933) <= a and not b;
    layer4_outputs(4934) <= a or b;
    layer4_outputs(4935) <= not a;
    layer4_outputs(4936) <= not b;
    layer4_outputs(4937) <= not a;
    layer4_outputs(4938) <= not (a or b);
    layer4_outputs(4939) <= a and b;
    layer4_outputs(4940) <= '0';
    layer4_outputs(4941) <= not a or b;
    layer4_outputs(4942) <= '1';
    layer4_outputs(4943) <= a;
    layer4_outputs(4944) <= b;
    layer4_outputs(4945) <= '0';
    layer4_outputs(4946) <= a and b;
    layer4_outputs(4947) <= not b or a;
    layer4_outputs(4948) <= b;
    layer4_outputs(4949) <= not (a or b);
    layer4_outputs(4950) <= '0';
    layer4_outputs(4951) <= a;
    layer4_outputs(4952) <= a;
    layer4_outputs(4953) <= not (a or b);
    layer4_outputs(4954) <= a;
    layer4_outputs(4955) <= b;
    layer4_outputs(4956) <= '0';
    layer4_outputs(4957) <= not b;
    layer4_outputs(4958) <= b and not a;
    layer4_outputs(4959) <= a;
    layer4_outputs(4960) <= not (a and b);
    layer4_outputs(4961) <= not a or b;
    layer4_outputs(4962) <= a and b;
    layer4_outputs(4963) <= a and not b;
    layer4_outputs(4964) <= not (a and b);
    layer4_outputs(4965) <= '0';
    layer4_outputs(4966) <= '0';
    layer4_outputs(4967) <= not b or a;
    layer4_outputs(4968) <= a or b;
    layer4_outputs(4969) <= a or b;
    layer4_outputs(4970) <= '0';
    layer4_outputs(4971) <= not (a or b);
    layer4_outputs(4972) <= not a or b;
    layer4_outputs(4973) <= not b;
    layer4_outputs(4974) <= not a;
    layer4_outputs(4975) <= b and not a;
    layer4_outputs(4976) <= b;
    layer4_outputs(4977) <= a and not b;
    layer4_outputs(4978) <= a and not b;
    layer4_outputs(4979) <= b;
    layer4_outputs(4980) <= not (a or b);
    layer4_outputs(4981) <= not a or b;
    layer4_outputs(4982) <= a xor b;
    layer4_outputs(4983) <= not a or b;
    layer4_outputs(4984) <= not a;
    layer4_outputs(4985) <= not (a xor b);
    layer4_outputs(4986) <= a and b;
    layer4_outputs(4987) <= a and not b;
    layer4_outputs(4988) <= not (a and b);
    layer4_outputs(4989) <= not b or a;
    layer4_outputs(4990) <= a or b;
    layer4_outputs(4991) <= b;
    layer4_outputs(4992) <= not a;
    layer4_outputs(4993) <= not a or b;
    layer4_outputs(4994) <= '0';
    layer4_outputs(4995) <= not a or b;
    layer4_outputs(4996) <= '1';
    layer4_outputs(4997) <= not (a or b);
    layer4_outputs(4998) <= b;
    layer4_outputs(4999) <= a or b;
    layer4_outputs(5000) <= '0';
    layer4_outputs(5001) <= a and not b;
    layer4_outputs(5002) <= a and not b;
    layer4_outputs(5003) <= not b or a;
    layer4_outputs(5004) <= not a;
    layer4_outputs(5005) <= not (a or b);
    layer4_outputs(5006) <= b;
    layer4_outputs(5007) <= a;
    layer4_outputs(5008) <= not a or b;
    layer4_outputs(5009) <= not a or b;
    layer4_outputs(5010) <= b and not a;
    layer4_outputs(5011) <= not (a xor b);
    layer4_outputs(5012) <= a;
    layer4_outputs(5013) <= b and not a;
    layer4_outputs(5014) <= not (a and b);
    layer4_outputs(5015) <= b;
    layer4_outputs(5016) <= a and not b;
    layer4_outputs(5017) <= b;
    layer4_outputs(5018) <= not b;
    layer4_outputs(5019) <= a and b;
    layer4_outputs(5020) <= '0';
    layer4_outputs(5021) <= a and not b;
    layer4_outputs(5022) <= b;
    layer4_outputs(5023) <= b and not a;
    layer4_outputs(5024) <= not (a or b);
    layer4_outputs(5025) <= b;
    layer4_outputs(5026) <= b;
    layer4_outputs(5027) <= not a;
    layer4_outputs(5028) <= b and not a;
    layer4_outputs(5029) <= a;
    layer4_outputs(5030) <= a and b;
    layer4_outputs(5031) <= b;
    layer4_outputs(5032) <= '1';
    layer4_outputs(5033) <= not b;
    layer4_outputs(5034) <= not b;
    layer4_outputs(5035) <= not b;
    layer4_outputs(5036) <= '0';
    layer4_outputs(5037) <= not b or a;
    layer4_outputs(5038) <= a;
    layer4_outputs(5039) <= '1';
    layer4_outputs(5040) <= not (a xor b);
    layer4_outputs(5041) <= not (a or b);
    layer4_outputs(5042) <= a and not b;
    layer4_outputs(5043) <= not b;
    layer4_outputs(5044) <= b;
    layer4_outputs(5045) <= not (a or b);
    layer4_outputs(5046) <= not b or a;
    layer4_outputs(5047) <= a;
    layer4_outputs(5048) <= not b;
    layer4_outputs(5049) <= a or b;
    layer4_outputs(5050) <= a and not b;
    layer4_outputs(5051) <= a and not b;
    layer4_outputs(5052) <= b;
    layer4_outputs(5053) <= '1';
    layer4_outputs(5054) <= '1';
    layer4_outputs(5055) <= '0';
    layer4_outputs(5056) <= b and not a;
    layer4_outputs(5057) <= a and b;
    layer4_outputs(5058) <= not a;
    layer4_outputs(5059) <= not a or b;
    layer4_outputs(5060) <= a;
    layer4_outputs(5061) <= a and not b;
    layer4_outputs(5062) <= not a;
    layer4_outputs(5063) <= b;
    layer4_outputs(5064) <= not a;
    layer4_outputs(5065) <= b and not a;
    layer4_outputs(5066) <= not (a and b);
    layer4_outputs(5067) <= b and not a;
    layer4_outputs(5068) <= not b or a;
    layer4_outputs(5069) <= a or b;
    layer4_outputs(5070) <= a or b;
    layer4_outputs(5071) <= '0';
    layer4_outputs(5072) <= b;
    layer4_outputs(5073) <= a and b;
    layer4_outputs(5074) <= a and not b;
    layer4_outputs(5075) <= not a;
    layer4_outputs(5076) <= not b or a;
    layer4_outputs(5077) <= a and b;
    layer4_outputs(5078) <= '0';
    layer4_outputs(5079) <= a;
    layer4_outputs(5080) <= not (a or b);
    layer4_outputs(5081) <= a and b;
    layer4_outputs(5082) <= not (a and b);
    layer4_outputs(5083) <= a and not b;
    layer4_outputs(5084) <= not b or a;
    layer4_outputs(5085) <= not b or a;
    layer4_outputs(5086) <= not b or a;
    layer4_outputs(5087) <= '1';
    layer4_outputs(5088) <= not b;
    layer4_outputs(5089) <= a and b;
    layer4_outputs(5090) <= a or b;
    layer4_outputs(5091) <= '0';
    layer4_outputs(5092) <= a and not b;
    layer4_outputs(5093) <= b;
    layer4_outputs(5094) <= b and not a;
    layer4_outputs(5095) <= '0';
    layer4_outputs(5096) <= a and not b;
    layer4_outputs(5097) <= not (a and b);
    layer4_outputs(5098) <= not a;
    layer4_outputs(5099) <= not (a and b);
    layer4_outputs(5100) <= a or b;
    layer4_outputs(5101) <= b and not a;
    layer4_outputs(5102) <= a and b;
    layer4_outputs(5103) <= not (a xor b);
    layer4_outputs(5104) <= b;
    layer4_outputs(5105) <= a and b;
    layer4_outputs(5106) <= not (a or b);
    layer4_outputs(5107) <= b and not a;
    layer4_outputs(5108) <= not a or b;
    layer4_outputs(5109) <= a and not b;
    layer4_outputs(5110) <= not (a and b);
    layer4_outputs(5111) <= a and not b;
    layer4_outputs(5112) <= not b;
    layer4_outputs(5113) <= a or b;
    layer4_outputs(5114) <= '1';
    layer4_outputs(5115) <= not (a and b);
    layer4_outputs(5116) <= a and b;
    layer4_outputs(5117) <= b;
    layer4_outputs(5118) <= a and not b;
    layer4_outputs(5119) <= not a or b;
    layer4_outputs(5120) <= a;
    layer4_outputs(5121) <= not a;
    layer4_outputs(5122) <= not (a or b);
    layer4_outputs(5123) <= not b or a;
    layer4_outputs(5124) <= b and not a;
    layer4_outputs(5125) <= '1';
    layer4_outputs(5126) <= '1';
    layer4_outputs(5127) <= a or b;
    layer4_outputs(5128) <= a and not b;
    layer4_outputs(5129) <= b and not a;
    layer4_outputs(5130) <= not a or b;
    layer4_outputs(5131) <= a and b;
    layer4_outputs(5132) <= a and b;
    layer4_outputs(5133) <= not a;
    layer4_outputs(5134) <= not b or a;
    layer4_outputs(5135) <= a;
    layer4_outputs(5136) <= not b;
    layer4_outputs(5137) <= not (a and b);
    layer4_outputs(5138) <= not b;
    layer4_outputs(5139) <= a and b;
    layer4_outputs(5140) <= '1';
    layer4_outputs(5141) <= a xor b;
    layer4_outputs(5142) <= a and not b;
    layer4_outputs(5143) <= not b or a;
    layer4_outputs(5144) <= not b;
    layer4_outputs(5145) <= a;
    layer4_outputs(5146) <= a and not b;
    layer4_outputs(5147) <= not (a and b);
    layer4_outputs(5148) <= a and not b;
    layer4_outputs(5149) <= a;
    layer4_outputs(5150) <= not (a and b);
    layer4_outputs(5151) <= a and b;
    layer4_outputs(5152) <= a xor b;
    layer4_outputs(5153) <= not b;
    layer4_outputs(5154) <= not b or a;
    layer4_outputs(5155) <= not (a or b);
    layer4_outputs(5156) <= not b;
    layer4_outputs(5157) <= not a;
    layer4_outputs(5158) <= not b;
    layer4_outputs(5159) <= a;
    layer4_outputs(5160) <= a or b;
    layer4_outputs(5161) <= a or b;
    layer4_outputs(5162) <= not (a and b);
    layer4_outputs(5163) <= a;
    layer4_outputs(5164) <= a and b;
    layer4_outputs(5165) <= b and not a;
    layer4_outputs(5166) <= not b;
    layer4_outputs(5167) <= a;
    layer4_outputs(5168) <= a and b;
    layer4_outputs(5169) <= a;
    layer4_outputs(5170) <= not (a and b);
    layer4_outputs(5171) <= a and b;
    layer4_outputs(5172) <= not (a or b);
    layer4_outputs(5173) <= a or b;
    layer4_outputs(5174) <= '0';
    layer4_outputs(5175) <= a;
    layer4_outputs(5176) <= a and not b;
    layer4_outputs(5177) <= '1';
    layer4_outputs(5178) <= not b or a;
    layer4_outputs(5179) <= not b;
    layer4_outputs(5180) <= not (a xor b);
    layer4_outputs(5181) <= not (a xor b);
    layer4_outputs(5182) <= b and not a;
    layer4_outputs(5183) <= not a;
    layer4_outputs(5184) <= not (a and b);
    layer4_outputs(5185) <= not (a and b);
    layer4_outputs(5186) <= b;
    layer4_outputs(5187) <= not a or b;
    layer4_outputs(5188) <= not (a and b);
    layer4_outputs(5189) <= not a or b;
    layer4_outputs(5190) <= b and not a;
    layer4_outputs(5191) <= not (a and b);
    layer4_outputs(5192) <= not (a or b);
    layer4_outputs(5193) <= a;
    layer4_outputs(5194) <= a and not b;
    layer4_outputs(5195) <= '0';
    layer4_outputs(5196) <= b;
    layer4_outputs(5197) <= b and not a;
    layer4_outputs(5198) <= a;
    layer4_outputs(5199) <= not (a or b);
    layer4_outputs(5200) <= not (a or b);
    layer4_outputs(5201) <= not b or a;
    layer4_outputs(5202) <= not (a and b);
    layer4_outputs(5203) <= b;
    layer4_outputs(5204) <= b;
    layer4_outputs(5205) <= not (a or b);
    layer4_outputs(5206) <= not b or a;
    layer4_outputs(5207) <= not b or a;
    layer4_outputs(5208) <= a and b;
    layer4_outputs(5209) <= a or b;
    layer4_outputs(5210) <= not (a and b);
    layer4_outputs(5211) <= a and not b;
    layer4_outputs(5212) <= not (a and b);
    layer4_outputs(5213) <= not (a and b);
    layer4_outputs(5214) <= not b or a;
    layer4_outputs(5215) <= a or b;
    layer4_outputs(5216) <= not (a and b);
    layer4_outputs(5217) <= not b;
    layer4_outputs(5218) <= a;
    layer4_outputs(5219) <= not a or b;
    layer4_outputs(5220) <= not b;
    layer4_outputs(5221) <= '0';
    layer4_outputs(5222) <= '1';
    layer4_outputs(5223) <= a xor b;
    layer4_outputs(5224) <= b;
    layer4_outputs(5225) <= not a or b;
    layer4_outputs(5226) <= a and not b;
    layer4_outputs(5227) <= not (a or b);
    layer4_outputs(5228) <= not b;
    layer4_outputs(5229) <= '1';
    layer4_outputs(5230) <= a and not b;
    layer4_outputs(5231) <= a;
    layer4_outputs(5232) <= a;
    layer4_outputs(5233) <= not a;
    layer4_outputs(5234) <= '1';
    layer4_outputs(5235) <= a xor b;
    layer4_outputs(5236) <= a and b;
    layer4_outputs(5237) <= not a;
    layer4_outputs(5238) <= a xor b;
    layer4_outputs(5239) <= a and b;
    layer4_outputs(5240) <= a;
    layer4_outputs(5241) <= b;
    layer4_outputs(5242) <= a xor b;
    layer4_outputs(5243) <= a or b;
    layer4_outputs(5244) <= not a or b;
    layer4_outputs(5245) <= a and not b;
    layer4_outputs(5246) <= not (a or b);
    layer4_outputs(5247) <= not a or b;
    layer4_outputs(5248) <= not b;
    layer4_outputs(5249) <= b;
    layer4_outputs(5250) <= a;
    layer4_outputs(5251) <= not a;
    layer4_outputs(5252) <= a and b;
    layer4_outputs(5253) <= not (a and b);
    layer4_outputs(5254) <= not b;
    layer4_outputs(5255) <= b and not a;
    layer4_outputs(5256) <= b;
    layer4_outputs(5257) <= not b;
    layer4_outputs(5258) <= not b or a;
    layer4_outputs(5259) <= b;
    layer4_outputs(5260) <= a and b;
    layer4_outputs(5261) <= not b;
    layer4_outputs(5262) <= not a or b;
    layer4_outputs(5263) <= not a or b;
    layer4_outputs(5264) <= b;
    layer4_outputs(5265) <= not b or a;
    layer4_outputs(5266) <= not (a and b);
    layer4_outputs(5267) <= not b;
    layer4_outputs(5268) <= not b;
    layer4_outputs(5269) <= not a;
    layer4_outputs(5270) <= a and not b;
    layer4_outputs(5271) <= not (a or b);
    layer4_outputs(5272) <= not b or a;
    layer4_outputs(5273) <= not a;
    layer4_outputs(5274) <= '1';
    layer4_outputs(5275) <= not (a or b);
    layer4_outputs(5276) <= b and not a;
    layer4_outputs(5277) <= a and not b;
    layer4_outputs(5278) <= b;
    layer4_outputs(5279) <= not a;
    layer4_outputs(5280) <= b and not a;
    layer4_outputs(5281) <= a and b;
    layer4_outputs(5282) <= a xor b;
    layer4_outputs(5283) <= '1';
    layer4_outputs(5284) <= a;
    layer4_outputs(5285) <= not b;
    layer4_outputs(5286) <= a or b;
    layer4_outputs(5287) <= not (a or b);
    layer4_outputs(5288) <= not b;
    layer4_outputs(5289) <= not (a and b);
    layer4_outputs(5290) <= not b or a;
    layer4_outputs(5291) <= a or b;
    layer4_outputs(5292) <= not a or b;
    layer4_outputs(5293) <= '1';
    layer4_outputs(5294) <= a and b;
    layer4_outputs(5295) <= b;
    layer4_outputs(5296) <= not b or a;
    layer4_outputs(5297) <= not a;
    layer4_outputs(5298) <= b;
    layer4_outputs(5299) <= b;
    layer4_outputs(5300) <= a and b;
    layer4_outputs(5301) <= a and not b;
    layer4_outputs(5302) <= not a or b;
    layer4_outputs(5303) <= a and not b;
    layer4_outputs(5304) <= a;
    layer4_outputs(5305) <= '1';
    layer4_outputs(5306) <= not b;
    layer4_outputs(5307) <= not a;
    layer4_outputs(5308) <= not (a and b);
    layer4_outputs(5309) <= not a;
    layer4_outputs(5310) <= a and not b;
    layer4_outputs(5311) <= not b or a;
    layer4_outputs(5312) <= not (a or b);
    layer4_outputs(5313) <= b;
    layer4_outputs(5314) <= a and b;
    layer4_outputs(5315) <= a or b;
    layer4_outputs(5316) <= '1';
    layer4_outputs(5317) <= b;
    layer4_outputs(5318) <= '1';
    layer4_outputs(5319) <= a;
    layer4_outputs(5320) <= a and not b;
    layer4_outputs(5321) <= '0';
    layer4_outputs(5322) <= a;
    layer4_outputs(5323) <= b;
    layer4_outputs(5324) <= '1';
    layer4_outputs(5325) <= b and not a;
    layer4_outputs(5326) <= not b or a;
    layer4_outputs(5327) <= a xor b;
    layer4_outputs(5328) <= not a or b;
    layer4_outputs(5329) <= not (a and b);
    layer4_outputs(5330) <= a and not b;
    layer4_outputs(5331) <= '1';
    layer4_outputs(5332) <= not b;
    layer4_outputs(5333) <= b;
    layer4_outputs(5334) <= b and not a;
    layer4_outputs(5335) <= '0';
    layer4_outputs(5336) <= not b;
    layer4_outputs(5337) <= not a or b;
    layer4_outputs(5338) <= b and not a;
    layer4_outputs(5339) <= not (a xor b);
    layer4_outputs(5340) <= a and b;
    layer4_outputs(5341) <= not b or a;
    layer4_outputs(5342) <= '0';
    layer4_outputs(5343) <= a and b;
    layer4_outputs(5344) <= '1';
    layer4_outputs(5345) <= not (a or b);
    layer4_outputs(5346) <= a;
    layer4_outputs(5347) <= not b;
    layer4_outputs(5348) <= a;
    layer4_outputs(5349) <= a or b;
    layer4_outputs(5350) <= not b or a;
    layer4_outputs(5351) <= a xor b;
    layer4_outputs(5352) <= not b;
    layer4_outputs(5353) <= not (a or b);
    layer4_outputs(5354) <= not b;
    layer4_outputs(5355) <= not (a or b);
    layer4_outputs(5356) <= a or b;
    layer4_outputs(5357) <= not (a xor b);
    layer4_outputs(5358) <= '1';
    layer4_outputs(5359) <= not a or b;
    layer4_outputs(5360) <= a xor b;
    layer4_outputs(5361) <= not b or a;
    layer4_outputs(5362) <= a and b;
    layer4_outputs(5363) <= '1';
    layer4_outputs(5364) <= a or b;
    layer4_outputs(5365) <= a and b;
    layer4_outputs(5366) <= a;
    layer4_outputs(5367) <= not (a and b);
    layer4_outputs(5368) <= not a;
    layer4_outputs(5369) <= not a or b;
    layer4_outputs(5370) <= not a or b;
    layer4_outputs(5371) <= b and not a;
    layer4_outputs(5372) <= '1';
    layer4_outputs(5373) <= not b;
    layer4_outputs(5374) <= not (a or b);
    layer4_outputs(5375) <= a;
    layer4_outputs(5376) <= not (a and b);
    layer4_outputs(5377) <= not a;
    layer4_outputs(5378) <= b;
    layer4_outputs(5379) <= '0';
    layer4_outputs(5380) <= a;
    layer4_outputs(5381) <= not a;
    layer4_outputs(5382) <= not b;
    layer4_outputs(5383) <= a and b;
    layer4_outputs(5384) <= '0';
    layer4_outputs(5385) <= not (a or b);
    layer4_outputs(5386) <= not a or b;
    layer4_outputs(5387) <= not a or b;
    layer4_outputs(5388) <= b;
    layer4_outputs(5389) <= not b or a;
    layer4_outputs(5390) <= a or b;
    layer4_outputs(5391) <= not (a xor b);
    layer4_outputs(5392) <= b;
    layer4_outputs(5393) <= not b or a;
    layer4_outputs(5394) <= '0';
    layer4_outputs(5395) <= not b;
    layer4_outputs(5396) <= a and not b;
    layer4_outputs(5397) <= b and not a;
    layer4_outputs(5398) <= not (a and b);
    layer4_outputs(5399) <= a;
    layer4_outputs(5400) <= b;
    layer4_outputs(5401) <= '0';
    layer4_outputs(5402) <= not (a and b);
    layer4_outputs(5403) <= not (a and b);
    layer4_outputs(5404) <= a;
    layer4_outputs(5405) <= not b or a;
    layer4_outputs(5406) <= a;
    layer4_outputs(5407) <= not a or b;
    layer4_outputs(5408) <= not (a and b);
    layer4_outputs(5409) <= '1';
    layer4_outputs(5410) <= not a;
    layer4_outputs(5411) <= not (a and b);
    layer4_outputs(5412) <= a and b;
    layer4_outputs(5413) <= '1';
    layer4_outputs(5414) <= b;
    layer4_outputs(5415) <= '0';
    layer4_outputs(5416) <= a;
    layer4_outputs(5417) <= not a;
    layer4_outputs(5418) <= a or b;
    layer4_outputs(5419) <= not b;
    layer4_outputs(5420) <= '0';
    layer4_outputs(5421) <= a and not b;
    layer4_outputs(5422) <= not (a and b);
    layer4_outputs(5423) <= not b;
    layer4_outputs(5424) <= not a;
    layer4_outputs(5425) <= not a or b;
    layer4_outputs(5426) <= not a;
    layer4_outputs(5427) <= b;
    layer4_outputs(5428) <= '0';
    layer4_outputs(5429) <= b and not a;
    layer4_outputs(5430) <= not a;
    layer4_outputs(5431) <= a or b;
    layer4_outputs(5432) <= b;
    layer4_outputs(5433) <= b and not a;
    layer4_outputs(5434) <= '1';
    layer4_outputs(5435) <= '1';
    layer4_outputs(5436) <= not (a xor b);
    layer4_outputs(5437) <= '1';
    layer4_outputs(5438) <= a;
    layer4_outputs(5439) <= not b;
    layer4_outputs(5440) <= not a;
    layer4_outputs(5441) <= b;
    layer4_outputs(5442) <= b;
    layer4_outputs(5443) <= a and not b;
    layer4_outputs(5444) <= not a or b;
    layer4_outputs(5445) <= b;
    layer4_outputs(5446) <= a or b;
    layer4_outputs(5447) <= b;
    layer4_outputs(5448) <= not a;
    layer4_outputs(5449) <= a and b;
    layer4_outputs(5450) <= '1';
    layer4_outputs(5451) <= not a;
    layer4_outputs(5452) <= not (a and b);
    layer4_outputs(5453) <= not a;
    layer4_outputs(5454) <= a or b;
    layer4_outputs(5455) <= not b;
    layer4_outputs(5456) <= a or b;
    layer4_outputs(5457) <= not a or b;
    layer4_outputs(5458) <= b and not a;
    layer4_outputs(5459) <= not (a or b);
    layer4_outputs(5460) <= '1';
    layer4_outputs(5461) <= not (a or b);
    layer4_outputs(5462) <= not b or a;
    layer4_outputs(5463) <= not b;
    layer4_outputs(5464) <= a and b;
    layer4_outputs(5465) <= not a or b;
    layer4_outputs(5466) <= a and b;
    layer4_outputs(5467) <= not b or a;
    layer4_outputs(5468) <= a;
    layer4_outputs(5469) <= b;
    layer4_outputs(5470) <= not a or b;
    layer4_outputs(5471) <= not a;
    layer4_outputs(5472) <= not (a and b);
    layer4_outputs(5473) <= a and b;
    layer4_outputs(5474) <= b;
    layer4_outputs(5475) <= a or b;
    layer4_outputs(5476) <= not b or a;
    layer4_outputs(5477) <= a and b;
    layer4_outputs(5478) <= a and b;
    layer4_outputs(5479) <= b and not a;
    layer4_outputs(5480) <= '1';
    layer4_outputs(5481) <= '1';
    layer4_outputs(5482) <= b and not a;
    layer4_outputs(5483) <= not b or a;
    layer4_outputs(5484) <= not (a and b);
    layer4_outputs(5485) <= a xor b;
    layer4_outputs(5486) <= a and not b;
    layer4_outputs(5487) <= not (a and b);
    layer4_outputs(5488) <= a and b;
    layer4_outputs(5489) <= a xor b;
    layer4_outputs(5490) <= not (a xor b);
    layer4_outputs(5491) <= a and not b;
    layer4_outputs(5492) <= not a;
    layer4_outputs(5493) <= a or b;
    layer4_outputs(5494) <= '1';
    layer4_outputs(5495) <= not (a and b);
    layer4_outputs(5496) <= not a;
    layer4_outputs(5497) <= a;
    layer4_outputs(5498) <= '1';
    layer4_outputs(5499) <= b;
    layer4_outputs(5500) <= not b or a;
    layer4_outputs(5501) <= not a or b;
    layer4_outputs(5502) <= not b;
    layer4_outputs(5503) <= not a;
    layer4_outputs(5504) <= a or b;
    layer4_outputs(5505) <= b and not a;
    layer4_outputs(5506) <= not (a or b);
    layer4_outputs(5507) <= a and not b;
    layer4_outputs(5508) <= a;
    layer4_outputs(5509) <= not a;
    layer4_outputs(5510) <= not (a and b);
    layer4_outputs(5511) <= not b;
    layer4_outputs(5512) <= a;
    layer4_outputs(5513) <= not (a and b);
    layer4_outputs(5514) <= not b or a;
    layer4_outputs(5515) <= a xor b;
    layer4_outputs(5516) <= a and b;
    layer4_outputs(5517) <= not a or b;
    layer4_outputs(5518) <= not b;
    layer4_outputs(5519) <= b and not a;
    layer4_outputs(5520) <= a and b;
    layer4_outputs(5521) <= b;
    layer4_outputs(5522) <= a;
    layer4_outputs(5523) <= not (a xor b);
    layer4_outputs(5524) <= not a;
    layer4_outputs(5525) <= not (a or b);
    layer4_outputs(5526) <= a and not b;
    layer4_outputs(5527) <= a and b;
    layer4_outputs(5528) <= not (a and b);
    layer4_outputs(5529) <= b;
    layer4_outputs(5530) <= not a;
    layer4_outputs(5531) <= not a or b;
    layer4_outputs(5532) <= not b or a;
    layer4_outputs(5533) <= not b;
    layer4_outputs(5534) <= not a;
    layer4_outputs(5535) <= a and b;
    layer4_outputs(5536) <= not b;
    layer4_outputs(5537) <= b;
    layer4_outputs(5538) <= not b or a;
    layer4_outputs(5539) <= not b or a;
    layer4_outputs(5540) <= '1';
    layer4_outputs(5541) <= not (a or b);
    layer4_outputs(5542) <= a and not b;
    layer4_outputs(5543) <= not b;
    layer4_outputs(5544) <= a and b;
    layer4_outputs(5545) <= '0';
    layer4_outputs(5546) <= b and not a;
    layer4_outputs(5547) <= not (a and b);
    layer4_outputs(5548) <= not (a or b);
    layer4_outputs(5549) <= '1';
    layer4_outputs(5550) <= not (a xor b);
    layer4_outputs(5551) <= not b or a;
    layer4_outputs(5552) <= a and not b;
    layer4_outputs(5553) <= not a;
    layer4_outputs(5554) <= not b;
    layer4_outputs(5555) <= a xor b;
    layer4_outputs(5556) <= '0';
    layer4_outputs(5557) <= not a or b;
    layer4_outputs(5558) <= a and not b;
    layer4_outputs(5559) <= not (a and b);
    layer4_outputs(5560) <= not a;
    layer4_outputs(5561) <= not a;
    layer4_outputs(5562) <= a and not b;
    layer4_outputs(5563) <= a or b;
    layer4_outputs(5564) <= a and b;
    layer4_outputs(5565) <= b and not a;
    layer4_outputs(5566) <= not (a or b);
    layer4_outputs(5567) <= a and not b;
    layer4_outputs(5568) <= not a;
    layer4_outputs(5569) <= not a or b;
    layer4_outputs(5570) <= a;
    layer4_outputs(5571) <= not a;
    layer4_outputs(5572) <= not a or b;
    layer4_outputs(5573) <= not (a and b);
    layer4_outputs(5574) <= a and b;
    layer4_outputs(5575) <= a;
    layer4_outputs(5576) <= '1';
    layer4_outputs(5577) <= a xor b;
    layer4_outputs(5578) <= a;
    layer4_outputs(5579) <= not (a or b);
    layer4_outputs(5580) <= a or b;
    layer4_outputs(5581) <= '0';
    layer4_outputs(5582) <= not (a xor b);
    layer4_outputs(5583) <= a and not b;
    layer4_outputs(5584) <= not (a xor b);
    layer4_outputs(5585) <= '0';
    layer4_outputs(5586) <= a and b;
    layer4_outputs(5587) <= not b;
    layer4_outputs(5588) <= b and not a;
    layer4_outputs(5589) <= a;
    layer4_outputs(5590) <= b;
    layer4_outputs(5591) <= a and not b;
    layer4_outputs(5592) <= not a or b;
    layer4_outputs(5593) <= b and not a;
    layer4_outputs(5594) <= b;
    layer4_outputs(5595) <= a and not b;
    layer4_outputs(5596) <= b;
    layer4_outputs(5597) <= b and not a;
    layer4_outputs(5598) <= b and not a;
    layer4_outputs(5599) <= not a or b;
    layer4_outputs(5600) <= b and not a;
    layer4_outputs(5601) <= b and not a;
    layer4_outputs(5602) <= '1';
    layer4_outputs(5603) <= not a;
    layer4_outputs(5604) <= not b;
    layer4_outputs(5605) <= not b;
    layer4_outputs(5606) <= not a or b;
    layer4_outputs(5607) <= not b;
    layer4_outputs(5608) <= a and b;
    layer4_outputs(5609) <= not a or b;
    layer4_outputs(5610) <= a and b;
    layer4_outputs(5611) <= a or b;
    layer4_outputs(5612) <= a and not b;
    layer4_outputs(5613) <= a and not b;
    layer4_outputs(5614) <= b;
    layer4_outputs(5615) <= b and not a;
    layer4_outputs(5616) <= a or b;
    layer4_outputs(5617) <= a and b;
    layer4_outputs(5618) <= not a;
    layer4_outputs(5619) <= not a;
    layer4_outputs(5620) <= b and not a;
    layer4_outputs(5621) <= '1';
    layer4_outputs(5622) <= a and not b;
    layer4_outputs(5623) <= b and not a;
    layer4_outputs(5624) <= a;
    layer4_outputs(5625) <= not a;
    layer4_outputs(5626) <= not a;
    layer4_outputs(5627) <= a and b;
    layer4_outputs(5628) <= not b;
    layer4_outputs(5629) <= b and not a;
    layer4_outputs(5630) <= not b or a;
    layer4_outputs(5631) <= a or b;
    layer4_outputs(5632) <= a and not b;
    layer4_outputs(5633) <= a xor b;
    layer4_outputs(5634) <= not a;
    layer4_outputs(5635) <= b and not a;
    layer4_outputs(5636) <= a or b;
    layer4_outputs(5637) <= '1';
    layer4_outputs(5638) <= not a;
    layer4_outputs(5639) <= not a;
    layer4_outputs(5640) <= a or b;
    layer4_outputs(5641) <= not a or b;
    layer4_outputs(5642) <= a and b;
    layer4_outputs(5643) <= a and b;
    layer4_outputs(5644) <= not (a and b);
    layer4_outputs(5645) <= not a;
    layer4_outputs(5646) <= not a or b;
    layer4_outputs(5647) <= a or b;
    layer4_outputs(5648) <= not (a xor b);
    layer4_outputs(5649) <= a and not b;
    layer4_outputs(5650) <= not a or b;
    layer4_outputs(5651) <= not (a or b);
    layer4_outputs(5652) <= a or b;
    layer4_outputs(5653) <= not (a xor b);
    layer4_outputs(5654) <= '1';
    layer4_outputs(5655) <= not b;
    layer4_outputs(5656) <= a or b;
    layer4_outputs(5657) <= b;
    layer4_outputs(5658) <= not b or a;
    layer4_outputs(5659) <= a;
    layer4_outputs(5660) <= not b;
    layer4_outputs(5661) <= not b or a;
    layer4_outputs(5662) <= b;
    layer4_outputs(5663) <= a and b;
    layer4_outputs(5664) <= a or b;
    layer4_outputs(5665) <= not (a and b);
    layer4_outputs(5666) <= not a or b;
    layer4_outputs(5667) <= '1';
    layer4_outputs(5668) <= a;
    layer4_outputs(5669) <= not a;
    layer4_outputs(5670) <= not a or b;
    layer4_outputs(5671) <= a and not b;
    layer4_outputs(5672) <= '0';
    layer4_outputs(5673) <= a xor b;
    layer4_outputs(5674) <= not a;
    layer4_outputs(5675) <= not b;
    layer4_outputs(5676) <= a xor b;
    layer4_outputs(5677) <= '1';
    layer4_outputs(5678) <= not (a and b);
    layer4_outputs(5679) <= b;
    layer4_outputs(5680) <= '1';
    layer4_outputs(5681) <= not b;
    layer4_outputs(5682) <= a;
    layer4_outputs(5683) <= a;
    layer4_outputs(5684) <= not a;
    layer4_outputs(5685) <= '1';
    layer4_outputs(5686) <= '0';
    layer4_outputs(5687) <= not (a and b);
    layer4_outputs(5688) <= a xor b;
    layer4_outputs(5689) <= not b or a;
    layer4_outputs(5690) <= not b;
    layer4_outputs(5691) <= b and not a;
    layer4_outputs(5692) <= not (a and b);
    layer4_outputs(5693) <= b and not a;
    layer4_outputs(5694) <= a and b;
    layer4_outputs(5695) <= not b;
    layer4_outputs(5696) <= b;
    layer4_outputs(5697) <= not a;
    layer4_outputs(5698) <= not b or a;
    layer4_outputs(5699) <= a;
    layer4_outputs(5700) <= not a;
    layer4_outputs(5701) <= '0';
    layer4_outputs(5702) <= not (a and b);
    layer4_outputs(5703) <= not b or a;
    layer4_outputs(5704) <= not (a or b);
    layer4_outputs(5705) <= b;
    layer4_outputs(5706) <= not b;
    layer4_outputs(5707) <= not (a xor b);
    layer4_outputs(5708) <= a and not b;
    layer4_outputs(5709) <= not a or b;
    layer4_outputs(5710) <= a or b;
    layer4_outputs(5711) <= not b or a;
    layer4_outputs(5712) <= b and not a;
    layer4_outputs(5713) <= b and not a;
    layer4_outputs(5714) <= b;
    layer4_outputs(5715) <= '0';
    layer4_outputs(5716) <= '0';
    layer4_outputs(5717) <= not a;
    layer4_outputs(5718) <= b and not a;
    layer4_outputs(5719) <= b;
    layer4_outputs(5720) <= not (a or b);
    layer4_outputs(5721) <= not a;
    layer4_outputs(5722) <= b and not a;
    layer4_outputs(5723) <= not a;
    layer4_outputs(5724) <= a and not b;
    layer4_outputs(5725) <= not (a or b);
    layer4_outputs(5726) <= b and not a;
    layer4_outputs(5727) <= b;
    layer4_outputs(5728) <= not (a and b);
    layer4_outputs(5729) <= not b;
    layer4_outputs(5730) <= b;
    layer4_outputs(5731) <= not a;
    layer4_outputs(5732) <= b;
    layer4_outputs(5733) <= a;
    layer4_outputs(5734) <= b;
    layer4_outputs(5735) <= a or b;
    layer4_outputs(5736) <= not a;
    layer4_outputs(5737) <= a and not b;
    layer4_outputs(5738) <= not (a xor b);
    layer4_outputs(5739) <= '1';
    layer4_outputs(5740) <= not (a or b);
    layer4_outputs(5741) <= '0';
    layer4_outputs(5742) <= not b;
    layer4_outputs(5743) <= b;
    layer4_outputs(5744) <= a;
    layer4_outputs(5745) <= not (a or b);
    layer4_outputs(5746) <= a or b;
    layer4_outputs(5747) <= a and not b;
    layer4_outputs(5748) <= a or b;
    layer4_outputs(5749) <= a xor b;
    layer4_outputs(5750) <= not b;
    layer4_outputs(5751) <= '0';
    layer4_outputs(5752) <= a;
    layer4_outputs(5753) <= not b or a;
    layer4_outputs(5754) <= not a or b;
    layer4_outputs(5755) <= not (a and b);
    layer4_outputs(5756) <= a;
    layer4_outputs(5757) <= not a;
    layer4_outputs(5758) <= not a;
    layer4_outputs(5759) <= a and b;
    layer4_outputs(5760) <= not (a xor b);
    layer4_outputs(5761) <= '0';
    layer4_outputs(5762) <= a and not b;
    layer4_outputs(5763) <= b;
    layer4_outputs(5764) <= '0';
    layer4_outputs(5765) <= a and not b;
    layer4_outputs(5766) <= a and not b;
    layer4_outputs(5767) <= '0';
    layer4_outputs(5768) <= not b or a;
    layer4_outputs(5769) <= a or b;
    layer4_outputs(5770) <= not (a and b);
    layer4_outputs(5771) <= a and not b;
    layer4_outputs(5772) <= a or b;
    layer4_outputs(5773) <= '0';
    layer4_outputs(5774) <= b and not a;
    layer4_outputs(5775) <= '0';
    layer4_outputs(5776) <= b and not a;
    layer4_outputs(5777) <= a or b;
    layer4_outputs(5778) <= not a or b;
    layer4_outputs(5779) <= not b;
    layer4_outputs(5780) <= a or b;
    layer4_outputs(5781) <= a and b;
    layer4_outputs(5782) <= not (a or b);
    layer4_outputs(5783) <= a;
    layer4_outputs(5784) <= not b or a;
    layer4_outputs(5785) <= a;
    layer4_outputs(5786) <= a;
    layer4_outputs(5787) <= a or b;
    layer4_outputs(5788) <= not (a and b);
    layer4_outputs(5789) <= not (a and b);
    layer4_outputs(5790) <= '0';
    layer4_outputs(5791) <= not b or a;
    layer4_outputs(5792) <= not b;
    layer4_outputs(5793) <= a and not b;
    layer4_outputs(5794) <= not b;
    layer4_outputs(5795) <= a and b;
    layer4_outputs(5796) <= b and not a;
    layer4_outputs(5797) <= not (a and b);
    layer4_outputs(5798) <= '1';
    layer4_outputs(5799) <= not b or a;
    layer4_outputs(5800) <= not a or b;
    layer4_outputs(5801) <= a xor b;
    layer4_outputs(5802) <= b and not a;
    layer4_outputs(5803) <= not (a or b);
    layer4_outputs(5804) <= not (a xor b);
    layer4_outputs(5805) <= a and b;
    layer4_outputs(5806) <= '1';
    layer4_outputs(5807) <= not b;
    layer4_outputs(5808) <= '0';
    layer4_outputs(5809) <= b;
    layer4_outputs(5810) <= '1';
    layer4_outputs(5811) <= a and b;
    layer4_outputs(5812) <= a and not b;
    layer4_outputs(5813) <= a and not b;
    layer4_outputs(5814) <= b;
    layer4_outputs(5815) <= a and b;
    layer4_outputs(5816) <= not a;
    layer4_outputs(5817) <= b;
    layer4_outputs(5818) <= not a or b;
    layer4_outputs(5819) <= not b or a;
    layer4_outputs(5820) <= a;
    layer4_outputs(5821) <= a or b;
    layer4_outputs(5822) <= not (a xor b);
    layer4_outputs(5823) <= not a or b;
    layer4_outputs(5824) <= a;
    layer4_outputs(5825) <= a or b;
    layer4_outputs(5826) <= not b;
    layer4_outputs(5827) <= not (a and b);
    layer4_outputs(5828) <= '0';
    layer4_outputs(5829) <= not b;
    layer4_outputs(5830) <= '1';
    layer4_outputs(5831) <= a and not b;
    layer4_outputs(5832) <= '1';
    layer4_outputs(5833) <= b;
    layer4_outputs(5834) <= b and not a;
    layer4_outputs(5835) <= not b;
    layer4_outputs(5836) <= not b;
    layer4_outputs(5837) <= b;
    layer4_outputs(5838) <= b and not a;
    layer4_outputs(5839) <= '1';
    layer4_outputs(5840) <= a xor b;
    layer4_outputs(5841) <= a and b;
    layer4_outputs(5842) <= '1';
    layer4_outputs(5843) <= b;
    layer4_outputs(5844) <= not (a or b);
    layer4_outputs(5845) <= not (a and b);
    layer4_outputs(5846) <= a and not b;
    layer4_outputs(5847) <= not (a or b);
    layer4_outputs(5848) <= a and b;
    layer4_outputs(5849) <= a;
    layer4_outputs(5850) <= b;
    layer4_outputs(5851) <= '1';
    layer4_outputs(5852) <= '1';
    layer4_outputs(5853) <= not b;
    layer4_outputs(5854) <= '0';
    layer4_outputs(5855) <= not a or b;
    layer4_outputs(5856) <= not b;
    layer4_outputs(5857) <= '0';
    layer4_outputs(5858) <= not a or b;
    layer4_outputs(5859) <= not (a and b);
    layer4_outputs(5860) <= not a or b;
    layer4_outputs(5861) <= a or b;
    layer4_outputs(5862) <= not (a or b);
    layer4_outputs(5863) <= not b;
    layer4_outputs(5864) <= not a;
    layer4_outputs(5865) <= a and b;
    layer4_outputs(5866) <= not b;
    layer4_outputs(5867) <= a xor b;
    layer4_outputs(5868) <= a xor b;
    layer4_outputs(5869) <= a and b;
    layer4_outputs(5870) <= b;
    layer4_outputs(5871) <= a and b;
    layer4_outputs(5872) <= not (a or b);
    layer4_outputs(5873) <= a and b;
    layer4_outputs(5874) <= not a or b;
    layer4_outputs(5875) <= not (a or b);
    layer4_outputs(5876) <= not (a or b);
    layer4_outputs(5877) <= not (a or b);
    layer4_outputs(5878) <= not (a xor b);
    layer4_outputs(5879) <= '1';
    layer4_outputs(5880) <= not b;
    layer4_outputs(5881) <= not (a or b);
    layer4_outputs(5882) <= a or b;
    layer4_outputs(5883) <= not a or b;
    layer4_outputs(5884) <= not b;
    layer4_outputs(5885) <= not b or a;
    layer4_outputs(5886) <= not (a or b);
    layer4_outputs(5887) <= b and not a;
    layer4_outputs(5888) <= not (a or b);
    layer4_outputs(5889) <= a and not b;
    layer4_outputs(5890) <= not a or b;
    layer4_outputs(5891) <= not b;
    layer4_outputs(5892) <= not (a and b);
    layer4_outputs(5893) <= b;
    layer4_outputs(5894) <= a or b;
    layer4_outputs(5895) <= a;
    layer4_outputs(5896) <= b;
    layer4_outputs(5897) <= not a;
    layer4_outputs(5898) <= '1';
    layer4_outputs(5899) <= a;
    layer4_outputs(5900) <= a and not b;
    layer4_outputs(5901) <= not a or b;
    layer4_outputs(5902) <= a and not b;
    layer4_outputs(5903) <= not (a and b);
    layer4_outputs(5904) <= not (a or b);
    layer4_outputs(5905) <= b;
    layer4_outputs(5906) <= b;
    layer4_outputs(5907) <= not a;
    layer4_outputs(5908) <= not (a or b);
    layer4_outputs(5909) <= not a;
    layer4_outputs(5910) <= a and b;
    layer4_outputs(5911) <= not (a and b);
    layer4_outputs(5912) <= not a;
    layer4_outputs(5913) <= not a;
    layer4_outputs(5914) <= not a;
    layer4_outputs(5915) <= a and b;
    layer4_outputs(5916) <= not b;
    layer4_outputs(5917) <= not (a or b);
    layer4_outputs(5918) <= not b;
    layer4_outputs(5919) <= not (a or b);
    layer4_outputs(5920) <= not (a or b);
    layer4_outputs(5921) <= not a;
    layer4_outputs(5922) <= not a or b;
    layer4_outputs(5923) <= a and b;
    layer4_outputs(5924) <= b;
    layer4_outputs(5925) <= not a;
    layer4_outputs(5926) <= not (a and b);
    layer4_outputs(5927) <= not b or a;
    layer4_outputs(5928) <= a;
    layer4_outputs(5929) <= a and not b;
    layer4_outputs(5930) <= a or b;
    layer4_outputs(5931) <= not b;
    layer4_outputs(5932) <= not (a and b);
    layer4_outputs(5933) <= b;
    layer4_outputs(5934) <= not a or b;
    layer4_outputs(5935) <= not b or a;
    layer4_outputs(5936) <= not a;
    layer4_outputs(5937) <= a or b;
    layer4_outputs(5938) <= a or b;
    layer4_outputs(5939) <= a;
    layer4_outputs(5940) <= '1';
    layer4_outputs(5941) <= '1';
    layer4_outputs(5942) <= a;
    layer4_outputs(5943) <= not (a or b);
    layer4_outputs(5944) <= not a;
    layer4_outputs(5945) <= not b;
    layer4_outputs(5946) <= '1';
    layer4_outputs(5947) <= not (a and b);
    layer4_outputs(5948) <= b and not a;
    layer4_outputs(5949) <= a or b;
    layer4_outputs(5950) <= a or b;
    layer4_outputs(5951) <= b;
    layer4_outputs(5952) <= not a or b;
    layer4_outputs(5953) <= b and not a;
    layer4_outputs(5954) <= b;
    layer4_outputs(5955) <= not a or b;
    layer4_outputs(5956) <= a or b;
    layer4_outputs(5957) <= a and b;
    layer4_outputs(5958) <= not b;
    layer4_outputs(5959) <= not b;
    layer4_outputs(5960) <= a;
    layer4_outputs(5961) <= not b;
    layer4_outputs(5962) <= '1';
    layer4_outputs(5963) <= a;
    layer4_outputs(5964) <= '1';
    layer4_outputs(5965) <= not a;
    layer4_outputs(5966) <= not (a and b);
    layer4_outputs(5967) <= not a;
    layer4_outputs(5968) <= not a or b;
    layer4_outputs(5969) <= b and not a;
    layer4_outputs(5970) <= not (a or b);
    layer4_outputs(5971) <= not a;
    layer4_outputs(5972) <= '0';
    layer4_outputs(5973) <= b;
    layer4_outputs(5974) <= '1';
    layer4_outputs(5975) <= not a or b;
    layer4_outputs(5976) <= not a or b;
    layer4_outputs(5977) <= not a;
    layer4_outputs(5978) <= a xor b;
    layer4_outputs(5979) <= not (a and b);
    layer4_outputs(5980) <= not b;
    layer4_outputs(5981) <= b and not a;
    layer4_outputs(5982) <= not (a or b);
    layer4_outputs(5983) <= not a;
    layer4_outputs(5984) <= not a;
    layer4_outputs(5985) <= a and not b;
    layer4_outputs(5986) <= a and not b;
    layer4_outputs(5987) <= a and b;
    layer4_outputs(5988) <= a;
    layer4_outputs(5989) <= '0';
    layer4_outputs(5990) <= b and not a;
    layer4_outputs(5991) <= a and b;
    layer4_outputs(5992) <= a xor b;
    layer4_outputs(5993) <= not (a or b);
    layer4_outputs(5994) <= b;
    layer4_outputs(5995) <= '0';
    layer4_outputs(5996) <= '1';
    layer4_outputs(5997) <= a and b;
    layer4_outputs(5998) <= a;
    layer4_outputs(5999) <= a or b;
    layer4_outputs(6000) <= a and b;
    layer4_outputs(6001) <= '0';
    layer4_outputs(6002) <= not (a and b);
    layer4_outputs(6003) <= not b;
    layer4_outputs(6004) <= not b;
    layer4_outputs(6005) <= not (a and b);
    layer4_outputs(6006) <= a and not b;
    layer4_outputs(6007) <= not a;
    layer4_outputs(6008) <= not a;
    layer4_outputs(6009) <= not b;
    layer4_outputs(6010) <= not b;
    layer4_outputs(6011) <= b and not a;
    layer4_outputs(6012) <= not (a or b);
    layer4_outputs(6013) <= not (a and b);
    layer4_outputs(6014) <= '1';
    layer4_outputs(6015) <= not b;
    layer4_outputs(6016) <= not (a or b);
    layer4_outputs(6017) <= b and not a;
    layer4_outputs(6018) <= a or b;
    layer4_outputs(6019) <= '1';
    layer4_outputs(6020) <= not (a or b);
    layer4_outputs(6021) <= a;
    layer4_outputs(6022) <= b;
    layer4_outputs(6023) <= not b;
    layer4_outputs(6024) <= a and b;
    layer4_outputs(6025) <= not (a or b);
    layer4_outputs(6026) <= a;
    layer4_outputs(6027) <= not (a or b);
    layer4_outputs(6028) <= not (a and b);
    layer4_outputs(6029) <= not b or a;
    layer4_outputs(6030) <= not a or b;
    layer4_outputs(6031) <= a;
    layer4_outputs(6032) <= a;
    layer4_outputs(6033) <= a and b;
    layer4_outputs(6034) <= not a;
    layer4_outputs(6035) <= not b;
    layer4_outputs(6036) <= not b;
    layer4_outputs(6037) <= a and b;
    layer4_outputs(6038) <= b and not a;
    layer4_outputs(6039) <= not (a and b);
    layer4_outputs(6040) <= not (a or b);
    layer4_outputs(6041) <= '1';
    layer4_outputs(6042) <= b and not a;
    layer4_outputs(6043) <= '1';
    layer4_outputs(6044) <= a and b;
    layer4_outputs(6045) <= not b;
    layer4_outputs(6046) <= a or b;
    layer4_outputs(6047) <= a;
    layer4_outputs(6048) <= not (a and b);
    layer4_outputs(6049) <= not b or a;
    layer4_outputs(6050) <= a and b;
    layer4_outputs(6051) <= not b or a;
    layer4_outputs(6052) <= not (a or b);
    layer4_outputs(6053) <= a and b;
    layer4_outputs(6054) <= not a or b;
    layer4_outputs(6055) <= not a or b;
    layer4_outputs(6056) <= a or b;
    layer4_outputs(6057) <= a and b;
    layer4_outputs(6058) <= not b;
    layer4_outputs(6059) <= not b or a;
    layer4_outputs(6060) <= not b;
    layer4_outputs(6061) <= b;
    layer4_outputs(6062) <= not a;
    layer4_outputs(6063) <= a and b;
    layer4_outputs(6064) <= a and b;
    layer4_outputs(6065) <= b and not a;
    layer4_outputs(6066) <= a or b;
    layer4_outputs(6067) <= not (a xor b);
    layer4_outputs(6068) <= a and not b;
    layer4_outputs(6069) <= not b;
    layer4_outputs(6070) <= b and not a;
    layer4_outputs(6071) <= a or b;
    layer4_outputs(6072) <= not (a or b);
    layer4_outputs(6073) <= not (a or b);
    layer4_outputs(6074) <= not a or b;
    layer4_outputs(6075) <= not b or a;
    layer4_outputs(6076) <= a and not b;
    layer4_outputs(6077) <= not a;
    layer4_outputs(6078) <= a and b;
    layer4_outputs(6079) <= a and not b;
    layer4_outputs(6080) <= not b;
    layer4_outputs(6081) <= '1';
    layer4_outputs(6082) <= a;
    layer4_outputs(6083) <= a and b;
    layer4_outputs(6084) <= a and b;
    layer4_outputs(6085) <= b;
    layer4_outputs(6086) <= a or b;
    layer4_outputs(6087) <= not (a xor b);
    layer4_outputs(6088) <= b;
    layer4_outputs(6089) <= a and b;
    layer4_outputs(6090) <= a and b;
    layer4_outputs(6091) <= not a or b;
    layer4_outputs(6092) <= not a or b;
    layer4_outputs(6093) <= '1';
    layer4_outputs(6094) <= not b;
    layer4_outputs(6095) <= not b or a;
    layer4_outputs(6096) <= b;
    layer4_outputs(6097) <= a and b;
    layer4_outputs(6098) <= a and not b;
    layer4_outputs(6099) <= not b;
    layer4_outputs(6100) <= a and not b;
    layer4_outputs(6101) <= b and not a;
    layer4_outputs(6102) <= '1';
    layer4_outputs(6103) <= not a;
    layer4_outputs(6104) <= a or b;
    layer4_outputs(6105) <= a and b;
    layer4_outputs(6106) <= b;
    layer4_outputs(6107) <= '1';
    layer4_outputs(6108) <= not a or b;
    layer4_outputs(6109) <= a and not b;
    layer4_outputs(6110) <= a or b;
    layer4_outputs(6111) <= not b;
    layer4_outputs(6112) <= a and b;
    layer4_outputs(6113) <= '1';
    layer4_outputs(6114) <= a and b;
    layer4_outputs(6115) <= not b;
    layer4_outputs(6116) <= b and not a;
    layer4_outputs(6117) <= not a or b;
    layer4_outputs(6118) <= b and not a;
    layer4_outputs(6119) <= b;
    layer4_outputs(6120) <= not a;
    layer4_outputs(6121) <= '0';
    layer4_outputs(6122) <= '0';
    layer4_outputs(6123) <= b;
    layer4_outputs(6124) <= a and b;
    layer4_outputs(6125) <= '1';
    layer4_outputs(6126) <= not b;
    layer4_outputs(6127) <= '1';
    layer4_outputs(6128) <= a;
    layer4_outputs(6129) <= not (a or b);
    layer4_outputs(6130) <= b and not a;
    layer4_outputs(6131) <= a and not b;
    layer4_outputs(6132) <= a or b;
    layer4_outputs(6133) <= not a or b;
    layer4_outputs(6134) <= not b;
    layer4_outputs(6135) <= not a;
    layer4_outputs(6136) <= a and b;
    layer4_outputs(6137) <= a xor b;
    layer4_outputs(6138) <= not a;
    layer4_outputs(6139) <= a xor b;
    layer4_outputs(6140) <= not (a xor b);
    layer4_outputs(6141) <= not b or a;
    layer4_outputs(6142) <= not (a and b);
    layer4_outputs(6143) <= not a;
    layer4_outputs(6144) <= not a;
    layer4_outputs(6145) <= a xor b;
    layer4_outputs(6146) <= not (a or b);
    layer4_outputs(6147) <= not b or a;
    layer4_outputs(6148) <= '1';
    layer4_outputs(6149) <= a or b;
    layer4_outputs(6150) <= not b;
    layer4_outputs(6151) <= not (a and b);
    layer4_outputs(6152) <= not a or b;
    layer4_outputs(6153) <= not a;
    layer4_outputs(6154) <= not a;
    layer4_outputs(6155) <= '1';
    layer4_outputs(6156) <= not b;
    layer4_outputs(6157) <= a or b;
    layer4_outputs(6158) <= not a;
    layer4_outputs(6159) <= a;
    layer4_outputs(6160) <= not (a and b);
    layer4_outputs(6161) <= not a;
    layer4_outputs(6162) <= a and b;
    layer4_outputs(6163) <= a and b;
    layer4_outputs(6164) <= not (a or b);
    layer4_outputs(6165) <= not b or a;
    layer4_outputs(6166) <= b;
    layer4_outputs(6167) <= a and not b;
    layer4_outputs(6168) <= not b;
    layer4_outputs(6169) <= a xor b;
    layer4_outputs(6170) <= a and not b;
    layer4_outputs(6171) <= not a or b;
    layer4_outputs(6172) <= not b;
    layer4_outputs(6173) <= a and b;
    layer4_outputs(6174) <= not (a and b);
    layer4_outputs(6175) <= not (a xor b);
    layer4_outputs(6176) <= a and b;
    layer4_outputs(6177) <= b;
    layer4_outputs(6178) <= b;
    layer4_outputs(6179) <= b and not a;
    layer4_outputs(6180) <= not (a or b);
    layer4_outputs(6181) <= not b;
    layer4_outputs(6182) <= not a;
    layer4_outputs(6183) <= b and not a;
    layer4_outputs(6184) <= not b;
    layer4_outputs(6185) <= not a;
    layer4_outputs(6186) <= not b or a;
    layer4_outputs(6187) <= not b or a;
    layer4_outputs(6188) <= a or b;
    layer4_outputs(6189) <= a xor b;
    layer4_outputs(6190) <= a;
    layer4_outputs(6191) <= a;
    layer4_outputs(6192) <= b;
    layer4_outputs(6193) <= not (a and b);
    layer4_outputs(6194) <= not b or a;
    layer4_outputs(6195) <= a and b;
    layer4_outputs(6196) <= a and b;
    layer4_outputs(6197) <= not (a and b);
    layer4_outputs(6198) <= not a or b;
    layer4_outputs(6199) <= a or b;
    layer4_outputs(6200) <= not a or b;
    layer4_outputs(6201) <= not (a or b);
    layer4_outputs(6202) <= a;
    layer4_outputs(6203) <= a and not b;
    layer4_outputs(6204) <= a and b;
    layer4_outputs(6205) <= not a or b;
    layer4_outputs(6206) <= a or b;
    layer4_outputs(6207) <= b;
    layer4_outputs(6208) <= not a;
    layer4_outputs(6209) <= b and not a;
    layer4_outputs(6210) <= not a;
    layer4_outputs(6211) <= b;
    layer4_outputs(6212) <= not b;
    layer4_outputs(6213) <= not a;
    layer4_outputs(6214) <= not a or b;
    layer4_outputs(6215) <= b;
    layer4_outputs(6216) <= b and not a;
    layer4_outputs(6217) <= not a;
    layer4_outputs(6218) <= a and b;
    layer4_outputs(6219) <= b;
    layer4_outputs(6220) <= b and not a;
    layer4_outputs(6221) <= b;
    layer4_outputs(6222) <= a or b;
    layer4_outputs(6223) <= b;
    layer4_outputs(6224) <= not (a and b);
    layer4_outputs(6225) <= a;
    layer4_outputs(6226) <= not (a xor b);
    layer4_outputs(6227) <= a and b;
    layer4_outputs(6228) <= a;
    layer4_outputs(6229) <= '1';
    layer4_outputs(6230) <= a and not b;
    layer4_outputs(6231) <= not (a and b);
    layer4_outputs(6232) <= a and b;
    layer4_outputs(6233) <= '0';
    layer4_outputs(6234) <= not b;
    layer4_outputs(6235) <= b;
    layer4_outputs(6236) <= not a or b;
    layer4_outputs(6237) <= not (a and b);
    layer4_outputs(6238) <= not a;
    layer4_outputs(6239) <= '0';
    layer4_outputs(6240) <= b;
    layer4_outputs(6241) <= not b or a;
    layer4_outputs(6242) <= not a or b;
    layer4_outputs(6243) <= not b or a;
    layer4_outputs(6244) <= '1';
    layer4_outputs(6245) <= b and not a;
    layer4_outputs(6246) <= not (a or b);
    layer4_outputs(6247) <= b;
    layer4_outputs(6248) <= a or b;
    layer4_outputs(6249) <= not (a and b);
    layer4_outputs(6250) <= b;
    layer4_outputs(6251) <= a xor b;
    layer4_outputs(6252) <= not b or a;
    layer4_outputs(6253) <= not (a and b);
    layer4_outputs(6254) <= b and not a;
    layer4_outputs(6255) <= not b;
    layer4_outputs(6256) <= a and b;
    layer4_outputs(6257) <= not (a and b);
    layer4_outputs(6258) <= b;
    layer4_outputs(6259) <= '1';
    layer4_outputs(6260) <= not a;
    layer4_outputs(6261) <= a xor b;
    layer4_outputs(6262) <= b and not a;
    layer4_outputs(6263) <= not b;
    layer4_outputs(6264) <= a and b;
    layer4_outputs(6265) <= not (a and b);
    layer4_outputs(6266) <= not (a xor b);
    layer4_outputs(6267) <= a and b;
    layer4_outputs(6268) <= b;
    layer4_outputs(6269) <= not a;
    layer4_outputs(6270) <= a and b;
    layer4_outputs(6271) <= '1';
    layer4_outputs(6272) <= not (a and b);
    layer4_outputs(6273) <= not (a and b);
    layer4_outputs(6274) <= not (a and b);
    layer4_outputs(6275) <= '1';
    layer4_outputs(6276) <= b and not a;
    layer4_outputs(6277) <= not (a xor b);
    layer4_outputs(6278) <= b and not a;
    layer4_outputs(6279) <= b;
    layer4_outputs(6280) <= not b;
    layer4_outputs(6281) <= not a;
    layer4_outputs(6282) <= not a or b;
    layer4_outputs(6283) <= a;
    layer4_outputs(6284) <= a or b;
    layer4_outputs(6285) <= a or b;
    layer4_outputs(6286) <= not (a and b);
    layer4_outputs(6287) <= a and not b;
    layer4_outputs(6288) <= a;
    layer4_outputs(6289) <= not b or a;
    layer4_outputs(6290) <= b;
    layer4_outputs(6291) <= b;
    layer4_outputs(6292) <= a and b;
    layer4_outputs(6293) <= a and not b;
    layer4_outputs(6294) <= a or b;
    layer4_outputs(6295) <= a;
    layer4_outputs(6296) <= a and b;
    layer4_outputs(6297) <= not (a xor b);
    layer4_outputs(6298) <= not a or b;
    layer4_outputs(6299) <= b;
    layer4_outputs(6300) <= not a or b;
    layer4_outputs(6301) <= a xor b;
    layer4_outputs(6302) <= not b;
    layer4_outputs(6303) <= not a or b;
    layer4_outputs(6304) <= '1';
    layer4_outputs(6305) <= not (a and b);
    layer4_outputs(6306) <= '0';
    layer4_outputs(6307) <= b;
    layer4_outputs(6308) <= not a or b;
    layer4_outputs(6309) <= not b or a;
    layer4_outputs(6310) <= not b;
    layer4_outputs(6311) <= a;
    layer4_outputs(6312) <= a and not b;
    layer4_outputs(6313) <= a and not b;
    layer4_outputs(6314) <= not a or b;
    layer4_outputs(6315) <= a and b;
    layer4_outputs(6316) <= '0';
    layer4_outputs(6317) <= b;
    layer4_outputs(6318) <= not a;
    layer4_outputs(6319) <= not a or b;
    layer4_outputs(6320) <= a or b;
    layer4_outputs(6321) <= not (a or b);
    layer4_outputs(6322) <= '0';
    layer4_outputs(6323) <= not b or a;
    layer4_outputs(6324) <= b and not a;
    layer4_outputs(6325) <= b and not a;
    layer4_outputs(6326) <= not (a or b);
    layer4_outputs(6327) <= not (a and b);
    layer4_outputs(6328) <= a and not b;
    layer4_outputs(6329) <= '0';
    layer4_outputs(6330) <= not a or b;
    layer4_outputs(6331) <= a and not b;
    layer4_outputs(6332) <= b;
    layer4_outputs(6333) <= a;
    layer4_outputs(6334) <= not a or b;
    layer4_outputs(6335) <= a or b;
    layer4_outputs(6336) <= not b or a;
    layer4_outputs(6337) <= not a or b;
    layer4_outputs(6338) <= not a;
    layer4_outputs(6339) <= a and b;
    layer4_outputs(6340) <= not (a or b);
    layer4_outputs(6341) <= a;
    layer4_outputs(6342) <= a xor b;
    layer4_outputs(6343) <= '1';
    layer4_outputs(6344) <= not a or b;
    layer4_outputs(6345) <= not (a or b);
    layer4_outputs(6346) <= not a;
    layer4_outputs(6347) <= not b;
    layer4_outputs(6348) <= not (a or b);
    layer4_outputs(6349) <= b and not a;
    layer4_outputs(6350) <= a;
    layer4_outputs(6351) <= not a;
    layer4_outputs(6352) <= a and b;
    layer4_outputs(6353) <= a;
    layer4_outputs(6354) <= not b or a;
    layer4_outputs(6355) <= a and b;
    layer4_outputs(6356) <= b;
    layer4_outputs(6357) <= '0';
    layer4_outputs(6358) <= '1';
    layer4_outputs(6359) <= '1';
    layer4_outputs(6360) <= a;
    layer4_outputs(6361) <= a and b;
    layer4_outputs(6362) <= not b;
    layer4_outputs(6363) <= '0';
    layer4_outputs(6364) <= not b;
    layer4_outputs(6365) <= not (a and b);
    layer4_outputs(6366) <= not b or a;
    layer4_outputs(6367) <= '1';
    layer4_outputs(6368) <= not (a or b);
    layer4_outputs(6369) <= not (a and b);
    layer4_outputs(6370) <= b and not a;
    layer4_outputs(6371) <= b and not a;
    layer4_outputs(6372) <= not b;
    layer4_outputs(6373) <= b;
    layer4_outputs(6374) <= a and not b;
    layer4_outputs(6375) <= a xor b;
    layer4_outputs(6376) <= not a;
    layer4_outputs(6377) <= a and not b;
    layer4_outputs(6378) <= not (a or b);
    layer4_outputs(6379) <= a and not b;
    layer4_outputs(6380) <= not (a xor b);
    layer4_outputs(6381) <= a;
    layer4_outputs(6382) <= not a or b;
    layer4_outputs(6383) <= a;
    layer4_outputs(6384) <= b;
    layer4_outputs(6385) <= b;
    layer4_outputs(6386) <= not a or b;
    layer4_outputs(6387) <= a and b;
    layer4_outputs(6388) <= not a;
    layer4_outputs(6389) <= a;
    layer4_outputs(6390) <= not a or b;
    layer4_outputs(6391) <= b and not a;
    layer4_outputs(6392) <= b;
    layer4_outputs(6393) <= not (a and b);
    layer4_outputs(6394) <= '1';
    layer4_outputs(6395) <= b;
    layer4_outputs(6396) <= a or b;
    layer4_outputs(6397) <= not a or b;
    layer4_outputs(6398) <= b;
    layer4_outputs(6399) <= a or b;
    layer4_outputs(6400) <= b;
    layer4_outputs(6401) <= '1';
    layer4_outputs(6402) <= not b;
    layer4_outputs(6403) <= a xor b;
    layer4_outputs(6404) <= a;
    layer4_outputs(6405) <= a and b;
    layer4_outputs(6406) <= not b;
    layer4_outputs(6407) <= not b;
    layer4_outputs(6408) <= b and not a;
    layer4_outputs(6409) <= a xor b;
    layer4_outputs(6410) <= not a;
    layer4_outputs(6411) <= a;
    layer4_outputs(6412) <= not (a or b);
    layer4_outputs(6413) <= not (a or b);
    layer4_outputs(6414) <= a;
    layer4_outputs(6415) <= a and not b;
    layer4_outputs(6416) <= not (a xor b);
    layer4_outputs(6417) <= a and not b;
    layer4_outputs(6418) <= a xor b;
    layer4_outputs(6419) <= b;
    layer4_outputs(6420) <= not a;
    layer4_outputs(6421) <= not (a or b);
    layer4_outputs(6422) <= a or b;
    layer4_outputs(6423) <= a;
    layer4_outputs(6424) <= not a or b;
    layer4_outputs(6425) <= not a or b;
    layer4_outputs(6426) <= b and not a;
    layer4_outputs(6427) <= b and not a;
    layer4_outputs(6428) <= not (a and b);
    layer4_outputs(6429) <= '0';
    layer4_outputs(6430) <= a and not b;
    layer4_outputs(6431) <= a and b;
    layer4_outputs(6432) <= a xor b;
    layer4_outputs(6433) <= not (a xor b);
    layer4_outputs(6434) <= not a;
    layer4_outputs(6435) <= '0';
    layer4_outputs(6436) <= not a or b;
    layer4_outputs(6437) <= b and not a;
    layer4_outputs(6438) <= not (a and b);
    layer4_outputs(6439) <= b and not a;
    layer4_outputs(6440) <= a or b;
    layer4_outputs(6441) <= not b or a;
    layer4_outputs(6442) <= not a;
    layer4_outputs(6443) <= not (a or b);
    layer4_outputs(6444) <= not (a or b);
    layer4_outputs(6445) <= a;
    layer4_outputs(6446) <= a and b;
    layer4_outputs(6447) <= a xor b;
    layer4_outputs(6448) <= not a or b;
    layer4_outputs(6449) <= a;
    layer4_outputs(6450) <= b;
    layer4_outputs(6451) <= not b or a;
    layer4_outputs(6452) <= b and not a;
    layer4_outputs(6453) <= '1';
    layer4_outputs(6454) <= b and not a;
    layer4_outputs(6455) <= '0';
    layer4_outputs(6456) <= not b;
    layer4_outputs(6457) <= not a or b;
    layer4_outputs(6458) <= a and not b;
    layer4_outputs(6459) <= not a;
    layer4_outputs(6460) <= not a;
    layer4_outputs(6461) <= not b;
    layer4_outputs(6462) <= a and not b;
    layer4_outputs(6463) <= a and b;
    layer4_outputs(6464) <= not a or b;
    layer4_outputs(6465) <= b;
    layer4_outputs(6466) <= not a or b;
    layer4_outputs(6467) <= not b;
    layer4_outputs(6468) <= a;
    layer4_outputs(6469) <= a and not b;
    layer4_outputs(6470) <= a or b;
    layer4_outputs(6471) <= a and not b;
    layer4_outputs(6472) <= not (a and b);
    layer4_outputs(6473) <= b and not a;
    layer4_outputs(6474) <= a and not b;
    layer4_outputs(6475) <= not a or b;
    layer4_outputs(6476) <= a;
    layer4_outputs(6477) <= a or b;
    layer4_outputs(6478) <= not a;
    layer4_outputs(6479) <= not b;
    layer4_outputs(6480) <= not b or a;
    layer4_outputs(6481) <= b;
    layer4_outputs(6482) <= a;
    layer4_outputs(6483) <= a;
    layer4_outputs(6484) <= '1';
    layer4_outputs(6485) <= a xor b;
    layer4_outputs(6486) <= '0';
    layer4_outputs(6487) <= a or b;
    layer4_outputs(6488) <= not a or b;
    layer4_outputs(6489) <= a xor b;
    layer4_outputs(6490) <= b;
    layer4_outputs(6491) <= not (a and b);
    layer4_outputs(6492) <= a and b;
    layer4_outputs(6493) <= a and not b;
    layer4_outputs(6494) <= b and not a;
    layer4_outputs(6495) <= not a or b;
    layer4_outputs(6496) <= not a;
    layer4_outputs(6497) <= not a or b;
    layer4_outputs(6498) <= not a;
    layer4_outputs(6499) <= a;
    layer4_outputs(6500) <= a and not b;
    layer4_outputs(6501) <= a or b;
    layer4_outputs(6502) <= not (a and b);
    layer4_outputs(6503) <= a and b;
    layer4_outputs(6504) <= a;
    layer4_outputs(6505) <= a;
    layer4_outputs(6506) <= a or b;
    layer4_outputs(6507) <= b and not a;
    layer4_outputs(6508) <= '1';
    layer4_outputs(6509) <= not (a and b);
    layer4_outputs(6510) <= a xor b;
    layer4_outputs(6511) <= not (a or b);
    layer4_outputs(6512) <= not (a or b);
    layer4_outputs(6513) <= not a;
    layer4_outputs(6514) <= '1';
    layer4_outputs(6515) <= not b or a;
    layer4_outputs(6516) <= '1';
    layer4_outputs(6517) <= a and not b;
    layer4_outputs(6518) <= a and b;
    layer4_outputs(6519) <= a or b;
    layer4_outputs(6520) <= not (a and b);
    layer4_outputs(6521) <= a;
    layer4_outputs(6522) <= not b;
    layer4_outputs(6523) <= '1';
    layer4_outputs(6524) <= a xor b;
    layer4_outputs(6525) <= b;
    layer4_outputs(6526) <= not b;
    layer4_outputs(6527) <= '0';
    layer4_outputs(6528) <= a and not b;
    layer4_outputs(6529) <= a and b;
    layer4_outputs(6530) <= not a;
    layer4_outputs(6531) <= a;
    layer4_outputs(6532) <= not (a xor b);
    layer4_outputs(6533) <= a;
    layer4_outputs(6534) <= not (a and b);
    layer4_outputs(6535) <= not b or a;
    layer4_outputs(6536) <= a;
    layer4_outputs(6537) <= not (a or b);
    layer4_outputs(6538) <= not a or b;
    layer4_outputs(6539) <= b;
    layer4_outputs(6540) <= '1';
    layer4_outputs(6541) <= b;
    layer4_outputs(6542) <= not b or a;
    layer4_outputs(6543) <= b and not a;
    layer4_outputs(6544) <= not (a xor b);
    layer4_outputs(6545) <= not a or b;
    layer4_outputs(6546) <= a and not b;
    layer4_outputs(6547) <= b and not a;
    layer4_outputs(6548) <= not b;
    layer4_outputs(6549) <= not (a and b);
    layer4_outputs(6550) <= '0';
    layer4_outputs(6551) <= not b or a;
    layer4_outputs(6552) <= '1';
    layer4_outputs(6553) <= '0';
    layer4_outputs(6554) <= a and not b;
    layer4_outputs(6555) <= b;
    layer4_outputs(6556) <= not b;
    layer4_outputs(6557) <= not (a or b);
    layer4_outputs(6558) <= a xor b;
    layer4_outputs(6559) <= not (a or b);
    layer4_outputs(6560) <= not b;
    layer4_outputs(6561) <= not b;
    layer4_outputs(6562) <= a or b;
    layer4_outputs(6563) <= not (a or b);
    layer4_outputs(6564) <= '0';
    layer4_outputs(6565) <= a or b;
    layer4_outputs(6566) <= not a or b;
    layer4_outputs(6567) <= not a or b;
    layer4_outputs(6568) <= not (a or b);
    layer4_outputs(6569) <= '0';
    layer4_outputs(6570) <= not (a xor b);
    layer4_outputs(6571) <= a and b;
    layer4_outputs(6572) <= a and not b;
    layer4_outputs(6573) <= not b or a;
    layer4_outputs(6574) <= a and not b;
    layer4_outputs(6575) <= not b or a;
    layer4_outputs(6576) <= b;
    layer4_outputs(6577) <= not b;
    layer4_outputs(6578) <= a and b;
    layer4_outputs(6579) <= a and b;
    layer4_outputs(6580) <= not (a or b);
    layer4_outputs(6581) <= '0';
    layer4_outputs(6582) <= a and not b;
    layer4_outputs(6583) <= not (a and b);
    layer4_outputs(6584) <= b and not a;
    layer4_outputs(6585) <= not (a and b);
    layer4_outputs(6586) <= b;
    layer4_outputs(6587) <= not b;
    layer4_outputs(6588) <= not (a and b);
    layer4_outputs(6589) <= not a;
    layer4_outputs(6590) <= not (a or b);
    layer4_outputs(6591) <= '0';
    layer4_outputs(6592) <= b and not a;
    layer4_outputs(6593) <= a and not b;
    layer4_outputs(6594) <= '0';
    layer4_outputs(6595) <= not a or b;
    layer4_outputs(6596) <= not a or b;
    layer4_outputs(6597) <= '1';
    layer4_outputs(6598) <= b;
    layer4_outputs(6599) <= b;
    layer4_outputs(6600) <= not (a or b);
    layer4_outputs(6601) <= not (a and b);
    layer4_outputs(6602) <= '1';
    layer4_outputs(6603) <= not a;
    layer4_outputs(6604) <= not a or b;
    layer4_outputs(6605) <= not b or a;
    layer4_outputs(6606) <= a or b;
    layer4_outputs(6607) <= not b;
    layer4_outputs(6608) <= not b or a;
    layer4_outputs(6609) <= '0';
    layer4_outputs(6610) <= '1';
    layer4_outputs(6611) <= b and not a;
    layer4_outputs(6612) <= not b or a;
    layer4_outputs(6613) <= not a;
    layer4_outputs(6614) <= a and not b;
    layer4_outputs(6615) <= b;
    layer4_outputs(6616) <= not (a or b);
    layer4_outputs(6617) <= a and not b;
    layer4_outputs(6618) <= b and not a;
    layer4_outputs(6619) <= not a;
    layer4_outputs(6620) <= a xor b;
    layer4_outputs(6621) <= a;
    layer4_outputs(6622) <= '0';
    layer4_outputs(6623) <= not a;
    layer4_outputs(6624) <= not (a and b);
    layer4_outputs(6625) <= a and not b;
    layer4_outputs(6626) <= not b;
    layer4_outputs(6627) <= b;
    layer4_outputs(6628) <= not (a or b);
    layer4_outputs(6629) <= b;
    layer4_outputs(6630) <= not a or b;
    layer4_outputs(6631) <= not b;
    layer4_outputs(6632) <= not b or a;
    layer4_outputs(6633) <= not a or b;
    layer4_outputs(6634) <= not b or a;
    layer4_outputs(6635) <= a or b;
    layer4_outputs(6636) <= '0';
    layer4_outputs(6637) <= b and not a;
    layer4_outputs(6638) <= not a;
    layer4_outputs(6639) <= not a;
    layer4_outputs(6640) <= not b;
    layer4_outputs(6641) <= b and not a;
    layer4_outputs(6642) <= a;
    layer4_outputs(6643) <= a;
    layer4_outputs(6644) <= a;
    layer4_outputs(6645) <= not a;
    layer4_outputs(6646) <= not b or a;
    layer4_outputs(6647) <= not (a and b);
    layer4_outputs(6648) <= not (a or b);
    layer4_outputs(6649) <= not a;
    layer4_outputs(6650) <= a and b;
    layer4_outputs(6651) <= a or b;
    layer4_outputs(6652) <= not b;
    layer4_outputs(6653) <= not b or a;
    layer4_outputs(6654) <= a;
    layer4_outputs(6655) <= not a;
    layer4_outputs(6656) <= not a;
    layer4_outputs(6657) <= a or b;
    layer4_outputs(6658) <= b and not a;
    layer4_outputs(6659) <= not b;
    layer4_outputs(6660) <= not b or a;
    layer4_outputs(6661) <= a;
    layer4_outputs(6662) <= b;
    layer4_outputs(6663) <= not (a and b);
    layer4_outputs(6664) <= a or b;
    layer4_outputs(6665) <= a or b;
    layer4_outputs(6666) <= '1';
    layer4_outputs(6667) <= b;
    layer4_outputs(6668) <= a;
    layer4_outputs(6669) <= not (a and b);
    layer4_outputs(6670) <= a or b;
    layer4_outputs(6671) <= b;
    layer4_outputs(6672) <= a;
    layer4_outputs(6673) <= not b or a;
    layer4_outputs(6674) <= a;
    layer4_outputs(6675) <= not b or a;
    layer4_outputs(6676) <= '1';
    layer4_outputs(6677) <= '0';
    layer4_outputs(6678) <= not a;
    layer4_outputs(6679) <= '0';
    layer4_outputs(6680) <= not b;
    layer4_outputs(6681) <= not b;
    layer4_outputs(6682) <= not (a or b);
    layer4_outputs(6683) <= b;
    layer4_outputs(6684) <= not (a and b);
    layer4_outputs(6685) <= b and not a;
    layer4_outputs(6686) <= b;
    layer4_outputs(6687) <= '1';
    layer4_outputs(6688) <= '1';
    layer4_outputs(6689) <= not b or a;
    layer4_outputs(6690) <= b;
    layer4_outputs(6691) <= not a;
    layer4_outputs(6692) <= not (a and b);
    layer4_outputs(6693) <= not (a and b);
    layer4_outputs(6694) <= not (a or b);
    layer4_outputs(6695) <= not (a and b);
    layer4_outputs(6696) <= a;
    layer4_outputs(6697) <= not a or b;
    layer4_outputs(6698) <= a and b;
    layer4_outputs(6699) <= a and b;
    layer4_outputs(6700) <= b and not a;
    layer4_outputs(6701) <= not b;
    layer4_outputs(6702) <= not a or b;
    layer4_outputs(6703) <= a;
    layer4_outputs(6704) <= not a or b;
    layer4_outputs(6705) <= b and not a;
    layer4_outputs(6706) <= a;
    layer4_outputs(6707) <= a and not b;
    layer4_outputs(6708) <= not a;
    layer4_outputs(6709) <= not a or b;
    layer4_outputs(6710) <= a and not b;
    layer4_outputs(6711) <= not a or b;
    layer4_outputs(6712) <= b and not a;
    layer4_outputs(6713) <= a;
    layer4_outputs(6714) <= a and b;
    layer4_outputs(6715) <= not (a or b);
    layer4_outputs(6716) <= a and not b;
    layer4_outputs(6717) <= '0';
    layer4_outputs(6718) <= not b or a;
    layer4_outputs(6719) <= not b;
    layer4_outputs(6720) <= b;
    layer4_outputs(6721) <= not a or b;
    layer4_outputs(6722) <= '0';
    layer4_outputs(6723) <= not (a or b);
    layer4_outputs(6724) <= not (a xor b);
    layer4_outputs(6725) <= not a;
    layer4_outputs(6726) <= not a;
    layer4_outputs(6727) <= not a or b;
    layer4_outputs(6728) <= not b or a;
    layer4_outputs(6729) <= not a or b;
    layer4_outputs(6730) <= not a or b;
    layer4_outputs(6731) <= '1';
    layer4_outputs(6732) <= not b or a;
    layer4_outputs(6733) <= b and not a;
    layer4_outputs(6734) <= a;
    layer4_outputs(6735) <= not a;
    layer4_outputs(6736) <= b and not a;
    layer4_outputs(6737) <= not a;
    layer4_outputs(6738) <= not (a xor b);
    layer4_outputs(6739) <= a and not b;
    layer4_outputs(6740) <= not b or a;
    layer4_outputs(6741) <= not b or a;
    layer4_outputs(6742) <= not b;
    layer4_outputs(6743) <= a and not b;
    layer4_outputs(6744) <= not a or b;
    layer4_outputs(6745) <= '0';
    layer4_outputs(6746) <= not b;
    layer4_outputs(6747) <= not b;
    layer4_outputs(6748) <= not b;
    layer4_outputs(6749) <= a xor b;
    layer4_outputs(6750) <= b;
    layer4_outputs(6751) <= '0';
    layer4_outputs(6752) <= a or b;
    layer4_outputs(6753) <= a;
    layer4_outputs(6754) <= a and b;
    layer4_outputs(6755) <= not (a xor b);
    layer4_outputs(6756) <= not b;
    layer4_outputs(6757) <= a and not b;
    layer4_outputs(6758) <= a and b;
    layer4_outputs(6759) <= a or b;
    layer4_outputs(6760) <= a or b;
    layer4_outputs(6761) <= a and not b;
    layer4_outputs(6762) <= b;
    layer4_outputs(6763) <= a and not b;
    layer4_outputs(6764) <= not (a and b);
    layer4_outputs(6765) <= a and not b;
    layer4_outputs(6766) <= a and b;
    layer4_outputs(6767) <= not a;
    layer4_outputs(6768) <= b;
    layer4_outputs(6769) <= a and not b;
    layer4_outputs(6770) <= not b;
    layer4_outputs(6771) <= b;
    layer4_outputs(6772) <= not (a or b);
    layer4_outputs(6773) <= not a or b;
    layer4_outputs(6774) <= a and b;
    layer4_outputs(6775) <= not (a xor b);
    layer4_outputs(6776) <= not b or a;
    layer4_outputs(6777) <= '0';
    layer4_outputs(6778) <= not (a and b);
    layer4_outputs(6779) <= not b;
    layer4_outputs(6780) <= a or b;
    layer4_outputs(6781) <= not a;
    layer4_outputs(6782) <= b and not a;
    layer4_outputs(6783) <= not (a and b);
    layer4_outputs(6784) <= not (a and b);
    layer4_outputs(6785) <= not a;
    layer4_outputs(6786) <= b;
    layer4_outputs(6787) <= not a;
    layer4_outputs(6788) <= not a;
    layer4_outputs(6789) <= b and not a;
    layer4_outputs(6790) <= b;
    layer4_outputs(6791) <= b and not a;
    layer4_outputs(6792) <= a;
    layer4_outputs(6793) <= a and b;
    layer4_outputs(6794) <= '0';
    layer4_outputs(6795) <= not b;
    layer4_outputs(6796) <= '0';
    layer4_outputs(6797) <= '1';
    layer4_outputs(6798) <= b;
    layer4_outputs(6799) <= not (a and b);
    layer4_outputs(6800) <= '0';
    layer4_outputs(6801) <= a or b;
    layer4_outputs(6802) <= not (a or b);
    layer4_outputs(6803) <= not b or a;
    layer4_outputs(6804) <= a or b;
    layer4_outputs(6805) <= '1';
    layer4_outputs(6806) <= a or b;
    layer4_outputs(6807) <= a and not b;
    layer4_outputs(6808) <= not (a and b);
    layer4_outputs(6809) <= not b;
    layer4_outputs(6810) <= not a;
    layer4_outputs(6811) <= b and not a;
    layer4_outputs(6812) <= a;
    layer4_outputs(6813) <= not b or a;
    layer4_outputs(6814) <= b and not a;
    layer4_outputs(6815) <= a and not b;
    layer4_outputs(6816) <= not (a and b);
    layer4_outputs(6817) <= a and not b;
    layer4_outputs(6818) <= a and b;
    layer4_outputs(6819) <= not a or b;
    layer4_outputs(6820) <= a and b;
    layer4_outputs(6821) <= '1';
    layer4_outputs(6822) <= a xor b;
    layer4_outputs(6823) <= a or b;
    layer4_outputs(6824) <= not a or b;
    layer4_outputs(6825) <= a or b;
    layer4_outputs(6826) <= not (a and b);
    layer4_outputs(6827) <= '0';
    layer4_outputs(6828) <= a;
    layer4_outputs(6829) <= not (a or b);
    layer4_outputs(6830) <= a;
    layer4_outputs(6831) <= a;
    layer4_outputs(6832) <= not b or a;
    layer4_outputs(6833) <= '0';
    layer4_outputs(6834) <= not b;
    layer4_outputs(6835) <= '0';
    layer4_outputs(6836) <= b;
    layer4_outputs(6837) <= a xor b;
    layer4_outputs(6838) <= a or b;
    layer4_outputs(6839) <= not a or b;
    layer4_outputs(6840) <= not b or a;
    layer4_outputs(6841) <= not b;
    layer4_outputs(6842) <= b;
    layer4_outputs(6843) <= a;
    layer4_outputs(6844) <= b;
    layer4_outputs(6845) <= not b or a;
    layer4_outputs(6846) <= not (a or b);
    layer4_outputs(6847) <= not (a xor b);
    layer4_outputs(6848) <= not (a and b);
    layer4_outputs(6849) <= a and not b;
    layer4_outputs(6850) <= a and b;
    layer4_outputs(6851) <= '1';
    layer4_outputs(6852) <= '1';
    layer4_outputs(6853) <= '1';
    layer4_outputs(6854) <= b;
    layer4_outputs(6855) <= '1';
    layer4_outputs(6856) <= not a or b;
    layer4_outputs(6857) <= not (a xor b);
    layer4_outputs(6858) <= a and b;
    layer4_outputs(6859) <= '1';
    layer4_outputs(6860) <= not b;
    layer4_outputs(6861) <= a;
    layer4_outputs(6862) <= b and not a;
    layer4_outputs(6863) <= not b or a;
    layer4_outputs(6864) <= not b or a;
    layer4_outputs(6865) <= not a or b;
    layer4_outputs(6866) <= a or b;
    layer4_outputs(6867) <= a and b;
    layer4_outputs(6868) <= not a or b;
    layer4_outputs(6869) <= a;
    layer4_outputs(6870) <= not (a or b);
    layer4_outputs(6871) <= '1';
    layer4_outputs(6872) <= '0';
    layer4_outputs(6873) <= not (a or b);
    layer4_outputs(6874) <= not b or a;
    layer4_outputs(6875) <= a;
    layer4_outputs(6876) <= a and not b;
    layer4_outputs(6877) <= not b;
    layer4_outputs(6878) <= a xor b;
    layer4_outputs(6879) <= not (a and b);
    layer4_outputs(6880) <= not (a and b);
    layer4_outputs(6881) <= not a;
    layer4_outputs(6882) <= not (a and b);
    layer4_outputs(6883) <= a and b;
    layer4_outputs(6884) <= b;
    layer4_outputs(6885) <= not a;
    layer4_outputs(6886) <= '1';
    layer4_outputs(6887) <= b;
    layer4_outputs(6888) <= not b or a;
    layer4_outputs(6889) <= '0';
    layer4_outputs(6890) <= not b;
    layer4_outputs(6891) <= not a;
    layer4_outputs(6892) <= not a;
    layer4_outputs(6893) <= b and not a;
    layer4_outputs(6894) <= b;
    layer4_outputs(6895) <= not a;
    layer4_outputs(6896) <= not a or b;
    layer4_outputs(6897) <= not b or a;
    layer4_outputs(6898) <= not b or a;
    layer4_outputs(6899) <= not b or a;
    layer4_outputs(6900) <= b and not a;
    layer4_outputs(6901) <= not a or b;
    layer4_outputs(6902) <= not (a or b);
    layer4_outputs(6903) <= '1';
    layer4_outputs(6904) <= a and b;
    layer4_outputs(6905) <= a or b;
    layer4_outputs(6906) <= not b or a;
    layer4_outputs(6907) <= a or b;
    layer4_outputs(6908) <= a and not b;
    layer4_outputs(6909) <= b and not a;
    layer4_outputs(6910) <= not a or b;
    layer4_outputs(6911) <= '1';
    layer4_outputs(6912) <= not b or a;
    layer4_outputs(6913) <= not (a xor b);
    layer4_outputs(6914) <= not b or a;
    layer4_outputs(6915) <= not (a and b);
    layer4_outputs(6916) <= a and b;
    layer4_outputs(6917) <= a and not b;
    layer4_outputs(6918) <= b;
    layer4_outputs(6919) <= not a;
    layer4_outputs(6920) <= not (a and b);
    layer4_outputs(6921) <= a and b;
    layer4_outputs(6922) <= not (a xor b);
    layer4_outputs(6923) <= not (a or b);
    layer4_outputs(6924) <= not b or a;
    layer4_outputs(6925) <= not a;
    layer4_outputs(6926) <= a or b;
    layer4_outputs(6927) <= b and not a;
    layer4_outputs(6928) <= a and not b;
    layer4_outputs(6929) <= a;
    layer4_outputs(6930) <= a and not b;
    layer4_outputs(6931) <= b;
    layer4_outputs(6932) <= '0';
    layer4_outputs(6933) <= a and b;
    layer4_outputs(6934) <= a or b;
    layer4_outputs(6935) <= '0';
    layer4_outputs(6936) <= a or b;
    layer4_outputs(6937) <= a or b;
    layer4_outputs(6938) <= a or b;
    layer4_outputs(6939) <= not b;
    layer4_outputs(6940) <= a;
    layer4_outputs(6941) <= '0';
    layer4_outputs(6942) <= '0';
    layer4_outputs(6943) <= a or b;
    layer4_outputs(6944) <= a and b;
    layer4_outputs(6945) <= a or b;
    layer4_outputs(6946) <= b;
    layer4_outputs(6947) <= not (a or b);
    layer4_outputs(6948) <= b;
    layer4_outputs(6949) <= not (a or b);
    layer4_outputs(6950) <= a and b;
    layer4_outputs(6951) <= not a;
    layer4_outputs(6952) <= a and not b;
    layer4_outputs(6953) <= a or b;
    layer4_outputs(6954) <= a;
    layer4_outputs(6955) <= b and not a;
    layer4_outputs(6956) <= b and not a;
    layer4_outputs(6957) <= a and not b;
    layer4_outputs(6958) <= a and not b;
    layer4_outputs(6959) <= '0';
    layer4_outputs(6960) <= '0';
    layer4_outputs(6961) <= a and b;
    layer4_outputs(6962) <= b;
    layer4_outputs(6963) <= not (a and b);
    layer4_outputs(6964) <= not (a or b);
    layer4_outputs(6965) <= not a or b;
    layer4_outputs(6966) <= not (a and b);
    layer4_outputs(6967) <= not a;
    layer4_outputs(6968) <= a xor b;
    layer4_outputs(6969) <= '0';
    layer4_outputs(6970) <= not (a or b);
    layer4_outputs(6971) <= a;
    layer4_outputs(6972) <= not (a xor b);
    layer4_outputs(6973) <= b;
    layer4_outputs(6974) <= '1';
    layer4_outputs(6975) <= not a or b;
    layer4_outputs(6976) <= a xor b;
    layer4_outputs(6977) <= '1';
    layer4_outputs(6978) <= not (a and b);
    layer4_outputs(6979) <= b and not a;
    layer4_outputs(6980) <= not (a and b);
    layer4_outputs(6981) <= not (a or b);
    layer4_outputs(6982) <= b and not a;
    layer4_outputs(6983) <= b and not a;
    layer4_outputs(6984) <= not a or b;
    layer4_outputs(6985) <= not (a or b);
    layer4_outputs(6986) <= not a;
    layer4_outputs(6987) <= a and b;
    layer4_outputs(6988) <= not a or b;
    layer4_outputs(6989) <= b and not a;
    layer4_outputs(6990) <= b and not a;
    layer4_outputs(6991) <= not (a or b);
    layer4_outputs(6992) <= not a or b;
    layer4_outputs(6993) <= a and b;
    layer4_outputs(6994) <= '1';
    layer4_outputs(6995) <= a and b;
    layer4_outputs(6996) <= b;
    layer4_outputs(6997) <= '1';
    layer4_outputs(6998) <= not b or a;
    layer4_outputs(6999) <= not a;
    layer4_outputs(7000) <= not (a or b);
    layer4_outputs(7001) <= not a;
    layer4_outputs(7002) <= not b or a;
    layer4_outputs(7003) <= a;
    layer4_outputs(7004) <= a;
    layer4_outputs(7005) <= a and not b;
    layer4_outputs(7006) <= b;
    layer4_outputs(7007) <= not b or a;
    layer4_outputs(7008) <= not (a or b);
    layer4_outputs(7009) <= a and b;
    layer4_outputs(7010) <= not (a or b);
    layer4_outputs(7011) <= a;
    layer4_outputs(7012) <= not (a or b);
    layer4_outputs(7013) <= not a;
    layer4_outputs(7014) <= '0';
    layer4_outputs(7015) <= not (a and b);
    layer4_outputs(7016) <= not a or b;
    layer4_outputs(7017) <= not a;
    layer4_outputs(7018) <= '0';
    layer4_outputs(7019) <= not a;
    layer4_outputs(7020) <= not b;
    layer4_outputs(7021) <= not b or a;
    layer4_outputs(7022) <= a xor b;
    layer4_outputs(7023) <= a and not b;
    layer4_outputs(7024) <= a;
    layer4_outputs(7025) <= not b or a;
    layer4_outputs(7026) <= not (a xor b);
    layer4_outputs(7027) <= b;
    layer4_outputs(7028) <= a and b;
    layer4_outputs(7029) <= not b;
    layer4_outputs(7030) <= not b or a;
    layer4_outputs(7031) <= not b or a;
    layer4_outputs(7032) <= not b;
    layer4_outputs(7033) <= not b or a;
    layer4_outputs(7034) <= not a or b;
    layer4_outputs(7035) <= not b;
    layer4_outputs(7036) <= '1';
    layer4_outputs(7037) <= a and b;
    layer4_outputs(7038) <= '1';
    layer4_outputs(7039) <= '0';
    layer4_outputs(7040) <= not a;
    layer4_outputs(7041) <= a xor b;
    layer4_outputs(7042) <= b;
    layer4_outputs(7043) <= '0';
    layer4_outputs(7044) <= '0';
    layer4_outputs(7045) <= b;
    layer4_outputs(7046) <= not a;
    layer4_outputs(7047) <= b;
    layer4_outputs(7048) <= not (a or b);
    layer4_outputs(7049) <= not (a and b);
    layer4_outputs(7050) <= a and b;
    layer4_outputs(7051) <= not a;
    layer4_outputs(7052) <= b;
    layer4_outputs(7053) <= a or b;
    layer4_outputs(7054) <= a;
    layer4_outputs(7055) <= not (a or b);
    layer4_outputs(7056) <= not b or a;
    layer4_outputs(7057) <= a or b;
    layer4_outputs(7058) <= a and not b;
    layer4_outputs(7059) <= not a or b;
    layer4_outputs(7060) <= a or b;
    layer4_outputs(7061) <= '1';
    layer4_outputs(7062) <= b;
    layer4_outputs(7063) <= a and not b;
    layer4_outputs(7064) <= b;
    layer4_outputs(7065) <= b and not a;
    layer4_outputs(7066) <= a and b;
    layer4_outputs(7067) <= b;
    layer4_outputs(7068) <= not b;
    layer4_outputs(7069) <= a or b;
    layer4_outputs(7070) <= not (a or b);
    layer4_outputs(7071) <= a and b;
    layer4_outputs(7072) <= '1';
    layer4_outputs(7073) <= not b or a;
    layer4_outputs(7074) <= '0';
    layer4_outputs(7075) <= not a or b;
    layer4_outputs(7076) <= a and b;
    layer4_outputs(7077) <= a and not b;
    layer4_outputs(7078) <= not (a or b);
    layer4_outputs(7079) <= a or b;
    layer4_outputs(7080) <= a or b;
    layer4_outputs(7081) <= b;
    layer4_outputs(7082) <= not a;
    layer4_outputs(7083) <= a and not b;
    layer4_outputs(7084) <= a xor b;
    layer4_outputs(7085) <= not a;
    layer4_outputs(7086) <= a or b;
    layer4_outputs(7087) <= '1';
    layer4_outputs(7088) <= not b;
    layer4_outputs(7089) <= not (a and b);
    layer4_outputs(7090) <= b and not a;
    layer4_outputs(7091) <= not (a and b);
    layer4_outputs(7092) <= a;
    layer4_outputs(7093) <= b;
    layer4_outputs(7094) <= not b;
    layer4_outputs(7095) <= b and not a;
    layer4_outputs(7096) <= not a or b;
    layer4_outputs(7097) <= a or b;
    layer4_outputs(7098) <= not (a and b);
    layer4_outputs(7099) <= not b;
    layer4_outputs(7100) <= a or b;
    layer4_outputs(7101) <= not (a or b);
    layer4_outputs(7102) <= not (a xor b);
    layer4_outputs(7103) <= b;
    layer4_outputs(7104) <= '1';
    layer4_outputs(7105) <= a or b;
    layer4_outputs(7106) <= not (a and b);
    layer4_outputs(7107) <= a or b;
    layer4_outputs(7108) <= a and b;
    layer4_outputs(7109) <= a;
    layer4_outputs(7110) <= not a;
    layer4_outputs(7111) <= not a or b;
    layer4_outputs(7112) <= not a;
    layer4_outputs(7113) <= not b;
    layer4_outputs(7114) <= not a or b;
    layer4_outputs(7115) <= a or b;
    layer4_outputs(7116) <= a or b;
    layer4_outputs(7117) <= b and not a;
    layer4_outputs(7118) <= a and b;
    layer4_outputs(7119) <= not a;
    layer4_outputs(7120) <= not (a xor b);
    layer4_outputs(7121) <= not a or b;
    layer4_outputs(7122) <= not a or b;
    layer4_outputs(7123) <= a or b;
    layer4_outputs(7124) <= a;
    layer4_outputs(7125) <= b and not a;
    layer4_outputs(7126) <= a;
    layer4_outputs(7127) <= not a;
    layer4_outputs(7128) <= not (a and b);
    layer4_outputs(7129) <= not a;
    layer4_outputs(7130) <= not (a or b);
    layer4_outputs(7131) <= a;
    layer4_outputs(7132) <= '0';
    layer4_outputs(7133) <= not (a and b);
    layer4_outputs(7134) <= a;
    layer4_outputs(7135) <= not (a or b);
    layer4_outputs(7136) <= not b or a;
    layer4_outputs(7137) <= '0';
    layer4_outputs(7138) <= b and not a;
    layer4_outputs(7139) <= b and not a;
    layer4_outputs(7140) <= not a or b;
    layer4_outputs(7141) <= not a or b;
    layer4_outputs(7142) <= a and not b;
    layer4_outputs(7143) <= b and not a;
    layer4_outputs(7144) <= a and b;
    layer4_outputs(7145) <= '0';
    layer4_outputs(7146) <= not a;
    layer4_outputs(7147) <= not (a or b);
    layer4_outputs(7148) <= not b or a;
    layer4_outputs(7149) <= not a or b;
    layer4_outputs(7150) <= a xor b;
    layer4_outputs(7151) <= not a;
    layer4_outputs(7152) <= not a or b;
    layer4_outputs(7153) <= a and not b;
    layer4_outputs(7154) <= not a;
    layer4_outputs(7155) <= a and not b;
    layer4_outputs(7156) <= not b;
    layer4_outputs(7157) <= a;
    layer4_outputs(7158) <= not a;
    layer4_outputs(7159) <= '0';
    layer4_outputs(7160) <= a or b;
    layer4_outputs(7161) <= b and not a;
    layer4_outputs(7162) <= a and b;
    layer4_outputs(7163) <= b;
    layer4_outputs(7164) <= not a;
    layer4_outputs(7165) <= not a;
    layer4_outputs(7166) <= not (a and b);
    layer4_outputs(7167) <= not (a and b);
    layer4_outputs(7168) <= not b or a;
    layer4_outputs(7169) <= a or b;
    layer4_outputs(7170) <= b;
    layer4_outputs(7171) <= a;
    layer4_outputs(7172) <= a;
    layer4_outputs(7173) <= not b;
    layer4_outputs(7174) <= a xor b;
    layer4_outputs(7175) <= not a;
    layer4_outputs(7176) <= a and b;
    layer4_outputs(7177) <= b;
    layer4_outputs(7178) <= not a;
    layer4_outputs(7179) <= not a or b;
    layer4_outputs(7180) <= not a or b;
    layer4_outputs(7181) <= a or b;
    layer4_outputs(7182) <= b and not a;
    layer4_outputs(7183) <= b and not a;
    layer4_outputs(7184) <= a or b;
    layer4_outputs(7185) <= a and b;
    layer4_outputs(7186) <= not (a and b);
    layer4_outputs(7187) <= b;
    layer4_outputs(7188) <= a;
    layer4_outputs(7189) <= b and not a;
    layer4_outputs(7190) <= '0';
    layer4_outputs(7191) <= b and not a;
    layer4_outputs(7192) <= not (a and b);
    layer4_outputs(7193) <= b;
    layer4_outputs(7194) <= not a or b;
    layer4_outputs(7195) <= a and not b;
    layer4_outputs(7196) <= not b;
    layer4_outputs(7197) <= '1';
    layer4_outputs(7198) <= not b or a;
    layer4_outputs(7199) <= '1';
    layer4_outputs(7200) <= not (a and b);
    layer4_outputs(7201) <= '0';
    layer4_outputs(7202) <= a;
    layer4_outputs(7203) <= not a or b;
    layer4_outputs(7204) <= '0';
    layer4_outputs(7205) <= not b;
    layer4_outputs(7206) <= b and not a;
    layer4_outputs(7207) <= b;
    layer4_outputs(7208) <= not a;
    layer4_outputs(7209) <= not b;
    layer4_outputs(7210) <= a and not b;
    layer4_outputs(7211) <= '1';
    layer4_outputs(7212) <= not b or a;
    layer4_outputs(7213) <= b;
    layer4_outputs(7214) <= b;
    layer4_outputs(7215) <= a;
    layer4_outputs(7216) <= not b or a;
    layer4_outputs(7217) <= a;
    layer4_outputs(7218) <= a and b;
    layer4_outputs(7219) <= not b or a;
    layer4_outputs(7220) <= not a;
    layer4_outputs(7221) <= not (a and b);
    layer4_outputs(7222) <= b;
    layer4_outputs(7223) <= not b;
    layer4_outputs(7224) <= a;
    layer4_outputs(7225) <= not (a xor b);
    layer4_outputs(7226) <= a and b;
    layer4_outputs(7227) <= a and not b;
    layer4_outputs(7228) <= not (a xor b);
    layer4_outputs(7229) <= '1';
    layer4_outputs(7230) <= not b;
    layer4_outputs(7231) <= '1';
    layer4_outputs(7232) <= a and b;
    layer4_outputs(7233) <= not a or b;
    layer4_outputs(7234) <= '0';
    layer4_outputs(7235) <= not a or b;
    layer4_outputs(7236) <= a and not b;
    layer4_outputs(7237) <= a and not b;
    layer4_outputs(7238) <= a;
    layer4_outputs(7239) <= a or b;
    layer4_outputs(7240) <= not b;
    layer4_outputs(7241) <= b;
    layer4_outputs(7242) <= a or b;
    layer4_outputs(7243) <= a or b;
    layer4_outputs(7244) <= not a;
    layer4_outputs(7245) <= not a;
    layer4_outputs(7246) <= a or b;
    layer4_outputs(7247) <= not (a xor b);
    layer4_outputs(7248) <= a or b;
    layer4_outputs(7249) <= a;
    layer4_outputs(7250) <= not b;
    layer4_outputs(7251) <= '1';
    layer4_outputs(7252) <= not a or b;
    layer4_outputs(7253) <= not (a and b);
    layer4_outputs(7254) <= not (a or b);
    layer4_outputs(7255) <= a or b;
    layer4_outputs(7256) <= a and b;
    layer4_outputs(7257) <= a or b;
    layer4_outputs(7258) <= a;
    layer4_outputs(7259) <= not a;
    layer4_outputs(7260) <= not a or b;
    layer4_outputs(7261) <= a and b;
    layer4_outputs(7262) <= a and not b;
    layer4_outputs(7263) <= a xor b;
    layer4_outputs(7264) <= not a;
    layer4_outputs(7265) <= not b or a;
    layer4_outputs(7266) <= a and b;
    layer4_outputs(7267) <= not (a and b);
    layer4_outputs(7268) <= not (a or b);
    layer4_outputs(7269) <= not a;
    layer4_outputs(7270) <= not (a or b);
    layer4_outputs(7271) <= not (a and b);
    layer4_outputs(7272) <= a or b;
    layer4_outputs(7273) <= a or b;
    layer4_outputs(7274) <= a and not b;
    layer4_outputs(7275) <= not b;
    layer4_outputs(7276) <= a and not b;
    layer4_outputs(7277) <= not (a xor b);
    layer4_outputs(7278) <= a or b;
    layer4_outputs(7279) <= not a or b;
    layer4_outputs(7280) <= not (a xor b);
    layer4_outputs(7281) <= not b or a;
    layer4_outputs(7282) <= not b;
    layer4_outputs(7283) <= a and not b;
    layer4_outputs(7284) <= not b;
    layer4_outputs(7285) <= not b;
    layer4_outputs(7286) <= a and not b;
    layer4_outputs(7287) <= not b;
    layer4_outputs(7288) <= a and not b;
    layer4_outputs(7289) <= a and b;
    layer4_outputs(7290) <= a and not b;
    layer4_outputs(7291) <= a;
    layer4_outputs(7292) <= b;
    layer4_outputs(7293) <= b and not a;
    layer4_outputs(7294) <= not a;
    layer4_outputs(7295) <= not b;
    layer4_outputs(7296) <= not a or b;
    layer4_outputs(7297) <= b;
    layer4_outputs(7298) <= not b;
    layer4_outputs(7299) <= a;
    layer4_outputs(7300) <= not b;
    layer4_outputs(7301) <= b;
    layer4_outputs(7302) <= not a;
    layer4_outputs(7303) <= not (a and b);
    layer4_outputs(7304) <= b;
    layer4_outputs(7305) <= b;
    layer4_outputs(7306) <= a and not b;
    layer4_outputs(7307) <= b and not a;
    layer4_outputs(7308) <= '1';
    layer4_outputs(7309) <= not (a and b);
    layer4_outputs(7310) <= '1';
    layer4_outputs(7311) <= not b or a;
    layer4_outputs(7312) <= a and not b;
    layer4_outputs(7313) <= not b or a;
    layer4_outputs(7314) <= not a;
    layer4_outputs(7315) <= a and b;
    layer4_outputs(7316) <= b and not a;
    layer4_outputs(7317) <= '0';
    layer4_outputs(7318) <= not a;
    layer4_outputs(7319) <= not (a and b);
    layer4_outputs(7320) <= not a;
    layer4_outputs(7321) <= a and not b;
    layer4_outputs(7322) <= not (a or b);
    layer4_outputs(7323) <= a and b;
    layer4_outputs(7324) <= b;
    layer4_outputs(7325) <= a and not b;
    layer4_outputs(7326) <= b;
    layer4_outputs(7327) <= not (a and b);
    layer4_outputs(7328) <= b;
    layer4_outputs(7329) <= a or b;
    layer4_outputs(7330) <= a or b;
    layer4_outputs(7331) <= not b;
    layer4_outputs(7332) <= a xor b;
    layer4_outputs(7333) <= not b or a;
    layer4_outputs(7334) <= not b;
    layer4_outputs(7335) <= a or b;
    layer4_outputs(7336) <= a;
    layer4_outputs(7337) <= a or b;
    layer4_outputs(7338) <= b;
    layer4_outputs(7339) <= b and not a;
    layer4_outputs(7340) <= not b or a;
    layer4_outputs(7341) <= not (a and b);
    layer4_outputs(7342) <= b;
    layer4_outputs(7343) <= '0';
    layer4_outputs(7344) <= b and not a;
    layer4_outputs(7345) <= a or b;
    layer4_outputs(7346) <= b and not a;
    layer4_outputs(7347) <= not a;
    layer4_outputs(7348) <= a and not b;
    layer4_outputs(7349) <= not (a and b);
    layer4_outputs(7350) <= a and b;
    layer4_outputs(7351) <= not b or a;
    layer4_outputs(7352) <= not (a and b);
    layer4_outputs(7353) <= b and not a;
    layer4_outputs(7354) <= not (a xor b);
    layer4_outputs(7355) <= '0';
    layer4_outputs(7356) <= b;
    layer4_outputs(7357) <= a and not b;
    layer4_outputs(7358) <= '0';
    layer4_outputs(7359) <= not b or a;
    layer4_outputs(7360) <= a or b;
    layer4_outputs(7361) <= not a;
    layer4_outputs(7362) <= a and b;
    layer4_outputs(7363) <= not (a and b);
    layer4_outputs(7364) <= a and not b;
    layer4_outputs(7365) <= a xor b;
    layer4_outputs(7366) <= not (a and b);
    layer4_outputs(7367) <= '0';
    layer4_outputs(7368) <= not (a or b);
    layer4_outputs(7369) <= not b;
    layer4_outputs(7370) <= not b;
    layer4_outputs(7371) <= not b or a;
    layer4_outputs(7372) <= not a or b;
    layer4_outputs(7373) <= not b or a;
    layer4_outputs(7374) <= a or b;
    layer4_outputs(7375) <= a;
    layer4_outputs(7376) <= '1';
    layer4_outputs(7377) <= not (a or b);
    layer4_outputs(7378) <= a and not b;
    layer4_outputs(7379) <= not a or b;
    layer4_outputs(7380) <= '1';
    layer4_outputs(7381) <= a or b;
    layer4_outputs(7382) <= not a;
    layer4_outputs(7383) <= not (a and b);
    layer4_outputs(7384) <= not b or a;
    layer4_outputs(7385) <= a and b;
    layer4_outputs(7386) <= a and not b;
    layer4_outputs(7387) <= not a or b;
    layer4_outputs(7388) <= '1';
    layer4_outputs(7389) <= b;
    layer4_outputs(7390) <= a or b;
    layer4_outputs(7391) <= not a;
    layer4_outputs(7392) <= not (a or b);
    layer4_outputs(7393) <= a and b;
    layer4_outputs(7394) <= b and not a;
    layer4_outputs(7395) <= not (a and b);
    layer4_outputs(7396) <= a xor b;
    layer4_outputs(7397) <= not b or a;
    layer4_outputs(7398) <= not (a and b);
    layer4_outputs(7399) <= not (a or b);
    layer4_outputs(7400) <= not (a or b);
    layer4_outputs(7401) <= b and not a;
    layer4_outputs(7402) <= a;
    layer4_outputs(7403) <= not (a and b);
    layer4_outputs(7404) <= a and not b;
    layer4_outputs(7405) <= '0';
    layer4_outputs(7406) <= b and not a;
    layer4_outputs(7407) <= b;
    layer4_outputs(7408) <= a xor b;
    layer4_outputs(7409) <= '1';
    layer4_outputs(7410) <= '0';
    layer4_outputs(7411) <= b;
    layer4_outputs(7412) <= not (a xor b);
    layer4_outputs(7413) <= not a or b;
    layer4_outputs(7414) <= not b or a;
    layer4_outputs(7415) <= a;
    layer4_outputs(7416) <= '1';
    layer4_outputs(7417) <= a;
    layer4_outputs(7418) <= '0';
    layer4_outputs(7419) <= not b;
    layer4_outputs(7420) <= a and b;
    layer4_outputs(7421) <= not b or a;
    layer4_outputs(7422) <= '1';
    layer4_outputs(7423) <= not b;
    layer4_outputs(7424) <= '1';
    layer4_outputs(7425) <= a and not b;
    layer4_outputs(7426) <= not (a and b);
    layer4_outputs(7427) <= not b or a;
    layer4_outputs(7428) <= b;
    layer4_outputs(7429) <= b and not a;
    layer4_outputs(7430) <= not (a or b);
    layer4_outputs(7431) <= a and b;
    layer4_outputs(7432) <= '0';
    layer4_outputs(7433) <= a;
    layer4_outputs(7434) <= a or b;
    layer4_outputs(7435) <= not (a and b);
    layer4_outputs(7436) <= b and not a;
    layer4_outputs(7437) <= not a;
    layer4_outputs(7438) <= not a or b;
    layer4_outputs(7439) <= b and not a;
    layer4_outputs(7440) <= a xor b;
    layer4_outputs(7441) <= not (a xor b);
    layer4_outputs(7442) <= a and b;
    layer4_outputs(7443) <= not a or b;
    layer4_outputs(7444) <= a or b;
    layer4_outputs(7445) <= a and not b;
    layer4_outputs(7446) <= not (a or b);
    layer4_outputs(7447) <= not a;
    layer4_outputs(7448) <= not a or b;
    layer4_outputs(7449) <= '1';
    layer4_outputs(7450) <= '0';
    layer4_outputs(7451) <= b;
    layer4_outputs(7452) <= not b;
    layer4_outputs(7453) <= b;
    layer4_outputs(7454) <= a or b;
    layer4_outputs(7455) <= not (a xor b);
    layer4_outputs(7456) <= b and not a;
    layer4_outputs(7457) <= a xor b;
    layer4_outputs(7458) <= a and not b;
    layer4_outputs(7459) <= a;
    layer4_outputs(7460) <= '0';
    layer4_outputs(7461) <= not (a or b);
    layer4_outputs(7462) <= not (a or b);
    layer4_outputs(7463) <= b and not a;
    layer4_outputs(7464) <= not (a and b);
    layer4_outputs(7465) <= not b;
    layer4_outputs(7466) <= b;
    layer4_outputs(7467) <= not a or b;
    layer4_outputs(7468) <= '1';
    layer4_outputs(7469) <= not a;
    layer4_outputs(7470) <= not (a or b);
    layer4_outputs(7471) <= '0';
    layer4_outputs(7472) <= not (a and b);
    layer4_outputs(7473) <= not b or a;
    layer4_outputs(7474) <= not (a or b);
    layer4_outputs(7475) <= a or b;
    layer4_outputs(7476) <= not (a xor b);
    layer4_outputs(7477) <= a or b;
    layer4_outputs(7478) <= not b or a;
    layer4_outputs(7479) <= not a;
    layer4_outputs(7480) <= not (a and b);
    layer4_outputs(7481) <= b;
    layer4_outputs(7482) <= b and not a;
    layer4_outputs(7483) <= a and not b;
    layer4_outputs(7484) <= not a;
    layer4_outputs(7485) <= '0';
    layer4_outputs(7486) <= '1';
    layer4_outputs(7487) <= b;
    layer4_outputs(7488) <= a or b;
    layer4_outputs(7489) <= a and b;
    layer4_outputs(7490) <= not a;
    layer4_outputs(7491) <= not b;
    layer4_outputs(7492) <= a or b;
    layer4_outputs(7493) <= a and not b;
    layer4_outputs(7494) <= not a;
    layer4_outputs(7495) <= b;
    layer4_outputs(7496) <= not b;
    layer4_outputs(7497) <= not a or b;
    layer4_outputs(7498) <= '1';
    layer4_outputs(7499) <= not (a or b);
    layer4_outputs(7500) <= not a or b;
    layer4_outputs(7501) <= a and not b;
    layer4_outputs(7502) <= a or b;
    layer4_outputs(7503) <= a and b;
    layer4_outputs(7504) <= a;
    layer4_outputs(7505) <= '0';
    layer4_outputs(7506) <= b;
    layer4_outputs(7507) <= a and b;
    layer4_outputs(7508) <= a or b;
    layer4_outputs(7509) <= b;
    layer4_outputs(7510) <= a and not b;
    layer4_outputs(7511) <= a or b;
    layer4_outputs(7512) <= not (a and b);
    layer4_outputs(7513) <= b;
    layer4_outputs(7514) <= not (a xor b);
    layer4_outputs(7515) <= not a;
    layer4_outputs(7516) <= not b;
    layer4_outputs(7517) <= '0';
    layer4_outputs(7518) <= a and not b;
    layer4_outputs(7519) <= a and not b;
    layer4_outputs(7520) <= b and not a;
    layer4_outputs(7521) <= not b;
    layer4_outputs(7522) <= not a or b;
    layer4_outputs(7523) <= b;
    layer4_outputs(7524) <= not (a and b);
    layer4_outputs(7525) <= b;
    layer4_outputs(7526) <= b;
    layer4_outputs(7527) <= a and not b;
    layer4_outputs(7528) <= '0';
    layer4_outputs(7529) <= b;
    layer4_outputs(7530) <= a and b;
    layer4_outputs(7531) <= not a or b;
    layer4_outputs(7532) <= b;
    layer4_outputs(7533) <= not b or a;
    layer4_outputs(7534) <= not (a xor b);
    layer4_outputs(7535) <= a and b;
    layer4_outputs(7536) <= a and b;
    layer4_outputs(7537) <= '1';
    layer4_outputs(7538) <= not (a or b);
    layer4_outputs(7539) <= a and not b;
    layer4_outputs(7540) <= a;
    layer4_outputs(7541) <= b and not a;
    layer4_outputs(7542) <= not (a or b);
    layer4_outputs(7543) <= not (a and b);
    layer4_outputs(7544) <= not a;
    layer4_outputs(7545) <= a and b;
    layer4_outputs(7546) <= b;
    layer4_outputs(7547) <= not a;
    layer4_outputs(7548) <= '1';
    layer4_outputs(7549) <= a or b;
    layer4_outputs(7550) <= b;
    layer4_outputs(7551) <= b;
    layer4_outputs(7552) <= b;
    layer4_outputs(7553) <= '0';
    layer4_outputs(7554) <= a and not b;
    layer4_outputs(7555) <= a or b;
    layer4_outputs(7556) <= a or b;
    layer4_outputs(7557) <= not a;
    layer4_outputs(7558) <= not a;
    layer4_outputs(7559) <= '0';
    layer4_outputs(7560) <= '0';
    layer4_outputs(7561) <= not (a or b);
    layer4_outputs(7562) <= a and b;
    layer4_outputs(7563) <= a xor b;
    layer4_outputs(7564) <= b and not a;
    layer4_outputs(7565) <= a and not b;
    layer4_outputs(7566) <= a and b;
    layer4_outputs(7567) <= a;
    layer4_outputs(7568) <= '0';
    layer4_outputs(7569) <= a;
    layer4_outputs(7570) <= not (a or b);
    layer4_outputs(7571) <= a;
    layer4_outputs(7572) <= not b or a;
    layer4_outputs(7573) <= b and not a;
    layer4_outputs(7574) <= not (a and b);
    layer4_outputs(7575) <= not b;
    layer4_outputs(7576) <= not b;
    layer4_outputs(7577) <= not a or b;
    layer4_outputs(7578) <= a and not b;
    layer4_outputs(7579) <= a or b;
    layer4_outputs(7580) <= a or b;
    layer4_outputs(7581) <= a;
    layer4_outputs(7582) <= '0';
    layer4_outputs(7583) <= b;
    layer4_outputs(7584) <= not a or b;
    layer4_outputs(7585) <= not a;
    layer4_outputs(7586) <= not a;
    layer4_outputs(7587) <= not (a and b);
    layer4_outputs(7588) <= a xor b;
    layer4_outputs(7589) <= not (a and b);
    layer4_outputs(7590) <= not a;
    layer4_outputs(7591) <= b;
    layer4_outputs(7592) <= a or b;
    layer4_outputs(7593) <= not (a or b);
    layer4_outputs(7594) <= not a;
    layer4_outputs(7595) <= not b or a;
    layer4_outputs(7596) <= '0';
    layer4_outputs(7597) <= not b;
    layer4_outputs(7598) <= a and b;
    layer4_outputs(7599) <= not (a and b);
    layer4_outputs(7600) <= b;
    layer4_outputs(7601) <= b and not a;
    layer4_outputs(7602) <= a and not b;
    layer4_outputs(7603) <= not a;
    layer4_outputs(7604) <= b;
    layer4_outputs(7605) <= a and not b;
    layer4_outputs(7606) <= not b;
    layer4_outputs(7607) <= not a or b;
    layer4_outputs(7608) <= '1';
    layer4_outputs(7609) <= not a or b;
    layer4_outputs(7610) <= not b;
    layer4_outputs(7611) <= b;
    layer4_outputs(7612) <= not b or a;
    layer4_outputs(7613) <= a or b;
    layer4_outputs(7614) <= a or b;
    layer4_outputs(7615) <= a or b;
    layer4_outputs(7616) <= not b;
    layer4_outputs(7617) <= not b;
    layer4_outputs(7618) <= not a or b;
    layer4_outputs(7619) <= not (a or b);
    layer4_outputs(7620) <= a;
    layer4_outputs(7621) <= b and not a;
    layer4_outputs(7622) <= a or b;
    layer4_outputs(7623) <= a and not b;
    layer4_outputs(7624) <= '0';
    layer4_outputs(7625) <= '0';
    layer4_outputs(7626) <= not a or b;
    layer4_outputs(7627) <= not (a and b);
    layer4_outputs(7628) <= a;
    layer4_outputs(7629) <= a;
    layer4_outputs(7630) <= not b or a;
    layer4_outputs(7631) <= b and not a;
    layer4_outputs(7632) <= a or b;
    layer4_outputs(7633) <= a and not b;
    layer4_outputs(7634) <= '1';
    layer4_outputs(7635) <= b and not a;
    layer4_outputs(7636) <= not b;
    layer4_outputs(7637) <= not a;
    layer4_outputs(7638) <= a or b;
    layer4_outputs(7639) <= not a or b;
    layer4_outputs(7640) <= not b;
    layer4_outputs(7641) <= not (a or b);
    layer4_outputs(7642) <= '1';
    layer4_outputs(7643) <= a or b;
    layer4_outputs(7644) <= a and not b;
    layer4_outputs(7645) <= not a or b;
    layer4_outputs(7646) <= a xor b;
    layer4_outputs(7647) <= not (a or b);
    layer4_outputs(7648) <= not b or a;
    layer4_outputs(7649) <= a or b;
    layer4_outputs(7650) <= not b;
    layer4_outputs(7651) <= b;
    layer4_outputs(7652) <= b and not a;
    layer4_outputs(7653) <= a;
    layer4_outputs(7654) <= b;
    layer4_outputs(7655) <= a and not b;
    layer4_outputs(7656) <= a;
    layer4_outputs(7657) <= not a or b;
    layer4_outputs(7658) <= a and b;
    layer4_outputs(7659) <= a and b;
    layer4_outputs(7660) <= '0';
    layer4_outputs(7661) <= not a;
    layer4_outputs(7662) <= a and not b;
    layer4_outputs(7663) <= b;
    layer4_outputs(7664) <= not a;
    layer4_outputs(7665) <= a;
    layer4_outputs(7666) <= a or b;
    layer4_outputs(7667) <= not b or a;
    layer4_outputs(7668) <= a and b;
    layer4_outputs(7669) <= a;
    layer4_outputs(7670) <= not b;
    layer4_outputs(7671) <= not (a and b);
    layer4_outputs(7672) <= a and b;
    layer4_outputs(7673) <= not a;
    layer4_outputs(7674) <= '1';
    layer4_outputs(7675) <= b and not a;
    layer4_outputs(7676) <= a or b;
    layer4_outputs(7677) <= not (a xor b);
    layer4_outputs(7678) <= a and b;
    layer4_outputs(7679) <= a and b;
    layer5_outputs(0) <= not b or a;
    layer5_outputs(1) <= not b;
    layer5_outputs(2) <= not a or b;
    layer5_outputs(3) <= not (a and b);
    layer5_outputs(4) <= a and not b;
    layer5_outputs(5) <= b and not a;
    layer5_outputs(6) <= not (a and b);
    layer5_outputs(7) <= b and not a;
    layer5_outputs(8) <= a and not b;
    layer5_outputs(9) <= not a or b;
    layer5_outputs(10) <= a or b;
    layer5_outputs(11) <= not (a and b);
    layer5_outputs(12) <= b and not a;
    layer5_outputs(13) <= a or b;
    layer5_outputs(14) <= b;
    layer5_outputs(15) <= b and not a;
    layer5_outputs(16) <= not a;
    layer5_outputs(17) <= not a or b;
    layer5_outputs(18) <= a and not b;
    layer5_outputs(19) <= a and b;
    layer5_outputs(20) <= a or b;
    layer5_outputs(21) <= a and b;
    layer5_outputs(22) <= a xor b;
    layer5_outputs(23) <= not (a xor b);
    layer5_outputs(24) <= a xor b;
    layer5_outputs(25) <= not b;
    layer5_outputs(26) <= not a or b;
    layer5_outputs(27) <= not (a or b);
    layer5_outputs(28) <= not a;
    layer5_outputs(29) <= not a;
    layer5_outputs(30) <= a or b;
    layer5_outputs(31) <= b and not a;
    layer5_outputs(32) <= b and not a;
    layer5_outputs(33) <= b and not a;
    layer5_outputs(34) <= a;
    layer5_outputs(35) <= not b or a;
    layer5_outputs(36) <= not b or a;
    layer5_outputs(37) <= a or b;
    layer5_outputs(38) <= not a;
    layer5_outputs(39) <= not b or a;
    layer5_outputs(40) <= not b;
    layer5_outputs(41) <= b;
    layer5_outputs(42) <= a and b;
    layer5_outputs(43) <= not b;
    layer5_outputs(44) <= b;
    layer5_outputs(45) <= not b;
    layer5_outputs(46) <= not a;
    layer5_outputs(47) <= b and not a;
    layer5_outputs(48) <= not (a and b);
    layer5_outputs(49) <= a or b;
    layer5_outputs(50) <= not (a and b);
    layer5_outputs(51) <= a or b;
    layer5_outputs(52) <= not b;
    layer5_outputs(53) <= '0';
    layer5_outputs(54) <= not a;
    layer5_outputs(55) <= a or b;
    layer5_outputs(56) <= not (a xor b);
    layer5_outputs(57) <= a;
    layer5_outputs(58) <= b and not a;
    layer5_outputs(59) <= b;
    layer5_outputs(60) <= b;
    layer5_outputs(61) <= '1';
    layer5_outputs(62) <= b;
    layer5_outputs(63) <= b;
    layer5_outputs(64) <= b;
    layer5_outputs(65) <= not a or b;
    layer5_outputs(66) <= not b;
    layer5_outputs(67) <= not (a or b);
    layer5_outputs(68) <= not a;
    layer5_outputs(69) <= a or b;
    layer5_outputs(70) <= not (a and b);
    layer5_outputs(71) <= b;
    layer5_outputs(72) <= not a;
    layer5_outputs(73) <= not a or b;
    layer5_outputs(74) <= a and b;
    layer5_outputs(75) <= a and b;
    layer5_outputs(76) <= a;
    layer5_outputs(77) <= not (a or b);
    layer5_outputs(78) <= a or b;
    layer5_outputs(79) <= b;
    layer5_outputs(80) <= a and b;
    layer5_outputs(81) <= a;
    layer5_outputs(82) <= a and not b;
    layer5_outputs(83) <= '1';
    layer5_outputs(84) <= a and b;
    layer5_outputs(85) <= a;
    layer5_outputs(86) <= not a;
    layer5_outputs(87) <= b and not a;
    layer5_outputs(88) <= a or b;
    layer5_outputs(89) <= not b;
    layer5_outputs(90) <= b;
    layer5_outputs(91) <= a and not b;
    layer5_outputs(92) <= b and not a;
    layer5_outputs(93) <= not a;
    layer5_outputs(94) <= a or b;
    layer5_outputs(95) <= not a;
    layer5_outputs(96) <= b and not a;
    layer5_outputs(97) <= b;
    layer5_outputs(98) <= a and not b;
    layer5_outputs(99) <= '0';
    layer5_outputs(100) <= not b;
    layer5_outputs(101) <= not b;
    layer5_outputs(102) <= not a or b;
    layer5_outputs(103) <= not a or b;
    layer5_outputs(104) <= not a;
    layer5_outputs(105) <= a;
    layer5_outputs(106) <= not (a or b);
    layer5_outputs(107) <= not b;
    layer5_outputs(108) <= not b;
    layer5_outputs(109) <= not a or b;
    layer5_outputs(110) <= a and b;
    layer5_outputs(111) <= a or b;
    layer5_outputs(112) <= not a;
    layer5_outputs(113) <= a xor b;
    layer5_outputs(114) <= a;
    layer5_outputs(115) <= a;
    layer5_outputs(116) <= a or b;
    layer5_outputs(117) <= not a or b;
    layer5_outputs(118) <= not (a xor b);
    layer5_outputs(119) <= not b or a;
    layer5_outputs(120) <= '1';
    layer5_outputs(121) <= b;
    layer5_outputs(122) <= not (a or b);
    layer5_outputs(123) <= a and not b;
    layer5_outputs(124) <= not b;
    layer5_outputs(125) <= a and not b;
    layer5_outputs(126) <= a;
    layer5_outputs(127) <= not (a xor b);
    layer5_outputs(128) <= not b or a;
    layer5_outputs(129) <= '0';
    layer5_outputs(130) <= a or b;
    layer5_outputs(131) <= a;
    layer5_outputs(132) <= not (a or b);
    layer5_outputs(133) <= a;
    layer5_outputs(134) <= not (a and b);
    layer5_outputs(135) <= b and not a;
    layer5_outputs(136) <= a xor b;
    layer5_outputs(137) <= not b;
    layer5_outputs(138) <= not a or b;
    layer5_outputs(139) <= not a;
    layer5_outputs(140) <= a and b;
    layer5_outputs(141) <= not b;
    layer5_outputs(142) <= not b or a;
    layer5_outputs(143) <= not a;
    layer5_outputs(144) <= not (a xor b);
    layer5_outputs(145) <= a xor b;
    layer5_outputs(146) <= a xor b;
    layer5_outputs(147) <= a xor b;
    layer5_outputs(148) <= not b or a;
    layer5_outputs(149) <= not b or a;
    layer5_outputs(150) <= a and b;
    layer5_outputs(151) <= not a;
    layer5_outputs(152) <= a and b;
    layer5_outputs(153) <= not b or a;
    layer5_outputs(154) <= b;
    layer5_outputs(155) <= not (a or b);
    layer5_outputs(156) <= a;
    layer5_outputs(157) <= not b;
    layer5_outputs(158) <= a and not b;
    layer5_outputs(159) <= b;
    layer5_outputs(160) <= not a;
    layer5_outputs(161) <= not b or a;
    layer5_outputs(162) <= '0';
    layer5_outputs(163) <= a or b;
    layer5_outputs(164) <= not b;
    layer5_outputs(165) <= a xor b;
    layer5_outputs(166) <= a or b;
    layer5_outputs(167) <= a and not b;
    layer5_outputs(168) <= b and not a;
    layer5_outputs(169) <= b and not a;
    layer5_outputs(170) <= not a or b;
    layer5_outputs(171) <= b;
    layer5_outputs(172) <= not (a and b);
    layer5_outputs(173) <= a and b;
    layer5_outputs(174) <= a xor b;
    layer5_outputs(175) <= b;
    layer5_outputs(176) <= not a;
    layer5_outputs(177) <= not (a or b);
    layer5_outputs(178) <= a and not b;
    layer5_outputs(179) <= not (a xor b);
    layer5_outputs(180) <= not (a xor b);
    layer5_outputs(181) <= not b;
    layer5_outputs(182) <= b and not a;
    layer5_outputs(183) <= not a or b;
    layer5_outputs(184) <= b;
    layer5_outputs(185) <= not b;
    layer5_outputs(186) <= not b or a;
    layer5_outputs(187) <= '0';
    layer5_outputs(188) <= not a or b;
    layer5_outputs(189) <= b and not a;
    layer5_outputs(190) <= a and b;
    layer5_outputs(191) <= b;
    layer5_outputs(192) <= not (a or b);
    layer5_outputs(193) <= not b;
    layer5_outputs(194) <= '0';
    layer5_outputs(195) <= not a;
    layer5_outputs(196) <= a;
    layer5_outputs(197) <= a and not b;
    layer5_outputs(198) <= a and b;
    layer5_outputs(199) <= a;
    layer5_outputs(200) <= not (a and b);
    layer5_outputs(201) <= '1';
    layer5_outputs(202) <= not (a and b);
    layer5_outputs(203) <= not (a and b);
    layer5_outputs(204) <= not b;
    layer5_outputs(205) <= a and b;
    layer5_outputs(206) <= b;
    layer5_outputs(207) <= a;
    layer5_outputs(208) <= b;
    layer5_outputs(209) <= not a or b;
    layer5_outputs(210) <= b and not a;
    layer5_outputs(211) <= not b;
    layer5_outputs(212) <= not a;
    layer5_outputs(213) <= a;
    layer5_outputs(214) <= '1';
    layer5_outputs(215) <= a or b;
    layer5_outputs(216) <= not a;
    layer5_outputs(217) <= not a;
    layer5_outputs(218) <= not a;
    layer5_outputs(219) <= not (a or b);
    layer5_outputs(220) <= not (a xor b);
    layer5_outputs(221) <= not a;
    layer5_outputs(222) <= a;
    layer5_outputs(223) <= b;
    layer5_outputs(224) <= not b;
    layer5_outputs(225) <= a and b;
    layer5_outputs(226) <= not a;
    layer5_outputs(227) <= not (a or b);
    layer5_outputs(228) <= not (a and b);
    layer5_outputs(229) <= a or b;
    layer5_outputs(230) <= a and not b;
    layer5_outputs(231) <= not (a and b);
    layer5_outputs(232) <= '0';
    layer5_outputs(233) <= not a;
    layer5_outputs(234) <= not a;
    layer5_outputs(235) <= b;
    layer5_outputs(236) <= a or b;
    layer5_outputs(237) <= '1';
    layer5_outputs(238) <= b;
    layer5_outputs(239) <= not (a and b);
    layer5_outputs(240) <= a and not b;
    layer5_outputs(241) <= not (a xor b);
    layer5_outputs(242) <= not b or a;
    layer5_outputs(243) <= a and b;
    layer5_outputs(244) <= not a;
    layer5_outputs(245) <= a;
    layer5_outputs(246) <= not b;
    layer5_outputs(247) <= not a;
    layer5_outputs(248) <= a or b;
    layer5_outputs(249) <= not a;
    layer5_outputs(250) <= not b;
    layer5_outputs(251) <= not a;
    layer5_outputs(252) <= a xor b;
    layer5_outputs(253) <= not b;
    layer5_outputs(254) <= not b;
    layer5_outputs(255) <= b;
    layer5_outputs(256) <= not (a and b);
    layer5_outputs(257) <= b;
    layer5_outputs(258) <= b;
    layer5_outputs(259) <= not b or a;
    layer5_outputs(260) <= not a;
    layer5_outputs(261) <= '1';
    layer5_outputs(262) <= not (a and b);
    layer5_outputs(263) <= not (a and b);
    layer5_outputs(264) <= '0';
    layer5_outputs(265) <= not b;
    layer5_outputs(266) <= not (a and b);
    layer5_outputs(267) <= a;
    layer5_outputs(268) <= a and not b;
    layer5_outputs(269) <= not a;
    layer5_outputs(270) <= not a;
    layer5_outputs(271) <= a and not b;
    layer5_outputs(272) <= not a or b;
    layer5_outputs(273) <= a and b;
    layer5_outputs(274) <= b;
    layer5_outputs(275) <= a or b;
    layer5_outputs(276) <= not a or b;
    layer5_outputs(277) <= '1';
    layer5_outputs(278) <= a;
    layer5_outputs(279) <= a xor b;
    layer5_outputs(280) <= not a;
    layer5_outputs(281) <= not (a and b);
    layer5_outputs(282) <= b and not a;
    layer5_outputs(283) <= b and not a;
    layer5_outputs(284) <= not b;
    layer5_outputs(285) <= not b or a;
    layer5_outputs(286) <= not (a xor b);
    layer5_outputs(287) <= not a or b;
    layer5_outputs(288) <= not a or b;
    layer5_outputs(289) <= not (a xor b);
    layer5_outputs(290) <= a and not b;
    layer5_outputs(291) <= a xor b;
    layer5_outputs(292) <= not a or b;
    layer5_outputs(293) <= a;
    layer5_outputs(294) <= a or b;
    layer5_outputs(295) <= a and b;
    layer5_outputs(296) <= b and not a;
    layer5_outputs(297) <= '1';
    layer5_outputs(298) <= a or b;
    layer5_outputs(299) <= a;
    layer5_outputs(300) <= a and b;
    layer5_outputs(301) <= not b;
    layer5_outputs(302) <= not b or a;
    layer5_outputs(303) <= b and not a;
    layer5_outputs(304) <= not (a and b);
    layer5_outputs(305) <= a and not b;
    layer5_outputs(306) <= a or b;
    layer5_outputs(307) <= b;
    layer5_outputs(308) <= not b;
    layer5_outputs(309) <= not a;
    layer5_outputs(310) <= a or b;
    layer5_outputs(311) <= '1';
    layer5_outputs(312) <= a or b;
    layer5_outputs(313) <= not a or b;
    layer5_outputs(314) <= not a or b;
    layer5_outputs(315) <= not b;
    layer5_outputs(316) <= a xor b;
    layer5_outputs(317) <= not (a and b);
    layer5_outputs(318) <= not a or b;
    layer5_outputs(319) <= '0';
    layer5_outputs(320) <= not (a or b);
    layer5_outputs(321) <= a;
    layer5_outputs(322) <= not a or b;
    layer5_outputs(323) <= not b;
    layer5_outputs(324) <= b;
    layer5_outputs(325) <= a and b;
    layer5_outputs(326) <= a and not b;
    layer5_outputs(327) <= b and not a;
    layer5_outputs(328) <= a;
    layer5_outputs(329) <= a and b;
    layer5_outputs(330) <= not b;
    layer5_outputs(331) <= b;
    layer5_outputs(332) <= a and not b;
    layer5_outputs(333) <= '1';
    layer5_outputs(334) <= a and b;
    layer5_outputs(335) <= a and not b;
    layer5_outputs(336) <= not b or a;
    layer5_outputs(337) <= '1';
    layer5_outputs(338) <= not a or b;
    layer5_outputs(339) <= '0';
    layer5_outputs(340) <= a;
    layer5_outputs(341) <= not b;
    layer5_outputs(342) <= a xor b;
    layer5_outputs(343) <= a or b;
    layer5_outputs(344) <= b and not a;
    layer5_outputs(345) <= not (a or b);
    layer5_outputs(346) <= '1';
    layer5_outputs(347) <= not a or b;
    layer5_outputs(348) <= a xor b;
    layer5_outputs(349) <= not a or b;
    layer5_outputs(350) <= b;
    layer5_outputs(351) <= '0';
    layer5_outputs(352) <= b;
    layer5_outputs(353) <= a;
    layer5_outputs(354) <= not a;
    layer5_outputs(355) <= b;
    layer5_outputs(356) <= a;
    layer5_outputs(357) <= not a;
    layer5_outputs(358) <= b and not a;
    layer5_outputs(359) <= not b or a;
    layer5_outputs(360) <= a or b;
    layer5_outputs(361) <= not (a or b);
    layer5_outputs(362) <= not a;
    layer5_outputs(363) <= not b or a;
    layer5_outputs(364) <= a and b;
    layer5_outputs(365) <= a and b;
    layer5_outputs(366) <= a and b;
    layer5_outputs(367) <= not a;
    layer5_outputs(368) <= a;
    layer5_outputs(369) <= a;
    layer5_outputs(370) <= a;
    layer5_outputs(371) <= a or b;
    layer5_outputs(372) <= a;
    layer5_outputs(373) <= a and b;
    layer5_outputs(374) <= not (a or b);
    layer5_outputs(375) <= not (a xor b);
    layer5_outputs(376) <= not b or a;
    layer5_outputs(377) <= b and not a;
    layer5_outputs(378) <= a or b;
    layer5_outputs(379) <= a;
    layer5_outputs(380) <= not a;
    layer5_outputs(381) <= b and not a;
    layer5_outputs(382) <= a;
    layer5_outputs(383) <= a xor b;
    layer5_outputs(384) <= not b;
    layer5_outputs(385) <= a xor b;
    layer5_outputs(386) <= '0';
    layer5_outputs(387) <= not (a xor b);
    layer5_outputs(388) <= a or b;
    layer5_outputs(389) <= not a or b;
    layer5_outputs(390) <= not b;
    layer5_outputs(391) <= not (a and b);
    layer5_outputs(392) <= a and b;
    layer5_outputs(393) <= a and b;
    layer5_outputs(394) <= not (a or b);
    layer5_outputs(395) <= not (a xor b);
    layer5_outputs(396) <= a and not b;
    layer5_outputs(397) <= b;
    layer5_outputs(398) <= a;
    layer5_outputs(399) <= b and not a;
    layer5_outputs(400) <= not a or b;
    layer5_outputs(401) <= '0';
    layer5_outputs(402) <= b and not a;
    layer5_outputs(403) <= not a or b;
    layer5_outputs(404) <= b;
    layer5_outputs(405) <= not b;
    layer5_outputs(406) <= '0';
    layer5_outputs(407) <= b;
    layer5_outputs(408) <= not (a and b);
    layer5_outputs(409) <= '0';
    layer5_outputs(410) <= b;
    layer5_outputs(411) <= not (a or b);
    layer5_outputs(412) <= not (a and b);
    layer5_outputs(413) <= '1';
    layer5_outputs(414) <= a or b;
    layer5_outputs(415) <= not (a and b);
    layer5_outputs(416) <= not a;
    layer5_outputs(417) <= b;
    layer5_outputs(418) <= b and not a;
    layer5_outputs(419) <= a xor b;
    layer5_outputs(420) <= b;
    layer5_outputs(421) <= not b;
    layer5_outputs(422) <= a or b;
    layer5_outputs(423) <= not (a and b);
    layer5_outputs(424) <= b and not a;
    layer5_outputs(425) <= not b or a;
    layer5_outputs(426) <= a or b;
    layer5_outputs(427) <= a and not b;
    layer5_outputs(428) <= not a or b;
    layer5_outputs(429) <= b;
    layer5_outputs(430) <= a or b;
    layer5_outputs(431) <= a and b;
    layer5_outputs(432) <= b and not a;
    layer5_outputs(433) <= '1';
    layer5_outputs(434) <= b;
    layer5_outputs(435) <= a and not b;
    layer5_outputs(436) <= b;
    layer5_outputs(437) <= b and not a;
    layer5_outputs(438) <= a xor b;
    layer5_outputs(439) <= a or b;
    layer5_outputs(440) <= not b or a;
    layer5_outputs(441) <= not a;
    layer5_outputs(442) <= not a;
    layer5_outputs(443) <= not a or b;
    layer5_outputs(444) <= '1';
    layer5_outputs(445) <= not b;
    layer5_outputs(446) <= a or b;
    layer5_outputs(447) <= not b or a;
    layer5_outputs(448) <= not b;
    layer5_outputs(449) <= a and not b;
    layer5_outputs(450) <= b and not a;
    layer5_outputs(451) <= '0';
    layer5_outputs(452) <= b;
    layer5_outputs(453) <= not b;
    layer5_outputs(454) <= '1';
    layer5_outputs(455) <= not (a or b);
    layer5_outputs(456) <= b and not a;
    layer5_outputs(457) <= not b;
    layer5_outputs(458) <= not (a or b);
    layer5_outputs(459) <= b;
    layer5_outputs(460) <= not (a xor b);
    layer5_outputs(461) <= '1';
    layer5_outputs(462) <= b;
    layer5_outputs(463) <= a and b;
    layer5_outputs(464) <= not b;
    layer5_outputs(465) <= b and not a;
    layer5_outputs(466) <= b;
    layer5_outputs(467) <= b;
    layer5_outputs(468) <= a and b;
    layer5_outputs(469) <= not a;
    layer5_outputs(470) <= not (a or b);
    layer5_outputs(471) <= not b;
    layer5_outputs(472) <= not a;
    layer5_outputs(473) <= b;
    layer5_outputs(474) <= not a;
    layer5_outputs(475) <= a;
    layer5_outputs(476) <= a and not b;
    layer5_outputs(477) <= not a;
    layer5_outputs(478) <= b and not a;
    layer5_outputs(479) <= a;
    layer5_outputs(480) <= not b or a;
    layer5_outputs(481) <= a;
    layer5_outputs(482) <= not a or b;
    layer5_outputs(483) <= not (a and b);
    layer5_outputs(484) <= not (a and b);
    layer5_outputs(485) <= not (a or b);
    layer5_outputs(486) <= not (a xor b);
    layer5_outputs(487) <= not b or a;
    layer5_outputs(488) <= a and b;
    layer5_outputs(489) <= not (a and b);
    layer5_outputs(490) <= not a;
    layer5_outputs(491) <= '1';
    layer5_outputs(492) <= a and not b;
    layer5_outputs(493) <= a or b;
    layer5_outputs(494) <= a and not b;
    layer5_outputs(495) <= not (a xor b);
    layer5_outputs(496) <= not b;
    layer5_outputs(497) <= not a or b;
    layer5_outputs(498) <= not b or a;
    layer5_outputs(499) <= not b or a;
    layer5_outputs(500) <= b;
    layer5_outputs(501) <= not (a xor b);
    layer5_outputs(502) <= not a;
    layer5_outputs(503) <= not a or b;
    layer5_outputs(504) <= '1';
    layer5_outputs(505) <= a and b;
    layer5_outputs(506) <= b;
    layer5_outputs(507) <= '1';
    layer5_outputs(508) <= not a;
    layer5_outputs(509) <= '1';
    layer5_outputs(510) <= a;
    layer5_outputs(511) <= not b;
    layer5_outputs(512) <= not a or b;
    layer5_outputs(513) <= a or b;
    layer5_outputs(514) <= not (a xor b);
    layer5_outputs(515) <= not a or b;
    layer5_outputs(516) <= not a or b;
    layer5_outputs(517) <= a and b;
    layer5_outputs(518) <= b;
    layer5_outputs(519) <= a and not b;
    layer5_outputs(520) <= not (a xor b);
    layer5_outputs(521) <= not a;
    layer5_outputs(522) <= not (a or b);
    layer5_outputs(523) <= a;
    layer5_outputs(524) <= a and not b;
    layer5_outputs(525) <= not b;
    layer5_outputs(526) <= a;
    layer5_outputs(527) <= not b or a;
    layer5_outputs(528) <= not (a and b);
    layer5_outputs(529) <= not a;
    layer5_outputs(530) <= not b;
    layer5_outputs(531) <= a or b;
    layer5_outputs(532) <= a;
    layer5_outputs(533) <= not a or b;
    layer5_outputs(534) <= b;
    layer5_outputs(535) <= b;
    layer5_outputs(536) <= a;
    layer5_outputs(537) <= a;
    layer5_outputs(538) <= not b or a;
    layer5_outputs(539) <= not (a and b);
    layer5_outputs(540) <= b and not a;
    layer5_outputs(541) <= not a;
    layer5_outputs(542) <= a or b;
    layer5_outputs(543) <= not b or a;
    layer5_outputs(544) <= not (a or b);
    layer5_outputs(545) <= not a;
    layer5_outputs(546) <= a and b;
    layer5_outputs(547) <= b;
    layer5_outputs(548) <= a and not b;
    layer5_outputs(549) <= a xor b;
    layer5_outputs(550) <= '0';
    layer5_outputs(551) <= not (a and b);
    layer5_outputs(552) <= not (a and b);
    layer5_outputs(553) <= a and b;
    layer5_outputs(554) <= b and not a;
    layer5_outputs(555) <= b and not a;
    layer5_outputs(556) <= not (a and b);
    layer5_outputs(557) <= not (a xor b);
    layer5_outputs(558) <= not b or a;
    layer5_outputs(559) <= not a or b;
    layer5_outputs(560) <= not b;
    layer5_outputs(561) <= '0';
    layer5_outputs(562) <= not a;
    layer5_outputs(563) <= not (a and b);
    layer5_outputs(564) <= a;
    layer5_outputs(565) <= not (a and b);
    layer5_outputs(566) <= b and not a;
    layer5_outputs(567) <= b;
    layer5_outputs(568) <= a;
    layer5_outputs(569) <= b and not a;
    layer5_outputs(570) <= not (a and b);
    layer5_outputs(571) <= a and not b;
    layer5_outputs(572) <= a;
    layer5_outputs(573) <= b;
    layer5_outputs(574) <= a;
    layer5_outputs(575) <= not a;
    layer5_outputs(576) <= '0';
    layer5_outputs(577) <= a and not b;
    layer5_outputs(578) <= '0';
    layer5_outputs(579) <= a;
    layer5_outputs(580) <= not b or a;
    layer5_outputs(581) <= not b;
    layer5_outputs(582) <= a;
    layer5_outputs(583) <= a;
    layer5_outputs(584) <= not (a and b);
    layer5_outputs(585) <= not (a or b);
    layer5_outputs(586) <= not b;
    layer5_outputs(587) <= a and not b;
    layer5_outputs(588) <= not (a or b);
    layer5_outputs(589) <= b and not a;
    layer5_outputs(590) <= a and not b;
    layer5_outputs(591) <= not b;
    layer5_outputs(592) <= not b;
    layer5_outputs(593) <= '0';
    layer5_outputs(594) <= b;
    layer5_outputs(595) <= a;
    layer5_outputs(596) <= not (a or b);
    layer5_outputs(597) <= b and not a;
    layer5_outputs(598) <= not a or b;
    layer5_outputs(599) <= not b or a;
    layer5_outputs(600) <= not b;
    layer5_outputs(601) <= not b;
    layer5_outputs(602) <= a;
    layer5_outputs(603) <= a and b;
    layer5_outputs(604) <= a;
    layer5_outputs(605) <= not a;
    layer5_outputs(606) <= a or b;
    layer5_outputs(607) <= b;
    layer5_outputs(608) <= a;
    layer5_outputs(609) <= not a;
    layer5_outputs(610) <= not (a or b);
    layer5_outputs(611) <= a;
    layer5_outputs(612) <= b;
    layer5_outputs(613) <= a;
    layer5_outputs(614) <= not b or a;
    layer5_outputs(615) <= a;
    layer5_outputs(616) <= not b;
    layer5_outputs(617) <= not (a xor b);
    layer5_outputs(618) <= not a;
    layer5_outputs(619) <= not b;
    layer5_outputs(620) <= '1';
    layer5_outputs(621) <= a or b;
    layer5_outputs(622) <= '0';
    layer5_outputs(623) <= a;
    layer5_outputs(624) <= not a or b;
    layer5_outputs(625) <= a xor b;
    layer5_outputs(626) <= a or b;
    layer5_outputs(627) <= not (a or b);
    layer5_outputs(628) <= not a;
    layer5_outputs(629) <= b and not a;
    layer5_outputs(630) <= not (a xor b);
    layer5_outputs(631) <= a and b;
    layer5_outputs(632) <= '1';
    layer5_outputs(633) <= '1';
    layer5_outputs(634) <= not (a or b);
    layer5_outputs(635) <= a;
    layer5_outputs(636) <= a;
    layer5_outputs(637) <= not b;
    layer5_outputs(638) <= '1';
    layer5_outputs(639) <= not b or a;
    layer5_outputs(640) <= b;
    layer5_outputs(641) <= a or b;
    layer5_outputs(642) <= not (a and b);
    layer5_outputs(643) <= b;
    layer5_outputs(644) <= not (a xor b);
    layer5_outputs(645) <= a xor b;
    layer5_outputs(646) <= a and not b;
    layer5_outputs(647) <= b and not a;
    layer5_outputs(648) <= '0';
    layer5_outputs(649) <= b;
    layer5_outputs(650) <= not a or b;
    layer5_outputs(651) <= not (a or b);
    layer5_outputs(652) <= b;
    layer5_outputs(653) <= not (a xor b);
    layer5_outputs(654) <= not b;
    layer5_outputs(655) <= a or b;
    layer5_outputs(656) <= not (a and b);
    layer5_outputs(657) <= not (a and b);
    layer5_outputs(658) <= not a;
    layer5_outputs(659) <= b;
    layer5_outputs(660) <= b and not a;
    layer5_outputs(661) <= not a or b;
    layer5_outputs(662) <= a xor b;
    layer5_outputs(663) <= not a;
    layer5_outputs(664) <= not (a and b);
    layer5_outputs(665) <= not (a or b);
    layer5_outputs(666) <= b;
    layer5_outputs(667) <= b and not a;
    layer5_outputs(668) <= not b;
    layer5_outputs(669) <= b;
    layer5_outputs(670) <= b;
    layer5_outputs(671) <= a;
    layer5_outputs(672) <= a and not b;
    layer5_outputs(673) <= not (a or b);
    layer5_outputs(674) <= not a;
    layer5_outputs(675) <= a and not b;
    layer5_outputs(676) <= not (a or b);
    layer5_outputs(677) <= a and not b;
    layer5_outputs(678) <= not (a or b);
    layer5_outputs(679) <= not b or a;
    layer5_outputs(680) <= a;
    layer5_outputs(681) <= a;
    layer5_outputs(682) <= '1';
    layer5_outputs(683) <= a;
    layer5_outputs(684) <= not a or b;
    layer5_outputs(685) <= a;
    layer5_outputs(686) <= not b or a;
    layer5_outputs(687) <= not a;
    layer5_outputs(688) <= b and not a;
    layer5_outputs(689) <= not a or b;
    layer5_outputs(690) <= not a;
    layer5_outputs(691) <= not (a and b);
    layer5_outputs(692) <= not a or b;
    layer5_outputs(693) <= not (a and b);
    layer5_outputs(694) <= not (a xor b);
    layer5_outputs(695) <= not (a or b);
    layer5_outputs(696) <= not (a and b);
    layer5_outputs(697) <= not (a or b);
    layer5_outputs(698) <= b;
    layer5_outputs(699) <= a or b;
    layer5_outputs(700) <= '0';
    layer5_outputs(701) <= b and not a;
    layer5_outputs(702) <= a and b;
    layer5_outputs(703) <= not (a and b);
    layer5_outputs(704) <= b;
    layer5_outputs(705) <= b and not a;
    layer5_outputs(706) <= not a;
    layer5_outputs(707) <= b;
    layer5_outputs(708) <= a or b;
    layer5_outputs(709) <= not b or a;
    layer5_outputs(710) <= not (a xor b);
    layer5_outputs(711) <= a and b;
    layer5_outputs(712) <= a and b;
    layer5_outputs(713) <= b;
    layer5_outputs(714) <= a or b;
    layer5_outputs(715) <= '0';
    layer5_outputs(716) <= a or b;
    layer5_outputs(717) <= not b;
    layer5_outputs(718) <= a or b;
    layer5_outputs(719) <= not (a and b);
    layer5_outputs(720) <= b and not a;
    layer5_outputs(721) <= not (a xor b);
    layer5_outputs(722) <= not a;
    layer5_outputs(723) <= '1';
    layer5_outputs(724) <= b and not a;
    layer5_outputs(725) <= a or b;
    layer5_outputs(726) <= a xor b;
    layer5_outputs(727) <= a and not b;
    layer5_outputs(728) <= a;
    layer5_outputs(729) <= '0';
    layer5_outputs(730) <= not b;
    layer5_outputs(731) <= a or b;
    layer5_outputs(732) <= a and b;
    layer5_outputs(733) <= not (a and b);
    layer5_outputs(734) <= not a or b;
    layer5_outputs(735) <= a or b;
    layer5_outputs(736) <= not a;
    layer5_outputs(737) <= a xor b;
    layer5_outputs(738) <= b and not a;
    layer5_outputs(739) <= a or b;
    layer5_outputs(740) <= a;
    layer5_outputs(741) <= a;
    layer5_outputs(742) <= not b;
    layer5_outputs(743) <= not (a and b);
    layer5_outputs(744) <= a;
    layer5_outputs(745) <= a;
    layer5_outputs(746) <= not b;
    layer5_outputs(747) <= not (a and b);
    layer5_outputs(748) <= not (a and b);
    layer5_outputs(749) <= not b;
    layer5_outputs(750) <= not (a xor b);
    layer5_outputs(751) <= not (a or b);
    layer5_outputs(752) <= not b or a;
    layer5_outputs(753) <= not (a xor b);
    layer5_outputs(754) <= not (a and b);
    layer5_outputs(755) <= not b;
    layer5_outputs(756) <= not a or b;
    layer5_outputs(757) <= a;
    layer5_outputs(758) <= b;
    layer5_outputs(759) <= not (a or b);
    layer5_outputs(760) <= not (a and b);
    layer5_outputs(761) <= a or b;
    layer5_outputs(762) <= not a;
    layer5_outputs(763) <= a and not b;
    layer5_outputs(764) <= a xor b;
    layer5_outputs(765) <= a and b;
    layer5_outputs(766) <= b;
    layer5_outputs(767) <= not a or b;
    layer5_outputs(768) <= b;
    layer5_outputs(769) <= a and b;
    layer5_outputs(770) <= '0';
    layer5_outputs(771) <= a and not b;
    layer5_outputs(772) <= not b;
    layer5_outputs(773) <= not b or a;
    layer5_outputs(774) <= b;
    layer5_outputs(775) <= not a;
    layer5_outputs(776) <= a and not b;
    layer5_outputs(777) <= not a or b;
    layer5_outputs(778) <= a;
    layer5_outputs(779) <= not (a xor b);
    layer5_outputs(780) <= not a;
    layer5_outputs(781) <= '1';
    layer5_outputs(782) <= a xor b;
    layer5_outputs(783) <= not a or b;
    layer5_outputs(784) <= not (a and b);
    layer5_outputs(785) <= not (a or b);
    layer5_outputs(786) <= not a or b;
    layer5_outputs(787) <= not (a or b);
    layer5_outputs(788) <= a;
    layer5_outputs(789) <= not b;
    layer5_outputs(790) <= not (a or b);
    layer5_outputs(791) <= not a;
    layer5_outputs(792) <= a and not b;
    layer5_outputs(793) <= a or b;
    layer5_outputs(794) <= not b or a;
    layer5_outputs(795) <= not b or a;
    layer5_outputs(796) <= '0';
    layer5_outputs(797) <= not b;
    layer5_outputs(798) <= b;
    layer5_outputs(799) <= not b or a;
    layer5_outputs(800) <= a;
    layer5_outputs(801) <= not b;
    layer5_outputs(802) <= '1';
    layer5_outputs(803) <= not a;
    layer5_outputs(804) <= a or b;
    layer5_outputs(805) <= '1';
    layer5_outputs(806) <= '1';
    layer5_outputs(807) <= not b;
    layer5_outputs(808) <= b;
    layer5_outputs(809) <= b and not a;
    layer5_outputs(810) <= b;
    layer5_outputs(811) <= a;
    layer5_outputs(812) <= b;
    layer5_outputs(813) <= not (a and b);
    layer5_outputs(814) <= a;
    layer5_outputs(815) <= a;
    layer5_outputs(816) <= '0';
    layer5_outputs(817) <= not a;
    layer5_outputs(818) <= not (a and b);
    layer5_outputs(819) <= not b;
    layer5_outputs(820) <= not (a xor b);
    layer5_outputs(821) <= not b;
    layer5_outputs(822) <= not (a xor b);
    layer5_outputs(823) <= not b;
    layer5_outputs(824) <= a and not b;
    layer5_outputs(825) <= a;
    layer5_outputs(826) <= b;
    layer5_outputs(827) <= a and not b;
    layer5_outputs(828) <= not a;
    layer5_outputs(829) <= b;
    layer5_outputs(830) <= a;
    layer5_outputs(831) <= '0';
    layer5_outputs(832) <= not a or b;
    layer5_outputs(833) <= '1';
    layer5_outputs(834) <= a;
    layer5_outputs(835) <= not b;
    layer5_outputs(836) <= not (a and b);
    layer5_outputs(837) <= a xor b;
    layer5_outputs(838) <= not a;
    layer5_outputs(839) <= a and not b;
    layer5_outputs(840) <= not a;
    layer5_outputs(841) <= a xor b;
    layer5_outputs(842) <= not a;
    layer5_outputs(843) <= not a;
    layer5_outputs(844) <= not a or b;
    layer5_outputs(845) <= not b;
    layer5_outputs(846) <= b;
    layer5_outputs(847) <= a or b;
    layer5_outputs(848) <= not a or b;
    layer5_outputs(849) <= a or b;
    layer5_outputs(850) <= a;
    layer5_outputs(851) <= a;
    layer5_outputs(852) <= not a or b;
    layer5_outputs(853) <= b;
    layer5_outputs(854) <= '1';
    layer5_outputs(855) <= b;
    layer5_outputs(856) <= b and not a;
    layer5_outputs(857) <= a;
    layer5_outputs(858) <= a and b;
    layer5_outputs(859) <= a and b;
    layer5_outputs(860) <= a;
    layer5_outputs(861) <= not a or b;
    layer5_outputs(862) <= a and b;
    layer5_outputs(863) <= a and b;
    layer5_outputs(864) <= not a;
    layer5_outputs(865) <= not b;
    layer5_outputs(866) <= a and b;
    layer5_outputs(867) <= not (a and b);
    layer5_outputs(868) <= not (a and b);
    layer5_outputs(869) <= a and b;
    layer5_outputs(870) <= a and b;
    layer5_outputs(871) <= not (a and b);
    layer5_outputs(872) <= not b or a;
    layer5_outputs(873) <= a and not b;
    layer5_outputs(874) <= b and not a;
    layer5_outputs(875) <= not (a and b);
    layer5_outputs(876) <= not a or b;
    layer5_outputs(877) <= not (a or b);
    layer5_outputs(878) <= a;
    layer5_outputs(879) <= not (a and b);
    layer5_outputs(880) <= '0';
    layer5_outputs(881) <= b and not a;
    layer5_outputs(882) <= b;
    layer5_outputs(883) <= a or b;
    layer5_outputs(884) <= a;
    layer5_outputs(885) <= not (a or b);
    layer5_outputs(886) <= '1';
    layer5_outputs(887) <= not b;
    layer5_outputs(888) <= not b;
    layer5_outputs(889) <= not b;
    layer5_outputs(890) <= b;
    layer5_outputs(891) <= not (a and b);
    layer5_outputs(892) <= not (a and b);
    layer5_outputs(893) <= a and not b;
    layer5_outputs(894) <= not a or b;
    layer5_outputs(895) <= not a;
    layer5_outputs(896) <= b;
    layer5_outputs(897) <= not b;
    layer5_outputs(898) <= a;
    layer5_outputs(899) <= not a or b;
    layer5_outputs(900) <= a;
    layer5_outputs(901) <= not (a or b);
    layer5_outputs(902) <= a and not b;
    layer5_outputs(903) <= a and not b;
    layer5_outputs(904) <= not b;
    layer5_outputs(905) <= not a or b;
    layer5_outputs(906) <= '0';
    layer5_outputs(907) <= b;
    layer5_outputs(908) <= a or b;
    layer5_outputs(909) <= not b;
    layer5_outputs(910) <= a or b;
    layer5_outputs(911) <= not a;
    layer5_outputs(912) <= not a or b;
    layer5_outputs(913) <= a or b;
    layer5_outputs(914) <= a or b;
    layer5_outputs(915) <= a;
    layer5_outputs(916) <= b;
    layer5_outputs(917) <= not (a xor b);
    layer5_outputs(918) <= b and not a;
    layer5_outputs(919) <= not (a or b);
    layer5_outputs(920) <= a or b;
    layer5_outputs(921) <= not a or b;
    layer5_outputs(922) <= a or b;
    layer5_outputs(923) <= not b or a;
    layer5_outputs(924) <= not a or b;
    layer5_outputs(925) <= a and b;
    layer5_outputs(926) <= not a or b;
    layer5_outputs(927) <= not (a and b);
    layer5_outputs(928) <= not a or b;
    layer5_outputs(929) <= not a or b;
    layer5_outputs(930) <= b;
    layer5_outputs(931) <= a and not b;
    layer5_outputs(932) <= a xor b;
    layer5_outputs(933) <= a and b;
    layer5_outputs(934) <= a and b;
    layer5_outputs(935) <= a;
    layer5_outputs(936) <= a;
    layer5_outputs(937) <= not b;
    layer5_outputs(938) <= not a;
    layer5_outputs(939) <= a and b;
    layer5_outputs(940) <= not (a xor b);
    layer5_outputs(941) <= b and not a;
    layer5_outputs(942) <= b and not a;
    layer5_outputs(943) <= not a or b;
    layer5_outputs(944) <= b;
    layer5_outputs(945) <= not a;
    layer5_outputs(946) <= a xor b;
    layer5_outputs(947) <= b;
    layer5_outputs(948) <= b;
    layer5_outputs(949) <= '0';
    layer5_outputs(950) <= not a;
    layer5_outputs(951) <= not a;
    layer5_outputs(952) <= not a;
    layer5_outputs(953) <= not a;
    layer5_outputs(954) <= not (a or b);
    layer5_outputs(955) <= not a;
    layer5_outputs(956) <= not (a or b);
    layer5_outputs(957) <= not b;
    layer5_outputs(958) <= not (a and b);
    layer5_outputs(959) <= not b or a;
    layer5_outputs(960) <= not (a or b);
    layer5_outputs(961) <= not (a or b);
    layer5_outputs(962) <= b;
    layer5_outputs(963) <= a and not b;
    layer5_outputs(964) <= a and b;
    layer5_outputs(965) <= a or b;
    layer5_outputs(966) <= b;
    layer5_outputs(967) <= not b or a;
    layer5_outputs(968) <= not (a xor b);
    layer5_outputs(969) <= b;
    layer5_outputs(970) <= a and not b;
    layer5_outputs(971) <= not b;
    layer5_outputs(972) <= not (a or b);
    layer5_outputs(973) <= b and not a;
    layer5_outputs(974) <= '1';
    layer5_outputs(975) <= a;
    layer5_outputs(976) <= not a;
    layer5_outputs(977) <= b;
    layer5_outputs(978) <= b;
    layer5_outputs(979) <= not a;
    layer5_outputs(980) <= a and not b;
    layer5_outputs(981) <= a and not b;
    layer5_outputs(982) <= a and b;
    layer5_outputs(983) <= a and b;
    layer5_outputs(984) <= '1';
    layer5_outputs(985) <= b;
    layer5_outputs(986) <= not (a and b);
    layer5_outputs(987) <= a;
    layer5_outputs(988) <= a or b;
    layer5_outputs(989) <= b and not a;
    layer5_outputs(990) <= not b;
    layer5_outputs(991) <= not (a and b);
    layer5_outputs(992) <= not (a xor b);
    layer5_outputs(993) <= not a;
    layer5_outputs(994) <= b;
    layer5_outputs(995) <= not b or a;
    layer5_outputs(996) <= a;
    layer5_outputs(997) <= not a;
    layer5_outputs(998) <= a and not b;
    layer5_outputs(999) <= a and not b;
    layer5_outputs(1000) <= not (a and b);
    layer5_outputs(1001) <= a xor b;
    layer5_outputs(1002) <= not (a xor b);
    layer5_outputs(1003) <= not b or a;
    layer5_outputs(1004) <= b;
    layer5_outputs(1005) <= not (a xor b);
    layer5_outputs(1006) <= a and b;
    layer5_outputs(1007) <= not (a or b);
    layer5_outputs(1008) <= not a;
    layer5_outputs(1009) <= not a or b;
    layer5_outputs(1010) <= not b;
    layer5_outputs(1011) <= b and not a;
    layer5_outputs(1012) <= not a;
    layer5_outputs(1013) <= '0';
    layer5_outputs(1014) <= b;
    layer5_outputs(1015) <= not a or b;
    layer5_outputs(1016) <= not (a xor b);
    layer5_outputs(1017) <= a and b;
    layer5_outputs(1018) <= not (a and b);
    layer5_outputs(1019) <= not a;
    layer5_outputs(1020) <= '0';
    layer5_outputs(1021) <= a or b;
    layer5_outputs(1022) <= a xor b;
    layer5_outputs(1023) <= not a or b;
    layer5_outputs(1024) <= not a;
    layer5_outputs(1025) <= not (a or b);
    layer5_outputs(1026) <= a or b;
    layer5_outputs(1027) <= not (a or b);
    layer5_outputs(1028) <= '1';
    layer5_outputs(1029) <= not a or b;
    layer5_outputs(1030) <= a or b;
    layer5_outputs(1031) <= not (a xor b);
    layer5_outputs(1032) <= a and b;
    layer5_outputs(1033) <= b;
    layer5_outputs(1034) <= a and not b;
    layer5_outputs(1035) <= not (a and b);
    layer5_outputs(1036) <= b;
    layer5_outputs(1037) <= '0';
    layer5_outputs(1038) <= '1';
    layer5_outputs(1039) <= not b or a;
    layer5_outputs(1040) <= not (a and b);
    layer5_outputs(1041) <= a;
    layer5_outputs(1042) <= not b;
    layer5_outputs(1043) <= b and not a;
    layer5_outputs(1044) <= not (a and b);
    layer5_outputs(1045) <= a and not b;
    layer5_outputs(1046) <= not b;
    layer5_outputs(1047) <= not (a xor b);
    layer5_outputs(1048) <= a xor b;
    layer5_outputs(1049) <= a xor b;
    layer5_outputs(1050) <= not b or a;
    layer5_outputs(1051) <= b and not a;
    layer5_outputs(1052) <= '1';
    layer5_outputs(1053) <= not (a and b);
    layer5_outputs(1054) <= not b or a;
    layer5_outputs(1055) <= not b or a;
    layer5_outputs(1056) <= not a or b;
    layer5_outputs(1057) <= '0';
    layer5_outputs(1058) <= not b or a;
    layer5_outputs(1059) <= a xor b;
    layer5_outputs(1060) <= not (a xor b);
    layer5_outputs(1061) <= a;
    layer5_outputs(1062) <= b and not a;
    layer5_outputs(1063) <= a or b;
    layer5_outputs(1064) <= b;
    layer5_outputs(1065) <= not (a or b);
    layer5_outputs(1066) <= a;
    layer5_outputs(1067) <= not b;
    layer5_outputs(1068) <= a;
    layer5_outputs(1069) <= a or b;
    layer5_outputs(1070) <= b;
    layer5_outputs(1071) <= a;
    layer5_outputs(1072) <= not b;
    layer5_outputs(1073) <= not a;
    layer5_outputs(1074) <= not b or a;
    layer5_outputs(1075) <= a or b;
    layer5_outputs(1076) <= b;
    layer5_outputs(1077) <= a and not b;
    layer5_outputs(1078) <= a and not b;
    layer5_outputs(1079) <= a;
    layer5_outputs(1080) <= a;
    layer5_outputs(1081) <= b and not a;
    layer5_outputs(1082) <= not b or a;
    layer5_outputs(1083) <= b;
    layer5_outputs(1084) <= a;
    layer5_outputs(1085) <= b and not a;
    layer5_outputs(1086) <= not (a and b);
    layer5_outputs(1087) <= '1';
    layer5_outputs(1088) <= a or b;
    layer5_outputs(1089) <= not a or b;
    layer5_outputs(1090) <= '0';
    layer5_outputs(1091) <= not a or b;
    layer5_outputs(1092) <= not (a and b);
    layer5_outputs(1093) <= not (a or b);
    layer5_outputs(1094) <= a;
    layer5_outputs(1095) <= b;
    layer5_outputs(1096) <= not b or a;
    layer5_outputs(1097) <= a and not b;
    layer5_outputs(1098) <= not a;
    layer5_outputs(1099) <= b and not a;
    layer5_outputs(1100) <= a;
    layer5_outputs(1101) <= not (a or b);
    layer5_outputs(1102) <= b;
    layer5_outputs(1103) <= not b;
    layer5_outputs(1104) <= b;
    layer5_outputs(1105) <= not (a and b);
    layer5_outputs(1106) <= a and b;
    layer5_outputs(1107) <= not b;
    layer5_outputs(1108) <= not b;
    layer5_outputs(1109) <= not a;
    layer5_outputs(1110) <= '1';
    layer5_outputs(1111) <= not (a or b);
    layer5_outputs(1112) <= a and not b;
    layer5_outputs(1113) <= a and not b;
    layer5_outputs(1114) <= a and b;
    layer5_outputs(1115) <= not (a or b);
    layer5_outputs(1116) <= not b or a;
    layer5_outputs(1117) <= not (a xor b);
    layer5_outputs(1118) <= a and not b;
    layer5_outputs(1119) <= a and b;
    layer5_outputs(1120) <= not (a and b);
    layer5_outputs(1121) <= not a;
    layer5_outputs(1122) <= not a;
    layer5_outputs(1123) <= '0';
    layer5_outputs(1124) <= '0';
    layer5_outputs(1125) <= not b;
    layer5_outputs(1126) <= a and not b;
    layer5_outputs(1127) <= not a or b;
    layer5_outputs(1128) <= a xor b;
    layer5_outputs(1129) <= not (a and b);
    layer5_outputs(1130) <= '1';
    layer5_outputs(1131) <= not b or a;
    layer5_outputs(1132) <= a or b;
    layer5_outputs(1133) <= a;
    layer5_outputs(1134) <= not a;
    layer5_outputs(1135) <= not b;
    layer5_outputs(1136) <= b and not a;
    layer5_outputs(1137) <= not b;
    layer5_outputs(1138) <= not b;
    layer5_outputs(1139) <= '1';
    layer5_outputs(1140) <= b;
    layer5_outputs(1141) <= not (a or b);
    layer5_outputs(1142) <= b;
    layer5_outputs(1143) <= a and b;
    layer5_outputs(1144) <= not (a xor b);
    layer5_outputs(1145) <= a or b;
    layer5_outputs(1146) <= not b;
    layer5_outputs(1147) <= a and b;
    layer5_outputs(1148) <= not (a xor b);
    layer5_outputs(1149) <= not (a and b);
    layer5_outputs(1150) <= not a or b;
    layer5_outputs(1151) <= not (a xor b);
    layer5_outputs(1152) <= a;
    layer5_outputs(1153) <= not (a or b);
    layer5_outputs(1154) <= a and not b;
    layer5_outputs(1155) <= '0';
    layer5_outputs(1156) <= not b;
    layer5_outputs(1157) <= not a;
    layer5_outputs(1158) <= not (a xor b);
    layer5_outputs(1159) <= not (a or b);
    layer5_outputs(1160) <= not a;
    layer5_outputs(1161) <= not b;
    layer5_outputs(1162) <= '0';
    layer5_outputs(1163) <= a and b;
    layer5_outputs(1164) <= b and not a;
    layer5_outputs(1165) <= b;
    layer5_outputs(1166) <= not (a and b);
    layer5_outputs(1167) <= not a or b;
    layer5_outputs(1168) <= a and b;
    layer5_outputs(1169) <= a and not b;
    layer5_outputs(1170) <= b and not a;
    layer5_outputs(1171) <= not a or b;
    layer5_outputs(1172) <= a and b;
    layer5_outputs(1173) <= b;
    layer5_outputs(1174) <= b;
    layer5_outputs(1175) <= not (a or b);
    layer5_outputs(1176) <= b;
    layer5_outputs(1177) <= not (a and b);
    layer5_outputs(1178) <= a and not b;
    layer5_outputs(1179) <= a;
    layer5_outputs(1180) <= not b;
    layer5_outputs(1181) <= not a;
    layer5_outputs(1182) <= '1';
    layer5_outputs(1183) <= not (a and b);
    layer5_outputs(1184) <= not (a and b);
    layer5_outputs(1185) <= b;
    layer5_outputs(1186) <= b;
    layer5_outputs(1187) <= not a;
    layer5_outputs(1188) <= a and not b;
    layer5_outputs(1189) <= b;
    layer5_outputs(1190) <= a xor b;
    layer5_outputs(1191) <= '1';
    layer5_outputs(1192) <= b;
    layer5_outputs(1193) <= a and not b;
    layer5_outputs(1194) <= a and not b;
    layer5_outputs(1195) <= a or b;
    layer5_outputs(1196) <= a and not b;
    layer5_outputs(1197) <= not (a or b);
    layer5_outputs(1198) <= not a;
    layer5_outputs(1199) <= b;
    layer5_outputs(1200) <= b and not a;
    layer5_outputs(1201) <= b and not a;
    layer5_outputs(1202) <= a and b;
    layer5_outputs(1203) <= a and b;
    layer5_outputs(1204) <= '1';
    layer5_outputs(1205) <= not a;
    layer5_outputs(1206) <= b and not a;
    layer5_outputs(1207) <= not b or a;
    layer5_outputs(1208) <= a and b;
    layer5_outputs(1209) <= not (a or b);
    layer5_outputs(1210) <= not b or a;
    layer5_outputs(1211) <= '0';
    layer5_outputs(1212) <= a;
    layer5_outputs(1213) <= not a;
    layer5_outputs(1214) <= a and not b;
    layer5_outputs(1215) <= a and not b;
    layer5_outputs(1216) <= not a;
    layer5_outputs(1217) <= not a or b;
    layer5_outputs(1218) <= not b;
    layer5_outputs(1219) <= a;
    layer5_outputs(1220) <= b;
    layer5_outputs(1221) <= not a;
    layer5_outputs(1222) <= '1';
    layer5_outputs(1223) <= a;
    layer5_outputs(1224) <= a and not b;
    layer5_outputs(1225) <= not b;
    layer5_outputs(1226) <= b;
    layer5_outputs(1227) <= not (a xor b);
    layer5_outputs(1228) <= not a;
    layer5_outputs(1229) <= not b or a;
    layer5_outputs(1230) <= not b;
    layer5_outputs(1231) <= not a;
    layer5_outputs(1232) <= not a;
    layer5_outputs(1233) <= a and not b;
    layer5_outputs(1234) <= not (a and b);
    layer5_outputs(1235) <= a xor b;
    layer5_outputs(1236) <= a;
    layer5_outputs(1237) <= not (a and b);
    layer5_outputs(1238) <= a xor b;
    layer5_outputs(1239) <= a and b;
    layer5_outputs(1240) <= not a;
    layer5_outputs(1241) <= b and not a;
    layer5_outputs(1242) <= a and not b;
    layer5_outputs(1243) <= not (a or b);
    layer5_outputs(1244) <= not a or b;
    layer5_outputs(1245) <= not a or b;
    layer5_outputs(1246) <= not a or b;
    layer5_outputs(1247) <= '1';
    layer5_outputs(1248) <= b;
    layer5_outputs(1249) <= b;
    layer5_outputs(1250) <= a and b;
    layer5_outputs(1251) <= not (a or b);
    layer5_outputs(1252) <= not a or b;
    layer5_outputs(1253) <= a;
    layer5_outputs(1254) <= a;
    layer5_outputs(1255) <= not (a xor b);
    layer5_outputs(1256) <= not a;
    layer5_outputs(1257) <= not (a xor b);
    layer5_outputs(1258) <= not a;
    layer5_outputs(1259) <= a or b;
    layer5_outputs(1260) <= not (a or b);
    layer5_outputs(1261) <= not (a or b);
    layer5_outputs(1262) <= not a or b;
    layer5_outputs(1263) <= not a or b;
    layer5_outputs(1264) <= a and b;
    layer5_outputs(1265) <= a or b;
    layer5_outputs(1266) <= not a or b;
    layer5_outputs(1267) <= not b or a;
    layer5_outputs(1268) <= a or b;
    layer5_outputs(1269) <= a and b;
    layer5_outputs(1270) <= not b or a;
    layer5_outputs(1271) <= a xor b;
    layer5_outputs(1272) <= not (a xor b);
    layer5_outputs(1273) <= not a;
    layer5_outputs(1274) <= not a or b;
    layer5_outputs(1275) <= not a;
    layer5_outputs(1276) <= not (a xor b);
    layer5_outputs(1277) <= not b or a;
    layer5_outputs(1278) <= not b or a;
    layer5_outputs(1279) <= '0';
    layer5_outputs(1280) <= a and b;
    layer5_outputs(1281) <= a or b;
    layer5_outputs(1282) <= not a or b;
    layer5_outputs(1283) <= a xor b;
    layer5_outputs(1284) <= a and not b;
    layer5_outputs(1285) <= not a or b;
    layer5_outputs(1286) <= b;
    layer5_outputs(1287) <= b and not a;
    layer5_outputs(1288) <= a or b;
    layer5_outputs(1289) <= b;
    layer5_outputs(1290) <= a;
    layer5_outputs(1291) <= not b or a;
    layer5_outputs(1292) <= not (a or b);
    layer5_outputs(1293) <= not b;
    layer5_outputs(1294) <= b and not a;
    layer5_outputs(1295) <= a and not b;
    layer5_outputs(1296) <= b;
    layer5_outputs(1297) <= a;
    layer5_outputs(1298) <= not b;
    layer5_outputs(1299) <= not (a and b);
    layer5_outputs(1300) <= b and not a;
    layer5_outputs(1301) <= not (a and b);
    layer5_outputs(1302) <= not a;
    layer5_outputs(1303) <= '1';
    layer5_outputs(1304) <= '0';
    layer5_outputs(1305) <= '1';
    layer5_outputs(1306) <= not b or a;
    layer5_outputs(1307) <= b and not a;
    layer5_outputs(1308) <= not (a and b);
    layer5_outputs(1309) <= not (a or b);
    layer5_outputs(1310) <= not b or a;
    layer5_outputs(1311) <= a;
    layer5_outputs(1312) <= b;
    layer5_outputs(1313) <= a and b;
    layer5_outputs(1314) <= b and not a;
    layer5_outputs(1315) <= a and b;
    layer5_outputs(1316) <= not (a xor b);
    layer5_outputs(1317) <= b and not a;
    layer5_outputs(1318) <= not a or b;
    layer5_outputs(1319) <= b and not a;
    layer5_outputs(1320) <= '1';
    layer5_outputs(1321) <= not a;
    layer5_outputs(1322) <= not (a xor b);
    layer5_outputs(1323) <= not a or b;
    layer5_outputs(1324) <= a and not b;
    layer5_outputs(1325) <= not (a and b);
    layer5_outputs(1326) <= a or b;
    layer5_outputs(1327) <= a and not b;
    layer5_outputs(1328) <= not a or b;
    layer5_outputs(1329) <= not (a xor b);
    layer5_outputs(1330) <= a and b;
    layer5_outputs(1331) <= a and not b;
    layer5_outputs(1332) <= '1';
    layer5_outputs(1333) <= a;
    layer5_outputs(1334) <= a or b;
    layer5_outputs(1335) <= not a;
    layer5_outputs(1336) <= b and not a;
    layer5_outputs(1337) <= not b;
    layer5_outputs(1338) <= not (a and b);
    layer5_outputs(1339) <= not b or a;
    layer5_outputs(1340) <= '0';
    layer5_outputs(1341) <= not (a or b);
    layer5_outputs(1342) <= a xor b;
    layer5_outputs(1343) <= a and b;
    layer5_outputs(1344) <= not a;
    layer5_outputs(1345) <= a;
    layer5_outputs(1346) <= not b or a;
    layer5_outputs(1347) <= not a;
    layer5_outputs(1348) <= b;
    layer5_outputs(1349) <= a and b;
    layer5_outputs(1350) <= '1';
    layer5_outputs(1351) <= a or b;
    layer5_outputs(1352) <= a;
    layer5_outputs(1353) <= not (a and b);
    layer5_outputs(1354) <= a and b;
    layer5_outputs(1355) <= a or b;
    layer5_outputs(1356) <= b;
    layer5_outputs(1357) <= not a;
    layer5_outputs(1358) <= a;
    layer5_outputs(1359) <= a and not b;
    layer5_outputs(1360) <= a and not b;
    layer5_outputs(1361) <= '0';
    layer5_outputs(1362) <= not (a and b);
    layer5_outputs(1363) <= a and b;
    layer5_outputs(1364) <= not a;
    layer5_outputs(1365) <= not b;
    layer5_outputs(1366) <= not b or a;
    layer5_outputs(1367) <= '0';
    layer5_outputs(1368) <= not a or b;
    layer5_outputs(1369) <= b and not a;
    layer5_outputs(1370) <= not b or a;
    layer5_outputs(1371) <= '1';
    layer5_outputs(1372) <= not (a or b);
    layer5_outputs(1373) <= a and not b;
    layer5_outputs(1374) <= not (a or b);
    layer5_outputs(1375) <= not a;
    layer5_outputs(1376) <= not a;
    layer5_outputs(1377) <= a or b;
    layer5_outputs(1378) <= a xor b;
    layer5_outputs(1379) <= b;
    layer5_outputs(1380) <= a;
    layer5_outputs(1381) <= not a or b;
    layer5_outputs(1382) <= not (a or b);
    layer5_outputs(1383) <= a and not b;
    layer5_outputs(1384) <= a and b;
    layer5_outputs(1385) <= a and not b;
    layer5_outputs(1386) <= '0';
    layer5_outputs(1387) <= a or b;
    layer5_outputs(1388) <= b and not a;
    layer5_outputs(1389) <= a or b;
    layer5_outputs(1390) <= '0';
    layer5_outputs(1391) <= a or b;
    layer5_outputs(1392) <= a and b;
    layer5_outputs(1393) <= b;
    layer5_outputs(1394) <= a and not b;
    layer5_outputs(1395) <= a and not b;
    layer5_outputs(1396) <= b;
    layer5_outputs(1397) <= '0';
    layer5_outputs(1398) <= '0';
    layer5_outputs(1399) <= a;
    layer5_outputs(1400) <= b;
    layer5_outputs(1401) <= not (a xor b);
    layer5_outputs(1402) <= a and b;
    layer5_outputs(1403) <= not (a and b);
    layer5_outputs(1404) <= a and not b;
    layer5_outputs(1405) <= a or b;
    layer5_outputs(1406) <= '0';
    layer5_outputs(1407) <= a;
    layer5_outputs(1408) <= a and b;
    layer5_outputs(1409) <= not (a and b);
    layer5_outputs(1410) <= not a or b;
    layer5_outputs(1411) <= a and b;
    layer5_outputs(1412) <= a;
    layer5_outputs(1413) <= not b;
    layer5_outputs(1414) <= a xor b;
    layer5_outputs(1415) <= not (a or b);
    layer5_outputs(1416) <= a or b;
    layer5_outputs(1417) <= not (a and b);
    layer5_outputs(1418) <= not b or a;
    layer5_outputs(1419) <= '1';
    layer5_outputs(1420) <= not a;
    layer5_outputs(1421) <= not a or b;
    layer5_outputs(1422) <= b;
    layer5_outputs(1423) <= a or b;
    layer5_outputs(1424) <= not b;
    layer5_outputs(1425) <= not b;
    layer5_outputs(1426) <= b;
    layer5_outputs(1427) <= not (a or b);
    layer5_outputs(1428) <= b;
    layer5_outputs(1429) <= b;
    layer5_outputs(1430) <= a and not b;
    layer5_outputs(1431) <= a;
    layer5_outputs(1432) <= a and not b;
    layer5_outputs(1433) <= not (a or b);
    layer5_outputs(1434) <= not a or b;
    layer5_outputs(1435) <= not a or b;
    layer5_outputs(1436) <= a or b;
    layer5_outputs(1437) <= b and not a;
    layer5_outputs(1438) <= a and b;
    layer5_outputs(1439) <= not (a or b);
    layer5_outputs(1440) <= a;
    layer5_outputs(1441) <= b;
    layer5_outputs(1442) <= not b or a;
    layer5_outputs(1443) <= not (a xor b);
    layer5_outputs(1444) <= a xor b;
    layer5_outputs(1445) <= b;
    layer5_outputs(1446) <= not (a and b);
    layer5_outputs(1447) <= b;
    layer5_outputs(1448) <= a;
    layer5_outputs(1449) <= not (a or b);
    layer5_outputs(1450) <= b and not a;
    layer5_outputs(1451) <= not b;
    layer5_outputs(1452) <= not (a xor b);
    layer5_outputs(1453) <= not a;
    layer5_outputs(1454) <= a xor b;
    layer5_outputs(1455) <= not b;
    layer5_outputs(1456) <= not (a and b);
    layer5_outputs(1457) <= b and not a;
    layer5_outputs(1458) <= a;
    layer5_outputs(1459) <= not b or a;
    layer5_outputs(1460) <= b;
    layer5_outputs(1461) <= '1';
    layer5_outputs(1462) <= not (a and b);
    layer5_outputs(1463) <= not a or b;
    layer5_outputs(1464) <= b and not a;
    layer5_outputs(1465) <= a and b;
    layer5_outputs(1466) <= a;
    layer5_outputs(1467) <= not a;
    layer5_outputs(1468) <= not a;
    layer5_outputs(1469) <= not a or b;
    layer5_outputs(1470) <= not a or b;
    layer5_outputs(1471) <= not b or a;
    layer5_outputs(1472) <= '1';
    layer5_outputs(1473) <= a and not b;
    layer5_outputs(1474) <= a or b;
    layer5_outputs(1475) <= not b;
    layer5_outputs(1476) <= a and b;
    layer5_outputs(1477) <= a and b;
    layer5_outputs(1478) <= not b;
    layer5_outputs(1479) <= not a;
    layer5_outputs(1480) <= '1';
    layer5_outputs(1481) <= b;
    layer5_outputs(1482) <= not b;
    layer5_outputs(1483) <= a and not b;
    layer5_outputs(1484) <= not a or b;
    layer5_outputs(1485) <= a xor b;
    layer5_outputs(1486) <= not a or b;
    layer5_outputs(1487) <= not (a xor b);
    layer5_outputs(1488) <= a and not b;
    layer5_outputs(1489) <= a and b;
    layer5_outputs(1490) <= a and b;
    layer5_outputs(1491) <= a;
    layer5_outputs(1492) <= not (a and b);
    layer5_outputs(1493) <= b;
    layer5_outputs(1494) <= b;
    layer5_outputs(1495) <= not (a or b);
    layer5_outputs(1496) <= not b;
    layer5_outputs(1497) <= not b;
    layer5_outputs(1498) <= not a;
    layer5_outputs(1499) <= a or b;
    layer5_outputs(1500) <= not a;
    layer5_outputs(1501) <= not a or b;
    layer5_outputs(1502) <= '1';
    layer5_outputs(1503) <= not b;
    layer5_outputs(1504) <= not b or a;
    layer5_outputs(1505) <= not b or a;
    layer5_outputs(1506) <= not (a and b);
    layer5_outputs(1507) <= b;
    layer5_outputs(1508) <= b and not a;
    layer5_outputs(1509) <= b and not a;
    layer5_outputs(1510) <= b;
    layer5_outputs(1511) <= not a;
    layer5_outputs(1512) <= not (a or b);
    layer5_outputs(1513) <= '1';
    layer5_outputs(1514) <= a and not b;
    layer5_outputs(1515) <= not (a or b);
    layer5_outputs(1516) <= not b or a;
    layer5_outputs(1517) <= not b;
    layer5_outputs(1518) <= not a;
    layer5_outputs(1519) <= '0';
    layer5_outputs(1520) <= not b or a;
    layer5_outputs(1521) <= a;
    layer5_outputs(1522) <= not (a and b);
    layer5_outputs(1523) <= a xor b;
    layer5_outputs(1524) <= not b or a;
    layer5_outputs(1525) <= a xor b;
    layer5_outputs(1526) <= b;
    layer5_outputs(1527) <= a and b;
    layer5_outputs(1528) <= not a;
    layer5_outputs(1529) <= not (a and b);
    layer5_outputs(1530) <= a;
    layer5_outputs(1531) <= not a;
    layer5_outputs(1532) <= not a;
    layer5_outputs(1533) <= a and not b;
    layer5_outputs(1534) <= a and not b;
    layer5_outputs(1535) <= not (a or b);
    layer5_outputs(1536) <= a;
    layer5_outputs(1537) <= not b or a;
    layer5_outputs(1538) <= not b;
    layer5_outputs(1539) <= not b;
    layer5_outputs(1540) <= not b or a;
    layer5_outputs(1541) <= not b or a;
    layer5_outputs(1542) <= a xor b;
    layer5_outputs(1543) <= a and b;
    layer5_outputs(1544) <= not (a or b);
    layer5_outputs(1545) <= a and not b;
    layer5_outputs(1546) <= b;
    layer5_outputs(1547) <= not (a and b);
    layer5_outputs(1548) <= not (a or b);
    layer5_outputs(1549) <= b;
    layer5_outputs(1550) <= not b or a;
    layer5_outputs(1551) <= not a or b;
    layer5_outputs(1552) <= a or b;
    layer5_outputs(1553) <= a;
    layer5_outputs(1554) <= b;
    layer5_outputs(1555) <= not b;
    layer5_outputs(1556) <= not a or b;
    layer5_outputs(1557) <= not (a and b);
    layer5_outputs(1558) <= '0';
    layer5_outputs(1559) <= a and not b;
    layer5_outputs(1560) <= not b;
    layer5_outputs(1561) <= a or b;
    layer5_outputs(1562) <= a and b;
    layer5_outputs(1563) <= b;
    layer5_outputs(1564) <= not a;
    layer5_outputs(1565) <= not a or b;
    layer5_outputs(1566) <= not (a or b);
    layer5_outputs(1567) <= not b;
    layer5_outputs(1568) <= '1';
    layer5_outputs(1569) <= '1';
    layer5_outputs(1570) <= a xor b;
    layer5_outputs(1571) <= not b or a;
    layer5_outputs(1572) <= a or b;
    layer5_outputs(1573) <= a or b;
    layer5_outputs(1574) <= a and not b;
    layer5_outputs(1575) <= a and not b;
    layer5_outputs(1576) <= '1';
    layer5_outputs(1577) <= b;
    layer5_outputs(1578) <= a and b;
    layer5_outputs(1579) <= b and not a;
    layer5_outputs(1580) <= a and not b;
    layer5_outputs(1581) <= not (a or b);
    layer5_outputs(1582) <= not (a and b);
    layer5_outputs(1583) <= '1';
    layer5_outputs(1584) <= a or b;
    layer5_outputs(1585) <= not (a xor b);
    layer5_outputs(1586) <= a;
    layer5_outputs(1587) <= not b or a;
    layer5_outputs(1588) <= b;
    layer5_outputs(1589) <= not b;
    layer5_outputs(1590) <= b;
    layer5_outputs(1591) <= a or b;
    layer5_outputs(1592) <= a;
    layer5_outputs(1593) <= '0';
    layer5_outputs(1594) <= not a or b;
    layer5_outputs(1595) <= a and not b;
    layer5_outputs(1596) <= a and b;
    layer5_outputs(1597) <= a and b;
    layer5_outputs(1598) <= b;
    layer5_outputs(1599) <= b;
    layer5_outputs(1600) <= a or b;
    layer5_outputs(1601) <= not a;
    layer5_outputs(1602) <= a and b;
    layer5_outputs(1603) <= '0';
    layer5_outputs(1604) <= not a;
    layer5_outputs(1605) <= a or b;
    layer5_outputs(1606) <= not a;
    layer5_outputs(1607) <= not a;
    layer5_outputs(1608) <= not b or a;
    layer5_outputs(1609) <= '0';
    layer5_outputs(1610) <= a xor b;
    layer5_outputs(1611) <= a xor b;
    layer5_outputs(1612) <= a and not b;
    layer5_outputs(1613) <= not b;
    layer5_outputs(1614) <= not a;
    layer5_outputs(1615) <= b and not a;
    layer5_outputs(1616) <= not (a xor b);
    layer5_outputs(1617) <= b;
    layer5_outputs(1618) <= not a;
    layer5_outputs(1619) <= b and not a;
    layer5_outputs(1620) <= not b or a;
    layer5_outputs(1621) <= b and not a;
    layer5_outputs(1622) <= not (a and b);
    layer5_outputs(1623) <= not (a or b);
    layer5_outputs(1624) <= a;
    layer5_outputs(1625) <= not (a and b);
    layer5_outputs(1626) <= '1';
    layer5_outputs(1627) <= not a;
    layer5_outputs(1628) <= not (a xor b);
    layer5_outputs(1629) <= not (a xor b);
    layer5_outputs(1630) <= not a;
    layer5_outputs(1631) <= a;
    layer5_outputs(1632) <= a;
    layer5_outputs(1633) <= not a or b;
    layer5_outputs(1634) <= b and not a;
    layer5_outputs(1635) <= '1';
    layer5_outputs(1636) <= not b or a;
    layer5_outputs(1637) <= not a;
    layer5_outputs(1638) <= not (a or b);
    layer5_outputs(1639) <= not b;
    layer5_outputs(1640) <= not (a and b);
    layer5_outputs(1641) <= not b or a;
    layer5_outputs(1642) <= b and not a;
    layer5_outputs(1643) <= a;
    layer5_outputs(1644) <= a or b;
    layer5_outputs(1645) <= b;
    layer5_outputs(1646) <= a and b;
    layer5_outputs(1647) <= a;
    layer5_outputs(1648) <= a or b;
    layer5_outputs(1649) <= a;
    layer5_outputs(1650) <= a;
    layer5_outputs(1651) <= a;
    layer5_outputs(1652) <= not b;
    layer5_outputs(1653) <= not a;
    layer5_outputs(1654) <= a or b;
    layer5_outputs(1655) <= a;
    layer5_outputs(1656) <= b;
    layer5_outputs(1657) <= not (a xor b);
    layer5_outputs(1658) <= b and not a;
    layer5_outputs(1659) <= not (a and b);
    layer5_outputs(1660) <= '0';
    layer5_outputs(1661) <= not a;
    layer5_outputs(1662) <= b;
    layer5_outputs(1663) <= not a or b;
    layer5_outputs(1664) <= not b;
    layer5_outputs(1665) <= a or b;
    layer5_outputs(1666) <= a and b;
    layer5_outputs(1667) <= not (a or b);
    layer5_outputs(1668) <= a xor b;
    layer5_outputs(1669) <= '0';
    layer5_outputs(1670) <= b;
    layer5_outputs(1671) <= b;
    layer5_outputs(1672) <= a;
    layer5_outputs(1673) <= not (a and b);
    layer5_outputs(1674) <= a;
    layer5_outputs(1675) <= not a;
    layer5_outputs(1676) <= a and b;
    layer5_outputs(1677) <= not a;
    layer5_outputs(1678) <= a and b;
    layer5_outputs(1679) <= a and b;
    layer5_outputs(1680) <= b and not a;
    layer5_outputs(1681) <= a;
    layer5_outputs(1682) <= not a;
    layer5_outputs(1683) <= not a or b;
    layer5_outputs(1684) <= not b;
    layer5_outputs(1685) <= not a or b;
    layer5_outputs(1686) <= not a;
    layer5_outputs(1687) <= a xor b;
    layer5_outputs(1688) <= not a;
    layer5_outputs(1689) <= not b or a;
    layer5_outputs(1690) <= not b;
    layer5_outputs(1691) <= not b;
    layer5_outputs(1692) <= not b or a;
    layer5_outputs(1693) <= not b;
    layer5_outputs(1694) <= not a or b;
    layer5_outputs(1695) <= a;
    layer5_outputs(1696) <= a xor b;
    layer5_outputs(1697) <= '1';
    layer5_outputs(1698) <= not a or b;
    layer5_outputs(1699) <= not a;
    layer5_outputs(1700) <= not (a or b);
    layer5_outputs(1701) <= b and not a;
    layer5_outputs(1702) <= not (a or b);
    layer5_outputs(1703) <= b;
    layer5_outputs(1704) <= not b or a;
    layer5_outputs(1705) <= '0';
    layer5_outputs(1706) <= a and not b;
    layer5_outputs(1707) <= a and not b;
    layer5_outputs(1708) <= not b;
    layer5_outputs(1709) <= not a;
    layer5_outputs(1710) <= '1';
    layer5_outputs(1711) <= not a;
    layer5_outputs(1712) <= not (a and b);
    layer5_outputs(1713) <= not a;
    layer5_outputs(1714) <= a;
    layer5_outputs(1715) <= not b;
    layer5_outputs(1716) <= not (a or b);
    layer5_outputs(1717) <= a;
    layer5_outputs(1718) <= not a or b;
    layer5_outputs(1719) <= not a;
    layer5_outputs(1720) <= not b or a;
    layer5_outputs(1721) <= not b or a;
    layer5_outputs(1722) <= not (a and b);
    layer5_outputs(1723) <= a xor b;
    layer5_outputs(1724) <= a;
    layer5_outputs(1725) <= a;
    layer5_outputs(1726) <= not a or b;
    layer5_outputs(1727) <= a xor b;
    layer5_outputs(1728) <= a;
    layer5_outputs(1729) <= not (a or b);
    layer5_outputs(1730) <= a;
    layer5_outputs(1731) <= a or b;
    layer5_outputs(1732) <= not a;
    layer5_outputs(1733) <= a and not b;
    layer5_outputs(1734) <= not (a and b);
    layer5_outputs(1735) <= b;
    layer5_outputs(1736) <= '0';
    layer5_outputs(1737) <= b;
    layer5_outputs(1738) <= not (a and b);
    layer5_outputs(1739) <= not b or a;
    layer5_outputs(1740) <= not (a or b);
    layer5_outputs(1741) <= a and b;
    layer5_outputs(1742) <= '0';
    layer5_outputs(1743) <= not (a and b);
    layer5_outputs(1744) <= not b or a;
    layer5_outputs(1745) <= a xor b;
    layer5_outputs(1746) <= a;
    layer5_outputs(1747) <= b and not a;
    layer5_outputs(1748) <= a and not b;
    layer5_outputs(1749) <= a and b;
    layer5_outputs(1750) <= not b or a;
    layer5_outputs(1751) <= '0';
    layer5_outputs(1752) <= a and not b;
    layer5_outputs(1753) <= not (a and b);
    layer5_outputs(1754) <= not a or b;
    layer5_outputs(1755) <= a xor b;
    layer5_outputs(1756) <= not a;
    layer5_outputs(1757) <= b;
    layer5_outputs(1758) <= b;
    layer5_outputs(1759) <= not a;
    layer5_outputs(1760) <= not (a or b);
    layer5_outputs(1761) <= not a or b;
    layer5_outputs(1762) <= not b;
    layer5_outputs(1763) <= not a;
    layer5_outputs(1764) <= not a;
    layer5_outputs(1765) <= a;
    layer5_outputs(1766) <= not a;
    layer5_outputs(1767) <= a and not b;
    layer5_outputs(1768) <= a and not b;
    layer5_outputs(1769) <= not a or b;
    layer5_outputs(1770) <= not b;
    layer5_outputs(1771) <= a and b;
    layer5_outputs(1772) <= a and b;
    layer5_outputs(1773) <= b;
    layer5_outputs(1774) <= b;
    layer5_outputs(1775) <= not (a and b);
    layer5_outputs(1776) <= b;
    layer5_outputs(1777) <= a xor b;
    layer5_outputs(1778) <= '1';
    layer5_outputs(1779) <= not (a or b);
    layer5_outputs(1780) <= not (a or b);
    layer5_outputs(1781) <= not b;
    layer5_outputs(1782) <= not b;
    layer5_outputs(1783) <= not (a xor b);
    layer5_outputs(1784) <= '0';
    layer5_outputs(1785) <= not b or a;
    layer5_outputs(1786) <= b;
    layer5_outputs(1787) <= not b or a;
    layer5_outputs(1788) <= a and not b;
    layer5_outputs(1789) <= a xor b;
    layer5_outputs(1790) <= not a;
    layer5_outputs(1791) <= not b;
    layer5_outputs(1792) <= a and b;
    layer5_outputs(1793) <= a and b;
    layer5_outputs(1794) <= not b;
    layer5_outputs(1795) <= a or b;
    layer5_outputs(1796) <= a and not b;
    layer5_outputs(1797) <= not (a or b);
    layer5_outputs(1798) <= b;
    layer5_outputs(1799) <= not b;
    layer5_outputs(1800) <= not b;
    layer5_outputs(1801) <= not b or a;
    layer5_outputs(1802) <= a;
    layer5_outputs(1803) <= not b;
    layer5_outputs(1804) <= not (a and b);
    layer5_outputs(1805) <= not a;
    layer5_outputs(1806) <= not (a or b);
    layer5_outputs(1807) <= b;
    layer5_outputs(1808) <= not a or b;
    layer5_outputs(1809) <= b;
    layer5_outputs(1810) <= b;
    layer5_outputs(1811) <= a;
    layer5_outputs(1812) <= b;
    layer5_outputs(1813) <= a xor b;
    layer5_outputs(1814) <= not b;
    layer5_outputs(1815) <= not (a or b);
    layer5_outputs(1816) <= a and not b;
    layer5_outputs(1817) <= a;
    layer5_outputs(1818) <= a;
    layer5_outputs(1819) <= not b;
    layer5_outputs(1820) <= not (a or b);
    layer5_outputs(1821) <= b;
    layer5_outputs(1822) <= a;
    layer5_outputs(1823) <= b;
    layer5_outputs(1824) <= not (a or b);
    layer5_outputs(1825) <= not a;
    layer5_outputs(1826) <= b;
    layer5_outputs(1827) <= a and b;
    layer5_outputs(1828) <= not a or b;
    layer5_outputs(1829) <= not a or b;
    layer5_outputs(1830) <= not (a or b);
    layer5_outputs(1831) <= not (a and b);
    layer5_outputs(1832) <= b and not a;
    layer5_outputs(1833) <= b and not a;
    layer5_outputs(1834) <= a;
    layer5_outputs(1835) <= a xor b;
    layer5_outputs(1836) <= not a or b;
    layer5_outputs(1837) <= b;
    layer5_outputs(1838) <= '0';
    layer5_outputs(1839) <= not (a and b);
    layer5_outputs(1840) <= not (a or b);
    layer5_outputs(1841) <= not a;
    layer5_outputs(1842) <= a;
    layer5_outputs(1843) <= b;
    layer5_outputs(1844) <= not (a or b);
    layer5_outputs(1845) <= b;
    layer5_outputs(1846) <= a and not b;
    layer5_outputs(1847) <= not a;
    layer5_outputs(1848) <= '0';
    layer5_outputs(1849) <= not a;
    layer5_outputs(1850) <= not a or b;
    layer5_outputs(1851) <= '1';
    layer5_outputs(1852) <= not b;
    layer5_outputs(1853) <= not a or b;
    layer5_outputs(1854) <= b;
    layer5_outputs(1855) <= b;
    layer5_outputs(1856) <= '1';
    layer5_outputs(1857) <= not a;
    layer5_outputs(1858) <= '1';
    layer5_outputs(1859) <= a and not b;
    layer5_outputs(1860) <= a and not b;
    layer5_outputs(1861) <= not (a xor b);
    layer5_outputs(1862) <= a and b;
    layer5_outputs(1863) <= not a;
    layer5_outputs(1864) <= b and not a;
    layer5_outputs(1865) <= a;
    layer5_outputs(1866) <= a or b;
    layer5_outputs(1867) <= not b;
    layer5_outputs(1868) <= b;
    layer5_outputs(1869) <= a and b;
    layer5_outputs(1870) <= not a;
    layer5_outputs(1871) <= not a;
    layer5_outputs(1872) <= b and not a;
    layer5_outputs(1873) <= not b;
    layer5_outputs(1874) <= not a;
    layer5_outputs(1875) <= a and b;
    layer5_outputs(1876) <= a and not b;
    layer5_outputs(1877) <= a xor b;
    layer5_outputs(1878) <= not b;
    layer5_outputs(1879) <= a and b;
    layer5_outputs(1880) <= a or b;
    layer5_outputs(1881) <= a and b;
    layer5_outputs(1882) <= '1';
    layer5_outputs(1883) <= b and not a;
    layer5_outputs(1884) <= '0';
    layer5_outputs(1885) <= not (a or b);
    layer5_outputs(1886) <= not b;
    layer5_outputs(1887) <= '1';
    layer5_outputs(1888) <= not a or b;
    layer5_outputs(1889) <= not b or a;
    layer5_outputs(1890) <= not a or b;
    layer5_outputs(1891) <= a or b;
    layer5_outputs(1892) <= b;
    layer5_outputs(1893) <= not b or a;
    layer5_outputs(1894) <= not (a and b);
    layer5_outputs(1895) <= not (a or b);
    layer5_outputs(1896) <= not b or a;
    layer5_outputs(1897) <= b;
    layer5_outputs(1898) <= not (a and b);
    layer5_outputs(1899) <= '0';
    layer5_outputs(1900) <= a or b;
    layer5_outputs(1901) <= a and not b;
    layer5_outputs(1902) <= a and not b;
    layer5_outputs(1903) <= '0';
    layer5_outputs(1904) <= not (a or b);
    layer5_outputs(1905) <= not a or b;
    layer5_outputs(1906) <= a and b;
    layer5_outputs(1907) <= b;
    layer5_outputs(1908) <= a and b;
    layer5_outputs(1909) <= b and not a;
    layer5_outputs(1910) <= a xor b;
    layer5_outputs(1911) <= not a or b;
    layer5_outputs(1912) <= a and b;
    layer5_outputs(1913) <= not a;
    layer5_outputs(1914) <= not (a or b);
    layer5_outputs(1915) <= not a or b;
    layer5_outputs(1916) <= a and b;
    layer5_outputs(1917) <= not a or b;
    layer5_outputs(1918) <= not b;
    layer5_outputs(1919) <= a and not b;
    layer5_outputs(1920) <= '0';
    layer5_outputs(1921) <= not (a or b);
    layer5_outputs(1922) <= a;
    layer5_outputs(1923) <= a xor b;
    layer5_outputs(1924) <= not a;
    layer5_outputs(1925) <= a and not b;
    layer5_outputs(1926) <= not a;
    layer5_outputs(1927) <= a and not b;
    layer5_outputs(1928) <= a or b;
    layer5_outputs(1929) <= not a;
    layer5_outputs(1930) <= a;
    layer5_outputs(1931) <= not (a and b);
    layer5_outputs(1932) <= not (a and b);
    layer5_outputs(1933) <= b;
    layer5_outputs(1934) <= b and not a;
    layer5_outputs(1935) <= not (a and b);
    layer5_outputs(1936) <= not (a and b);
    layer5_outputs(1937) <= not b;
    layer5_outputs(1938) <= a xor b;
    layer5_outputs(1939) <= b;
    layer5_outputs(1940) <= b;
    layer5_outputs(1941) <= not b;
    layer5_outputs(1942) <= a and not b;
    layer5_outputs(1943) <= not a;
    layer5_outputs(1944) <= a and b;
    layer5_outputs(1945) <= b and not a;
    layer5_outputs(1946) <= a and b;
    layer5_outputs(1947) <= not a;
    layer5_outputs(1948) <= a;
    layer5_outputs(1949) <= '0';
    layer5_outputs(1950) <= not b or a;
    layer5_outputs(1951) <= not (a or b);
    layer5_outputs(1952) <= b;
    layer5_outputs(1953) <= b and not a;
    layer5_outputs(1954) <= '1';
    layer5_outputs(1955) <= not a;
    layer5_outputs(1956) <= a xor b;
    layer5_outputs(1957) <= not (a or b);
    layer5_outputs(1958) <= a and not b;
    layer5_outputs(1959) <= a;
    layer5_outputs(1960) <= not b;
    layer5_outputs(1961) <= a;
    layer5_outputs(1962) <= a and b;
    layer5_outputs(1963) <= b;
    layer5_outputs(1964) <= a and not b;
    layer5_outputs(1965) <= not b;
    layer5_outputs(1966) <= a and not b;
    layer5_outputs(1967) <= not (a and b);
    layer5_outputs(1968) <= '1';
    layer5_outputs(1969) <= '1';
    layer5_outputs(1970) <= not a;
    layer5_outputs(1971) <= not a;
    layer5_outputs(1972) <= not (a xor b);
    layer5_outputs(1973) <= not (a or b);
    layer5_outputs(1974) <= a or b;
    layer5_outputs(1975) <= not (a or b);
    layer5_outputs(1976) <= a and not b;
    layer5_outputs(1977) <= a and b;
    layer5_outputs(1978) <= not a or b;
    layer5_outputs(1979) <= a;
    layer5_outputs(1980) <= not b;
    layer5_outputs(1981) <= a and b;
    layer5_outputs(1982) <= not a;
    layer5_outputs(1983) <= a and b;
    layer5_outputs(1984) <= not (a or b);
    layer5_outputs(1985) <= a or b;
    layer5_outputs(1986) <= '0';
    layer5_outputs(1987) <= a and b;
    layer5_outputs(1988) <= not b;
    layer5_outputs(1989) <= not (a and b);
    layer5_outputs(1990) <= not (a or b);
    layer5_outputs(1991) <= a and b;
    layer5_outputs(1992) <= a and not b;
    layer5_outputs(1993) <= a xor b;
    layer5_outputs(1994) <= not (a and b);
    layer5_outputs(1995) <= not b or a;
    layer5_outputs(1996) <= a and b;
    layer5_outputs(1997) <= not b;
    layer5_outputs(1998) <= a;
    layer5_outputs(1999) <= not a or b;
    layer5_outputs(2000) <= b;
    layer5_outputs(2001) <= '0';
    layer5_outputs(2002) <= not b;
    layer5_outputs(2003) <= not (a and b);
    layer5_outputs(2004) <= not (a and b);
    layer5_outputs(2005) <= '1';
    layer5_outputs(2006) <= '1';
    layer5_outputs(2007) <= b;
    layer5_outputs(2008) <= a;
    layer5_outputs(2009) <= a and b;
    layer5_outputs(2010) <= not a;
    layer5_outputs(2011) <= not b;
    layer5_outputs(2012) <= b;
    layer5_outputs(2013) <= not a;
    layer5_outputs(2014) <= not (a and b);
    layer5_outputs(2015) <= '1';
    layer5_outputs(2016) <= not b or a;
    layer5_outputs(2017) <= b;
    layer5_outputs(2018) <= not (a and b);
    layer5_outputs(2019) <= not b or a;
    layer5_outputs(2020) <= not (a or b);
    layer5_outputs(2021) <= not (a xor b);
    layer5_outputs(2022) <= not b or a;
    layer5_outputs(2023) <= a and b;
    layer5_outputs(2024) <= not b or a;
    layer5_outputs(2025) <= a and not b;
    layer5_outputs(2026) <= '1';
    layer5_outputs(2027) <= not b;
    layer5_outputs(2028) <= not a;
    layer5_outputs(2029) <= a xor b;
    layer5_outputs(2030) <= not a;
    layer5_outputs(2031) <= '1';
    layer5_outputs(2032) <= not b;
    layer5_outputs(2033) <= not a or b;
    layer5_outputs(2034) <= b;
    layer5_outputs(2035) <= not b or a;
    layer5_outputs(2036) <= not b or a;
    layer5_outputs(2037) <= a xor b;
    layer5_outputs(2038) <= '1';
    layer5_outputs(2039) <= b and not a;
    layer5_outputs(2040) <= a;
    layer5_outputs(2041) <= a xor b;
    layer5_outputs(2042) <= a;
    layer5_outputs(2043) <= not (a xor b);
    layer5_outputs(2044) <= a and not b;
    layer5_outputs(2045) <= a and not b;
    layer5_outputs(2046) <= a;
    layer5_outputs(2047) <= not (a and b);
    layer5_outputs(2048) <= not (a and b);
    layer5_outputs(2049) <= b;
    layer5_outputs(2050) <= not a;
    layer5_outputs(2051) <= a and not b;
    layer5_outputs(2052) <= '1';
    layer5_outputs(2053) <= not b;
    layer5_outputs(2054) <= not a;
    layer5_outputs(2055) <= a xor b;
    layer5_outputs(2056) <= not a;
    layer5_outputs(2057) <= a or b;
    layer5_outputs(2058) <= a or b;
    layer5_outputs(2059) <= not (a or b);
    layer5_outputs(2060) <= not (a and b);
    layer5_outputs(2061) <= not a or b;
    layer5_outputs(2062) <= not b;
    layer5_outputs(2063) <= a or b;
    layer5_outputs(2064) <= '0';
    layer5_outputs(2065) <= a xor b;
    layer5_outputs(2066) <= b and not a;
    layer5_outputs(2067) <= not (a and b);
    layer5_outputs(2068) <= b;
    layer5_outputs(2069) <= not a or b;
    layer5_outputs(2070) <= b and not a;
    layer5_outputs(2071) <= not (a and b);
    layer5_outputs(2072) <= not a;
    layer5_outputs(2073) <= not b;
    layer5_outputs(2074) <= '0';
    layer5_outputs(2075) <= a or b;
    layer5_outputs(2076) <= not (a or b);
    layer5_outputs(2077) <= b and not a;
    layer5_outputs(2078) <= not (a or b);
    layer5_outputs(2079) <= b;
    layer5_outputs(2080) <= not (a or b);
    layer5_outputs(2081) <= not a;
    layer5_outputs(2082) <= '0';
    layer5_outputs(2083) <= not a or b;
    layer5_outputs(2084) <= a or b;
    layer5_outputs(2085) <= not (a and b);
    layer5_outputs(2086) <= not a;
    layer5_outputs(2087) <= '1';
    layer5_outputs(2088) <= a or b;
    layer5_outputs(2089) <= a and b;
    layer5_outputs(2090) <= '0';
    layer5_outputs(2091) <= not b;
    layer5_outputs(2092) <= a;
    layer5_outputs(2093) <= not (a xor b);
    layer5_outputs(2094) <= a;
    layer5_outputs(2095) <= '0';
    layer5_outputs(2096) <= not (a and b);
    layer5_outputs(2097) <= a and b;
    layer5_outputs(2098) <= not a;
    layer5_outputs(2099) <= not b or a;
    layer5_outputs(2100) <= b;
    layer5_outputs(2101) <= b;
    layer5_outputs(2102) <= not a or b;
    layer5_outputs(2103) <= a xor b;
    layer5_outputs(2104) <= a;
    layer5_outputs(2105) <= a or b;
    layer5_outputs(2106) <= b;
    layer5_outputs(2107) <= b and not a;
    layer5_outputs(2108) <= not b or a;
    layer5_outputs(2109) <= not b;
    layer5_outputs(2110) <= a;
    layer5_outputs(2111) <= not a or b;
    layer5_outputs(2112) <= b and not a;
    layer5_outputs(2113) <= b and not a;
    layer5_outputs(2114) <= not (a xor b);
    layer5_outputs(2115) <= a and not b;
    layer5_outputs(2116) <= not (a xor b);
    layer5_outputs(2117) <= not (a and b);
    layer5_outputs(2118) <= not (a or b);
    layer5_outputs(2119) <= not b;
    layer5_outputs(2120) <= '0';
    layer5_outputs(2121) <= not b;
    layer5_outputs(2122) <= not a or b;
    layer5_outputs(2123) <= a and b;
    layer5_outputs(2124) <= not b or a;
    layer5_outputs(2125) <= not (a and b);
    layer5_outputs(2126) <= not (a and b);
    layer5_outputs(2127) <= a;
    layer5_outputs(2128) <= not a or b;
    layer5_outputs(2129) <= b;
    layer5_outputs(2130) <= b;
    layer5_outputs(2131) <= not (a and b);
    layer5_outputs(2132) <= b;
    layer5_outputs(2133) <= not (a and b);
    layer5_outputs(2134) <= not (a and b);
    layer5_outputs(2135) <= not b or a;
    layer5_outputs(2136) <= not (a xor b);
    layer5_outputs(2137) <= not a;
    layer5_outputs(2138) <= not (a or b);
    layer5_outputs(2139) <= not (a or b);
    layer5_outputs(2140) <= a;
    layer5_outputs(2141) <= not a or b;
    layer5_outputs(2142) <= not (a or b);
    layer5_outputs(2143) <= not b or a;
    layer5_outputs(2144) <= a;
    layer5_outputs(2145) <= a xor b;
    layer5_outputs(2146) <= not b;
    layer5_outputs(2147) <= b and not a;
    layer5_outputs(2148) <= a xor b;
    layer5_outputs(2149) <= '1';
    layer5_outputs(2150) <= not (a and b);
    layer5_outputs(2151) <= a and b;
    layer5_outputs(2152) <= not (a or b);
    layer5_outputs(2153) <= b and not a;
    layer5_outputs(2154) <= not a;
    layer5_outputs(2155) <= not (a or b);
    layer5_outputs(2156) <= not b;
    layer5_outputs(2157) <= a and b;
    layer5_outputs(2158) <= a;
    layer5_outputs(2159) <= not b;
    layer5_outputs(2160) <= a;
    layer5_outputs(2161) <= a xor b;
    layer5_outputs(2162) <= not b or a;
    layer5_outputs(2163) <= not (a or b);
    layer5_outputs(2164) <= a or b;
    layer5_outputs(2165) <= not b or a;
    layer5_outputs(2166) <= not b;
    layer5_outputs(2167) <= not a or b;
    layer5_outputs(2168) <= not (a or b);
    layer5_outputs(2169) <= b;
    layer5_outputs(2170) <= '1';
    layer5_outputs(2171) <= not a;
    layer5_outputs(2172) <= a;
    layer5_outputs(2173) <= a xor b;
    layer5_outputs(2174) <= not a;
    layer5_outputs(2175) <= b;
    layer5_outputs(2176) <= not a;
    layer5_outputs(2177) <= not (a or b);
    layer5_outputs(2178) <= not b;
    layer5_outputs(2179) <= a xor b;
    layer5_outputs(2180) <= b;
    layer5_outputs(2181) <= not (a and b);
    layer5_outputs(2182) <= '0';
    layer5_outputs(2183) <= not a;
    layer5_outputs(2184) <= not a;
    layer5_outputs(2185) <= a and b;
    layer5_outputs(2186) <= a xor b;
    layer5_outputs(2187) <= a and not b;
    layer5_outputs(2188) <= a or b;
    layer5_outputs(2189) <= b and not a;
    layer5_outputs(2190) <= a or b;
    layer5_outputs(2191) <= not a;
    layer5_outputs(2192) <= not b;
    layer5_outputs(2193) <= a or b;
    layer5_outputs(2194) <= b and not a;
    layer5_outputs(2195) <= a or b;
    layer5_outputs(2196) <= b and not a;
    layer5_outputs(2197) <= a and b;
    layer5_outputs(2198) <= not (a or b);
    layer5_outputs(2199) <= not (a xor b);
    layer5_outputs(2200) <= a and b;
    layer5_outputs(2201) <= a xor b;
    layer5_outputs(2202) <= not a;
    layer5_outputs(2203) <= '1';
    layer5_outputs(2204) <= not b;
    layer5_outputs(2205) <= not b;
    layer5_outputs(2206) <= not (a xor b);
    layer5_outputs(2207) <= a;
    layer5_outputs(2208) <= a xor b;
    layer5_outputs(2209) <= b and not a;
    layer5_outputs(2210) <= not b;
    layer5_outputs(2211) <= b and not a;
    layer5_outputs(2212) <= a and not b;
    layer5_outputs(2213) <= b;
    layer5_outputs(2214) <= not (a or b);
    layer5_outputs(2215) <= not (a or b);
    layer5_outputs(2216) <= a xor b;
    layer5_outputs(2217) <= not a or b;
    layer5_outputs(2218) <= b and not a;
    layer5_outputs(2219) <= a xor b;
    layer5_outputs(2220) <= not a;
    layer5_outputs(2221) <= not b or a;
    layer5_outputs(2222) <= b and not a;
    layer5_outputs(2223) <= b and not a;
    layer5_outputs(2224) <= a and b;
    layer5_outputs(2225) <= '0';
    layer5_outputs(2226) <= b;
    layer5_outputs(2227) <= not a or b;
    layer5_outputs(2228) <= a xor b;
    layer5_outputs(2229) <= not (a xor b);
    layer5_outputs(2230) <= not a;
    layer5_outputs(2231) <= not a or b;
    layer5_outputs(2232) <= not b or a;
    layer5_outputs(2233) <= not a or b;
    layer5_outputs(2234) <= not b or a;
    layer5_outputs(2235) <= a;
    layer5_outputs(2236) <= not (a and b);
    layer5_outputs(2237) <= a or b;
    layer5_outputs(2238) <= not b or a;
    layer5_outputs(2239) <= not a or b;
    layer5_outputs(2240) <= not (a and b);
    layer5_outputs(2241) <= not b or a;
    layer5_outputs(2242) <= not a or b;
    layer5_outputs(2243) <= a xor b;
    layer5_outputs(2244) <= '0';
    layer5_outputs(2245) <= a;
    layer5_outputs(2246) <= not b;
    layer5_outputs(2247) <= not (a xor b);
    layer5_outputs(2248) <= a and b;
    layer5_outputs(2249) <= not b;
    layer5_outputs(2250) <= a or b;
    layer5_outputs(2251) <= b;
    layer5_outputs(2252) <= b;
    layer5_outputs(2253) <= a and not b;
    layer5_outputs(2254) <= b;
    layer5_outputs(2255) <= not b;
    layer5_outputs(2256) <= b;
    layer5_outputs(2257) <= not (a xor b);
    layer5_outputs(2258) <= not b;
    layer5_outputs(2259) <= not b;
    layer5_outputs(2260) <= b and not a;
    layer5_outputs(2261) <= a and b;
    layer5_outputs(2262) <= '1';
    layer5_outputs(2263) <= not a;
    layer5_outputs(2264) <= a and b;
    layer5_outputs(2265) <= not (a xor b);
    layer5_outputs(2266) <= a;
    layer5_outputs(2267) <= not (a and b);
    layer5_outputs(2268) <= not (a xor b);
    layer5_outputs(2269) <= not (a xor b);
    layer5_outputs(2270) <= b and not a;
    layer5_outputs(2271) <= not (a and b);
    layer5_outputs(2272) <= not b or a;
    layer5_outputs(2273) <= b;
    layer5_outputs(2274) <= not (a or b);
    layer5_outputs(2275) <= not a or b;
    layer5_outputs(2276) <= not b;
    layer5_outputs(2277) <= b and not a;
    layer5_outputs(2278) <= not b or a;
    layer5_outputs(2279) <= b;
    layer5_outputs(2280) <= a;
    layer5_outputs(2281) <= a;
    layer5_outputs(2282) <= a;
    layer5_outputs(2283) <= '0';
    layer5_outputs(2284) <= a xor b;
    layer5_outputs(2285) <= not (a and b);
    layer5_outputs(2286) <= not a or b;
    layer5_outputs(2287) <= '1';
    layer5_outputs(2288) <= not (a and b);
    layer5_outputs(2289) <= not a or b;
    layer5_outputs(2290) <= not (a or b);
    layer5_outputs(2291) <= not a or b;
    layer5_outputs(2292) <= b and not a;
    layer5_outputs(2293) <= '0';
    layer5_outputs(2294) <= a;
    layer5_outputs(2295) <= b and not a;
    layer5_outputs(2296) <= not a;
    layer5_outputs(2297) <= not a;
    layer5_outputs(2298) <= a;
    layer5_outputs(2299) <= a xor b;
    layer5_outputs(2300) <= a and b;
    layer5_outputs(2301) <= b;
    layer5_outputs(2302) <= a or b;
    layer5_outputs(2303) <= a;
    layer5_outputs(2304) <= not b;
    layer5_outputs(2305) <= not a;
    layer5_outputs(2306) <= a or b;
    layer5_outputs(2307) <= not a or b;
    layer5_outputs(2308) <= b;
    layer5_outputs(2309) <= a or b;
    layer5_outputs(2310) <= b;
    layer5_outputs(2311) <= a or b;
    layer5_outputs(2312) <= not a;
    layer5_outputs(2313) <= not a;
    layer5_outputs(2314) <= b and not a;
    layer5_outputs(2315) <= not a or b;
    layer5_outputs(2316) <= a and not b;
    layer5_outputs(2317) <= not a;
    layer5_outputs(2318) <= a;
    layer5_outputs(2319) <= not a or b;
    layer5_outputs(2320) <= b;
    layer5_outputs(2321) <= '1';
    layer5_outputs(2322) <= not (a or b);
    layer5_outputs(2323) <= '1';
    layer5_outputs(2324) <= a;
    layer5_outputs(2325) <= not a or b;
    layer5_outputs(2326) <= not (a or b);
    layer5_outputs(2327) <= not (a and b);
    layer5_outputs(2328) <= not a;
    layer5_outputs(2329) <= not a;
    layer5_outputs(2330) <= not (a xor b);
    layer5_outputs(2331) <= a and b;
    layer5_outputs(2332) <= not b;
    layer5_outputs(2333) <= a or b;
    layer5_outputs(2334) <= not (a and b);
    layer5_outputs(2335) <= a xor b;
    layer5_outputs(2336) <= not b or a;
    layer5_outputs(2337) <= not a;
    layer5_outputs(2338) <= '0';
    layer5_outputs(2339) <= a or b;
    layer5_outputs(2340) <= a and b;
    layer5_outputs(2341) <= '0';
    layer5_outputs(2342) <= a and not b;
    layer5_outputs(2343) <= not b or a;
    layer5_outputs(2344) <= not a;
    layer5_outputs(2345) <= a;
    layer5_outputs(2346) <= b;
    layer5_outputs(2347) <= a or b;
    layer5_outputs(2348) <= b and not a;
    layer5_outputs(2349) <= b;
    layer5_outputs(2350) <= not b;
    layer5_outputs(2351) <= a and b;
    layer5_outputs(2352) <= b and not a;
    layer5_outputs(2353) <= not (a xor b);
    layer5_outputs(2354) <= a;
    layer5_outputs(2355) <= not (a or b);
    layer5_outputs(2356) <= a and b;
    layer5_outputs(2357) <= not a;
    layer5_outputs(2358) <= not (a or b);
    layer5_outputs(2359) <= not a;
    layer5_outputs(2360) <= not b;
    layer5_outputs(2361) <= not a or b;
    layer5_outputs(2362) <= a and not b;
    layer5_outputs(2363) <= not (a and b);
    layer5_outputs(2364) <= b;
    layer5_outputs(2365) <= not b;
    layer5_outputs(2366) <= '0';
    layer5_outputs(2367) <= not a or b;
    layer5_outputs(2368) <= a;
    layer5_outputs(2369) <= a and not b;
    layer5_outputs(2370) <= not a or b;
    layer5_outputs(2371) <= not (a and b);
    layer5_outputs(2372) <= a;
    layer5_outputs(2373) <= a xor b;
    layer5_outputs(2374) <= not b or a;
    layer5_outputs(2375) <= b;
    layer5_outputs(2376) <= not b;
    layer5_outputs(2377) <= not a;
    layer5_outputs(2378) <= a;
    layer5_outputs(2379) <= b;
    layer5_outputs(2380) <= not a or b;
    layer5_outputs(2381) <= not b or a;
    layer5_outputs(2382) <= a and not b;
    layer5_outputs(2383) <= not (a xor b);
    layer5_outputs(2384) <= not a;
    layer5_outputs(2385) <= not b or a;
    layer5_outputs(2386) <= b and not a;
    layer5_outputs(2387) <= not a;
    layer5_outputs(2388) <= a or b;
    layer5_outputs(2389) <= not a or b;
    layer5_outputs(2390) <= a and b;
    layer5_outputs(2391) <= not (a and b);
    layer5_outputs(2392) <= not (a or b);
    layer5_outputs(2393) <= a or b;
    layer5_outputs(2394) <= '0';
    layer5_outputs(2395) <= not (a xor b);
    layer5_outputs(2396) <= not (a xor b);
    layer5_outputs(2397) <= not a;
    layer5_outputs(2398) <= '0';
    layer5_outputs(2399) <= not b;
    layer5_outputs(2400) <= a or b;
    layer5_outputs(2401) <= not b or a;
    layer5_outputs(2402) <= a;
    layer5_outputs(2403) <= b and not a;
    layer5_outputs(2404) <= a;
    layer5_outputs(2405) <= not b or a;
    layer5_outputs(2406) <= a and b;
    layer5_outputs(2407) <= not (a or b);
    layer5_outputs(2408) <= not b or a;
    layer5_outputs(2409) <= not b;
    layer5_outputs(2410) <= b and not a;
    layer5_outputs(2411) <= a and not b;
    layer5_outputs(2412) <= a and b;
    layer5_outputs(2413) <= a or b;
    layer5_outputs(2414) <= not (a or b);
    layer5_outputs(2415) <= not a or b;
    layer5_outputs(2416) <= not (a or b);
    layer5_outputs(2417) <= not b;
    layer5_outputs(2418) <= b;
    layer5_outputs(2419) <= '1';
    layer5_outputs(2420) <= a xor b;
    layer5_outputs(2421) <= b;
    layer5_outputs(2422) <= a and not b;
    layer5_outputs(2423) <= a xor b;
    layer5_outputs(2424) <= not b;
    layer5_outputs(2425) <= not a or b;
    layer5_outputs(2426) <= b;
    layer5_outputs(2427) <= not a or b;
    layer5_outputs(2428) <= a or b;
    layer5_outputs(2429) <= '1';
    layer5_outputs(2430) <= '1';
    layer5_outputs(2431) <= not (a and b);
    layer5_outputs(2432) <= not (a or b);
    layer5_outputs(2433) <= '0';
    layer5_outputs(2434) <= b;
    layer5_outputs(2435) <= not (a or b);
    layer5_outputs(2436) <= '1';
    layer5_outputs(2437) <= a or b;
    layer5_outputs(2438) <= not b;
    layer5_outputs(2439) <= not b;
    layer5_outputs(2440) <= not (a or b);
    layer5_outputs(2441) <= not (a or b);
    layer5_outputs(2442) <= '1';
    layer5_outputs(2443) <= not b;
    layer5_outputs(2444) <= '1';
    layer5_outputs(2445) <= not a or b;
    layer5_outputs(2446) <= a and b;
    layer5_outputs(2447) <= b and not a;
    layer5_outputs(2448) <= a and b;
    layer5_outputs(2449) <= not a or b;
    layer5_outputs(2450) <= not (a or b);
    layer5_outputs(2451) <= '0';
    layer5_outputs(2452) <= a or b;
    layer5_outputs(2453) <= b;
    layer5_outputs(2454) <= not b;
    layer5_outputs(2455) <= not b;
    layer5_outputs(2456) <= not a;
    layer5_outputs(2457) <= not a or b;
    layer5_outputs(2458) <= a xor b;
    layer5_outputs(2459) <= not (a and b);
    layer5_outputs(2460) <= b and not a;
    layer5_outputs(2461) <= not (a and b);
    layer5_outputs(2462) <= '1';
    layer5_outputs(2463) <= a;
    layer5_outputs(2464) <= '0';
    layer5_outputs(2465) <= a or b;
    layer5_outputs(2466) <= a and not b;
    layer5_outputs(2467) <= not a or b;
    layer5_outputs(2468) <= b;
    layer5_outputs(2469) <= '0';
    layer5_outputs(2470) <= b;
    layer5_outputs(2471) <= not a or b;
    layer5_outputs(2472) <= a;
    layer5_outputs(2473) <= not b or a;
    layer5_outputs(2474) <= not b;
    layer5_outputs(2475) <= not (a and b);
    layer5_outputs(2476) <= not a or b;
    layer5_outputs(2477) <= a xor b;
    layer5_outputs(2478) <= a xor b;
    layer5_outputs(2479) <= a and b;
    layer5_outputs(2480) <= not (a or b);
    layer5_outputs(2481) <= a or b;
    layer5_outputs(2482) <= not (a and b);
    layer5_outputs(2483) <= not a or b;
    layer5_outputs(2484) <= not b;
    layer5_outputs(2485) <= b;
    layer5_outputs(2486) <= a;
    layer5_outputs(2487) <= not a;
    layer5_outputs(2488) <= a xor b;
    layer5_outputs(2489) <= a or b;
    layer5_outputs(2490) <= a or b;
    layer5_outputs(2491) <= a;
    layer5_outputs(2492) <= b and not a;
    layer5_outputs(2493) <= not (a xor b);
    layer5_outputs(2494) <= not (a or b);
    layer5_outputs(2495) <= '0';
    layer5_outputs(2496) <= a or b;
    layer5_outputs(2497) <= a and b;
    layer5_outputs(2498) <= '1';
    layer5_outputs(2499) <= not b;
    layer5_outputs(2500) <= '1';
    layer5_outputs(2501) <= not (a and b);
    layer5_outputs(2502) <= b and not a;
    layer5_outputs(2503) <= not a;
    layer5_outputs(2504) <= a or b;
    layer5_outputs(2505) <= not a;
    layer5_outputs(2506) <= b;
    layer5_outputs(2507) <= not a or b;
    layer5_outputs(2508) <= not (a and b);
    layer5_outputs(2509) <= a and not b;
    layer5_outputs(2510) <= not b or a;
    layer5_outputs(2511) <= a and b;
    layer5_outputs(2512) <= not a;
    layer5_outputs(2513) <= b;
    layer5_outputs(2514) <= b;
    layer5_outputs(2515) <= '1';
    layer5_outputs(2516) <= not (a and b);
    layer5_outputs(2517) <= a and b;
    layer5_outputs(2518) <= b and not a;
    layer5_outputs(2519) <= not (a or b);
    layer5_outputs(2520) <= a;
    layer5_outputs(2521) <= not b;
    layer5_outputs(2522) <= a and b;
    layer5_outputs(2523) <= not a;
    layer5_outputs(2524) <= a;
    layer5_outputs(2525) <= '1';
    layer5_outputs(2526) <= a and not b;
    layer5_outputs(2527) <= a xor b;
    layer5_outputs(2528) <= '1';
    layer5_outputs(2529) <= b;
    layer5_outputs(2530) <= a;
    layer5_outputs(2531) <= not a or b;
    layer5_outputs(2532) <= not b or a;
    layer5_outputs(2533) <= not a or b;
    layer5_outputs(2534) <= b;
    layer5_outputs(2535) <= a;
    layer5_outputs(2536) <= not a;
    layer5_outputs(2537) <= '1';
    layer5_outputs(2538) <= not (a and b);
    layer5_outputs(2539) <= b;
    layer5_outputs(2540) <= not b;
    layer5_outputs(2541) <= not a;
    layer5_outputs(2542) <= not a;
    layer5_outputs(2543) <= a and not b;
    layer5_outputs(2544) <= a and not b;
    layer5_outputs(2545) <= not b;
    layer5_outputs(2546) <= b;
    layer5_outputs(2547) <= b and not a;
    layer5_outputs(2548) <= not a or b;
    layer5_outputs(2549) <= not (a xor b);
    layer5_outputs(2550) <= a;
    layer5_outputs(2551) <= not b or a;
    layer5_outputs(2552) <= a or b;
    layer5_outputs(2553) <= not a;
    layer5_outputs(2554) <= a and not b;
    layer5_outputs(2555) <= not (a and b);
    layer5_outputs(2556) <= not a;
    layer5_outputs(2557) <= b;
    layer5_outputs(2558) <= not (a and b);
    layer5_outputs(2559) <= b;
    layer5_outputs(2560) <= not b or a;
    layer5_outputs(2561) <= not a;
    layer5_outputs(2562) <= b and not a;
    layer5_outputs(2563) <= not (a and b);
    layer5_outputs(2564) <= a xor b;
    layer5_outputs(2565) <= b;
    layer5_outputs(2566) <= b and not a;
    layer5_outputs(2567) <= not a;
    layer5_outputs(2568) <= not (a and b);
    layer5_outputs(2569) <= b;
    layer5_outputs(2570) <= a xor b;
    layer5_outputs(2571) <= '1';
    layer5_outputs(2572) <= not a;
    layer5_outputs(2573) <= not a or b;
    layer5_outputs(2574) <= '1';
    layer5_outputs(2575) <= not (a or b);
    layer5_outputs(2576) <= b;
    layer5_outputs(2577) <= not a or b;
    layer5_outputs(2578) <= a xor b;
    layer5_outputs(2579) <= a and b;
    layer5_outputs(2580) <= a and b;
    layer5_outputs(2581) <= not b or a;
    layer5_outputs(2582) <= not (a and b);
    layer5_outputs(2583) <= b;
    layer5_outputs(2584) <= not a;
    layer5_outputs(2585) <= a;
    layer5_outputs(2586) <= b;
    layer5_outputs(2587) <= not a;
    layer5_outputs(2588) <= not b or a;
    layer5_outputs(2589) <= not (a xor b);
    layer5_outputs(2590) <= not (a and b);
    layer5_outputs(2591) <= not (a or b);
    layer5_outputs(2592) <= a;
    layer5_outputs(2593) <= '0';
    layer5_outputs(2594) <= a xor b;
    layer5_outputs(2595) <= b and not a;
    layer5_outputs(2596) <= not a or b;
    layer5_outputs(2597) <= b;
    layer5_outputs(2598) <= a;
    layer5_outputs(2599) <= not b or a;
    layer5_outputs(2600) <= not a;
    layer5_outputs(2601) <= b;
    layer5_outputs(2602) <= not a;
    layer5_outputs(2603) <= not b;
    layer5_outputs(2604) <= not a;
    layer5_outputs(2605) <= not b;
    layer5_outputs(2606) <= '0';
    layer5_outputs(2607) <= not b or a;
    layer5_outputs(2608) <= b;
    layer5_outputs(2609) <= a or b;
    layer5_outputs(2610) <= not a or b;
    layer5_outputs(2611) <= not b or a;
    layer5_outputs(2612) <= not (a xor b);
    layer5_outputs(2613) <= not b;
    layer5_outputs(2614) <= not a;
    layer5_outputs(2615) <= not b;
    layer5_outputs(2616) <= a;
    layer5_outputs(2617) <= not a or b;
    layer5_outputs(2618) <= not (a or b);
    layer5_outputs(2619) <= not (a xor b);
    layer5_outputs(2620) <= b;
    layer5_outputs(2621) <= '1';
    layer5_outputs(2622) <= a xor b;
    layer5_outputs(2623) <= b;
    layer5_outputs(2624) <= not b;
    layer5_outputs(2625) <= a and b;
    layer5_outputs(2626) <= a;
    layer5_outputs(2627) <= a or b;
    layer5_outputs(2628) <= a and b;
    layer5_outputs(2629) <= a xor b;
    layer5_outputs(2630) <= b;
    layer5_outputs(2631) <= a and b;
    layer5_outputs(2632) <= a;
    layer5_outputs(2633) <= not b;
    layer5_outputs(2634) <= b and not a;
    layer5_outputs(2635) <= a or b;
    layer5_outputs(2636) <= not b;
    layer5_outputs(2637) <= b;
    layer5_outputs(2638) <= not a;
    layer5_outputs(2639) <= b;
    layer5_outputs(2640) <= a;
    layer5_outputs(2641) <= not a or b;
    layer5_outputs(2642) <= not (a or b);
    layer5_outputs(2643) <= not (a and b);
    layer5_outputs(2644) <= a;
    layer5_outputs(2645) <= not (a or b);
    layer5_outputs(2646) <= not (a or b);
    layer5_outputs(2647) <= b and not a;
    layer5_outputs(2648) <= a and b;
    layer5_outputs(2649) <= b;
    layer5_outputs(2650) <= a or b;
    layer5_outputs(2651) <= not b or a;
    layer5_outputs(2652) <= not b;
    layer5_outputs(2653) <= not b or a;
    layer5_outputs(2654) <= b;
    layer5_outputs(2655) <= b and not a;
    layer5_outputs(2656) <= a;
    layer5_outputs(2657) <= not (a or b);
    layer5_outputs(2658) <= b and not a;
    layer5_outputs(2659) <= not (a or b);
    layer5_outputs(2660) <= a xor b;
    layer5_outputs(2661) <= a;
    layer5_outputs(2662) <= not b;
    layer5_outputs(2663) <= not a;
    layer5_outputs(2664) <= b and not a;
    layer5_outputs(2665) <= not a;
    layer5_outputs(2666) <= a and not b;
    layer5_outputs(2667) <= not b;
    layer5_outputs(2668) <= not a;
    layer5_outputs(2669) <= not (a or b);
    layer5_outputs(2670) <= not a or b;
    layer5_outputs(2671) <= a xor b;
    layer5_outputs(2672) <= b;
    layer5_outputs(2673) <= a and not b;
    layer5_outputs(2674) <= not b;
    layer5_outputs(2675) <= a and b;
    layer5_outputs(2676) <= b;
    layer5_outputs(2677) <= not b;
    layer5_outputs(2678) <= b;
    layer5_outputs(2679) <= a;
    layer5_outputs(2680) <= not b;
    layer5_outputs(2681) <= a;
    layer5_outputs(2682) <= a;
    layer5_outputs(2683) <= not b or a;
    layer5_outputs(2684) <= not (a and b);
    layer5_outputs(2685) <= a or b;
    layer5_outputs(2686) <= a and b;
    layer5_outputs(2687) <= '1';
    layer5_outputs(2688) <= '1';
    layer5_outputs(2689) <= not a or b;
    layer5_outputs(2690) <= a xor b;
    layer5_outputs(2691) <= a and not b;
    layer5_outputs(2692) <= b and not a;
    layer5_outputs(2693) <= not (a xor b);
    layer5_outputs(2694) <= a and b;
    layer5_outputs(2695) <= not a;
    layer5_outputs(2696) <= a and b;
    layer5_outputs(2697) <= not a;
    layer5_outputs(2698) <= not a or b;
    layer5_outputs(2699) <= a and b;
    layer5_outputs(2700) <= a and b;
    layer5_outputs(2701) <= b and not a;
    layer5_outputs(2702) <= not a;
    layer5_outputs(2703) <= a and not b;
    layer5_outputs(2704) <= a;
    layer5_outputs(2705) <= a and not b;
    layer5_outputs(2706) <= b and not a;
    layer5_outputs(2707) <= a or b;
    layer5_outputs(2708) <= not a or b;
    layer5_outputs(2709) <= not (a or b);
    layer5_outputs(2710) <= b;
    layer5_outputs(2711) <= '0';
    layer5_outputs(2712) <= a or b;
    layer5_outputs(2713) <= b;
    layer5_outputs(2714) <= not a or b;
    layer5_outputs(2715) <= not (a or b);
    layer5_outputs(2716) <= not a;
    layer5_outputs(2717) <= not (a and b);
    layer5_outputs(2718) <= '0';
    layer5_outputs(2719) <= not (a and b);
    layer5_outputs(2720) <= a;
    layer5_outputs(2721) <= a and b;
    layer5_outputs(2722) <= not a;
    layer5_outputs(2723) <= '0';
    layer5_outputs(2724) <= a or b;
    layer5_outputs(2725) <= '0';
    layer5_outputs(2726) <= a;
    layer5_outputs(2727) <= a and b;
    layer5_outputs(2728) <= a;
    layer5_outputs(2729) <= '1';
    layer5_outputs(2730) <= a and not b;
    layer5_outputs(2731) <= not a;
    layer5_outputs(2732) <= not b or a;
    layer5_outputs(2733) <= a and b;
    layer5_outputs(2734) <= not (a xor b);
    layer5_outputs(2735) <= a;
    layer5_outputs(2736) <= a;
    layer5_outputs(2737) <= not b;
    layer5_outputs(2738) <= not (a xor b);
    layer5_outputs(2739) <= a;
    layer5_outputs(2740) <= '0';
    layer5_outputs(2741) <= a xor b;
    layer5_outputs(2742) <= not b;
    layer5_outputs(2743) <= a and b;
    layer5_outputs(2744) <= '1';
    layer5_outputs(2745) <= not b or a;
    layer5_outputs(2746) <= b;
    layer5_outputs(2747) <= a;
    layer5_outputs(2748) <= b;
    layer5_outputs(2749) <= '1';
    layer5_outputs(2750) <= a or b;
    layer5_outputs(2751) <= a or b;
    layer5_outputs(2752) <= a xor b;
    layer5_outputs(2753) <= a and not b;
    layer5_outputs(2754) <= not b;
    layer5_outputs(2755) <= not a or b;
    layer5_outputs(2756) <= '0';
    layer5_outputs(2757) <= a;
    layer5_outputs(2758) <= not (a and b);
    layer5_outputs(2759) <= a xor b;
    layer5_outputs(2760) <= a and not b;
    layer5_outputs(2761) <= b;
    layer5_outputs(2762) <= b;
    layer5_outputs(2763) <= a or b;
    layer5_outputs(2764) <= b and not a;
    layer5_outputs(2765) <= not (a and b);
    layer5_outputs(2766) <= a;
    layer5_outputs(2767) <= not b or a;
    layer5_outputs(2768) <= a and not b;
    layer5_outputs(2769) <= a or b;
    layer5_outputs(2770) <= not b;
    layer5_outputs(2771) <= a and not b;
    layer5_outputs(2772) <= not a;
    layer5_outputs(2773) <= not a or b;
    layer5_outputs(2774) <= '0';
    layer5_outputs(2775) <= not b;
    layer5_outputs(2776) <= not (a and b);
    layer5_outputs(2777) <= a and b;
    layer5_outputs(2778) <= a and not b;
    layer5_outputs(2779) <= b;
    layer5_outputs(2780) <= not (a and b);
    layer5_outputs(2781) <= a xor b;
    layer5_outputs(2782) <= b and not a;
    layer5_outputs(2783) <= a and b;
    layer5_outputs(2784) <= not b or a;
    layer5_outputs(2785) <= not a;
    layer5_outputs(2786) <= not (a and b);
    layer5_outputs(2787) <= not a;
    layer5_outputs(2788) <= a and b;
    layer5_outputs(2789) <= a;
    layer5_outputs(2790) <= not b;
    layer5_outputs(2791) <= a and b;
    layer5_outputs(2792) <= b;
    layer5_outputs(2793) <= b;
    layer5_outputs(2794) <= not b or a;
    layer5_outputs(2795) <= a or b;
    layer5_outputs(2796) <= '1';
    layer5_outputs(2797) <= a or b;
    layer5_outputs(2798) <= a and not b;
    layer5_outputs(2799) <= not b or a;
    layer5_outputs(2800) <= a xor b;
    layer5_outputs(2801) <= not b or a;
    layer5_outputs(2802) <= not b or a;
    layer5_outputs(2803) <= a xor b;
    layer5_outputs(2804) <= not b or a;
    layer5_outputs(2805) <= not (a and b);
    layer5_outputs(2806) <= a or b;
    layer5_outputs(2807) <= a;
    layer5_outputs(2808) <= a xor b;
    layer5_outputs(2809) <= not a or b;
    layer5_outputs(2810) <= a xor b;
    layer5_outputs(2811) <= b;
    layer5_outputs(2812) <= not a or b;
    layer5_outputs(2813) <= not b;
    layer5_outputs(2814) <= not b or a;
    layer5_outputs(2815) <= a and b;
    layer5_outputs(2816) <= not a;
    layer5_outputs(2817) <= not a;
    layer5_outputs(2818) <= not (a and b);
    layer5_outputs(2819) <= not (a xor b);
    layer5_outputs(2820) <= a or b;
    layer5_outputs(2821) <= not b;
    layer5_outputs(2822) <= b;
    layer5_outputs(2823) <= not a or b;
    layer5_outputs(2824) <= a and not b;
    layer5_outputs(2825) <= not b or a;
    layer5_outputs(2826) <= not b or a;
    layer5_outputs(2827) <= not b or a;
    layer5_outputs(2828) <= a and not b;
    layer5_outputs(2829) <= not a or b;
    layer5_outputs(2830) <= not (a xor b);
    layer5_outputs(2831) <= b and not a;
    layer5_outputs(2832) <= b;
    layer5_outputs(2833) <= not a or b;
    layer5_outputs(2834) <= a or b;
    layer5_outputs(2835) <= not (a or b);
    layer5_outputs(2836) <= b;
    layer5_outputs(2837) <= a and not b;
    layer5_outputs(2838) <= not (a xor b);
    layer5_outputs(2839) <= not (a or b);
    layer5_outputs(2840) <= a;
    layer5_outputs(2841) <= a;
    layer5_outputs(2842) <= a and b;
    layer5_outputs(2843) <= '1';
    layer5_outputs(2844) <= b and not a;
    layer5_outputs(2845) <= '0';
    layer5_outputs(2846) <= not (a and b);
    layer5_outputs(2847) <= b and not a;
    layer5_outputs(2848) <= not b or a;
    layer5_outputs(2849) <= b and not a;
    layer5_outputs(2850) <= not b;
    layer5_outputs(2851) <= b and not a;
    layer5_outputs(2852) <= not a or b;
    layer5_outputs(2853) <= a or b;
    layer5_outputs(2854) <= not (a or b);
    layer5_outputs(2855) <= b;
    layer5_outputs(2856) <= a and not b;
    layer5_outputs(2857) <= a;
    layer5_outputs(2858) <= b;
    layer5_outputs(2859) <= a;
    layer5_outputs(2860) <= a and not b;
    layer5_outputs(2861) <= not (a or b);
    layer5_outputs(2862) <= b;
    layer5_outputs(2863) <= b;
    layer5_outputs(2864) <= a or b;
    layer5_outputs(2865) <= not a or b;
    layer5_outputs(2866) <= not a or b;
    layer5_outputs(2867) <= not (a or b);
    layer5_outputs(2868) <= not b;
    layer5_outputs(2869) <= '1';
    layer5_outputs(2870) <= b;
    layer5_outputs(2871) <= a and b;
    layer5_outputs(2872) <= a and b;
    layer5_outputs(2873) <= not b;
    layer5_outputs(2874) <= not (a or b);
    layer5_outputs(2875) <= not (a and b);
    layer5_outputs(2876) <= b;
    layer5_outputs(2877) <= a and not b;
    layer5_outputs(2878) <= not b;
    layer5_outputs(2879) <= a;
    layer5_outputs(2880) <= not (a or b);
    layer5_outputs(2881) <= b and not a;
    layer5_outputs(2882) <= b;
    layer5_outputs(2883) <= a and not b;
    layer5_outputs(2884) <= a;
    layer5_outputs(2885) <= b and not a;
    layer5_outputs(2886) <= not (a and b);
    layer5_outputs(2887) <= not (a or b);
    layer5_outputs(2888) <= a or b;
    layer5_outputs(2889) <= not (a xor b);
    layer5_outputs(2890) <= b and not a;
    layer5_outputs(2891) <= a and b;
    layer5_outputs(2892) <= not a;
    layer5_outputs(2893) <= not (a or b);
    layer5_outputs(2894) <= '1';
    layer5_outputs(2895) <= not a or b;
    layer5_outputs(2896) <= not (a xor b);
    layer5_outputs(2897) <= a and b;
    layer5_outputs(2898) <= not a;
    layer5_outputs(2899) <= not a;
    layer5_outputs(2900) <= b;
    layer5_outputs(2901) <= not (a and b);
    layer5_outputs(2902) <= '0';
    layer5_outputs(2903) <= a xor b;
    layer5_outputs(2904) <= not a or b;
    layer5_outputs(2905) <= b and not a;
    layer5_outputs(2906) <= not (a or b);
    layer5_outputs(2907) <= not (a xor b);
    layer5_outputs(2908) <= not b;
    layer5_outputs(2909) <= not b;
    layer5_outputs(2910) <= not a;
    layer5_outputs(2911) <= not a or b;
    layer5_outputs(2912) <= not b;
    layer5_outputs(2913) <= not (a or b);
    layer5_outputs(2914) <= not b;
    layer5_outputs(2915) <= not a;
    layer5_outputs(2916) <= a or b;
    layer5_outputs(2917) <= not (a xor b);
    layer5_outputs(2918) <= not (a and b);
    layer5_outputs(2919) <= b and not a;
    layer5_outputs(2920) <= b;
    layer5_outputs(2921) <= not a;
    layer5_outputs(2922) <= '0';
    layer5_outputs(2923) <= a and b;
    layer5_outputs(2924) <= not (a and b);
    layer5_outputs(2925) <= not a;
    layer5_outputs(2926) <= not b or a;
    layer5_outputs(2927) <= a;
    layer5_outputs(2928) <= a or b;
    layer5_outputs(2929) <= b and not a;
    layer5_outputs(2930) <= a xor b;
    layer5_outputs(2931) <= b;
    layer5_outputs(2932) <= not (a or b);
    layer5_outputs(2933) <= '1';
    layer5_outputs(2934) <= a;
    layer5_outputs(2935) <= not b;
    layer5_outputs(2936) <= not a;
    layer5_outputs(2937) <= not (a xor b);
    layer5_outputs(2938) <= not b or a;
    layer5_outputs(2939) <= not (a xor b);
    layer5_outputs(2940) <= a xor b;
    layer5_outputs(2941) <= '1';
    layer5_outputs(2942) <= b and not a;
    layer5_outputs(2943) <= b;
    layer5_outputs(2944) <= a;
    layer5_outputs(2945) <= not a or b;
    layer5_outputs(2946) <= not a;
    layer5_outputs(2947) <= a xor b;
    layer5_outputs(2948) <= not b or a;
    layer5_outputs(2949) <= '1';
    layer5_outputs(2950) <= not a;
    layer5_outputs(2951) <= a or b;
    layer5_outputs(2952) <= a;
    layer5_outputs(2953) <= a and not b;
    layer5_outputs(2954) <= not (a and b);
    layer5_outputs(2955) <= b and not a;
    layer5_outputs(2956) <= a or b;
    layer5_outputs(2957) <= a and not b;
    layer5_outputs(2958) <= not (a and b);
    layer5_outputs(2959) <= a and not b;
    layer5_outputs(2960) <= a xor b;
    layer5_outputs(2961) <= not b;
    layer5_outputs(2962) <= not (a xor b);
    layer5_outputs(2963) <= a;
    layer5_outputs(2964) <= not (a or b);
    layer5_outputs(2965) <= '1';
    layer5_outputs(2966) <= b and not a;
    layer5_outputs(2967) <= not (a or b);
    layer5_outputs(2968) <= not b or a;
    layer5_outputs(2969) <= not a;
    layer5_outputs(2970) <= not a;
    layer5_outputs(2971) <= b;
    layer5_outputs(2972) <= not b or a;
    layer5_outputs(2973) <= a and b;
    layer5_outputs(2974) <= not a;
    layer5_outputs(2975) <= a or b;
    layer5_outputs(2976) <= not (a and b);
    layer5_outputs(2977) <= a;
    layer5_outputs(2978) <= not a;
    layer5_outputs(2979) <= a;
    layer5_outputs(2980) <= a;
    layer5_outputs(2981) <= '0';
    layer5_outputs(2982) <= a and not b;
    layer5_outputs(2983) <= '0';
    layer5_outputs(2984) <= not (a or b);
    layer5_outputs(2985) <= b and not a;
    layer5_outputs(2986) <= a;
    layer5_outputs(2987) <= not b;
    layer5_outputs(2988) <= a xor b;
    layer5_outputs(2989) <= '1';
    layer5_outputs(2990) <= '1';
    layer5_outputs(2991) <= b and not a;
    layer5_outputs(2992) <= not a;
    layer5_outputs(2993) <= not a or b;
    layer5_outputs(2994) <= not a;
    layer5_outputs(2995) <= '0';
    layer5_outputs(2996) <= not a;
    layer5_outputs(2997) <= a or b;
    layer5_outputs(2998) <= b and not a;
    layer5_outputs(2999) <= not a;
    layer5_outputs(3000) <= a;
    layer5_outputs(3001) <= b;
    layer5_outputs(3002) <= b and not a;
    layer5_outputs(3003) <= not b or a;
    layer5_outputs(3004) <= b;
    layer5_outputs(3005) <= not a or b;
    layer5_outputs(3006) <= b and not a;
    layer5_outputs(3007) <= a and b;
    layer5_outputs(3008) <= not a;
    layer5_outputs(3009) <= not b or a;
    layer5_outputs(3010) <= a;
    layer5_outputs(3011) <= not a;
    layer5_outputs(3012) <= not b or a;
    layer5_outputs(3013) <= a and b;
    layer5_outputs(3014) <= a and b;
    layer5_outputs(3015) <= a;
    layer5_outputs(3016) <= not a;
    layer5_outputs(3017) <= not b;
    layer5_outputs(3018) <= b and not a;
    layer5_outputs(3019) <= '0';
    layer5_outputs(3020) <= not b;
    layer5_outputs(3021) <= not a or b;
    layer5_outputs(3022) <= b;
    layer5_outputs(3023) <= not (a or b);
    layer5_outputs(3024) <= a and not b;
    layer5_outputs(3025) <= not a;
    layer5_outputs(3026) <= a;
    layer5_outputs(3027) <= a and b;
    layer5_outputs(3028) <= b;
    layer5_outputs(3029) <= not b;
    layer5_outputs(3030) <= a xor b;
    layer5_outputs(3031) <= a xor b;
    layer5_outputs(3032) <= a and not b;
    layer5_outputs(3033) <= not (a and b);
    layer5_outputs(3034) <= not b;
    layer5_outputs(3035) <= a or b;
    layer5_outputs(3036) <= not (a and b);
    layer5_outputs(3037) <= not (a xor b);
    layer5_outputs(3038) <= not b;
    layer5_outputs(3039) <= not b or a;
    layer5_outputs(3040) <= a or b;
    layer5_outputs(3041) <= a and not b;
    layer5_outputs(3042) <= not a;
    layer5_outputs(3043) <= not b or a;
    layer5_outputs(3044) <= not b;
    layer5_outputs(3045) <= b and not a;
    layer5_outputs(3046) <= not a or b;
    layer5_outputs(3047) <= not (a or b);
    layer5_outputs(3048) <= not b;
    layer5_outputs(3049) <= '0';
    layer5_outputs(3050) <= not b or a;
    layer5_outputs(3051) <= not b;
    layer5_outputs(3052) <= not b;
    layer5_outputs(3053) <= not (a or b);
    layer5_outputs(3054) <= not b or a;
    layer5_outputs(3055) <= b and not a;
    layer5_outputs(3056) <= a xor b;
    layer5_outputs(3057) <= '0';
    layer5_outputs(3058) <= not (a and b);
    layer5_outputs(3059) <= b;
    layer5_outputs(3060) <= not (a and b);
    layer5_outputs(3061) <= a xor b;
    layer5_outputs(3062) <= not a;
    layer5_outputs(3063) <= not b;
    layer5_outputs(3064) <= not b or a;
    layer5_outputs(3065) <= a and not b;
    layer5_outputs(3066) <= b;
    layer5_outputs(3067) <= a and b;
    layer5_outputs(3068) <= not (a or b);
    layer5_outputs(3069) <= not b or a;
    layer5_outputs(3070) <= '1';
    layer5_outputs(3071) <= not a or b;
    layer5_outputs(3072) <= not b or a;
    layer5_outputs(3073) <= not b;
    layer5_outputs(3074) <= not a;
    layer5_outputs(3075) <= not a or b;
    layer5_outputs(3076) <= not b;
    layer5_outputs(3077) <= not (a or b);
    layer5_outputs(3078) <= b;
    layer5_outputs(3079) <= not (a or b);
    layer5_outputs(3080) <= b;
    layer5_outputs(3081) <= b and not a;
    layer5_outputs(3082) <= a and b;
    layer5_outputs(3083) <= a xor b;
    layer5_outputs(3084) <= not a;
    layer5_outputs(3085) <= not a or b;
    layer5_outputs(3086) <= a and b;
    layer5_outputs(3087) <= a;
    layer5_outputs(3088) <= not a;
    layer5_outputs(3089) <= not (a xor b);
    layer5_outputs(3090) <= not a;
    layer5_outputs(3091) <= a and not b;
    layer5_outputs(3092) <= '1';
    layer5_outputs(3093) <= a or b;
    layer5_outputs(3094) <= not a or b;
    layer5_outputs(3095) <= a;
    layer5_outputs(3096) <= a;
    layer5_outputs(3097) <= a;
    layer5_outputs(3098) <= not (a or b);
    layer5_outputs(3099) <= b and not a;
    layer5_outputs(3100) <= a or b;
    layer5_outputs(3101) <= a;
    layer5_outputs(3102) <= not (a or b);
    layer5_outputs(3103) <= not (a or b);
    layer5_outputs(3104) <= a;
    layer5_outputs(3105) <= b;
    layer5_outputs(3106) <= a or b;
    layer5_outputs(3107) <= not b;
    layer5_outputs(3108) <= '0';
    layer5_outputs(3109) <= b;
    layer5_outputs(3110) <= not a;
    layer5_outputs(3111) <= b;
    layer5_outputs(3112) <= a xor b;
    layer5_outputs(3113) <= a;
    layer5_outputs(3114) <= b and not a;
    layer5_outputs(3115) <= b;
    layer5_outputs(3116) <= not a;
    layer5_outputs(3117) <= not (a or b);
    layer5_outputs(3118) <= not (a or b);
    layer5_outputs(3119) <= b and not a;
    layer5_outputs(3120) <= b and not a;
    layer5_outputs(3121) <= not b;
    layer5_outputs(3122) <= not b or a;
    layer5_outputs(3123) <= a xor b;
    layer5_outputs(3124) <= '1';
    layer5_outputs(3125) <= a xor b;
    layer5_outputs(3126) <= a;
    layer5_outputs(3127) <= not a;
    layer5_outputs(3128) <= b;
    layer5_outputs(3129) <= b;
    layer5_outputs(3130) <= b;
    layer5_outputs(3131) <= b;
    layer5_outputs(3132) <= a or b;
    layer5_outputs(3133) <= not b;
    layer5_outputs(3134) <= not a;
    layer5_outputs(3135) <= '0';
    layer5_outputs(3136) <= '0';
    layer5_outputs(3137) <= b;
    layer5_outputs(3138) <= a;
    layer5_outputs(3139) <= not b or a;
    layer5_outputs(3140) <= '1';
    layer5_outputs(3141) <= not (a and b);
    layer5_outputs(3142) <= b and not a;
    layer5_outputs(3143) <= not b;
    layer5_outputs(3144) <= a;
    layer5_outputs(3145) <= not (a or b);
    layer5_outputs(3146) <= a and not b;
    layer5_outputs(3147) <= not (a and b);
    layer5_outputs(3148) <= not a or b;
    layer5_outputs(3149) <= not (a and b);
    layer5_outputs(3150) <= b and not a;
    layer5_outputs(3151) <= not b or a;
    layer5_outputs(3152) <= a;
    layer5_outputs(3153) <= not a;
    layer5_outputs(3154) <= not (a or b);
    layer5_outputs(3155) <= a and not b;
    layer5_outputs(3156) <= not a;
    layer5_outputs(3157) <= a or b;
    layer5_outputs(3158) <= a and not b;
    layer5_outputs(3159) <= a and not b;
    layer5_outputs(3160) <= a xor b;
    layer5_outputs(3161) <= not a or b;
    layer5_outputs(3162) <= b;
    layer5_outputs(3163) <= not a;
    layer5_outputs(3164) <= a and not b;
    layer5_outputs(3165) <= not a;
    layer5_outputs(3166) <= not b;
    layer5_outputs(3167) <= b;
    layer5_outputs(3168) <= b and not a;
    layer5_outputs(3169) <= not b or a;
    layer5_outputs(3170) <= not a;
    layer5_outputs(3171) <= not (a and b);
    layer5_outputs(3172) <= a and b;
    layer5_outputs(3173) <= '0';
    layer5_outputs(3174) <= not a;
    layer5_outputs(3175) <= not b;
    layer5_outputs(3176) <= a or b;
    layer5_outputs(3177) <= not b or a;
    layer5_outputs(3178) <= not (a xor b);
    layer5_outputs(3179) <= not a;
    layer5_outputs(3180) <= not b;
    layer5_outputs(3181) <= '1';
    layer5_outputs(3182) <= b and not a;
    layer5_outputs(3183) <= a or b;
    layer5_outputs(3184) <= not b;
    layer5_outputs(3185) <= not b;
    layer5_outputs(3186) <= a and b;
    layer5_outputs(3187) <= not a;
    layer5_outputs(3188) <= a and b;
    layer5_outputs(3189) <= not a;
    layer5_outputs(3190) <= not a or b;
    layer5_outputs(3191) <= a;
    layer5_outputs(3192) <= b and not a;
    layer5_outputs(3193) <= '0';
    layer5_outputs(3194) <= not a or b;
    layer5_outputs(3195) <= a and not b;
    layer5_outputs(3196) <= b;
    layer5_outputs(3197) <= a and b;
    layer5_outputs(3198) <= not (a or b);
    layer5_outputs(3199) <= a and b;
    layer5_outputs(3200) <= not (a xor b);
    layer5_outputs(3201) <= a or b;
    layer5_outputs(3202) <= not (a or b);
    layer5_outputs(3203) <= not (a or b);
    layer5_outputs(3204) <= a and b;
    layer5_outputs(3205) <= a;
    layer5_outputs(3206) <= not b;
    layer5_outputs(3207) <= '0';
    layer5_outputs(3208) <= a;
    layer5_outputs(3209) <= not (a or b);
    layer5_outputs(3210) <= '0';
    layer5_outputs(3211) <= b;
    layer5_outputs(3212) <= not (a and b);
    layer5_outputs(3213) <= a and not b;
    layer5_outputs(3214) <= not (a and b);
    layer5_outputs(3215) <= not (a or b);
    layer5_outputs(3216) <= b and not a;
    layer5_outputs(3217) <= not (a or b);
    layer5_outputs(3218) <= b;
    layer5_outputs(3219) <= not (a and b);
    layer5_outputs(3220) <= not (a and b);
    layer5_outputs(3221) <= '0';
    layer5_outputs(3222) <= not a;
    layer5_outputs(3223) <= not b;
    layer5_outputs(3224) <= a or b;
    layer5_outputs(3225) <= not (a or b);
    layer5_outputs(3226) <= b;
    layer5_outputs(3227) <= a and b;
    layer5_outputs(3228) <= not b or a;
    layer5_outputs(3229) <= a and not b;
    layer5_outputs(3230) <= a and b;
    layer5_outputs(3231) <= '0';
    layer5_outputs(3232) <= not a or b;
    layer5_outputs(3233) <= b;
    layer5_outputs(3234) <= a xor b;
    layer5_outputs(3235) <= b;
    layer5_outputs(3236) <= '1';
    layer5_outputs(3237) <= a;
    layer5_outputs(3238) <= a or b;
    layer5_outputs(3239) <= b;
    layer5_outputs(3240) <= a and not b;
    layer5_outputs(3241) <= not (a or b);
    layer5_outputs(3242) <= not (a and b);
    layer5_outputs(3243) <= not (a or b);
    layer5_outputs(3244) <= not (a and b);
    layer5_outputs(3245) <= not a;
    layer5_outputs(3246) <= a and b;
    layer5_outputs(3247) <= a and b;
    layer5_outputs(3248) <= not b;
    layer5_outputs(3249) <= not a or b;
    layer5_outputs(3250) <= not (a or b);
    layer5_outputs(3251) <= not (a or b);
    layer5_outputs(3252) <= not b;
    layer5_outputs(3253) <= not (a and b);
    layer5_outputs(3254) <= not (a or b);
    layer5_outputs(3255) <= not a;
    layer5_outputs(3256) <= a;
    layer5_outputs(3257) <= not b or a;
    layer5_outputs(3258) <= a and not b;
    layer5_outputs(3259) <= a xor b;
    layer5_outputs(3260) <= b and not a;
    layer5_outputs(3261) <= b;
    layer5_outputs(3262) <= not (a or b);
    layer5_outputs(3263) <= not (a and b);
    layer5_outputs(3264) <= not (a and b);
    layer5_outputs(3265) <= '0';
    layer5_outputs(3266) <= not a;
    layer5_outputs(3267) <= '1';
    layer5_outputs(3268) <= not a or b;
    layer5_outputs(3269) <= not a or b;
    layer5_outputs(3270) <= a and not b;
    layer5_outputs(3271) <= a or b;
    layer5_outputs(3272) <= a and b;
    layer5_outputs(3273) <= not b;
    layer5_outputs(3274) <= not b;
    layer5_outputs(3275) <= not (a or b);
    layer5_outputs(3276) <= not (a xor b);
    layer5_outputs(3277) <= a xor b;
    layer5_outputs(3278) <= not a or b;
    layer5_outputs(3279) <= a;
    layer5_outputs(3280) <= not a;
    layer5_outputs(3281) <= a;
    layer5_outputs(3282) <= not (a and b);
    layer5_outputs(3283) <= a and b;
    layer5_outputs(3284) <= not b;
    layer5_outputs(3285) <= '0';
    layer5_outputs(3286) <= a;
    layer5_outputs(3287) <= not b;
    layer5_outputs(3288) <= a and b;
    layer5_outputs(3289) <= a;
    layer5_outputs(3290) <= a and not b;
    layer5_outputs(3291) <= not (a and b);
    layer5_outputs(3292) <= a and b;
    layer5_outputs(3293) <= a;
    layer5_outputs(3294) <= b and not a;
    layer5_outputs(3295) <= not b;
    layer5_outputs(3296) <= a or b;
    layer5_outputs(3297) <= not b;
    layer5_outputs(3298) <= '1';
    layer5_outputs(3299) <= not b or a;
    layer5_outputs(3300) <= a and b;
    layer5_outputs(3301) <= a and not b;
    layer5_outputs(3302) <= a;
    layer5_outputs(3303) <= not (a or b);
    layer5_outputs(3304) <= '1';
    layer5_outputs(3305) <= not b;
    layer5_outputs(3306) <= b and not a;
    layer5_outputs(3307) <= not b or a;
    layer5_outputs(3308) <= not b or a;
    layer5_outputs(3309) <= a;
    layer5_outputs(3310) <= a and b;
    layer5_outputs(3311) <= a;
    layer5_outputs(3312) <= not a;
    layer5_outputs(3313) <= a;
    layer5_outputs(3314) <= b;
    layer5_outputs(3315) <= not b;
    layer5_outputs(3316) <= b;
    layer5_outputs(3317) <= a and b;
    layer5_outputs(3318) <= b;
    layer5_outputs(3319) <= a xor b;
    layer5_outputs(3320) <= a;
    layer5_outputs(3321) <= not b;
    layer5_outputs(3322) <= b and not a;
    layer5_outputs(3323) <= not a or b;
    layer5_outputs(3324) <= a;
    layer5_outputs(3325) <= not a;
    layer5_outputs(3326) <= a and not b;
    layer5_outputs(3327) <= a and not b;
    layer5_outputs(3328) <= not b;
    layer5_outputs(3329) <= not (a and b);
    layer5_outputs(3330) <= not a;
    layer5_outputs(3331) <= not a;
    layer5_outputs(3332) <= not a;
    layer5_outputs(3333) <= not (a and b);
    layer5_outputs(3334) <= a and b;
    layer5_outputs(3335) <= not a or b;
    layer5_outputs(3336) <= a;
    layer5_outputs(3337) <= a and not b;
    layer5_outputs(3338) <= not a;
    layer5_outputs(3339) <= not b;
    layer5_outputs(3340) <= b;
    layer5_outputs(3341) <= b;
    layer5_outputs(3342) <= b;
    layer5_outputs(3343) <= not a or b;
    layer5_outputs(3344) <= not (a xor b);
    layer5_outputs(3345) <= b and not a;
    layer5_outputs(3346) <= not (a and b);
    layer5_outputs(3347) <= a and not b;
    layer5_outputs(3348) <= a and b;
    layer5_outputs(3349) <= not b;
    layer5_outputs(3350) <= a and b;
    layer5_outputs(3351) <= not (a xor b);
    layer5_outputs(3352) <= not (a or b);
    layer5_outputs(3353) <= b;
    layer5_outputs(3354) <= not (a or b);
    layer5_outputs(3355) <= not b or a;
    layer5_outputs(3356) <= not a or b;
    layer5_outputs(3357) <= a;
    layer5_outputs(3358) <= not (a or b);
    layer5_outputs(3359) <= a;
    layer5_outputs(3360) <= b;
    layer5_outputs(3361) <= not b or a;
    layer5_outputs(3362) <= a;
    layer5_outputs(3363) <= b;
    layer5_outputs(3364) <= b;
    layer5_outputs(3365) <= not (a and b);
    layer5_outputs(3366) <= not (a or b);
    layer5_outputs(3367) <= not a;
    layer5_outputs(3368) <= not a or b;
    layer5_outputs(3369) <= not a or b;
    layer5_outputs(3370) <= a and b;
    layer5_outputs(3371) <= a or b;
    layer5_outputs(3372) <= a and b;
    layer5_outputs(3373) <= not (a or b);
    layer5_outputs(3374) <= not a or b;
    layer5_outputs(3375) <= not b;
    layer5_outputs(3376) <= not b or a;
    layer5_outputs(3377) <= b;
    layer5_outputs(3378) <= not a or b;
    layer5_outputs(3379) <= a;
    layer5_outputs(3380) <= not b or a;
    layer5_outputs(3381) <= a xor b;
    layer5_outputs(3382) <= not (a and b);
    layer5_outputs(3383) <= not a or b;
    layer5_outputs(3384) <= b and not a;
    layer5_outputs(3385) <= not (a xor b);
    layer5_outputs(3386) <= not (a or b);
    layer5_outputs(3387) <= not a or b;
    layer5_outputs(3388) <= not (a xor b);
    layer5_outputs(3389) <= not (a and b);
    layer5_outputs(3390) <= not (a or b);
    layer5_outputs(3391) <= not (a or b);
    layer5_outputs(3392) <= not b or a;
    layer5_outputs(3393) <= not a;
    layer5_outputs(3394) <= not b or a;
    layer5_outputs(3395) <= not a;
    layer5_outputs(3396) <= not b or a;
    layer5_outputs(3397) <= not a;
    layer5_outputs(3398) <= b;
    layer5_outputs(3399) <= a and b;
    layer5_outputs(3400) <= a;
    layer5_outputs(3401) <= not a;
    layer5_outputs(3402) <= not (a and b);
    layer5_outputs(3403) <= a and b;
    layer5_outputs(3404) <= '1';
    layer5_outputs(3405) <= a and not b;
    layer5_outputs(3406) <= a and not b;
    layer5_outputs(3407) <= not (a and b);
    layer5_outputs(3408) <= not a or b;
    layer5_outputs(3409) <= a or b;
    layer5_outputs(3410) <= b;
    layer5_outputs(3411) <= not (a xor b);
    layer5_outputs(3412) <= a and b;
    layer5_outputs(3413) <= '0';
    layer5_outputs(3414) <= not a;
    layer5_outputs(3415) <= not b or a;
    layer5_outputs(3416) <= '0';
    layer5_outputs(3417) <= b and not a;
    layer5_outputs(3418) <= b and not a;
    layer5_outputs(3419) <= a or b;
    layer5_outputs(3420) <= not a;
    layer5_outputs(3421) <= a and b;
    layer5_outputs(3422) <= not a;
    layer5_outputs(3423) <= a or b;
    layer5_outputs(3424) <= a;
    layer5_outputs(3425) <= a xor b;
    layer5_outputs(3426) <= '0';
    layer5_outputs(3427) <= a and b;
    layer5_outputs(3428) <= b and not a;
    layer5_outputs(3429) <= not a;
    layer5_outputs(3430) <= not a;
    layer5_outputs(3431) <= not b or a;
    layer5_outputs(3432) <= not (a and b);
    layer5_outputs(3433) <= a and b;
    layer5_outputs(3434) <= not a or b;
    layer5_outputs(3435) <= b;
    layer5_outputs(3436) <= not (a and b);
    layer5_outputs(3437) <= a and b;
    layer5_outputs(3438) <= a;
    layer5_outputs(3439) <= not a;
    layer5_outputs(3440) <= b and not a;
    layer5_outputs(3441) <= not (a and b);
    layer5_outputs(3442) <= not a;
    layer5_outputs(3443) <= not b;
    layer5_outputs(3444) <= not a or b;
    layer5_outputs(3445) <= b;
    layer5_outputs(3446) <= not (a or b);
    layer5_outputs(3447) <= b;
    layer5_outputs(3448) <= not (a and b);
    layer5_outputs(3449) <= not (a xor b);
    layer5_outputs(3450) <= a and b;
    layer5_outputs(3451) <= a and b;
    layer5_outputs(3452) <= a or b;
    layer5_outputs(3453) <= '1';
    layer5_outputs(3454) <= not b;
    layer5_outputs(3455) <= a and not b;
    layer5_outputs(3456) <= not a or b;
    layer5_outputs(3457) <= a xor b;
    layer5_outputs(3458) <= a and not b;
    layer5_outputs(3459) <= a and not b;
    layer5_outputs(3460) <= '1';
    layer5_outputs(3461) <= not a;
    layer5_outputs(3462) <= '0';
    layer5_outputs(3463) <= a or b;
    layer5_outputs(3464) <= not a or b;
    layer5_outputs(3465) <= a xor b;
    layer5_outputs(3466) <= not b or a;
    layer5_outputs(3467) <= '1';
    layer5_outputs(3468) <= not a or b;
    layer5_outputs(3469) <= a or b;
    layer5_outputs(3470) <= not b or a;
    layer5_outputs(3471) <= not (a xor b);
    layer5_outputs(3472) <= a or b;
    layer5_outputs(3473) <= not a or b;
    layer5_outputs(3474) <= not a;
    layer5_outputs(3475) <= a or b;
    layer5_outputs(3476) <= '0';
    layer5_outputs(3477) <= a and not b;
    layer5_outputs(3478) <= not b;
    layer5_outputs(3479) <= a;
    layer5_outputs(3480) <= b and not a;
    layer5_outputs(3481) <= b;
    layer5_outputs(3482) <= not (a and b);
    layer5_outputs(3483) <= not b or a;
    layer5_outputs(3484) <= not a;
    layer5_outputs(3485) <= not a;
    layer5_outputs(3486) <= b;
    layer5_outputs(3487) <= '0';
    layer5_outputs(3488) <= a or b;
    layer5_outputs(3489) <= b and not a;
    layer5_outputs(3490) <= b and not a;
    layer5_outputs(3491) <= not b;
    layer5_outputs(3492) <= not (a and b);
    layer5_outputs(3493) <= b;
    layer5_outputs(3494) <= not b;
    layer5_outputs(3495) <= a and not b;
    layer5_outputs(3496) <= not b;
    layer5_outputs(3497) <= '1';
    layer5_outputs(3498) <= a;
    layer5_outputs(3499) <= a or b;
    layer5_outputs(3500) <= '0';
    layer5_outputs(3501) <= '1';
    layer5_outputs(3502) <= not b;
    layer5_outputs(3503) <= not (a and b);
    layer5_outputs(3504) <= not b;
    layer5_outputs(3505) <= not (a and b);
    layer5_outputs(3506) <= a and b;
    layer5_outputs(3507) <= not b or a;
    layer5_outputs(3508) <= a or b;
    layer5_outputs(3509) <= a;
    layer5_outputs(3510) <= a xor b;
    layer5_outputs(3511) <= a and not b;
    layer5_outputs(3512) <= not a or b;
    layer5_outputs(3513) <= not b or a;
    layer5_outputs(3514) <= not a or b;
    layer5_outputs(3515) <= not b or a;
    layer5_outputs(3516) <= not b or a;
    layer5_outputs(3517) <= b and not a;
    layer5_outputs(3518) <= a or b;
    layer5_outputs(3519) <= not b or a;
    layer5_outputs(3520) <= a;
    layer5_outputs(3521) <= a and not b;
    layer5_outputs(3522) <= not a;
    layer5_outputs(3523) <= '1';
    layer5_outputs(3524) <= a xor b;
    layer5_outputs(3525) <= not a or b;
    layer5_outputs(3526) <= a and not b;
    layer5_outputs(3527) <= a or b;
    layer5_outputs(3528) <= a;
    layer5_outputs(3529) <= not a or b;
    layer5_outputs(3530) <= b;
    layer5_outputs(3531) <= a and not b;
    layer5_outputs(3532) <= not a or b;
    layer5_outputs(3533) <= not a or b;
    layer5_outputs(3534) <= a and b;
    layer5_outputs(3535) <= a;
    layer5_outputs(3536) <= b;
    layer5_outputs(3537) <= not (a or b);
    layer5_outputs(3538) <= b;
    layer5_outputs(3539) <= not b;
    layer5_outputs(3540) <= not b;
    layer5_outputs(3541) <= not (a and b);
    layer5_outputs(3542) <= a;
    layer5_outputs(3543) <= b;
    layer5_outputs(3544) <= not a;
    layer5_outputs(3545) <= not (a xor b);
    layer5_outputs(3546) <= not (a or b);
    layer5_outputs(3547) <= '1';
    layer5_outputs(3548) <= b and not a;
    layer5_outputs(3549) <= not a or b;
    layer5_outputs(3550) <= not (a or b);
    layer5_outputs(3551) <= not (a and b);
    layer5_outputs(3552) <= a or b;
    layer5_outputs(3553) <= not b or a;
    layer5_outputs(3554) <= a and not b;
    layer5_outputs(3555) <= not b or a;
    layer5_outputs(3556) <= a and b;
    layer5_outputs(3557) <= not a or b;
    layer5_outputs(3558) <= a and not b;
    layer5_outputs(3559) <= not (a and b);
    layer5_outputs(3560) <= a;
    layer5_outputs(3561) <= a and b;
    layer5_outputs(3562) <= b;
    layer5_outputs(3563) <= '1';
    layer5_outputs(3564) <= '1';
    layer5_outputs(3565) <= not (a and b);
    layer5_outputs(3566) <= a or b;
    layer5_outputs(3567) <= not b;
    layer5_outputs(3568) <= not a;
    layer5_outputs(3569) <= not a;
    layer5_outputs(3570) <= a xor b;
    layer5_outputs(3571) <= not a;
    layer5_outputs(3572) <= not b or a;
    layer5_outputs(3573) <= a and b;
    layer5_outputs(3574) <= not (a and b);
    layer5_outputs(3575) <= '0';
    layer5_outputs(3576) <= not a or b;
    layer5_outputs(3577) <= a and not b;
    layer5_outputs(3578) <= b;
    layer5_outputs(3579) <= b;
    layer5_outputs(3580) <= not a;
    layer5_outputs(3581) <= a and not b;
    layer5_outputs(3582) <= a;
    layer5_outputs(3583) <= a xor b;
    layer5_outputs(3584) <= not b or a;
    layer5_outputs(3585) <= b and not a;
    layer5_outputs(3586) <= not b or a;
    layer5_outputs(3587) <= not a;
    layer5_outputs(3588) <= not a;
    layer5_outputs(3589) <= a;
    layer5_outputs(3590) <= not a or b;
    layer5_outputs(3591) <= not b;
    layer5_outputs(3592) <= b and not a;
    layer5_outputs(3593) <= not (a and b);
    layer5_outputs(3594) <= not a or b;
    layer5_outputs(3595) <= a or b;
    layer5_outputs(3596) <= not a or b;
    layer5_outputs(3597) <= b;
    layer5_outputs(3598) <= a and b;
    layer5_outputs(3599) <= a or b;
    layer5_outputs(3600) <= b;
    layer5_outputs(3601) <= not (a xor b);
    layer5_outputs(3602) <= not (a and b);
    layer5_outputs(3603) <= not a;
    layer5_outputs(3604) <= b;
    layer5_outputs(3605) <= b;
    layer5_outputs(3606) <= not a or b;
    layer5_outputs(3607) <= not b;
    layer5_outputs(3608) <= a;
    layer5_outputs(3609) <= not b or a;
    layer5_outputs(3610) <= not b;
    layer5_outputs(3611) <= b and not a;
    layer5_outputs(3612) <= not (a or b);
    layer5_outputs(3613) <= a and not b;
    layer5_outputs(3614) <= not a;
    layer5_outputs(3615) <= a and not b;
    layer5_outputs(3616) <= b and not a;
    layer5_outputs(3617) <= not b or a;
    layer5_outputs(3618) <= not a;
    layer5_outputs(3619) <= a;
    layer5_outputs(3620) <= not (a or b);
    layer5_outputs(3621) <= not a;
    layer5_outputs(3622) <= b and not a;
    layer5_outputs(3623) <= not (a and b);
    layer5_outputs(3624) <= a xor b;
    layer5_outputs(3625) <= not b;
    layer5_outputs(3626) <= '1';
    layer5_outputs(3627) <= b and not a;
    layer5_outputs(3628) <= not (a and b);
    layer5_outputs(3629) <= not b;
    layer5_outputs(3630) <= b;
    layer5_outputs(3631) <= a or b;
    layer5_outputs(3632) <= a xor b;
    layer5_outputs(3633) <= not b;
    layer5_outputs(3634) <= not (a and b);
    layer5_outputs(3635) <= not b or a;
    layer5_outputs(3636) <= b;
    layer5_outputs(3637) <= not a or b;
    layer5_outputs(3638) <= a;
    layer5_outputs(3639) <= a or b;
    layer5_outputs(3640) <= a xor b;
    layer5_outputs(3641) <= a;
    layer5_outputs(3642) <= not b;
    layer5_outputs(3643) <= a;
    layer5_outputs(3644) <= a or b;
    layer5_outputs(3645) <= b;
    layer5_outputs(3646) <= a and b;
    layer5_outputs(3647) <= not (a or b);
    layer5_outputs(3648) <= b;
    layer5_outputs(3649) <= a;
    layer5_outputs(3650) <= not b or a;
    layer5_outputs(3651) <= a;
    layer5_outputs(3652) <= b;
    layer5_outputs(3653) <= b and not a;
    layer5_outputs(3654) <= '1';
    layer5_outputs(3655) <= not (a or b);
    layer5_outputs(3656) <= a and b;
    layer5_outputs(3657) <= not b or a;
    layer5_outputs(3658) <= a and b;
    layer5_outputs(3659) <= b and not a;
    layer5_outputs(3660) <= not (a and b);
    layer5_outputs(3661) <= a;
    layer5_outputs(3662) <= not a or b;
    layer5_outputs(3663) <= not a or b;
    layer5_outputs(3664) <= not a or b;
    layer5_outputs(3665) <= not (a or b);
    layer5_outputs(3666) <= a and not b;
    layer5_outputs(3667) <= '0';
    layer5_outputs(3668) <= not (a and b);
    layer5_outputs(3669) <= not (a and b);
    layer5_outputs(3670) <= '0';
    layer5_outputs(3671) <= a or b;
    layer5_outputs(3672) <= a or b;
    layer5_outputs(3673) <= '1';
    layer5_outputs(3674) <= '0';
    layer5_outputs(3675) <= not (a and b);
    layer5_outputs(3676) <= a and b;
    layer5_outputs(3677) <= not a;
    layer5_outputs(3678) <= not b;
    layer5_outputs(3679) <= not a or b;
    layer5_outputs(3680) <= not b;
    layer5_outputs(3681) <= b;
    layer5_outputs(3682) <= a and not b;
    layer5_outputs(3683) <= a or b;
    layer5_outputs(3684) <= a xor b;
    layer5_outputs(3685) <= not (a or b);
    layer5_outputs(3686) <= a and b;
    layer5_outputs(3687) <= a or b;
    layer5_outputs(3688) <= not a;
    layer5_outputs(3689) <= not a or b;
    layer5_outputs(3690) <= not b or a;
    layer5_outputs(3691) <= b and not a;
    layer5_outputs(3692) <= not b or a;
    layer5_outputs(3693) <= '1';
    layer5_outputs(3694) <= a and not b;
    layer5_outputs(3695) <= not b;
    layer5_outputs(3696) <= a xor b;
    layer5_outputs(3697) <= not a;
    layer5_outputs(3698) <= '1';
    layer5_outputs(3699) <= not (a xor b);
    layer5_outputs(3700) <= a and b;
    layer5_outputs(3701) <= not b or a;
    layer5_outputs(3702) <= not b or a;
    layer5_outputs(3703) <= a and not b;
    layer5_outputs(3704) <= a and not b;
    layer5_outputs(3705) <= a or b;
    layer5_outputs(3706) <= a xor b;
    layer5_outputs(3707) <= a;
    layer5_outputs(3708) <= a;
    layer5_outputs(3709) <= not (a and b);
    layer5_outputs(3710) <= a;
    layer5_outputs(3711) <= b;
    layer5_outputs(3712) <= b and not a;
    layer5_outputs(3713) <= b;
    layer5_outputs(3714) <= b;
    layer5_outputs(3715) <= not b or a;
    layer5_outputs(3716) <= a;
    layer5_outputs(3717) <= a;
    layer5_outputs(3718) <= a xor b;
    layer5_outputs(3719) <= not (a and b);
    layer5_outputs(3720) <= not (a xor b);
    layer5_outputs(3721) <= not (a xor b);
    layer5_outputs(3722) <= not (a or b);
    layer5_outputs(3723) <= b and not a;
    layer5_outputs(3724) <= not a;
    layer5_outputs(3725) <= a;
    layer5_outputs(3726) <= not (a or b);
    layer5_outputs(3727) <= not b or a;
    layer5_outputs(3728) <= not b;
    layer5_outputs(3729) <= b and not a;
    layer5_outputs(3730) <= not b;
    layer5_outputs(3731) <= a and b;
    layer5_outputs(3732) <= not a or b;
    layer5_outputs(3733) <= not (a xor b);
    layer5_outputs(3734) <= b and not a;
    layer5_outputs(3735) <= b;
    layer5_outputs(3736) <= a and not b;
    layer5_outputs(3737) <= a;
    layer5_outputs(3738) <= not b or a;
    layer5_outputs(3739) <= a or b;
    layer5_outputs(3740) <= not (a and b);
    layer5_outputs(3741) <= not (a and b);
    layer5_outputs(3742) <= '0';
    layer5_outputs(3743) <= a and not b;
    layer5_outputs(3744) <= not a or b;
    layer5_outputs(3745) <= b and not a;
    layer5_outputs(3746) <= not (a and b);
    layer5_outputs(3747) <= a;
    layer5_outputs(3748) <= not b or a;
    layer5_outputs(3749) <= a and not b;
    layer5_outputs(3750) <= not a or b;
    layer5_outputs(3751) <= not b or a;
    layer5_outputs(3752) <= a;
    layer5_outputs(3753) <= a or b;
    layer5_outputs(3754) <= '1';
    layer5_outputs(3755) <= not b;
    layer5_outputs(3756) <= not (a and b);
    layer5_outputs(3757) <= not (a or b);
    layer5_outputs(3758) <= b;
    layer5_outputs(3759) <= not a;
    layer5_outputs(3760) <= b;
    layer5_outputs(3761) <= a xor b;
    layer5_outputs(3762) <= a;
    layer5_outputs(3763) <= a and not b;
    layer5_outputs(3764) <= not (a and b);
    layer5_outputs(3765) <= a;
    layer5_outputs(3766) <= not (a xor b);
    layer5_outputs(3767) <= not (a or b);
    layer5_outputs(3768) <= b and not a;
    layer5_outputs(3769) <= a;
    layer5_outputs(3770) <= not b or a;
    layer5_outputs(3771) <= not a or b;
    layer5_outputs(3772) <= not a or b;
    layer5_outputs(3773) <= not (a and b);
    layer5_outputs(3774) <= not b;
    layer5_outputs(3775) <= b;
    layer5_outputs(3776) <= not a;
    layer5_outputs(3777) <= a and not b;
    layer5_outputs(3778) <= not b;
    layer5_outputs(3779) <= not a;
    layer5_outputs(3780) <= not a;
    layer5_outputs(3781) <= not b;
    layer5_outputs(3782) <= b;
    layer5_outputs(3783) <= not (a xor b);
    layer5_outputs(3784) <= not (a or b);
    layer5_outputs(3785) <= a;
    layer5_outputs(3786) <= a or b;
    layer5_outputs(3787) <= not a or b;
    layer5_outputs(3788) <= not (a and b);
    layer5_outputs(3789) <= a and not b;
    layer5_outputs(3790) <= '1';
    layer5_outputs(3791) <= a xor b;
    layer5_outputs(3792) <= not b or a;
    layer5_outputs(3793) <= a and not b;
    layer5_outputs(3794) <= a;
    layer5_outputs(3795) <= not a;
    layer5_outputs(3796) <= not b;
    layer5_outputs(3797) <= not a;
    layer5_outputs(3798) <= a and not b;
    layer5_outputs(3799) <= not a;
    layer5_outputs(3800) <= not a;
    layer5_outputs(3801) <= not b;
    layer5_outputs(3802) <= b and not a;
    layer5_outputs(3803) <= a xor b;
    layer5_outputs(3804) <= not a or b;
    layer5_outputs(3805) <= not (a or b);
    layer5_outputs(3806) <= not (a and b);
    layer5_outputs(3807) <= b;
    layer5_outputs(3808) <= a or b;
    layer5_outputs(3809) <= not a or b;
    layer5_outputs(3810) <= a and b;
    layer5_outputs(3811) <= not (a xor b);
    layer5_outputs(3812) <= a xor b;
    layer5_outputs(3813) <= b and not a;
    layer5_outputs(3814) <= b;
    layer5_outputs(3815) <= not (a and b);
    layer5_outputs(3816) <= b;
    layer5_outputs(3817) <= a or b;
    layer5_outputs(3818) <= '0';
    layer5_outputs(3819) <= a or b;
    layer5_outputs(3820) <= '0';
    layer5_outputs(3821) <= '0';
    layer5_outputs(3822) <= not a or b;
    layer5_outputs(3823) <= a and not b;
    layer5_outputs(3824) <= not b or a;
    layer5_outputs(3825) <= b and not a;
    layer5_outputs(3826) <= '1';
    layer5_outputs(3827) <= b and not a;
    layer5_outputs(3828) <= b and not a;
    layer5_outputs(3829) <= b;
    layer5_outputs(3830) <= not (a and b);
    layer5_outputs(3831) <= not a or b;
    layer5_outputs(3832) <= not b;
    layer5_outputs(3833) <= a or b;
    layer5_outputs(3834) <= a and b;
    layer5_outputs(3835) <= not a or b;
    layer5_outputs(3836) <= not a;
    layer5_outputs(3837) <= a or b;
    layer5_outputs(3838) <= not (a or b);
    layer5_outputs(3839) <= not (a and b);
    layer5_outputs(3840) <= b;
    layer5_outputs(3841) <= b;
    layer5_outputs(3842) <= b and not a;
    layer5_outputs(3843) <= a and b;
    layer5_outputs(3844) <= a and b;
    layer5_outputs(3845) <= b;
    layer5_outputs(3846) <= not a;
    layer5_outputs(3847) <= not (a or b);
    layer5_outputs(3848) <= b and not a;
    layer5_outputs(3849) <= not b;
    layer5_outputs(3850) <= b;
    layer5_outputs(3851) <= a;
    layer5_outputs(3852) <= not b;
    layer5_outputs(3853) <= not b or a;
    layer5_outputs(3854) <= not (a and b);
    layer5_outputs(3855) <= a and b;
    layer5_outputs(3856) <= not (a or b);
    layer5_outputs(3857) <= a and b;
    layer5_outputs(3858) <= a or b;
    layer5_outputs(3859) <= not a or b;
    layer5_outputs(3860) <= not (a or b);
    layer5_outputs(3861) <= '1';
    layer5_outputs(3862) <= a;
    layer5_outputs(3863) <= a;
    layer5_outputs(3864) <= '1';
    layer5_outputs(3865) <= '0';
    layer5_outputs(3866) <= b and not a;
    layer5_outputs(3867) <= a;
    layer5_outputs(3868) <= b and not a;
    layer5_outputs(3869) <= not (a or b);
    layer5_outputs(3870) <= '1';
    layer5_outputs(3871) <= not b;
    layer5_outputs(3872) <= a or b;
    layer5_outputs(3873) <= not b;
    layer5_outputs(3874) <= b;
    layer5_outputs(3875) <= a and not b;
    layer5_outputs(3876) <= not (a and b);
    layer5_outputs(3877) <= a;
    layer5_outputs(3878) <= a and b;
    layer5_outputs(3879) <= a and not b;
    layer5_outputs(3880) <= a and not b;
    layer5_outputs(3881) <= not (a xor b);
    layer5_outputs(3882) <= a or b;
    layer5_outputs(3883) <= not (a and b);
    layer5_outputs(3884) <= not (a and b);
    layer5_outputs(3885) <= not a or b;
    layer5_outputs(3886) <= a and b;
    layer5_outputs(3887) <= a and not b;
    layer5_outputs(3888) <= a or b;
    layer5_outputs(3889) <= not b;
    layer5_outputs(3890) <= not a;
    layer5_outputs(3891) <= not (a or b);
    layer5_outputs(3892) <= a and b;
    layer5_outputs(3893) <= '0';
    layer5_outputs(3894) <= a and not b;
    layer5_outputs(3895) <= b and not a;
    layer5_outputs(3896) <= '1';
    layer5_outputs(3897) <= a;
    layer5_outputs(3898) <= a;
    layer5_outputs(3899) <= not b;
    layer5_outputs(3900) <= '1';
    layer5_outputs(3901) <= a;
    layer5_outputs(3902) <= b;
    layer5_outputs(3903) <= not (a xor b);
    layer5_outputs(3904) <= a or b;
    layer5_outputs(3905) <= a xor b;
    layer5_outputs(3906) <= not (a and b);
    layer5_outputs(3907) <= b;
    layer5_outputs(3908) <= not a;
    layer5_outputs(3909) <= a;
    layer5_outputs(3910) <= b and not a;
    layer5_outputs(3911) <= not (a and b);
    layer5_outputs(3912) <= '1';
    layer5_outputs(3913) <= not (a xor b);
    layer5_outputs(3914) <= not a;
    layer5_outputs(3915) <= '0';
    layer5_outputs(3916) <= a and b;
    layer5_outputs(3917) <= not b;
    layer5_outputs(3918) <= b;
    layer5_outputs(3919) <= a;
    layer5_outputs(3920) <= a and not b;
    layer5_outputs(3921) <= not a or b;
    layer5_outputs(3922) <= not b or a;
    layer5_outputs(3923) <= not (a xor b);
    layer5_outputs(3924) <= '1';
    layer5_outputs(3925) <= a or b;
    layer5_outputs(3926) <= not (a and b);
    layer5_outputs(3927) <= '0';
    layer5_outputs(3928) <= a and not b;
    layer5_outputs(3929) <= not (a xor b);
    layer5_outputs(3930) <= not b;
    layer5_outputs(3931) <= a;
    layer5_outputs(3932) <= a xor b;
    layer5_outputs(3933) <= '0';
    layer5_outputs(3934) <= a and not b;
    layer5_outputs(3935) <= not b;
    layer5_outputs(3936) <= a and not b;
    layer5_outputs(3937) <= a and not b;
    layer5_outputs(3938) <= not b or a;
    layer5_outputs(3939) <= b;
    layer5_outputs(3940) <= '0';
    layer5_outputs(3941) <= not b or a;
    layer5_outputs(3942) <= not (a or b);
    layer5_outputs(3943) <= not a or b;
    layer5_outputs(3944) <= '1';
    layer5_outputs(3945) <= not (a and b);
    layer5_outputs(3946) <= '1';
    layer5_outputs(3947) <= a and b;
    layer5_outputs(3948) <= not (a or b);
    layer5_outputs(3949) <= not (a or b);
    layer5_outputs(3950) <= b and not a;
    layer5_outputs(3951) <= not b or a;
    layer5_outputs(3952) <= a and b;
    layer5_outputs(3953) <= not a or b;
    layer5_outputs(3954) <= '0';
    layer5_outputs(3955) <= not b;
    layer5_outputs(3956) <= not (a xor b);
    layer5_outputs(3957) <= not (a and b);
    layer5_outputs(3958) <= a and b;
    layer5_outputs(3959) <= not (a or b);
    layer5_outputs(3960) <= not (a or b);
    layer5_outputs(3961) <= '1';
    layer5_outputs(3962) <= not b or a;
    layer5_outputs(3963) <= a;
    layer5_outputs(3964) <= not a;
    layer5_outputs(3965) <= not a or b;
    layer5_outputs(3966) <= b and not a;
    layer5_outputs(3967) <= not (a and b);
    layer5_outputs(3968) <= a;
    layer5_outputs(3969) <= not a;
    layer5_outputs(3970) <= a;
    layer5_outputs(3971) <= not b;
    layer5_outputs(3972) <= b and not a;
    layer5_outputs(3973) <= a and not b;
    layer5_outputs(3974) <= a and not b;
    layer5_outputs(3975) <= not b;
    layer5_outputs(3976) <= not a;
    layer5_outputs(3977) <= not b or a;
    layer5_outputs(3978) <= not a or b;
    layer5_outputs(3979) <= '0';
    layer5_outputs(3980) <= b and not a;
    layer5_outputs(3981) <= not b or a;
    layer5_outputs(3982) <= a;
    layer5_outputs(3983) <= not b;
    layer5_outputs(3984) <= '0';
    layer5_outputs(3985) <= not (a xor b);
    layer5_outputs(3986) <= a;
    layer5_outputs(3987) <= not a;
    layer5_outputs(3988) <= not b or a;
    layer5_outputs(3989) <= a and not b;
    layer5_outputs(3990) <= a;
    layer5_outputs(3991) <= b;
    layer5_outputs(3992) <= '1';
    layer5_outputs(3993) <= '1';
    layer5_outputs(3994) <= not (a xor b);
    layer5_outputs(3995) <= not b;
    layer5_outputs(3996) <= a or b;
    layer5_outputs(3997) <= a and b;
    layer5_outputs(3998) <= not b or a;
    layer5_outputs(3999) <= a and not b;
    layer5_outputs(4000) <= not b;
    layer5_outputs(4001) <= '1';
    layer5_outputs(4002) <= not a or b;
    layer5_outputs(4003) <= a and b;
    layer5_outputs(4004) <= a;
    layer5_outputs(4005) <= b;
    layer5_outputs(4006) <= not (a or b);
    layer5_outputs(4007) <= a xor b;
    layer5_outputs(4008) <= '1';
    layer5_outputs(4009) <= not a or b;
    layer5_outputs(4010) <= a or b;
    layer5_outputs(4011) <= not (a and b);
    layer5_outputs(4012) <= a and b;
    layer5_outputs(4013) <= '1';
    layer5_outputs(4014) <= a and not b;
    layer5_outputs(4015) <= b;
    layer5_outputs(4016) <= a;
    layer5_outputs(4017) <= not b;
    layer5_outputs(4018) <= not b;
    layer5_outputs(4019) <= not a;
    layer5_outputs(4020) <= not b;
    layer5_outputs(4021) <= b and not a;
    layer5_outputs(4022) <= not (a or b);
    layer5_outputs(4023) <= a;
    layer5_outputs(4024) <= not b;
    layer5_outputs(4025) <= not (a and b);
    layer5_outputs(4026) <= a or b;
    layer5_outputs(4027) <= not a or b;
    layer5_outputs(4028) <= '0';
    layer5_outputs(4029) <= a and not b;
    layer5_outputs(4030) <= not a;
    layer5_outputs(4031) <= a xor b;
    layer5_outputs(4032) <= a and not b;
    layer5_outputs(4033) <= not a;
    layer5_outputs(4034) <= not b;
    layer5_outputs(4035) <= a and not b;
    layer5_outputs(4036) <= '1';
    layer5_outputs(4037) <= a and not b;
    layer5_outputs(4038) <= not a or b;
    layer5_outputs(4039) <= a and not b;
    layer5_outputs(4040) <= a xor b;
    layer5_outputs(4041) <= not a or b;
    layer5_outputs(4042) <= b and not a;
    layer5_outputs(4043) <= a and b;
    layer5_outputs(4044) <= not a;
    layer5_outputs(4045) <= not (a and b);
    layer5_outputs(4046) <= a xor b;
    layer5_outputs(4047) <= b and not a;
    layer5_outputs(4048) <= b and not a;
    layer5_outputs(4049) <= not b or a;
    layer5_outputs(4050) <= not a or b;
    layer5_outputs(4051) <= a and not b;
    layer5_outputs(4052) <= a and not b;
    layer5_outputs(4053) <= not (a and b);
    layer5_outputs(4054) <= not (a or b);
    layer5_outputs(4055) <= not a or b;
    layer5_outputs(4056) <= a;
    layer5_outputs(4057) <= b;
    layer5_outputs(4058) <= '1';
    layer5_outputs(4059) <= not (a xor b);
    layer5_outputs(4060) <= b;
    layer5_outputs(4061) <= not a;
    layer5_outputs(4062) <= '0';
    layer5_outputs(4063) <= not (a or b);
    layer5_outputs(4064) <= b and not a;
    layer5_outputs(4065) <= '0';
    layer5_outputs(4066) <= a and not b;
    layer5_outputs(4067) <= a;
    layer5_outputs(4068) <= a;
    layer5_outputs(4069) <= b and not a;
    layer5_outputs(4070) <= not (a or b);
    layer5_outputs(4071) <= not (a xor b);
    layer5_outputs(4072) <= not b;
    layer5_outputs(4073) <= not (a or b);
    layer5_outputs(4074) <= a and not b;
    layer5_outputs(4075) <= '0';
    layer5_outputs(4076) <= not (a or b);
    layer5_outputs(4077) <= b;
    layer5_outputs(4078) <= b and not a;
    layer5_outputs(4079) <= b;
    layer5_outputs(4080) <= a and b;
    layer5_outputs(4081) <= not b or a;
    layer5_outputs(4082) <= not b;
    layer5_outputs(4083) <= b;
    layer5_outputs(4084) <= a;
    layer5_outputs(4085) <= a xor b;
    layer5_outputs(4086) <= not a or b;
    layer5_outputs(4087) <= a and not b;
    layer5_outputs(4088) <= a and b;
    layer5_outputs(4089) <= not (a and b);
    layer5_outputs(4090) <= a and b;
    layer5_outputs(4091) <= b;
    layer5_outputs(4092) <= not b or a;
    layer5_outputs(4093) <= '1';
    layer5_outputs(4094) <= not a;
    layer5_outputs(4095) <= b;
    layer5_outputs(4096) <= b;
    layer5_outputs(4097) <= not a or b;
    layer5_outputs(4098) <= a;
    layer5_outputs(4099) <= not a;
    layer5_outputs(4100) <= not a or b;
    layer5_outputs(4101) <= not (a or b);
    layer5_outputs(4102) <= not b or a;
    layer5_outputs(4103) <= not b;
    layer5_outputs(4104) <= b and not a;
    layer5_outputs(4105) <= b;
    layer5_outputs(4106) <= a and not b;
    layer5_outputs(4107) <= b and not a;
    layer5_outputs(4108) <= b;
    layer5_outputs(4109) <= not b;
    layer5_outputs(4110) <= b and not a;
    layer5_outputs(4111) <= a or b;
    layer5_outputs(4112) <= a;
    layer5_outputs(4113) <= not a;
    layer5_outputs(4114) <= not (a or b);
    layer5_outputs(4115) <= a and not b;
    layer5_outputs(4116) <= not a;
    layer5_outputs(4117) <= a and b;
    layer5_outputs(4118) <= not a;
    layer5_outputs(4119) <= b;
    layer5_outputs(4120) <= a;
    layer5_outputs(4121) <= not a;
    layer5_outputs(4122) <= a;
    layer5_outputs(4123) <= not a or b;
    layer5_outputs(4124) <= a and b;
    layer5_outputs(4125) <= not a;
    layer5_outputs(4126) <= '0';
    layer5_outputs(4127) <= a and b;
    layer5_outputs(4128) <= a or b;
    layer5_outputs(4129) <= not (a xor b);
    layer5_outputs(4130) <= not a or b;
    layer5_outputs(4131) <= not a;
    layer5_outputs(4132) <= a xor b;
    layer5_outputs(4133) <= not b or a;
    layer5_outputs(4134) <= not b or a;
    layer5_outputs(4135) <= a and b;
    layer5_outputs(4136) <= not (a xor b);
    layer5_outputs(4137) <= a or b;
    layer5_outputs(4138) <= a;
    layer5_outputs(4139) <= a and not b;
    layer5_outputs(4140) <= b;
    layer5_outputs(4141) <= not a;
    layer5_outputs(4142) <= a;
    layer5_outputs(4143) <= not b;
    layer5_outputs(4144) <= '1';
    layer5_outputs(4145) <= a;
    layer5_outputs(4146) <= not b or a;
    layer5_outputs(4147) <= a or b;
    layer5_outputs(4148) <= not b or a;
    layer5_outputs(4149) <= not b;
    layer5_outputs(4150) <= a and b;
    layer5_outputs(4151) <= not b;
    layer5_outputs(4152) <= a and b;
    layer5_outputs(4153) <= b and not a;
    layer5_outputs(4154) <= '1';
    layer5_outputs(4155) <= a and b;
    layer5_outputs(4156) <= b;
    layer5_outputs(4157) <= a;
    layer5_outputs(4158) <= a or b;
    layer5_outputs(4159) <= not a;
    layer5_outputs(4160) <= not b or a;
    layer5_outputs(4161) <= a and b;
    layer5_outputs(4162) <= not b;
    layer5_outputs(4163) <= not b or a;
    layer5_outputs(4164) <= '1';
    layer5_outputs(4165) <= not (a or b);
    layer5_outputs(4166) <= '0';
    layer5_outputs(4167) <= a and b;
    layer5_outputs(4168) <= b;
    layer5_outputs(4169) <= '0';
    layer5_outputs(4170) <= not b or a;
    layer5_outputs(4171) <= not a;
    layer5_outputs(4172) <= not a;
    layer5_outputs(4173) <= not b or a;
    layer5_outputs(4174) <= not (a and b);
    layer5_outputs(4175) <= a or b;
    layer5_outputs(4176) <= b;
    layer5_outputs(4177) <= '1';
    layer5_outputs(4178) <= not a;
    layer5_outputs(4179) <= b and not a;
    layer5_outputs(4180) <= a xor b;
    layer5_outputs(4181) <= b and not a;
    layer5_outputs(4182) <= b;
    layer5_outputs(4183) <= a or b;
    layer5_outputs(4184) <= a;
    layer5_outputs(4185) <= not b or a;
    layer5_outputs(4186) <= a or b;
    layer5_outputs(4187) <= a and not b;
    layer5_outputs(4188) <= not a or b;
    layer5_outputs(4189) <= b;
    layer5_outputs(4190) <= not (a xor b);
    layer5_outputs(4191) <= a and not b;
    layer5_outputs(4192) <= not a;
    layer5_outputs(4193) <= not b or a;
    layer5_outputs(4194) <= not (a and b);
    layer5_outputs(4195) <= not b or a;
    layer5_outputs(4196) <= a and not b;
    layer5_outputs(4197) <= b;
    layer5_outputs(4198) <= b and not a;
    layer5_outputs(4199) <= a or b;
    layer5_outputs(4200) <= not b or a;
    layer5_outputs(4201) <= not b;
    layer5_outputs(4202) <= not (a and b);
    layer5_outputs(4203) <= not a;
    layer5_outputs(4204) <= not b;
    layer5_outputs(4205) <= not (a or b);
    layer5_outputs(4206) <= not b or a;
    layer5_outputs(4207) <= '1';
    layer5_outputs(4208) <= a and b;
    layer5_outputs(4209) <= not b;
    layer5_outputs(4210) <= not (a or b);
    layer5_outputs(4211) <= not (a xor b);
    layer5_outputs(4212) <= not b;
    layer5_outputs(4213) <= not (a or b);
    layer5_outputs(4214) <= not (a and b);
    layer5_outputs(4215) <= not (a or b);
    layer5_outputs(4216) <= a or b;
    layer5_outputs(4217) <= not a or b;
    layer5_outputs(4218) <= not b or a;
    layer5_outputs(4219) <= not a;
    layer5_outputs(4220) <= not b or a;
    layer5_outputs(4221) <= a;
    layer5_outputs(4222) <= b and not a;
    layer5_outputs(4223) <= b and not a;
    layer5_outputs(4224) <= a or b;
    layer5_outputs(4225) <= b;
    layer5_outputs(4226) <= a and not b;
    layer5_outputs(4227) <= not b;
    layer5_outputs(4228) <= not a;
    layer5_outputs(4229) <= not a or b;
    layer5_outputs(4230) <= a or b;
    layer5_outputs(4231) <= a or b;
    layer5_outputs(4232) <= not a;
    layer5_outputs(4233) <= a and not b;
    layer5_outputs(4234) <= not a;
    layer5_outputs(4235) <= '0';
    layer5_outputs(4236) <= a and b;
    layer5_outputs(4237) <= a or b;
    layer5_outputs(4238) <= a xor b;
    layer5_outputs(4239) <= a and not b;
    layer5_outputs(4240) <= not (a xor b);
    layer5_outputs(4241) <= not (a or b);
    layer5_outputs(4242) <= '0';
    layer5_outputs(4243) <= not b;
    layer5_outputs(4244) <= a;
    layer5_outputs(4245) <= a and b;
    layer5_outputs(4246) <= a;
    layer5_outputs(4247) <= a;
    layer5_outputs(4248) <= not b;
    layer5_outputs(4249) <= not (a and b);
    layer5_outputs(4250) <= not a or b;
    layer5_outputs(4251) <= not (a and b);
    layer5_outputs(4252) <= not a;
    layer5_outputs(4253) <= not b;
    layer5_outputs(4254) <= not b or a;
    layer5_outputs(4255) <= not a;
    layer5_outputs(4256) <= b;
    layer5_outputs(4257) <= a;
    layer5_outputs(4258) <= a and not b;
    layer5_outputs(4259) <= not a;
    layer5_outputs(4260) <= not (a and b);
    layer5_outputs(4261) <= a and b;
    layer5_outputs(4262) <= a;
    layer5_outputs(4263) <= not b;
    layer5_outputs(4264) <= not (a and b);
    layer5_outputs(4265) <= b;
    layer5_outputs(4266) <= not a or b;
    layer5_outputs(4267) <= not (a and b);
    layer5_outputs(4268) <= not (a and b);
    layer5_outputs(4269) <= a xor b;
    layer5_outputs(4270) <= not b;
    layer5_outputs(4271) <= b and not a;
    layer5_outputs(4272) <= '0';
    layer5_outputs(4273) <= b;
    layer5_outputs(4274) <= not (a xor b);
    layer5_outputs(4275) <= not b;
    layer5_outputs(4276) <= '0';
    layer5_outputs(4277) <= a and b;
    layer5_outputs(4278) <= not a;
    layer5_outputs(4279) <= not (a and b);
    layer5_outputs(4280) <= not a or b;
    layer5_outputs(4281) <= a and b;
    layer5_outputs(4282) <= b and not a;
    layer5_outputs(4283) <= not b;
    layer5_outputs(4284) <= a or b;
    layer5_outputs(4285) <= a xor b;
    layer5_outputs(4286) <= '0';
    layer5_outputs(4287) <= b and not a;
    layer5_outputs(4288) <= not b or a;
    layer5_outputs(4289) <= a;
    layer5_outputs(4290) <= b and not a;
    layer5_outputs(4291) <= not b;
    layer5_outputs(4292) <= a or b;
    layer5_outputs(4293) <= a;
    layer5_outputs(4294) <= not b;
    layer5_outputs(4295) <= b;
    layer5_outputs(4296) <= not a;
    layer5_outputs(4297) <= a or b;
    layer5_outputs(4298) <= not a;
    layer5_outputs(4299) <= a xor b;
    layer5_outputs(4300) <= not b;
    layer5_outputs(4301) <= not (a and b);
    layer5_outputs(4302) <= a;
    layer5_outputs(4303) <= b and not a;
    layer5_outputs(4304) <= b;
    layer5_outputs(4305) <= b and not a;
    layer5_outputs(4306) <= a xor b;
    layer5_outputs(4307) <= '1';
    layer5_outputs(4308) <= not b;
    layer5_outputs(4309) <= not a;
    layer5_outputs(4310) <= a;
    layer5_outputs(4311) <= a;
    layer5_outputs(4312) <= b and not a;
    layer5_outputs(4313) <= a or b;
    layer5_outputs(4314) <= not (a and b);
    layer5_outputs(4315) <= not b;
    layer5_outputs(4316) <= '1';
    layer5_outputs(4317) <= not (a xor b);
    layer5_outputs(4318) <= not b or a;
    layer5_outputs(4319) <= not b;
    layer5_outputs(4320) <= a or b;
    layer5_outputs(4321) <= a and not b;
    layer5_outputs(4322) <= not b;
    layer5_outputs(4323) <= not (a xor b);
    layer5_outputs(4324) <= a;
    layer5_outputs(4325) <= a or b;
    layer5_outputs(4326) <= a xor b;
    layer5_outputs(4327) <= not b or a;
    layer5_outputs(4328) <= not a;
    layer5_outputs(4329) <= a;
    layer5_outputs(4330) <= '0';
    layer5_outputs(4331) <= a;
    layer5_outputs(4332) <= not b;
    layer5_outputs(4333) <= a or b;
    layer5_outputs(4334) <= a;
    layer5_outputs(4335) <= not (a xor b);
    layer5_outputs(4336) <= not (a or b);
    layer5_outputs(4337) <= b;
    layer5_outputs(4338) <= '0';
    layer5_outputs(4339) <= not a;
    layer5_outputs(4340) <= a;
    layer5_outputs(4341) <= a xor b;
    layer5_outputs(4342) <= not a or b;
    layer5_outputs(4343) <= not b or a;
    layer5_outputs(4344) <= a;
    layer5_outputs(4345) <= a or b;
    layer5_outputs(4346) <= not (a and b);
    layer5_outputs(4347) <= b;
    layer5_outputs(4348) <= not a or b;
    layer5_outputs(4349) <= a or b;
    layer5_outputs(4350) <= not (a xor b);
    layer5_outputs(4351) <= b and not a;
    layer5_outputs(4352) <= not (a xor b);
    layer5_outputs(4353) <= b;
    layer5_outputs(4354) <= not a;
    layer5_outputs(4355) <= a and not b;
    layer5_outputs(4356) <= b;
    layer5_outputs(4357) <= '1';
    layer5_outputs(4358) <= not b;
    layer5_outputs(4359) <= not (a and b);
    layer5_outputs(4360) <= a or b;
    layer5_outputs(4361) <= not (a or b);
    layer5_outputs(4362) <= not b;
    layer5_outputs(4363) <= not (a or b);
    layer5_outputs(4364) <= b and not a;
    layer5_outputs(4365) <= a and b;
    layer5_outputs(4366) <= b;
    layer5_outputs(4367) <= not b;
    layer5_outputs(4368) <= a and b;
    layer5_outputs(4369) <= not a;
    layer5_outputs(4370) <= not a;
    layer5_outputs(4371) <= a and not b;
    layer5_outputs(4372) <= b and not a;
    layer5_outputs(4373) <= a or b;
    layer5_outputs(4374) <= a or b;
    layer5_outputs(4375) <= a or b;
    layer5_outputs(4376) <= b;
    layer5_outputs(4377) <= not (a or b);
    layer5_outputs(4378) <= '0';
    layer5_outputs(4379) <= not b;
    layer5_outputs(4380) <= not (a and b);
    layer5_outputs(4381) <= a;
    layer5_outputs(4382) <= a;
    layer5_outputs(4383) <= not (a and b);
    layer5_outputs(4384) <= not a;
    layer5_outputs(4385) <= a;
    layer5_outputs(4386) <= not b;
    layer5_outputs(4387) <= b;
    layer5_outputs(4388) <= b;
    layer5_outputs(4389) <= a and not b;
    layer5_outputs(4390) <= a;
    layer5_outputs(4391) <= b;
    layer5_outputs(4392) <= not b;
    layer5_outputs(4393) <= '0';
    layer5_outputs(4394) <= a or b;
    layer5_outputs(4395) <= not (a and b);
    layer5_outputs(4396) <= not b or a;
    layer5_outputs(4397) <= a or b;
    layer5_outputs(4398) <= a and not b;
    layer5_outputs(4399) <= not (a or b);
    layer5_outputs(4400) <= a and not b;
    layer5_outputs(4401) <= not b;
    layer5_outputs(4402) <= a;
    layer5_outputs(4403) <= a;
    layer5_outputs(4404) <= not (a and b);
    layer5_outputs(4405) <= b;
    layer5_outputs(4406) <= not (a and b);
    layer5_outputs(4407) <= not (a or b);
    layer5_outputs(4408) <= not a or b;
    layer5_outputs(4409) <= a xor b;
    layer5_outputs(4410) <= not a or b;
    layer5_outputs(4411) <= a xor b;
    layer5_outputs(4412) <= a or b;
    layer5_outputs(4413) <= a;
    layer5_outputs(4414) <= not (a and b);
    layer5_outputs(4415) <= b and not a;
    layer5_outputs(4416) <= a and b;
    layer5_outputs(4417) <= b;
    layer5_outputs(4418) <= not (a xor b);
    layer5_outputs(4419) <= not (a and b);
    layer5_outputs(4420) <= not b or a;
    layer5_outputs(4421) <= not (a or b);
    layer5_outputs(4422) <= a and b;
    layer5_outputs(4423) <= '1';
    layer5_outputs(4424) <= a and not b;
    layer5_outputs(4425) <= a xor b;
    layer5_outputs(4426) <= not (a and b);
    layer5_outputs(4427) <= not a;
    layer5_outputs(4428) <= b and not a;
    layer5_outputs(4429) <= '0';
    layer5_outputs(4430) <= not b;
    layer5_outputs(4431) <= a;
    layer5_outputs(4432) <= a or b;
    layer5_outputs(4433) <= a or b;
    layer5_outputs(4434) <= b;
    layer5_outputs(4435) <= a;
    layer5_outputs(4436) <= not a;
    layer5_outputs(4437) <= not b or a;
    layer5_outputs(4438) <= b and not a;
    layer5_outputs(4439) <= not (a or b);
    layer5_outputs(4440) <= not (a or b);
    layer5_outputs(4441) <= not (a or b);
    layer5_outputs(4442) <= a and b;
    layer5_outputs(4443) <= a;
    layer5_outputs(4444) <= not (a or b);
    layer5_outputs(4445) <= b and not a;
    layer5_outputs(4446) <= a;
    layer5_outputs(4447) <= not (a and b);
    layer5_outputs(4448) <= not a or b;
    layer5_outputs(4449) <= a or b;
    layer5_outputs(4450) <= not b;
    layer5_outputs(4451) <= not a or b;
    layer5_outputs(4452) <= not (a or b);
    layer5_outputs(4453) <= a and b;
    layer5_outputs(4454) <= not b;
    layer5_outputs(4455) <= not b;
    layer5_outputs(4456) <= a and not b;
    layer5_outputs(4457) <= not b;
    layer5_outputs(4458) <= not (a xor b);
    layer5_outputs(4459) <= a;
    layer5_outputs(4460) <= a;
    layer5_outputs(4461) <= a and not b;
    layer5_outputs(4462) <= b;
    layer5_outputs(4463) <= not (a or b);
    layer5_outputs(4464) <= a and not b;
    layer5_outputs(4465) <= a xor b;
    layer5_outputs(4466) <= not a;
    layer5_outputs(4467) <= b;
    layer5_outputs(4468) <= not a;
    layer5_outputs(4469) <= '0';
    layer5_outputs(4470) <= not b or a;
    layer5_outputs(4471) <= a xor b;
    layer5_outputs(4472) <= a;
    layer5_outputs(4473) <= '1';
    layer5_outputs(4474) <= not a;
    layer5_outputs(4475) <= a;
    layer5_outputs(4476) <= a and not b;
    layer5_outputs(4477) <= b;
    layer5_outputs(4478) <= b;
    layer5_outputs(4479) <= '0';
    layer5_outputs(4480) <= not (a and b);
    layer5_outputs(4481) <= not a or b;
    layer5_outputs(4482) <= b and not a;
    layer5_outputs(4483) <= not (a and b);
    layer5_outputs(4484) <= not b or a;
    layer5_outputs(4485) <= a or b;
    layer5_outputs(4486) <= not b;
    layer5_outputs(4487) <= '1';
    layer5_outputs(4488) <= not b;
    layer5_outputs(4489) <= a;
    layer5_outputs(4490) <= not (a and b);
    layer5_outputs(4491) <= b;
    layer5_outputs(4492) <= not (a or b);
    layer5_outputs(4493) <= not a;
    layer5_outputs(4494) <= '0';
    layer5_outputs(4495) <= '0';
    layer5_outputs(4496) <= b;
    layer5_outputs(4497) <= a or b;
    layer5_outputs(4498) <= not (a xor b);
    layer5_outputs(4499) <= b;
    layer5_outputs(4500) <= not a;
    layer5_outputs(4501) <= '1';
    layer5_outputs(4502) <= a or b;
    layer5_outputs(4503) <= b;
    layer5_outputs(4504) <= not a;
    layer5_outputs(4505) <= a;
    layer5_outputs(4506) <= a or b;
    layer5_outputs(4507) <= not a;
    layer5_outputs(4508) <= a;
    layer5_outputs(4509) <= a and b;
    layer5_outputs(4510) <= not (a xor b);
    layer5_outputs(4511) <= a xor b;
    layer5_outputs(4512) <= a xor b;
    layer5_outputs(4513) <= a;
    layer5_outputs(4514) <= not b;
    layer5_outputs(4515) <= a xor b;
    layer5_outputs(4516) <= not a;
    layer5_outputs(4517) <= not a or b;
    layer5_outputs(4518) <= b and not a;
    layer5_outputs(4519) <= a;
    layer5_outputs(4520) <= a xor b;
    layer5_outputs(4521) <= a or b;
    layer5_outputs(4522) <= not b or a;
    layer5_outputs(4523) <= not a;
    layer5_outputs(4524) <= '1';
    layer5_outputs(4525) <= not a;
    layer5_outputs(4526) <= not b or a;
    layer5_outputs(4527) <= a;
    layer5_outputs(4528) <= not a;
    layer5_outputs(4529) <= a;
    layer5_outputs(4530) <= '0';
    layer5_outputs(4531) <= a;
    layer5_outputs(4532) <= b and not a;
    layer5_outputs(4533) <= not a;
    layer5_outputs(4534) <= '1';
    layer5_outputs(4535) <= a and b;
    layer5_outputs(4536) <= a;
    layer5_outputs(4537) <= b;
    layer5_outputs(4538) <= a and not b;
    layer5_outputs(4539) <= a;
    layer5_outputs(4540) <= a;
    layer5_outputs(4541) <= b;
    layer5_outputs(4542) <= not b;
    layer5_outputs(4543) <= a;
    layer5_outputs(4544) <= b and not a;
    layer5_outputs(4545) <= not b or a;
    layer5_outputs(4546) <= not a or b;
    layer5_outputs(4547) <= b and not a;
    layer5_outputs(4548) <= a and not b;
    layer5_outputs(4549) <= '1';
    layer5_outputs(4550) <= not a or b;
    layer5_outputs(4551) <= not b;
    layer5_outputs(4552) <= not a;
    layer5_outputs(4553) <= a;
    layer5_outputs(4554) <= not a;
    layer5_outputs(4555) <= not (a and b);
    layer5_outputs(4556) <= not (a xor b);
    layer5_outputs(4557) <= b;
    layer5_outputs(4558) <= b;
    layer5_outputs(4559) <= b;
    layer5_outputs(4560) <= not (a xor b);
    layer5_outputs(4561) <= b;
    layer5_outputs(4562) <= not (a and b);
    layer5_outputs(4563) <= '1';
    layer5_outputs(4564) <= not b or a;
    layer5_outputs(4565) <= not a;
    layer5_outputs(4566) <= '0';
    layer5_outputs(4567) <= a or b;
    layer5_outputs(4568) <= not a or b;
    layer5_outputs(4569) <= not (a xor b);
    layer5_outputs(4570) <= not b;
    layer5_outputs(4571) <= not a or b;
    layer5_outputs(4572) <= a;
    layer5_outputs(4573) <= a;
    layer5_outputs(4574) <= a xor b;
    layer5_outputs(4575) <= b;
    layer5_outputs(4576) <= not a;
    layer5_outputs(4577) <= not (a or b);
    layer5_outputs(4578) <= a;
    layer5_outputs(4579) <= a or b;
    layer5_outputs(4580) <= b and not a;
    layer5_outputs(4581) <= a and b;
    layer5_outputs(4582) <= a;
    layer5_outputs(4583) <= not b;
    layer5_outputs(4584) <= a xor b;
    layer5_outputs(4585) <= a or b;
    layer5_outputs(4586) <= a or b;
    layer5_outputs(4587) <= not a;
    layer5_outputs(4588) <= not a;
    layer5_outputs(4589) <= not (a or b);
    layer5_outputs(4590) <= not b;
    layer5_outputs(4591) <= not (a or b);
    layer5_outputs(4592) <= a and not b;
    layer5_outputs(4593) <= not (a and b);
    layer5_outputs(4594) <= not b or a;
    layer5_outputs(4595) <= a and b;
    layer5_outputs(4596) <= b and not a;
    layer5_outputs(4597) <= not b;
    layer5_outputs(4598) <= not a or b;
    layer5_outputs(4599) <= '0';
    layer5_outputs(4600) <= not a;
    layer5_outputs(4601) <= not a or b;
    layer5_outputs(4602) <= a or b;
    layer5_outputs(4603) <= not (a or b);
    layer5_outputs(4604) <= a or b;
    layer5_outputs(4605) <= not (a xor b);
    layer5_outputs(4606) <= b and not a;
    layer5_outputs(4607) <= not (a and b);
    layer5_outputs(4608) <= not a or b;
    layer5_outputs(4609) <= '1';
    layer5_outputs(4610) <= a;
    layer5_outputs(4611) <= a and b;
    layer5_outputs(4612) <= not a;
    layer5_outputs(4613) <= not (a xor b);
    layer5_outputs(4614) <= a;
    layer5_outputs(4615) <= '0';
    layer5_outputs(4616) <= not (a xor b);
    layer5_outputs(4617) <= a xor b;
    layer5_outputs(4618) <= not b;
    layer5_outputs(4619) <= a and b;
    layer5_outputs(4620) <= not a or b;
    layer5_outputs(4621) <= not a or b;
    layer5_outputs(4622) <= not b;
    layer5_outputs(4623) <= a and b;
    layer5_outputs(4624) <= '1';
    layer5_outputs(4625) <= not b;
    layer5_outputs(4626) <= b and not a;
    layer5_outputs(4627) <= not a or b;
    layer5_outputs(4628) <= not (a xor b);
    layer5_outputs(4629) <= not a;
    layer5_outputs(4630) <= '0';
    layer5_outputs(4631) <= not a or b;
    layer5_outputs(4632) <= not (a xor b);
    layer5_outputs(4633) <= b;
    layer5_outputs(4634) <= b and not a;
    layer5_outputs(4635) <= not a or b;
    layer5_outputs(4636) <= not a;
    layer5_outputs(4637) <= not a;
    layer5_outputs(4638) <= not a;
    layer5_outputs(4639) <= a and b;
    layer5_outputs(4640) <= a and not b;
    layer5_outputs(4641) <= '1';
    layer5_outputs(4642) <= not a or b;
    layer5_outputs(4643) <= a;
    layer5_outputs(4644) <= not b or a;
    layer5_outputs(4645) <= a;
    layer5_outputs(4646) <= not (a and b);
    layer5_outputs(4647) <= not b;
    layer5_outputs(4648) <= a;
    layer5_outputs(4649) <= a or b;
    layer5_outputs(4650) <= not (a or b);
    layer5_outputs(4651) <= not b or a;
    layer5_outputs(4652) <= a;
    layer5_outputs(4653) <= not a or b;
    layer5_outputs(4654) <= not (a xor b);
    layer5_outputs(4655) <= a;
    layer5_outputs(4656) <= a and not b;
    layer5_outputs(4657) <= b and not a;
    layer5_outputs(4658) <= b and not a;
    layer5_outputs(4659) <= b;
    layer5_outputs(4660) <= a;
    layer5_outputs(4661) <= b and not a;
    layer5_outputs(4662) <= not a;
    layer5_outputs(4663) <= a and not b;
    layer5_outputs(4664) <= '0';
    layer5_outputs(4665) <= a and not b;
    layer5_outputs(4666) <= not b or a;
    layer5_outputs(4667) <= '1';
    layer5_outputs(4668) <= a and not b;
    layer5_outputs(4669) <= b and not a;
    layer5_outputs(4670) <= not b;
    layer5_outputs(4671) <= not b or a;
    layer5_outputs(4672) <= a or b;
    layer5_outputs(4673) <= b;
    layer5_outputs(4674) <= a or b;
    layer5_outputs(4675) <= a;
    layer5_outputs(4676) <= a and not b;
    layer5_outputs(4677) <= not a;
    layer5_outputs(4678) <= not (a and b);
    layer5_outputs(4679) <= not a;
    layer5_outputs(4680) <= not a or b;
    layer5_outputs(4681) <= not (a or b);
    layer5_outputs(4682) <= '0';
    layer5_outputs(4683) <= not a;
    layer5_outputs(4684) <= not b;
    layer5_outputs(4685) <= a and not b;
    layer5_outputs(4686) <= '0';
    layer5_outputs(4687) <= not b or a;
    layer5_outputs(4688) <= not a;
    layer5_outputs(4689) <= '1';
    layer5_outputs(4690) <= a xor b;
    layer5_outputs(4691) <= a;
    layer5_outputs(4692) <= not b;
    layer5_outputs(4693) <= not b;
    layer5_outputs(4694) <= b and not a;
    layer5_outputs(4695) <= a or b;
    layer5_outputs(4696) <= not (a or b);
    layer5_outputs(4697) <= not a;
    layer5_outputs(4698) <= a and not b;
    layer5_outputs(4699) <= not a or b;
    layer5_outputs(4700) <= b and not a;
    layer5_outputs(4701) <= a;
    layer5_outputs(4702) <= not a;
    layer5_outputs(4703) <= not b;
    layer5_outputs(4704) <= not (a xor b);
    layer5_outputs(4705) <= not a or b;
    layer5_outputs(4706) <= a and not b;
    layer5_outputs(4707) <= not (a or b);
    layer5_outputs(4708) <= not a or b;
    layer5_outputs(4709) <= not b or a;
    layer5_outputs(4710) <= a and not b;
    layer5_outputs(4711) <= b and not a;
    layer5_outputs(4712) <= a;
    layer5_outputs(4713) <= a xor b;
    layer5_outputs(4714) <= not (a or b);
    layer5_outputs(4715) <= a and not b;
    layer5_outputs(4716) <= a and not b;
    layer5_outputs(4717) <= not a;
    layer5_outputs(4718) <= a and b;
    layer5_outputs(4719) <= not b;
    layer5_outputs(4720) <= not a or b;
    layer5_outputs(4721) <= not (a and b);
    layer5_outputs(4722) <= a and b;
    layer5_outputs(4723) <= '0';
    layer5_outputs(4724) <= '1';
    layer5_outputs(4725) <= a and not b;
    layer5_outputs(4726) <= '1';
    layer5_outputs(4727) <= not b;
    layer5_outputs(4728) <= '1';
    layer5_outputs(4729) <= not a;
    layer5_outputs(4730) <= not (a and b);
    layer5_outputs(4731) <= not (a xor b);
    layer5_outputs(4732) <= not a or b;
    layer5_outputs(4733) <= '0';
    layer5_outputs(4734) <= a;
    layer5_outputs(4735) <= b;
    layer5_outputs(4736) <= not (a and b);
    layer5_outputs(4737) <= not a;
    layer5_outputs(4738) <= not a;
    layer5_outputs(4739) <= not a or b;
    layer5_outputs(4740) <= not (a xor b);
    layer5_outputs(4741) <= a or b;
    layer5_outputs(4742) <= not a or b;
    layer5_outputs(4743) <= a or b;
    layer5_outputs(4744) <= not b;
    layer5_outputs(4745) <= not a or b;
    layer5_outputs(4746) <= not (a or b);
    layer5_outputs(4747) <= not b;
    layer5_outputs(4748) <= b and not a;
    layer5_outputs(4749) <= not a or b;
    layer5_outputs(4750) <= not (a or b);
    layer5_outputs(4751) <= not a;
    layer5_outputs(4752) <= not (a and b);
    layer5_outputs(4753) <= a xor b;
    layer5_outputs(4754) <= not (a or b);
    layer5_outputs(4755) <= a and not b;
    layer5_outputs(4756) <= not (a and b);
    layer5_outputs(4757) <= a;
    layer5_outputs(4758) <= b and not a;
    layer5_outputs(4759) <= '0';
    layer5_outputs(4760) <= not (a or b);
    layer5_outputs(4761) <= a;
    layer5_outputs(4762) <= '1';
    layer5_outputs(4763) <= a or b;
    layer5_outputs(4764) <= '0';
    layer5_outputs(4765) <= a and not b;
    layer5_outputs(4766) <= not a or b;
    layer5_outputs(4767) <= not a;
    layer5_outputs(4768) <= b and not a;
    layer5_outputs(4769) <= b;
    layer5_outputs(4770) <= '1';
    layer5_outputs(4771) <= a;
    layer5_outputs(4772) <= '0';
    layer5_outputs(4773) <= '1';
    layer5_outputs(4774) <= not b or a;
    layer5_outputs(4775) <= not a or b;
    layer5_outputs(4776) <= '1';
    layer5_outputs(4777) <= b;
    layer5_outputs(4778) <= a;
    layer5_outputs(4779) <= not (a xor b);
    layer5_outputs(4780) <= a xor b;
    layer5_outputs(4781) <= '0';
    layer5_outputs(4782) <= not (a xor b);
    layer5_outputs(4783) <= a and not b;
    layer5_outputs(4784) <= not a;
    layer5_outputs(4785) <= not (a and b);
    layer5_outputs(4786) <= a or b;
    layer5_outputs(4787) <= not a;
    layer5_outputs(4788) <= a;
    layer5_outputs(4789) <= not (a or b);
    layer5_outputs(4790) <= '1';
    layer5_outputs(4791) <= not (a and b);
    layer5_outputs(4792) <= b and not a;
    layer5_outputs(4793) <= not b or a;
    layer5_outputs(4794) <= not b;
    layer5_outputs(4795) <= a;
    layer5_outputs(4796) <= not (a and b);
    layer5_outputs(4797) <= a or b;
    layer5_outputs(4798) <= not a;
    layer5_outputs(4799) <= b and not a;
    layer5_outputs(4800) <= not (a or b);
    layer5_outputs(4801) <= b;
    layer5_outputs(4802) <= a xor b;
    layer5_outputs(4803) <= not a or b;
    layer5_outputs(4804) <= a;
    layer5_outputs(4805) <= a and b;
    layer5_outputs(4806) <= not b;
    layer5_outputs(4807) <= not (a and b);
    layer5_outputs(4808) <= not b;
    layer5_outputs(4809) <= a;
    layer5_outputs(4810) <= a xor b;
    layer5_outputs(4811) <= a and b;
    layer5_outputs(4812) <= a;
    layer5_outputs(4813) <= b and not a;
    layer5_outputs(4814) <= b;
    layer5_outputs(4815) <= '1';
    layer5_outputs(4816) <= not a;
    layer5_outputs(4817) <= not b;
    layer5_outputs(4818) <= a xor b;
    layer5_outputs(4819) <= not (a or b);
    layer5_outputs(4820) <= not a;
    layer5_outputs(4821) <= not b or a;
    layer5_outputs(4822) <= not b;
    layer5_outputs(4823) <= b;
    layer5_outputs(4824) <= a;
    layer5_outputs(4825) <= a xor b;
    layer5_outputs(4826) <= b and not a;
    layer5_outputs(4827) <= not (a and b);
    layer5_outputs(4828) <= not (a and b);
    layer5_outputs(4829) <= not (a and b);
    layer5_outputs(4830) <= b and not a;
    layer5_outputs(4831) <= b and not a;
    layer5_outputs(4832) <= not a;
    layer5_outputs(4833) <= '1';
    layer5_outputs(4834) <= '0';
    layer5_outputs(4835) <= '0';
    layer5_outputs(4836) <= not (a xor b);
    layer5_outputs(4837) <= not a or b;
    layer5_outputs(4838) <= a and b;
    layer5_outputs(4839) <= not a;
    layer5_outputs(4840) <= b;
    layer5_outputs(4841) <= b and not a;
    layer5_outputs(4842) <= not b;
    layer5_outputs(4843) <= not b or a;
    layer5_outputs(4844) <= not (a and b);
    layer5_outputs(4845) <= not (a xor b);
    layer5_outputs(4846) <= '0';
    layer5_outputs(4847) <= not b;
    layer5_outputs(4848) <= a;
    layer5_outputs(4849) <= a and not b;
    layer5_outputs(4850) <= not a or b;
    layer5_outputs(4851) <= not a or b;
    layer5_outputs(4852) <= '1';
    layer5_outputs(4853) <= a or b;
    layer5_outputs(4854) <= '1';
    layer5_outputs(4855) <= not a;
    layer5_outputs(4856) <= b;
    layer5_outputs(4857) <= not a;
    layer5_outputs(4858) <= a;
    layer5_outputs(4859) <= '0';
    layer5_outputs(4860) <= not a;
    layer5_outputs(4861) <= a and b;
    layer5_outputs(4862) <= b;
    layer5_outputs(4863) <= not b;
    layer5_outputs(4864) <= not (a and b);
    layer5_outputs(4865) <= b;
    layer5_outputs(4866) <= b and not a;
    layer5_outputs(4867) <= not b;
    layer5_outputs(4868) <= a and b;
    layer5_outputs(4869) <= a;
    layer5_outputs(4870) <= '0';
    layer5_outputs(4871) <= a;
    layer5_outputs(4872) <= not b;
    layer5_outputs(4873) <= not b;
    layer5_outputs(4874) <= b;
    layer5_outputs(4875) <= '1';
    layer5_outputs(4876) <= not a;
    layer5_outputs(4877) <= not b;
    layer5_outputs(4878) <= not (a xor b);
    layer5_outputs(4879) <= a;
    layer5_outputs(4880) <= b;
    layer5_outputs(4881) <= not (a or b);
    layer5_outputs(4882) <= b and not a;
    layer5_outputs(4883) <= not a;
    layer5_outputs(4884) <= not (a or b);
    layer5_outputs(4885) <= not b or a;
    layer5_outputs(4886) <= a xor b;
    layer5_outputs(4887) <= a or b;
    layer5_outputs(4888) <= not b or a;
    layer5_outputs(4889) <= a or b;
    layer5_outputs(4890) <= not a;
    layer5_outputs(4891) <= not a;
    layer5_outputs(4892) <= a and not b;
    layer5_outputs(4893) <= not b;
    layer5_outputs(4894) <= a and not b;
    layer5_outputs(4895) <= a;
    layer5_outputs(4896) <= not (a or b);
    layer5_outputs(4897) <= not b;
    layer5_outputs(4898) <= a;
    layer5_outputs(4899) <= b;
    layer5_outputs(4900) <= a and b;
    layer5_outputs(4901) <= a;
    layer5_outputs(4902) <= b and not a;
    layer5_outputs(4903) <= not (a and b);
    layer5_outputs(4904) <= not b;
    layer5_outputs(4905) <= not (a and b);
    layer5_outputs(4906) <= a and not b;
    layer5_outputs(4907) <= not a;
    layer5_outputs(4908) <= b;
    layer5_outputs(4909) <= not a;
    layer5_outputs(4910) <= b and not a;
    layer5_outputs(4911) <= not b;
    layer5_outputs(4912) <= a;
    layer5_outputs(4913) <= not (a xor b);
    layer5_outputs(4914) <= not (a or b);
    layer5_outputs(4915) <= a;
    layer5_outputs(4916) <= b;
    layer5_outputs(4917) <= a xor b;
    layer5_outputs(4918) <= a and not b;
    layer5_outputs(4919) <= b;
    layer5_outputs(4920) <= not (a or b);
    layer5_outputs(4921) <= a and b;
    layer5_outputs(4922) <= not a;
    layer5_outputs(4923) <= not (a or b);
    layer5_outputs(4924) <= a xor b;
    layer5_outputs(4925) <= not (a and b);
    layer5_outputs(4926) <= a or b;
    layer5_outputs(4927) <= a;
    layer5_outputs(4928) <= not b or a;
    layer5_outputs(4929) <= not a;
    layer5_outputs(4930) <= a and not b;
    layer5_outputs(4931) <= a and b;
    layer5_outputs(4932) <= not (a xor b);
    layer5_outputs(4933) <= b and not a;
    layer5_outputs(4934) <= b;
    layer5_outputs(4935) <= b and not a;
    layer5_outputs(4936) <= '0';
    layer5_outputs(4937) <= a or b;
    layer5_outputs(4938) <= a xor b;
    layer5_outputs(4939) <= not (a xor b);
    layer5_outputs(4940) <= not a;
    layer5_outputs(4941) <= a or b;
    layer5_outputs(4942) <= not a;
    layer5_outputs(4943) <= a and b;
    layer5_outputs(4944) <= a or b;
    layer5_outputs(4945) <= not b;
    layer5_outputs(4946) <= a xor b;
    layer5_outputs(4947) <= a and b;
    layer5_outputs(4948) <= not b;
    layer5_outputs(4949) <= b;
    layer5_outputs(4950) <= a;
    layer5_outputs(4951) <= a and not b;
    layer5_outputs(4952) <= not (a xor b);
    layer5_outputs(4953) <= not a or b;
    layer5_outputs(4954) <= not a or b;
    layer5_outputs(4955) <= not b or a;
    layer5_outputs(4956) <= not a;
    layer5_outputs(4957) <= b and not a;
    layer5_outputs(4958) <= not (a and b);
    layer5_outputs(4959) <= '0';
    layer5_outputs(4960) <= not b;
    layer5_outputs(4961) <= not (a or b);
    layer5_outputs(4962) <= a xor b;
    layer5_outputs(4963) <= a and not b;
    layer5_outputs(4964) <= not b or a;
    layer5_outputs(4965) <= not b or a;
    layer5_outputs(4966) <= not b;
    layer5_outputs(4967) <= not b or a;
    layer5_outputs(4968) <= '1';
    layer5_outputs(4969) <= a and not b;
    layer5_outputs(4970) <= a and b;
    layer5_outputs(4971) <= a and b;
    layer5_outputs(4972) <= not a;
    layer5_outputs(4973) <= not a;
    layer5_outputs(4974) <= a;
    layer5_outputs(4975) <= b and not a;
    layer5_outputs(4976) <= not a or b;
    layer5_outputs(4977) <= not a or b;
    layer5_outputs(4978) <= b;
    layer5_outputs(4979) <= a and b;
    layer5_outputs(4980) <= b;
    layer5_outputs(4981) <= a;
    layer5_outputs(4982) <= b;
    layer5_outputs(4983) <= a xor b;
    layer5_outputs(4984) <= not a or b;
    layer5_outputs(4985) <= not a;
    layer5_outputs(4986) <= not a or b;
    layer5_outputs(4987) <= not b;
    layer5_outputs(4988) <= a;
    layer5_outputs(4989) <= '1';
    layer5_outputs(4990) <= not b;
    layer5_outputs(4991) <= not b or a;
    layer5_outputs(4992) <= not b;
    layer5_outputs(4993) <= not (a or b);
    layer5_outputs(4994) <= not a or b;
    layer5_outputs(4995) <= a and b;
    layer5_outputs(4996) <= b and not a;
    layer5_outputs(4997) <= not (a or b);
    layer5_outputs(4998) <= b;
    layer5_outputs(4999) <= '0';
    layer5_outputs(5000) <= not (a or b);
    layer5_outputs(5001) <= a or b;
    layer5_outputs(5002) <= not a or b;
    layer5_outputs(5003) <= not (a and b);
    layer5_outputs(5004) <= '1';
    layer5_outputs(5005) <= a and not b;
    layer5_outputs(5006) <= a;
    layer5_outputs(5007) <= not (a xor b);
    layer5_outputs(5008) <= '0';
    layer5_outputs(5009) <= not (a and b);
    layer5_outputs(5010) <= not (a and b);
    layer5_outputs(5011) <= a xor b;
    layer5_outputs(5012) <= a and b;
    layer5_outputs(5013) <= not (a xor b);
    layer5_outputs(5014) <= b and not a;
    layer5_outputs(5015) <= not (a or b);
    layer5_outputs(5016) <= not (a or b);
    layer5_outputs(5017) <= not (a xor b);
    layer5_outputs(5018) <= a or b;
    layer5_outputs(5019) <= a or b;
    layer5_outputs(5020) <= not b or a;
    layer5_outputs(5021) <= a and b;
    layer5_outputs(5022) <= '0';
    layer5_outputs(5023) <= a or b;
    layer5_outputs(5024) <= a and b;
    layer5_outputs(5025) <= a;
    layer5_outputs(5026) <= a;
    layer5_outputs(5027) <= b and not a;
    layer5_outputs(5028) <= a and b;
    layer5_outputs(5029) <= '1';
    layer5_outputs(5030) <= '0';
    layer5_outputs(5031) <= a and not b;
    layer5_outputs(5032) <= a;
    layer5_outputs(5033) <= a or b;
    layer5_outputs(5034) <= not (a xor b);
    layer5_outputs(5035) <= not b or a;
    layer5_outputs(5036) <= '1';
    layer5_outputs(5037) <= b;
    layer5_outputs(5038) <= not b or a;
    layer5_outputs(5039) <= b;
    layer5_outputs(5040) <= b;
    layer5_outputs(5041) <= a or b;
    layer5_outputs(5042) <= not a;
    layer5_outputs(5043) <= a or b;
    layer5_outputs(5044) <= a and b;
    layer5_outputs(5045) <= a or b;
    layer5_outputs(5046) <= a;
    layer5_outputs(5047) <= not b;
    layer5_outputs(5048) <= a or b;
    layer5_outputs(5049) <= b;
    layer5_outputs(5050) <= not a;
    layer5_outputs(5051) <= not (a xor b);
    layer5_outputs(5052) <= '0';
    layer5_outputs(5053) <= a;
    layer5_outputs(5054) <= a;
    layer5_outputs(5055) <= not b;
    layer5_outputs(5056) <= a;
    layer5_outputs(5057) <= not a;
    layer5_outputs(5058) <= not a or b;
    layer5_outputs(5059) <= not b;
    layer5_outputs(5060) <= a and b;
    layer5_outputs(5061) <= b and not a;
    layer5_outputs(5062) <= a and not b;
    layer5_outputs(5063) <= not (a and b);
    layer5_outputs(5064) <= '1';
    layer5_outputs(5065) <= not b or a;
    layer5_outputs(5066) <= a;
    layer5_outputs(5067) <= not (a xor b);
    layer5_outputs(5068) <= a;
    layer5_outputs(5069) <= a or b;
    layer5_outputs(5070) <= '0';
    layer5_outputs(5071) <= b;
    layer5_outputs(5072) <= a and b;
    layer5_outputs(5073) <= not a;
    layer5_outputs(5074) <= b;
    layer5_outputs(5075) <= not b or a;
    layer5_outputs(5076) <= not b or a;
    layer5_outputs(5077) <= not a;
    layer5_outputs(5078) <= '0';
    layer5_outputs(5079) <= b and not a;
    layer5_outputs(5080) <= '0';
    layer5_outputs(5081) <= a and b;
    layer5_outputs(5082) <= not b;
    layer5_outputs(5083) <= not b;
    layer5_outputs(5084) <= not a;
    layer5_outputs(5085) <= a or b;
    layer5_outputs(5086) <= not b;
    layer5_outputs(5087) <= b;
    layer5_outputs(5088) <= '1';
    layer5_outputs(5089) <= b and not a;
    layer5_outputs(5090) <= a or b;
    layer5_outputs(5091) <= not b;
    layer5_outputs(5092) <= a and not b;
    layer5_outputs(5093) <= not b;
    layer5_outputs(5094) <= b and not a;
    layer5_outputs(5095) <= a;
    layer5_outputs(5096) <= b and not a;
    layer5_outputs(5097) <= not a or b;
    layer5_outputs(5098) <= a or b;
    layer5_outputs(5099) <= not b;
    layer5_outputs(5100) <= b and not a;
    layer5_outputs(5101) <= a or b;
    layer5_outputs(5102) <= a;
    layer5_outputs(5103) <= not (a or b);
    layer5_outputs(5104) <= b;
    layer5_outputs(5105) <= not b or a;
    layer5_outputs(5106) <= a or b;
    layer5_outputs(5107) <= a or b;
    layer5_outputs(5108) <= a;
    layer5_outputs(5109) <= b and not a;
    layer5_outputs(5110) <= b;
    layer5_outputs(5111) <= b and not a;
    layer5_outputs(5112) <= not b or a;
    layer5_outputs(5113) <= a and not b;
    layer5_outputs(5114) <= b;
    layer5_outputs(5115) <= b;
    layer5_outputs(5116) <= a or b;
    layer5_outputs(5117) <= not b;
    layer5_outputs(5118) <= a;
    layer5_outputs(5119) <= a;
    layer5_outputs(5120) <= not a;
    layer5_outputs(5121) <= '0';
    layer5_outputs(5122) <= a;
    layer5_outputs(5123) <= not b or a;
    layer5_outputs(5124) <= b;
    layer5_outputs(5125) <= not (a and b);
    layer5_outputs(5126) <= b and not a;
    layer5_outputs(5127) <= not b or a;
    layer5_outputs(5128) <= not a;
    layer5_outputs(5129) <= '0';
    layer5_outputs(5130) <= not b;
    layer5_outputs(5131) <= not a;
    layer5_outputs(5132) <= a and b;
    layer5_outputs(5133) <= '1';
    layer5_outputs(5134) <= '0';
    layer5_outputs(5135) <= b;
    layer5_outputs(5136) <= not b;
    layer5_outputs(5137) <= not a;
    layer5_outputs(5138) <= not (a and b);
    layer5_outputs(5139) <= not b;
    layer5_outputs(5140) <= not (a xor b);
    layer5_outputs(5141) <= b and not a;
    layer5_outputs(5142) <= a;
    layer5_outputs(5143) <= not (a and b);
    layer5_outputs(5144) <= not (a or b);
    layer5_outputs(5145) <= not b or a;
    layer5_outputs(5146) <= b;
    layer5_outputs(5147) <= not b;
    layer5_outputs(5148) <= not b or a;
    layer5_outputs(5149) <= b;
    layer5_outputs(5150) <= b;
    layer5_outputs(5151) <= not (a xor b);
    layer5_outputs(5152) <= not b;
    layer5_outputs(5153) <= not b;
    layer5_outputs(5154) <= not (a and b);
    layer5_outputs(5155) <= a and not b;
    layer5_outputs(5156) <= '1';
    layer5_outputs(5157) <= not (a or b);
    layer5_outputs(5158) <= not b;
    layer5_outputs(5159) <= not a;
    layer5_outputs(5160) <= not a;
    layer5_outputs(5161) <= a;
    layer5_outputs(5162) <= not (a or b);
    layer5_outputs(5163) <= not b;
    layer5_outputs(5164) <= not a or b;
    layer5_outputs(5165) <= b;
    layer5_outputs(5166) <= not a;
    layer5_outputs(5167) <= not b;
    layer5_outputs(5168) <= not b or a;
    layer5_outputs(5169) <= b;
    layer5_outputs(5170) <= not a;
    layer5_outputs(5171) <= b and not a;
    layer5_outputs(5172) <= '1';
    layer5_outputs(5173) <= a or b;
    layer5_outputs(5174) <= b;
    layer5_outputs(5175) <= '0';
    layer5_outputs(5176) <= a;
    layer5_outputs(5177) <= b;
    layer5_outputs(5178) <= not b;
    layer5_outputs(5179) <= not b or a;
    layer5_outputs(5180) <= a and b;
    layer5_outputs(5181) <= a and b;
    layer5_outputs(5182) <= not (a or b);
    layer5_outputs(5183) <= not a;
    layer5_outputs(5184) <= not (a or b);
    layer5_outputs(5185) <= not a or b;
    layer5_outputs(5186) <= not b or a;
    layer5_outputs(5187) <= '0';
    layer5_outputs(5188) <= not a;
    layer5_outputs(5189) <= not (a and b);
    layer5_outputs(5190) <= not b or a;
    layer5_outputs(5191) <= '0';
    layer5_outputs(5192) <= not b or a;
    layer5_outputs(5193) <= a and not b;
    layer5_outputs(5194) <= not a;
    layer5_outputs(5195) <= a;
    layer5_outputs(5196) <= not b;
    layer5_outputs(5197) <= '0';
    layer5_outputs(5198) <= not (a and b);
    layer5_outputs(5199) <= not b or a;
    layer5_outputs(5200) <= not b;
    layer5_outputs(5201) <= not (a xor b);
    layer5_outputs(5202) <= not b;
    layer5_outputs(5203) <= a;
    layer5_outputs(5204) <= b;
    layer5_outputs(5205) <= not (a or b);
    layer5_outputs(5206) <= not a;
    layer5_outputs(5207) <= a xor b;
    layer5_outputs(5208) <= not b;
    layer5_outputs(5209) <= not (a and b);
    layer5_outputs(5210) <= not b;
    layer5_outputs(5211) <= a;
    layer5_outputs(5212) <= a;
    layer5_outputs(5213) <= not a or b;
    layer5_outputs(5214) <= not (a and b);
    layer5_outputs(5215) <= not (a xor b);
    layer5_outputs(5216) <= b;
    layer5_outputs(5217) <= '0';
    layer5_outputs(5218) <= a or b;
    layer5_outputs(5219) <= b;
    layer5_outputs(5220) <= a;
    layer5_outputs(5221) <= not a;
    layer5_outputs(5222) <= not (a or b);
    layer5_outputs(5223) <= not (a and b);
    layer5_outputs(5224) <= b;
    layer5_outputs(5225) <= not (a or b);
    layer5_outputs(5226) <= not (a or b);
    layer5_outputs(5227) <= a and b;
    layer5_outputs(5228) <= a and b;
    layer5_outputs(5229) <= a and b;
    layer5_outputs(5230) <= b;
    layer5_outputs(5231) <= not a;
    layer5_outputs(5232) <= b;
    layer5_outputs(5233) <= not a or b;
    layer5_outputs(5234) <= not (a and b);
    layer5_outputs(5235) <= a or b;
    layer5_outputs(5236) <= not a or b;
    layer5_outputs(5237) <= a and b;
    layer5_outputs(5238) <= not (a or b);
    layer5_outputs(5239) <= not b;
    layer5_outputs(5240) <= a and not b;
    layer5_outputs(5241) <= '0';
    layer5_outputs(5242) <= not a;
    layer5_outputs(5243) <= a xor b;
    layer5_outputs(5244) <= a and b;
    layer5_outputs(5245) <= a and b;
    layer5_outputs(5246) <= not a or b;
    layer5_outputs(5247) <= a or b;
    layer5_outputs(5248) <= a or b;
    layer5_outputs(5249) <= not a;
    layer5_outputs(5250) <= not a or b;
    layer5_outputs(5251) <= b and not a;
    layer5_outputs(5252) <= a;
    layer5_outputs(5253) <= not (a and b);
    layer5_outputs(5254) <= a or b;
    layer5_outputs(5255) <= not (a and b);
    layer5_outputs(5256) <= a;
    layer5_outputs(5257) <= not b;
    layer5_outputs(5258) <= a and b;
    layer5_outputs(5259) <= not a;
    layer5_outputs(5260) <= b;
    layer5_outputs(5261) <= not (a xor b);
    layer5_outputs(5262) <= not b or a;
    layer5_outputs(5263) <= b;
    layer5_outputs(5264) <= b;
    layer5_outputs(5265) <= not a;
    layer5_outputs(5266) <= not (a or b);
    layer5_outputs(5267) <= a and not b;
    layer5_outputs(5268) <= not b;
    layer5_outputs(5269) <= not (a or b);
    layer5_outputs(5270) <= a or b;
    layer5_outputs(5271) <= '1';
    layer5_outputs(5272) <= b;
    layer5_outputs(5273) <= b;
    layer5_outputs(5274) <= a and not b;
    layer5_outputs(5275) <= '0';
    layer5_outputs(5276) <= not a;
    layer5_outputs(5277) <= not a or b;
    layer5_outputs(5278) <= '1';
    layer5_outputs(5279) <= b;
    layer5_outputs(5280) <= not b or a;
    layer5_outputs(5281) <= b and not a;
    layer5_outputs(5282) <= a and not b;
    layer5_outputs(5283) <= not a;
    layer5_outputs(5284) <= b and not a;
    layer5_outputs(5285) <= a and not b;
    layer5_outputs(5286) <= not (a and b);
    layer5_outputs(5287) <= a and b;
    layer5_outputs(5288) <= not (a or b);
    layer5_outputs(5289) <= a xor b;
    layer5_outputs(5290) <= b;
    layer5_outputs(5291) <= not a;
    layer5_outputs(5292) <= not a;
    layer5_outputs(5293) <= not a;
    layer5_outputs(5294) <= not a;
    layer5_outputs(5295) <= not a;
    layer5_outputs(5296) <= a;
    layer5_outputs(5297) <= a or b;
    layer5_outputs(5298) <= a or b;
    layer5_outputs(5299) <= not a;
    layer5_outputs(5300) <= not a;
    layer5_outputs(5301) <= a;
    layer5_outputs(5302) <= a xor b;
    layer5_outputs(5303) <= a or b;
    layer5_outputs(5304) <= a;
    layer5_outputs(5305) <= not b or a;
    layer5_outputs(5306) <= not (a xor b);
    layer5_outputs(5307) <= not a;
    layer5_outputs(5308) <= a;
    layer5_outputs(5309) <= not (a and b);
    layer5_outputs(5310) <= a or b;
    layer5_outputs(5311) <= a and not b;
    layer5_outputs(5312) <= a;
    layer5_outputs(5313) <= a and not b;
    layer5_outputs(5314) <= not a;
    layer5_outputs(5315) <= not a;
    layer5_outputs(5316) <= not b or a;
    layer5_outputs(5317) <= not a;
    layer5_outputs(5318) <= a xor b;
    layer5_outputs(5319) <= b;
    layer5_outputs(5320) <= not a;
    layer5_outputs(5321) <= a xor b;
    layer5_outputs(5322) <= not b;
    layer5_outputs(5323) <= not (a or b);
    layer5_outputs(5324) <= not (a or b);
    layer5_outputs(5325) <= a or b;
    layer5_outputs(5326) <= a and b;
    layer5_outputs(5327) <= a and b;
    layer5_outputs(5328) <= b;
    layer5_outputs(5329) <= a or b;
    layer5_outputs(5330) <= not b or a;
    layer5_outputs(5331) <= b;
    layer5_outputs(5332) <= not a;
    layer5_outputs(5333) <= b and not a;
    layer5_outputs(5334) <= a and b;
    layer5_outputs(5335) <= not a or b;
    layer5_outputs(5336) <= a or b;
    layer5_outputs(5337) <= not a or b;
    layer5_outputs(5338) <= b;
    layer5_outputs(5339) <= a xor b;
    layer5_outputs(5340) <= b and not a;
    layer5_outputs(5341) <= a or b;
    layer5_outputs(5342) <= '0';
    layer5_outputs(5343) <= a xor b;
    layer5_outputs(5344) <= b and not a;
    layer5_outputs(5345) <= a and not b;
    layer5_outputs(5346) <= b;
    layer5_outputs(5347) <= a;
    layer5_outputs(5348) <= not (a and b);
    layer5_outputs(5349) <= b;
    layer5_outputs(5350) <= '1';
    layer5_outputs(5351) <= a and not b;
    layer5_outputs(5352) <= a and not b;
    layer5_outputs(5353) <= b and not a;
    layer5_outputs(5354) <= '1';
    layer5_outputs(5355) <= a;
    layer5_outputs(5356) <= not (a or b);
    layer5_outputs(5357) <= a or b;
    layer5_outputs(5358) <= a and b;
    layer5_outputs(5359) <= a and not b;
    layer5_outputs(5360) <= b;
    layer5_outputs(5361) <= b;
    layer5_outputs(5362) <= a and not b;
    layer5_outputs(5363) <= a and b;
    layer5_outputs(5364) <= not (a or b);
    layer5_outputs(5365) <= a;
    layer5_outputs(5366) <= not a;
    layer5_outputs(5367) <= b;
    layer5_outputs(5368) <= b;
    layer5_outputs(5369) <= a and b;
    layer5_outputs(5370) <= not a;
    layer5_outputs(5371) <= not b;
    layer5_outputs(5372) <= not a;
    layer5_outputs(5373) <= a or b;
    layer5_outputs(5374) <= not b or a;
    layer5_outputs(5375) <= not b or a;
    layer5_outputs(5376) <= not b;
    layer5_outputs(5377) <= a and not b;
    layer5_outputs(5378) <= b;
    layer5_outputs(5379) <= not a;
    layer5_outputs(5380) <= not a or b;
    layer5_outputs(5381) <= not (a and b);
    layer5_outputs(5382) <= not a;
    layer5_outputs(5383) <= not b or a;
    layer5_outputs(5384) <= not b or a;
    layer5_outputs(5385) <= not b or a;
    layer5_outputs(5386) <= not (a or b);
    layer5_outputs(5387) <= b and not a;
    layer5_outputs(5388) <= a xor b;
    layer5_outputs(5389) <= a xor b;
    layer5_outputs(5390) <= a and not b;
    layer5_outputs(5391) <= not (a or b);
    layer5_outputs(5392) <= a and not b;
    layer5_outputs(5393) <= a and b;
    layer5_outputs(5394) <= '1';
    layer5_outputs(5395) <= not (a or b);
    layer5_outputs(5396) <= not a;
    layer5_outputs(5397) <= not b;
    layer5_outputs(5398) <= a and b;
    layer5_outputs(5399) <= not (a and b);
    layer5_outputs(5400) <= b and not a;
    layer5_outputs(5401) <= not (a and b);
    layer5_outputs(5402) <= not a;
    layer5_outputs(5403) <= not b;
    layer5_outputs(5404) <= not b or a;
    layer5_outputs(5405) <= a;
    layer5_outputs(5406) <= not (a or b);
    layer5_outputs(5407) <= a and not b;
    layer5_outputs(5408) <= a xor b;
    layer5_outputs(5409) <= not b;
    layer5_outputs(5410) <= not (a xor b);
    layer5_outputs(5411) <= not a;
    layer5_outputs(5412) <= a;
    layer5_outputs(5413) <= not b;
    layer5_outputs(5414) <= b;
    layer5_outputs(5415) <= not b;
    layer5_outputs(5416) <= not b;
    layer5_outputs(5417) <= not (a and b);
    layer5_outputs(5418) <= not a;
    layer5_outputs(5419) <= b;
    layer5_outputs(5420) <= a;
    layer5_outputs(5421) <= '0';
    layer5_outputs(5422) <= '1';
    layer5_outputs(5423) <= not b or a;
    layer5_outputs(5424) <= not (a xor b);
    layer5_outputs(5425) <= a and b;
    layer5_outputs(5426) <= '1';
    layer5_outputs(5427) <= not b or a;
    layer5_outputs(5428) <= b;
    layer5_outputs(5429) <= not a;
    layer5_outputs(5430) <= not (a xor b);
    layer5_outputs(5431) <= b;
    layer5_outputs(5432) <= not a;
    layer5_outputs(5433) <= b;
    layer5_outputs(5434) <= not (a or b);
    layer5_outputs(5435) <= not b;
    layer5_outputs(5436) <= a and b;
    layer5_outputs(5437) <= '0';
    layer5_outputs(5438) <= not a or b;
    layer5_outputs(5439) <= a and b;
    layer5_outputs(5440) <= a xor b;
    layer5_outputs(5441) <= not b or a;
    layer5_outputs(5442) <= not a or b;
    layer5_outputs(5443) <= a;
    layer5_outputs(5444) <= a xor b;
    layer5_outputs(5445) <= b and not a;
    layer5_outputs(5446) <= b and not a;
    layer5_outputs(5447) <= a and b;
    layer5_outputs(5448) <= b;
    layer5_outputs(5449) <= not (a or b);
    layer5_outputs(5450) <= a;
    layer5_outputs(5451) <= not b or a;
    layer5_outputs(5452) <= not b or a;
    layer5_outputs(5453) <= b and not a;
    layer5_outputs(5454) <= a and b;
    layer5_outputs(5455) <= not b;
    layer5_outputs(5456) <= not (a and b);
    layer5_outputs(5457) <= '1';
    layer5_outputs(5458) <= a and not b;
    layer5_outputs(5459) <= a or b;
    layer5_outputs(5460) <= a and not b;
    layer5_outputs(5461) <= a xor b;
    layer5_outputs(5462) <= b;
    layer5_outputs(5463) <= '1';
    layer5_outputs(5464) <= not (a and b);
    layer5_outputs(5465) <= '1';
    layer5_outputs(5466) <= '0';
    layer5_outputs(5467) <= a xor b;
    layer5_outputs(5468) <= not (a or b);
    layer5_outputs(5469) <= not b or a;
    layer5_outputs(5470) <= a;
    layer5_outputs(5471) <= not a;
    layer5_outputs(5472) <= a and b;
    layer5_outputs(5473) <= a;
    layer5_outputs(5474) <= a;
    layer5_outputs(5475) <= not (a or b);
    layer5_outputs(5476) <= b;
    layer5_outputs(5477) <= a;
    layer5_outputs(5478) <= not b;
    layer5_outputs(5479) <= a and not b;
    layer5_outputs(5480) <= not (a xor b);
    layer5_outputs(5481) <= not (a and b);
    layer5_outputs(5482) <= not b or a;
    layer5_outputs(5483) <= b and not a;
    layer5_outputs(5484) <= not (a or b);
    layer5_outputs(5485) <= not b or a;
    layer5_outputs(5486) <= not b;
    layer5_outputs(5487) <= b;
    layer5_outputs(5488) <= a;
    layer5_outputs(5489) <= a;
    layer5_outputs(5490) <= a and b;
    layer5_outputs(5491) <= not a or b;
    layer5_outputs(5492) <= a;
    layer5_outputs(5493) <= not (a and b);
    layer5_outputs(5494) <= not (a xor b);
    layer5_outputs(5495) <= a and b;
    layer5_outputs(5496) <= not a;
    layer5_outputs(5497) <= a or b;
    layer5_outputs(5498) <= not (a and b);
    layer5_outputs(5499) <= not a;
    layer5_outputs(5500) <= not b or a;
    layer5_outputs(5501) <= not (a or b);
    layer5_outputs(5502) <= a;
    layer5_outputs(5503) <= '1';
    layer5_outputs(5504) <= b;
    layer5_outputs(5505) <= a or b;
    layer5_outputs(5506) <= not a or b;
    layer5_outputs(5507) <= '0';
    layer5_outputs(5508) <= not (a or b);
    layer5_outputs(5509) <= b and not a;
    layer5_outputs(5510) <= a;
    layer5_outputs(5511) <= not (a and b);
    layer5_outputs(5512) <= a or b;
    layer5_outputs(5513) <= not b;
    layer5_outputs(5514) <= not a or b;
    layer5_outputs(5515) <= not a or b;
    layer5_outputs(5516) <= b;
    layer5_outputs(5517) <= a;
    layer5_outputs(5518) <= not a;
    layer5_outputs(5519) <= not b or a;
    layer5_outputs(5520) <= not a;
    layer5_outputs(5521) <= a;
    layer5_outputs(5522) <= not a or b;
    layer5_outputs(5523) <= a;
    layer5_outputs(5524) <= a;
    layer5_outputs(5525) <= not b or a;
    layer5_outputs(5526) <= a or b;
    layer5_outputs(5527) <= not (a and b);
    layer5_outputs(5528) <= not b or a;
    layer5_outputs(5529) <= a;
    layer5_outputs(5530) <= not (a or b);
    layer5_outputs(5531) <= not a;
    layer5_outputs(5532) <= b;
    layer5_outputs(5533) <= a and not b;
    layer5_outputs(5534) <= a xor b;
    layer5_outputs(5535) <= not (a and b);
    layer5_outputs(5536) <= '1';
    layer5_outputs(5537) <= not (a and b);
    layer5_outputs(5538) <= b;
    layer5_outputs(5539) <= not b;
    layer5_outputs(5540) <= not a or b;
    layer5_outputs(5541) <= b and not a;
    layer5_outputs(5542) <= not b;
    layer5_outputs(5543) <= not a or b;
    layer5_outputs(5544) <= '0';
    layer5_outputs(5545) <= a xor b;
    layer5_outputs(5546) <= not b;
    layer5_outputs(5547) <= b;
    layer5_outputs(5548) <= not b;
    layer5_outputs(5549) <= not b or a;
    layer5_outputs(5550) <= not b or a;
    layer5_outputs(5551) <= b;
    layer5_outputs(5552) <= a xor b;
    layer5_outputs(5553) <= a;
    layer5_outputs(5554) <= b;
    layer5_outputs(5555) <= b and not a;
    layer5_outputs(5556) <= not (a or b);
    layer5_outputs(5557) <= a;
    layer5_outputs(5558) <= '0';
    layer5_outputs(5559) <= not a or b;
    layer5_outputs(5560) <= a xor b;
    layer5_outputs(5561) <= b;
    layer5_outputs(5562) <= not a or b;
    layer5_outputs(5563) <= a;
    layer5_outputs(5564) <= not b;
    layer5_outputs(5565) <= not (a or b);
    layer5_outputs(5566) <= not (a or b);
    layer5_outputs(5567) <= b and not a;
    layer5_outputs(5568) <= not (a xor b);
    layer5_outputs(5569) <= not (a and b);
    layer5_outputs(5570) <= a;
    layer5_outputs(5571) <= not b;
    layer5_outputs(5572) <= a;
    layer5_outputs(5573) <= not a or b;
    layer5_outputs(5574) <= b and not a;
    layer5_outputs(5575) <= a or b;
    layer5_outputs(5576) <= not a;
    layer5_outputs(5577) <= not b or a;
    layer5_outputs(5578) <= '0';
    layer5_outputs(5579) <= a and b;
    layer5_outputs(5580) <= a;
    layer5_outputs(5581) <= a or b;
    layer5_outputs(5582) <= '1';
    layer5_outputs(5583) <= a;
    layer5_outputs(5584) <= a or b;
    layer5_outputs(5585) <= a and not b;
    layer5_outputs(5586) <= not b;
    layer5_outputs(5587) <= b;
    layer5_outputs(5588) <= '1';
    layer5_outputs(5589) <= not b or a;
    layer5_outputs(5590) <= b;
    layer5_outputs(5591) <= not (a and b);
    layer5_outputs(5592) <= b;
    layer5_outputs(5593) <= a or b;
    layer5_outputs(5594) <= a and not b;
    layer5_outputs(5595) <= a and b;
    layer5_outputs(5596) <= not (a xor b);
    layer5_outputs(5597) <= not b;
    layer5_outputs(5598) <= a;
    layer5_outputs(5599) <= not (a or b);
    layer5_outputs(5600) <= a xor b;
    layer5_outputs(5601) <= b;
    layer5_outputs(5602) <= not a or b;
    layer5_outputs(5603) <= a and not b;
    layer5_outputs(5604) <= b and not a;
    layer5_outputs(5605) <= a;
    layer5_outputs(5606) <= '1';
    layer5_outputs(5607) <= not a or b;
    layer5_outputs(5608) <= a and not b;
    layer5_outputs(5609) <= not (a or b);
    layer5_outputs(5610) <= a and b;
    layer5_outputs(5611) <= not a or b;
    layer5_outputs(5612) <= a xor b;
    layer5_outputs(5613) <= not b;
    layer5_outputs(5614) <= a or b;
    layer5_outputs(5615) <= '0';
    layer5_outputs(5616) <= not a;
    layer5_outputs(5617) <= a;
    layer5_outputs(5618) <= not (a and b);
    layer5_outputs(5619) <= not a;
    layer5_outputs(5620) <= not (a and b);
    layer5_outputs(5621) <= a and not b;
    layer5_outputs(5622) <= '1';
    layer5_outputs(5623) <= not (a xor b);
    layer5_outputs(5624) <= b and not a;
    layer5_outputs(5625) <= not b;
    layer5_outputs(5626) <= not b or a;
    layer5_outputs(5627) <= '1';
    layer5_outputs(5628) <= not a or b;
    layer5_outputs(5629) <= not (a or b);
    layer5_outputs(5630) <= a and not b;
    layer5_outputs(5631) <= not a or b;
    layer5_outputs(5632) <= b;
    layer5_outputs(5633) <= not (a and b);
    layer5_outputs(5634) <= not a;
    layer5_outputs(5635) <= not a or b;
    layer5_outputs(5636) <= not b;
    layer5_outputs(5637) <= not b or a;
    layer5_outputs(5638) <= not (a and b);
    layer5_outputs(5639) <= not (a or b);
    layer5_outputs(5640) <= '0';
    layer5_outputs(5641) <= not (a or b);
    layer5_outputs(5642) <= '1';
    layer5_outputs(5643) <= not a;
    layer5_outputs(5644) <= a xor b;
    layer5_outputs(5645) <= not a;
    layer5_outputs(5646) <= not a;
    layer5_outputs(5647) <= b and not a;
    layer5_outputs(5648) <= not (a xor b);
    layer5_outputs(5649) <= a;
    layer5_outputs(5650) <= a or b;
    layer5_outputs(5651) <= a and b;
    layer5_outputs(5652) <= a;
    layer5_outputs(5653) <= not a or b;
    layer5_outputs(5654) <= not (a and b);
    layer5_outputs(5655) <= not a;
    layer5_outputs(5656) <= a and b;
    layer5_outputs(5657) <= b and not a;
    layer5_outputs(5658) <= '0';
    layer5_outputs(5659) <= a or b;
    layer5_outputs(5660) <= a and b;
    layer5_outputs(5661) <= b;
    layer5_outputs(5662) <= not (a and b);
    layer5_outputs(5663) <= not b;
    layer5_outputs(5664) <= not b or a;
    layer5_outputs(5665) <= a;
    layer5_outputs(5666) <= a and not b;
    layer5_outputs(5667) <= a;
    layer5_outputs(5668) <= not b or a;
    layer5_outputs(5669) <= not a;
    layer5_outputs(5670) <= a and b;
    layer5_outputs(5671) <= not b;
    layer5_outputs(5672) <= a xor b;
    layer5_outputs(5673) <= not a;
    layer5_outputs(5674) <= a or b;
    layer5_outputs(5675) <= not b or a;
    layer5_outputs(5676) <= a or b;
    layer5_outputs(5677) <= '1';
    layer5_outputs(5678) <= not a;
    layer5_outputs(5679) <= not b;
    layer5_outputs(5680) <= a;
    layer5_outputs(5681) <= a and b;
    layer5_outputs(5682) <= '1';
    layer5_outputs(5683) <= '1';
    layer5_outputs(5684) <= a and b;
    layer5_outputs(5685) <= a and b;
    layer5_outputs(5686) <= not b;
    layer5_outputs(5687) <= a or b;
    layer5_outputs(5688) <= a and not b;
    layer5_outputs(5689) <= a and b;
    layer5_outputs(5690) <= a;
    layer5_outputs(5691) <= not b or a;
    layer5_outputs(5692) <= a;
    layer5_outputs(5693) <= not b or a;
    layer5_outputs(5694) <= a and b;
    layer5_outputs(5695) <= not (a and b);
    layer5_outputs(5696) <= b;
    layer5_outputs(5697) <= not (a xor b);
    layer5_outputs(5698) <= a or b;
    layer5_outputs(5699) <= b and not a;
    layer5_outputs(5700) <= not (a or b);
    layer5_outputs(5701) <= '0';
    layer5_outputs(5702) <= a;
    layer5_outputs(5703) <= not a;
    layer5_outputs(5704) <= not (a and b);
    layer5_outputs(5705) <= not b or a;
    layer5_outputs(5706) <= not a;
    layer5_outputs(5707) <= '0';
    layer5_outputs(5708) <= a and b;
    layer5_outputs(5709) <= not (a xor b);
    layer5_outputs(5710) <= a;
    layer5_outputs(5711) <= a or b;
    layer5_outputs(5712) <= not b;
    layer5_outputs(5713) <= not b;
    layer5_outputs(5714) <= b and not a;
    layer5_outputs(5715) <= not b;
    layer5_outputs(5716) <= a xor b;
    layer5_outputs(5717) <= not b or a;
    layer5_outputs(5718) <= a and b;
    layer5_outputs(5719) <= not (a xor b);
    layer5_outputs(5720) <= a xor b;
    layer5_outputs(5721) <= a xor b;
    layer5_outputs(5722) <= not (a or b);
    layer5_outputs(5723) <= not a;
    layer5_outputs(5724) <= a;
    layer5_outputs(5725) <= b;
    layer5_outputs(5726) <= not (a xor b);
    layer5_outputs(5727) <= a and not b;
    layer5_outputs(5728) <= a and not b;
    layer5_outputs(5729) <= a xor b;
    layer5_outputs(5730) <= not b or a;
    layer5_outputs(5731) <= not b or a;
    layer5_outputs(5732) <= a;
    layer5_outputs(5733) <= '0';
    layer5_outputs(5734) <= not b or a;
    layer5_outputs(5735) <= a and not b;
    layer5_outputs(5736) <= b;
    layer5_outputs(5737) <= not a;
    layer5_outputs(5738) <= a and not b;
    layer5_outputs(5739) <= not b;
    layer5_outputs(5740) <= b;
    layer5_outputs(5741) <= b;
    layer5_outputs(5742) <= '0';
    layer5_outputs(5743) <= a and b;
    layer5_outputs(5744) <= not a;
    layer5_outputs(5745) <= not a or b;
    layer5_outputs(5746) <= b;
    layer5_outputs(5747) <= not (a or b);
    layer5_outputs(5748) <= '0';
    layer5_outputs(5749) <= not b;
    layer5_outputs(5750) <= not (a xor b);
    layer5_outputs(5751) <= '0';
    layer5_outputs(5752) <= b and not a;
    layer5_outputs(5753) <= a and not b;
    layer5_outputs(5754) <= b;
    layer5_outputs(5755) <= '0';
    layer5_outputs(5756) <= '0';
    layer5_outputs(5757) <= a and b;
    layer5_outputs(5758) <= not (a xor b);
    layer5_outputs(5759) <= a and not b;
    layer5_outputs(5760) <= a and b;
    layer5_outputs(5761) <= not (a or b);
    layer5_outputs(5762) <= a and b;
    layer5_outputs(5763) <= not b or a;
    layer5_outputs(5764) <= not a;
    layer5_outputs(5765) <= a;
    layer5_outputs(5766) <= not a;
    layer5_outputs(5767) <= a and b;
    layer5_outputs(5768) <= not (a xor b);
    layer5_outputs(5769) <= not (a and b);
    layer5_outputs(5770) <= b;
    layer5_outputs(5771) <= b;
    layer5_outputs(5772) <= a and not b;
    layer5_outputs(5773) <= not b;
    layer5_outputs(5774) <= a or b;
    layer5_outputs(5775) <= a and b;
    layer5_outputs(5776) <= not (a or b);
    layer5_outputs(5777) <= a or b;
    layer5_outputs(5778) <= not (a and b);
    layer5_outputs(5779) <= a or b;
    layer5_outputs(5780) <= not b or a;
    layer5_outputs(5781) <= a;
    layer5_outputs(5782) <= not b or a;
    layer5_outputs(5783) <= not (a and b);
    layer5_outputs(5784) <= a;
    layer5_outputs(5785) <= '1';
    layer5_outputs(5786) <= not b;
    layer5_outputs(5787) <= a and b;
    layer5_outputs(5788) <= not (a xor b);
    layer5_outputs(5789) <= b;
    layer5_outputs(5790) <= not a or b;
    layer5_outputs(5791) <= b;
    layer5_outputs(5792) <= '0';
    layer5_outputs(5793) <= not b;
    layer5_outputs(5794) <= not b;
    layer5_outputs(5795) <= a and b;
    layer5_outputs(5796) <= a and not b;
    layer5_outputs(5797) <= a and not b;
    layer5_outputs(5798) <= not (a and b);
    layer5_outputs(5799) <= a or b;
    layer5_outputs(5800) <= not a;
    layer5_outputs(5801) <= a and not b;
    layer5_outputs(5802) <= a xor b;
    layer5_outputs(5803) <= not a or b;
    layer5_outputs(5804) <= not (a or b);
    layer5_outputs(5805) <= b;
    layer5_outputs(5806) <= not (a xor b);
    layer5_outputs(5807) <= not (a and b);
    layer5_outputs(5808) <= b and not a;
    layer5_outputs(5809) <= a and b;
    layer5_outputs(5810) <= not (a xor b);
    layer5_outputs(5811) <= not b or a;
    layer5_outputs(5812) <= not b;
    layer5_outputs(5813) <= not b;
    layer5_outputs(5814) <= a;
    layer5_outputs(5815) <= not b or a;
    layer5_outputs(5816) <= '0';
    layer5_outputs(5817) <= not a or b;
    layer5_outputs(5818) <= not b;
    layer5_outputs(5819) <= a and not b;
    layer5_outputs(5820) <= a and not b;
    layer5_outputs(5821) <= b;
    layer5_outputs(5822) <= not a;
    layer5_outputs(5823) <= b and not a;
    layer5_outputs(5824) <= b and not a;
    layer5_outputs(5825) <= '0';
    layer5_outputs(5826) <= not (a xor b);
    layer5_outputs(5827) <= a;
    layer5_outputs(5828) <= not b;
    layer5_outputs(5829) <= not a or b;
    layer5_outputs(5830) <= not a;
    layer5_outputs(5831) <= a and b;
    layer5_outputs(5832) <= a;
    layer5_outputs(5833) <= b and not a;
    layer5_outputs(5834) <= b and not a;
    layer5_outputs(5835) <= not a or b;
    layer5_outputs(5836) <= not a;
    layer5_outputs(5837) <= a or b;
    layer5_outputs(5838) <= b;
    layer5_outputs(5839) <= not (a xor b);
    layer5_outputs(5840) <= a;
    layer5_outputs(5841) <= a and not b;
    layer5_outputs(5842) <= not b or a;
    layer5_outputs(5843) <= not a;
    layer5_outputs(5844) <= a and b;
    layer5_outputs(5845) <= not (a or b);
    layer5_outputs(5846) <= not a;
    layer5_outputs(5847) <= a and not b;
    layer5_outputs(5848) <= b and not a;
    layer5_outputs(5849) <= not (a and b);
    layer5_outputs(5850) <= not (a or b);
    layer5_outputs(5851) <= a and b;
    layer5_outputs(5852) <= a and not b;
    layer5_outputs(5853) <= not (a xor b);
    layer5_outputs(5854) <= a and not b;
    layer5_outputs(5855) <= not (a or b);
    layer5_outputs(5856) <= not (a and b);
    layer5_outputs(5857) <= a or b;
    layer5_outputs(5858) <= a and not b;
    layer5_outputs(5859) <= a or b;
    layer5_outputs(5860) <= a and not b;
    layer5_outputs(5861) <= a or b;
    layer5_outputs(5862) <= not a;
    layer5_outputs(5863) <= '0';
    layer5_outputs(5864) <= a;
    layer5_outputs(5865) <= '0';
    layer5_outputs(5866) <= not a;
    layer5_outputs(5867) <= a;
    layer5_outputs(5868) <= a or b;
    layer5_outputs(5869) <= a;
    layer5_outputs(5870) <= not a;
    layer5_outputs(5871) <= a and b;
    layer5_outputs(5872) <= b and not a;
    layer5_outputs(5873) <= a;
    layer5_outputs(5874) <= a;
    layer5_outputs(5875) <= a or b;
    layer5_outputs(5876) <= not a;
    layer5_outputs(5877) <= not b or a;
    layer5_outputs(5878) <= b and not a;
    layer5_outputs(5879) <= b and not a;
    layer5_outputs(5880) <= a;
    layer5_outputs(5881) <= not b;
    layer5_outputs(5882) <= not a;
    layer5_outputs(5883) <= '0';
    layer5_outputs(5884) <= b and not a;
    layer5_outputs(5885) <= a xor b;
    layer5_outputs(5886) <= not a or b;
    layer5_outputs(5887) <= '0';
    layer5_outputs(5888) <= '1';
    layer5_outputs(5889) <= a xor b;
    layer5_outputs(5890) <= not b;
    layer5_outputs(5891) <= a and b;
    layer5_outputs(5892) <= not b;
    layer5_outputs(5893) <= a or b;
    layer5_outputs(5894) <= '0';
    layer5_outputs(5895) <= a or b;
    layer5_outputs(5896) <= a xor b;
    layer5_outputs(5897) <= b;
    layer5_outputs(5898) <= b and not a;
    layer5_outputs(5899) <= b and not a;
    layer5_outputs(5900) <= not a;
    layer5_outputs(5901) <= not (a and b);
    layer5_outputs(5902) <= a or b;
    layer5_outputs(5903) <= b;
    layer5_outputs(5904) <= b and not a;
    layer5_outputs(5905) <= a and b;
    layer5_outputs(5906) <= not b or a;
    layer5_outputs(5907) <= b;
    layer5_outputs(5908) <= not a;
    layer5_outputs(5909) <= not (a xor b);
    layer5_outputs(5910) <= '1';
    layer5_outputs(5911) <= not b;
    layer5_outputs(5912) <= '0';
    layer5_outputs(5913) <= b and not a;
    layer5_outputs(5914) <= not b or a;
    layer5_outputs(5915) <= b and not a;
    layer5_outputs(5916) <= a or b;
    layer5_outputs(5917) <= not (a and b);
    layer5_outputs(5918) <= not (a and b);
    layer5_outputs(5919) <= not (a or b);
    layer5_outputs(5920) <= not b;
    layer5_outputs(5921) <= a xor b;
    layer5_outputs(5922) <= b and not a;
    layer5_outputs(5923) <= a and not b;
    layer5_outputs(5924) <= b;
    layer5_outputs(5925) <= not a or b;
    layer5_outputs(5926) <= '1';
    layer5_outputs(5927) <= not (a and b);
    layer5_outputs(5928) <= b;
    layer5_outputs(5929) <= not a;
    layer5_outputs(5930) <= a or b;
    layer5_outputs(5931) <= not a;
    layer5_outputs(5932) <= b and not a;
    layer5_outputs(5933) <= not b;
    layer5_outputs(5934) <= not b or a;
    layer5_outputs(5935) <= '0';
    layer5_outputs(5936) <= not (a or b);
    layer5_outputs(5937) <= a and b;
    layer5_outputs(5938) <= a or b;
    layer5_outputs(5939) <= a and b;
    layer5_outputs(5940) <= a;
    layer5_outputs(5941) <= a and b;
    layer5_outputs(5942) <= b;
    layer5_outputs(5943) <= not a or b;
    layer5_outputs(5944) <= not b or a;
    layer5_outputs(5945) <= not a;
    layer5_outputs(5946) <= b and not a;
    layer5_outputs(5947) <= not b or a;
    layer5_outputs(5948) <= not a;
    layer5_outputs(5949) <= not b;
    layer5_outputs(5950) <= not a or b;
    layer5_outputs(5951) <= b;
    layer5_outputs(5952) <= a;
    layer5_outputs(5953) <= a and b;
    layer5_outputs(5954) <= not a or b;
    layer5_outputs(5955) <= a and b;
    layer5_outputs(5956) <= not a;
    layer5_outputs(5957) <= not a or b;
    layer5_outputs(5958) <= b;
    layer5_outputs(5959) <= '0';
    layer5_outputs(5960) <= not a;
    layer5_outputs(5961) <= not a or b;
    layer5_outputs(5962) <= a;
    layer5_outputs(5963) <= a;
    layer5_outputs(5964) <= not a;
    layer5_outputs(5965) <= a and b;
    layer5_outputs(5966) <= a;
    layer5_outputs(5967) <= b;
    layer5_outputs(5968) <= a or b;
    layer5_outputs(5969) <= a;
    layer5_outputs(5970) <= not b;
    layer5_outputs(5971) <= b and not a;
    layer5_outputs(5972) <= a or b;
    layer5_outputs(5973) <= not b;
    layer5_outputs(5974) <= b;
    layer5_outputs(5975) <= b;
    layer5_outputs(5976) <= a or b;
    layer5_outputs(5977) <= b;
    layer5_outputs(5978) <= not b;
    layer5_outputs(5979) <= a and b;
    layer5_outputs(5980) <= not (a and b);
    layer5_outputs(5981) <= b;
    layer5_outputs(5982) <= not (a xor b);
    layer5_outputs(5983) <= a and not b;
    layer5_outputs(5984) <= not b;
    layer5_outputs(5985) <= not (a and b);
    layer5_outputs(5986) <= not a;
    layer5_outputs(5987) <= not (a or b);
    layer5_outputs(5988) <= not (a or b);
    layer5_outputs(5989) <= b and not a;
    layer5_outputs(5990) <= not a or b;
    layer5_outputs(5991) <= not (a and b);
    layer5_outputs(5992) <= a or b;
    layer5_outputs(5993) <= not a;
    layer5_outputs(5994) <= not a;
    layer5_outputs(5995) <= a and b;
    layer5_outputs(5996) <= a;
    layer5_outputs(5997) <= not a or b;
    layer5_outputs(5998) <= a and b;
    layer5_outputs(5999) <= a and not b;
    layer5_outputs(6000) <= a and not b;
    layer5_outputs(6001) <= not (a and b);
    layer5_outputs(6002) <= not a or b;
    layer5_outputs(6003) <= a and not b;
    layer5_outputs(6004) <= not a or b;
    layer5_outputs(6005) <= not b;
    layer5_outputs(6006) <= not b or a;
    layer5_outputs(6007) <= not (a or b);
    layer5_outputs(6008) <= b;
    layer5_outputs(6009) <= not a or b;
    layer5_outputs(6010) <= not a;
    layer5_outputs(6011) <= not (a and b);
    layer5_outputs(6012) <= not (a or b);
    layer5_outputs(6013) <= not a;
    layer5_outputs(6014) <= a;
    layer5_outputs(6015) <= not (a and b);
    layer5_outputs(6016) <= a;
    layer5_outputs(6017) <= a or b;
    layer5_outputs(6018) <= '0';
    layer5_outputs(6019) <= b;
    layer5_outputs(6020) <= a and not b;
    layer5_outputs(6021) <= not b;
    layer5_outputs(6022) <= a xor b;
    layer5_outputs(6023) <= a xor b;
    layer5_outputs(6024) <= a;
    layer5_outputs(6025) <= b and not a;
    layer5_outputs(6026) <= a xor b;
    layer5_outputs(6027) <= not (a or b);
    layer5_outputs(6028) <= not b;
    layer5_outputs(6029) <= not a;
    layer5_outputs(6030) <= a and not b;
    layer5_outputs(6031) <= a;
    layer5_outputs(6032) <= not b;
    layer5_outputs(6033) <= '1';
    layer5_outputs(6034) <= b and not a;
    layer5_outputs(6035) <= a and not b;
    layer5_outputs(6036) <= not a or b;
    layer5_outputs(6037) <= not a;
    layer5_outputs(6038) <= not b or a;
    layer5_outputs(6039) <= a or b;
    layer5_outputs(6040) <= a or b;
    layer5_outputs(6041) <= a and b;
    layer5_outputs(6042) <= a xor b;
    layer5_outputs(6043) <= a and b;
    layer5_outputs(6044) <= a;
    layer5_outputs(6045) <= a and b;
    layer5_outputs(6046) <= not b or a;
    layer5_outputs(6047) <= not b or a;
    layer5_outputs(6048) <= a and b;
    layer5_outputs(6049) <= not a;
    layer5_outputs(6050) <= not b;
    layer5_outputs(6051) <= '0';
    layer5_outputs(6052) <= not (a or b);
    layer5_outputs(6053) <= not a or b;
    layer5_outputs(6054) <= not a;
    layer5_outputs(6055) <= not (a or b);
    layer5_outputs(6056) <= b;
    layer5_outputs(6057) <= a xor b;
    layer5_outputs(6058) <= a;
    layer5_outputs(6059) <= not a;
    layer5_outputs(6060) <= '1';
    layer5_outputs(6061) <= a;
    layer5_outputs(6062) <= not a or b;
    layer5_outputs(6063) <= not b;
    layer5_outputs(6064) <= a and b;
    layer5_outputs(6065) <= not (a and b);
    layer5_outputs(6066) <= not a;
    layer5_outputs(6067) <= not a;
    layer5_outputs(6068) <= not b;
    layer5_outputs(6069) <= not a;
    layer5_outputs(6070) <= not b or a;
    layer5_outputs(6071) <= not a;
    layer5_outputs(6072) <= not b or a;
    layer5_outputs(6073) <= not (a and b);
    layer5_outputs(6074) <= not (a and b);
    layer5_outputs(6075) <= a xor b;
    layer5_outputs(6076) <= a xor b;
    layer5_outputs(6077) <= '1';
    layer5_outputs(6078) <= not b;
    layer5_outputs(6079) <= not a;
    layer5_outputs(6080) <= a;
    layer5_outputs(6081) <= not b;
    layer5_outputs(6082) <= not b or a;
    layer5_outputs(6083) <= not b;
    layer5_outputs(6084) <= a;
    layer5_outputs(6085) <= not a;
    layer5_outputs(6086) <= not b;
    layer5_outputs(6087) <= '0';
    layer5_outputs(6088) <= not b or a;
    layer5_outputs(6089) <= a or b;
    layer5_outputs(6090) <= not a or b;
    layer5_outputs(6091) <= not b;
    layer5_outputs(6092) <= not a or b;
    layer5_outputs(6093) <= a and not b;
    layer5_outputs(6094) <= a;
    layer5_outputs(6095) <= not b;
    layer5_outputs(6096) <= not b;
    layer5_outputs(6097) <= b and not a;
    layer5_outputs(6098) <= not (a and b);
    layer5_outputs(6099) <= a and not b;
    layer5_outputs(6100) <= not (a or b);
    layer5_outputs(6101) <= a and b;
    layer5_outputs(6102) <= b;
    layer5_outputs(6103) <= not a;
    layer5_outputs(6104) <= not b or a;
    layer5_outputs(6105) <= not (a and b);
    layer5_outputs(6106) <= not b;
    layer5_outputs(6107) <= not a;
    layer5_outputs(6108) <= not b or a;
    layer5_outputs(6109) <= not a;
    layer5_outputs(6110) <= '1';
    layer5_outputs(6111) <= a;
    layer5_outputs(6112) <= '1';
    layer5_outputs(6113) <= not b or a;
    layer5_outputs(6114) <= not b;
    layer5_outputs(6115) <= b;
    layer5_outputs(6116) <= a and b;
    layer5_outputs(6117) <= a xor b;
    layer5_outputs(6118) <= a and not b;
    layer5_outputs(6119) <= not b or a;
    layer5_outputs(6120) <= a or b;
    layer5_outputs(6121) <= not (a and b);
    layer5_outputs(6122) <= not b or a;
    layer5_outputs(6123) <= not (a and b);
    layer5_outputs(6124) <= b;
    layer5_outputs(6125) <= not a;
    layer5_outputs(6126) <= a and b;
    layer5_outputs(6127) <= not a or b;
    layer5_outputs(6128) <= not b;
    layer5_outputs(6129) <= not a;
    layer5_outputs(6130) <= not a or b;
    layer5_outputs(6131) <= b and not a;
    layer5_outputs(6132) <= a;
    layer5_outputs(6133) <= not b or a;
    layer5_outputs(6134) <= a;
    layer5_outputs(6135) <= a and not b;
    layer5_outputs(6136) <= '1';
    layer5_outputs(6137) <= b and not a;
    layer5_outputs(6138) <= not b or a;
    layer5_outputs(6139) <= '0';
    layer5_outputs(6140) <= a and b;
    layer5_outputs(6141) <= a and b;
    layer5_outputs(6142) <= not a or b;
    layer5_outputs(6143) <= not (a and b);
    layer5_outputs(6144) <= b;
    layer5_outputs(6145) <= b;
    layer5_outputs(6146) <= not (a and b);
    layer5_outputs(6147) <= a and b;
    layer5_outputs(6148) <= not a;
    layer5_outputs(6149) <= b and not a;
    layer5_outputs(6150) <= a and not b;
    layer5_outputs(6151) <= not (a or b);
    layer5_outputs(6152) <= not (a or b);
    layer5_outputs(6153) <= b;
    layer5_outputs(6154) <= not a or b;
    layer5_outputs(6155) <= b;
    layer5_outputs(6156) <= b;
    layer5_outputs(6157) <= not (a or b);
    layer5_outputs(6158) <= b and not a;
    layer5_outputs(6159) <= not b;
    layer5_outputs(6160) <= not b;
    layer5_outputs(6161) <= not a;
    layer5_outputs(6162) <= not a;
    layer5_outputs(6163) <= a and not b;
    layer5_outputs(6164) <= not b;
    layer5_outputs(6165) <= b and not a;
    layer5_outputs(6166) <= b;
    layer5_outputs(6167) <= a xor b;
    layer5_outputs(6168) <= a and b;
    layer5_outputs(6169) <= not a;
    layer5_outputs(6170) <= a;
    layer5_outputs(6171) <= not a or b;
    layer5_outputs(6172) <= b and not a;
    layer5_outputs(6173) <= b and not a;
    layer5_outputs(6174) <= a or b;
    layer5_outputs(6175) <= not b;
    layer5_outputs(6176) <= not (a and b);
    layer5_outputs(6177) <= a xor b;
    layer5_outputs(6178) <= '1';
    layer5_outputs(6179) <= a;
    layer5_outputs(6180) <= not (a and b);
    layer5_outputs(6181) <= '1';
    layer5_outputs(6182) <= b;
    layer5_outputs(6183) <= not b;
    layer5_outputs(6184) <= not b;
    layer5_outputs(6185) <= '0';
    layer5_outputs(6186) <= not a;
    layer5_outputs(6187) <= b and not a;
    layer5_outputs(6188) <= not a;
    layer5_outputs(6189) <= b;
    layer5_outputs(6190) <= not b or a;
    layer5_outputs(6191) <= not (a and b);
    layer5_outputs(6192) <= a and b;
    layer5_outputs(6193) <= b and not a;
    layer5_outputs(6194) <= not b;
    layer5_outputs(6195) <= not b;
    layer5_outputs(6196) <= a;
    layer5_outputs(6197) <= not b or a;
    layer5_outputs(6198) <= '0';
    layer5_outputs(6199) <= a;
    layer5_outputs(6200) <= not (a or b);
    layer5_outputs(6201) <= b and not a;
    layer5_outputs(6202) <= a and not b;
    layer5_outputs(6203) <= a xor b;
    layer5_outputs(6204) <= a and not b;
    layer5_outputs(6205) <= a or b;
    layer5_outputs(6206) <= '0';
    layer5_outputs(6207) <= b;
    layer5_outputs(6208) <= not a;
    layer5_outputs(6209) <= not a;
    layer5_outputs(6210) <= not a or b;
    layer5_outputs(6211) <= a and b;
    layer5_outputs(6212) <= a and not b;
    layer5_outputs(6213) <= b and not a;
    layer5_outputs(6214) <= a and not b;
    layer5_outputs(6215) <= '1';
    layer5_outputs(6216) <= a and b;
    layer5_outputs(6217) <= not a;
    layer5_outputs(6218) <= not b;
    layer5_outputs(6219) <= '0';
    layer5_outputs(6220) <= not a;
    layer5_outputs(6221) <= not (a and b);
    layer5_outputs(6222) <= not (a and b);
    layer5_outputs(6223) <= not (a xor b);
    layer5_outputs(6224) <= b and not a;
    layer5_outputs(6225) <= a or b;
    layer5_outputs(6226) <= a and not b;
    layer5_outputs(6227) <= a;
    layer5_outputs(6228) <= b;
    layer5_outputs(6229) <= not a or b;
    layer5_outputs(6230) <= not a;
    layer5_outputs(6231) <= not b;
    layer5_outputs(6232) <= not (a xor b);
    layer5_outputs(6233) <= a xor b;
    layer5_outputs(6234) <= b and not a;
    layer5_outputs(6235) <= a;
    layer5_outputs(6236) <= a xor b;
    layer5_outputs(6237) <= a xor b;
    layer5_outputs(6238) <= a or b;
    layer5_outputs(6239) <= not (a xor b);
    layer5_outputs(6240) <= a xor b;
    layer5_outputs(6241) <= not (a and b);
    layer5_outputs(6242) <= b;
    layer5_outputs(6243) <= a and b;
    layer5_outputs(6244) <= b;
    layer5_outputs(6245) <= b;
    layer5_outputs(6246) <= not b;
    layer5_outputs(6247) <= not (a and b);
    layer5_outputs(6248) <= not b;
    layer5_outputs(6249) <= not a;
    layer5_outputs(6250) <= a or b;
    layer5_outputs(6251) <= not a;
    layer5_outputs(6252) <= a or b;
    layer5_outputs(6253) <= '0';
    layer5_outputs(6254) <= a or b;
    layer5_outputs(6255) <= not a;
    layer5_outputs(6256) <= not b or a;
    layer5_outputs(6257) <= not (a or b);
    layer5_outputs(6258) <= a;
    layer5_outputs(6259) <= not b or a;
    layer5_outputs(6260) <= not b or a;
    layer5_outputs(6261) <= a or b;
    layer5_outputs(6262) <= not b or a;
    layer5_outputs(6263) <= a and b;
    layer5_outputs(6264) <= a or b;
    layer5_outputs(6265) <= not (a or b);
    layer5_outputs(6266) <= not a;
    layer5_outputs(6267) <= not (a xor b);
    layer5_outputs(6268) <= a;
    layer5_outputs(6269) <= not (a and b);
    layer5_outputs(6270) <= b and not a;
    layer5_outputs(6271) <= a and not b;
    layer5_outputs(6272) <= not (a or b);
    layer5_outputs(6273) <= b;
    layer5_outputs(6274) <= a and b;
    layer5_outputs(6275) <= '0';
    layer5_outputs(6276) <= b;
    layer5_outputs(6277) <= not a or b;
    layer5_outputs(6278) <= not a;
    layer5_outputs(6279) <= b;
    layer5_outputs(6280) <= b;
    layer5_outputs(6281) <= not a;
    layer5_outputs(6282) <= not b or a;
    layer5_outputs(6283) <= not b;
    layer5_outputs(6284) <= a or b;
    layer5_outputs(6285) <= '0';
    layer5_outputs(6286) <= not (a and b);
    layer5_outputs(6287) <= not a;
    layer5_outputs(6288) <= not (a xor b);
    layer5_outputs(6289) <= not a;
    layer5_outputs(6290) <= not (a xor b);
    layer5_outputs(6291) <= b;
    layer5_outputs(6292) <= not (a xor b);
    layer5_outputs(6293) <= '0';
    layer5_outputs(6294) <= a or b;
    layer5_outputs(6295) <= not b or a;
    layer5_outputs(6296) <= not (a xor b);
    layer5_outputs(6297) <= a and b;
    layer5_outputs(6298) <= b;
    layer5_outputs(6299) <= b;
    layer5_outputs(6300) <= a;
    layer5_outputs(6301) <= not b;
    layer5_outputs(6302) <= b and not a;
    layer5_outputs(6303) <= b and not a;
    layer5_outputs(6304) <= not a;
    layer5_outputs(6305) <= '1';
    layer5_outputs(6306) <= a and b;
    layer5_outputs(6307) <= not b;
    layer5_outputs(6308) <= b;
    layer5_outputs(6309) <= not (a and b);
    layer5_outputs(6310) <= not a;
    layer5_outputs(6311) <= a and b;
    layer5_outputs(6312) <= a and not b;
    layer5_outputs(6313) <= not (a or b);
    layer5_outputs(6314) <= '0';
    layer5_outputs(6315) <= '0';
    layer5_outputs(6316) <= not a;
    layer5_outputs(6317) <= not b;
    layer5_outputs(6318) <= not b;
    layer5_outputs(6319) <= not a;
    layer5_outputs(6320) <= not a or b;
    layer5_outputs(6321) <= b and not a;
    layer5_outputs(6322) <= a;
    layer5_outputs(6323) <= '0';
    layer5_outputs(6324) <= not a or b;
    layer5_outputs(6325) <= b;
    layer5_outputs(6326) <= b;
    layer5_outputs(6327) <= not b or a;
    layer5_outputs(6328) <= not a;
    layer5_outputs(6329) <= b and not a;
    layer5_outputs(6330) <= a or b;
    layer5_outputs(6331) <= '0';
    layer5_outputs(6332) <= b and not a;
    layer5_outputs(6333) <= a;
    layer5_outputs(6334) <= not (a xor b);
    layer5_outputs(6335) <= not b;
    layer5_outputs(6336) <= '0';
    layer5_outputs(6337) <= not a;
    layer5_outputs(6338) <= a and b;
    layer5_outputs(6339) <= not (a or b);
    layer5_outputs(6340) <= not a;
    layer5_outputs(6341) <= b and not a;
    layer5_outputs(6342) <= not b or a;
    layer5_outputs(6343) <= a or b;
    layer5_outputs(6344) <= b and not a;
    layer5_outputs(6345) <= b;
    layer5_outputs(6346) <= not (a and b);
    layer5_outputs(6347) <= b;
    layer5_outputs(6348) <= b and not a;
    layer5_outputs(6349) <= a;
    layer5_outputs(6350) <= a and not b;
    layer5_outputs(6351) <= not b;
    layer5_outputs(6352) <= not b;
    layer5_outputs(6353) <= '1';
    layer5_outputs(6354) <= a and not b;
    layer5_outputs(6355) <= not a or b;
    layer5_outputs(6356) <= not b or a;
    layer5_outputs(6357) <= not b or a;
    layer5_outputs(6358) <= a;
    layer5_outputs(6359) <= a and not b;
    layer5_outputs(6360) <= a xor b;
    layer5_outputs(6361) <= not (a and b);
    layer5_outputs(6362) <= not b;
    layer5_outputs(6363) <= not (a or b);
    layer5_outputs(6364) <= b and not a;
    layer5_outputs(6365) <= '1';
    layer5_outputs(6366) <= not b;
    layer5_outputs(6367) <= not (a or b);
    layer5_outputs(6368) <= a or b;
    layer5_outputs(6369) <= not (a or b);
    layer5_outputs(6370) <= a and not b;
    layer5_outputs(6371) <= not b or a;
    layer5_outputs(6372) <= a and b;
    layer5_outputs(6373) <= b and not a;
    layer5_outputs(6374) <= not (a and b);
    layer5_outputs(6375) <= a and not b;
    layer5_outputs(6376) <= '1';
    layer5_outputs(6377) <= a;
    layer5_outputs(6378) <= not a or b;
    layer5_outputs(6379) <= a;
    layer5_outputs(6380) <= not b;
    layer5_outputs(6381) <= a and b;
    layer5_outputs(6382) <= a or b;
    layer5_outputs(6383) <= b and not a;
    layer5_outputs(6384) <= not a;
    layer5_outputs(6385) <= not (a xor b);
    layer5_outputs(6386) <= not b or a;
    layer5_outputs(6387) <= b and not a;
    layer5_outputs(6388) <= not b;
    layer5_outputs(6389) <= not b;
    layer5_outputs(6390) <= a;
    layer5_outputs(6391) <= b;
    layer5_outputs(6392) <= '1';
    layer5_outputs(6393) <= '0';
    layer5_outputs(6394) <= not a;
    layer5_outputs(6395) <= not (a or b);
    layer5_outputs(6396) <= not a or b;
    layer5_outputs(6397) <= a and not b;
    layer5_outputs(6398) <= '1';
    layer5_outputs(6399) <= a;
    layer5_outputs(6400) <= not b;
    layer5_outputs(6401) <= b;
    layer5_outputs(6402) <= not a;
    layer5_outputs(6403) <= not a or b;
    layer5_outputs(6404) <= a;
    layer5_outputs(6405) <= b;
    layer5_outputs(6406) <= a;
    layer5_outputs(6407) <= a;
    layer5_outputs(6408) <= b;
    layer5_outputs(6409) <= a;
    layer5_outputs(6410) <= not b;
    layer5_outputs(6411) <= '0';
    layer5_outputs(6412) <= not b or a;
    layer5_outputs(6413) <= a or b;
    layer5_outputs(6414) <= '0';
    layer5_outputs(6415) <= b and not a;
    layer5_outputs(6416) <= not (a and b);
    layer5_outputs(6417) <= '1';
    layer5_outputs(6418) <= a and not b;
    layer5_outputs(6419) <= not a or b;
    layer5_outputs(6420) <= a and not b;
    layer5_outputs(6421) <= not a;
    layer5_outputs(6422) <= a xor b;
    layer5_outputs(6423) <= not (a or b);
    layer5_outputs(6424) <= '1';
    layer5_outputs(6425) <= not a or b;
    layer5_outputs(6426) <= not b or a;
    layer5_outputs(6427) <= not b;
    layer5_outputs(6428) <= a and not b;
    layer5_outputs(6429) <= not a or b;
    layer5_outputs(6430) <= b;
    layer5_outputs(6431) <= '0';
    layer5_outputs(6432) <= not b;
    layer5_outputs(6433) <= not b or a;
    layer5_outputs(6434) <= a and b;
    layer5_outputs(6435) <= not a;
    layer5_outputs(6436) <= b;
    layer5_outputs(6437) <= a and not b;
    layer5_outputs(6438) <= b and not a;
    layer5_outputs(6439) <= '0';
    layer5_outputs(6440) <= a and b;
    layer5_outputs(6441) <= '0';
    layer5_outputs(6442) <= not b;
    layer5_outputs(6443) <= a and b;
    layer5_outputs(6444) <= not (a or b);
    layer5_outputs(6445) <= '1';
    layer5_outputs(6446) <= not (a or b);
    layer5_outputs(6447) <= not b or a;
    layer5_outputs(6448) <= b;
    layer5_outputs(6449) <= not b;
    layer5_outputs(6450) <= a or b;
    layer5_outputs(6451) <= not (a and b);
    layer5_outputs(6452) <= not a;
    layer5_outputs(6453) <= a or b;
    layer5_outputs(6454) <= not b or a;
    layer5_outputs(6455) <= not b;
    layer5_outputs(6456) <= b;
    layer5_outputs(6457) <= a or b;
    layer5_outputs(6458) <= a;
    layer5_outputs(6459) <= a or b;
    layer5_outputs(6460) <= b;
    layer5_outputs(6461) <= a xor b;
    layer5_outputs(6462) <= not b;
    layer5_outputs(6463) <= a;
    layer5_outputs(6464) <= not a;
    layer5_outputs(6465) <= not b or a;
    layer5_outputs(6466) <= a;
    layer5_outputs(6467) <= a and not b;
    layer5_outputs(6468) <= a and not b;
    layer5_outputs(6469) <= b;
    layer5_outputs(6470) <= a or b;
    layer5_outputs(6471) <= not (a xor b);
    layer5_outputs(6472) <= not b;
    layer5_outputs(6473) <= b and not a;
    layer5_outputs(6474) <= b and not a;
    layer5_outputs(6475) <= a or b;
    layer5_outputs(6476) <= b and not a;
    layer5_outputs(6477) <= not b;
    layer5_outputs(6478) <= a;
    layer5_outputs(6479) <= b;
    layer5_outputs(6480) <= '1';
    layer5_outputs(6481) <= not (a and b);
    layer5_outputs(6482) <= b;
    layer5_outputs(6483) <= not a;
    layer5_outputs(6484) <= '1';
    layer5_outputs(6485) <= '0';
    layer5_outputs(6486) <= a and b;
    layer5_outputs(6487) <= a;
    layer5_outputs(6488) <= b;
    layer5_outputs(6489) <= '0';
    layer5_outputs(6490) <= not a;
    layer5_outputs(6491) <= a;
    layer5_outputs(6492) <= not (a or b);
    layer5_outputs(6493) <= not b or a;
    layer5_outputs(6494) <= a;
    layer5_outputs(6495) <= not b or a;
    layer5_outputs(6496) <= not b;
    layer5_outputs(6497) <= not (a and b);
    layer5_outputs(6498) <= not a or b;
    layer5_outputs(6499) <= not a or b;
    layer5_outputs(6500) <= a;
    layer5_outputs(6501) <= a or b;
    layer5_outputs(6502) <= a xor b;
    layer5_outputs(6503) <= a and b;
    layer5_outputs(6504) <= not b;
    layer5_outputs(6505) <= b;
    layer5_outputs(6506) <= b;
    layer5_outputs(6507) <= not b;
    layer5_outputs(6508) <= a;
    layer5_outputs(6509) <= a or b;
    layer5_outputs(6510) <= not a;
    layer5_outputs(6511) <= a;
    layer5_outputs(6512) <= a;
    layer5_outputs(6513) <= a and not b;
    layer5_outputs(6514) <= not (a or b);
    layer5_outputs(6515) <= b;
    layer5_outputs(6516) <= not b;
    layer5_outputs(6517) <= a xor b;
    layer5_outputs(6518) <= a and not b;
    layer5_outputs(6519) <= '1';
    layer5_outputs(6520) <= not a or b;
    layer5_outputs(6521) <= b;
    layer5_outputs(6522) <= not a;
    layer5_outputs(6523) <= not (a or b);
    layer5_outputs(6524) <= not (a xor b);
    layer5_outputs(6525) <= '0';
    layer5_outputs(6526) <= a;
    layer5_outputs(6527) <= a;
    layer5_outputs(6528) <= not (a and b);
    layer5_outputs(6529) <= a or b;
    layer5_outputs(6530) <= not (a and b);
    layer5_outputs(6531) <= a;
    layer5_outputs(6532) <= a xor b;
    layer5_outputs(6533) <= a;
    layer5_outputs(6534) <= a or b;
    layer5_outputs(6535) <= a or b;
    layer5_outputs(6536) <= not (a or b);
    layer5_outputs(6537) <= a;
    layer5_outputs(6538) <= b and not a;
    layer5_outputs(6539) <= '1';
    layer5_outputs(6540) <= b and not a;
    layer5_outputs(6541) <= b and not a;
    layer5_outputs(6542) <= not b or a;
    layer5_outputs(6543) <= not a or b;
    layer5_outputs(6544) <= not a or b;
    layer5_outputs(6545) <= not (a and b);
    layer5_outputs(6546) <= '1';
    layer5_outputs(6547) <= '1';
    layer5_outputs(6548) <= not (a or b);
    layer5_outputs(6549) <= not b;
    layer5_outputs(6550) <= a and b;
    layer5_outputs(6551) <= a or b;
    layer5_outputs(6552) <= a;
    layer5_outputs(6553) <= not b;
    layer5_outputs(6554) <= not a;
    layer5_outputs(6555) <= a or b;
    layer5_outputs(6556) <= not a or b;
    layer5_outputs(6557) <= a;
    layer5_outputs(6558) <= a and b;
    layer5_outputs(6559) <= a;
    layer5_outputs(6560) <= a and b;
    layer5_outputs(6561) <= b and not a;
    layer5_outputs(6562) <= not b;
    layer5_outputs(6563) <= a and b;
    layer5_outputs(6564) <= not (a or b);
    layer5_outputs(6565) <= a;
    layer5_outputs(6566) <= not b;
    layer5_outputs(6567) <= '1';
    layer5_outputs(6568) <= b;
    layer5_outputs(6569) <= not a or b;
    layer5_outputs(6570) <= a and not b;
    layer5_outputs(6571) <= not a;
    layer5_outputs(6572) <= not b or a;
    layer5_outputs(6573) <= '1';
    layer5_outputs(6574) <= a;
    layer5_outputs(6575) <= a;
    layer5_outputs(6576) <= not a or b;
    layer5_outputs(6577) <= a or b;
    layer5_outputs(6578) <= a and not b;
    layer5_outputs(6579) <= a and b;
    layer5_outputs(6580) <= a;
    layer5_outputs(6581) <= b and not a;
    layer5_outputs(6582) <= not (a or b);
    layer5_outputs(6583) <= a and b;
    layer5_outputs(6584) <= a and not b;
    layer5_outputs(6585) <= not b;
    layer5_outputs(6586) <= a;
    layer5_outputs(6587) <= a and not b;
    layer5_outputs(6588) <= '0';
    layer5_outputs(6589) <= not b or a;
    layer5_outputs(6590) <= not (a xor b);
    layer5_outputs(6591) <= not a or b;
    layer5_outputs(6592) <= b;
    layer5_outputs(6593) <= a or b;
    layer5_outputs(6594) <= a;
    layer5_outputs(6595) <= not a or b;
    layer5_outputs(6596) <= a and not b;
    layer5_outputs(6597) <= '1';
    layer5_outputs(6598) <= b;
    layer5_outputs(6599) <= b;
    layer5_outputs(6600) <= b;
    layer5_outputs(6601) <= not (a or b);
    layer5_outputs(6602) <= '0';
    layer5_outputs(6603) <= not b;
    layer5_outputs(6604) <= b;
    layer5_outputs(6605) <= not (a and b);
    layer5_outputs(6606) <= a and b;
    layer5_outputs(6607) <= not (a and b);
    layer5_outputs(6608) <= a and not b;
    layer5_outputs(6609) <= a;
    layer5_outputs(6610) <= not b;
    layer5_outputs(6611) <= a and not b;
    layer5_outputs(6612) <= not a or b;
    layer5_outputs(6613) <= a and not b;
    layer5_outputs(6614) <= b;
    layer5_outputs(6615) <= a and not b;
    layer5_outputs(6616) <= not a;
    layer5_outputs(6617) <= a;
    layer5_outputs(6618) <= a or b;
    layer5_outputs(6619) <= b;
    layer5_outputs(6620) <= not a;
    layer5_outputs(6621) <= a or b;
    layer5_outputs(6622) <= not (a and b);
    layer5_outputs(6623) <= b;
    layer5_outputs(6624) <= not b;
    layer5_outputs(6625) <= b and not a;
    layer5_outputs(6626) <= a;
    layer5_outputs(6627) <= not (a and b);
    layer5_outputs(6628) <= not a or b;
    layer5_outputs(6629) <= b;
    layer5_outputs(6630) <= a;
    layer5_outputs(6631) <= a or b;
    layer5_outputs(6632) <= a or b;
    layer5_outputs(6633) <= not (a or b);
    layer5_outputs(6634) <= a xor b;
    layer5_outputs(6635) <= a or b;
    layer5_outputs(6636) <= '0';
    layer5_outputs(6637) <= a and b;
    layer5_outputs(6638) <= not (a and b);
    layer5_outputs(6639) <= not a;
    layer5_outputs(6640) <= a;
    layer5_outputs(6641) <= not b;
    layer5_outputs(6642) <= a;
    layer5_outputs(6643) <= a;
    layer5_outputs(6644) <= a;
    layer5_outputs(6645) <= not (a xor b);
    layer5_outputs(6646) <= not a or b;
    layer5_outputs(6647) <= not a;
    layer5_outputs(6648) <= a and not b;
    layer5_outputs(6649) <= not b;
    layer5_outputs(6650) <= not a or b;
    layer5_outputs(6651) <= not a;
    layer5_outputs(6652) <= '1';
    layer5_outputs(6653) <= a and not b;
    layer5_outputs(6654) <= a and b;
    layer5_outputs(6655) <= not (a xor b);
    layer5_outputs(6656) <= not (a and b);
    layer5_outputs(6657) <= not a;
    layer5_outputs(6658) <= not (a and b);
    layer5_outputs(6659) <= a or b;
    layer5_outputs(6660) <= not (a or b);
    layer5_outputs(6661) <= a and not b;
    layer5_outputs(6662) <= '1';
    layer5_outputs(6663) <= not b or a;
    layer5_outputs(6664) <= '1';
    layer5_outputs(6665) <= a or b;
    layer5_outputs(6666) <= b and not a;
    layer5_outputs(6667) <= not (a or b);
    layer5_outputs(6668) <= not (a xor b);
    layer5_outputs(6669) <= a or b;
    layer5_outputs(6670) <= not (a xor b);
    layer5_outputs(6671) <= b and not a;
    layer5_outputs(6672) <= not b;
    layer5_outputs(6673) <= b;
    layer5_outputs(6674) <= a and b;
    layer5_outputs(6675) <= a or b;
    layer5_outputs(6676) <= not b or a;
    layer5_outputs(6677) <= a and not b;
    layer5_outputs(6678) <= not b or a;
    layer5_outputs(6679) <= a and not b;
    layer5_outputs(6680) <= '1';
    layer5_outputs(6681) <= not (a and b);
    layer5_outputs(6682) <= not (a and b);
    layer5_outputs(6683) <= b;
    layer5_outputs(6684) <= a and b;
    layer5_outputs(6685) <= a and not b;
    layer5_outputs(6686) <= b;
    layer5_outputs(6687) <= not b or a;
    layer5_outputs(6688) <= '0';
    layer5_outputs(6689) <= a or b;
    layer5_outputs(6690) <= a;
    layer5_outputs(6691) <= a or b;
    layer5_outputs(6692) <= not b or a;
    layer5_outputs(6693) <= '1';
    layer5_outputs(6694) <= a;
    layer5_outputs(6695) <= not b or a;
    layer5_outputs(6696) <= not (a xor b);
    layer5_outputs(6697) <= not (a xor b);
    layer5_outputs(6698) <= not (a or b);
    layer5_outputs(6699) <= a and b;
    layer5_outputs(6700) <= not a or b;
    layer5_outputs(6701) <= b and not a;
    layer5_outputs(6702) <= a;
    layer5_outputs(6703) <= '1';
    layer5_outputs(6704) <= '1';
    layer5_outputs(6705) <= a and not b;
    layer5_outputs(6706) <= b;
    layer5_outputs(6707) <= not (a and b);
    layer5_outputs(6708) <= not (a xor b);
    layer5_outputs(6709) <= '1';
    layer5_outputs(6710) <= b and not a;
    layer5_outputs(6711) <= b and not a;
    layer5_outputs(6712) <= b;
    layer5_outputs(6713) <= not a or b;
    layer5_outputs(6714) <= not b;
    layer5_outputs(6715) <= b and not a;
    layer5_outputs(6716) <= a or b;
    layer5_outputs(6717) <= not (a xor b);
    layer5_outputs(6718) <= '1';
    layer5_outputs(6719) <= not (a and b);
    layer5_outputs(6720) <= not (a or b);
    layer5_outputs(6721) <= a xor b;
    layer5_outputs(6722) <= b;
    layer5_outputs(6723) <= not a or b;
    layer5_outputs(6724) <= a and b;
    layer5_outputs(6725) <= not b;
    layer5_outputs(6726) <= a xor b;
    layer5_outputs(6727) <= b;
    layer5_outputs(6728) <= a or b;
    layer5_outputs(6729) <= not (a and b);
    layer5_outputs(6730) <= a;
    layer5_outputs(6731) <= a;
    layer5_outputs(6732) <= a xor b;
    layer5_outputs(6733) <= not b;
    layer5_outputs(6734) <= not a or b;
    layer5_outputs(6735) <= not (a or b);
    layer5_outputs(6736) <= not a;
    layer5_outputs(6737) <= not b or a;
    layer5_outputs(6738) <= not (a and b);
    layer5_outputs(6739) <= not b;
    layer5_outputs(6740) <= not b;
    layer5_outputs(6741) <= b and not a;
    layer5_outputs(6742) <= not b;
    layer5_outputs(6743) <= not b;
    layer5_outputs(6744) <= not b;
    layer5_outputs(6745) <= b;
    layer5_outputs(6746) <= a and b;
    layer5_outputs(6747) <= not (a and b);
    layer5_outputs(6748) <= b;
    layer5_outputs(6749) <= b;
    layer5_outputs(6750) <= not (a and b);
    layer5_outputs(6751) <= '1';
    layer5_outputs(6752) <= not b;
    layer5_outputs(6753) <= not (a xor b);
    layer5_outputs(6754) <= '1';
    layer5_outputs(6755) <= b and not a;
    layer5_outputs(6756) <= not b;
    layer5_outputs(6757) <= not (a xor b);
    layer5_outputs(6758) <= a xor b;
    layer5_outputs(6759) <= a and b;
    layer5_outputs(6760) <= a;
    layer5_outputs(6761) <= not b;
    layer5_outputs(6762) <= a and not b;
    layer5_outputs(6763) <= not a;
    layer5_outputs(6764) <= not b;
    layer5_outputs(6765) <= b;
    layer5_outputs(6766) <= not b or a;
    layer5_outputs(6767) <= not a or b;
    layer5_outputs(6768) <= '1';
    layer5_outputs(6769) <= not (a xor b);
    layer5_outputs(6770) <= not a or b;
    layer5_outputs(6771) <= a and not b;
    layer5_outputs(6772) <= not b or a;
    layer5_outputs(6773) <= b;
    layer5_outputs(6774) <= not a or b;
    layer5_outputs(6775) <= not a or b;
    layer5_outputs(6776) <= a and b;
    layer5_outputs(6777) <= not a;
    layer5_outputs(6778) <= b;
    layer5_outputs(6779) <= not (a and b);
    layer5_outputs(6780) <= a xor b;
    layer5_outputs(6781) <= a and not b;
    layer5_outputs(6782) <= not (a or b);
    layer5_outputs(6783) <= a;
    layer5_outputs(6784) <= a and not b;
    layer5_outputs(6785) <= '1';
    layer5_outputs(6786) <= a xor b;
    layer5_outputs(6787) <= a and not b;
    layer5_outputs(6788) <= a;
    layer5_outputs(6789) <= not a;
    layer5_outputs(6790) <= not a;
    layer5_outputs(6791) <= a and not b;
    layer5_outputs(6792) <= a and b;
    layer5_outputs(6793) <= not (a or b);
    layer5_outputs(6794) <= not a;
    layer5_outputs(6795) <= a and not b;
    layer5_outputs(6796) <= '0';
    layer5_outputs(6797) <= not (a and b);
    layer5_outputs(6798) <= a;
    layer5_outputs(6799) <= b;
    layer5_outputs(6800) <= '0';
    layer5_outputs(6801) <= a xor b;
    layer5_outputs(6802) <= not (a and b);
    layer5_outputs(6803) <= a and b;
    layer5_outputs(6804) <= b and not a;
    layer5_outputs(6805) <= not a;
    layer5_outputs(6806) <= a and b;
    layer5_outputs(6807) <= '1';
    layer5_outputs(6808) <= not a;
    layer5_outputs(6809) <= b and not a;
    layer5_outputs(6810) <= not b;
    layer5_outputs(6811) <= a and not b;
    layer5_outputs(6812) <= a;
    layer5_outputs(6813) <= b;
    layer5_outputs(6814) <= not (a xor b);
    layer5_outputs(6815) <= a and b;
    layer5_outputs(6816) <= a or b;
    layer5_outputs(6817) <= not (a or b);
    layer5_outputs(6818) <= '1';
    layer5_outputs(6819) <= not (a and b);
    layer5_outputs(6820) <= b;
    layer5_outputs(6821) <= '0';
    layer5_outputs(6822) <= '1';
    layer5_outputs(6823) <= not a or b;
    layer5_outputs(6824) <= not a or b;
    layer5_outputs(6825) <= not (a or b);
    layer5_outputs(6826) <= not b;
    layer5_outputs(6827) <= not (a xor b);
    layer5_outputs(6828) <= not b or a;
    layer5_outputs(6829) <= not b;
    layer5_outputs(6830) <= not (a or b);
    layer5_outputs(6831) <= not b or a;
    layer5_outputs(6832) <= b and not a;
    layer5_outputs(6833) <= not a or b;
    layer5_outputs(6834) <= a and b;
    layer5_outputs(6835) <= not (a or b);
    layer5_outputs(6836) <= a and b;
    layer5_outputs(6837) <= not a;
    layer5_outputs(6838) <= not (a xor b);
    layer5_outputs(6839) <= not (a and b);
    layer5_outputs(6840) <= a xor b;
    layer5_outputs(6841) <= not (a or b);
    layer5_outputs(6842) <= not a or b;
    layer5_outputs(6843) <= a and b;
    layer5_outputs(6844) <= a and b;
    layer5_outputs(6845) <= not a;
    layer5_outputs(6846) <= not a;
    layer5_outputs(6847) <= a and b;
    layer5_outputs(6848) <= a and not b;
    layer5_outputs(6849) <= '1';
    layer5_outputs(6850) <= b;
    layer5_outputs(6851) <= not b;
    layer5_outputs(6852) <= a or b;
    layer5_outputs(6853) <= a or b;
    layer5_outputs(6854) <= '1';
    layer5_outputs(6855) <= b;
    layer5_outputs(6856) <= a and b;
    layer5_outputs(6857) <= b;
    layer5_outputs(6858) <= not (a and b);
    layer5_outputs(6859) <= not (a or b);
    layer5_outputs(6860) <= not b or a;
    layer5_outputs(6861) <= not a;
    layer5_outputs(6862) <= a;
    layer5_outputs(6863) <= b and not a;
    layer5_outputs(6864) <= not b or a;
    layer5_outputs(6865) <= a xor b;
    layer5_outputs(6866) <= a xor b;
    layer5_outputs(6867) <= not a or b;
    layer5_outputs(6868) <= b and not a;
    layer5_outputs(6869) <= a and not b;
    layer5_outputs(6870) <= a;
    layer5_outputs(6871) <= not a or b;
    layer5_outputs(6872) <= b and not a;
    layer5_outputs(6873) <= a and b;
    layer5_outputs(6874) <= not b;
    layer5_outputs(6875) <= not b;
    layer5_outputs(6876) <= not a;
    layer5_outputs(6877) <= not a;
    layer5_outputs(6878) <= not (a xor b);
    layer5_outputs(6879) <= not a;
    layer5_outputs(6880) <= not a;
    layer5_outputs(6881) <= a and b;
    layer5_outputs(6882) <= a;
    layer5_outputs(6883) <= not b;
    layer5_outputs(6884) <= not a or b;
    layer5_outputs(6885) <= not b;
    layer5_outputs(6886) <= not (a or b);
    layer5_outputs(6887) <= not b or a;
    layer5_outputs(6888) <= b and not a;
    layer5_outputs(6889) <= not a;
    layer5_outputs(6890) <= '1';
    layer5_outputs(6891) <= b;
    layer5_outputs(6892) <= a and not b;
    layer5_outputs(6893) <= b and not a;
    layer5_outputs(6894) <= a xor b;
    layer5_outputs(6895) <= not b;
    layer5_outputs(6896) <= a or b;
    layer5_outputs(6897) <= not (a and b);
    layer5_outputs(6898) <= not b;
    layer5_outputs(6899) <= not (a or b);
    layer5_outputs(6900) <= not a;
    layer5_outputs(6901) <= not (a xor b);
    layer5_outputs(6902) <= a and b;
    layer5_outputs(6903) <= b;
    layer5_outputs(6904) <= a or b;
    layer5_outputs(6905) <= a;
    layer5_outputs(6906) <= b and not a;
    layer5_outputs(6907) <= not b;
    layer5_outputs(6908) <= a and b;
    layer5_outputs(6909) <= not a;
    layer5_outputs(6910) <= a;
    layer5_outputs(6911) <= not (a and b);
    layer5_outputs(6912) <= not (a and b);
    layer5_outputs(6913) <= not a;
    layer5_outputs(6914) <= a;
    layer5_outputs(6915) <= not a;
    layer5_outputs(6916) <= b;
    layer5_outputs(6917) <= not b;
    layer5_outputs(6918) <= b;
    layer5_outputs(6919) <= b;
    layer5_outputs(6920) <= not (a xor b);
    layer5_outputs(6921) <= a and b;
    layer5_outputs(6922) <= a and b;
    layer5_outputs(6923) <= not (a and b);
    layer5_outputs(6924) <= not (a or b);
    layer5_outputs(6925) <= not a or b;
    layer5_outputs(6926) <= a and b;
    layer5_outputs(6927) <= a;
    layer5_outputs(6928) <= a and not b;
    layer5_outputs(6929) <= not a or b;
    layer5_outputs(6930) <= not (a and b);
    layer5_outputs(6931) <= not b or a;
    layer5_outputs(6932) <= a;
    layer5_outputs(6933) <= a and b;
    layer5_outputs(6934) <= not (a or b);
    layer5_outputs(6935) <= not (a or b);
    layer5_outputs(6936) <= '0';
    layer5_outputs(6937) <= '1';
    layer5_outputs(6938) <= not a;
    layer5_outputs(6939) <= not b or a;
    layer5_outputs(6940) <= b and not a;
    layer5_outputs(6941) <= a or b;
    layer5_outputs(6942) <= not (a and b);
    layer5_outputs(6943) <= a xor b;
    layer5_outputs(6944) <= a xor b;
    layer5_outputs(6945) <= a xor b;
    layer5_outputs(6946) <= b and not a;
    layer5_outputs(6947) <= not a or b;
    layer5_outputs(6948) <= a;
    layer5_outputs(6949) <= a and not b;
    layer5_outputs(6950) <= not (a and b);
    layer5_outputs(6951) <= b;
    layer5_outputs(6952) <= a;
    layer5_outputs(6953) <= a;
    layer5_outputs(6954) <= not (a or b);
    layer5_outputs(6955) <= a or b;
    layer5_outputs(6956) <= a;
    layer5_outputs(6957) <= not b;
    layer5_outputs(6958) <= a and b;
    layer5_outputs(6959) <= b and not a;
    layer5_outputs(6960) <= not a;
    layer5_outputs(6961) <= a and not b;
    layer5_outputs(6962) <= not b;
    layer5_outputs(6963) <= b and not a;
    layer5_outputs(6964) <= a and not b;
    layer5_outputs(6965) <= not b;
    layer5_outputs(6966) <= not a or b;
    layer5_outputs(6967) <= '1';
    layer5_outputs(6968) <= '0';
    layer5_outputs(6969) <= a;
    layer5_outputs(6970) <= not a or b;
    layer5_outputs(6971) <= not b;
    layer5_outputs(6972) <= a and b;
    layer5_outputs(6973) <= '1';
    layer5_outputs(6974) <= a;
    layer5_outputs(6975) <= not b or a;
    layer5_outputs(6976) <= b;
    layer5_outputs(6977) <= not (a xor b);
    layer5_outputs(6978) <= a;
    layer5_outputs(6979) <= a and b;
    layer5_outputs(6980) <= not b;
    layer5_outputs(6981) <= a;
    layer5_outputs(6982) <= '1';
    layer5_outputs(6983) <= not (a and b);
    layer5_outputs(6984) <= not a;
    layer5_outputs(6985) <= a;
    layer5_outputs(6986) <= a and not b;
    layer5_outputs(6987) <= a or b;
    layer5_outputs(6988) <= b;
    layer5_outputs(6989) <= not b or a;
    layer5_outputs(6990) <= not (a and b);
    layer5_outputs(6991) <= not (a xor b);
    layer5_outputs(6992) <= b and not a;
    layer5_outputs(6993) <= a and not b;
    layer5_outputs(6994) <= a and not b;
    layer5_outputs(6995) <= b;
    layer5_outputs(6996) <= a or b;
    layer5_outputs(6997) <= '0';
    layer5_outputs(6998) <= not (a and b);
    layer5_outputs(6999) <= a xor b;
    layer5_outputs(7000) <= a and not b;
    layer5_outputs(7001) <= not b;
    layer5_outputs(7002) <= a;
    layer5_outputs(7003) <= not (a xor b);
    layer5_outputs(7004) <= b;
    layer5_outputs(7005) <= a;
    layer5_outputs(7006) <= not a;
    layer5_outputs(7007) <= not a;
    layer5_outputs(7008) <= not b or a;
    layer5_outputs(7009) <= not b or a;
    layer5_outputs(7010) <= not b;
    layer5_outputs(7011) <= not (a or b);
    layer5_outputs(7012) <= b and not a;
    layer5_outputs(7013) <= not (a or b);
    layer5_outputs(7014) <= not a;
    layer5_outputs(7015) <= a and not b;
    layer5_outputs(7016) <= not (a and b);
    layer5_outputs(7017) <= not (a xor b);
    layer5_outputs(7018) <= a;
    layer5_outputs(7019) <= b and not a;
    layer5_outputs(7020) <= b and not a;
    layer5_outputs(7021) <= not (a and b);
    layer5_outputs(7022) <= a or b;
    layer5_outputs(7023) <= '0';
    layer5_outputs(7024) <= not a;
    layer5_outputs(7025) <= not b;
    layer5_outputs(7026) <= not a;
    layer5_outputs(7027) <= a and not b;
    layer5_outputs(7028) <= not b;
    layer5_outputs(7029) <= a and not b;
    layer5_outputs(7030) <= not (a xor b);
    layer5_outputs(7031) <= not a or b;
    layer5_outputs(7032) <= a or b;
    layer5_outputs(7033) <= not a;
    layer5_outputs(7034) <= '1';
    layer5_outputs(7035) <= b and not a;
    layer5_outputs(7036) <= not a;
    layer5_outputs(7037) <= a xor b;
    layer5_outputs(7038) <= a;
    layer5_outputs(7039) <= not b or a;
    layer5_outputs(7040) <= a;
    layer5_outputs(7041) <= a and b;
    layer5_outputs(7042) <= not a;
    layer5_outputs(7043) <= a or b;
    layer5_outputs(7044) <= a and b;
    layer5_outputs(7045) <= '1';
    layer5_outputs(7046) <= a and not b;
    layer5_outputs(7047) <= '1';
    layer5_outputs(7048) <= not a;
    layer5_outputs(7049) <= b;
    layer5_outputs(7050) <= a xor b;
    layer5_outputs(7051) <= not a;
    layer5_outputs(7052) <= not a;
    layer5_outputs(7053) <= b;
    layer5_outputs(7054) <= a and not b;
    layer5_outputs(7055) <= a;
    layer5_outputs(7056) <= not (a xor b);
    layer5_outputs(7057) <= not a or b;
    layer5_outputs(7058) <= not b or a;
    layer5_outputs(7059) <= not (a or b);
    layer5_outputs(7060) <= a or b;
    layer5_outputs(7061) <= a and not b;
    layer5_outputs(7062) <= '0';
    layer5_outputs(7063) <= b;
    layer5_outputs(7064) <= a xor b;
    layer5_outputs(7065) <= a or b;
    layer5_outputs(7066) <= not (a xor b);
    layer5_outputs(7067) <= a and not b;
    layer5_outputs(7068) <= '1';
    layer5_outputs(7069) <= '1';
    layer5_outputs(7070) <= not a;
    layer5_outputs(7071) <= not b or a;
    layer5_outputs(7072) <= b and not a;
    layer5_outputs(7073) <= a or b;
    layer5_outputs(7074) <= b;
    layer5_outputs(7075) <= a and not b;
    layer5_outputs(7076) <= b and not a;
    layer5_outputs(7077) <= not a or b;
    layer5_outputs(7078) <= not a or b;
    layer5_outputs(7079) <= not (a and b);
    layer5_outputs(7080) <= not b or a;
    layer5_outputs(7081) <= b;
    layer5_outputs(7082) <= b;
    layer5_outputs(7083) <= a;
    layer5_outputs(7084) <= a;
    layer5_outputs(7085) <= a and b;
    layer5_outputs(7086) <= not b or a;
    layer5_outputs(7087) <= not a;
    layer5_outputs(7088) <= not a;
    layer5_outputs(7089) <= not (a or b);
    layer5_outputs(7090) <= '1';
    layer5_outputs(7091) <= a;
    layer5_outputs(7092) <= a and b;
    layer5_outputs(7093) <= b;
    layer5_outputs(7094) <= a or b;
    layer5_outputs(7095) <= a and b;
    layer5_outputs(7096) <= not a;
    layer5_outputs(7097) <= not (a and b);
    layer5_outputs(7098) <= a xor b;
    layer5_outputs(7099) <= a;
    layer5_outputs(7100) <= a or b;
    layer5_outputs(7101) <= a and b;
    layer5_outputs(7102) <= b;
    layer5_outputs(7103) <= a xor b;
    layer5_outputs(7104) <= b;
    layer5_outputs(7105) <= '1';
    layer5_outputs(7106) <= a;
    layer5_outputs(7107) <= '0';
    layer5_outputs(7108) <= '1';
    layer5_outputs(7109) <= '0';
    layer5_outputs(7110) <= a and b;
    layer5_outputs(7111) <= a xor b;
    layer5_outputs(7112) <= a or b;
    layer5_outputs(7113) <= a;
    layer5_outputs(7114) <= b and not a;
    layer5_outputs(7115) <= a and not b;
    layer5_outputs(7116) <= b;
    layer5_outputs(7117) <= not a;
    layer5_outputs(7118) <= not b;
    layer5_outputs(7119) <= a and b;
    layer5_outputs(7120) <= a or b;
    layer5_outputs(7121) <= not (a and b);
    layer5_outputs(7122) <= not (a or b);
    layer5_outputs(7123) <= a and b;
    layer5_outputs(7124) <= a and not b;
    layer5_outputs(7125) <= a xor b;
    layer5_outputs(7126) <= a;
    layer5_outputs(7127) <= a;
    layer5_outputs(7128) <= a xor b;
    layer5_outputs(7129) <= a and b;
    layer5_outputs(7130) <= not (a or b);
    layer5_outputs(7131) <= not a;
    layer5_outputs(7132) <= a and b;
    layer5_outputs(7133) <= a and b;
    layer5_outputs(7134) <= b;
    layer5_outputs(7135) <= not a or b;
    layer5_outputs(7136) <= not a;
    layer5_outputs(7137) <= not (a or b);
    layer5_outputs(7138) <= not b or a;
    layer5_outputs(7139) <= a and b;
    layer5_outputs(7140) <= not a or b;
    layer5_outputs(7141) <= b;
    layer5_outputs(7142) <= b;
    layer5_outputs(7143) <= b;
    layer5_outputs(7144) <= '0';
    layer5_outputs(7145) <= not a or b;
    layer5_outputs(7146) <= a or b;
    layer5_outputs(7147) <= a and b;
    layer5_outputs(7148) <= '1';
    layer5_outputs(7149) <= not a;
    layer5_outputs(7150) <= not b;
    layer5_outputs(7151) <= not (a and b);
    layer5_outputs(7152) <= a and b;
    layer5_outputs(7153) <= not (a or b);
    layer5_outputs(7154) <= a and b;
    layer5_outputs(7155) <= a;
    layer5_outputs(7156) <= b;
    layer5_outputs(7157) <= not (a or b);
    layer5_outputs(7158) <= not b;
    layer5_outputs(7159) <= '1';
    layer5_outputs(7160) <= a and not b;
    layer5_outputs(7161) <= '0';
    layer5_outputs(7162) <= a and b;
    layer5_outputs(7163) <= b and not a;
    layer5_outputs(7164) <= a xor b;
    layer5_outputs(7165) <= not a;
    layer5_outputs(7166) <= a and not b;
    layer5_outputs(7167) <= a and not b;
    layer5_outputs(7168) <= not b;
    layer5_outputs(7169) <= b and not a;
    layer5_outputs(7170) <= not a or b;
    layer5_outputs(7171) <= '1';
    layer5_outputs(7172) <= '0';
    layer5_outputs(7173) <= b and not a;
    layer5_outputs(7174) <= not a;
    layer5_outputs(7175) <= not a or b;
    layer5_outputs(7176) <= a and b;
    layer5_outputs(7177) <= not (a xor b);
    layer5_outputs(7178) <= a and not b;
    layer5_outputs(7179) <= not (a or b);
    layer5_outputs(7180) <= a and b;
    layer5_outputs(7181) <= not b or a;
    layer5_outputs(7182) <= a;
    layer5_outputs(7183) <= not a;
    layer5_outputs(7184) <= a and not b;
    layer5_outputs(7185) <= not a or b;
    layer5_outputs(7186) <= not a or b;
    layer5_outputs(7187) <= not b;
    layer5_outputs(7188) <= not (a or b);
    layer5_outputs(7189) <= not b;
    layer5_outputs(7190) <= a and b;
    layer5_outputs(7191) <= not a;
    layer5_outputs(7192) <= not a or b;
    layer5_outputs(7193) <= '1';
    layer5_outputs(7194) <= b;
    layer5_outputs(7195) <= a or b;
    layer5_outputs(7196) <= a;
    layer5_outputs(7197) <= not b;
    layer5_outputs(7198) <= not a or b;
    layer5_outputs(7199) <= not (a and b);
    layer5_outputs(7200) <= not a;
    layer5_outputs(7201) <= not b or a;
    layer5_outputs(7202) <= not b;
    layer5_outputs(7203) <= not (a and b);
    layer5_outputs(7204) <= a and not b;
    layer5_outputs(7205) <= not (a xor b);
    layer5_outputs(7206) <= not a;
    layer5_outputs(7207) <= not a or b;
    layer5_outputs(7208) <= not b or a;
    layer5_outputs(7209) <= a xor b;
    layer5_outputs(7210) <= a xor b;
    layer5_outputs(7211) <= a and b;
    layer5_outputs(7212) <= a;
    layer5_outputs(7213) <= not b or a;
    layer5_outputs(7214) <= not b;
    layer5_outputs(7215) <= not (a and b);
    layer5_outputs(7216) <= a or b;
    layer5_outputs(7217) <= a and b;
    layer5_outputs(7218) <= not b or a;
    layer5_outputs(7219) <= a;
    layer5_outputs(7220) <= a and not b;
    layer5_outputs(7221) <= a or b;
    layer5_outputs(7222) <= not b or a;
    layer5_outputs(7223) <= a;
    layer5_outputs(7224) <= not b;
    layer5_outputs(7225) <= b;
    layer5_outputs(7226) <= not (a and b);
    layer5_outputs(7227) <= a;
    layer5_outputs(7228) <= a xor b;
    layer5_outputs(7229) <= a and not b;
    layer5_outputs(7230) <= a;
    layer5_outputs(7231) <= b;
    layer5_outputs(7232) <= a xor b;
    layer5_outputs(7233) <= a;
    layer5_outputs(7234) <= not b;
    layer5_outputs(7235) <= not (a and b);
    layer5_outputs(7236) <= not (a and b);
    layer5_outputs(7237) <= not b;
    layer5_outputs(7238) <= not b or a;
    layer5_outputs(7239) <= b and not a;
    layer5_outputs(7240) <= not (a and b);
    layer5_outputs(7241) <= not b;
    layer5_outputs(7242) <= b and not a;
    layer5_outputs(7243) <= a and b;
    layer5_outputs(7244) <= a;
    layer5_outputs(7245) <= not (a and b);
    layer5_outputs(7246) <= not (a and b);
    layer5_outputs(7247) <= not a or b;
    layer5_outputs(7248) <= a;
    layer5_outputs(7249) <= not (a or b);
    layer5_outputs(7250) <= a and not b;
    layer5_outputs(7251) <= not (a and b);
    layer5_outputs(7252) <= not a;
    layer5_outputs(7253) <= b;
    layer5_outputs(7254) <= a or b;
    layer5_outputs(7255) <= not b;
    layer5_outputs(7256) <= not a;
    layer5_outputs(7257) <= not b;
    layer5_outputs(7258) <= '1';
    layer5_outputs(7259) <= not (a xor b);
    layer5_outputs(7260) <= a or b;
    layer5_outputs(7261) <= not (a and b);
    layer5_outputs(7262) <= a xor b;
    layer5_outputs(7263) <= not a or b;
    layer5_outputs(7264) <= not b or a;
    layer5_outputs(7265) <= a;
    layer5_outputs(7266) <= not (a or b);
    layer5_outputs(7267) <= '1';
    layer5_outputs(7268) <= '1';
    layer5_outputs(7269) <= not a;
    layer5_outputs(7270) <= '0';
    layer5_outputs(7271) <= not a or b;
    layer5_outputs(7272) <= not (a or b);
    layer5_outputs(7273) <= not a or b;
    layer5_outputs(7274) <= '1';
    layer5_outputs(7275) <= not a;
    layer5_outputs(7276) <= not b;
    layer5_outputs(7277) <= b and not a;
    layer5_outputs(7278) <= not a;
    layer5_outputs(7279) <= a;
    layer5_outputs(7280) <= not b;
    layer5_outputs(7281) <= not (a or b);
    layer5_outputs(7282) <= not a or b;
    layer5_outputs(7283) <= a or b;
    layer5_outputs(7284) <= a;
    layer5_outputs(7285) <= a and not b;
    layer5_outputs(7286) <= not (a and b);
    layer5_outputs(7287) <= not a or b;
    layer5_outputs(7288) <= not a;
    layer5_outputs(7289) <= b;
    layer5_outputs(7290) <= not b;
    layer5_outputs(7291) <= not (a or b);
    layer5_outputs(7292) <= not b;
    layer5_outputs(7293) <= not a;
    layer5_outputs(7294) <= b;
    layer5_outputs(7295) <= a and b;
    layer5_outputs(7296) <= a and b;
    layer5_outputs(7297) <= b and not a;
    layer5_outputs(7298) <= '0';
    layer5_outputs(7299) <= '0';
    layer5_outputs(7300) <= not (a or b);
    layer5_outputs(7301) <= not b or a;
    layer5_outputs(7302) <= not b or a;
    layer5_outputs(7303) <= not a;
    layer5_outputs(7304) <= '0';
    layer5_outputs(7305) <= not a;
    layer5_outputs(7306) <= '0';
    layer5_outputs(7307) <= not b or a;
    layer5_outputs(7308) <= a and b;
    layer5_outputs(7309) <= a and not b;
    layer5_outputs(7310) <= b and not a;
    layer5_outputs(7311) <= not b or a;
    layer5_outputs(7312) <= a and not b;
    layer5_outputs(7313) <= not (a or b);
    layer5_outputs(7314) <= a;
    layer5_outputs(7315) <= not (a xor b);
    layer5_outputs(7316) <= b and not a;
    layer5_outputs(7317) <= not b;
    layer5_outputs(7318) <= a and not b;
    layer5_outputs(7319) <= not (a and b);
    layer5_outputs(7320) <= b and not a;
    layer5_outputs(7321) <= not b;
    layer5_outputs(7322) <= a xor b;
    layer5_outputs(7323) <= not (a and b);
    layer5_outputs(7324) <= a;
    layer5_outputs(7325) <= not (a and b);
    layer5_outputs(7326) <= a and b;
    layer5_outputs(7327) <= not (a xor b);
    layer5_outputs(7328) <= '1';
    layer5_outputs(7329) <= '0';
    layer5_outputs(7330) <= a and not b;
    layer5_outputs(7331) <= b;
    layer5_outputs(7332) <= a;
    layer5_outputs(7333) <= b;
    layer5_outputs(7334) <= not b;
    layer5_outputs(7335) <= not b or a;
    layer5_outputs(7336) <= b and not a;
    layer5_outputs(7337) <= not (a and b);
    layer5_outputs(7338) <= not a or b;
    layer5_outputs(7339) <= b;
    layer5_outputs(7340) <= not (a and b);
    layer5_outputs(7341) <= a;
    layer5_outputs(7342) <= not a;
    layer5_outputs(7343) <= a and b;
    layer5_outputs(7344) <= not a;
    layer5_outputs(7345) <= a;
    layer5_outputs(7346) <= a xor b;
    layer5_outputs(7347) <= not a or b;
    layer5_outputs(7348) <= not (a and b);
    layer5_outputs(7349) <= a;
    layer5_outputs(7350) <= not b or a;
    layer5_outputs(7351) <= not b or a;
    layer5_outputs(7352) <= a;
    layer5_outputs(7353) <= a and b;
    layer5_outputs(7354) <= a and not b;
    layer5_outputs(7355) <= not (a and b);
    layer5_outputs(7356) <= '0';
    layer5_outputs(7357) <= b and not a;
    layer5_outputs(7358) <= '1';
    layer5_outputs(7359) <= not a or b;
    layer5_outputs(7360) <= not (a or b);
    layer5_outputs(7361) <= b and not a;
    layer5_outputs(7362) <= b;
    layer5_outputs(7363) <= not a or b;
    layer5_outputs(7364) <= b and not a;
    layer5_outputs(7365) <= not (a xor b);
    layer5_outputs(7366) <= not (a xor b);
    layer5_outputs(7367) <= not b or a;
    layer5_outputs(7368) <= not b or a;
    layer5_outputs(7369) <= not (a and b);
    layer5_outputs(7370) <= '1';
    layer5_outputs(7371) <= b and not a;
    layer5_outputs(7372) <= '0';
    layer5_outputs(7373) <= not a;
    layer5_outputs(7374) <= not a;
    layer5_outputs(7375) <= a and not b;
    layer5_outputs(7376) <= b and not a;
    layer5_outputs(7377) <= '0';
    layer5_outputs(7378) <= a xor b;
    layer5_outputs(7379) <= not a or b;
    layer5_outputs(7380) <= b;
    layer5_outputs(7381) <= not a or b;
    layer5_outputs(7382) <= not a;
    layer5_outputs(7383) <= a and not b;
    layer5_outputs(7384) <= b;
    layer5_outputs(7385) <= b;
    layer5_outputs(7386) <= a;
    layer5_outputs(7387) <= not b;
    layer5_outputs(7388) <= not (a and b);
    layer5_outputs(7389) <= not a;
    layer5_outputs(7390) <= a and not b;
    layer5_outputs(7391) <= not b or a;
    layer5_outputs(7392) <= b and not a;
    layer5_outputs(7393) <= not a or b;
    layer5_outputs(7394) <= not b;
    layer5_outputs(7395) <= not (a and b);
    layer5_outputs(7396) <= a;
    layer5_outputs(7397) <= not a or b;
    layer5_outputs(7398) <= a or b;
    layer5_outputs(7399) <= a and not b;
    layer5_outputs(7400) <= not b or a;
    layer5_outputs(7401) <= b;
    layer5_outputs(7402) <= b;
    layer5_outputs(7403) <= a and b;
    layer5_outputs(7404) <= not a;
    layer5_outputs(7405) <= not b or a;
    layer5_outputs(7406) <= not a;
    layer5_outputs(7407) <= not b;
    layer5_outputs(7408) <= b;
    layer5_outputs(7409) <= not b or a;
    layer5_outputs(7410) <= a or b;
    layer5_outputs(7411) <= a;
    layer5_outputs(7412) <= a and b;
    layer5_outputs(7413) <= '0';
    layer5_outputs(7414) <= a and not b;
    layer5_outputs(7415) <= not (a and b);
    layer5_outputs(7416) <= not b;
    layer5_outputs(7417) <= not a or b;
    layer5_outputs(7418) <= b and not a;
    layer5_outputs(7419) <= not a;
    layer5_outputs(7420) <= not (a or b);
    layer5_outputs(7421) <= a or b;
    layer5_outputs(7422) <= not (a and b);
    layer5_outputs(7423) <= b;
    layer5_outputs(7424) <= '1';
    layer5_outputs(7425) <= '0';
    layer5_outputs(7426) <= not (a or b);
    layer5_outputs(7427) <= a or b;
    layer5_outputs(7428) <= not (a and b);
    layer5_outputs(7429) <= b and not a;
    layer5_outputs(7430) <= a;
    layer5_outputs(7431) <= not (a or b);
    layer5_outputs(7432) <= not (a xor b);
    layer5_outputs(7433) <= b and not a;
    layer5_outputs(7434) <= a;
    layer5_outputs(7435) <= not b;
    layer5_outputs(7436) <= a;
    layer5_outputs(7437) <= b and not a;
    layer5_outputs(7438) <= b;
    layer5_outputs(7439) <= b and not a;
    layer5_outputs(7440) <= a;
    layer5_outputs(7441) <= '0';
    layer5_outputs(7442) <= not a;
    layer5_outputs(7443) <= a or b;
    layer5_outputs(7444) <= '0';
    layer5_outputs(7445) <= b and not a;
    layer5_outputs(7446) <= not (a and b);
    layer5_outputs(7447) <= b and not a;
    layer5_outputs(7448) <= not a or b;
    layer5_outputs(7449) <= a and not b;
    layer5_outputs(7450) <= not a or b;
    layer5_outputs(7451) <= not a;
    layer5_outputs(7452) <= not a or b;
    layer5_outputs(7453) <= not a;
    layer5_outputs(7454) <= not a;
    layer5_outputs(7455) <= not b;
    layer5_outputs(7456) <= '0';
    layer5_outputs(7457) <= not (a or b);
    layer5_outputs(7458) <= not b;
    layer5_outputs(7459) <= a and not b;
    layer5_outputs(7460) <= a;
    layer5_outputs(7461) <= a;
    layer5_outputs(7462) <= a;
    layer5_outputs(7463) <= not a or b;
    layer5_outputs(7464) <= a;
    layer5_outputs(7465) <= not (a or b);
    layer5_outputs(7466) <= b;
    layer5_outputs(7467) <= a xor b;
    layer5_outputs(7468) <= a and b;
    layer5_outputs(7469) <= not (a and b);
    layer5_outputs(7470) <= not a;
    layer5_outputs(7471) <= a and not b;
    layer5_outputs(7472) <= a and b;
    layer5_outputs(7473) <= not b;
    layer5_outputs(7474) <= not (a and b);
    layer5_outputs(7475) <= '0';
    layer5_outputs(7476) <= a;
    layer5_outputs(7477) <= '1';
    layer5_outputs(7478) <= not (a and b);
    layer5_outputs(7479) <= b;
    layer5_outputs(7480) <= b;
    layer5_outputs(7481) <= a and b;
    layer5_outputs(7482) <= a xor b;
    layer5_outputs(7483) <= b;
    layer5_outputs(7484) <= not (a xor b);
    layer5_outputs(7485) <= not a;
    layer5_outputs(7486) <= a;
    layer5_outputs(7487) <= b and not a;
    layer5_outputs(7488) <= not a;
    layer5_outputs(7489) <= not b or a;
    layer5_outputs(7490) <= a;
    layer5_outputs(7491) <= not (a and b);
    layer5_outputs(7492) <= a;
    layer5_outputs(7493) <= not b;
    layer5_outputs(7494) <= a or b;
    layer5_outputs(7495) <= b;
    layer5_outputs(7496) <= not (a or b);
    layer5_outputs(7497) <= not b or a;
    layer5_outputs(7498) <= not b;
    layer5_outputs(7499) <= not a or b;
    layer5_outputs(7500) <= '0';
    layer5_outputs(7501) <= a and not b;
    layer5_outputs(7502) <= not a;
    layer5_outputs(7503) <= not (a xor b);
    layer5_outputs(7504) <= not a;
    layer5_outputs(7505) <= b;
    layer5_outputs(7506) <= a and b;
    layer5_outputs(7507) <= a and not b;
    layer5_outputs(7508) <= not (a xor b);
    layer5_outputs(7509) <= a or b;
    layer5_outputs(7510) <= a or b;
    layer5_outputs(7511) <= not a;
    layer5_outputs(7512) <= not b;
    layer5_outputs(7513) <= not a;
    layer5_outputs(7514) <= not a or b;
    layer5_outputs(7515) <= '1';
    layer5_outputs(7516) <= '1';
    layer5_outputs(7517) <= b and not a;
    layer5_outputs(7518) <= not (a and b);
    layer5_outputs(7519) <= a;
    layer5_outputs(7520) <= a and b;
    layer5_outputs(7521) <= not b or a;
    layer5_outputs(7522) <= a;
    layer5_outputs(7523) <= not a or b;
    layer5_outputs(7524) <= not (a or b);
    layer5_outputs(7525) <= not (a xor b);
    layer5_outputs(7526) <= a;
    layer5_outputs(7527) <= not (a or b);
    layer5_outputs(7528) <= not a or b;
    layer5_outputs(7529) <= a and b;
    layer5_outputs(7530) <= a and not b;
    layer5_outputs(7531) <= not b;
    layer5_outputs(7532) <= not b;
    layer5_outputs(7533) <= not a;
    layer5_outputs(7534) <= b and not a;
    layer5_outputs(7535) <= a;
    layer5_outputs(7536) <= not a or b;
    layer5_outputs(7537) <= a and b;
    layer5_outputs(7538) <= not (a and b);
    layer5_outputs(7539) <= a and not b;
    layer5_outputs(7540) <= a;
    layer5_outputs(7541) <= not (a and b);
    layer5_outputs(7542) <= not (a or b);
    layer5_outputs(7543) <= not (a xor b);
    layer5_outputs(7544) <= b;
    layer5_outputs(7545) <= b;
    layer5_outputs(7546) <= a and not b;
    layer5_outputs(7547) <= b;
    layer5_outputs(7548) <= not b;
    layer5_outputs(7549) <= '0';
    layer5_outputs(7550) <= '0';
    layer5_outputs(7551) <= b and not a;
    layer5_outputs(7552) <= not (a or b);
    layer5_outputs(7553) <= a and b;
    layer5_outputs(7554) <= not (a xor b);
    layer5_outputs(7555) <= not a or b;
    layer5_outputs(7556) <= a and b;
    layer5_outputs(7557) <= '0';
    layer5_outputs(7558) <= '0';
    layer5_outputs(7559) <= b and not a;
    layer5_outputs(7560) <= b;
    layer5_outputs(7561) <= a;
    layer5_outputs(7562) <= not (a or b);
    layer5_outputs(7563) <= not (a or b);
    layer5_outputs(7564) <= a or b;
    layer5_outputs(7565) <= a and not b;
    layer5_outputs(7566) <= a and b;
    layer5_outputs(7567) <= b and not a;
    layer5_outputs(7568) <= a;
    layer5_outputs(7569) <= not (a or b);
    layer5_outputs(7570) <= not b or a;
    layer5_outputs(7571) <= not b;
    layer5_outputs(7572) <= a and b;
    layer5_outputs(7573) <= '1';
    layer5_outputs(7574) <= '0';
    layer5_outputs(7575) <= not b or a;
    layer5_outputs(7576) <= not (a or b);
    layer5_outputs(7577) <= not (a or b);
    layer5_outputs(7578) <= a or b;
    layer5_outputs(7579) <= '0';
    layer5_outputs(7580) <= not (a or b);
    layer5_outputs(7581) <= b;
    layer5_outputs(7582) <= b and not a;
    layer5_outputs(7583) <= '1';
    layer5_outputs(7584) <= not b or a;
    layer5_outputs(7585) <= not (a and b);
    layer5_outputs(7586) <= b and not a;
    layer5_outputs(7587) <= not a or b;
    layer5_outputs(7588) <= b;
    layer5_outputs(7589) <= not b or a;
    layer5_outputs(7590) <= not a;
    layer5_outputs(7591) <= a xor b;
    layer5_outputs(7592) <= not a or b;
    layer5_outputs(7593) <= not a;
    layer5_outputs(7594) <= a;
    layer5_outputs(7595) <= not b or a;
    layer5_outputs(7596) <= a or b;
    layer5_outputs(7597) <= not (a xor b);
    layer5_outputs(7598) <= a and not b;
    layer5_outputs(7599) <= not (a and b);
    layer5_outputs(7600) <= not a;
    layer5_outputs(7601) <= a and not b;
    layer5_outputs(7602) <= a;
    layer5_outputs(7603) <= not a;
    layer5_outputs(7604) <= b and not a;
    layer5_outputs(7605) <= '0';
    layer5_outputs(7606) <= not (a or b);
    layer5_outputs(7607) <= '0';
    layer5_outputs(7608) <= not a;
    layer5_outputs(7609) <= not b;
    layer5_outputs(7610) <= a;
    layer5_outputs(7611) <= a xor b;
    layer5_outputs(7612) <= not b or a;
    layer5_outputs(7613) <= not a;
    layer5_outputs(7614) <= a or b;
    layer5_outputs(7615) <= not a or b;
    layer5_outputs(7616) <= a;
    layer5_outputs(7617) <= not a;
    layer5_outputs(7618) <= a and not b;
    layer5_outputs(7619) <= b and not a;
    layer5_outputs(7620) <= not (a xor b);
    layer5_outputs(7621) <= a and not b;
    layer5_outputs(7622) <= not a;
    layer5_outputs(7623) <= a or b;
    layer5_outputs(7624) <= not (a and b);
    layer5_outputs(7625) <= b and not a;
    layer5_outputs(7626) <= not b;
    layer5_outputs(7627) <= a and b;
    layer5_outputs(7628) <= a xor b;
    layer5_outputs(7629) <= b and not a;
    layer5_outputs(7630) <= not a or b;
    layer5_outputs(7631) <= not (a and b);
    layer5_outputs(7632) <= a and b;
    layer5_outputs(7633) <= not (a or b);
    layer5_outputs(7634) <= a;
    layer5_outputs(7635) <= not a;
    layer5_outputs(7636) <= not (a or b);
    layer5_outputs(7637) <= not a;
    layer5_outputs(7638) <= a;
    layer5_outputs(7639) <= not b;
    layer5_outputs(7640) <= a and b;
    layer5_outputs(7641) <= not a;
    layer5_outputs(7642) <= b and not a;
    layer5_outputs(7643) <= not a;
    layer5_outputs(7644) <= not b;
    layer5_outputs(7645) <= not (a or b);
    layer5_outputs(7646) <= not a or b;
    layer5_outputs(7647) <= not a;
    layer5_outputs(7648) <= not (a and b);
    layer5_outputs(7649) <= not b or a;
    layer5_outputs(7650) <= not (a and b);
    layer5_outputs(7651) <= a;
    layer5_outputs(7652) <= not (a or b);
    layer5_outputs(7653) <= a;
    layer5_outputs(7654) <= not a;
    layer5_outputs(7655) <= b;
    layer5_outputs(7656) <= not a;
    layer5_outputs(7657) <= a and not b;
    layer5_outputs(7658) <= a or b;
    layer5_outputs(7659) <= not a or b;
    layer5_outputs(7660) <= a;
    layer5_outputs(7661) <= '0';
    layer5_outputs(7662) <= '1';
    layer5_outputs(7663) <= not a;
    layer5_outputs(7664) <= not a or b;
    layer5_outputs(7665) <= not a;
    layer5_outputs(7666) <= not b or a;
    layer5_outputs(7667) <= not (a or b);
    layer5_outputs(7668) <= a xor b;
    layer5_outputs(7669) <= not b or a;
    layer5_outputs(7670) <= not a or b;
    layer5_outputs(7671) <= b;
    layer5_outputs(7672) <= a and b;
    layer5_outputs(7673) <= not b;
    layer5_outputs(7674) <= a or b;
    layer5_outputs(7675) <= b;
    layer5_outputs(7676) <= not b;
    layer5_outputs(7677) <= not b;
    layer5_outputs(7678) <= not (a or b);
    layer5_outputs(7679) <= a;
    layer6_outputs(0) <= a and b;
    layer6_outputs(1) <= b;
    layer6_outputs(2) <= a;
    layer6_outputs(3) <= b;
    layer6_outputs(4) <= not b;
    layer6_outputs(5) <= a and not b;
    layer6_outputs(6) <= not b;
    layer6_outputs(7) <= not b;
    layer6_outputs(8) <= not a;
    layer6_outputs(9) <= not (a and b);
    layer6_outputs(10) <= a and b;
    layer6_outputs(11) <= b;
    layer6_outputs(12) <= not a or b;
    layer6_outputs(13) <= a and not b;
    layer6_outputs(14) <= not b or a;
    layer6_outputs(15) <= not (a or b);
    layer6_outputs(16) <= a;
    layer6_outputs(17) <= not (a or b);
    layer6_outputs(18) <= b;
    layer6_outputs(19) <= b;
    layer6_outputs(20) <= a xor b;
    layer6_outputs(21) <= a and b;
    layer6_outputs(22) <= not b;
    layer6_outputs(23) <= a;
    layer6_outputs(24) <= a;
    layer6_outputs(25) <= a and not b;
    layer6_outputs(26) <= not (a or b);
    layer6_outputs(27) <= a;
    layer6_outputs(28) <= not a or b;
    layer6_outputs(29) <= not a;
    layer6_outputs(30) <= not b;
    layer6_outputs(31) <= a and b;
    layer6_outputs(32) <= not a;
    layer6_outputs(33) <= b;
    layer6_outputs(34) <= b;
    layer6_outputs(35) <= not (a xor b);
    layer6_outputs(36) <= '1';
    layer6_outputs(37) <= b;
    layer6_outputs(38) <= not (a xor b);
    layer6_outputs(39) <= not (a or b);
    layer6_outputs(40) <= a;
    layer6_outputs(41) <= not (a and b);
    layer6_outputs(42) <= a xor b;
    layer6_outputs(43) <= not a;
    layer6_outputs(44) <= not b or a;
    layer6_outputs(45) <= not b;
    layer6_outputs(46) <= not b or a;
    layer6_outputs(47) <= not b or a;
    layer6_outputs(48) <= a and b;
    layer6_outputs(49) <= not (a and b);
    layer6_outputs(50) <= not a;
    layer6_outputs(51) <= not a;
    layer6_outputs(52) <= not (a xor b);
    layer6_outputs(53) <= a and b;
    layer6_outputs(54) <= a or b;
    layer6_outputs(55) <= not a;
    layer6_outputs(56) <= a xor b;
    layer6_outputs(57) <= not a or b;
    layer6_outputs(58) <= not b;
    layer6_outputs(59) <= b and not a;
    layer6_outputs(60) <= a;
    layer6_outputs(61) <= a and not b;
    layer6_outputs(62) <= not (a and b);
    layer6_outputs(63) <= not a;
    layer6_outputs(64) <= not (a xor b);
    layer6_outputs(65) <= a;
    layer6_outputs(66) <= not b;
    layer6_outputs(67) <= '1';
    layer6_outputs(68) <= a or b;
    layer6_outputs(69) <= a and not b;
    layer6_outputs(70) <= '1';
    layer6_outputs(71) <= a and b;
    layer6_outputs(72) <= a;
    layer6_outputs(73) <= b;
    layer6_outputs(74) <= '0';
    layer6_outputs(75) <= not (a and b);
    layer6_outputs(76) <= not (a or b);
    layer6_outputs(77) <= b;
    layer6_outputs(78) <= not (a or b);
    layer6_outputs(79) <= a and b;
    layer6_outputs(80) <= a and not b;
    layer6_outputs(81) <= not b or a;
    layer6_outputs(82) <= not a;
    layer6_outputs(83) <= a;
    layer6_outputs(84) <= b;
    layer6_outputs(85) <= not a;
    layer6_outputs(86) <= b and not a;
    layer6_outputs(87) <= not (a or b);
    layer6_outputs(88) <= b;
    layer6_outputs(89) <= not a;
    layer6_outputs(90) <= not a or b;
    layer6_outputs(91) <= a;
    layer6_outputs(92) <= b and not a;
    layer6_outputs(93) <= not (a or b);
    layer6_outputs(94) <= not a or b;
    layer6_outputs(95) <= b and not a;
    layer6_outputs(96) <= '0';
    layer6_outputs(97) <= not a;
    layer6_outputs(98) <= not a or b;
    layer6_outputs(99) <= not (a xor b);
    layer6_outputs(100) <= not a or b;
    layer6_outputs(101) <= not a;
    layer6_outputs(102) <= not a;
    layer6_outputs(103) <= not a or b;
    layer6_outputs(104) <= a xor b;
    layer6_outputs(105) <= not a or b;
    layer6_outputs(106) <= not a;
    layer6_outputs(107) <= not (a xor b);
    layer6_outputs(108) <= a;
    layer6_outputs(109) <= a and not b;
    layer6_outputs(110) <= b;
    layer6_outputs(111) <= a xor b;
    layer6_outputs(112) <= not a;
    layer6_outputs(113) <= a xor b;
    layer6_outputs(114) <= b;
    layer6_outputs(115) <= not (a xor b);
    layer6_outputs(116) <= b;
    layer6_outputs(117) <= a and b;
    layer6_outputs(118) <= not (a xor b);
    layer6_outputs(119) <= not a or b;
    layer6_outputs(120) <= not (a and b);
    layer6_outputs(121) <= not a;
    layer6_outputs(122) <= a and b;
    layer6_outputs(123) <= not b;
    layer6_outputs(124) <= b and not a;
    layer6_outputs(125) <= '0';
    layer6_outputs(126) <= b;
    layer6_outputs(127) <= not b;
    layer6_outputs(128) <= not b;
    layer6_outputs(129) <= not b;
    layer6_outputs(130) <= not b or a;
    layer6_outputs(131) <= a and b;
    layer6_outputs(132) <= not (a or b);
    layer6_outputs(133) <= b;
    layer6_outputs(134) <= a or b;
    layer6_outputs(135) <= not b or a;
    layer6_outputs(136) <= a or b;
    layer6_outputs(137) <= b and not a;
    layer6_outputs(138) <= not a or b;
    layer6_outputs(139) <= not b;
    layer6_outputs(140) <= a;
    layer6_outputs(141) <= b;
    layer6_outputs(142) <= a;
    layer6_outputs(143) <= not b or a;
    layer6_outputs(144) <= not b;
    layer6_outputs(145) <= a or b;
    layer6_outputs(146) <= a and not b;
    layer6_outputs(147) <= a;
    layer6_outputs(148) <= not a or b;
    layer6_outputs(149) <= not a;
    layer6_outputs(150) <= '0';
    layer6_outputs(151) <= a and b;
    layer6_outputs(152) <= '0';
    layer6_outputs(153) <= not (a or b);
    layer6_outputs(154) <= a and b;
    layer6_outputs(155) <= a or b;
    layer6_outputs(156) <= b;
    layer6_outputs(157) <= not a or b;
    layer6_outputs(158) <= not a;
    layer6_outputs(159) <= not b or a;
    layer6_outputs(160) <= not (a or b);
    layer6_outputs(161) <= not b or a;
    layer6_outputs(162) <= not a;
    layer6_outputs(163) <= b and not a;
    layer6_outputs(164) <= a or b;
    layer6_outputs(165) <= a and b;
    layer6_outputs(166) <= a and not b;
    layer6_outputs(167) <= b and not a;
    layer6_outputs(168) <= not b;
    layer6_outputs(169) <= b;
    layer6_outputs(170) <= b;
    layer6_outputs(171) <= not a;
    layer6_outputs(172) <= a or b;
    layer6_outputs(173) <= not (a xor b);
    layer6_outputs(174) <= not a or b;
    layer6_outputs(175) <= not b or a;
    layer6_outputs(176) <= b;
    layer6_outputs(177) <= not (a xor b);
    layer6_outputs(178) <= not (a xor b);
    layer6_outputs(179) <= '1';
    layer6_outputs(180) <= not a;
    layer6_outputs(181) <= not b;
    layer6_outputs(182) <= '1';
    layer6_outputs(183) <= '1';
    layer6_outputs(184) <= not b;
    layer6_outputs(185) <= not b;
    layer6_outputs(186) <= a and b;
    layer6_outputs(187) <= not (a and b);
    layer6_outputs(188) <= not a;
    layer6_outputs(189) <= not a or b;
    layer6_outputs(190) <= b;
    layer6_outputs(191) <= b and not a;
    layer6_outputs(192) <= a and b;
    layer6_outputs(193) <= a;
    layer6_outputs(194) <= b and not a;
    layer6_outputs(195) <= not b;
    layer6_outputs(196) <= not b;
    layer6_outputs(197) <= a;
    layer6_outputs(198) <= not (a and b);
    layer6_outputs(199) <= not b;
    layer6_outputs(200) <= b;
    layer6_outputs(201) <= b;
    layer6_outputs(202) <= '1';
    layer6_outputs(203) <= not b;
    layer6_outputs(204) <= b;
    layer6_outputs(205) <= not (a or b);
    layer6_outputs(206) <= '0';
    layer6_outputs(207) <= not (a or b);
    layer6_outputs(208) <= a and b;
    layer6_outputs(209) <= b;
    layer6_outputs(210) <= not a;
    layer6_outputs(211) <= not (a or b);
    layer6_outputs(212) <= a and b;
    layer6_outputs(213) <= a and not b;
    layer6_outputs(214) <= a;
    layer6_outputs(215) <= not (a or b);
    layer6_outputs(216) <= a;
    layer6_outputs(217) <= not b or a;
    layer6_outputs(218) <= not a;
    layer6_outputs(219) <= '1';
    layer6_outputs(220) <= not b;
    layer6_outputs(221) <= a;
    layer6_outputs(222) <= not (a and b);
    layer6_outputs(223) <= a and b;
    layer6_outputs(224) <= not b;
    layer6_outputs(225) <= not b;
    layer6_outputs(226) <= a xor b;
    layer6_outputs(227) <= a and not b;
    layer6_outputs(228) <= not (a xor b);
    layer6_outputs(229) <= a;
    layer6_outputs(230) <= b;
    layer6_outputs(231) <= b;
    layer6_outputs(232) <= a and not b;
    layer6_outputs(233) <= not b or a;
    layer6_outputs(234) <= not (a xor b);
    layer6_outputs(235) <= '0';
    layer6_outputs(236) <= not a;
    layer6_outputs(237) <= not (a or b);
    layer6_outputs(238) <= a xor b;
    layer6_outputs(239) <= b and not a;
    layer6_outputs(240) <= not (a or b);
    layer6_outputs(241) <= '0';
    layer6_outputs(242) <= not (a and b);
    layer6_outputs(243) <= not (a xor b);
    layer6_outputs(244) <= not a;
    layer6_outputs(245) <= a and b;
    layer6_outputs(246) <= b and not a;
    layer6_outputs(247) <= a;
    layer6_outputs(248) <= not (a xor b);
    layer6_outputs(249) <= b;
    layer6_outputs(250) <= '0';
    layer6_outputs(251) <= a;
    layer6_outputs(252) <= not a;
    layer6_outputs(253) <= not (a xor b);
    layer6_outputs(254) <= not a;
    layer6_outputs(255) <= not b;
    layer6_outputs(256) <= b;
    layer6_outputs(257) <= a and not b;
    layer6_outputs(258) <= not b;
    layer6_outputs(259) <= not (a or b);
    layer6_outputs(260) <= a;
    layer6_outputs(261) <= b;
    layer6_outputs(262) <= b;
    layer6_outputs(263) <= not b;
    layer6_outputs(264) <= not a;
    layer6_outputs(265) <= a;
    layer6_outputs(266) <= a xor b;
    layer6_outputs(267) <= not (a and b);
    layer6_outputs(268) <= a;
    layer6_outputs(269) <= b;
    layer6_outputs(270) <= not a;
    layer6_outputs(271) <= not a;
    layer6_outputs(272) <= a;
    layer6_outputs(273) <= a or b;
    layer6_outputs(274) <= a and b;
    layer6_outputs(275) <= a;
    layer6_outputs(276) <= a and not b;
    layer6_outputs(277) <= not (a and b);
    layer6_outputs(278) <= not (a xor b);
    layer6_outputs(279) <= '1';
    layer6_outputs(280) <= not (a or b);
    layer6_outputs(281) <= b;
    layer6_outputs(282) <= not b or a;
    layer6_outputs(283) <= not (a or b);
    layer6_outputs(284) <= not a or b;
    layer6_outputs(285) <= a or b;
    layer6_outputs(286) <= not a;
    layer6_outputs(287) <= a and b;
    layer6_outputs(288) <= not b;
    layer6_outputs(289) <= not (a and b);
    layer6_outputs(290) <= not a;
    layer6_outputs(291) <= b;
    layer6_outputs(292) <= not a;
    layer6_outputs(293) <= a;
    layer6_outputs(294) <= not b;
    layer6_outputs(295) <= a or b;
    layer6_outputs(296) <= not b;
    layer6_outputs(297) <= not (a and b);
    layer6_outputs(298) <= not (a or b);
    layer6_outputs(299) <= a;
    layer6_outputs(300) <= a xor b;
    layer6_outputs(301) <= not a or b;
    layer6_outputs(302) <= not a or b;
    layer6_outputs(303) <= not (a and b);
    layer6_outputs(304) <= a;
    layer6_outputs(305) <= not b;
    layer6_outputs(306) <= a and b;
    layer6_outputs(307) <= a and b;
    layer6_outputs(308) <= not a;
    layer6_outputs(309) <= a;
    layer6_outputs(310) <= not b or a;
    layer6_outputs(311) <= a and b;
    layer6_outputs(312) <= not (a and b);
    layer6_outputs(313) <= not a or b;
    layer6_outputs(314) <= not (a xor b);
    layer6_outputs(315) <= '1';
    layer6_outputs(316) <= a xor b;
    layer6_outputs(317) <= b;
    layer6_outputs(318) <= a or b;
    layer6_outputs(319) <= not (a or b);
    layer6_outputs(320) <= a;
    layer6_outputs(321) <= not a;
    layer6_outputs(322) <= a;
    layer6_outputs(323) <= not b;
    layer6_outputs(324) <= not b;
    layer6_outputs(325) <= a xor b;
    layer6_outputs(326) <= not b;
    layer6_outputs(327) <= not (a and b);
    layer6_outputs(328) <= not b;
    layer6_outputs(329) <= a and b;
    layer6_outputs(330) <= not a;
    layer6_outputs(331) <= not b or a;
    layer6_outputs(332) <= not b or a;
    layer6_outputs(333) <= not (a or b);
    layer6_outputs(334) <= b and not a;
    layer6_outputs(335) <= b;
    layer6_outputs(336) <= not a or b;
    layer6_outputs(337) <= '0';
    layer6_outputs(338) <= not a or b;
    layer6_outputs(339) <= not a;
    layer6_outputs(340) <= not (a xor b);
    layer6_outputs(341) <= a and not b;
    layer6_outputs(342) <= b;
    layer6_outputs(343) <= b;
    layer6_outputs(344) <= not b;
    layer6_outputs(345) <= not a;
    layer6_outputs(346) <= a and not b;
    layer6_outputs(347) <= a;
    layer6_outputs(348) <= b and not a;
    layer6_outputs(349) <= not a;
    layer6_outputs(350) <= a and not b;
    layer6_outputs(351) <= a;
    layer6_outputs(352) <= not a;
    layer6_outputs(353) <= a or b;
    layer6_outputs(354) <= b and not a;
    layer6_outputs(355) <= '1';
    layer6_outputs(356) <= '0';
    layer6_outputs(357) <= not a;
    layer6_outputs(358) <= b;
    layer6_outputs(359) <= not a;
    layer6_outputs(360) <= a and not b;
    layer6_outputs(361) <= not (a or b);
    layer6_outputs(362) <= a;
    layer6_outputs(363) <= '0';
    layer6_outputs(364) <= not b;
    layer6_outputs(365) <= not (a or b);
    layer6_outputs(366) <= a and not b;
    layer6_outputs(367) <= b and not a;
    layer6_outputs(368) <= not b or a;
    layer6_outputs(369) <= not b;
    layer6_outputs(370) <= a and not b;
    layer6_outputs(371) <= not (a and b);
    layer6_outputs(372) <= b;
    layer6_outputs(373) <= not (a and b);
    layer6_outputs(374) <= b;
    layer6_outputs(375) <= not a;
    layer6_outputs(376) <= not b;
    layer6_outputs(377) <= not (a or b);
    layer6_outputs(378) <= a;
    layer6_outputs(379) <= not b or a;
    layer6_outputs(380) <= not a or b;
    layer6_outputs(381) <= a;
    layer6_outputs(382) <= a;
    layer6_outputs(383) <= a or b;
    layer6_outputs(384) <= a or b;
    layer6_outputs(385) <= b;
    layer6_outputs(386) <= a and not b;
    layer6_outputs(387) <= not b or a;
    layer6_outputs(388) <= not (a or b);
    layer6_outputs(389) <= not b or a;
    layer6_outputs(390) <= not (a xor b);
    layer6_outputs(391) <= b;
    layer6_outputs(392) <= b and not a;
    layer6_outputs(393) <= not (a xor b);
    layer6_outputs(394) <= b;
    layer6_outputs(395) <= a or b;
    layer6_outputs(396) <= a or b;
    layer6_outputs(397) <= not a;
    layer6_outputs(398) <= not a;
    layer6_outputs(399) <= b and not a;
    layer6_outputs(400) <= not b;
    layer6_outputs(401) <= not a or b;
    layer6_outputs(402) <= not b or a;
    layer6_outputs(403) <= a xor b;
    layer6_outputs(404) <= '1';
    layer6_outputs(405) <= not b or a;
    layer6_outputs(406) <= not a;
    layer6_outputs(407) <= not (a or b);
    layer6_outputs(408) <= not (a xor b);
    layer6_outputs(409) <= b;
    layer6_outputs(410) <= a xor b;
    layer6_outputs(411) <= a and b;
    layer6_outputs(412) <= '1';
    layer6_outputs(413) <= not b or a;
    layer6_outputs(414) <= a or b;
    layer6_outputs(415) <= a and b;
    layer6_outputs(416) <= a and not b;
    layer6_outputs(417) <= not b;
    layer6_outputs(418) <= not (a and b);
    layer6_outputs(419) <= a and not b;
    layer6_outputs(420) <= not b;
    layer6_outputs(421) <= a;
    layer6_outputs(422) <= a;
    layer6_outputs(423) <= not (a xor b);
    layer6_outputs(424) <= a and b;
    layer6_outputs(425) <= b;
    layer6_outputs(426) <= not a;
    layer6_outputs(427) <= b and not a;
    layer6_outputs(428) <= not a;
    layer6_outputs(429) <= a xor b;
    layer6_outputs(430) <= b and not a;
    layer6_outputs(431) <= b;
    layer6_outputs(432) <= '0';
    layer6_outputs(433) <= not a;
    layer6_outputs(434) <= b;
    layer6_outputs(435) <= not b;
    layer6_outputs(436) <= b and not a;
    layer6_outputs(437) <= a and b;
    layer6_outputs(438) <= not (a and b);
    layer6_outputs(439) <= a or b;
    layer6_outputs(440) <= '0';
    layer6_outputs(441) <= not a or b;
    layer6_outputs(442) <= b;
    layer6_outputs(443) <= b;
    layer6_outputs(444) <= a and not b;
    layer6_outputs(445) <= not (a and b);
    layer6_outputs(446) <= b;
    layer6_outputs(447) <= not a;
    layer6_outputs(448) <= not a;
    layer6_outputs(449) <= not (a and b);
    layer6_outputs(450) <= a and b;
    layer6_outputs(451) <= b;
    layer6_outputs(452) <= a;
    layer6_outputs(453) <= not a;
    layer6_outputs(454) <= not (a or b);
    layer6_outputs(455) <= '0';
    layer6_outputs(456) <= not a;
    layer6_outputs(457) <= not a;
    layer6_outputs(458) <= not a or b;
    layer6_outputs(459) <= a or b;
    layer6_outputs(460) <= a xor b;
    layer6_outputs(461) <= a;
    layer6_outputs(462) <= a;
    layer6_outputs(463) <= not (a or b);
    layer6_outputs(464) <= not b or a;
    layer6_outputs(465) <= a;
    layer6_outputs(466) <= a and not b;
    layer6_outputs(467) <= not (a or b);
    layer6_outputs(468) <= b;
    layer6_outputs(469) <= not b or a;
    layer6_outputs(470) <= a and not b;
    layer6_outputs(471) <= a or b;
    layer6_outputs(472) <= not b or a;
    layer6_outputs(473) <= a;
    layer6_outputs(474) <= a xor b;
    layer6_outputs(475) <= not a;
    layer6_outputs(476) <= a xor b;
    layer6_outputs(477) <= b;
    layer6_outputs(478) <= a;
    layer6_outputs(479) <= not (a or b);
    layer6_outputs(480) <= not (a or b);
    layer6_outputs(481) <= b;
    layer6_outputs(482) <= b and not a;
    layer6_outputs(483) <= not b;
    layer6_outputs(484) <= a and b;
    layer6_outputs(485) <= a and b;
    layer6_outputs(486) <= b;
    layer6_outputs(487) <= not b or a;
    layer6_outputs(488) <= not b;
    layer6_outputs(489) <= '0';
    layer6_outputs(490) <= a;
    layer6_outputs(491) <= not a or b;
    layer6_outputs(492) <= b;
    layer6_outputs(493) <= b;
    layer6_outputs(494) <= a and not b;
    layer6_outputs(495) <= a or b;
    layer6_outputs(496) <= b;
    layer6_outputs(497) <= a and not b;
    layer6_outputs(498) <= not b or a;
    layer6_outputs(499) <= a;
    layer6_outputs(500) <= a;
    layer6_outputs(501) <= b;
    layer6_outputs(502) <= b;
    layer6_outputs(503) <= not a;
    layer6_outputs(504) <= a and not b;
    layer6_outputs(505) <= a and b;
    layer6_outputs(506) <= a and not b;
    layer6_outputs(507) <= not (a or b);
    layer6_outputs(508) <= a xor b;
    layer6_outputs(509) <= not a;
    layer6_outputs(510) <= not b;
    layer6_outputs(511) <= b;
    layer6_outputs(512) <= a;
    layer6_outputs(513) <= b and not a;
    layer6_outputs(514) <= not b;
    layer6_outputs(515) <= not a;
    layer6_outputs(516) <= '1';
    layer6_outputs(517) <= not (a or b);
    layer6_outputs(518) <= b;
    layer6_outputs(519) <= not a;
    layer6_outputs(520) <= a or b;
    layer6_outputs(521) <= a xor b;
    layer6_outputs(522) <= a xor b;
    layer6_outputs(523) <= not (a and b);
    layer6_outputs(524) <= a;
    layer6_outputs(525) <= a xor b;
    layer6_outputs(526) <= a;
    layer6_outputs(527) <= not (a and b);
    layer6_outputs(528) <= a or b;
    layer6_outputs(529) <= not a;
    layer6_outputs(530) <= not (a xor b);
    layer6_outputs(531) <= not a or b;
    layer6_outputs(532) <= not (a xor b);
    layer6_outputs(533) <= not b;
    layer6_outputs(534) <= a or b;
    layer6_outputs(535) <= not a;
    layer6_outputs(536) <= b;
    layer6_outputs(537) <= b;
    layer6_outputs(538) <= not b or a;
    layer6_outputs(539) <= not (a xor b);
    layer6_outputs(540) <= not b;
    layer6_outputs(541) <= a and not b;
    layer6_outputs(542) <= not (a xor b);
    layer6_outputs(543) <= not a;
    layer6_outputs(544) <= not a or b;
    layer6_outputs(545) <= a;
    layer6_outputs(546) <= '0';
    layer6_outputs(547) <= not b or a;
    layer6_outputs(548) <= b;
    layer6_outputs(549) <= a xor b;
    layer6_outputs(550) <= not b;
    layer6_outputs(551) <= not (a xor b);
    layer6_outputs(552) <= a and b;
    layer6_outputs(553) <= not a or b;
    layer6_outputs(554) <= b;
    layer6_outputs(555) <= not (a and b);
    layer6_outputs(556) <= not b;
    layer6_outputs(557) <= a or b;
    layer6_outputs(558) <= not (a xor b);
    layer6_outputs(559) <= not (a and b);
    layer6_outputs(560) <= a xor b;
    layer6_outputs(561) <= a or b;
    layer6_outputs(562) <= not (a and b);
    layer6_outputs(563) <= not (a or b);
    layer6_outputs(564) <= b and not a;
    layer6_outputs(565) <= not b;
    layer6_outputs(566) <= not (a xor b);
    layer6_outputs(567) <= a and b;
    layer6_outputs(568) <= b;
    layer6_outputs(569) <= not a;
    layer6_outputs(570) <= '0';
    layer6_outputs(571) <= not a;
    layer6_outputs(572) <= not a or b;
    layer6_outputs(573) <= not (a and b);
    layer6_outputs(574) <= not a or b;
    layer6_outputs(575) <= a and b;
    layer6_outputs(576) <= not a or b;
    layer6_outputs(577) <= not (a or b);
    layer6_outputs(578) <= '0';
    layer6_outputs(579) <= not b;
    layer6_outputs(580) <= not (a and b);
    layer6_outputs(581) <= '1';
    layer6_outputs(582) <= not a or b;
    layer6_outputs(583) <= a;
    layer6_outputs(584) <= not a;
    layer6_outputs(585) <= a;
    layer6_outputs(586) <= not b or a;
    layer6_outputs(587) <= not (a xor b);
    layer6_outputs(588) <= a;
    layer6_outputs(589) <= b;
    layer6_outputs(590) <= b and not a;
    layer6_outputs(591) <= b and not a;
    layer6_outputs(592) <= a and b;
    layer6_outputs(593) <= not (a and b);
    layer6_outputs(594) <= a and not b;
    layer6_outputs(595) <= not a;
    layer6_outputs(596) <= not a;
    layer6_outputs(597) <= '1';
    layer6_outputs(598) <= '0';
    layer6_outputs(599) <= not a or b;
    layer6_outputs(600) <= b;
    layer6_outputs(601) <= not (a xor b);
    layer6_outputs(602) <= not b;
    layer6_outputs(603) <= not b or a;
    layer6_outputs(604) <= a xor b;
    layer6_outputs(605) <= b and not a;
    layer6_outputs(606) <= not b;
    layer6_outputs(607) <= not (a and b);
    layer6_outputs(608) <= not b;
    layer6_outputs(609) <= b and not a;
    layer6_outputs(610) <= not b or a;
    layer6_outputs(611) <= '0';
    layer6_outputs(612) <= not b;
    layer6_outputs(613) <= a;
    layer6_outputs(614) <= not a;
    layer6_outputs(615) <= not b or a;
    layer6_outputs(616) <= not a or b;
    layer6_outputs(617) <= not a;
    layer6_outputs(618) <= not a or b;
    layer6_outputs(619) <= b;
    layer6_outputs(620) <= a or b;
    layer6_outputs(621) <= not (a or b);
    layer6_outputs(622) <= '0';
    layer6_outputs(623) <= a;
    layer6_outputs(624) <= not a;
    layer6_outputs(625) <= not (a and b);
    layer6_outputs(626) <= b and not a;
    layer6_outputs(627) <= b;
    layer6_outputs(628) <= b;
    layer6_outputs(629) <= a;
    layer6_outputs(630) <= not (a and b);
    layer6_outputs(631) <= b;
    layer6_outputs(632) <= a and not b;
    layer6_outputs(633) <= a or b;
    layer6_outputs(634) <= a;
    layer6_outputs(635) <= a;
    layer6_outputs(636) <= a or b;
    layer6_outputs(637) <= a;
    layer6_outputs(638) <= a and b;
    layer6_outputs(639) <= a and b;
    layer6_outputs(640) <= not a;
    layer6_outputs(641) <= not a;
    layer6_outputs(642) <= '1';
    layer6_outputs(643) <= not a;
    layer6_outputs(644) <= b;
    layer6_outputs(645) <= not (a and b);
    layer6_outputs(646) <= not (a or b);
    layer6_outputs(647) <= a or b;
    layer6_outputs(648) <= a and b;
    layer6_outputs(649) <= b;
    layer6_outputs(650) <= '0';
    layer6_outputs(651) <= '0';
    layer6_outputs(652) <= b and not a;
    layer6_outputs(653) <= a;
    layer6_outputs(654) <= not b;
    layer6_outputs(655) <= b and not a;
    layer6_outputs(656) <= a;
    layer6_outputs(657) <= not b or a;
    layer6_outputs(658) <= b;
    layer6_outputs(659) <= not a or b;
    layer6_outputs(660) <= not b or a;
    layer6_outputs(661) <= a or b;
    layer6_outputs(662) <= not a;
    layer6_outputs(663) <= not b;
    layer6_outputs(664) <= a or b;
    layer6_outputs(665) <= a;
    layer6_outputs(666) <= '1';
    layer6_outputs(667) <= '1';
    layer6_outputs(668) <= not a or b;
    layer6_outputs(669) <= not a or b;
    layer6_outputs(670) <= not (a or b);
    layer6_outputs(671) <= not (a xor b);
    layer6_outputs(672) <= not a;
    layer6_outputs(673) <= not b or a;
    layer6_outputs(674) <= not (a xor b);
    layer6_outputs(675) <= b and not a;
    layer6_outputs(676) <= not a;
    layer6_outputs(677) <= not a;
    layer6_outputs(678) <= not a or b;
    layer6_outputs(679) <= a and not b;
    layer6_outputs(680) <= not (a and b);
    layer6_outputs(681) <= a;
    layer6_outputs(682) <= not b or a;
    layer6_outputs(683) <= '1';
    layer6_outputs(684) <= a or b;
    layer6_outputs(685) <= not (a or b);
    layer6_outputs(686) <= a;
    layer6_outputs(687) <= not (a xor b);
    layer6_outputs(688) <= not (a or b);
    layer6_outputs(689) <= a and not b;
    layer6_outputs(690) <= b and not a;
    layer6_outputs(691) <= not (a and b);
    layer6_outputs(692) <= not (a or b);
    layer6_outputs(693) <= b;
    layer6_outputs(694) <= not b or a;
    layer6_outputs(695) <= not b;
    layer6_outputs(696) <= b and not a;
    layer6_outputs(697) <= b and not a;
    layer6_outputs(698) <= not (a and b);
    layer6_outputs(699) <= b;
    layer6_outputs(700) <= '0';
    layer6_outputs(701) <= not (a and b);
    layer6_outputs(702) <= not b;
    layer6_outputs(703) <= '1';
    layer6_outputs(704) <= b;
    layer6_outputs(705) <= a;
    layer6_outputs(706) <= not (a xor b);
    layer6_outputs(707) <= b;
    layer6_outputs(708) <= not (a and b);
    layer6_outputs(709) <= not a;
    layer6_outputs(710) <= b;
    layer6_outputs(711) <= b;
    layer6_outputs(712) <= a;
    layer6_outputs(713) <= a or b;
    layer6_outputs(714) <= b;
    layer6_outputs(715) <= a;
    layer6_outputs(716) <= a and not b;
    layer6_outputs(717) <= not b;
    layer6_outputs(718) <= not b or a;
    layer6_outputs(719) <= not b or a;
    layer6_outputs(720) <= not a;
    layer6_outputs(721) <= b;
    layer6_outputs(722) <= not (a or b);
    layer6_outputs(723) <= a;
    layer6_outputs(724) <= a;
    layer6_outputs(725) <= b;
    layer6_outputs(726) <= not b;
    layer6_outputs(727) <= a and b;
    layer6_outputs(728) <= b;
    layer6_outputs(729) <= a xor b;
    layer6_outputs(730) <= b;
    layer6_outputs(731) <= not (a xor b);
    layer6_outputs(732) <= b and not a;
    layer6_outputs(733) <= b and not a;
    layer6_outputs(734) <= not b or a;
    layer6_outputs(735) <= a;
    layer6_outputs(736) <= b and not a;
    layer6_outputs(737) <= not (a and b);
    layer6_outputs(738) <= not a;
    layer6_outputs(739) <= not (a or b);
    layer6_outputs(740) <= not b;
    layer6_outputs(741) <= a or b;
    layer6_outputs(742) <= not a or b;
    layer6_outputs(743) <= not (a and b);
    layer6_outputs(744) <= b;
    layer6_outputs(745) <= a;
    layer6_outputs(746) <= a and not b;
    layer6_outputs(747) <= not a;
    layer6_outputs(748) <= a or b;
    layer6_outputs(749) <= not a;
    layer6_outputs(750) <= not a;
    layer6_outputs(751) <= not b or a;
    layer6_outputs(752) <= not (a xor b);
    layer6_outputs(753) <= not a;
    layer6_outputs(754) <= not (a xor b);
    layer6_outputs(755) <= a and not b;
    layer6_outputs(756) <= not b or a;
    layer6_outputs(757) <= b;
    layer6_outputs(758) <= a;
    layer6_outputs(759) <= not (a and b);
    layer6_outputs(760) <= not a;
    layer6_outputs(761) <= a or b;
    layer6_outputs(762) <= '0';
    layer6_outputs(763) <= not b or a;
    layer6_outputs(764) <= not a;
    layer6_outputs(765) <= not b;
    layer6_outputs(766) <= a;
    layer6_outputs(767) <= a;
    layer6_outputs(768) <= a and b;
    layer6_outputs(769) <= not b;
    layer6_outputs(770) <= a or b;
    layer6_outputs(771) <= not b;
    layer6_outputs(772) <= a or b;
    layer6_outputs(773) <= not a or b;
    layer6_outputs(774) <= a or b;
    layer6_outputs(775) <= b and not a;
    layer6_outputs(776) <= not a or b;
    layer6_outputs(777) <= not (a and b);
    layer6_outputs(778) <= a or b;
    layer6_outputs(779) <= a xor b;
    layer6_outputs(780) <= a;
    layer6_outputs(781) <= a and not b;
    layer6_outputs(782) <= not a;
    layer6_outputs(783) <= a and b;
    layer6_outputs(784) <= a;
    layer6_outputs(785) <= not a or b;
    layer6_outputs(786) <= '1';
    layer6_outputs(787) <= a and not b;
    layer6_outputs(788) <= a;
    layer6_outputs(789) <= a and not b;
    layer6_outputs(790) <= a xor b;
    layer6_outputs(791) <= not (a or b);
    layer6_outputs(792) <= a xor b;
    layer6_outputs(793) <= not b;
    layer6_outputs(794) <= b and not a;
    layer6_outputs(795) <= '0';
    layer6_outputs(796) <= b;
    layer6_outputs(797) <= b;
    layer6_outputs(798) <= a or b;
    layer6_outputs(799) <= '0';
    layer6_outputs(800) <= not (a xor b);
    layer6_outputs(801) <= not a;
    layer6_outputs(802) <= a and not b;
    layer6_outputs(803) <= '0';
    layer6_outputs(804) <= '1';
    layer6_outputs(805) <= a or b;
    layer6_outputs(806) <= '0';
    layer6_outputs(807) <= not b or a;
    layer6_outputs(808) <= not (a xor b);
    layer6_outputs(809) <= not (a or b);
    layer6_outputs(810) <= not (a xor b);
    layer6_outputs(811) <= a and b;
    layer6_outputs(812) <= not (a xor b);
    layer6_outputs(813) <= not (a or b);
    layer6_outputs(814) <= b and not a;
    layer6_outputs(815) <= a and b;
    layer6_outputs(816) <= not a or b;
    layer6_outputs(817) <= a and not b;
    layer6_outputs(818) <= '1';
    layer6_outputs(819) <= b;
    layer6_outputs(820) <= '1';
    layer6_outputs(821) <= not a;
    layer6_outputs(822) <= not b or a;
    layer6_outputs(823) <= '1';
    layer6_outputs(824) <= b;
    layer6_outputs(825) <= not a;
    layer6_outputs(826) <= a or b;
    layer6_outputs(827) <= b and not a;
    layer6_outputs(828) <= a and not b;
    layer6_outputs(829) <= not a or b;
    layer6_outputs(830) <= not (a and b);
    layer6_outputs(831) <= a;
    layer6_outputs(832) <= b;
    layer6_outputs(833) <= not b or a;
    layer6_outputs(834) <= not a;
    layer6_outputs(835) <= not b or a;
    layer6_outputs(836) <= not a;
    layer6_outputs(837) <= b;
    layer6_outputs(838) <= a and not b;
    layer6_outputs(839) <= b and not a;
    layer6_outputs(840) <= not (a and b);
    layer6_outputs(841) <= not b;
    layer6_outputs(842) <= not a;
    layer6_outputs(843) <= not a;
    layer6_outputs(844) <= a;
    layer6_outputs(845) <= b;
    layer6_outputs(846) <= not a or b;
    layer6_outputs(847) <= b;
    layer6_outputs(848) <= b;
    layer6_outputs(849) <= not b;
    layer6_outputs(850) <= a xor b;
    layer6_outputs(851) <= not b;
    layer6_outputs(852) <= not (a xor b);
    layer6_outputs(853) <= a and not b;
    layer6_outputs(854) <= a and not b;
    layer6_outputs(855) <= a;
    layer6_outputs(856) <= not b or a;
    layer6_outputs(857) <= not b;
    layer6_outputs(858) <= a xor b;
    layer6_outputs(859) <= a and not b;
    layer6_outputs(860) <= not b;
    layer6_outputs(861) <= a or b;
    layer6_outputs(862) <= not (a and b);
    layer6_outputs(863) <= not b or a;
    layer6_outputs(864) <= a;
    layer6_outputs(865) <= not b;
    layer6_outputs(866) <= not (a and b);
    layer6_outputs(867) <= a or b;
    layer6_outputs(868) <= b and not a;
    layer6_outputs(869) <= not (a xor b);
    layer6_outputs(870) <= not (a xor b);
    layer6_outputs(871) <= a xor b;
    layer6_outputs(872) <= a and b;
    layer6_outputs(873) <= a;
    layer6_outputs(874) <= not b;
    layer6_outputs(875) <= a;
    layer6_outputs(876) <= '1';
    layer6_outputs(877) <= not b;
    layer6_outputs(878) <= not a;
    layer6_outputs(879) <= a and not b;
    layer6_outputs(880) <= b;
    layer6_outputs(881) <= a;
    layer6_outputs(882) <= a and not b;
    layer6_outputs(883) <= '0';
    layer6_outputs(884) <= b;
    layer6_outputs(885) <= not b or a;
    layer6_outputs(886) <= '1';
    layer6_outputs(887) <= a;
    layer6_outputs(888) <= not b or a;
    layer6_outputs(889) <= a;
    layer6_outputs(890) <= not b;
    layer6_outputs(891) <= a;
    layer6_outputs(892) <= a;
    layer6_outputs(893) <= not a;
    layer6_outputs(894) <= not a;
    layer6_outputs(895) <= a or b;
    layer6_outputs(896) <= not b;
    layer6_outputs(897) <= not a;
    layer6_outputs(898) <= b;
    layer6_outputs(899) <= a;
    layer6_outputs(900) <= a;
    layer6_outputs(901) <= b;
    layer6_outputs(902) <= b;
    layer6_outputs(903) <= a xor b;
    layer6_outputs(904) <= not (a xor b);
    layer6_outputs(905) <= a;
    layer6_outputs(906) <= not a or b;
    layer6_outputs(907) <= not (a xor b);
    layer6_outputs(908) <= not a;
    layer6_outputs(909) <= b;
    layer6_outputs(910) <= not b;
    layer6_outputs(911) <= not a or b;
    layer6_outputs(912) <= b;
    layer6_outputs(913) <= '0';
    layer6_outputs(914) <= a or b;
    layer6_outputs(915) <= not (a xor b);
    layer6_outputs(916) <= not (a and b);
    layer6_outputs(917) <= b;
    layer6_outputs(918) <= a and b;
    layer6_outputs(919) <= b and not a;
    layer6_outputs(920) <= not a;
    layer6_outputs(921) <= not (a or b);
    layer6_outputs(922) <= a xor b;
    layer6_outputs(923) <= a;
    layer6_outputs(924) <= a;
    layer6_outputs(925) <= not b;
    layer6_outputs(926) <= a and not b;
    layer6_outputs(927) <= a;
    layer6_outputs(928) <= a and not b;
    layer6_outputs(929) <= a and b;
    layer6_outputs(930) <= not b or a;
    layer6_outputs(931) <= not a;
    layer6_outputs(932) <= b and not a;
    layer6_outputs(933) <= not a;
    layer6_outputs(934) <= a or b;
    layer6_outputs(935) <= b;
    layer6_outputs(936) <= not a or b;
    layer6_outputs(937) <= a or b;
    layer6_outputs(938) <= not b or a;
    layer6_outputs(939) <= not a;
    layer6_outputs(940) <= '0';
    layer6_outputs(941) <= a;
    layer6_outputs(942) <= not b;
    layer6_outputs(943) <= '0';
    layer6_outputs(944) <= a;
    layer6_outputs(945) <= not a;
    layer6_outputs(946) <= not a or b;
    layer6_outputs(947) <= not b;
    layer6_outputs(948) <= a and b;
    layer6_outputs(949) <= not a;
    layer6_outputs(950) <= not b;
    layer6_outputs(951) <= not (a or b);
    layer6_outputs(952) <= b;
    layer6_outputs(953) <= not (a or b);
    layer6_outputs(954) <= not (a xor b);
    layer6_outputs(955) <= a;
    layer6_outputs(956) <= not a;
    layer6_outputs(957) <= b and not a;
    layer6_outputs(958) <= not (a and b);
    layer6_outputs(959) <= a and b;
    layer6_outputs(960) <= b;
    layer6_outputs(961) <= not a or b;
    layer6_outputs(962) <= a or b;
    layer6_outputs(963) <= b;
    layer6_outputs(964) <= '1';
    layer6_outputs(965) <= a;
    layer6_outputs(966) <= a or b;
    layer6_outputs(967) <= b;
    layer6_outputs(968) <= a xor b;
    layer6_outputs(969) <= not a;
    layer6_outputs(970) <= not (a xor b);
    layer6_outputs(971) <= not a or b;
    layer6_outputs(972) <= a and b;
    layer6_outputs(973) <= '1';
    layer6_outputs(974) <= b and not a;
    layer6_outputs(975) <= a and b;
    layer6_outputs(976) <= not b;
    layer6_outputs(977) <= not (a or b);
    layer6_outputs(978) <= not a or b;
    layer6_outputs(979) <= not a or b;
    layer6_outputs(980) <= a and b;
    layer6_outputs(981) <= not a;
    layer6_outputs(982) <= b;
    layer6_outputs(983) <= not (a xor b);
    layer6_outputs(984) <= not a;
    layer6_outputs(985) <= b;
    layer6_outputs(986) <= a or b;
    layer6_outputs(987) <= b;
    layer6_outputs(988) <= a and not b;
    layer6_outputs(989) <= not b;
    layer6_outputs(990) <= not a;
    layer6_outputs(991) <= '1';
    layer6_outputs(992) <= a;
    layer6_outputs(993) <= a and not b;
    layer6_outputs(994) <= not a;
    layer6_outputs(995) <= '0';
    layer6_outputs(996) <= a and b;
    layer6_outputs(997) <= b and not a;
    layer6_outputs(998) <= '0';
    layer6_outputs(999) <= not (a xor b);
    layer6_outputs(1000) <= a or b;
    layer6_outputs(1001) <= not a or b;
    layer6_outputs(1002) <= not a or b;
    layer6_outputs(1003) <= not b or a;
    layer6_outputs(1004) <= a and b;
    layer6_outputs(1005) <= '1';
    layer6_outputs(1006) <= not (a xor b);
    layer6_outputs(1007) <= not a;
    layer6_outputs(1008) <= '0';
    layer6_outputs(1009) <= not a;
    layer6_outputs(1010) <= not b;
    layer6_outputs(1011) <= b;
    layer6_outputs(1012) <= '0';
    layer6_outputs(1013) <= b and not a;
    layer6_outputs(1014) <= not (a xor b);
    layer6_outputs(1015) <= a or b;
    layer6_outputs(1016) <= not (a or b);
    layer6_outputs(1017) <= a or b;
    layer6_outputs(1018) <= b;
    layer6_outputs(1019) <= not (a or b);
    layer6_outputs(1020) <= not a;
    layer6_outputs(1021) <= not b;
    layer6_outputs(1022) <= a or b;
    layer6_outputs(1023) <= '0';
    layer6_outputs(1024) <= not b;
    layer6_outputs(1025) <= b;
    layer6_outputs(1026) <= not b or a;
    layer6_outputs(1027) <= not a or b;
    layer6_outputs(1028) <= not b or a;
    layer6_outputs(1029) <= not a or b;
    layer6_outputs(1030) <= b;
    layer6_outputs(1031) <= a or b;
    layer6_outputs(1032) <= not b;
    layer6_outputs(1033) <= not b;
    layer6_outputs(1034) <= not b;
    layer6_outputs(1035) <= not (a or b);
    layer6_outputs(1036) <= not (a xor b);
    layer6_outputs(1037) <= not b;
    layer6_outputs(1038) <= not b;
    layer6_outputs(1039) <= a and not b;
    layer6_outputs(1040) <= b;
    layer6_outputs(1041) <= '0';
    layer6_outputs(1042) <= not (a xor b);
    layer6_outputs(1043) <= '1';
    layer6_outputs(1044) <= not a;
    layer6_outputs(1045) <= a;
    layer6_outputs(1046) <= a xor b;
    layer6_outputs(1047) <= a or b;
    layer6_outputs(1048) <= not (a xor b);
    layer6_outputs(1049) <= a;
    layer6_outputs(1050) <= b;
    layer6_outputs(1051) <= not a;
    layer6_outputs(1052) <= a;
    layer6_outputs(1053) <= not (a or b);
    layer6_outputs(1054) <= a;
    layer6_outputs(1055) <= not (a and b);
    layer6_outputs(1056) <= not (a or b);
    layer6_outputs(1057) <= a and b;
    layer6_outputs(1058) <= '0';
    layer6_outputs(1059) <= '0';
    layer6_outputs(1060) <= b;
    layer6_outputs(1061) <= not a;
    layer6_outputs(1062) <= a;
    layer6_outputs(1063) <= not (a or b);
    layer6_outputs(1064) <= b and not a;
    layer6_outputs(1065) <= not (a or b);
    layer6_outputs(1066) <= not b;
    layer6_outputs(1067) <= a xor b;
    layer6_outputs(1068) <= not (a or b);
    layer6_outputs(1069) <= not b;
    layer6_outputs(1070) <= a or b;
    layer6_outputs(1071) <= a and b;
    layer6_outputs(1072) <= a xor b;
    layer6_outputs(1073) <= a or b;
    layer6_outputs(1074) <= a;
    layer6_outputs(1075) <= '1';
    layer6_outputs(1076) <= a xor b;
    layer6_outputs(1077) <= not a;
    layer6_outputs(1078) <= not a;
    layer6_outputs(1079) <= not b;
    layer6_outputs(1080) <= not (a xor b);
    layer6_outputs(1081) <= a and b;
    layer6_outputs(1082) <= a;
    layer6_outputs(1083) <= b and not a;
    layer6_outputs(1084) <= not (a or b);
    layer6_outputs(1085) <= '0';
    layer6_outputs(1086) <= not (a or b);
    layer6_outputs(1087) <= not b;
    layer6_outputs(1088) <= not (a or b);
    layer6_outputs(1089) <= a xor b;
    layer6_outputs(1090) <= b and not a;
    layer6_outputs(1091) <= a and not b;
    layer6_outputs(1092) <= not (a or b);
    layer6_outputs(1093) <= a or b;
    layer6_outputs(1094) <= b;
    layer6_outputs(1095) <= not (a and b);
    layer6_outputs(1096) <= a and not b;
    layer6_outputs(1097) <= b and not a;
    layer6_outputs(1098) <= b;
    layer6_outputs(1099) <= a and not b;
    layer6_outputs(1100) <= not b or a;
    layer6_outputs(1101) <= '0';
    layer6_outputs(1102) <= not b;
    layer6_outputs(1103) <= not a or b;
    layer6_outputs(1104) <= not a;
    layer6_outputs(1105) <= b;
    layer6_outputs(1106) <= not b;
    layer6_outputs(1107) <= '0';
    layer6_outputs(1108) <= a xor b;
    layer6_outputs(1109) <= not (a and b);
    layer6_outputs(1110) <= not b;
    layer6_outputs(1111) <= a or b;
    layer6_outputs(1112) <= a;
    layer6_outputs(1113) <= a;
    layer6_outputs(1114) <= not a;
    layer6_outputs(1115) <= b;
    layer6_outputs(1116) <= not a or b;
    layer6_outputs(1117) <= not a;
    layer6_outputs(1118) <= not a;
    layer6_outputs(1119) <= b;
    layer6_outputs(1120) <= b and not a;
    layer6_outputs(1121) <= b;
    layer6_outputs(1122) <= not (a or b);
    layer6_outputs(1123) <= not b;
    layer6_outputs(1124) <= not (a xor b);
    layer6_outputs(1125) <= a xor b;
    layer6_outputs(1126) <= a xor b;
    layer6_outputs(1127) <= a and not b;
    layer6_outputs(1128) <= not (a and b);
    layer6_outputs(1129) <= a;
    layer6_outputs(1130) <= '1';
    layer6_outputs(1131) <= b;
    layer6_outputs(1132) <= not b;
    layer6_outputs(1133) <= not a;
    layer6_outputs(1134) <= a;
    layer6_outputs(1135) <= not a or b;
    layer6_outputs(1136) <= not b or a;
    layer6_outputs(1137) <= a or b;
    layer6_outputs(1138) <= not a;
    layer6_outputs(1139) <= b;
    layer6_outputs(1140) <= a and not b;
    layer6_outputs(1141) <= not (a or b);
    layer6_outputs(1142) <= a and b;
    layer6_outputs(1143) <= not b or a;
    layer6_outputs(1144) <= not (a or b);
    layer6_outputs(1145) <= not b;
    layer6_outputs(1146) <= not a;
    layer6_outputs(1147) <= a and not b;
    layer6_outputs(1148) <= a and b;
    layer6_outputs(1149) <= a xor b;
    layer6_outputs(1150) <= a and b;
    layer6_outputs(1151) <= not a;
    layer6_outputs(1152) <= a xor b;
    layer6_outputs(1153) <= not a;
    layer6_outputs(1154) <= '1';
    layer6_outputs(1155) <= b and not a;
    layer6_outputs(1156) <= not (a and b);
    layer6_outputs(1157) <= b;
    layer6_outputs(1158) <= a xor b;
    layer6_outputs(1159) <= a and not b;
    layer6_outputs(1160) <= not a;
    layer6_outputs(1161) <= not a or b;
    layer6_outputs(1162) <= not a or b;
    layer6_outputs(1163) <= not b or a;
    layer6_outputs(1164) <= not b;
    layer6_outputs(1165) <= b;
    layer6_outputs(1166) <= b;
    layer6_outputs(1167) <= not b;
    layer6_outputs(1168) <= not b or a;
    layer6_outputs(1169) <= a xor b;
    layer6_outputs(1170) <= not a;
    layer6_outputs(1171) <= not b;
    layer6_outputs(1172) <= a or b;
    layer6_outputs(1173) <= not b;
    layer6_outputs(1174) <= a;
    layer6_outputs(1175) <= b;
    layer6_outputs(1176) <= not b;
    layer6_outputs(1177) <= '0';
    layer6_outputs(1178) <= not b;
    layer6_outputs(1179) <= not b or a;
    layer6_outputs(1180) <= not b;
    layer6_outputs(1181) <= not b;
    layer6_outputs(1182) <= not b;
    layer6_outputs(1183) <= not b;
    layer6_outputs(1184) <= not b;
    layer6_outputs(1185) <= not a or b;
    layer6_outputs(1186) <= not b;
    layer6_outputs(1187) <= a or b;
    layer6_outputs(1188) <= a;
    layer6_outputs(1189) <= not a or b;
    layer6_outputs(1190) <= not (a xor b);
    layer6_outputs(1191) <= not (a and b);
    layer6_outputs(1192) <= not b;
    layer6_outputs(1193) <= a xor b;
    layer6_outputs(1194) <= a or b;
    layer6_outputs(1195) <= not a or b;
    layer6_outputs(1196) <= a and b;
    layer6_outputs(1197) <= not a or b;
    layer6_outputs(1198) <= not b;
    layer6_outputs(1199) <= a and b;
    layer6_outputs(1200) <= a xor b;
    layer6_outputs(1201) <= '1';
    layer6_outputs(1202) <= a and not b;
    layer6_outputs(1203) <= not b or a;
    layer6_outputs(1204) <= not b or a;
    layer6_outputs(1205) <= a xor b;
    layer6_outputs(1206) <= a or b;
    layer6_outputs(1207) <= b;
    layer6_outputs(1208) <= b;
    layer6_outputs(1209) <= a and not b;
    layer6_outputs(1210) <= a and not b;
    layer6_outputs(1211) <= '1';
    layer6_outputs(1212) <= not (a and b);
    layer6_outputs(1213) <= not (a or b);
    layer6_outputs(1214) <= not (a xor b);
    layer6_outputs(1215) <= a;
    layer6_outputs(1216) <= a or b;
    layer6_outputs(1217) <= b;
    layer6_outputs(1218) <= not (a xor b);
    layer6_outputs(1219) <= a;
    layer6_outputs(1220) <= b;
    layer6_outputs(1221) <= a;
    layer6_outputs(1222) <= not (a and b);
    layer6_outputs(1223) <= a xor b;
    layer6_outputs(1224) <= a and not b;
    layer6_outputs(1225) <= not a;
    layer6_outputs(1226) <= b;
    layer6_outputs(1227) <= not (a or b);
    layer6_outputs(1228) <= not (a and b);
    layer6_outputs(1229) <= not b;
    layer6_outputs(1230) <= a;
    layer6_outputs(1231) <= '0';
    layer6_outputs(1232) <= b and not a;
    layer6_outputs(1233) <= not a or b;
    layer6_outputs(1234) <= not (a and b);
    layer6_outputs(1235) <= a and b;
    layer6_outputs(1236) <= not b;
    layer6_outputs(1237) <= not a;
    layer6_outputs(1238) <= not a or b;
    layer6_outputs(1239) <= not a or b;
    layer6_outputs(1240) <= not (a and b);
    layer6_outputs(1241) <= not b or a;
    layer6_outputs(1242) <= a;
    layer6_outputs(1243) <= not b;
    layer6_outputs(1244) <= not a;
    layer6_outputs(1245) <= not b;
    layer6_outputs(1246) <= not (a xor b);
    layer6_outputs(1247) <= not a;
    layer6_outputs(1248) <= a and not b;
    layer6_outputs(1249) <= a and not b;
    layer6_outputs(1250) <= b and not a;
    layer6_outputs(1251) <= b;
    layer6_outputs(1252) <= b;
    layer6_outputs(1253) <= b;
    layer6_outputs(1254) <= a;
    layer6_outputs(1255) <= a and not b;
    layer6_outputs(1256) <= a xor b;
    layer6_outputs(1257) <= '1';
    layer6_outputs(1258) <= not (a or b);
    layer6_outputs(1259) <= not b or a;
    layer6_outputs(1260) <= a and not b;
    layer6_outputs(1261) <= b and not a;
    layer6_outputs(1262) <= not b or a;
    layer6_outputs(1263) <= '0';
    layer6_outputs(1264) <= b;
    layer6_outputs(1265) <= b and not a;
    layer6_outputs(1266) <= b;
    layer6_outputs(1267) <= b;
    layer6_outputs(1268) <= a and b;
    layer6_outputs(1269) <= not a;
    layer6_outputs(1270) <= not b or a;
    layer6_outputs(1271) <= b and not a;
    layer6_outputs(1272) <= not a;
    layer6_outputs(1273) <= not b or a;
    layer6_outputs(1274) <= a;
    layer6_outputs(1275) <= a xor b;
    layer6_outputs(1276) <= a;
    layer6_outputs(1277) <= a;
    layer6_outputs(1278) <= b;
    layer6_outputs(1279) <= not a;
    layer6_outputs(1280) <= not a or b;
    layer6_outputs(1281) <= not b;
    layer6_outputs(1282) <= a xor b;
    layer6_outputs(1283) <= a and not b;
    layer6_outputs(1284) <= a;
    layer6_outputs(1285) <= b and not a;
    layer6_outputs(1286) <= a and not b;
    layer6_outputs(1287) <= not b;
    layer6_outputs(1288) <= a;
    layer6_outputs(1289) <= '1';
    layer6_outputs(1290) <= b;
    layer6_outputs(1291) <= a;
    layer6_outputs(1292) <= not a;
    layer6_outputs(1293) <= not b;
    layer6_outputs(1294) <= not b;
    layer6_outputs(1295) <= not a or b;
    layer6_outputs(1296) <= a and b;
    layer6_outputs(1297) <= not b or a;
    layer6_outputs(1298) <= b;
    layer6_outputs(1299) <= b and not a;
    layer6_outputs(1300) <= a and b;
    layer6_outputs(1301) <= a;
    layer6_outputs(1302) <= not (a xor b);
    layer6_outputs(1303) <= not a or b;
    layer6_outputs(1304) <= b and not a;
    layer6_outputs(1305) <= not b or a;
    layer6_outputs(1306) <= a;
    layer6_outputs(1307) <= not b;
    layer6_outputs(1308) <= not b;
    layer6_outputs(1309) <= not (a and b);
    layer6_outputs(1310) <= a;
    layer6_outputs(1311) <= '0';
    layer6_outputs(1312) <= not (a and b);
    layer6_outputs(1313) <= not b;
    layer6_outputs(1314) <= not a or b;
    layer6_outputs(1315) <= not b;
    layer6_outputs(1316) <= a;
    layer6_outputs(1317) <= a and not b;
    layer6_outputs(1318) <= b;
    layer6_outputs(1319) <= a and b;
    layer6_outputs(1320) <= not b or a;
    layer6_outputs(1321) <= not (a and b);
    layer6_outputs(1322) <= a and b;
    layer6_outputs(1323) <= not (a and b);
    layer6_outputs(1324) <= a and b;
    layer6_outputs(1325) <= not (a and b);
    layer6_outputs(1326) <= not b;
    layer6_outputs(1327) <= '0';
    layer6_outputs(1328) <= b;
    layer6_outputs(1329) <= not (a xor b);
    layer6_outputs(1330) <= b;
    layer6_outputs(1331) <= a and not b;
    layer6_outputs(1332) <= a or b;
    layer6_outputs(1333) <= not (a xor b);
    layer6_outputs(1334) <= not (a and b);
    layer6_outputs(1335) <= not a or b;
    layer6_outputs(1336) <= not (a and b);
    layer6_outputs(1337) <= a or b;
    layer6_outputs(1338) <= a and not b;
    layer6_outputs(1339) <= not a;
    layer6_outputs(1340) <= b and not a;
    layer6_outputs(1341) <= a and not b;
    layer6_outputs(1342) <= not a or b;
    layer6_outputs(1343) <= a;
    layer6_outputs(1344) <= '0';
    layer6_outputs(1345) <= not (a xor b);
    layer6_outputs(1346) <= '0';
    layer6_outputs(1347) <= a xor b;
    layer6_outputs(1348) <= a;
    layer6_outputs(1349) <= not (a and b);
    layer6_outputs(1350) <= not a;
    layer6_outputs(1351) <= b and not a;
    layer6_outputs(1352) <= '1';
    layer6_outputs(1353) <= b;
    layer6_outputs(1354) <= a xor b;
    layer6_outputs(1355) <= not b;
    layer6_outputs(1356) <= not (a or b);
    layer6_outputs(1357) <= b and not a;
    layer6_outputs(1358) <= not a or b;
    layer6_outputs(1359) <= not a or b;
    layer6_outputs(1360) <= not a or b;
    layer6_outputs(1361) <= a;
    layer6_outputs(1362) <= not a;
    layer6_outputs(1363) <= a;
    layer6_outputs(1364) <= not a;
    layer6_outputs(1365) <= not b;
    layer6_outputs(1366) <= a xor b;
    layer6_outputs(1367) <= b;
    layer6_outputs(1368) <= not b;
    layer6_outputs(1369) <= b;
    layer6_outputs(1370) <= '0';
    layer6_outputs(1371) <= '1';
    layer6_outputs(1372) <= b;
    layer6_outputs(1373) <= not b;
    layer6_outputs(1374) <= '1';
    layer6_outputs(1375) <= a or b;
    layer6_outputs(1376) <= a xor b;
    layer6_outputs(1377) <= a and not b;
    layer6_outputs(1378) <= b and not a;
    layer6_outputs(1379) <= not b;
    layer6_outputs(1380) <= a or b;
    layer6_outputs(1381) <= a and not b;
    layer6_outputs(1382) <= not a;
    layer6_outputs(1383) <= '0';
    layer6_outputs(1384) <= not (a or b);
    layer6_outputs(1385) <= b;
    layer6_outputs(1386) <= not a;
    layer6_outputs(1387) <= not b;
    layer6_outputs(1388) <= not (a and b);
    layer6_outputs(1389) <= a;
    layer6_outputs(1390) <= '0';
    layer6_outputs(1391) <= '0';
    layer6_outputs(1392) <= a xor b;
    layer6_outputs(1393) <= not b;
    layer6_outputs(1394) <= not a;
    layer6_outputs(1395) <= a;
    layer6_outputs(1396) <= not (a and b);
    layer6_outputs(1397) <= not b;
    layer6_outputs(1398) <= b and not a;
    layer6_outputs(1399) <= not b;
    layer6_outputs(1400) <= not a;
    layer6_outputs(1401) <= a;
    layer6_outputs(1402) <= not b or a;
    layer6_outputs(1403) <= b and not a;
    layer6_outputs(1404) <= a xor b;
    layer6_outputs(1405) <= a;
    layer6_outputs(1406) <= not a or b;
    layer6_outputs(1407) <= b;
    layer6_outputs(1408) <= not (a and b);
    layer6_outputs(1409) <= not (a xor b);
    layer6_outputs(1410) <= b;
    layer6_outputs(1411) <= not (a xor b);
    layer6_outputs(1412) <= not (a and b);
    layer6_outputs(1413) <= a;
    layer6_outputs(1414) <= a;
    layer6_outputs(1415) <= a and not b;
    layer6_outputs(1416) <= a;
    layer6_outputs(1417) <= b;
    layer6_outputs(1418) <= not (a xor b);
    layer6_outputs(1419) <= a xor b;
    layer6_outputs(1420) <= not a;
    layer6_outputs(1421) <= not a or b;
    layer6_outputs(1422) <= b;
    layer6_outputs(1423) <= not b;
    layer6_outputs(1424) <= a;
    layer6_outputs(1425) <= a and b;
    layer6_outputs(1426) <= b;
    layer6_outputs(1427) <= a;
    layer6_outputs(1428) <= not a;
    layer6_outputs(1429) <= not (a xor b);
    layer6_outputs(1430) <= not a;
    layer6_outputs(1431) <= not a;
    layer6_outputs(1432) <= a;
    layer6_outputs(1433) <= not a or b;
    layer6_outputs(1434) <= not b;
    layer6_outputs(1435) <= a;
    layer6_outputs(1436) <= a and b;
    layer6_outputs(1437) <= not a or b;
    layer6_outputs(1438) <= not a;
    layer6_outputs(1439) <= not (a xor b);
    layer6_outputs(1440) <= b;
    layer6_outputs(1441) <= a;
    layer6_outputs(1442) <= not a or b;
    layer6_outputs(1443) <= a or b;
    layer6_outputs(1444) <= a;
    layer6_outputs(1445) <= a and not b;
    layer6_outputs(1446) <= a and not b;
    layer6_outputs(1447) <= b and not a;
    layer6_outputs(1448) <= not a or b;
    layer6_outputs(1449) <= not a or b;
    layer6_outputs(1450) <= not a;
    layer6_outputs(1451) <= not (a xor b);
    layer6_outputs(1452) <= a xor b;
    layer6_outputs(1453) <= a;
    layer6_outputs(1454) <= a or b;
    layer6_outputs(1455) <= not b or a;
    layer6_outputs(1456) <= not b or a;
    layer6_outputs(1457) <= not (a and b);
    layer6_outputs(1458) <= a and b;
    layer6_outputs(1459) <= a and not b;
    layer6_outputs(1460) <= not (a or b);
    layer6_outputs(1461) <= b and not a;
    layer6_outputs(1462) <= '0';
    layer6_outputs(1463) <= not b;
    layer6_outputs(1464) <= not (a and b);
    layer6_outputs(1465) <= a xor b;
    layer6_outputs(1466) <= not b;
    layer6_outputs(1467) <= a;
    layer6_outputs(1468) <= a;
    layer6_outputs(1469) <= '0';
    layer6_outputs(1470) <= not b;
    layer6_outputs(1471) <= not b;
    layer6_outputs(1472) <= '1';
    layer6_outputs(1473) <= a or b;
    layer6_outputs(1474) <= not (a xor b);
    layer6_outputs(1475) <= a and b;
    layer6_outputs(1476) <= not a;
    layer6_outputs(1477) <= a;
    layer6_outputs(1478) <= a xor b;
    layer6_outputs(1479) <= '1';
    layer6_outputs(1480) <= a xor b;
    layer6_outputs(1481) <= b;
    layer6_outputs(1482) <= not (a or b);
    layer6_outputs(1483) <= a and b;
    layer6_outputs(1484) <= not b;
    layer6_outputs(1485) <= not b or a;
    layer6_outputs(1486) <= a or b;
    layer6_outputs(1487) <= not a;
    layer6_outputs(1488) <= a and not b;
    layer6_outputs(1489) <= not a;
    layer6_outputs(1490) <= b;
    layer6_outputs(1491) <= not a or b;
    layer6_outputs(1492) <= not a or b;
    layer6_outputs(1493) <= not a;
    layer6_outputs(1494) <= '1';
    layer6_outputs(1495) <= not b or a;
    layer6_outputs(1496) <= not b or a;
    layer6_outputs(1497) <= not a;
    layer6_outputs(1498) <= not (a and b);
    layer6_outputs(1499) <= a or b;
    layer6_outputs(1500) <= a and b;
    layer6_outputs(1501) <= not a or b;
    layer6_outputs(1502) <= not (a or b);
    layer6_outputs(1503) <= b;
    layer6_outputs(1504) <= b;
    layer6_outputs(1505) <= b and not a;
    layer6_outputs(1506) <= a;
    layer6_outputs(1507) <= not a;
    layer6_outputs(1508) <= not (a and b);
    layer6_outputs(1509) <= not b or a;
    layer6_outputs(1510) <= '1';
    layer6_outputs(1511) <= b and not a;
    layer6_outputs(1512) <= not (a and b);
    layer6_outputs(1513) <= b and not a;
    layer6_outputs(1514) <= not a or b;
    layer6_outputs(1515) <= b and not a;
    layer6_outputs(1516) <= a or b;
    layer6_outputs(1517) <= a and b;
    layer6_outputs(1518) <= a;
    layer6_outputs(1519) <= b;
    layer6_outputs(1520) <= not a or b;
    layer6_outputs(1521) <= '1';
    layer6_outputs(1522) <= a and b;
    layer6_outputs(1523) <= not a;
    layer6_outputs(1524) <= not b or a;
    layer6_outputs(1525) <= a and not b;
    layer6_outputs(1526) <= b;
    layer6_outputs(1527) <= a and not b;
    layer6_outputs(1528) <= not a;
    layer6_outputs(1529) <= a and b;
    layer6_outputs(1530) <= not a;
    layer6_outputs(1531) <= not b;
    layer6_outputs(1532) <= not b;
    layer6_outputs(1533) <= a;
    layer6_outputs(1534) <= not (a xor b);
    layer6_outputs(1535) <= not b or a;
    layer6_outputs(1536) <= a;
    layer6_outputs(1537) <= a xor b;
    layer6_outputs(1538) <= b;
    layer6_outputs(1539) <= a or b;
    layer6_outputs(1540) <= a and not b;
    layer6_outputs(1541) <= not b or a;
    layer6_outputs(1542) <= not a;
    layer6_outputs(1543) <= b;
    layer6_outputs(1544) <= not b or a;
    layer6_outputs(1545) <= a xor b;
    layer6_outputs(1546) <= a and not b;
    layer6_outputs(1547) <= a xor b;
    layer6_outputs(1548) <= not a;
    layer6_outputs(1549) <= a xor b;
    layer6_outputs(1550) <= a;
    layer6_outputs(1551) <= not a or b;
    layer6_outputs(1552) <= not a;
    layer6_outputs(1553) <= '0';
    layer6_outputs(1554) <= not (a or b);
    layer6_outputs(1555) <= a and not b;
    layer6_outputs(1556) <= a or b;
    layer6_outputs(1557) <= a;
    layer6_outputs(1558) <= not a;
    layer6_outputs(1559) <= b;
    layer6_outputs(1560) <= not a or b;
    layer6_outputs(1561) <= '1';
    layer6_outputs(1562) <= a;
    layer6_outputs(1563) <= not (a and b);
    layer6_outputs(1564) <= a or b;
    layer6_outputs(1565) <= b;
    layer6_outputs(1566) <= b and not a;
    layer6_outputs(1567) <= not b;
    layer6_outputs(1568) <= not b;
    layer6_outputs(1569) <= not b or a;
    layer6_outputs(1570) <= b and not a;
    layer6_outputs(1571) <= a;
    layer6_outputs(1572) <= not (a or b);
    layer6_outputs(1573) <= a or b;
    layer6_outputs(1574) <= a;
    layer6_outputs(1575) <= a;
    layer6_outputs(1576) <= b and not a;
    layer6_outputs(1577) <= not a;
    layer6_outputs(1578) <= a and b;
    layer6_outputs(1579) <= not b;
    layer6_outputs(1580) <= a;
    layer6_outputs(1581) <= b;
    layer6_outputs(1582) <= not b;
    layer6_outputs(1583) <= not a;
    layer6_outputs(1584) <= b;
    layer6_outputs(1585) <= '1';
    layer6_outputs(1586) <= a;
    layer6_outputs(1587) <= b;
    layer6_outputs(1588) <= a xor b;
    layer6_outputs(1589) <= b;
    layer6_outputs(1590) <= b;
    layer6_outputs(1591) <= not b;
    layer6_outputs(1592) <= not b;
    layer6_outputs(1593) <= b;
    layer6_outputs(1594) <= not (a and b);
    layer6_outputs(1595) <= not a;
    layer6_outputs(1596) <= b;
    layer6_outputs(1597) <= not a;
    layer6_outputs(1598) <= not b;
    layer6_outputs(1599) <= a;
    layer6_outputs(1600) <= a xor b;
    layer6_outputs(1601) <= b;
    layer6_outputs(1602) <= not b;
    layer6_outputs(1603) <= not (a and b);
    layer6_outputs(1604) <= not a or b;
    layer6_outputs(1605) <= not a;
    layer6_outputs(1606) <= b;
    layer6_outputs(1607) <= a and not b;
    layer6_outputs(1608) <= b;
    layer6_outputs(1609) <= not b;
    layer6_outputs(1610) <= a and b;
    layer6_outputs(1611) <= a and not b;
    layer6_outputs(1612) <= not a or b;
    layer6_outputs(1613) <= a and not b;
    layer6_outputs(1614) <= a;
    layer6_outputs(1615) <= not (a and b);
    layer6_outputs(1616) <= a and not b;
    layer6_outputs(1617) <= b;
    layer6_outputs(1618) <= not (a and b);
    layer6_outputs(1619) <= not b or a;
    layer6_outputs(1620) <= not b;
    layer6_outputs(1621) <= not b;
    layer6_outputs(1622) <= a;
    layer6_outputs(1623) <= a and b;
    layer6_outputs(1624) <= not a;
    layer6_outputs(1625) <= not a;
    layer6_outputs(1626) <= a;
    layer6_outputs(1627) <= b and not a;
    layer6_outputs(1628) <= a and not b;
    layer6_outputs(1629) <= a;
    layer6_outputs(1630) <= not b or a;
    layer6_outputs(1631) <= not (a and b);
    layer6_outputs(1632) <= not b;
    layer6_outputs(1633) <= a xor b;
    layer6_outputs(1634) <= not a;
    layer6_outputs(1635) <= not (a or b);
    layer6_outputs(1636) <= b and not a;
    layer6_outputs(1637) <= not b;
    layer6_outputs(1638) <= a;
    layer6_outputs(1639) <= a and not b;
    layer6_outputs(1640) <= not b;
    layer6_outputs(1641) <= not (a and b);
    layer6_outputs(1642) <= b;
    layer6_outputs(1643) <= b;
    layer6_outputs(1644) <= a xor b;
    layer6_outputs(1645) <= a and b;
    layer6_outputs(1646) <= a or b;
    layer6_outputs(1647) <= not b;
    layer6_outputs(1648) <= a or b;
    layer6_outputs(1649) <= b;
    layer6_outputs(1650) <= b and not a;
    layer6_outputs(1651) <= not b;
    layer6_outputs(1652) <= not (a or b);
    layer6_outputs(1653) <= '0';
    layer6_outputs(1654) <= not (a and b);
    layer6_outputs(1655) <= not b or a;
    layer6_outputs(1656) <= a or b;
    layer6_outputs(1657) <= not (a xor b);
    layer6_outputs(1658) <= not a;
    layer6_outputs(1659) <= a and b;
    layer6_outputs(1660) <= not b;
    layer6_outputs(1661) <= a xor b;
    layer6_outputs(1662) <= not a;
    layer6_outputs(1663) <= a or b;
    layer6_outputs(1664) <= a xor b;
    layer6_outputs(1665) <= not b;
    layer6_outputs(1666) <= not (a or b);
    layer6_outputs(1667) <= a and b;
    layer6_outputs(1668) <= a;
    layer6_outputs(1669) <= not (a xor b);
    layer6_outputs(1670) <= a xor b;
    layer6_outputs(1671) <= not (a or b);
    layer6_outputs(1672) <= b;
    layer6_outputs(1673) <= a and b;
    layer6_outputs(1674) <= '0';
    layer6_outputs(1675) <= a xor b;
    layer6_outputs(1676) <= not a;
    layer6_outputs(1677) <= a and b;
    layer6_outputs(1678) <= a xor b;
    layer6_outputs(1679) <= not b or a;
    layer6_outputs(1680) <= not b;
    layer6_outputs(1681) <= not a;
    layer6_outputs(1682) <= a xor b;
    layer6_outputs(1683) <= b and not a;
    layer6_outputs(1684) <= not (a and b);
    layer6_outputs(1685) <= a or b;
    layer6_outputs(1686) <= a and not b;
    layer6_outputs(1687) <= not b or a;
    layer6_outputs(1688) <= b;
    layer6_outputs(1689) <= not (a or b);
    layer6_outputs(1690) <= a and b;
    layer6_outputs(1691) <= b;
    layer6_outputs(1692) <= a xor b;
    layer6_outputs(1693) <= a;
    layer6_outputs(1694) <= not b or a;
    layer6_outputs(1695) <= not b;
    layer6_outputs(1696) <= not b or a;
    layer6_outputs(1697) <= not (a and b);
    layer6_outputs(1698) <= not a;
    layer6_outputs(1699) <= '1';
    layer6_outputs(1700) <= not (a or b);
    layer6_outputs(1701) <= not (a and b);
    layer6_outputs(1702) <= not (a xor b);
    layer6_outputs(1703) <= b and not a;
    layer6_outputs(1704) <= b;
    layer6_outputs(1705) <= a and b;
    layer6_outputs(1706) <= a and b;
    layer6_outputs(1707) <= a and not b;
    layer6_outputs(1708) <= not a;
    layer6_outputs(1709) <= not a or b;
    layer6_outputs(1710) <= b;
    layer6_outputs(1711) <= not (a or b);
    layer6_outputs(1712) <= a;
    layer6_outputs(1713) <= not a;
    layer6_outputs(1714) <= not (a xor b);
    layer6_outputs(1715) <= not (a or b);
    layer6_outputs(1716) <= not b;
    layer6_outputs(1717) <= not b;
    layer6_outputs(1718) <= not b or a;
    layer6_outputs(1719) <= not b;
    layer6_outputs(1720) <= a xor b;
    layer6_outputs(1721) <= not a;
    layer6_outputs(1722) <= a xor b;
    layer6_outputs(1723) <= a xor b;
    layer6_outputs(1724) <= a and not b;
    layer6_outputs(1725) <= not b or a;
    layer6_outputs(1726) <= a;
    layer6_outputs(1727) <= a;
    layer6_outputs(1728) <= not (a and b);
    layer6_outputs(1729) <= not b;
    layer6_outputs(1730) <= b and not a;
    layer6_outputs(1731) <= b;
    layer6_outputs(1732) <= a or b;
    layer6_outputs(1733) <= not a;
    layer6_outputs(1734) <= not b;
    layer6_outputs(1735) <= not (a and b);
    layer6_outputs(1736) <= a;
    layer6_outputs(1737) <= not a;
    layer6_outputs(1738) <= not a or b;
    layer6_outputs(1739) <= not b;
    layer6_outputs(1740) <= a;
    layer6_outputs(1741) <= not b;
    layer6_outputs(1742) <= not b or a;
    layer6_outputs(1743) <= a and b;
    layer6_outputs(1744) <= not b;
    layer6_outputs(1745) <= not a;
    layer6_outputs(1746) <= a xor b;
    layer6_outputs(1747) <= a and not b;
    layer6_outputs(1748) <= a;
    layer6_outputs(1749) <= b;
    layer6_outputs(1750) <= b;
    layer6_outputs(1751) <= not a;
    layer6_outputs(1752) <= a or b;
    layer6_outputs(1753) <= not b;
    layer6_outputs(1754) <= not a or b;
    layer6_outputs(1755) <= not a or b;
    layer6_outputs(1756) <= b and not a;
    layer6_outputs(1757) <= a and b;
    layer6_outputs(1758) <= not a;
    layer6_outputs(1759) <= not b or a;
    layer6_outputs(1760) <= b;
    layer6_outputs(1761) <= b;
    layer6_outputs(1762) <= not b;
    layer6_outputs(1763) <= a;
    layer6_outputs(1764) <= a or b;
    layer6_outputs(1765) <= not a;
    layer6_outputs(1766) <= a or b;
    layer6_outputs(1767) <= a and not b;
    layer6_outputs(1768) <= a and not b;
    layer6_outputs(1769) <= not (a or b);
    layer6_outputs(1770) <= not (a and b);
    layer6_outputs(1771) <= a;
    layer6_outputs(1772) <= not (a xor b);
    layer6_outputs(1773) <= b;
    layer6_outputs(1774) <= a and not b;
    layer6_outputs(1775) <= not b;
    layer6_outputs(1776) <= a xor b;
    layer6_outputs(1777) <= not a;
    layer6_outputs(1778) <= not a or b;
    layer6_outputs(1779) <= not (a or b);
    layer6_outputs(1780) <= not b;
    layer6_outputs(1781) <= not a;
    layer6_outputs(1782) <= a;
    layer6_outputs(1783) <= a;
    layer6_outputs(1784) <= a xor b;
    layer6_outputs(1785) <= a;
    layer6_outputs(1786) <= not a;
    layer6_outputs(1787) <= not (a and b);
    layer6_outputs(1788) <= not a;
    layer6_outputs(1789) <= not b;
    layer6_outputs(1790) <= b;
    layer6_outputs(1791) <= b;
    layer6_outputs(1792) <= not a;
    layer6_outputs(1793) <= a;
    layer6_outputs(1794) <= not (a xor b);
    layer6_outputs(1795) <= b;
    layer6_outputs(1796) <= not b;
    layer6_outputs(1797) <= not (a xor b);
    layer6_outputs(1798) <= a xor b;
    layer6_outputs(1799) <= not a or b;
    layer6_outputs(1800) <= not (a or b);
    layer6_outputs(1801) <= not a or b;
    layer6_outputs(1802) <= not b;
    layer6_outputs(1803) <= a xor b;
    layer6_outputs(1804) <= b;
    layer6_outputs(1805) <= b;
    layer6_outputs(1806) <= b;
    layer6_outputs(1807) <= not a;
    layer6_outputs(1808) <= '0';
    layer6_outputs(1809) <= a or b;
    layer6_outputs(1810) <= not b or a;
    layer6_outputs(1811) <= not b;
    layer6_outputs(1812) <= not (a xor b);
    layer6_outputs(1813) <= a and b;
    layer6_outputs(1814) <= not (a and b);
    layer6_outputs(1815) <= not (a or b);
    layer6_outputs(1816) <= not b or a;
    layer6_outputs(1817) <= b and not a;
    layer6_outputs(1818) <= not a;
    layer6_outputs(1819) <= b;
    layer6_outputs(1820) <= not a;
    layer6_outputs(1821) <= not a;
    layer6_outputs(1822) <= not a;
    layer6_outputs(1823) <= a and not b;
    layer6_outputs(1824) <= '0';
    layer6_outputs(1825) <= not a;
    layer6_outputs(1826) <= not b or a;
    layer6_outputs(1827) <= a and not b;
    layer6_outputs(1828) <= not a or b;
    layer6_outputs(1829) <= a or b;
    layer6_outputs(1830) <= a;
    layer6_outputs(1831) <= not (a xor b);
    layer6_outputs(1832) <= a;
    layer6_outputs(1833) <= not a;
    layer6_outputs(1834) <= not a or b;
    layer6_outputs(1835) <= a xor b;
    layer6_outputs(1836) <= not b;
    layer6_outputs(1837) <= not (a or b);
    layer6_outputs(1838) <= not b or a;
    layer6_outputs(1839) <= not b;
    layer6_outputs(1840) <= not (a xor b);
    layer6_outputs(1841) <= '1';
    layer6_outputs(1842) <= not a;
    layer6_outputs(1843) <= b;
    layer6_outputs(1844) <= a;
    layer6_outputs(1845) <= a or b;
    layer6_outputs(1846) <= a xor b;
    layer6_outputs(1847) <= a and not b;
    layer6_outputs(1848) <= not a;
    layer6_outputs(1849) <= a xor b;
    layer6_outputs(1850) <= not b;
    layer6_outputs(1851) <= not (a xor b);
    layer6_outputs(1852) <= not b;
    layer6_outputs(1853) <= '1';
    layer6_outputs(1854) <= not (a and b);
    layer6_outputs(1855) <= not (a or b);
    layer6_outputs(1856) <= a and b;
    layer6_outputs(1857) <= a xor b;
    layer6_outputs(1858) <= b and not a;
    layer6_outputs(1859) <= '1';
    layer6_outputs(1860) <= b and not a;
    layer6_outputs(1861) <= not (a or b);
    layer6_outputs(1862) <= b;
    layer6_outputs(1863) <= not b;
    layer6_outputs(1864) <= b and not a;
    layer6_outputs(1865) <= not a;
    layer6_outputs(1866) <= not (a and b);
    layer6_outputs(1867) <= b;
    layer6_outputs(1868) <= b;
    layer6_outputs(1869) <= not b;
    layer6_outputs(1870) <= '1';
    layer6_outputs(1871) <= not a or b;
    layer6_outputs(1872) <= not a;
    layer6_outputs(1873) <= not a;
    layer6_outputs(1874) <= '1';
    layer6_outputs(1875) <= not (a and b);
    layer6_outputs(1876) <= a;
    layer6_outputs(1877) <= a;
    layer6_outputs(1878) <= not a;
    layer6_outputs(1879) <= '1';
    layer6_outputs(1880) <= not (a and b);
    layer6_outputs(1881) <= b and not a;
    layer6_outputs(1882) <= a;
    layer6_outputs(1883) <= not (a xor b);
    layer6_outputs(1884) <= a xor b;
    layer6_outputs(1885) <= not b or a;
    layer6_outputs(1886) <= not (a or b);
    layer6_outputs(1887) <= b and not a;
    layer6_outputs(1888) <= a and not b;
    layer6_outputs(1889) <= a xor b;
    layer6_outputs(1890) <= not b;
    layer6_outputs(1891) <= a and b;
    layer6_outputs(1892) <= not (a and b);
    layer6_outputs(1893) <= b;
    layer6_outputs(1894) <= b;
    layer6_outputs(1895) <= not b or a;
    layer6_outputs(1896) <= not (a or b);
    layer6_outputs(1897) <= not (a xor b);
    layer6_outputs(1898) <= b;
    layer6_outputs(1899) <= b;
    layer6_outputs(1900) <= not a;
    layer6_outputs(1901) <= not b;
    layer6_outputs(1902) <= a or b;
    layer6_outputs(1903) <= not (a and b);
    layer6_outputs(1904) <= not b;
    layer6_outputs(1905) <= not a;
    layer6_outputs(1906) <= not (a xor b);
    layer6_outputs(1907) <= b and not a;
    layer6_outputs(1908) <= not b;
    layer6_outputs(1909) <= b;
    layer6_outputs(1910) <= a and not b;
    layer6_outputs(1911) <= a or b;
    layer6_outputs(1912) <= b;
    layer6_outputs(1913) <= not b or a;
    layer6_outputs(1914) <= a and not b;
    layer6_outputs(1915) <= not a or b;
    layer6_outputs(1916) <= not b;
    layer6_outputs(1917) <= not b;
    layer6_outputs(1918) <= a;
    layer6_outputs(1919) <= a and b;
    layer6_outputs(1920) <= not (a xor b);
    layer6_outputs(1921) <= not (a or b);
    layer6_outputs(1922) <= a and not b;
    layer6_outputs(1923) <= not a;
    layer6_outputs(1924) <= b and not a;
    layer6_outputs(1925) <= not b or a;
    layer6_outputs(1926) <= not (a or b);
    layer6_outputs(1927) <= '0';
    layer6_outputs(1928) <= b and not a;
    layer6_outputs(1929) <= b and not a;
    layer6_outputs(1930) <= '1';
    layer6_outputs(1931) <= '0';
    layer6_outputs(1932) <= a;
    layer6_outputs(1933) <= not (a and b);
    layer6_outputs(1934) <= b and not a;
    layer6_outputs(1935) <= not (a or b);
    layer6_outputs(1936) <= not b;
    layer6_outputs(1937) <= not b;
    layer6_outputs(1938) <= not b;
    layer6_outputs(1939) <= a xor b;
    layer6_outputs(1940) <= not b;
    layer6_outputs(1941) <= b;
    layer6_outputs(1942) <= a and not b;
    layer6_outputs(1943) <= not b;
    layer6_outputs(1944) <= not (a xor b);
    layer6_outputs(1945) <= not a or b;
    layer6_outputs(1946) <= a;
    layer6_outputs(1947) <= not (a and b);
    layer6_outputs(1948) <= a and b;
    layer6_outputs(1949) <= not a;
    layer6_outputs(1950) <= a;
    layer6_outputs(1951) <= not (a and b);
    layer6_outputs(1952) <= not b;
    layer6_outputs(1953) <= a or b;
    layer6_outputs(1954) <= a xor b;
    layer6_outputs(1955) <= b and not a;
    layer6_outputs(1956) <= b and not a;
    layer6_outputs(1957) <= not a or b;
    layer6_outputs(1958) <= not (a and b);
    layer6_outputs(1959) <= not (a xor b);
    layer6_outputs(1960) <= not (a xor b);
    layer6_outputs(1961) <= a and not b;
    layer6_outputs(1962) <= not (a and b);
    layer6_outputs(1963) <= not (a xor b);
    layer6_outputs(1964) <= not b or a;
    layer6_outputs(1965) <= b;
    layer6_outputs(1966) <= b;
    layer6_outputs(1967) <= '1';
    layer6_outputs(1968) <= not a or b;
    layer6_outputs(1969) <= b and not a;
    layer6_outputs(1970) <= a and not b;
    layer6_outputs(1971) <= not b;
    layer6_outputs(1972) <= a;
    layer6_outputs(1973) <= a;
    layer6_outputs(1974) <= not (a or b);
    layer6_outputs(1975) <= not (a or b);
    layer6_outputs(1976) <= not b or a;
    layer6_outputs(1977) <= a;
    layer6_outputs(1978) <= b;
    layer6_outputs(1979) <= '1';
    layer6_outputs(1980) <= a;
    layer6_outputs(1981) <= a and not b;
    layer6_outputs(1982) <= '0';
    layer6_outputs(1983) <= a;
    layer6_outputs(1984) <= a and not b;
    layer6_outputs(1985) <= b and not a;
    layer6_outputs(1986) <= not b;
    layer6_outputs(1987) <= a and b;
    layer6_outputs(1988) <= not b;
    layer6_outputs(1989) <= not a;
    layer6_outputs(1990) <= a;
    layer6_outputs(1991) <= not a or b;
    layer6_outputs(1992) <= not a or b;
    layer6_outputs(1993) <= a;
    layer6_outputs(1994) <= not b or a;
    layer6_outputs(1995) <= not b;
    layer6_outputs(1996) <= not (a xor b);
    layer6_outputs(1997) <= not a;
    layer6_outputs(1998) <= not b or a;
    layer6_outputs(1999) <= a;
    layer6_outputs(2000) <= not (a xor b);
    layer6_outputs(2001) <= not a;
    layer6_outputs(2002) <= a;
    layer6_outputs(2003) <= b;
    layer6_outputs(2004) <= a;
    layer6_outputs(2005) <= not b or a;
    layer6_outputs(2006) <= not a;
    layer6_outputs(2007) <= a;
    layer6_outputs(2008) <= a xor b;
    layer6_outputs(2009) <= a and b;
    layer6_outputs(2010) <= a and b;
    layer6_outputs(2011) <= a and not b;
    layer6_outputs(2012) <= not a or b;
    layer6_outputs(2013) <= a and not b;
    layer6_outputs(2014) <= b;
    layer6_outputs(2015) <= b;
    layer6_outputs(2016) <= not a;
    layer6_outputs(2017) <= not b;
    layer6_outputs(2018) <= not a;
    layer6_outputs(2019) <= a and not b;
    layer6_outputs(2020) <= not a;
    layer6_outputs(2021) <= not (a xor b);
    layer6_outputs(2022) <= a or b;
    layer6_outputs(2023) <= a and b;
    layer6_outputs(2024) <= a xor b;
    layer6_outputs(2025) <= a;
    layer6_outputs(2026) <= not a;
    layer6_outputs(2027) <= not b;
    layer6_outputs(2028) <= a and not b;
    layer6_outputs(2029) <= not (a or b);
    layer6_outputs(2030) <= a or b;
    layer6_outputs(2031) <= not (a or b);
    layer6_outputs(2032) <= not b;
    layer6_outputs(2033) <= '0';
    layer6_outputs(2034) <= not (a and b);
    layer6_outputs(2035) <= not (a and b);
    layer6_outputs(2036) <= b;
    layer6_outputs(2037) <= not a;
    layer6_outputs(2038) <= a or b;
    layer6_outputs(2039) <= not b;
    layer6_outputs(2040) <= a or b;
    layer6_outputs(2041) <= not b;
    layer6_outputs(2042) <= not a or b;
    layer6_outputs(2043) <= b;
    layer6_outputs(2044) <= a xor b;
    layer6_outputs(2045) <= not (a and b);
    layer6_outputs(2046) <= not (a and b);
    layer6_outputs(2047) <= not a;
    layer6_outputs(2048) <= not b;
    layer6_outputs(2049) <= not (a or b);
    layer6_outputs(2050) <= not a;
    layer6_outputs(2051) <= b;
    layer6_outputs(2052) <= a;
    layer6_outputs(2053) <= a and b;
    layer6_outputs(2054) <= a;
    layer6_outputs(2055) <= a and b;
    layer6_outputs(2056) <= not (a xor b);
    layer6_outputs(2057) <= not a or b;
    layer6_outputs(2058) <= a or b;
    layer6_outputs(2059) <= not b;
    layer6_outputs(2060) <= not b or a;
    layer6_outputs(2061) <= b;
    layer6_outputs(2062) <= a;
    layer6_outputs(2063) <= b and not a;
    layer6_outputs(2064) <= not (a xor b);
    layer6_outputs(2065) <= a;
    layer6_outputs(2066) <= not (a xor b);
    layer6_outputs(2067) <= not b or a;
    layer6_outputs(2068) <= a;
    layer6_outputs(2069) <= not a;
    layer6_outputs(2070) <= a and b;
    layer6_outputs(2071) <= b;
    layer6_outputs(2072) <= b;
    layer6_outputs(2073) <= b;
    layer6_outputs(2074) <= b;
    layer6_outputs(2075) <= b;
    layer6_outputs(2076) <= a;
    layer6_outputs(2077) <= a;
    layer6_outputs(2078) <= a;
    layer6_outputs(2079) <= a and b;
    layer6_outputs(2080) <= not (a and b);
    layer6_outputs(2081) <= not b;
    layer6_outputs(2082) <= not (a or b);
    layer6_outputs(2083) <= not a;
    layer6_outputs(2084) <= not b or a;
    layer6_outputs(2085) <= b;
    layer6_outputs(2086) <= not (a xor b);
    layer6_outputs(2087) <= a or b;
    layer6_outputs(2088) <= not a;
    layer6_outputs(2089) <= b and not a;
    layer6_outputs(2090) <= not a;
    layer6_outputs(2091) <= not b or a;
    layer6_outputs(2092) <= not a;
    layer6_outputs(2093) <= a;
    layer6_outputs(2094) <= not b;
    layer6_outputs(2095) <= not b;
    layer6_outputs(2096) <= b and not a;
    layer6_outputs(2097) <= not b or a;
    layer6_outputs(2098) <= not a;
    layer6_outputs(2099) <= not b;
    layer6_outputs(2100) <= a and not b;
    layer6_outputs(2101) <= a xor b;
    layer6_outputs(2102) <= not b;
    layer6_outputs(2103) <= b and not a;
    layer6_outputs(2104) <= a;
    layer6_outputs(2105) <= not a or b;
    layer6_outputs(2106) <= a and b;
    layer6_outputs(2107) <= b;
    layer6_outputs(2108) <= not b;
    layer6_outputs(2109) <= not a;
    layer6_outputs(2110) <= a;
    layer6_outputs(2111) <= not (a or b);
    layer6_outputs(2112) <= b;
    layer6_outputs(2113) <= not (a or b);
    layer6_outputs(2114) <= not a;
    layer6_outputs(2115) <= not (a or b);
    layer6_outputs(2116) <= not a or b;
    layer6_outputs(2117) <= not (a or b);
    layer6_outputs(2118) <= not b;
    layer6_outputs(2119) <= '1';
    layer6_outputs(2120) <= a xor b;
    layer6_outputs(2121) <= not (a xor b);
    layer6_outputs(2122) <= not a;
    layer6_outputs(2123) <= a or b;
    layer6_outputs(2124) <= a xor b;
    layer6_outputs(2125) <= not a;
    layer6_outputs(2126) <= not b;
    layer6_outputs(2127) <= not (a and b);
    layer6_outputs(2128) <= a;
    layer6_outputs(2129) <= a;
    layer6_outputs(2130) <= '1';
    layer6_outputs(2131) <= not (a and b);
    layer6_outputs(2132) <= b;
    layer6_outputs(2133) <= not b or a;
    layer6_outputs(2134) <= not (a xor b);
    layer6_outputs(2135) <= a or b;
    layer6_outputs(2136) <= a and not b;
    layer6_outputs(2137) <= not (a and b);
    layer6_outputs(2138) <= a and b;
    layer6_outputs(2139) <= not b or a;
    layer6_outputs(2140) <= a;
    layer6_outputs(2141) <= not b or a;
    layer6_outputs(2142) <= not a;
    layer6_outputs(2143) <= a or b;
    layer6_outputs(2144) <= b and not a;
    layer6_outputs(2145) <= a xor b;
    layer6_outputs(2146) <= not (a or b);
    layer6_outputs(2147) <= not a or b;
    layer6_outputs(2148) <= not b or a;
    layer6_outputs(2149) <= b;
    layer6_outputs(2150) <= a;
    layer6_outputs(2151) <= not a;
    layer6_outputs(2152) <= not (a and b);
    layer6_outputs(2153) <= not a;
    layer6_outputs(2154) <= not a or b;
    layer6_outputs(2155) <= b and not a;
    layer6_outputs(2156) <= not b;
    layer6_outputs(2157) <= a xor b;
    layer6_outputs(2158) <= '1';
    layer6_outputs(2159) <= b and not a;
    layer6_outputs(2160) <= not (a or b);
    layer6_outputs(2161) <= a and b;
    layer6_outputs(2162) <= a or b;
    layer6_outputs(2163) <= a or b;
    layer6_outputs(2164) <= not b;
    layer6_outputs(2165) <= not (a xor b);
    layer6_outputs(2166) <= a and b;
    layer6_outputs(2167) <= b and not a;
    layer6_outputs(2168) <= b;
    layer6_outputs(2169) <= a or b;
    layer6_outputs(2170) <= not (a and b);
    layer6_outputs(2171) <= not (a or b);
    layer6_outputs(2172) <= b;
    layer6_outputs(2173) <= b;
    layer6_outputs(2174) <= not a or b;
    layer6_outputs(2175) <= not b;
    layer6_outputs(2176) <= a;
    layer6_outputs(2177) <= not (a xor b);
    layer6_outputs(2178) <= not (a or b);
    layer6_outputs(2179) <= not b;
    layer6_outputs(2180) <= not a;
    layer6_outputs(2181) <= '1';
    layer6_outputs(2182) <= not b;
    layer6_outputs(2183) <= not a;
    layer6_outputs(2184) <= not (a xor b);
    layer6_outputs(2185) <= not (a and b);
    layer6_outputs(2186) <= a;
    layer6_outputs(2187) <= not b;
    layer6_outputs(2188) <= a or b;
    layer6_outputs(2189) <= b;
    layer6_outputs(2190) <= not a;
    layer6_outputs(2191) <= not a;
    layer6_outputs(2192) <= not b;
    layer6_outputs(2193) <= a xor b;
    layer6_outputs(2194) <= a or b;
    layer6_outputs(2195) <= not a;
    layer6_outputs(2196) <= not b;
    layer6_outputs(2197) <= not b or a;
    layer6_outputs(2198) <= not (a or b);
    layer6_outputs(2199) <= a and b;
    layer6_outputs(2200) <= not a;
    layer6_outputs(2201) <= not a or b;
    layer6_outputs(2202) <= a;
    layer6_outputs(2203) <= not (a and b);
    layer6_outputs(2204) <= not a or b;
    layer6_outputs(2205) <= a;
    layer6_outputs(2206) <= not (a or b);
    layer6_outputs(2207) <= not b;
    layer6_outputs(2208) <= not b;
    layer6_outputs(2209) <= a;
    layer6_outputs(2210) <= '1';
    layer6_outputs(2211) <= not a;
    layer6_outputs(2212) <= not a;
    layer6_outputs(2213) <= b;
    layer6_outputs(2214) <= a and b;
    layer6_outputs(2215) <= '1';
    layer6_outputs(2216) <= not a;
    layer6_outputs(2217) <= not a;
    layer6_outputs(2218) <= a;
    layer6_outputs(2219) <= a and not b;
    layer6_outputs(2220) <= a and not b;
    layer6_outputs(2221) <= not a or b;
    layer6_outputs(2222) <= a or b;
    layer6_outputs(2223) <= b;
    layer6_outputs(2224) <= not b;
    layer6_outputs(2225) <= b;
    layer6_outputs(2226) <= a xor b;
    layer6_outputs(2227) <= not (a and b);
    layer6_outputs(2228) <= not b;
    layer6_outputs(2229) <= not (a xor b);
    layer6_outputs(2230) <= not b;
    layer6_outputs(2231) <= a xor b;
    layer6_outputs(2232) <= not a or b;
    layer6_outputs(2233) <= not (a or b);
    layer6_outputs(2234) <= a;
    layer6_outputs(2235) <= not b;
    layer6_outputs(2236) <= a and b;
    layer6_outputs(2237) <= not b or a;
    layer6_outputs(2238) <= b and not a;
    layer6_outputs(2239) <= b;
    layer6_outputs(2240) <= not (a or b);
    layer6_outputs(2241) <= a and b;
    layer6_outputs(2242) <= a or b;
    layer6_outputs(2243) <= a xor b;
    layer6_outputs(2244) <= not (a xor b);
    layer6_outputs(2245) <= a or b;
    layer6_outputs(2246) <= '0';
    layer6_outputs(2247) <= not (a xor b);
    layer6_outputs(2248) <= '1';
    layer6_outputs(2249) <= a or b;
    layer6_outputs(2250) <= not b;
    layer6_outputs(2251) <= a xor b;
    layer6_outputs(2252) <= b;
    layer6_outputs(2253) <= not (a and b);
    layer6_outputs(2254) <= a and not b;
    layer6_outputs(2255) <= a and not b;
    layer6_outputs(2256) <= a or b;
    layer6_outputs(2257) <= b;
    layer6_outputs(2258) <= '0';
    layer6_outputs(2259) <= a xor b;
    layer6_outputs(2260) <= '0';
    layer6_outputs(2261) <= b and not a;
    layer6_outputs(2262) <= not b;
    layer6_outputs(2263) <= not (a and b);
    layer6_outputs(2264) <= a xor b;
    layer6_outputs(2265) <= not (a xor b);
    layer6_outputs(2266) <= b;
    layer6_outputs(2267) <= not a;
    layer6_outputs(2268) <= b and not a;
    layer6_outputs(2269) <= not a;
    layer6_outputs(2270) <= not a;
    layer6_outputs(2271) <= not a or b;
    layer6_outputs(2272) <= not (a and b);
    layer6_outputs(2273) <= not (a and b);
    layer6_outputs(2274) <= a xor b;
    layer6_outputs(2275) <= a;
    layer6_outputs(2276) <= not b;
    layer6_outputs(2277) <= not b;
    layer6_outputs(2278) <= a;
    layer6_outputs(2279) <= not a or b;
    layer6_outputs(2280) <= b and not a;
    layer6_outputs(2281) <= not a;
    layer6_outputs(2282) <= not b;
    layer6_outputs(2283) <= b and not a;
    layer6_outputs(2284) <= a xor b;
    layer6_outputs(2285) <= b and not a;
    layer6_outputs(2286) <= b;
    layer6_outputs(2287) <= not a;
    layer6_outputs(2288) <= b;
    layer6_outputs(2289) <= not b or a;
    layer6_outputs(2290) <= not (a or b);
    layer6_outputs(2291) <= not (a xor b);
    layer6_outputs(2292) <= b and not a;
    layer6_outputs(2293) <= b;
    layer6_outputs(2294) <= a or b;
    layer6_outputs(2295) <= not (a or b);
    layer6_outputs(2296) <= a or b;
    layer6_outputs(2297) <= not (a or b);
    layer6_outputs(2298) <= not b;
    layer6_outputs(2299) <= '1';
    layer6_outputs(2300) <= not (a xor b);
    layer6_outputs(2301) <= not (a and b);
    layer6_outputs(2302) <= not b;
    layer6_outputs(2303) <= a or b;
    layer6_outputs(2304) <= b and not a;
    layer6_outputs(2305) <= not a or b;
    layer6_outputs(2306) <= not (a and b);
    layer6_outputs(2307) <= b and not a;
    layer6_outputs(2308) <= a xor b;
    layer6_outputs(2309) <= not a;
    layer6_outputs(2310) <= not (a and b);
    layer6_outputs(2311) <= b and not a;
    layer6_outputs(2312) <= a and not b;
    layer6_outputs(2313) <= a and not b;
    layer6_outputs(2314) <= not b;
    layer6_outputs(2315) <= a;
    layer6_outputs(2316) <= a;
    layer6_outputs(2317) <= b;
    layer6_outputs(2318) <= b and not a;
    layer6_outputs(2319) <= a;
    layer6_outputs(2320) <= not a or b;
    layer6_outputs(2321) <= b and not a;
    layer6_outputs(2322) <= not (a xor b);
    layer6_outputs(2323) <= not b or a;
    layer6_outputs(2324) <= a and not b;
    layer6_outputs(2325) <= a xor b;
    layer6_outputs(2326) <= not a or b;
    layer6_outputs(2327) <= a xor b;
    layer6_outputs(2328) <= not (a xor b);
    layer6_outputs(2329) <= a or b;
    layer6_outputs(2330) <= a xor b;
    layer6_outputs(2331) <= a and b;
    layer6_outputs(2332) <= not b;
    layer6_outputs(2333) <= a and not b;
    layer6_outputs(2334) <= a;
    layer6_outputs(2335) <= not a or b;
    layer6_outputs(2336) <= not a;
    layer6_outputs(2337) <= not a or b;
    layer6_outputs(2338) <= not a;
    layer6_outputs(2339) <= a;
    layer6_outputs(2340) <= b;
    layer6_outputs(2341) <= not (a xor b);
    layer6_outputs(2342) <= not a or b;
    layer6_outputs(2343) <= not (a xor b);
    layer6_outputs(2344) <= a and not b;
    layer6_outputs(2345) <= '0';
    layer6_outputs(2346) <= a or b;
    layer6_outputs(2347) <= a xor b;
    layer6_outputs(2348) <= not (a or b);
    layer6_outputs(2349) <= a xor b;
    layer6_outputs(2350) <= '0';
    layer6_outputs(2351) <= b;
    layer6_outputs(2352) <= not a;
    layer6_outputs(2353) <= a;
    layer6_outputs(2354) <= a xor b;
    layer6_outputs(2355) <= '1';
    layer6_outputs(2356) <= b and not a;
    layer6_outputs(2357) <= not b;
    layer6_outputs(2358) <= a;
    layer6_outputs(2359) <= not b;
    layer6_outputs(2360) <= a and not b;
    layer6_outputs(2361) <= a;
    layer6_outputs(2362) <= a and not b;
    layer6_outputs(2363) <= not b;
    layer6_outputs(2364) <= b and not a;
    layer6_outputs(2365) <= not (a or b);
    layer6_outputs(2366) <= not a;
    layer6_outputs(2367) <= b and not a;
    layer6_outputs(2368) <= a and not b;
    layer6_outputs(2369) <= b and not a;
    layer6_outputs(2370) <= not (a and b);
    layer6_outputs(2371) <= not a;
    layer6_outputs(2372) <= a or b;
    layer6_outputs(2373) <= a or b;
    layer6_outputs(2374) <= not (a xor b);
    layer6_outputs(2375) <= not a or b;
    layer6_outputs(2376) <= a;
    layer6_outputs(2377) <= not (a or b);
    layer6_outputs(2378) <= a;
    layer6_outputs(2379) <= not b;
    layer6_outputs(2380) <= not (a xor b);
    layer6_outputs(2381) <= b and not a;
    layer6_outputs(2382) <= a and b;
    layer6_outputs(2383) <= a xor b;
    layer6_outputs(2384) <= not b;
    layer6_outputs(2385) <= a and not b;
    layer6_outputs(2386) <= not (a or b);
    layer6_outputs(2387) <= not b or a;
    layer6_outputs(2388) <= a or b;
    layer6_outputs(2389) <= not b;
    layer6_outputs(2390) <= not b;
    layer6_outputs(2391) <= a and b;
    layer6_outputs(2392) <= a and b;
    layer6_outputs(2393) <= not (a and b);
    layer6_outputs(2394) <= b;
    layer6_outputs(2395) <= not a;
    layer6_outputs(2396) <= not (a and b);
    layer6_outputs(2397) <= not (a xor b);
    layer6_outputs(2398) <= not (a and b);
    layer6_outputs(2399) <= not (a or b);
    layer6_outputs(2400) <= not a;
    layer6_outputs(2401) <= not (a or b);
    layer6_outputs(2402) <= not a;
    layer6_outputs(2403) <= a or b;
    layer6_outputs(2404) <= not a;
    layer6_outputs(2405) <= not (a xor b);
    layer6_outputs(2406) <= a;
    layer6_outputs(2407) <= not b or a;
    layer6_outputs(2408) <= b;
    layer6_outputs(2409) <= not (a xor b);
    layer6_outputs(2410) <= a;
    layer6_outputs(2411) <= not (a xor b);
    layer6_outputs(2412) <= a or b;
    layer6_outputs(2413) <= a and b;
    layer6_outputs(2414) <= a xor b;
    layer6_outputs(2415) <= a;
    layer6_outputs(2416) <= b and not a;
    layer6_outputs(2417) <= not a or b;
    layer6_outputs(2418) <= a;
    layer6_outputs(2419) <= not a;
    layer6_outputs(2420) <= not a;
    layer6_outputs(2421) <= not a;
    layer6_outputs(2422) <= a;
    layer6_outputs(2423) <= a and not b;
    layer6_outputs(2424) <= '0';
    layer6_outputs(2425) <= not a or b;
    layer6_outputs(2426) <= a or b;
    layer6_outputs(2427) <= a and not b;
    layer6_outputs(2428) <= not b or a;
    layer6_outputs(2429) <= a;
    layer6_outputs(2430) <= not a;
    layer6_outputs(2431) <= not (a and b);
    layer6_outputs(2432) <= a or b;
    layer6_outputs(2433) <= b and not a;
    layer6_outputs(2434) <= not (a or b);
    layer6_outputs(2435) <= a and b;
    layer6_outputs(2436) <= not (a or b);
    layer6_outputs(2437) <= b;
    layer6_outputs(2438) <= a;
    layer6_outputs(2439) <= not b or a;
    layer6_outputs(2440) <= not b;
    layer6_outputs(2441) <= not b or a;
    layer6_outputs(2442) <= a xor b;
    layer6_outputs(2443) <= a;
    layer6_outputs(2444) <= b;
    layer6_outputs(2445) <= not (a xor b);
    layer6_outputs(2446) <= b and not a;
    layer6_outputs(2447) <= '0';
    layer6_outputs(2448) <= a xor b;
    layer6_outputs(2449) <= not b;
    layer6_outputs(2450) <= '1';
    layer6_outputs(2451) <= a or b;
    layer6_outputs(2452) <= not a or b;
    layer6_outputs(2453) <= a and b;
    layer6_outputs(2454) <= b and not a;
    layer6_outputs(2455) <= b and not a;
    layer6_outputs(2456) <= not (a xor b);
    layer6_outputs(2457) <= not (a or b);
    layer6_outputs(2458) <= a xor b;
    layer6_outputs(2459) <= not b;
    layer6_outputs(2460) <= a xor b;
    layer6_outputs(2461) <= a or b;
    layer6_outputs(2462) <= a xor b;
    layer6_outputs(2463) <= b and not a;
    layer6_outputs(2464) <= b;
    layer6_outputs(2465) <= not b;
    layer6_outputs(2466) <= not (a and b);
    layer6_outputs(2467) <= not b;
    layer6_outputs(2468) <= b and not a;
    layer6_outputs(2469) <= a;
    layer6_outputs(2470) <= a;
    layer6_outputs(2471) <= '1';
    layer6_outputs(2472) <= not (a or b);
    layer6_outputs(2473) <= not (a or b);
    layer6_outputs(2474) <= a;
    layer6_outputs(2475) <= a or b;
    layer6_outputs(2476) <= not a or b;
    layer6_outputs(2477) <= not b;
    layer6_outputs(2478) <= not a;
    layer6_outputs(2479) <= not a;
    layer6_outputs(2480) <= not b;
    layer6_outputs(2481) <= a and b;
    layer6_outputs(2482) <= not b;
    layer6_outputs(2483) <= not b or a;
    layer6_outputs(2484) <= a or b;
    layer6_outputs(2485) <= b;
    layer6_outputs(2486) <= b and not a;
    layer6_outputs(2487) <= b and not a;
    layer6_outputs(2488) <= a xor b;
    layer6_outputs(2489) <= a and b;
    layer6_outputs(2490) <= b;
    layer6_outputs(2491) <= b and not a;
    layer6_outputs(2492) <= b;
    layer6_outputs(2493) <= a;
    layer6_outputs(2494) <= not (a or b);
    layer6_outputs(2495) <= not (a xor b);
    layer6_outputs(2496) <= not (a and b);
    layer6_outputs(2497) <= not b;
    layer6_outputs(2498) <= b and not a;
    layer6_outputs(2499) <= not b;
    layer6_outputs(2500) <= not b or a;
    layer6_outputs(2501) <= not (a and b);
    layer6_outputs(2502) <= b;
    layer6_outputs(2503) <= a;
    layer6_outputs(2504) <= '1';
    layer6_outputs(2505) <= a and b;
    layer6_outputs(2506) <= a xor b;
    layer6_outputs(2507) <= a and not b;
    layer6_outputs(2508) <= a or b;
    layer6_outputs(2509) <= not b;
    layer6_outputs(2510) <= a and not b;
    layer6_outputs(2511) <= a or b;
    layer6_outputs(2512) <= not b;
    layer6_outputs(2513) <= a;
    layer6_outputs(2514) <= b and not a;
    layer6_outputs(2515) <= b;
    layer6_outputs(2516) <= not b or a;
    layer6_outputs(2517) <= a;
    layer6_outputs(2518) <= a or b;
    layer6_outputs(2519) <= b;
    layer6_outputs(2520) <= not (a xor b);
    layer6_outputs(2521) <= not b;
    layer6_outputs(2522) <= not (a xor b);
    layer6_outputs(2523) <= not b;
    layer6_outputs(2524) <= a and b;
    layer6_outputs(2525) <= not (a and b);
    layer6_outputs(2526) <= a xor b;
    layer6_outputs(2527) <= not a or b;
    layer6_outputs(2528) <= not b or a;
    layer6_outputs(2529) <= b and not a;
    layer6_outputs(2530) <= not a;
    layer6_outputs(2531) <= not a;
    layer6_outputs(2532) <= not (a or b);
    layer6_outputs(2533) <= not a or b;
    layer6_outputs(2534) <= not (a or b);
    layer6_outputs(2535) <= a;
    layer6_outputs(2536) <= not a or b;
    layer6_outputs(2537) <= not (a or b);
    layer6_outputs(2538) <= not (a xor b);
    layer6_outputs(2539) <= a or b;
    layer6_outputs(2540) <= b;
    layer6_outputs(2541) <= not (a or b);
    layer6_outputs(2542) <= not b or a;
    layer6_outputs(2543) <= a xor b;
    layer6_outputs(2544) <= a and b;
    layer6_outputs(2545) <= not (a or b);
    layer6_outputs(2546) <= not (a xor b);
    layer6_outputs(2547) <= a and b;
    layer6_outputs(2548) <= a xor b;
    layer6_outputs(2549) <= not (a or b);
    layer6_outputs(2550) <= not b or a;
    layer6_outputs(2551) <= not b or a;
    layer6_outputs(2552) <= b and not a;
    layer6_outputs(2553) <= not a;
    layer6_outputs(2554) <= b and not a;
    layer6_outputs(2555) <= not b;
    layer6_outputs(2556) <= not a;
    layer6_outputs(2557) <= a;
    layer6_outputs(2558) <= b;
    layer6_outputs(2559) <= not a;
    layer6_outputs(2560) <= not b;
    layer6_outputs(2561) <= not a or b;
    layer6_outputs(2562) <= not b or a;
    layer6_outputs(2563) <= not (a or b);
    layer6_outputs(2564) <= b;
    layer6_outputs(2565) <= b and not a;
    layer6_outputs(2566) <= a and b;
    layer6_outputs(2567) <= not (a xor b);
    layer6_outputs(2568) <= not (a xor b);
    layer6_outputs(2569) <= a and not b;
    layer6_outputs(2570) <= a xor b;
    layer6_outputs(2571) <= a and b;
    layer6_outputs(2572) <= not a;
    layer6_outputs(2573) <= a;
    layer6_outputs(2574) <= not a;
    layer6_outputs(2575) <= '0';
    layer6_outputs(2576) <= not b or a;
    layer6_outputs(2577) <= b and not a;
    layer6_outputs(2578) <= not (a and b);
    layer6_outputs(2579) <= b;
    layer6_outputs(2580) <= a and b;
    layer6_outputs(2581) <= a and not b;
    layer6_outputs(2582) <= not a or b;
    layer6_outputs(2583) <= a and not b;
    layer6_outputs(2584) <= not b;
    layer6_outputs(2585) <= a xor b;
    layer6_outputs(2586) <= a and not b;
    layer6_outputs(2587) <= b;
    layer6_outputs(2588) <= not b;
    layer6_outputs(2589) <= not b;
    layer6_outputs(2590) <= not (a xor b);
    layer6_outputs(2591) <= not a or b;
    layer6_outputs(2592) <= not b or a;
    layer6_outputs(2593) <= not (a or b);
    layer6_outputs(2594) <= a and not b;
    layer6_outputs(2595) <= not b;
    layer6_outputs(2596) <= not b;
    layer6_outputs(2597) <= b;
    layer6_outputs(2598) <= a and b;
    layer6_outputs(2599) <= a and not b;
    layer6_outputs(2600) <= a;
    layer6_outputs(2601) <= not (a or b);
    layer6_outputs(2602) <= '1';
    layer6_outputs(2603) <= not (a and b);
    layer6_outputs(2604) <= a and b;
    layer6_outputs(2605) <= not b or a;
    layer6_outputs(2606) <= not b;
    layer6_outputs(2607) <= b;
    layer6_outputs(2608) <= a and not b;
    layer6_outputs(2609) <= not (a xor b);
    layer6_outputs(2610) <= not a or b;
    layer6_outputs(2611) <= a or b;
    layer6_outputs(2612) <= a and b;
    layer6_outputs(2613) <= b and not a;
    layer6_outputs(2614) <= b and not a;
    layer6_outputs(2615) <= not b;
    layer6_outputs(2616) <= b and not a;
    layer6_outputs(2617) <= not a;
    layer6_outputs(2618) <= not (a and b);
    layer6_outputs(2619) <= not (a or b);
    layer6_outputs(2620) <= a xor b;
    layer6_outputs(2621) <= a xor b;
    layer6_outputs(2622) <= a or b;
    layer6_outputs(2623) <= a xor b;
    layer6_outputs(2624) <= a;
    layer6_outputs(2625) <= b;
    layer6_outputs(2626) <= b and not a;
    layer6_outputs(2627) <= b;
    layer6_outputs(2628) <= a xor b;
    layer6_outputs(2629) <= b and not a;
    layer6_outputs(2630) <= not (a xor b);
    layer6_outputs(2631) <= not b or a;
    layer6_outputs(2632) <= a;
    layer6_outputs(2633) <= a and not b;
    layer6_outputs(2634) <= a and not b;
    layer6_outputs(2635) <= not (a and b);
    layer6_outputs(2636) <= a or b;
    layer6_outputs(2637) <= a and not b;
    layer6_outputs(2638) <= not b;
    layer6_outputs(2639) <= not (a and b);
    layer6_outputs(2640) <= not b or a;
    layer6_outputs(2641) <= not a or b;
    layer6_outputs(2642) <= a;
    layer6_outputs(2643) <= not b;
    layer6_outputs(2644) <= a and b;
    layer6_outputs(2645) <= a xor b;
    layer6_outputs(2646) <= not (a or b);
    layer6_outputs(2647) <= not (a and b);
    layer6_outputs(2648) <= not (a or b);
    layer6_outputs(2649) <= '0';
    layer6_outputs(2650) <= b;
    layer6_outputs(2651) <= a;
    layer6_outputs(2652) <= not a or b;
    layer6_outputs(2653) <= not a;
    layer6_outputs(2654) <= a xor b;
    layer6_outputs(2655) <= not (a and b);
    layer6_outputs(2656) <= not a;
    layer6_outputs(2657) <= not a;
    layer6_outputs(2658) <= b;
    layer6_outputs(2659) <= not a or b;
    layer6_outputs(2660) <= not a;
    layer6_outputs(2661) <= not a;
    layer6_outputs(2662) <= not b;
    layer6_outputs(2663) <= not a;
    layer6_outputs(2664) <= not a;
    layer6_outputs(2665) <= b;
    layer6_outputs(2666) <= not (a xor b);
    layer6_outputs(2667) <= not b;
    layer6_outputs(2668) <= a and not b;
    layer6_outputs(2669) <= a and not b;
    layer6_outputs(2670) <= a;
    layer6_outputs(2671) <= a and not b;
    layer6_outputs(2672) <= not a;
    layer6_outputs(2673) <= not b;
    layer6_outputs(2674) <= not a;
    layer6_outputs(2675) <= not (a and b);
    layer6_outputs(2676) <= not (a and b);
    layer6_outputs(2677) <= a and not b;
    layer6_outputs(2678) <= a;
    layer6_outputs(2679) <= b;
    layer6_outputs(2680) <= a;
    layer6_outputs(2681) <= not a;
    layer6_outputs(2682) <= a or b;
    layer6_outputs(2683) <= not a or b;
    layer6_outputs(2684) <= not (a or b);
    layer6_outputs(2685) <= a xor b;
    layer6_outputs(2686) <= not b;
    layer6_outputs(2687) <= not b;
    layer6_outputs(2688) <= not b;
    layer6_outputs(2689) <= not a;
    layer6_outputs(2690) <= not a;
    layer6_outputs(2691) <= a;
    layer6_outputs(2692) <= a and b;
    layer6_outputs(2693) <= a;
    layer6_outputs(2694) <= a and not b;
    layer6_outputs(2695) <= not a or b;
    layer6_outputs(2696) <= b;
    layer6_outputs(2697) <= not b or a;
    layer6_outputs(2698) <= not b;
    layer6_outputs(2699) <= b;
    layer6_outputs(2700) <= a xor b;
    layer6_outputs(2701) <= a and b;
    layer6_outputs(2702) <= b;
    layer6_outputs(2703) <= b;
    layer6_outputs(2704) <= not a;
    layer6_outputs(2705) <= not (a xor b);
    layer6_outputs(2706) <= a and b;
    layer6_outputs(2707) <= not b or a;
    layer6_outputs(2708) <= not (a or b);
    layer6_outputs(2709) <= not b or a;
    layer6_outputs(2710) <= not (a xor b);
    layer6_outputs(2711) <= a xor b;
    layer6_outputs(2712) <= a;
    layer6_outputs(2713) <= a;
    layer6_outputs(2714) <= not b;
    layer6_outputs(2715) <= b and not a;
    layer6_outputs(2716) <= a and b;
    layer6_outputs(2717) <= a and not b;
    layer6_outputs(2718) <= b;
    layer6_outputs(2719) <= a xor b;
    layer6_outputs(2720) <= not a;
    layer6_outputs(2721) <= a or b;
    layer6_outputs(2722) <= not (a xor b);
    layer6_outputs(2723) <= not a;
    layer6_outputs(2724) <= not a or b;
    layer6_outputs(2725) <= a xor b;
    layer6_outputs(2726) <= b;
    layer6_outputs(2727) <= a xor b;
    layer6_outputs(2728) <= b;
    layer6_outputs(2729) <= not a or b;
    layer6_outputs(2730) <= not (a or b);
    layer6_outputs(2731) <= not b;
    layer6_outputs(2732) <= b and not a;
    layer6_outputs(2733) <= b;
    layer6_outputs(2734) <= not a or b;
    layer6_outputs(2735) <= not (a and b);
    layer6_outputs(2736) <= a;
    layer6_outputs(2737) <= b and not a;
    layer6_outputs(2738) <= not a or b;
    layer6_outputs(2739) <= not (a or b);
    layer6_outputs(2740) <= a or b;
    layer6_outputs(2741) <= not b;
    layer6_outputs(2742) <= not (a and b);
    layer6_outputs(2743) <= not b;
    layer6_outputs(2744) <= not (a xor b);
    layer6_outputs(2745) <= a;
    layer6_outputs(2746) <= not a;
    layer6_outputs(2747) <= b;
    layer6_outputs(2748) <= '1';
    layer6_outputs(2749) <= b and not a;
    layer6_outputs(2750) <= not b or a;
    layer6_outputs(2751) <= a;
    layer6_outputs(2752) <= a;
    layer6_outputs(2753) <= b;
    layer6_outputs(2754) <= a and not b;
    layer6_outputs(2755) <= not b;
    layer6_outputs(2756) <= b;
    layer6_outputs(2757) <= '1';
    layer6_outputs(2758) <= not b;
    layer6_outputs(2759) <= not a;
    layer6_outputs(2760) <= a or b;
    layer6_outputs(2761) <= b;
    layer6_outputs(2762) <= b;
    layer6_outputs(2763) <= not a or b;
    layer6_outputs(2764) <= b;
    layer6_outputs(2765) <= not (a or b);
    layer6_outputs(2766) <= not b;
    layer6_outputs(2767) <= b and not a;
    layer6_outputs(2768) <= a xor b;
    layer6_outputs(2769) <= not a or b;
    layer6_outputs(2770) <= a xor b;
    layer6_outputs(2771) <= b;
    layer6_outputs(2772) <= not a or b;
    layer6_outputs(2773) <= not (a or b);
    layer6_outputs(2774) <= a or b;
    layer6_outputs(2775) <= b;
    layer6_outputs(2776) <= b;
    layer6_outputs(2777) <= '1';
    layer6_outputs(2778) <= not (a and b);
    layer6_outputs(2779) <= not b;
    layer6_outputs(2780) <= not (a or b);
    layer6_outputs(2781) <= a and b;
    layer6_outputs(2782) <= b and not a;
    layer6_outputs(2783) <= not (a or b);
    layer6_outputs(2784) <= not a;
    layer6_outputs(2785) <= not b or a;
    layer6_outputs(2786) <= a or b;
    layer6_outputs(2787) <= not (a and b);
    layer6_outputs(2788) <= a;
    layer6_outputs(2789) <= not (a or b);
    layer6_outputs(2790) <= not a or b;
    layer6_outputs(2791) <= b;
    layer6_outputs(2792) <= '1';
    layer6_outputs(2793) <= b and not a;
    layer6_outputs(2794) <= a;
    layer6_outputs(2795) <= b and not a;
    layer6_outputs(2796) <= a and not b;
    layer6_outputs(2797) <= a or b;
    layer6_outputs(2798) <= b and not a;
    layer6_outputs(2799) <= b;
    layer6_outputs(2800) <= a and b;
    layer6_outputs(2801) <= not (a and b);
    layer6_outputs(2802) <= not (a or b);
    layer6_outputs(2803) <= not (a xor b);
    layer6_outputs(2804) <= '1';
    layer6_outputs(2805) <= not a;
    layer6_outputs(2806) <= not a or b;
    layer6_outputs(2807) <= not (a and b);
    layer6_outputs(2808) <= b;
    layer6_outputs(2809) <= not a or b;
    layer6_outputs(2810) <= not a or b;
    layer6_outputs(2811) <= a xor b;
    layer6_outputs(2812) <= b and not a;
    layer6_outputs(2813) <= a xor b;
    layer6_outputs(2814) <= not a or b;
    layer6_outputs(2815) <= a;
    layer6_outputs(2816) <= a or b;
    layer6_outputs(2817) <= not b or a;
    layer6_outputs(2818) <= not a or b;
    layer6_outputs(2819) <= a and not b;
    layer6_outputs(2820) <= not b or a;
    layer6_outputs(2821) <= a and b;
    layer6_outputs(2822) <= not b;
    layer6_outputs(2823) <= b;
    layer6_outputs(2824) <= not (a xor b);
    layer6_outputs(2825) <= not a or b;
    layer6_outputs(2826) <= b;
    layer6_outputs(2827) <= '1';
    layer6_outputs(2828) <= not a or b;
    layer6_outputs(2829) <= not b;
    layer6_outputs(2830) <= a and b;
    layer6_outputs(2831) <= a and b;
    layer6_outputs(2832) <= not a;
    layer6_outputs(2833) <= b;
    layer6_outputs(2834) <= not b or a;
    layer6_outputs(2835) <= not a or b;
    layer6_outputs(2836) <= not a;
    layer6_outputs(2837) <= a and b;
    layer6_outputs(2838) <= not (a xor b);
    layer6_outputs(2839) <= a and b;
    layer6_outputs(2840) <= not a;
    layer6_outputs(2841) <= not b;
    layer6_outputs(2842) <= not (a and b);
    layer6_outputs(2843) <= '0';
    layer6_outputs(2844) <= a;
    layer6_outputs(2845) <= a and not b;
    layer6_outputs(2846) <= not a;
    layer6_outputs(2847) <= not b;
    layer6_outputs(2848) <= not (a and b);
    layer6_outputs(2849) <= not b;
    layer6_outputs(2850) <= b;
    layer6_outputs(2851) <= b;
    layer6_outputs(2852) <= a xor b;
    layer6_outputs(2853) <= not a or b;
    layer6_outputs(2854) <= a;
    layer6_outputs(2855) <= not (a xor b);
    layer6_outputs(2856) <= a and not b;
    layer6_outputs(2857) <= not a or b;
    layer6_outputs(2858) <= not b or a;
    layer6_outputs(2859) <= not (a or b);
    layer6_outputs(2860) <= a and not b;
    layer6_outputs(2861) <= a and b;
    layer6_outputs(2862) <= not a or b;
    layer6_outputs(2863) <= not a or b;
    layer6_outputs(2864) <= a;
    layer6_outputs(2865) <= not b;
    layer6_outputs(2866) <= not a;
    layer6_outputs(2867) <= not a;
    layer6_outputs(2868) <= not b;
    layer6_outputs(2869) <= not a;
    layer6_outputs(2870) <= '0';
    layer6_outputs(2871) <= a or b;
    layer6_outputs(2872) <= a;
    layer6_outputs(2873) <= '1';
    layer6_outputs(2874) <= a and not b;
    layer6_outputs(2875) <= not b or a;
    layer6_outputs(2876) <= not a or b;
    layer6_outputs(2877) <= not a or b;
    layer6_outputs(2878) <= not a;
    layer6_outputs(2879) <= b;
    layer6_outputs(2880) <= not (a and b);
    layer6_outputs(2881) <= a and not b;
    layer6_outputs(2882) <= not (a and b);
    layer6_outputs(2883) <= not b;
    layer6_outputs(2884) <= b;
    layer6_outputs(2885) <= not b;
    layer6_outputs(2886) <= not a or b;
    layer6_outputs(2887) <= a xor b;
    layer6_outputs(2888) <= not (a xor b);
    layer6_outputs(2889) <= a;
    layer6_outputs(2890) <= not a or b;
    layer6_outputs(2891) <= '0';
    layer6_outputs(2892) <= a or b;
    layer6_outputs(2893) <= not b;
    layer6_outputs(2894) <= not (a or b);
    layer6_outputs(2895) <= b;
    layer6_outputs(2896) <= not b;
    layer6_outputs(2897) <= b and not a;
    layer6_outputs(2898) <= a;
    layer6_outputs(2899) <= a xor b;
    layer6_outputs(2900) <= not a;
    layer6_outputs(2901) <= a or b;
    layer6_outputs(2902) <= not b or a;
    layer6_outputs(2903) <= a;
    layer6_outputs(2904) <= b and not a;
    layer6_outputs(2905) <= not b or a;
    layer6_outputs(2906) <= '0';
    layer6_outputs(2907) <= a xor b;
    layer6_outputs(2908) <= not (a and b);
    layer6_outputs(2909) <= b;
    layer6_outputs(2910) <= not b or a;
    layer6_outputs(2911) <= not (a or b);
    layer6_outputs(2912) <= '0';
    layer6_outputs(2913) <= b;
    layer6_outputs(2914) <= b and not a;
    layer6_outputs(2915) <= a or b;
    layer6_outputs(2916) <= a and b;
    layer6_outputs(2917) <= not (a and b);
    layer6_outputs(2918) <= a and not b;
    layer6_outputs(2919) <= b;
    layer6_outputs(2920) <= not b;
    layer6_outputs(2921) <= not a;
    layer6_outputs(2922) <= a xor b;
    layer6_outputs(2923) <= not a;
    layer6_outputs(2924) <= a;
    layer6_outputs(2925) <= not b;
    layer6_outputs(2926) <= a xor b;
    layer6_outputs(2927) <= not a;
    layer6_outputs(2928) <= not b or a;
    layer6_outputs(2929) <= not (a and b);
    layer6_outputs(2930) <= not a;
    layer6_outputs(2931) <= not b;
    layer6_outputs(2932) <= a and b;
    layer6_outputs(2933) <= not (a and b);
    layer6_outputs(2934) <= not (a or b);
    layer6_outputs(2935) <= not (a or b);
    layer6_outputs(2936) <= not a;
    layer6_outputs(2937) <= b and not a;
    layer6_outputs(2938) <= b;
    layer6_outputs(2939) <= not (a xor b);
    layer6_outputs(2940) <= not (a xor b);
    layer6_outputs(2941) <= not (a and b);
    layer6_outputs(2942) <= not b;
    layer6_outputs(2943) <= not b or a;
    layer6_outputs(2944) <= not a or b;
    layer6_outputs(2945) <= not b;
    layer6_outputs(2946) <= a;
    layer6_outputs(2947) <= not (a xor b);
    layer6_outputs(2948) <= not (a or b);
    layer6_outputs(2949) <= not b;
    layer6_outputs(2950) <= not (a and b);
    layer6_outputs(2951) <= not (a and b);
    layer6_outputs(2952) <= not a or b;
    layer6_outputs(2953) <= not (a or b);
    layer6_outputs(2954) <= a and b;
    layer6_outputs(2955) <= not a or b;
    layer6_outputs(2956) <= a;
    layer6_outputs(2957) <= not a;
    layer6_outputs(2958) <= not (a xor b);
    layer6_outputs(2959) <= not a or b;
    layer6_outputs(2960) <= not b;
    layer6_outputs(2961) <= a;
    layer6_outputs(2962) <= a or b;
    layer6_outputs(2963) <= not a or b;
    layer6_outputs(2964) <= not a;
    layer6_outputs(2965) <= a and not b;
    layer6_outputs(2966) <= a;
    layer6_outputs(2967) <= not b or a;
    layer6_outputs(2968) <= not a;
    layer6_outputs(2969) <= '0';
    layer6_outputs(2970) <= not a or b;
    layer6_outputs(2971) <= not b;
    layer6_outputs(2972) <= a or b;
    layer6_outputs(2973) <= not b;
    layer6_outputs(2974) <= not (a or b);
    layer6_outputs(2975) <= not b;
    layer6_outputs(2976) <= not b;
    layer6_outputs(2977) <= a;
    layer6_outputs(2978) <= b;
    layer6_outputs(2979) <= not b;
    layer6_outputs(2980) <= b and not a;
    layer6_outputs(2981) <= not b;
    layer6_outputs(2982) <= a and b;
    layer6_outputs(2983) <= not a;
    layer6_outputs(2984) <= not a or b;
    layer6_outputs(2985) <= not b;
    layer6_outputs(2986) <= not b;
    layer6_outputs(2987) <= not a;
    layer6_outputs(2988) <= not b;
    layer6_outputs(2989) <= a;
    layer6_outputs(2990) <= not (a and b);
    layer6_outputs(2991) <= not (a and b);
    layer6_outputs(2992) <= a xor b;
    layer6_outputs(2993) <= not (a and b);
    layer6_outputs(2994) <= a or b;
    layer6_outputs(2995) <= not a or b;
    layer6_outputs(2996) <= not a;
    layer6_outputs(2997) <= '0';
    layer6_outputs(2998) <= b;
    layer6_outputs(2999) <= not (a or b);
    layer6_outputs(3000) <= not (a or b);
    layer6_outputs(3001) <= a xor b;
    layer6_outputs(3002) <= a and b;
    layer6_outputs(3003) <= a and b;
    layer6_outputs(3004) <= not a;
    layer6_outputs(3005) <= a and b;
    layer6_outputs(3006) <= not b or a;
    layer6_outputs(3007) <= not a or b;
    layer6_outputs(3008) <= b and not a;
    layer6_outputs(3009) <= b;
    layer6_outputs(3010) <= a or b;
    layer6_outputs(3011) <= not a;
    layer6_outputs(3012) <= a and not b;
    layer6_outputs(3013) <= b;
    layer6_outputs(3014) <= b and not a;
    layer6_outputs(3015) <= a or b;
    layer6_outputs(3016) <= not (a or b);
    layer6_outputs(3017) <= not a;
    layer6_outputs(3018) <= '1';
    layer6_outputs(3019) <= not a;
    layer6_outputs(3020) <= not (a and b);
    layer6_outputs(3021) <= not a;
    layer6_outputs(3022) <= b;
    layer6_outputs(3023) <= a;
    layer6_outputs(3024) <= a;
    layer6_outputs(3025) <= not a;
    layer6_outputs(3026) <= '0';
    layer6_outputs(3027) <= not b;
    layer6_outputs(3028) <= a;
    layer6_outputs(3029) <= b;
    layer6_outputs(3030) <= not a or b;
    layer6_outputs(3031) <= b and not a;
    layer6_outputs(3032) <= not a;
    layer6_outputs(3033) <= a or b;
    layer6_outputs(3034) <= a or b;
    layer6_outputs(3035) <= not a;
    layer6_outputs(3036) <= not a;
    layer6_outputs(3037) <= not a;
    layer6_outputs(3038) <= not b or a;
    layer6_outputs(3039) <= not b;
    layer6_outputs(3040) <= not a or b;
    layer6_outputs(3041) <= not (a xor b);
    layer6_outputs(3042) <= not a or b;
    layer6_outputs(3043) <= not a or b;
    layer6_outputs(3044) <= a;
    layer6_outputs(3045) <= a or b;
    layer6_outputs(3046) <= a or b;
    layer6_outputs(3047) <= a;
    layer6_outputs(3048) <= '1';
    layer6_outputs(3049) <= a xor b;
    layer6_outputs(3050) <= b and not a;
    layer6_outputs(3051) <= b;
    layer6_outputs(3052) <= not b;
    layer6_outputs(3053) <= not b;
    layer6_outputs(3054) <= a and not b;
    layer6_outputs(3055) <= a;
    layer6_outputs(3056) <= a and not b;
    layer6_outputs(3057) <= not a;
    layer6_outputs(3058) <= '1';
    layer6_outputs(3059) <= b and not a;
    layer6_outputs(3060) <= not (a xor b);
    layer6_outputs(3061) <= not b;
    layer6_outputs(3062) <= not a;
    layer6_outputs(3063) <= not b;
    layer6_outputs(3064) <= not b;
    layer6_outputs(3065) <= a and b;
    layer6_outputs(3066) <= a;
    layer6_outputs(3067) <= a and not b;
    layer6_outputs(3068) <= not a;
    layer6_outputs(3069) <= b;
    layer6_outputs(3070) <= not a or b;
    layer6_outputs(3071) <= not a;
    layer6_outputs(3072) <= not (a or b);
    layer6_outputs(3073) <= not (a and b);
    layer6_outputs(3074) <= b;
    layer6_outputs(3075) <= b;
    layer6_outputs(3076) <= not (a and b);
    layer6_outputs(3077) <= not (a and b);
    layer6_outputs(3078) <= not (a and b);
    layer6_outputs(3079) <= not (a xor b);
    layer6_outputs(3080) <= a xor b;
    layer6_outputs(3081) <= a;
    layer6_outputs(3082) <= b;
    layer6_outputs(3083) <= b;
    layer6_outputs(3084) <= a;
    layer6_outputs(3085) <= b;
    layer6_outputs(3086) <= a xor b;
    layer6_outputs(3087) <= not b or a;
    layer6_outputs(3088) <= b and not a;
    layer6_outputs(3089) <= not b or a;
    layer6_outputs(3090) <= not b or a;
    layer6_outputs(3091) <= not (a or b);
    layer6_outputs(3092) <= not (a or b);
    layer6_outputs(3093) <= b and not a;
    layer6_outputs(3094) <= a;
    layer6_outputs(3095) <= a;
    layer6_outputs(3096) <= b;
    layer6_outputs(3097) <= not (a or b);
    layer6_outputs(3098) <= a and not b;
    layer6_outputs(3099) <= a;
    layer6_outputs(3100) <= b and not a;
    layer6_outputs(3101) <= not a or b;
    layer6_outputs(3102) <= not a or b;
    layer6_outputs(3103) <= b;
    layer6_outputs(3104) <= a;
    layer6_outputs(3105) <= not (a and b);
    layer6_outputs(3106) <= not b or a;
    layer6_outputs(3107) <= not b;
    layer6_outputs(3108) <= b and not a;
    layer6_outputs(3109) <= not (a xor b);
    layer6_outputs(3110) <= a xor b;
    layer6_outputs(3111) <= a xor b;
    layer6_outputs(3112) <= not (a and b);
    layer6_outputs(3113) <= not a;
    layer6_outputs(3114) <= not b;
    layer6_outputs(3115) <= a;
    layer6_outputs(3116) <= not a;
    layer6_outputs(3117) <= '0';
    layer6_outputs(3118) <= not a;
    layer6_outputs(3119) <= not a;
    layer6_outputs(3120) <= a and b;
    layer6_outputs(3121) <= b and not a;
    layer6_outputs(3122) <= not a or b;
    layer6_outputs(3123) <= not (a xor b);
    layer6_outputs(3124) <= not b;
    layer6_outputs(3125) <= not b or a;
    layer6_outputs(3126) <= b and not a;
    layer6_outputs(3127) <= not (a or b);
    layer6_outputs(3128) <= not (a xor b);
    layer6_outputs(3129) <= b and not a;
    layer6_outputs(3130) <= not b;
    layer6_outputs(3131) <= not b;
    layer6_outputs(3132) <= a;
    layer6_outputs(3133) <= not (a and b);
    layer6_outputs(3134) <= not a;
    layer6_outputs(3135) <= not a;
    layer6_outputs(3136) <= b;
    layer6_outputs(3137) <= not b;
    layer6_outputs(3138) <= a or b;
    layer6_outputs(3139) <= not b or a;
    layer6_outputs(3140) <= b;
    layer6_outputs(3141) <= not (a and b);
    layer6_outputs(3142) <= not b or a;
    layer6_outputs(3143) <= b;
    layer6_outputs(3144) <= not (a and b);
    layer6_outputs(3145) <= a;
    layer6_outputs(3146) <= not b;
    layer6_outputs(3147) <= a xor b;
    layer6_outputs(3148) <= not b;
    layer6_outputs(3149) <= not a;
    layer6_outputs(3150) <= a xor b;
    layer6_outputs(3151) <= a and b;
    layer6_outputs(3152) <= '1';
    layer6_outputs(3153) <= not (a or b);
    layer6_outputs(3154) <= not (a and b);
    layer6_outputs(3155) <= b and not a;
    layer6_outputs(3156) <= a;
    layer6_outputs(3157) <= a or b;
    layer6_outputs(3158) <= a;
    layer6_outputs(3159) <= not (a and b);
    layer6_outputs(3160) <= b;
    layer6_outputs(3161) <= not b;
    layer6_outputs(3162) <= b;
    layer6_outputs(3163) <= '0';
    layer6_outputs(3164) <= a;
    layer6_outputs(3165) <= not b or a;
    layer6_outputs(3166) <= a xor b;
    layer6_outputs(3167) <= not a or b;
    layer6_outputs(3168) <= not b;
    layer6_outputs(3169) <= not (a and b);
    layer6_outputs(3170) <= b;
    layer6_outputs(3171) <= a or b;
    layer6_outputs(3172) <= b and not a;
    layer6_outputs(3173) <= a xor b;
    layer6_outputs(3174) <= not a;
    layer6_outputs(3175) <= not a;
    layer6_outputs(3176) <= not a or b;
    layer6_outputs(3177) <= a and not b;
    layer6_outputs(3178) <= a or b;
    layer6_outputs(3179) <= a;
    layer6_outputs(3180) <= a xor b;
    layer6_outputs(3181) <= a or b;
    layer6_outputs(3182) <= b and not a;
    layer6_outputs(3183) <= a;
    layer6_outputs(3184) <= a;
    layer6_outputs(3185) <= a and not b;
    layer6_outputs(3186) <= a;
    layer6_outputs(3187) <= a;
    layer6_outputs(3188) <= not b;
    layer6_outputs(3189) <= not b or a;
    layer6_outputs(3190) <= not b or a;
    layer6_outputs(3191) <= not a;
    layer6_outputs(3192) <= not b;
    layer6_outputs(3193) <= not (a or b);
    layer6_outputs(3194) <= not (a or b);
    layer6_outputs(3195) <= not b;
    layer6_outputs(3196) <= not a;
    layer6_outputs(3197) <= a;
    layer6_outputs(3198) <= not (a or b);
    layer6_outputs(3199) <= '0';
    layer6_outputs(3200) <= a;
    layer6_outputs(3201) <= not b or a;
    layer6_outputs(3202) <= not (a and b);
    layer6_outputs(3203) <= '1';
    layer6_outputs(3204) <= a and not b;
    layer6_outputs(3205) <= a;
    layer6_outputs(3206) <= a and b;
    layer6_outputs(3207) <= a xor b;
    layer6_outputs(3208) <= not (a xor b);
    layer6_outputs(3209) <= a xor b;
    layer6_outputs(3210) <= not a;
    layer6_outputs(3211) <= not a;
    layer6_outputs(3212) <= not b;
    layer6_outputs(3213) <= a;
    layer6_outputs(3214) <= not b or a;
    layer6_outputs(3215) <= not b;
    layer6_outputs(3216) <= not b;
    layer6_outputs(3217) <= a xor b;
    layer6_outputs(3218) <= a and not b;
    layer6_outputs(3219) <= not a;
    layer6_outputs(3220) <= not a;
    layer6_outputs(3221) <= not (a or b);
    layer6_outputs(3222) <= not (a xor b);
    layer6_outputs(3223) <= not a;
    layer6_outputs(3224) <= '1';
    layer6_outputs(3225) <= b;
    layer6_outputs(3226) <= a;
    layer6_outputs(3227) <= a and not b;
    layer6_outputs(3228) <= not (a xor b);
    layer6_outputs(3229) <= not (a and b);
    layer6_outputs(3230) <= b;
    layer6_outputs(3231) <= a and not b;
    layer6_outputs(3232) <= not b;
    layer6_outputs(3233) <= a;
    layer6_outputs(3234) <= b and not a;
    layer6_outputs(3235) <= not a or b;
    layer6_outputs(3236) <= not (a or b);
    layer6_outputs(3237) <= not a or b;
    layer6_outputs(3238) <= not a;
    layer6_outputs(3239) <= not (a xor b);
    layer6_outputs(3240) <= a and not b;
    layer6_outputs(3241) <= not b or a;
    layer6_outputs(3242) <= b;
    layer6_outputs(3243) <= b;
    layer6_outputs(3244) <= a and not b;
    layer6_outputs(3245) <= a and not b;
    layer6_outputs(3246) <= not (a and b);
    layer6_outputs(3247) <= b and not a;
    layer6_outputs(3248) <= a;
    layer6_outputs(3249) <= '0';
    layer6_outputs(3250) <= b;
    layer6_outputs(3251) <= b and not a;
    layer6_outputs(3252) <= not b or a;
    layer6_outputs(3253) <= b;
    layer6_outputs(3254) <= not (a and b);
    layer6_outputs(3255) <= not (a and b);
    layer6_outputs(3256) <= a;
    layer6_outputs(3257) <= not b;
    layer6_outputs(3258) <= '1';
    layer6_outputs(3259) <= not b;
    layer6_outputs(3260) <= a or b;
    layer6_outputs(3261) <= not (a and b);
    layer6_outputs(3262) <= b;
    layer6_outputs(3263) <= not (a or b);
    layer6_outputs(3264) <= not b or a;
    layer6_outputs(3265) <= a or b;
    layer6_outputs(3266) <= not (a xor b);
    layer6_outputs(3267) <= a and b;
    layer6_outputs(3268) <= not a;
    layer6_outputs(3269) <= a and b;
    layer6_outputs(3270) <= not a;
    layer6_outputs(3271) <= not a or b;
    layer6_outputs(3272) <= not (a xor b);
    layer6_outputs(3273) <= not b;
    layer6_outputs(3274) <= not (a or b);
    layer6_outputs(3275) <= a and b;
    layer6_outputs(3276) <= not b;
    layer6_outputs(3277) <= a and not b;
    layer6_outputs(3278) <= not b or a;
    layer6_outputs(3279) <= not b;
    layer6_outputs(3280) <= not a;
    layer6_outputs(3281) <= a;
    layer6_outputs(3282) <= not (a and b);
    layer6_outputs(3283) <= a and b;
    layer6_outputs(3284) <= a or b;
    layer6_outputs(3285) <= not (a or b);
    layer6_outputs(3286) <= a and b;
    layer6_outputs(3287) <= a;
    layer6_outputs(3288) <= a;
    layer6_outputs(3289) <= '1';
    layer6_outputs(3290) <= a;
    layer6_outputs(3291) <= '1';
    layer6_outputs(3292) <= a;
    layer6_outputs(3293) <= a or b;
    layer6_outputs(3294) <= not (a and b);
    layer6_outputs(3295) <= b and not a;
    layer6_outputs(3296) <= a or b;
    layer6_outputs(3297) <= not a;
    layer6_outputs(3298) <= a xor b;
    layer6_outputs(3299) <= a and b;
    layer6_outputs(3300) <= not (a xor b);
    layer6_outputs(3301) <= a and b;
    layer6_outputs(3302) <= not a;
    layer6_outputs(3303) <= a or b;
    layer6_outputs(3304) <= a;
    layer6_outputs(3305) <= b;
    layer6_outputs(3306) <= a and b;
    layer6_outputs(3307) <= not (a and b);
    layer6_outputs(3308) <= a and b;
    layer6_outputs(3309) <= a xor b;
    layer6_outputs(3310) <= not a;
    layer6_outputs(3311) <= not b;
    layer6_outputs(3312) <= a and not b;
    layer6_outputs(3313) <= a xor b;
    layer6_outputs(3314) <= '0';
    layer6_outputs(3315) <= '0';
    layer6_outputs(3316) <= a;
    layer6_outputs(3317) <= not (a or b);
    layer6_outputs(3318) <= '0';
    layer6_outputs(3319) <= b;
    layer6_outputs(3320) <= '1';
    layer6_outputs(3321) <= a and not b;
    layer6_outputs(3322) <= '1';
    layer6_outputs(3323) <= not b or a;
    layer6_outputs(3324) <= a;
    layer6_outputs(3325) <= a;
    layer6_outputs(3326) <= a and b;
    layer6_outputs(3327) <= a and not b;
    layer6_outputs(3328) <= not a;
    layer6_outputs(3329) <= a and not b;
    layer6_outputs(3330) <= not a;
    layer6_outputs(3331) <= a and b;
    layer6_outputs(3332) <= not b;
    layer6_outputs(3333) <= a;
    layer6_outputs(3334) <= not b;
    layer6_outputs(3335) <= b;
    layer6_outputs(3336) <= not (a or b);
    layer6_outputs(3337) <= not a;
    layer6_outputs(3338) <= not b or a;
    layer6_outputs(3339) <= not (a or b);
    layer6_outputs(3340) <= not b;
    layer6_outputs(3341) <= not a;
    layer6_outputs(3342) <= '0';
    layer6_outputs(3343) <= a and not b;
    layer6_outputs(3344) <= not (a and b);
    layer6_outputs(3345) <= not (a and b);
    layer6_outputs(3346) <= a and b;
    layer6_outputs(3347) <= a and b;
    layer6_outputs(3348) <= b;
    layer6_outputs(3349) <= '0';
    layer6_outputs(3350) <= a and not b;
    layer6_outputs(3351) <= not (a or b);
    layer6_outputs(3352) <= not (a or b);
    layer6_outputs(3353) <= '1';
    layer6_outputs(3354) <= not a;
    layer6_outputs(3355) <= a;
    layer6_outputs(3356) <= not a;
    layer6_outputs(3357) <= not b or a;
    layer6_outputs(3358) <= a;
    layer6_outputs(3359) <= not (a or b);
    layer6_outputs(3360) <= not (a and b);
    layer6_outputs(3361) <= not a or b;
    layer6_outputs(3362) <= not a or b;
    layer6_outputs(3363) <= a and b;
    layer6_outputs(3364) <= a;
    layer6_outputs(3365) <= not (a and b);
    layer6_outputs(3366) <= not b or a;
    layer6_outputs(3367) <= a or b;
    layer6_outputs(3368) <= b;
    layer6_outputs(3369) <= not (a and b);
    layer6_outputs(3370) <= b;
    layer6_outputs(3371) <= not b;
    layer6_outputs(3372) <= b and not a;
    layer6_outputs(3373) <= '1';
    layer6_outputs(3374) <= not (a and b);
    layer6_outputs(3375) <= not b;
    layer6_outputs(3376) <= '1';
    layer6_outputs(3377) <= not (a or b);
    layer6_outputs(3378) <= '1';
    layer6_outputs(3379) <= a;
    layer6_outputs(3380) <= b and not a;
    layer6_outputs(3381) <= a or b;
    layer6_outputs(3382) <= not a;
    layer6_outputs(3383) <= not a;
    layer6_outputs(3384) <= not a;
    layer6_outputs(3385) <= not (a xor b);
    layer6_outputs(3386) <= a or b;
    layer6_outputs(3387) <= not b or a;
    layer6_outputs(3388) <= a and not b;
    layer6_outputs(3389) <= not b;
    layer6_outputs(3390) <= a and b;
    layer6_outputs(3391) <= a xor b;
    layer6_outputs(3392) <= not (a xor b);
    layer6_outputs(3393) <= not b or a;
    layer6_outputs(3394) <= a and b;
    layer6_outputs(3395) <= a;
    layer6_outputs(3396) <= not (a or b);
    layer6_outputs(3397) <= a;
    layer6_outputs(3398) <= not b;
    layer6_outputs(3399) <= not b;
    layer6_outputs(3400) <= a;
    layer6_outputs(3401) <= a and b;
    layer6_outputs(3402) <= b;
    layer6_outputs(3403) <= not (a and b);
    layer6_outputs(3404) <= a and b;
    layer6_outputs(3405) <= not a;
    layer6_outputs(3406) <= a and not b;
    layer6_outputs(3407) <= b;
    layer6_outputs(3408) <= not a;
    layer6_outputs(3409) <= b and not a;
    layer6_outputs(3410) <= b;
    layer6_outputs(3411) <= not b or a;
    layer6_outputs(3412) <= not a;
    layer6_outputs(3413) <= not a or b;
    layer6_outputs(3414) <= a;
    layer6_outputs(3415) <= a;
    layer6_outputs(3416) <= not a;
    layer6_outputs(3417) <= not a;
    layer6_outputs(3418) <= a and b;
    layer6_outputs(3419) <= a or b;
    layer6_outputs(3420) <= not a;
    layer6_outputs(3421) <= not (a or b);
    layer6_outputs(3422) <= a xor b;
    layer6_outputs(3423) <= not (a xor b);
    layer6_outputs(3424) <= b;
    layer6_outputs(3425) <= not a;
    layer6_outputs(3426) <= b;
    layer6_outputs(3427) <= a xor b;
    layer6_outputs(3428) <= a;
    layer6_outputs(3429) <= not a;
    layer6_outputs(3430) <= not a;
    layer6_outputs(3431) <= not a or b;
    layer6_outputs(3432) <= a xor b;
    layer6_outputs(3433) <= not b;
    layer6_outputs(3434) <= not (a or b);
    layer6_outputs(3435) <= not b or a;
    layer6_outputs(3436) <= b;
    layer6_outputs(3437) <= a or b;
    layer6_outputs(3438) <= a and not b;
    layer6_outputs(3439) <= not a;
    layer6_outputs(3440) <= b;
    layer6_outputs(3441) <= a or b;
    layer6_outputs(3442) <= not a;
    layer6_outputs(3443) <= not b;
    layer6_outputs(3444) <= b;
    layer6_outputs(3445) <= not a or b;
    layer6_outputs(3446) <= not a;
    layer6_outputs(3447) <= not a;
    layer6_outputs(3448) <= not b;
    layer6_outputs(3449) <= a and b;
    layer6_outputs(3450) <= b and not a;
    layer6_outputs(3451) <= a xor b;
    layer6_outputs(3452) <= not b;
    layer6_outputs(3453) <= b;
    layer6_outputs(3454) <= a;
    layer6_outputs(3455) <= not b;
    layer6_outputs(3456) <= not (a or b);
    layer6_outputs(3457) <= b;
    layer6_outputs(3458) <= not (a or b);
    layer6_outputs(3459) <= a and b;
    layer6_outputs(3460) <= not b;
    layer6_outputs(3461) <= a;
    layer6_outputs(3462) <= not a;
    layer6_outputs(3463) <= b;
    layer6_outputs(3464) <= a and not b;
    layer6_outputs(3465) <= '1';
    layer6_outputs(3466) <= not a;
    layer6_outputs(3467) <= not (a and b);
    layer6_outputs(3468) <= a or b;
    layer6_outputs(3469) <= b;
    layer6_outputs(3470) <= b and not a;
    layer6_outputs(3471) <= not a;
    layer6_outputs(3472) <= not a;
    layer6_outputs(3473) <= not b;
    layer6_outputs(3474) <= not b;
    layer6_outputs(3475) <= a or b;
    layer6_outputs(3476) <= not (a xor b);
    layer6_outputs(3477) <= a;
    layer6_outputs(3478) <= a xor b;
    layer6_outputs(3479) <= b;
    layer6_outputs(3480) <= not (a xor b);
    layer6_outputs(3481) <= not (a and b);
    layer6_outputs(3482) <= a;
    layer6_outputs(3483) <= a xor b;
    layer6_outputs(3484) <= not a;
    layer6_outputs(3485) <= not a;
    layer6_outputs(3486) <= not b;
    layer6_outputs(3487) <= '0';
    layer6_outputs(3488) <= not b;
    layer6_outputs(3489) <= a or b;
    layer6_outputs(3490) <= not a;
    layer6_outputs(3491) <= not b;
    layer6_outputs(3492) <= not a;
    layer6_outputs(3493) <= b;
    layer6_outputs(3494) <= b and not a;
    layer6_outputs(3495) <= not b or a;
    layer6_outputs(3496) <= not b;
    layer6_outputs(3497) <= a;
    layer6_outputs(3498) <= a;
    layer6_outputs(3499) <= a;
    layer6_outputs(3500) <= b;
    layer6_outputs(3501) <= a;
    layer6_outputs(3502) <= b;
    layer6_outputs(3503) <= not (a xor b);
    layer6_outputs(3504) <= not b;
    layer6_outputs(3505) <= a;
    layer6_outputs(3506) <= b;
    layer6_outputs(3507) <= a;
    layer6_outputs(3508) <= a or b;
    layer6_outputs(3509) <= b and not a;
    layer6_outputs(3510) <= not (a or b);
    layer6_outputs(3511) <= a or b;
    layer6_outputs(3512) <= not (a and b);
    layer6_outputs(3513) <= a and not b;
    layer6_outputs(3514) <= not (a or b);
    layer6_outputs(3515) <= b;
    layer6_outputs(3516) <= not b or a;
    layer6_outputs(3517) <= a or b;
    layer6_outputs(3518) <= not (a or b);
    layer6_outputs(3519) <= not b or a;
    layer6_outputs(3520) <= a and not b;
    layer6_outputs(3521) <= not a;
    layer6_outputs(3522) <= not b;
    layer6_outputs(3523) <= b and not a;
    layer6_outputs(3524) <= not b;
    layer6_outputs(3525) <= not (a and b);
    layer6_outputs(3526) <= a and not b;
    layer6_outputs(3527) <= a;
    layer6_outputs(3528) <= a;
    layer6_outputs(3529) <= a and not b;
    layer6_outputs(3530) <= a xor b;
    layer6_outputs(3531) <= '1';
    layer6_outputs(3532) <= not b or a;
    layer6_outputs(3533) <= not b or a;
    layer6_outputs(3534) <= not b;
    layer6_outputs(3535) <= a and not b;
    layer6_outputs(3536) <= not (a xor b);
    layer6_outputs(3537) <= a and not b;
    layer6_outputs(3538) <= not a or b;
    layer6_outputs(3539) <= not a;
    layer6_outputs(3540) <= a and not b;
    layer6_outputs(3541) <= not a or b;
    layer6_outputs(3542) <= not a;
    layer6_outputs(3543) <= b;
    layer6_outputs(3544) <= not b;
    layer6_outputs(3545) <= b and not a;
    layer6_outputs(3546) <= not a or b;
    layer6_outputs(3547) <= b;
    layer6_outputs(3548) <= b;
    layer6_outputs(3549) <= a xor b;
    layer6_outputs(3550) <= b;
    layer6_outputs(3551) <= not a;
    layer6_outputs(3552) <= not (a xor b);
    layer6_outputs(3553) <= a;
    layer6_outputs(3554) <= not (a or b);
    layer6_outputs(3555) <= not (a xor b);
    layer6_outputs(3556) <= not b or a;
    layer6_outputs(3557) <= a and b;
    layer6_outputs(3558) <= not b;
    layer6_outputs(3559) <= not (a or b);
    layer6_outputs(3560) <= not (a or b);
    layer6_outputs(3561) <= not b;
    layer6_outputs(3562) <= a and not b;
    layer6_outputs(3563) <= b;
    layer6_outputs(3564) <= not a or b;
    layer6_outputs(3565) <= not b;
    layer6_outputs(3566) <= not b or a;
    layer6_outputs(3567) <= a;
    layer6_outputs(3568) <= a and not b;
    layer6_outputs(3569) <= not b;
    layer6_outputs(3570) <= not (a or b);
    layer6_outputs(3571) <= b and not a;
    layer6_outputs(3572) <= not (a or b);
    layer6_outputs(3573) <= not b or a;
    layer6_outputs(3574) <= not (a xor b);
    layer6_outputs(3575) <= not (a xor b);
    layer6_outputs(3576) <= a or b;
    layer6_outputs(3577) <= not b or a;
    layer6_outputs(3578) <= a and b;
    layer6_outputs(3579) <= a and not b;
    layer6_outputs(3580) <= '0';
    layer6_outputs(3581) <= not b;
    layer6_outputs(3582) <= not (a or b);
    layer6_outputs(3583) <= b;
    layer6_outputs(3584) <= not b;
    layer6_outputs(3585) <= a;
    layer6_outputs(3586) <= a or b;
    layer6_outputs(3587) <= not (a or b);
    layer6_outputs(3588) <= not a;
    layer6_outputs(3589) <= '1';
    layer6_outputs(3590) <= a or b;
    layer6_outputs(3591) <= not (a and b);
    layer6_outputs(3592) <= not (a xor b);
    layer6_outputs(3593) <= not a or b;
    layer6_outputs(3594) <= not (a and b);
    layer6_outputs(3595) <= not a;
    layer6_outputs(3596) <= not (a or b);
    layer6_outputs(3597) <= a or b;
    layer6_outputs(3598) <= not a;
    layer6_outputs(3599) <= not a or b;
    layer6_outputs(3600) <= a or b;
    layer6_outputs(3601) <= not b or a;
    layer6_outputs(3602) <= not a;
    layer6_outputs(3603) <= b;
    layer6_outputs(3604) <= a;
    layer6_outputs(3605) <= a and b;
    layer6_outputs(3606) <= not (a and b);
    layer6_outputs(3607) <= a xor b;
    layer6_outputs(3608) <= not (a and b);
    layer6_outputs(3609) <= b and not a;
    layer6_outputs(3610) <= b;
    layer6_outputs(3611) <= a and b;
    layer6_outputs(3612) <= not (a xor b);
    layer6_outputs(3613) <= b and not a;
    layer6_outputs(3614) <= b;
    layer6_outputs(3615) <= b;
    layer6_outputs(3616) <= not a or b;
    layer6_outputs(3617) <= b and not a;
    layer6_outputs(3618) <= not a;
    layer6_outputs(3619) <= b;
    layer6_outputs(3620) <= not (a xor b);
    layer6_outputs(3621) <= not b;
    layer6_outputs(3622) <= not (a xor b);
    layer6_outputs(3623) <= a xor b;
    layer6_outputs(3624) <= not b;
    layer6_outputs(3625) <= not a or b;
    layer6_outputs(3626) <= not a or b;
    layer6_outputs(3627) <= a and not b;
    layer6_outputs(3628) <= a or b;
    layer6_outputs(3629) <= not b;
    layer6_outputs(3630) <= a;
    layer6_outputs(3631) <= a and b;
    layer6_outputs(3632) <= not (a or b);
    layer6_outputs(3633) <= a;
    layer6_outputs(3634) <= not a;
    layer6_outputs(3635) <= not (a xor b);
    layer6_outputs(3636) <= not (a and b);
    layer6_outputs(3637) <= not a;
    layer6_outputs(3638) <= not a;
    layer6_outputs(3639) <= a and b;
    layer6_outputs(3640) <= not a or b;
    layer6_outputs(3641) <= not b;
    layer6_outputs(3642) <= not b;
    layer6_outputs(3643) <= not (a xor b);
    layer6_outputs(3644) <= b;
    layer6_outputs(3645) <= a;
    layer6_outputs(3646) <= not (a or b);
    layer6_outputs(3647) <= a and b;
    layer6_outputs(3648) <= b;
    layer6_outputs(3649) <= '1';
    layer6_outputs(3650) <= not a;
    layer6_outputs(3651) <= a xor b;
    layer6_outputs(3652) <= a;
    layer6_outputs(3653) <= a and b;
    layer6_outputs(3654) <= not (a and b);
    layer6_outputs(3655) <= not (a and b);
    layer6_outputs(3656) <= not a or b;
    layer6_outputs(3657) <= a and not b;
    layer6_outputs(3658) <= a and not b;
    layer6_outputs(3659) <= b;
    layer6_outputs(3660) <= a or b;
    layer6_outputs(3661) <= not b or a;
    layer6_outputs(3662) <= a and not b;
    layer6_outputs(3663) <= not a;
    layer6_outputs(3664) <= a and not b;
    layer6_outputs(3665) <= a;
    layer6_outputs(3666) <= not a;
    layer6_outputs(3667) <= not (a or b);
    layer6_outputs(3668) <= a;
    layer6_outputs(3669) <= not (a or b);
    layer6_outputs(3670) <= not (a and b);
    layer6_outputs(3671) <= b;
    layer6_outputs(3672) <= '1';
    layer6_outputs(3673) <= '0';
    layer6_outputs(3674) <= not a or b;
    layer6_outputs(3675) <= b;
    layer6_outputs(3676) <= not a;
    layer6_outputs(3677) <= a xor b;
    layer6_outputs(3678) <= a;
    layer6_outputs(3679) <= not a;
    layer6_outputs(3680) <= not (a xor b);
    layer6_outputs(3681) <= not a or b;
    layer6_outputs(3682) <= b;
    layer6_outputs(3683) <= not a;
    layer6_outputs(3684) <= b and not a;
    layer6_outputs(3685) <= a and b;
    layer6_outputs(3686) <= b and not a;
    layer6_outputs(3687) <= a;
    layer6_outputs(3688) <= not b or a;
    layer6_outputs(3689) <= b and not a;
    layer6_outputs(3690) <= a and b;
    layer6_outputs(3691) <= not a or b;
    layer6_outputs(3692) <= not b or a;
    layer6_outputs(3693) <= a and not b;
    layer6_outputs(3694) <= '0';
    layer6_outputs(3695) <= a and not b;
    layer6_outputs(3696) <= a;
    layer6_outputs(3697) <= '1';
    layer6_outputs(3698) <= a xor b;
    layer6_outputs(3699) <= b and not a;
    layer6_outputs(3700) <= not (a or b);
    layer6_outputs(3701) <= not (a or b);
    layer6_outputs(3702) <= not (a or b);
    layer6_outputs(3703) <= b and not a;
    layer6_outputs(3704) <= not b;
    layer6_outputs(3705) <= a xor b;
    layer6_outputs(3706) <= not b or a;
    layer6_outputs(3707) <= not b;
    layer6_outputs(3708) <= not (a xor b);
    layer6_outputs(3709) <= a;
    layer6_outputs(3710) <= a;
    layer6_outputs(3711) <= b;
    layer6_outputs(3712) <= not b or a;
    layer6_outputs(3713) <= a xor b;
    layer6_outputs(3714) <= not a or b;
    layer6_outputs(3715) <= a;
    layer6_outputs(3716) <= a;
    layer6_outputs(3717) <= a and b;
    layer6_outputs(3718) <= not a;
    layer6_outputs(3719) <= not b;
    layer6_outputs(3720) <= b and not a;
    layer6_outputs(3721) <= b and not a;
    layer6_outputs(3722) <= not b or a;
    layer6_outputs(3723) <= b and not a;
    layer6_outputs(3724) <= not b or a;
    layer6_outputs(3725) <= not a;
    layer6_outputs(3726) <= b and not a;
    layer6_outputs(3727) <= not (a and b);
    layer6_outputs(3728) <= not b or a;
    layer6_outputs(3729) <= not b;
    layer6_outputs(3730) <= a;
    layer6_outputs(3731) <= not b;
    layer6_outputs(3732) <= not (a xor b);
    layer6_outputs(3733) <= not (a and b);
    layer6_outputs(3734) <= not a;
    layer6_outputs(3735) <= a or b;
    layer6_outputs(3736) <= not b;
    layer6_outputs(3737) <= not (a and b);
    layer6_outputs(3738) <= a and b;
    layer6_outputs(3739) <= b and not a;
    layer6_outputs(3740) <= a and not b;
    layer6_outputs(3741) <= a;
    layer6_outputs(3742) <= not a;
    layer6_outputs(3743) <= a and not b;
    layer6_outputs(3744) <= not a;
    layer6_outputs(3745) <= not (a and b);
    layer6_outputs(3746) <= b;
    layer6_outputs(3747) <= a or b;
    layer6_outputs(3748) <= not a;
    layer6_outputs(3749) <= b;
    layer6_outputs(3750) <= not a;
    layer6_outputs(3751) <= not (a or b);
    layer6_outputs(3752) <= a xor b;
    layer6_outputs(3753) <= a;
    layer6_outputs(3754) <= a and b;
    layer6_outputs(3755) <= not a or b;
    layer6_outputs(3756) <= a and b;
    layer6_outputs(3757) <= a and not b;
    layer6_outputs(3758) <= not (a xor b);
    layer6_outputs(3759) <= a and b;
    layer6_outputs(3760) <= '1';
    layer6_outputs(3761) <= not a or b;
    layer6_outputs(3762) <= a xor b;
    layer6_outputs(3763) <= '1';
    layer6_outputs(3764) <= a and b;
    layer6_outputs(3765) <= a and b;
    layer6_outputs(3766) <= not (a xor b);
    layer6_outputs(3767) <= not a or b;
    layer6_outputs(3768) <= not (a or b);
    layer6_outputs(3769) <= a or b;
    layer6_outputs(3770) <= a or b;
    layer6_outputs(3771) <= not (a xor b);
    layer6_outputs(3772) <= not b or a;
    layer6_outputs(3773) <= b;
    layer6_outputs(3774) <= a and not b;
    layer6_outputs(3775) <= b and not a;
    layer6_outputs(3776) <= b;
    layer6_outputs(3777) <= a and not b;
    layer6_outputs(3778) <= b;
    layer6_outputs(3779) <= a or b;
    layer6_outputs(3780) <= b;
    layer6_outputs(3781) <= not b or a;
    layer6_outputs(3782) <= not (a and b);
    layer6_outputs(3783) <= a;
    layer6_outputs(3784) <= not a;
    layer6_outputs(3785) <= b and not a;
    layer6_outputs(3786) <= a and b;
    layer6_outputs(3787) <= not a;
    layer6_outputs(3788) <= not b;
    layer6_outputs(3789) <= a and not b;
    layer6_outputs(3790) <= a or b;
    layer6_outputs(3791) <= b;
    layer6_outputs(3792) <= not (a or b);
    layer6_outputs(3793) <= a or b;
    layer6_outputs(3794) <= a or b;
    layer6_outputs(3795) <= not b or a;
    layer6_outputs(3796) <= not a;
    layer6_outputs(3797) <= b;
    layer6_outputs(3798) <= a;
    layer6_outputs(3799) <= not a or b;
    layer6_outputs(3800) <= not b or a;
    layer6_outputs(3801) <= a and b;
    layer6_outputs(3802) <= not a or b;
    layer6_outputs(3803) <= a;
    layer6_outputs(3804) <= a or b;
    layer6_outputs(3805) <= not a;
    layer6_outputs(3806) <= a xor b;
    layer6_outputs(3807) <= not a or b;
    layer6_outputs(3808) <= not (a and b);
    layer6_outputs(3809) <= b;
    layer6_outputs(3810) <= a or b;
    layer6_outputs(3811) <= not a;
    layer6_outputs(3812) <= not b;
    layer6_outputs(3813) <= not b;
    layer6_outputs(3814) <= a;
    layer6_outputs(3815) <= not a or b;
    layer6_outputs(3816) <= a;
    layer6_outputs(3817) <= a or b;
    layer6_outputs(3818) <= not (a or b);
    layer6_outputs(3819) <= a and not b;
    layer6_outputs(3820) <= not b;
    layer6_outputs(3821) <= a xor b;
    layer6_outputs(3822) <= not a or b;
    layer6_outputs(3823) <= a;
    layer6_outputs(3824) <= not (a or b);
    layer6_outputs(3825) <= b;
    layer6_outputs(3826) <= '1';
    layer6_outputs(3827) <= b and not a;
    layer6_outputs(3828) <= not a;
    layer6_outputs(3829) <= a and not b;
    layer6_outputs(3830) <= not b;
    layer6_outputs(3831) <= a xor b;
    layer6_outputs(3832) <= not b or a;
    layer6_outputs(3833) <= a or b;
    layer6_outputs(3834) <= '0';
    layer6_outputs(3835) <= a and not b;
    layer6_outputs(3836) <= not (a xor b);
    layer6_outputs(3837) <= not (a or b);
    layer6_outputs(3838) <= a and b;
    layer6_outputs(3839) <= not a;
    layer6_outputs(3840) <= '1';
    layer6_outputs(3841) <= not a or b;
    layer6_outputs(3842) <= not b or a;
    layer6_outputs(3843) <= a and not b;
    layer6_outputs(3844) <= not b;
    layer6_outputs(3845) <= not a;
    layer6_outputs(3846) <= not b;
    layer6_outputs(3847) <= a;
    layer6_outputs(3848) <= a and b;
    layer6_outputs(3849) <= a;
    layer6_outputs(3850) <= not a;
    layer6_outputs(3851) <= a;
    layer6_outputs(3852) <= a or b;
    layer6_outputs(3853) <= a and b;
    layer6_outputs(3854) <= not b or a;
    layer6_outputs(3855) <= not a;
    layer6_outputs(3856) <= not (a and b);
    layer6_outputs(3857) <= not a or b;
    layer6_outputs(3858) <= b;
    layer6_outputs(3859) <= a and b;
    layer6_outputs(3860) <= not b or a;
    layer6_outputs(3861) <= b;
    layer6_outputs(3862) <= a or b;
    layer6_outputs(3863) <= b and not a;
    layer6_outputs(3864) <= b and not a;
    layer6_outputs(3865) <= not b;
    layer6_outputs(3866) <= a and b;
    layer6_outputs(3867) <= a and b;
    layer6_outputs(3868) <= a xor b;
    layer6_outputs(3869) <= b and not a;
    layer6_outputs(3870) <= a or b;
    layer6_outputs(3871) <= not (a or b);
    layer6_outputs(3872) <= not (a or b);
    layer6_outputs(3873) <= b and not a;
    layer6_outputs(3874) <= not (a or b);
    layer6_outputs(3875) <= a and b;
    layer6_outputs(3876) <= '1';
    layer6_outputs(3877) <= not b or a;
    layer6_outputs(3878) <= not b or a;
    layer6_outputs(3879) <= a xor b;
    layer6_outputs(3880) <= a xor b;
    layer6_outputs(3881) <= not a;
    layer6_outputs(3882) <= not b or a;
    layer6_outputs(3883) <= not b or a;
    layer6_outputs(3884) <= not (a xor b);
    layer6_outputs(3885) <= not b;
    layer6_outputs(3886) <= a;
    layer6_outputs(3887) <= not (a and b);
    layer6_outputs(3888) <= not a;
    layer6_outputs(3889) <= not (a or b);
    layer6_outputs(3890) <= not a;
    layer6_outputs(3891) <= a or b;
    layer6_outputs(3892) <= not b;
    layer6_outputs(3893) <= a and b;
    layer6_outputs(3894) <= a and b;
    layer6_outputs(3895) <= not b;
    layer6_outputs(3896) <= not a;
    layer6_outputs(3897) <= a and not b;
    layer6_outputs(3898) <= not b;
    layer6_outputs(3899) <= not b or a;
    layer6_outputs(3900) <= a or b;
    layer6_outputs(3901) <= b;
    layer6_outputs(3902) <= not a or b;
    layer6_outputs(3903) <= a and not b;
    layer6_outputs(3904) <= not a or b;
    layer6_outputs(3905) <= a xor b;
    layer6_outputs(3906) <= a or b;
    layer6_outputs(3907) <= a;
    layer6_outputs(3908) <= b and not a;
    layer6_outputs(3909) <= not b;
    layer6_outputs(3910) <= not a;
    layer6_outputs(3911) <= b;
    layer6_outputs(3912) <= not b;
    layer6_outputs(3913) <= b and not a;
    layer6_outputs(3914) <= a;
    layer6_outputs(3915) <= not b;
    layer6_outputs(3916) <= not b;
    layer6_outputs(3917) <= not (a or b);
    layer6_outputs(3918) <= b;
    layer6_outputs(3919) <= not a or b;
    layer6_outputs(3920) <= b;
    layer6_outputs(3921) <= '0';
    layer6_outputs(3922) <= a xor b;
    layer6_outputs(3923) <= not (a and b);
    layer6_outputs(3924) <= '0';
    layer6_outputs(3925) <= a or b;
    layer6_outputs(3926) <= a;
    layer6_outputs(3927) <= not (a and b);
    layer6_outputs(3928) <= a xor b;
    layer6_outputs(3929) <= not b;
    layer6_outputs(3930) <= not a;
    layer6_outputs(3931) <= not (a and b);
    layer6_outputs(3932) <= a and not b;
    layer6_outputs(3933) <= a and not b;
    layer6_outputs(3934) <= not (a and b);
    layer6_outputs(3935) <= not (a or b);
    layer6_outputs(3936) <= a and not b;
    layer6_outputs(3937) <= a;
    layer6_outputs(3938) <= a;
    layer6_outputs(3939) <= not a;
    layer6_outputs(3940) <= not b or a;
    layer6_outputs(3941) <= b and not a;
    layer6_outputs(3942) <= a and not b;
    layer6_outputs(3943) <= not (a and b);
    layer6_outputs(3944) <= a;
    layer6_outputs(3945) <= not b;
    layer6_outputs(3946) <= b;
    layer6_outputs(3947) <= a and b;
    layer6_outputs(3948) <= not (a and b);
    layer6_outputs(3949) <= a or b;
    layer6_outputs(3950) <= a xor b;
    layer6_outputs(3951) <= not (a and b);
    layer6_outputs(3952) <= a and b;
    layer6_outputs(3953) <= not (a and b);
    layer6_outputs(3954) <= '0';
    layer6_outputs(3955) <= not a;
    layer6_outputs(3956) <= not b;
    layer6_outputs(3957) <= a xor b;
    layer6_outputs(3958) <= not b or a;
    layer6_outputs(3959) <= not b;
    layer6_outputs(3960) <= not (a xor b);
    layer6_outputs(3961) <= not a;
    layer6_outputs(3962) <= not a;
    layer6_outputs(3963) <= a or b;
    layer6_outputs(3964) <= b;
    layer6_outputs(3965) <= a xor b;
    layer6_outputs(3966) <= a and b;
    layer6_outputs(3967) <= not a;
    layer6_outputs(3968) <= not (a xor b);
    layer6_outputs(3969) <= a;
    layer6_outputs(3970) <= a and not b;
    layer6_outputs(3971) <= not b or a;
    layer6_outputs(3972) <= b;
    layer6_outputs(3973) <= not a or b;
    layer6_outputs(3974) <= not (a and b);
    layer6_outputs(3975) <= not (a and b);
    layer6_outputs(3976) <= not (a and b);
    layer6_outputs(3977) <= a and not b;
    layer6_outputs(3978) <= b;
    layer6_outputs(3979) <= not b or a;
    layer6_outputs(3980) <= a or b;
    layer6_outputs(3981) <= a or b;
    layer6_outputs(3982) <= a and b;
    layer6_outputs(3983) <= not b;
    layer6_outputs(3984) <= a;
    layer6_outputs(3985) <= b and not a;
    layer6_outputs(3986) <= a and not b;
    layer6_outputs(3987) <= a and b;
    layer6_outputs(3988) <= a;
    layer6_outputs(3989) <= not b;
    layer6_outputs(3990) <= a and b;
    layer6_outputs(3991) <= not b or a;
    layer6_outputs(3992) <= not b;
    layer6_outputs(3993) <= not a;
    layer6_outputs(3994) <= '0';
    layer6_outputs(3995) <= a xor b;
    layer6_outputs(3996) <= not b or a;
    layer6_outputs(3997) <= not a or b;
    layer6_outputs(3998) <= b and not a;
    layer6_outputs(3999) <= not a;
    layer6_outputs(4000) <= not b or a;
    layer6_outputs(4001) <= not (a and b);
    layer6_outputs(4002) <= b;
    layer6_outputs(4003) <= not b;
    layer6_outputs(4004) <= not b or a;
    layer6_outputs(4005) <= not b or a;
    layer6_outputs(4006) <= '1';
    layer6_outputs(4007) <= a;
    layer6_outputs(4008) <= '0';
    layer6_outputs(4009) <= not (a and b);
    layer6_outputs(4010) <= a or b;
    layer6_outputs(4011) <= a;
    layer6_outputs(4012) <= a and b;
    layer6_outputs(4013) <= not a;
    layer6_outputs(4014) <= b and not a;
    layer6_outputs(4015) <= b;
    layer6_outputs(4016) <= '0';
    layer6_outputs(4017) <= not (a or b);
    layer6_outputs(4018) <= a or b;
    layer6_outputs(4019) <= a;
    layer6_outputs(4020) <= not a;
    layer6_outputs(4021) <= not b or a;
    layer6_outputs(4022) <= b;
    layer6_outputs(4023) <= not (a xor b);
    layer6_outputs(4024) <= a;
    layer6_outputs(4025) <= not b;
    layer6_outputs(4026) <= a;
    layer6_outputs(4027) <= not a;
    layer6_outputs(4028) <= not b or a;
    layer6_outputs(4029) <= a;
    layer6_outputs(4030) <= b and not a;
    layer6_outputs(4031) <= not b;
    layer6_outputs(4032) <= not b;
    layer6_outputs(4033) <= a;
    layer6_outputs(4034) <= a xor b;
    layer6_outputs(4035) <= '0';
    layer6_outputs(4036) <= not a;
    layer6_outputs(4037) <= not a or b;
    layer6_outputs(4038) <= not (a and b);
    layer6_outputs(4039) <= a;
    layer6_outputs(4040) <= '1';
    layer6_outputs(4041) <= b and not a;
    layer6_outputs(4042) <= b and not a;
    layer6_outputs(4043) <= not (a or b);
    layer6_outputs(4044) <= not (a xor b);
    layer6_outputs(4045) <= a and not b;
    layer6_outputs(4046) <= b;
    layer6_outputs(4047) <= not a;
    layer6_outputs(4048) <= a;
    layer6_outputs(4049) <= not b;
    layer6_outputs(4050) <= not b or a;
    layer6_outputs(4051) <= not a;
    layer6_outputs(4052) <= a;
    layer6_outputs(4053) <= not a;
    layer6_outputs(4054) <= b;
    layer6_outputs(4055) <= a and not b;
    layer6_outputs(4056) <= b;
    layer6_outputs(4057) <= b;
    layer6_outputs(4058) <= not a;
    layer6_outputs(4059) <= not b or a;
    layer6_outputs(4060) <= not b;
    layer6_outputs(4061) <= not (a and b);
    layer6_outputs(4062) <= not a;
    layer6_outputs(4063) <= not a;
    layer6_outputs(4064) <= not a;
    layer6_outputs(4065) <= a and b;
    layer6_outputs(4066) <= b;
    layer6_outputs(4067) <= not (a and b);
    layer6_outputs(4068) <= a xor b;
    layer6_outputs(4069) <= b;
    layer6_outputs(4070) <= not b;
    layer6_outputs(4071) <= a or b;
    layer6_outputs(4072) <= a and b;
    layer6_outputs(4073) <= a;
    layer6_outputs(4074) <= not a or b;
    layer6_outputs(4075) <= not (a or b);
    layer6_outputs(4076) <= b;
    layer6_outputs(4077) <= not (a xor b);
    layer6_outputs(4078) <= not (a and b);
    layer6_outputs(4079) <= not (a and b);
    layer6_outputs(4080) <= a or b;
    layer6_outputs(4081) <= b;
    layer6_outputs(4082) <= b;
    layer6_outputs(4083) <= not (a or b);
    layer6_outputs(4084) <= a and b;
    layer6_outputs(4085) <= a and b;
    layer6_outputs(4086) <= not a;
    layer6_outputs(4087) <= b;
    layer6_outputs(4088) <= a and not b;
    layer6_outputs(4089) <= not b or a;
    layer6_outputs(4090) <= b;
    layer6_outputs(4091) <= not a or b;
    layer6_outputs(4092) <= b;
    layer6_outputs(4093) <= not (a or b);
    layer6_outputs(4094) <= a and not b;
    layer6_outputs(4095) <= not (a and b);
    layer6_outputs(4096) <= a or b;
    layer6_outputs(4097) <= a xor b;
    layer6_outputs(4098) <= not a;
    layer6_outputs(4099) <= not (a and b);
    layer6_outputs(4100) <= not b;
    layer6_outputs(4101) <= a or b;
    layer6_outputs(4102) <= not b;
    layer6_outputs(4103) <= not a;
    layer6_outputs(4104) <= not (a or b);
    layer6_outputs(4105) <= not (a or b);
    layer6_outputs(4106) <= a;
    layer6_outputs(4107) <= not (a xor b);
    layer6_outputs(4108) <= a xor b;
    layer6_outputs(4109) <= not (a or b);
    layer6_outputs(4110) <= not a;
    layer6_outputs(4111) <= not (a or b);
    layer6_outputs(4112) <= a or b;
    layer6_outputs(4113) <= a;
    layer6_outputs(4114) <= not b;
    layer6_outputs(4115) <= not b;
    layer6_outputs(4116) <= not a;
    layer6_outputs(4117) <= not a;
    layer6_outputs(4118) <= a xor b;
    layer6_outputs(4119) <= not (a xor b);
    layer6_outputs(4120) <= not (a or b);
    layer6_outputs(4121) <= a or b;
    layer6_outputs(4122) <= a and b;
    layer6_outputs(4123) <= not (a and b);
    layer6_outputs(4124) <= not a;
    layer6_outputs(4125) <= not b or a;
    layer6_outputs(4126) <= not b or a;
    layer6_outputs(4127) <= a or b;
    layer6_outputs(4128) <= not a;
    layer6_outputs(4129) <= b;
    layer6_outputs(4130) <= b and not a;
    layer6_outputs(4131) <= not a;
    layer6_outputs(4132) <= a and b;
    layer6_outputs(4133) <= not b;
    layer6_outputs(4134) <= not b;
    layer6_outputs(4135) <= not a;
    layer6_outputs(4136) <= b;
    layer6_outputs(4137) <= a;
    layer6_outputs(4138) <= a xor b;
    layer6_outputs(4139) <= not a or b;
    layer6_outputs(4140) <= b and not a;
    layer6_outputs(4141) <= b and not a;
    layer6_outputs(4142) <= not a or b;
    layer6_outputs(4143) <= not a;
    layer6_outputs(4144) <= b;
    layer6_outputs(4145) <= not b or a;
    layer6_outputs(4146) <= not b or a;
    layer6_outputs(4147) <= a;
    layer6_outputs(4148) <= a xor b;
    layer6_outputs(4149) <= not a;
    layer6_outputs(4150) <= not (a or b);
    layer6_outputs(4151) <= a and b;
    layer6_outputs(4152) <= not b;
    layer6_outputs(4153) <= '0';
    layer6_outputs(4154) <= '1';
    layer6_outputs(4155) <= not a;
    layer6_outputs(4156) <= a and b;
    layer6_outputs(4157) <= b and not a;
    layer6_outputs(4158) <= b;
    layer6_outputs(4159) <= b;
    layer6_outputs(4160) <= a and not b;
    layer6_outputs(4161) <= a;
    layer6_outputs(4162) <= not a;
    layer6_outputs(4163) <= not b;
    layer6_outputs(4164) <= a;
    layer6_outputs(4165) <= not (a and b);
    layer6_outputs(4166) <= not (a or b);
    layer6_outputs(4167) <= not (a or b);
    layer6_outputs(4168) <= not (a and b);
    layer6_outputs(4169) <= not (a and b);
    layer6_outputs(4170) <= b and not a;
    layer6_outputs(4171) <= a xor b;
    layer6_outputs(4172) <= a;
    layer6_outputs(4173) <= not b or a;
    layer6_outputs(4174) <= not (a or b);
    layer6_outputs(4175) <= not a;
    layer6_outputs(4176) <= not (a and b);
    layer6_outputs(4177) <= not a;
    layer6_outputs(4178) <= a or b;
    layer6_outputs(4179) <= not (a or b);
    layer6_outputs(4180) <= b and not a;
    layer6_outputs(4181) <= not (a or b);
    layer6_outputs(4182) <= not b or a;
    layer6_outputs(4183) <= b;
    layer6_outputs(4184) <= a xor b;
    layer6_outputs(4185) <= a and not b;
    layer6_outputs(4186) <= a xor b;
    layer6_outputs(4187) <= b;
    layer6_outputs(4188) <= a or b;
    layer6_outputs(4189) <= a or b;
    layer6_outputs(4190) <= not (a or b);
    layer6_outputs(4191) <= b;
    layer6_outputs(4192) <= not a;
    layer6_outputs(4193) <= not b;
    layer6_outputs(4194) <= not b;
    layer6_outputs(4195) <= not (a xor b);
    layer6_outputs(4196) <= a or b;
    layer6_outputs(4197) <= not a or b;
    layer6_outputs(4198) <= not a;
    layer6_outputs(4199) <= not b;
    layer6_outputs(4200) <= a;
    layer6_outputs(4201) <= not (a or b);
    layer6_outputs(4202) <= a and b;
    layer6_outputs(4203) <= a and not b;
    layer6_outputs(4204) <= a and b;
    layer6_outputs(4205) <= a and b;
    layer6_outputs(4206) <= not (a or b);
    layer6_outputs(4207) <= not a;
    layer6_outputs(4208) <= not a;
    layer6_outputs(4209) <= '0';
    layer6_outputs(4210) <= a and b;
    layer6_outputs(4211) <= a and not b;
    layer6_outputs(4212) <= a and b;
    layer6_outputs(4213) <= not (a xor b);
    layer6_outputs(4214) <= a;
    layer6_outputs(4215) <= not a;
    layer6_outputs(4216) <= not (a or b);
    layer6_outputs(4217) <= not a;
    layer6_outputs(4218) <= not (a xor b);
    layer6_outputs(4219) <= not (a or b);
    layer6_outputs(4220) <= not (a xor b);
    layer6_outputs(4221) <= a;
    layer6_outputs(4222) <= a xor b;
    layer6_outputs(4223) <= not b or a;
    layer6_outputs(4224) <= b and not a;
    layer6_outputs(4225) <= a and not b;
    layer6_outputs(4226) <= not b;
    layer6_outputs(4227) <= not b;
    layer6_outputs(4228) <= not a;
    layer6_outputs(4229) <= not (a or b);
    layer6_outputs(4230) <= b;
    layer6_outputs(4231) <= not b;
    layer6_outputs(4232) <= '1';
    layer6_outputs(4233) <= a;
    layer6_outputs(4234) <= not b or a;
    layer6_outputs(4235) <= not a;
    layer6_outputs(4236) <= not (a xor b);
    layer6_outputs(4237) <= not a;
    layer6_outputs(4238) <= a;
    layer6_outputs(4239) <= b;
    layer6_outputs(4240) <= a;
    layer6_outputs(4241) <= not b or a;
    layer6_outputs(4242) <= not (a and b);
    layer6_outputs(4243) <= b;
    layer6_outputs(4244) <= not a or b;
    layer6_outputs(4245) <= not (a xor b);
    layer6_outputs(4246) <= a or b;
    layer6_outputs(4247) <= a xor b;
    layer6_outputs(4248) <= b and not a;
    layer6_outputs(4249) <= a;
    layer6_outputs(4250) <= a xor b;
    layer6_outputs(4251) <= not b;
    layer6_outputs(4252) <= not a;
    layer6_outputs(4253) <= not (a xor b);
    layer6_outputs(4254) <= not a;
    layer6_outputs(4255) <= a and b;
    layer6_outputs(4256) <= not a;
    layer6_outputs(4257) <= b;
    layer6_outputs(4258) <= not (a and b);
    layer6_outputs(4259) <= not (a xor b);
    layer6_outputs(4260) <= a;
    layer6_outputs(4261) <= not a;
    layer6_outputs(4262) <= a xor b;
    layer6_outputs(4263) <= a or b;
    layer6_outputs(4264) <= not (a xor b);
    layer6_outputs(4265) <= a and not b;
    layer6_outputs(4266) <= not b or a;
    layer6_outputs(4267) <= not b or a;
    layer6_outputs(4268) <= a;
    layer6_outputs(4269) <= not (a or b);
    layer6_outputs(4270) <= not a;
    layer6_outputs(4271) <= not (a and b);
    layer6_outputs(4272) <= not a;
    layer6_outputs(4273) <= not a;
    layer6_outputs(4274) <= b and not a;
    layer6_outputs(4275) <= not b or a;
    layer6_outputs(4276) <= a and b;
    layer6_outputs(4277) <= a or b;
    layer6_outputs(4278) <= b;
    layer6_outputs(4279) <= b;
    layer6_outputs(4280) <= b;
    layer6_outputs(4281) <= b;
    layer6_outputs(4282) <= a or b;
    layer6_outputs(4283) <= not a or b;
    layer6_outputs(4284) <= a or b;
    layer6_outputs(4285) <= not (a and b);
    layer6_outputs(4286) <= a;
    layer6_outputs(4287) <= a and b;
    layer6_outputs(4288) <= not b;
    layer6_outputs(4289) <= b;
    layer6_outputs(4290) <= a and b;
    layer6_outputs(4291) <= not (a or b);
    layer6_outputs(4292) <= not b;
    layer6_outputs(4293) <= not (a or b);
    layer6_outputs(4294) <= a and b;
    layer6_outputs(4295) <= not a;
    layer6_outputs(4296) <= not (a or b);
    layer6_outputs(4297) <= a;
    layer6_outputs(4298) <= not b;
    layer6_outputs(4299) <= b;
    layer6_outputs(4300) <= not b;
    layer6_outputs(4301) <= not (a and b);
    layer6_outputs(4302) <= not a;
    layer6_outputs(4303) <= not b;
    layer6_outputs(4304) <= a xor b;
    layer6_outputs(4305) <= a and not b;
    layer6_outputs(4306) <= '0';
    layer6_outputs(4307) <= b;
    layer6_outputs(4308) <= b;
    layer6_outputs(4309) <= b;
    layer6_outputs(4310) <= a and not b;
    layer6_outputs(4311) <= a xor b;
    layer6_outputs(4312) <= not a;
    layer6_outputs(4313) <= not a or b;
    layer6_outputs(4314) <= '1';
    layer6_outputs(4315) <= '0';
    layer6_outputs(4316) <= not a;
    layer6_outputs(4317) <= '0';
    layer6_outputs(4318) <= a;
    layer6_outputs(4319) <= not a;
    layer6_outputs(4320) <= a and not b;
    layer6_outputs(4321) <= not (a or b);
    layer6_outputs(4322) <= not a;
    layer6_outputs(4323) <= a and b;
    layer6_outputs(4324) <= not b or a;
    layer6_outputs(4325) <= b;
    layer6_outputs(4326) <= not b;
    layer6_outputs(4327) <= not a;
    layer6_outputs(4328) <= not a;
    layer6_outputs(4329) <= not a or b;
    layer6_outputs(4330) <= not b;
    layer6_outputs(4331) <= b;
    layer6_outputs(4332) <= not b;
    layer6_outputs(4333) <= b;
    layer6_outputs(4334) <= b;
    layer6_outputs(4335) <= not b;
    layer6_outputs(4336) <= not a or b;
    layer6_outputs(4337) <= b;
    layer6_outputs(4338) <= not b;
    layer6_outputs(4339) <= not b or a;
    layer6_outputs(4340) <= not (a or b);
    layer6_outputs(4341) <= b and not a;
    layer6_outputs(4342) <= not b;
    layer6_outputs(4343) <= '0';
    layer6_outputs(4344) <= a and b;
    layer6_outputs(4345) <= not a;
    layer6_outputs(4346) <= not (a or b);
    layer6_outputs(4347) <= a;
    layer6_outputs(4348) <= not (a or b);
    layer6_outputs(4349) <= not b or a;
    layer6_outputs(4350) <= not a or b;
    layer6_outputs(4351) <= not (a or b);
    layer6_outputs(4352) <= a and b;
    layer6_outputs(4353) <= a or b;
    layer6_outputs(4354) <= not (a or b);
    layer6_outputs(4355) <= not (a or b);
    layer6_outputs(4356) <= b;
    layer6_outputs(4357) <= a and b;
    layer6_outputs(4358) <= not (a xor b);
    layer6_outputs(4359) <= a and b;
    layer6_outputs(4360) <= b and not a;
    layer6_outputs(4361) <= not a;
    layer6_outputs(4362) <= not a;
    layer6_outputs(4363) <= b;
    layer6_outputs(4364) <= not a;
    layer6_outputs(4365) <= '0';
    layer6_outputs(4366) <= b;
    layer6_outputs(4367) <= a xor b;
    layer6_outputs(4368) <= a;
    layer6_outputs(4369) <= b and not a;
    layer6_outputs(4370) <= not b;
    layer6_outputs(4371) <= a and not b;
    layer6_outputs(4372) <= not (a or b);
    layer6_outputs(4373) <= a xor b;
    layer6_outputs(4374) <= a;
    layer6_outputs(4375) <= a or b;
    layer6_outputs(4376) <= b and not a;
    layer6_outputs(4377) <= not b or a;
    layer6_outputs(4378) <= a and b;
    layer6_outputs(4379) <= not a;
    layer6_outputs(4380) <= not b;
    layer6_outputs(4381) <= not b or a;
    layer6_outputs(4382) <= not (a xor b);
    layer6_outputs(4383) <= not b;
    layer6_outputs(4384) <= b and not a;
    layer6_outputs(4385) <= a and not b;
    layer6_outputs(4386) <= not (a and b);
    layer6_outputs(4387) <= a and not b;
    layer6_outputs(4388) <= not (a or b);
    layer6_outputs(4389) <= not (a xor b);
    layer6_outputs(4390) <= a;
    layer6_outputs(4391) <= b;
    layer6_outputs(4392) <= b;
    layer6_outputs(4393) <= b;
    layer6_outputs(4394) <= b;
    layer6_outputs(4395) <= a and not b;
    layer6_outputs(4396) <= a and b;
    layer6_outputs(4397) <= not b;
    layer6_outputs(4398) <= not b;
    layer6_outputs(4399) <= '0';
    layer6_outputs(4400) <= not a;
    layer6_outputs(4401) <= a;
    layer6_outputs(4402) <= a and not b;
    layer6_outputs(4403) <= not (a and b);
    layer6_outputs(4404) <= not a;
    layer6_outputs(4405) <= '0';
    layer6_outputs(4406) <= a xor b;
    layer6_outputs(4407) <= '1';
    layer6_outputs(4408) <= not b;
    layer6_outputs(4409) <= a and b;
    layer6_outputs(4410) <= not (a or b);
    layer6_outputs(4411) <= not b;
    layer6_outputs(4412) <= b;
    layer6_outputs(4413) <= a and b;
    layer6_outputs(4414) <= a;
    layer6_outputs(4415) <= a and b;
    layer6_outputs(4416) <= a;
    layer6_outputs(4417) <= not b or a;
    layer6_outputs(4418) <= not b or a;
    layer6_outputs(4419) <= a xor b;
    layer6_outputs(4420) <= not b;
    layer6_outputs(4421) <= not (a or b);
    layer6_outputs(4422) <= not (a or b);
    layer6_outputs(4423) <= a;
    layer6_outputs(4424) <= a or b;
    layer6_outputs(4425) <= not (a and b);
    layer6_outputs(4426) <= not b;
    layer6_outputs(4427) <= not (a or b);
    layer6_outputs(4428) <= a;
    layer6_outputs(4429) <= '0';
    layer6_outputs(4430) <= not b;
    layer6_outputs(4431) <= not b;
    layer6_outputs(4432) <= not (a and b);
    layer6_outputs(4433) <= b;
    layer6_outputs(4434) <= a xor b;
    layer6_outputs(4435) <= not a;
    layer6_outputs(4436) <= not a or b;
    layer6_outputs(4437) <= not (a and b);
    layer6_outputs(4438) <= b;
    layer6_outputs(4439) <= b;
    layer6_outputs(4440) <= a xor b;
    layer6_outputs(4441) <= b;
    layer6_outputs(4442) <= a;
    layer6_outputs(4443) <= b;
    layer6_outputs(4444) <= not (a and b);
    layer6_outputs(4445) <= a or b;
    layer6_outputs(4446) <= not b or a;
    layer6_outputs(4447) <= a;
    layer6_outputs(4448) <= not b or a;
    layer6_outputs(4449) <= not (a and b);
    layer6_outputs(4450) <= not a;
    layer6_outputs(4451) <= b;
    layer6_outputs(4452) <= '0';
    layer6_outputs(4453) <= a;
    layer6_outputs(4454) <= not (a and b);
    layer6_outputs(4455) <= b;
    layer6_outputs(4456) <= a or b;
    layer6_outputs(4457) <= a;
    layer6_outputs(4458) <= not a;
    layer6_outputs(4459) <= a;
    layer6_outputs(4460) <= b;
    layer6_outputs(4461) <= not b;
    layer6_outputs(4462) <= not (a or b);
    layer6_outputs(4463) <= not a or b;
    layer6_outputs(4464) <= a and b;
    layer6_outputs(4465) <= a;
    layer6_outputs(4466) <= a or b;
    layer6_outputs(4467) <= a or b;
    layer6_outputs(4468) <= not b;
    layer6_outputs(4469) <= b;
    layer6_outputs(4470) <= b and not a;
    layer6_outputs(4471) <= not (a xor b);
    layer6_outputs(4472) <= not (a xor b);
    layer6_outputs(4473) <= a;
    layer6_outputs(4474) <= a;
    layer6_outputs(4475) <= b;
    layer6_outputs(4476) <= not b or a;
    layer6_outputs(4477) <= not b or a;
    layer6_outputs(4478) <= not (a xor b);
    layer6_outputs(4479) <= not b;
    layer6_outputs(4480) <= b;
    layer6_outputs(4481) <= a;
    layer6_outputs(4482) <= not b;
    layer6_outputs(4483) <= not a;
    layer6_outputs(4484) <= '0';
    layer6_outputs(4485) <= a;
    layer6_outputs(4486) <= a;
    layer6_outputs(4487) <= a or b;
    layer6_outputs(4488) <= not a;
    layer6_outputs(4489) <= not (a xor b);
    layer6_outputs(4490) <= b;
    layer6_outputs(4491) <= not a or b;
    layer6_outputs(4492) <= not b;
    layer6_outputs(4493) <= a;
    layer6_outputs(4494) <= not a or b;
    layer6_outputs(4495) <= not b;
    layer6_outputs(4496) <= not (a or b);
    layer6_outputs(4497) <= '0';
    layer6_outputs(4498) <= not b;
    layer6_outputs(4499) <= a;
    layer6_outputs(4500) <= a and not b;
    layer6_outputs(4501) <= b;
    layer6_outputs(4502) <= not b or a;
    layer6_outputs(4503) <= b;
    layer6_outputs(4504) <= b and not a;
    layer6_outputs(4505) <= not b or a;
    layer6_outputs(4506) <= '1';
    layer6_outputs(4507) <= not (a or b);
    layer6_outputs(4508) <= b;
    layer6_outputs(4509) <= not (a and b);
    layer6_outputs(4510) <= b;
    layer6_outputs(4511) <= a;
    layer6_outputs(4512) <= not (a and b);
    layer6_outputs(4513) <= a and b;
    layer6_outputs(4514) <= not b;
    layer6_outputs(4515) <= b;
    layer6_outputs(4516) <= not b;
    layer6_outputs(4517) <= not b;
    layer6_outputs(4518) <= not b;
    layer6_outputs(4519) <= not b;
    layer6_outputs(4520) <= a xor b;
    layer6_outputs(4521) <= not a or b;
    layer6_outputs(4522) <= a;
    layer6_outputs(4523) <= b and not a;
    layer6_outputs(4524) <= not (a or b);
    layer6_outputs(4525) <= not (a xor b);
    layer6_outputs(4526) <= a;
    layer6_outputs(4527) <= not a;
    layer6_outputs(4528) <= a;
    layer6_outputs(4529) <= b;
    layer6_outputs(4530) <= a and not b;
    layer6_outputs(4531) <= not b;
    layer6_outputs(4532) <= not a;
    layer6_outputs(4533) <= a;
    layer6_outputs(4534) <= '1';
    layer6_outputs(4535) <= a;
    layer6_outputs(4536) <= not a or b;
    layer6_outputs(4537) <= a;
    layer6_outputs(4538) <= b and not a;
    layer6_outputs(4539) <= b and not a;
    layer6_outputs(4540) <= not (a xor b);
    layer6_outputs(4541) <= not (a or b);
    layer6_outputs(4542) <= not (a or b);
    layer6_outputs(4543) <= not b or a;
    layer6_outputs(4544) <= a;
    layer6_outputs(4545) <= b;
    layer6_outputs(4546) <= not a or b;
    layer6_outputs(4547) <= a and b;
    layer6_outputs(4548) <= not b or a;
    layer6_outputs(4549) <= not b or a;
    layer6_outputs(4550) <= not a;
    layer6_outputs(4551) <= not b;
    layer6_outputs(4552) <= b;
    layer6_outputs(4553) <= not (a or b);
    layer6_outputs(4554) <= a;
    layer6_outputs(4555) <= a;
    layer6_outputs(4556) <= not (a and b);
    layer6_outputs(4557) <= not b or a;
    layer6_outputs(4558) <= b;
    layer6_outputs(4559) <= b and not a;
    layer6_outputs(4560) <= b;
    layer6_outputs(4561) <= not b;
    layer6_outputs(4562) <= not b;
    layer6_outputs(4563) <= a;
    layer6_outputs(4564) <= a and not b;
    layer6_outputs(4565) <= a xor b;
    layer6_outputs(4566) <= '0';
    layer6_outputs(4567) <= a;
    layer6_outputs(4568) <= not (a or b);
    layer6_outputs(4569) <= not a or b;
    layer6_outputs(4570) <= not (a xor b);
    layer6_outputs(4571) <= not b;
    layer6_outputs(4572) <= b;
    layer6_outputs(4573) <= a;
    layer6_outputs(4574) <= not b;
    layer6_outputs(4575) <= not (a and b);
    layer6_outputs(4576) <= not b or a;
    layer6_outputs(4577) <= a and not b;
    layer6_outputs(4578) <= not a;
    layer6_outputs(4579) <= not (a and b);
    layer6_outputs(4580) <= a and b;
    layer6_outputs(4581) <= not a;
    layer6_outputs(4582) <= a or b;
    layer6_outputs(4583) <= a and b;
    layer6_outputs(4584) <= not b or a;
    layer6_outputs(4585) <= not (a and b);
    layer6_outputs(4586) <= a or b;
    layer6_outputs(4587) <= not (a xor b);
    layer6_outputs(4588) <= not b;
    layer6_outputs(4589) <= not a or b;
    layer6_outputs(4590) <= not b;
    layer6_outputs(4591) <= '0';
    layer6_outputs(4592) <= not b;
    layer6_outputs(4593) <= not b;
    layer6_outputs(4594) <= not (a xor b);
    layer6_outputs(4595) <= not (a and b);
    layer6_outputs(4596) <= '0';
    layer6_outputs(4597) <= not (a and b);
    layer6_outputs(4598) <= '1';
    layer6_outputs(4599) <= b;
    layer6_outputs(4600) <= not b;
    layer6_outputs(4601) <= a and not b;
    layer6_outputs(4602) <= not a or b;
    layer6_outputs(4603) <= not a;
    layer6_outputs(4604) <= b;
    layer6_outputs(4605) <= a;
    layer6_outputs(4606) <= a or b;
    layer6_outputs(4607) <= not (a or b);
    layer6_outputs(4608) <= not a;
    layer6_outputs(4609) <= not b or a;
    layer6_outputs(4610) <= not a;
    layer6_outputs(4611) <= a;
    layer6_outputs(4612) <= not b;
    layer6_outputs(4613) <= a xor b;
    layer6_outputs(4614) <= not a;
    layer6_outputs(4615) <= a;
    layer6_outputs(4616) <= a;
    layer6_outputs(4617) <= b;
    layer6_outputs(4618) <= a and b;
    layer6_outputs(4619) <= not a;
    layer6_outputs(4620) <= not (a xor b);
    layer6_outputs(4621) <= '1';
    layer6_outputs(4622) <= b;
    layer6_outputs(4623) <= '1';
    layer6_outputs(4624) <= a and b;
    layer6_outputs(4625) <= not a;
    layer6_outputs(4626) <= not (a xor b);
    layer6_outputs(4627) <= not (a xor b);
    layer6_outputs(4628) <= not a or b;
    layer6_outputs(4629) <= a;
    layer6_outputs(4630) <= not (a xor b);
    layer6_outputs(4631) <= b and not a;
    layer6_outputs(4632) <= b;
    layer6_outputs(4633) <= not b;
    layer6_outputs(4634) <= a;
    layer6_outputs(4635) <= not a;
    layer6_outputs(4636) <= not a;
    layer6_outputs(4637) <= a and b;
    layer6_outputs(4638) <= a or b;
    layer6_outputs(4639) <= a;
    layer6_outputs(4640) <= not b or a;
    layer6_outputs(4641) <= b and not a;
    layer6_outputs(4642) <= a and not b;
    layer6_outputs(4643) <= a and b;
    layer6_outputs(4644) <= a and not b;
    layer6_outputs(4645) <= a and not b;
    layer6_outputs(4646) <= not b or a;
    layer6_outputs(4647) <= not b or a;
    layer6_outputs(4648) <= a;
    layer6_outputs(4649) <= '0';
    layer6_outputs(4650) <= b;
    layer6_outputs(4651) <= not a;
    layer6_outputs(4652) <= a and not b;
    layer6_outputs(4653) <= not (a or b);
    layer6_outputs(4654) <= not (a or b);
    layer6_outputs(4655) <= a and b;
    layer6_outputs(4656) <= b;
    layer6_outputs(4657) <= not b;
    layer6_outputs(4658) <= a and not b;
    layer6_outputs(4659) <= a or b;
    layer6_outputs(4660) <= not (a xor b);
    layer6_outputs(4661) <= not a or b;
    layer6_outputs(4662) <= not (a or b);
    layer6_outputs(4663) <= not b or a;
    layer6_outputs(4664) <= not b;
    layer6_outputs(4665) <= b and not a;
    layer6_outputs(4666) <= not b;
    layer6_outputs(4667) <= a;
    layer6_outputs(4668) <= not a;
    layer6_outputs(4669) <= a;
    layer6_outputs(4670) <= a and not b;
    layer6_outputs(4671) <= not b or a;
    layer6_outputs(4672) <= b and not a;
    layer6_outputs(4673) <= not a or b;
    layer6_outputs(4674) <= not (a and b);
    layer6_outputs(4675) <= not (a xor b);
    layer6_outputs(4676) <= not b;
    layer6_outputs(4677) <= a and not b;
    layer6_outputs(4678) <= not a;
    layer6_outputs(4679) <= not b;
    layer6_outputs(4680) <= b;
    layer6_outputs(4681) <= a;
    layer6_outputs(4682) <= not b;
    layer6_outputs(4683) <= not a or b;
    layer6_outputs(4684) <= b;
    layer6_outputs(4685) <= a;
    layer6_outputs(4686) <= not a;
    layer6_outputs(4687) <= b and not a;
    layer6_outputs(4688) <= b;
    layer6_outputs(4689) <= '0';
    layer6_outputs(4690) <= not (a or b);
    layer6_outputs(4691) <= not a;
    layer6_outputs(4692) <= not b;
    layer6_outputs(4693) <= not (a xor b);
    layer6_outputs(4694) <= not a or b;
    layer6_outputs(4695) <= a;
    layer6_outputs(4696) <= a;
    layer6_outputs(4697) <= a and b;
    layer6_outputs(4698) <= '0';
    layer6_outputs(4699) <= a;
    layer6_outputs(4700) <= '0';
    layer6_outputs(4701) <= b and not a;
    layer6_outputs(4702) <= a;
    layer6_outputs(4703) <= a and not b;
    layer6_outputs(4704) <= a or b;
    layer6_outputs(4705) <= not b;
    layer6_outputs(4706) <= not a;
    layer6_outputs(4707) <= not a;
    layer6_outputs(4708) <= not a;
    layer6_outputs(4709) <= a;
    layer6_outputs(4710) <= a or b;
    layer6_outputs(4711) <= not a or b;
    layer6_outputs(4712) <= not (a xor b);
    layer6_outputs(4713) <= a or b;
    layer6_outputs(4714) <= a xor b;
    layer6_outputs(4715) <= a and b;
    layer6_outputs(4716) <= b and not a;
    layer6_outputs(4717) <= a and b;
    layer6_outputs(4718) <= a or b;
    layer6_outputs(4719) <= b;
    layer6_outputs(4720) <= not a;
    layer6_outputs(4721) <= not (a xor b);
    layer6_outputs(4722) <= not b;
    layer6_outputs(4723) <= not (a or b);
    layer6_outputs(4724) <= not (a xor b);
    layer6_outputs(4725) <= a;
    layer6_outputs(4726) <= a and not b;
    layer6_outputs(4727) <= not a or b;
    layer6_outputs(4728) <= not a;
    layer6_outputs(4729) <= not b or a;
    layer6_outputs(4730) <= '1';
    layer6_outputs(4731) <= not (a xor b);
    layer6_outputs(4732) <= not (a xor b);
    layer6_outputs(4733) <= not a;
    layer6_outputs(4734) <= not b;
    layer6_outputs(4735) <= not a or b;
    layer6_outputs(4736) <= not (a and b);
    layer6_outputs(4737) <= not (a and b);
    layer6_outputs(4738) <= a;
    layer6_outputs(4739) <= a or b;
    layer6_outputs(4740) <= b and not a;
    layer6_outputs(4741) <= not a or b;
    layer6_outputs(4742) <= a;
    layer6_outputs(4743) <= not a;
    layer6_outputs(4744) <= not (a or b);
    layer6_outputs(4745) <= not b or a;
    layer6_outputs(4746) <= a;
    layer6_outputs(4747) <= a;
    layer6_outputs(4748) <= not a;
    layer6_outputs(4749) <= not (a or b);
    layer6_outputs(4750) <= b;
    layer6_outputs(4751) <= not b;
    layer6_outputs(4752) <= not a;
    layer6_outputs(4753) <= a or b;
    layer6_outputs(4754) <= b and not a;
    layer6_outputs(4755) <= not b;
    layer6_outputs(4756) <= b and not a;
    layer6_outputs(4757) <= not b;
    layer6_outputs(4758) <= a and not b;
    layer6_outputs(4759) <= not a;
    layer6_outputs(4760) <= a and not b;
    layer6_outputs(4761) <= a and not b;
    layer6_outputs(4762) <= a;
    layer6_outputs(4763) <= not (a xor b);
    layer6_outputs(4764) <= a and b;
    layer6_outputs(4765) <= a;
    layer6_outputs(4766) <= b and not a;
    layer6_outputs(4767) <= not a;
    layer6_outputs(4768) <= b and not a;
    layer6_outputs(4769) <= not b;
    layer6_outputs(4770) <= not b or a;
    layer6_outputs(4771) <= a and b;
    layer6_outputs(4772) <= not a or b;
    layer6_outputs(4773) <= a or b;
    layer6_outputs(4774) <= '0';
    layer6_outputs(4775) <= not (a xor b);
    layer6_outputs(4776) <= not a or b;
    layer6_outputs(4777) <= a and not b;
    layer6_outputs(4778) <= not b or a;
    layer6_outputs(4779) <= not a;
    layer6_outputs(4780) <= a xor b;
    layer6_outputs(4781) <= a;
    layer6_outputs(4782) <= not a or b;
    layer6_outputs(4783) <= a xor b;
    layer6_outputs(4784) <= not (a or b);
    layer6_outputs(4785) <= '0';
    layer6_outputs(4786) <= not b or a;
    layer6_outputs(4787) <= b and not a;
    layer6_outputs(4788) <= not a or b;
    layer6_outputs(4789) <= not b;
    layer6_outputs(4790) <= a xor b;
    layer6_outputs(4791) <= not b or a;
    layer6_outputs(4792) <= not (a or b);
    layer6_outputs(4793) <= a xor b;
    layer6_outputs(4794) <= b;
    layer6_outputs(4795) <= not b or a;
    layer6_outputs(4796) <= not a;
    layer6_outputs(4797) <= not a;
    layer6_outputs(4798) <= a xor b;
    layer6_outputs(4799) <= not b or a;
    layer6_outputs(4800) <= not b or a;
    layer6_outputs(4801) <= a;
    layer6_outputs(4802) <= not a;
    layer6_outputs(4803) <= b;
    layer6_outputs(4804) <= a and b;
    layer6_outputs(4805) <= a and not b;
    layer6_outputs(4806) <= not (a xor b);
    layer6_outputs(4807) <= not a;
    layer6_outputs(4808) <= a and not b;
    layer6_outputs(4809) <= '0';
    layer6_outputs(4810) <= not a;
    layer6_outputs(4811) <= not b;
    layer6_outputs(4812) <= b;
    layer6_outputs(4813) <= a or b;
    layer6_outputs(4814) <= b;
    layer6_outputs(4815) <= not a;
    layer6_outputs(4816) <= '1';
    layer6_outputs(4817) <= a and not b;
    layer6_outputs(4818) <= b and not a;
    layer6_outputs(4819) <= a xor b;
    layer6_outputs(4820) <= b;
    layer6_outputs(4821) <= b;
    layer6_outputs(4822) <= not (a xor b);
    layer6_outputs(4823) <= not (a or b);
    layer6_outputs(4824) <= not (a xor b);
    layer6_outputs(4825) <= a and b;
    layer6_outputs(4826) <= a xor b;
    layer6_outputs(4827) <= not (a xor b);
    layer6_outputs(4828) <= not b;
    layer6_outputs(4829) <= a xor b;
    layer6_outputs(4830) <= a and not b;
    layer6_outputs(4831) <= a and b;
    layer6_outputs(4832) <= a xor b;
    layer6_outputs(4833) <= a and not b;
    layer6_outputs(4834) <= not b;
    layer6_outputs(4835) <= b and not a;
    layer6_outputs(4836) <= a and b;
    layer6_outputs(4837) <= '1';
    layer6_outputs(4838) <= not a or b;
    layer6_outputs(4839) <= a or b;
    layer6_outputs(4840) <= not (a and b);
    layer6_outputs(4841) <= b and not a;
    layer6_outputs(4842) <= '0';
    layer6_outputs(4843) <= a;
    layer6_outputs(4844) <= not b;
    layer6_outputs(4845) <= not (a xor b);
    layer6_outputs(4846) <= not b or a;
    layer6_outputs(4847) <= b and not a;
    layer6_outputs(4848) <= b and not a;
    layer6_outputs(4849) <= not b or a;
    layer6_outputs(4850) <= a and b;
    layer6_outputs(4851) <= not a;
    layer6_outputs(4852) <= not a or b;
    layer6_outputs(4853) <= a and not b;
    layer6_outputs(4854) <= not b;
    layer6_outputs(4855) <= not (a and b);
    layer6_outputs(4856) <= not a;
    layer6_outputs(4857) <= '1';
    layer6_outputs(4858) <= a xor b;
    layer6_outputs(4859) <= a and not b;
    layer6_outputs(4860) <= not b;
    layer6_outputs(4861) <= not a;
    layer6_outputs(4862) <= a;
    layer6_outputs(4863) <= b;
    layer6_outputs(4864) <= not (a and b);
    layer6_outputs(4865) <= not a;
    layer6_outputs(4866) <= a and b;
    layer6_outputs(4867) <= '0';
    layer6_outputs(4868) <= not b;
    layer6_outputs(4869) <= not a;
    layer6_outputs(4870) <= b and not a;
    layer6_outputs(4871) <= b;
    layer6_outputs(4872) <= a and not b;
    layer6_outputs(4873) <= a and not b;
    layer6_outputs(4874) <= not a or b;
    layer6_outputs(4875) <= a;
    layer6_outputs(4876) <= a and b;
    layer6_outputs(4877) <= not a;
    layer6_outputs(4878) <= not (a xor b);
    layer6_outputs(4879) <= b and not a;
    layer6_outputs(4880) <= a;
    layer6_outputs(4881) <= not a;
    layer6_outputs(4882) <= not (a and b);
    layer6_outputs(4883) <= a;
    layer6_outputs(4884) <= not b;
    layer6_outputs(4885) <= b and not a;
    layer6_outputs(4886) <= not a;
    layer6_outputs(4887) <= b;
    layer6_outputs(4888) <= not b;
    layer6_outputs(4889) <= b;
    layer6_outputs(4890) <= not (a or b);
    layer6_outputs(4891) <= not a;
    layer6_outputs(4892) <= not b or a;
    layer6_outputs(4893) <= b;
    layer6_outputs(4894) <= b;
    layer6_outputs(4895) <= a and b;
    layer6_outputs(4896) <= a xor b;
    layer6_outputs(4897) <= a;
    layer6_outputs(4898) <= a;
    layer6_outputs(4899) <= not b or a;
    layer6_outputs(4900) <= not (a and b);
    layer6_outputs(4901) <= a and not b;
    layer6_outputs(4902) <= not (a xor b);
    layer6_outputs(4903) <= a and not b;
    layer6_outputs(4904) <= a or b;
    layer6_outputs(4905) <= not a;
    layer6_outputs(4906) <= not a or b;
    layer6_outputs(4907) <= not (a xor b);
    layer6_outputs(4908) <= a;
    layer6_outputs(4909) <= not (a xor b);
    layer6_outputs(4910) <= not (a and b);
    layer6_outputs(4911) <= not a or b;
    layer6_outputs(4912) <= not b or a;
    layer6_outputs(4913) <= not b;
    layer6_outputs(4914) <= not a;
    layer6_outputs(4915) <= '1';
    layer6_outputs(4916) <= b and not a;
    layer6_outputs(4917) <= a and not b;
    layer6_outputs(4918) <= not b;
    layer6_outputs(4919) <= '1';
    layer6_outputs(4920) <= b and not a;
    layer6_outputs(4921) <= not (a xor b);
    layer6_outputs(4922) <= not a;
    layer6_outputs(4923) <= not (a or b);
    layer6_outputs(4924) <= not b or a;
    layer6_outputs(4925) <= not (a xor b);
    layer6_outputs(4926) <= a;
    layer6_outputs(4927) <= not b or a;
    layer6_outputs(4928) <= b and not a;
    layer6_outputs(4929) <= a and not b;
    layer6_outputs(4930) <= not a;
    layer6_outputs(4931) <= a and b;
    layer6_outputs(4932) <= a and b;
    layer6_outputs(4933) <= not (a or b);
    layer6_outputs(4934) <= b;
    layer6_outputs(4935) <= b;
    layer6_outputs(4936) <= b;
    layer6_outputs(4937) <= not b;
    layer6_outputs(4938) <= not (a and b);
    layer6_outputs(4939) <= not (a or b);
    layer6_outputs(4940) <= not b;
    layer6_outputs(4941) <= a and not b;
    layer6_outputs(4942) <= b and not a;
    layer6_outputs(4943) <= not a;
    layer6_outputs(4944) <= not (a and b);
    layer6_outputs(4945) <= not b;
    layer6_outputs(4946) <= not b;
    layer6_outputs(4947) <= not a or b;
    layer6_outputs(4948) <= a and not b;
    layer6_outputs(4949) <= b;
    layer6_outputs(4950) <= not b or a;
    layer6_outputs(4951) <= not b;
    layer6_outputs(4952) <= not b;
    layer6_outputs(4953) <= not a;
    layer6_outputs(4954) <= b and not a;
    layer6_outputs(4955) <= not a or b;
    layer6_outputs(4956) <= a;
    layer6_outputs(4957) <= a xor b;
    layer6_outputs(4958) <= b and not a;
    layer6_outputs(4959) <= not b;
    layer6_outputs(4960) <= not b;
    layer6_outputs(4961) <= a and b;
    layer6_outputs(4962) <= b and not a;
    layer6_outputs(4963) <= a or b;
    layer6_outputs(4964) <= a;
    layer6_outputs(4965) <= a or b;
    layer6_outputs(4966) <= a;
    layer6_outputs(4967) <= not a or b;
    layer6_outputs(4968) <= a and b;
    layer6_outputs(4969) <= '1';
    layer6_outputs(4970) <= a and not b;
    layer6_outputs(4971) <= not a or b;
    layer6_outputs(4972) <= a and b;
    layer6_outputs(4973) <= not a or b;
    layer6_outputs(4974) <= b;
    layer6_outputs(4975) <= not a or b;
    layer6_outputs(4976) <= a and not b;
    layer6_outputs(4977) <= not b or a;
    layer6_outputs(4978) <= not (a or b);
    layer6_outputs(4979) <= not b;
    layer6_outputs(4980) <= not (a and b);
    layer6_outputs(4981) <= not (a xor b);
    layer6_outputs(4982) <= not b;
    layer6_outputs(4983) <= not (a and b);
    layer6_outputs(4984) <= not b;
    layer6_outputs(4985) <= b;
    layer6_outputs(4986) <= not a;
    layer6_outputs(4987) <= not b;
    layer6_outputs(4988) <= not a;
    layer6_outputs(4989) <= a;
    layer6_outputs(4990) <= a xor b;
    layer6_outputs(4991) <= b and not a;
    layer6_outputs(4992) <= b and not a;
    layer6_outputs(4993) <= not a;
    layer6_outputs(4994) <= a and b;
    layer6_outputs(4995) <= a xor b;
    layer6_outputs(4996) <= a and not b;
    layer6_outputs(4997) <= not (a and b);
    layer6_outputs(4998) <= a xor b;
    layer6_outputs(4999) <= a and not b;
    layer6_outputs(5000) <= not (a xor b);
    layer6_outputs(5001) <= b and not a;
    layer6_outputs(5002) <= not (a xor b);
    layer6_outputs(5003) <= b;
    layer6_outputs(5004) <= a and not b;
    layer6_outputs(5005) <= b;
    layer6_outputs(5006) <= not (a and b);
    layer6_outputs(5007) <= b and not a;
    layer6_outputs(5008) <= not (a and b);
    layer6_outputs(5009) <= not a or b;
    layer6_outputs(5010) <= not b;
    layer6_outputs(5011) <= not (a xor b);
    layer6_outputs(5012) <= b;
    layer6_outputs(5013) <= b;
    layer6_outputs(5014) <= not b;
    layer6_outputs(5015) <= a and b;
    layer6_outputs(5016) <= b;
    layer6_outputs(5017) <= not b;
    layer6_outputs(5018) <= not a;
    layer6_outputs(5019) <= not b;
    layer6_outputs(5020) <= not (a xor b);
    layer6_outputs(5021) <= not b or a;
    layer6_outputs(5022) <= not a;
    layer6_outputs(5023) <= a xor b;
    layer6_outputs(5024) <= not b or a;
    layer6_outputs(5025) <= not a;
    layer6_outputs(5026) <= '0';
    layer6_outputs(5027) <= a xor b;
    layer6_outputs(5028) <= not b or a;
    layer6_outputs(5029) <= not (a or b);
    layer6_outputs(5030) <= not a;
    layer6_outputs(5031) <= not a;
    layer6_outputs(5032) <= not a;
    layer6_outputs(5033) <= not (a xor b);
    layer6_outputs(5034) <= a;
    layer6_outputs(5035) <= a and b;
    layer6_outputs(5036) <= not (a or b);
    layer6_outputs(5037) <= not a or b;
    layer6_outputs(5038) <= not b;
    layer6_outputs(5039) <= a or b;
    layer6_outputs(5040) <= not a or b;
    layer6_outputs(5041) <= not a or b;
    layer6_outputs(5042) <= not b or a;
    layer6_outputs(5043) <= not a;
    layer6_outputs(5044) <= not (a xor b);
    layer6_outputs(5045) <= a;
    layer6_outputs(5046) <= a xor b;
    layer6_outputs(5047) <= a;
    layer6_outputs(5048) <= a and b;
    layer6_outputs(5049) <= b and not a;
    layer6_outputs(5050) <= not b or a;
    layer6_outputs(5051) <= not (a and b);
    layer6_outputs(5052) <= a or b;
    layer6_outputs(5053) <= b;
    layer6_outputs(5054) <= not b or a;
    layer6_outputs(5055) <= not (a xor b);
    layer6_outputs(5056) <= not b;
    layer6_outputs(5057) <= not (a or b);
    layer6_outputs(5058) <= a;
    layer6_outputs(5059) <= not (a or b);
    layer6_outputs(5060) <= not (a and b);
    layer6_outputs(5061) <= not a;
    layer6_outputs(5062) <= not (a or b);
    layer6_outputs(5063) <= not b or a;
    layer6_outputs(5064) <= a and not b;
    layer6_outputs(5065) <= not (a or b);
    layer6_outputs(5066) <= not a or b;
    layer6_outputs(5067) <= a and not b;
    layer6_outputs(5068) <= a;
    layer6_outputs(5069) <= a and not b;
    layer6_outputs(5070) <= a and b;
    layer6_outputs(5071) <= not b or a;
    layer6_outputs(5072) <= not b;
    layer6_outputs(5073) <= not (a xor b);
    layer6_outputs(5074) <= b;
    layer6_outputs(5075) <= not (a and b);
    layer6_outputs(5076) <= a;
    layer6_outputs(5077) <= not a or b;
    layer6_outputs(5078) <= not b;
    layer6_outputs(5079) <= a;
    layer6_outputs(5080) <= not (a xor b);
    layer6_outputs(5081) <= b;
    layer6_outputs(5082) <= not b;
    layer6_outputs(5083) <= not (a and b);
    layer6_outputs(5084) <= '1';
    layer6_outputs(5085) <= a or b;
    layer6_outputs(5086) <= a and b;
    layer6_outputs(5087) <= a and b;
    layer6_outputs(5088) <= b;
    layer6_outputs(5089) <= not (a xor b);
    layer6_outputs(5090) <= a;
    layer6_outputs(5091) <= not a or b;
    layer6_outputs(5092) <= a;
    layer6_outputs(5093) <= not a;
    layer6_outputs(5094) <= not a;
    layer6_outputs(5095) <= not b;
    layer6_outputs(5096) <= a or b;
    layer6_outputs(5097) <= not b;
    layer6_outputs(5098) <= not b;
    layer6_outputs(5099) <= not a or b;
    layer6_outputs(5100) <= a xor b;
    layer6_outputs(5101) <= a or b;
    layer6_outputs(5102) <= not (a or b);
    layer6_outputs(5103) <= not a;
    layer6_outputs(5104) <= a xor b;
    layer6_outputs(5105) <= not (a and b);
    layer6_outputs(5106) <= b and not a;
    layer6_outputs(5107) <= not (a xor b);
    layer6_outputs(5108) <= '0';
    layer6_outputs(5109) <= not b or a;
    layer6_outputs(5110) <= b;
    layer6_outputs(5111) <= a or b;
    layer6_outputs(5112) <= '0';
    layer6_outputs(5113) <= a and b;
    layer6_outputs(5114) <= not (a and b);
    layer6_outputs(5115) <= '0';
    layer6_outputs(5116) <= not a;
    layer6_outputs(5117) <= b;
    layer6_outputs(5118) <= b and not a;
    layer6_outputs(5119) <= b and not a;
    layer6_outputs(5120) <= b;
    layer6_outputs(5121) <= a and b;
    layer6_outputs(5122) <= a;
    layer6_outputs(5123) <= not b;
    layer6_outputs(5124) <= a and not b;
    layer6_outputs(5125) <= b and not a;
    layer6_outputs(5126) <= a or b;
    layer6_outputs(5127) <= not a;
    layer6_outputs(5128) <= b;
    layer6_outputs(5129) <= not b;
    layer6_outputs(5130) <= a and b;
    layer6_outputs(5131) <= not a or b;
    layer6_outputs(5132) <= not a or b;
    layer6_outputs(5133) <= not (a or b);
    layer6_outputs(5134) <= not a;
    layer6_outputs(5135) <= a xor b;
    layer6_outputs(5136) <= a;
    layer6_outputs(5137) <= b and not a;
    layer6_outputs(5138) <= a;
    layer6_outputs(5139) <= not (a or b);
    layer6_outputs(5140) <= a xor b;
    layer6_outputs(5141) <= a;
    layer6_outputs(5142) <= b and not a;
    layer6_outputs(5143) <= not (a or b);
    layer6_outputs(5144) <= a and not b;
    layer6_outputs(5145) <= not b or a;
    layer6_outputs(5146) <= not b;
    layer6_outputs(5147) <= a;
    layer6_outputs(5148) <= not (a xor b);
    layer6_outputs(5149) <= a or b;
    layer6_outputs(5150) <= a and b;
    layer6_outputs(5151) <= a or b;
    layer6_outputs(5152) <= not a;
    layer6_outputs(5153) <= a or b;
    layer6_outputs(5154) <= b;
    layer6_outputs(5155) <= not a;
    layer6_outputs(5156) <= a and b;
    layer6_outputs(5157) <= b;
    layer6_outputs(5158) <= not (a or b);
    layer6_outputs(5159) <= not b or a;
    layer6_outputs(5160) <= not a or b;
    layer6_outputs(5161) <= not (a xor b);
    layer6_outputs(5162) <= not (a xor b);
    layer6_outputs(5163) <= a and b;
    layer6_outputs(5164) <= a;
    layer6_outputs(5165) <= a xor b;
    layer6_outputs(5166) <= '1';
    layer6_outputs(5167) <= not b;
    layer6_outputs(5168) <= not b or a;
    layer6_outputs(5169) <= not b or a;
    layer6_outputs(5170) <= a or b;
    layer6_outputs(5171) <= b and not a;
    layer6_outputs(5172) <= a or b;
    layer6_outputs(5173) <= b and not a;
    layer6_outputs(5174) <= b and not a;
    layer6_outputs(5175) <= a and not b;
    layer6_outputs(5176) <= not b;
    layer6_outputs(5177) <= a;
    layer6_outputs(5178) <= b and not a;
    layer6_outputs(5179) <= not (a or b);
    layer6_outputs(5180) <= a;
    layer6_outputs(5181) <= a or b;
    layer6_outputs(5182) <= not b;
    layer6_outputs(5183) <= not b;
    layer6_outputs(5184) <= '1';
    layer6_outputs(5185) <= not (a or b);
    layer6_outputs(5186) <= a and not b;
    layer6_outputs(5187) <= a xor b;
    layer6_outputs(5188) <= not a or b;
    layer6_outputs(5189) <= b;
    layer6_outputs(5190) <= a and b;
    layer6_outputs(5191) <= a;
    layer6_outputs(5192) <= '1';
    layer6_outputs(5193) <= not (a xor b);
    layer6_outputs(5194) <= a or b;
    layer6_outputs(5195) <= not (a or b);
    layer6_outputs(5196) <= a;
    layer6_outputs(5197) <= a or b;
    layer6_outputs(5198) <= not a or b;
    layer6_outputs(5199) <= not a or b;
    layer6_outputs(5200) <= b;
    layer6_outputs(5201) <= not (a and b);
    layer6_outputs(5202) <= b;
    layer6_outputs(5203) <= a and b;
    layer6_outputs(5204) <= b;
    layer6_outputs(5205) <= not a or b;
    layer6_outputs(5206) <= not b or a;
    layer6_outputs(5207) <= not a;
    layer6_outputs(5208) <= not a;
    layer6_outputs(5209) <= a;
    layer6_outputs(5210) <= not (a and b);
    layer6_outputs(5211) <= not (a and b);
    layer6_outputs(5212) <= not a;
    layer6_outputs(5213) <= not a;
    layer6_outputs(5214) <= a or b;
    layer6_outputs(5215) <= not a or b;
    layer6_outputs(5216) <= not (a and b);
    layer6_outputs(5217) <= not b;
    layer6_outputs(5218) <= a;
    layer6_outputs(5219) <= a and b;
    layer6_outputs(5220) <= b;
    layer6_outputs(5221) <= a or b;
    layer6_outputs(5222) <= b;
    layer6_outputs(5223) <= not (a and b);
    layer6_outputs(5224) <= a;
    layer6_outputs(5225) <= not a or b;
    layer6_outputs(5226) <= not b;
    layer6_outputs(5227) <= not a or b;
    layer6_outputs(5228) <= '0';
    layer6_outputs(5229) <= not a;
    layer6_outputs(5230) <= a or b;
    layer6_outputs(5231) <= b;
    layer6_outputs(5232) <= not a or b;
    layer6_outputs(5233) <= a;
    layer6_outputs(5234) <= not b;
    layer6_outputs(5235) <= '0';
    layer6_outputs(5236) <= not (a or b);
    layer6_outputs(5237) <= not (a or b);
    layer6_outputs(5238) <= '1';
    layer6_outputs(5239) <= not a;
    layer6_outputs(5240) <= a and b;
    layer6_outputs(5241) <= a;
    layer6_outputs(5242) <= a and not b;
    layer6_outputs(5243) <= a xor b;
    layer6_outputs(5244) <= b;
    layer6_outputs(5245) <= not (a or b);
    layer6_outputs(5246) <= '1';
    layer6_outputs(5247) <= not a;
    layer6_outputs(5248) <= not a;
    layer6_outputs(5249) <= a;
    layer6_outputs(5250) <= a;
    layer6_outputs(5251) <= not b or a;
    layer6_outputs(5252) <= a;
    layer6_outputs(5253) <= not (a and b);
    layer6_outputs(5254) <= not a or b;
    layer6_outputs(5255) <= not (a and b);
    layer6_outputs(5256) <= a;
    layer6_outputs(5257) <= not a;
    layer6_outputs(5258) <= not a or b;
    layer6_outputs(5259) <= not a or b;
    layer6_outputs(5260) <= '1';
    layer6_outputs(5261) <= a;
    layer6_outputs(5262) <= b;
    layer6_outputs(5263) <= not b;
    layer6_outputs(5264) <= not a;
    layer6_outputs(5265) <= '0';
    layer6_outputs(5266) <= a and not b;
    layer6_outputs(5267) <= not a or b;
    layer6_outputs(5268) <= not b;
    layer6_outputs(5269) <= not (a xor b);
    layer6_outputs(5270) <= a and not b;
    layer6_outputs(5271) <= not b or a;
    layer6_outputs(5272) <= not a;
    layer6_outputs(5273) <= a;
    layer6_outputs(5274) <= not (a or b);
    layer6_outputs(5275) <= not a or b;
    layer6_outputs(5276) <= not (a and b);
    layer6_outputs(5277) <= a or b;
    layer6_outputs(5278) <= not (a xor b);
    layer6_outputs(5279) <= not b or a;
    layer6_outputs(5280) <= '0';
    layer6_outputs(5281) <= a xor b;
    layer6_outputs(5282) <= not b or a;
    layer6_outputs(5283) <= not b or a;
    layer6_outputs(5284) <= not a or b;
    layer6_outputs(5285) <= not b;
    layer6_outputs(5286) <= not b or a;
    layer6_outputs(5287) <= b;
    layer6_outputs(5288) <= not b or a;
    layer6_outputs(5289) <= '0';
    layer6_outputs(5290) <= a or b;
    layer6_outputs(5291) <= not b;
    layer6_outputs(5292) <= a;
    layer6_outputs(5293) <= not a or b;
    layer6_outputs(5294) <= a xor b;
    layer6_outputs(5295) <= a or b;
    layer6_outputs(5296) <= not a;
    layer6_outputs(5297) <= not a or b;
    layer6_outputs(5298) <= not (a or b);
    layer6_outputs(5299) <= not a;
    layer6_outputs(5300) <= a and b;
    layer6_outputs(5301) <= a;
    layer6_outputs(5302) <= not a or b;
    layer6_outputs(5303) <= not (a xor b);
    layer6_outputs(5304) <= b;
    layer6_outputs(5305) <= not (a or b);
    layer6_outputs(5306) <= not (a or b);
    layer6_outputs(5307) <= a;
    layer6_outputs(5308) <= not a;
    layer6_outputs(5309) <= not a;
    layer6_outputs(5310) <= not (a and b);
    layer6_outputs(5311) <= a;
    layer6_outputs(5312) <= a and b;
    layer6_outputs(5313) <= not b;
    layer6_outputs(5314) <= not b or a;
    layer6_outputs(5315) <= '0';
    layer6_outputs(5316) <= b and not a;
    layer6_outputs(5317) <= not b or a;
    layer6_outputs(5318) <= b and not a;
    layer6_outputs(5319) <= a xor b;
    layer6_outputs(5320) <= '0';
    layer6_outputs(5321) <= b;
    layer6_outputs(5322) <= b;
    layer6_outputs(5323) <= not b;
    layer6_outputs(5324) <= not (a and b);
    layer6_outputs(5325) <= '0';
    layer6_outputs(5326) <= a;
    layer6_outputs(5327) <= not a;
    layer6_outputs(5328) <= not b or a;
    layer6_outputs(5329) <= b;
    layer6_outputs(5330) <= a or b;
    layer6_outputs(5331) <= not a;
    layer6_outputs(5332) <= not (a or b);
    layer6_outputs(5333) <= a xor b;
    layer6_outputs(5334) <= a;
    layer6_outputs(5335) <= not a;
    layer6_outputs(5336) <= not (a or b);
    layer6_outputs(5337) <= not (a xor b);
    layer6_outputs(5338) <= b and not a;
    layer6_outputs(5339) <= b;
    layer6_outputs(5340) <= a xor b;
    layer6_outputs(5341) <= a;
    layer6_outputs(5342) <= a or b;
    layer6_outputs(5343) <= not a;
    layer6_outputs(5344) <= b and not a;
    layer6_outputs(5345) <= a and not b;
    layer6_outputs(5346) <= not b;
    layer6_outputs(5347) <= a or b;
    layer6_outputs(5348) <= a or b;
    layer6_outputs(5349) <= not (a and b);
    layer6_outputs(5350) <= not (a and b);
    layer6_outputs(5351) <= not (a and b);
    layer6_outputs(5352) <= not (a and b);
    layer6_outputs(5353) <= a;
    layer6_outputs(5354) <= not b or a;
    layer6_outputs(5355) <= '1';
    layer6_outputs(5356) <= a xor b;
    layer6_outputs(5357) <= not b or a;
    layer6_outputs(5358) <= a or b;
    layer6_outputs(5359) <= a or b;
    layer6_outputs(5360) <= not (a xor b);
    layer6_outputs(5361) <= not b;
    layer6_outputs(5362) <= a and not b;
    layer6_outputs(5363) <= not b or a;
    layer6_outputs(5364) <= not b;
    layer6_outputs(5365) <= not (a and b);
    layer6_outputs(5366) <= a;
    layer6_outputs(5367) <= not a or b;
    layer6_outputs(5368) <= not b or a;
    layer6_outputs(5369) <= not (a or b);
    layer6_outputs(5370) <= a xor b;
    layer6_outputs(5371) <= b and not a;
    layer6_outputs(5372) <= b and not a;
    layer6_outputs(5373) <= not b;
    layer6_outputs(5374) <= not (a or b);
    layer6_outputs(5375) <= a or b;
    layer6_outputs(5376) <= not a or b;
    layer6_outputs(5377) <= a or b;
    layer6_outputs(5378) <= not a;
    layer6_outputs(5379) <= a and not b;
    layer6_outputs(5380) <= a or b;
    layer6_outputs(5381) <= a xor b;
    layer6_outputs(5382) <= a;
    layer6_outputs(5383) <= b;
    layer6_outputs(5384) <= b;
    layer6_outputs(5385) <= b;
    layer6_outputs(5386) <= a;
    layer6_outputs(5387) <= a xor b;
    layer6_outputs(5388) <= not a;
    layer6_outputs(5389) <= '1';
    layer6_outputs(5390) <= not (a xor b);
    layer6_outputs(5391) <= b and not a;
    layer6_outputs(5392) <= not b or a;
    layer6_outputs(5393) <= b and not a;
    layer6_outputs(5394) <= not a;
    layer6_outputs(5395) <= a and not b;
    layer6_outputs(5396) <= not b or a;
    layer6_outputs(5397) <= a and not b;
    layer6_outputs(5398) <= '1';
    layer6_outputs(5399) <= not a or b;
    layer6_outputs(5400) <= a;
    layer6_outputs(5401) <= a and not b;
    layer6_outputs(5402) <= not a;
    layer6_outputs(5403) <= not (a and b);
    layer6_outputs(5404) <= not b;
    layer6_outputs(5405) <= not b;
    layer6_outputs(5406) <= b;
    layer6_outputs(5407) <= not a or b;
    layer6_outputs(5408) <= b;
    layer6_outputs(5409) <= not a;
    layer6_outputs(5410) <= not b;
    layer6_outputs(5411) <= not (a or b);
    layer6_outputs(5412) <= a and not b;
    layer6_outputs(5413) <= a and not b;
    layer6_outputs(5414) <= a xor b;
    layer6_outputs(5415) <= not a;
    layer6_outputs(5416) <= not (a xor b);
    layer6_outputs(5417) <= not a or b;
    layer6_outputs(5418) <= a and not b;
    layer6_outputs(5419) <= a xor b;
    layer6_outputs(5420) <= a or b;
    layer6_outputs(5421) <= b;
    layer6_outputs(5422) <= a or b;
    layer6_outputs(5423) <= b;
    layer6_outputs(5424) <= not b or a;
    layer6_outputs(5425) <= a;
    layer6_outputs(5426) <= a or b;
    layer6_outputs(5427) <= a xor b;
    layer6_outputs(5428) <= not b;
    layer6_outputs(5429) <= not (a or b);
    layer6_outputs(5430) <= a and not b;
    layer6_outputs(5431) <= b and not a;
    layer6_outputs(5432) <= a;
    layer6_outputs(5433) <= a xor b;
    layer6_outputs(5434) <= not a;
    layer6_outputs(5435) <= not (a and b);
    layer6_outputs(5436) <= not (a xor b);
    layer6_outputs(5437) <= a xor b;
    layer6_outputs(5438) <= a;
    layer6_outputs(5439) <= a;
    layer6_outputs(5440) <= b and not a;
    layer6_outputs(5441) <= not a or b;
    layer6_outputs(5442) <= not a;
    layer6_outputs(5443) <= not a or b;
    layer6_outputs(5444) <= b and not a;
    layer6_outputs(5445) <= not a or b;
    layer6_outputs(5446) <= a;
    layer6_outputs(5447) <= b;
    layer6_outputs(5448) <= not b;
    layer6_outputs(5449) <= b;
    layer6_outputs(5450) <= b;
    layer6_outputs(5451) <= not a or b;
    layer6_outputs(5452) <= not a or b;
    layer6_outputs(5453) <= a;
    layer6_outputs(5454) <= not b;
    layer6_outputs(5455) <= not (a and b);
    layer6_outputs(5456) <= not a;
    layer6_outputs(5457) <= a;
    layer6_outputs(5458) <= a and b;
    layer6_outputs(5459) <= not a;
    layer6_outputs(5460) <= not a or b;
    layer6_outputs(5461) <= b;
    layer6_outputs(5462) <= not a or b;
    layer6_outputs(5463) <= a and b;
    layer6_outputs(5464) <= a or b;
    layer6_outputs(5465) <= not a;
    layer6_outputs(5466) <= a;
    layer6_outputs(5467) <= a;
    layer6_outputs(5468) <= a or b;
    layer6_outputs(5469) <= b;
    layer6_outputs(5470) <= not a or b;
    layer6_outputs(5471) <= not b;
    layer6_outputs(5472) <= not b or a;
    layer6_outputs(5473) <= not (a xor b);
    layer6_outputs(5474) <= '1';
    layer6_outputs(5475) <= a;
    layer6_outputs(5476) <= a or b;
    layer6_outputs(5477) <= not a or b;
    layer6_outputs(5478) <= a or b;
    layer6_outputs(5479) <= a and b;
    layer6_outputs(5480) <= a xor b;
    layer6_outputs(5481) <= b and not a;
    layer6_outputs(5482) <= not a;
    layer6_outputs(5483) <= a;
    layer6_outputs(5484) <= b;
    layer6_outputs(5485) <= a;
    layer6_outputs(5486) <= a or b;
    layer6_outputs(5487) <= not a;
    layer6_outputs(5488) <= a and not b;
    layer6_outputs(5489) <= not b;
    layer6_outputs(5490) <= a;
    layer6_outputs(5491) <= not a;
    layer6_outputs(5492) <= not a or b;
    layer6_outputs(5493) <= not (a or b);
    layer6_outputs(5494) <= not (a xor b);
    layer6_outputs(5495) <= not b or a;
    layer6_outputs(5496) <= not (a and b);
    layer6_outputs(5497) <= not a;
    layer6_outputs(5498) <= not a;
    layer6_outputs(5499) <= b and not a;
    layer6_outputs(5500) <= b;
    layer6_outputs(5501) <= not b or a;
    layer6_outputs(5502) <= '0';
    layer6_outputs(5503) <= not b;
    layer6_outputs(5504) <= b and not a;
    layer6_outputs(5505) <= not a;
    layer6_outputs(5506) <= b and not a;
    layer6_outputs(5507) <= not b;
    layer6_outputs(5508) <= a and b;
    layer6_outputs(5509) <= a or b;
    layer6_outputs(5510) <= a xor b;
    layer6_outputs(5511) <= a;
    layer6_outputs(5512) <= '0';
    layer6_outputs(5513) <= b and not a;
    layer6_outputs(5514) <= not a;
    layer6_outputs(5515) <= not a or b;
    layer6_outputs(5516) <= a and not b;
    layer6_outputs(5517) <= not b;
    layer6_outputs(5518) <= a and not b;
    layer6_outputs(5519) <= a;
    layer6_outputs(5520) <= not b;
    layer6_outputs(5521) <= a;
    layer6_outputs(5522) <= a;
    layer6_outputs(5523) <= b;
    layer6_outputs(5524) <= not a or b;
    layer6_outputs(5525) <= b and not a;
    layer6_outputs(5526) <= a or b;
    layer6_outputs(5527) <= not b;
    layer6_outputs(5528) <= not b or a;
    layer6_outputs(5529) <= a;
    layer6_outputs(5530) <= '1';
    layer6_outputs(5531) <= not b or a;
    layer6_outputs(5532) <= not a or b;
    layer6_outputs(5533) <= a and not b;
    layer6_outputs(5534) <= not (a or b);
    layer6_outputs(5535) <= not b;
    layer6_outputs(5536) <= a;
    layer6_outputs(5537) <= a and not b;
    layer6_outputs(5538) <= not a;
    layer6_outputs(5539) <= not b or a;
    layer6_outputs(5540) <= a;
    layer6_outputs(5541) <= b and not a;
    layer6_outputs(5542) <= a xor b;
    layer6_outputs(5543) <= a and b;
    layer6_outputs(5544) <= not b;
    layer6_outputs(5545) <= a or b;
    layer6_outputs(5546) <= b and not a;
    layer6_outputs(5547) <= not a;
    layer6_outputs(5548) <= b;
    layer6_outputs(5549) <= not b;
    layer6_outputs(5550) <= not b;
    layer6_outputs(5551) <= not b;
    layer6_outputs(5552) <= not (a and b);
    layer6_outputs(5553) <= a xor b;
    layer6_outputs(5554) <= not a or b;
    layer6_outputs(5555) <= a;
    layer6_outputs(5556) <= not (a or b);
    layer6_outputs(5557) <= a or b;
    layer6_outputs(5558) <= b;
    layer6_outputs(5559) <= not b or a;
    layer6_outputs(5560) <= a;
    layer6_outputs(5561) <= b;
    layer6_outputs(5562) <= a;
    layer6_outputs(5563) <= a and not b;
    layer6_outputs(5564) <= a xor b;
    layer6_outputs(5565) <= not (a xor b);
    layer6_outputs(5566) <= a;
    layer6_outputs(5567) <= b;
    layer6_outputs(5568) <= '0';
    layer6_outputs(5569) <= not (a and b);
    layer6_outputs(5570) <= not b;
    layer6_outputs(5571) <= not b;
    layer6_outputs(5572) <= not (a or b);
    layer6_outputs(5573) <= not a or b;
    layer6_outputs(5574) <= not b;
    layer6_outputs(5575) <= b;
    layer6_outputs(5576) <= not (a or b);
    layer6_outputs(5577) <= not (a or b);
    layer6_outputs(5578) <= not a or b;
    layer6_outputs(5579) <= not (a or b);
    layer6_outputs(5580) <= not (a xor b);
    layer6_outputs(5581) <= not (a or b);
    layer6_outputs(5582) <= b;
    layer6_outputs(5583) <= not b;
    layer6_outputs(5584) <= not b;
    layer6_outputs(5585) <= not a;
    layer6_outputs(5586) <= a and not b;
    layer6_outputs(5587) <= not (a or b);
    layer6_outputs(5588) <= a and not b;
    layer6_outputs(5589) <= a and not b;
    layer6_outputs(5590) <= not (a xor b);
    layer6_outputs(5591) <= a and b;
    layer6_outputs(5592) <= not (a or b);
    layer6_outputs(5593) <= a;
    layer6_outputs(5594) <= '0';
    layer6_outputs(5595) <= not b;
    layer6_outputs(5596) <= not (a or b);
    layer6_outputs(5597) <= a and not b;
    layer6_outputs(5598) <= not (a or b);
    layer6_outputs(5599) <= not (a xor b);
    layer6_outputs(5600) <= a;
    layer6_outputs(5601) <= not b or a;
    layer6_outputs(5602) <= '0';
    layer6_outputs(5603) <= b;
    layer6_outputs(5604) <= not b;
    layer6_outputs(5605) <= a;
    layer6_outputs(5606) <= not (a or b);
    layer6_outputs(5607) <= a xor b;
    layer6_outputs(5608) <= not a;
    layer6_outputs(5609) <= not (a or b);
    layer6_outputs(5610) <= '1';
    layer6_outputs(5611) <= b;
    layer6_outputs(5612) <= not b or a;
    layer6_outputs(5613) <= b;
    layer6_outputs(5614) <= not (a or b);
    layer6_outputs(5615) <= not b or a;
    layer6_outputs(5616) <= a or b;
    layer6_outputs(5617) <= b;
    layer6_outputs(5618) <= b;
    layer6_outputs(5619) <= not (a or b);
    layer6_outputs(5620) <= '1';
    layer6_outputs(5621) <= not a or b;
    layer6_outputs(5622) <= '1';
    layer6_outputs(5623) <= not b;
    layer6_outputs(5624) <= not b;
    layer6_outputs(5625) <= a xor b;
    layer6_outputs(5626) <= not a;
    layer6_outputs(5627) <= '0';
    layer6_outputs(5628) <= not a or b;
    layer6_outputs(5629) <= not (a and b);
    layer6_outputs(5630) <= not b or a;
    layer6_outputs(5631) <= not a;
    layer6_outputs(5632) <= not a or b;
    layer6_outputs(5633) <= a;
    layer6_outputs(5634) <= b;
    layer6_outputs(5635) <= a or b;
    layer6_outputs(5636) <= '0';
    layer6_outputs(5637) <= not a;
    layer6_outputs(5638) <= b;
    layer6_outputs(5639) <= not a or b;
    layer6_outputs(5640) <= a xor b;
    layer6_outputs(5641) <= not (a and b);
    layer6_outputs(5642) <= not (a xor b);
    layer6_outputs(5643) <= a or b;
    layer6_outputs(5644) <= a and b;
    layer6_outputs(5645) <= not a;
    layer6_outputs(5646) <= a and not b;
    layer6_outputs(5647) <= a;
    layer6_outputs(5648) <= b;
    layer6_outputs(5649) <= not (a and b);
    layer6_outputs(5650) <= b;
    layer6_outputs(5651) <= b and not a;
    layer6_outputs(5652) <= not (a xor b);
    layer6_outputs(5653) <= '0';
    layer6_outputs(5654) <= not (a and b);
    layer6_outputs(5655) <= a and b;
    layer6_outputs(5656) <= a xor b;
    layer6_outputs(5657) <= a;
    layer6_outputs(5658) <= not (a xor b);
    layer6_outputs(5659) <= not b;
    layer6_outputs(5660) <= b;
    layer6_outputs(5661) <= not (a xor b);
    layer6_outputs(5662) <= not a;
    layer6_outputs(5663) <= not (a and b);
    layer6_outputs(5664) <= not a;
    layer6_outputs(5665) <= a;
    layer6_outputs(5666) <= not b;
    layer6_outputs(5667) <= not b or a;
    layer6_outputs(5668) <= not (a or b);
    layer6_outputs(5669) <= a and not b;
    layer6_outputs(5670) <= b;
    layer6_outputs(5671) <= b and not a;
    layer6_outputs(5672) <= not a;
    layer6_outputs(5673) <= a and b;
    layer6_outputs(5674) <= not b;
    layer6_outputs(5675) <= a and b;
    layer6_outputs(5676) <= not (a and b);
    layer6_outputs(5677) <= not a or b;
    layer6_outputs(5678) <= a or b;
    layer6_outputs(5679) <= not b;
    layer6_outputs(5680) <= a and not b;
    layer6_outputs(5681) <= not b;
    layer6_outputs(5682) <= a and not b;
    layer6_outputs(5683) <= not a or b;
    layer6_outputs(5684) <= '1';
    layer6_outputs(5685) <= a or b;
    layer6_outputs(5686) <= not (a or b);
    layer6_outputs(5687) <= a or b;
    layer6_outputs(5688) <= not (a or b);
    layer6_outputs(5689) <= a;
    layer6_outputs(5690) <= a and not b;
    layer6_outputs(5691) <= a;
    layer6_outputs(5692) <= a xor b;
    layer6_outputs(5693) <= a and b;
    layer6_outputs(5694) <= a or b;
    layer6_outputs(5695) <= not a;
    layer6_outputs(5696) <= a and b;
    layer6_outputs(5697) <= a and b;
    layer6_outputs(5698) <= a;
    layer6_outputs(5699) <= not a or b;
    layer6_outputs(5700) <= not b or a;
    layer6_outputs(5701) <= a;
    layer6_outputs(5702) <= a or b;
    layer6_outputs(5703) <= a and not b;
    layer6_outputs(5704) <= not (a xor b);
    layer6_outputs(5705) <= not (a and b);
    layer6_outputs(5706) <= b and not a;
    layer6_outputs(5707) <= not a;
    layer6_outputs(5708) <= not b;
    layer6_outputs(5709) <= a or b;
    layer6_outputs(5710) <= b;
    layer6_outputs(5711) <= a;
    layer6_outputs(5712) <= not (a xor b);
    layer6_outputs(5713) <= b and not a;
    layer6_outputs(5714) <= a or b;
    layer6_outputs(5715) <= a;
    layer6_outputs(5716) <= a;
    layer6_outputs(5717) <= a and not b;
    layer6_outputs(5718) <= not a;
    layer6_outputs(5719) <= a;
    layer6_outputs(5720) <= a and not b;
    layer6_outputs(5721) <= not a or b;
    layer6_outputs(5722) <= a and not b;
    layer6_outputs(5723) <= not b;
    layer6_outputs(5724) <= not (a or b);
    layer6_outputs(5725) <= a and not b;
    layer6_outputs(5726) <= not b or a;
    layer6_outputs(5727) <= not b;
    layer6_outputs(5728) <= not b or a;
    layer6_outputs(5729) <= b and not a;
    layer6_outputs(5730) <= not b;
    layer6_outputs(5731) <= b;
    layer6_outputs(5732) <= not (a and b);
    layer6_outputs(5733) <= not (a or b);
    layer6_outputs(5734) <= b;
    layer6_outputs(5735) <= '1';
    layer6_outputs(5736) <= b;
    layer6_outputs(5737) <= not a;
    layer6_outputs(5738) <= a or b;
    layer6_outputs(5739) <= a and not b;
    layer6_outputs(5740) <= a;
    layer6_outputs(5741) <= not (a or b);
    layer6_outputs(5742) <= a and b;
    layer6_outputs(5743) <= a or b;
    layer6_outputs(5744) <= a and not b;
    layer6_outputs(5745) <= not b;
    layer6_outputs(5746) <= not (a and b);
    layer6_outputs(5747) <= a or b;
    layer6_outputs(5748) <= '0';
    layer6_outputs(5749) <= not (a xor b);
    layer6_outputs(5750) <= not a;
    layer6_outputs(5751) <= not a or b;
    layer6_outputs(5752) <= not a;
    layer6_outputs(5753) <= not a or b;
    layer6_outputs(5754) <= b and not a;
    layer6_outputs(5755) <= not a or b;
    layer6_outputs(5756) <= b and not a;
    layer6_outputs(5757) <= '1';
    layer6_outputs(5758) <= '0';
    layer6_outputs(5759) <= a xor b;
    layer6_outputs(5760) <= not a;
    layer6_outputs(5761) <= a;
    layer6_outputs(5762) <= not b;
    layer6_outputs(5763) <= not a;
    layer6_outputs(5764) <= b;
    layer6_outputs(5765) <= '0';
    layer6_outputs(5766) <= not b;
    layer6_outputs(5767) <= a or b;
    layer6_outputs(5768) <= not b or a;
    layer6_outputs(5769) <= b;
    layer6_outputs(5770) <= not (a and b);
    layer6_outputs(5771) <= a and b;
    layer6_outputs(5772) <= b;
    layer6_outputs(5773) <= a or b;
    layer6_outputs(5774) <= not (a xor b);
    layer6_outputs(5775) <= not (a and b);
    layer6_outputs(5776) <= b and not a;
    layer6_outputs(5777) <= not (a or b);
    layer6_outputs(5778) <= not b or a;
    layer6_outputs(5779) <= not a;
    layer6_outputs(5780) <= a;
    layer6_outputs(5781) <= '1';
    layer6_outputs(5782) <= b;
    layer6_outputs(5783) <= not b or a;
    layer6_outputs(5784) <= a or b;
    layer6_outputs(5785) <= not a;
    layer6_outputs(5786) <= a and b;
    layer6_outputs(5787) <= b and not a;
    layer6_outputs(5788) <= not a;
    layer6_outputs(5789) <= not a;
    layer6_outputs(5790) <= b;
    layer6_outputs(5791) <= not (a or b);
    layer6_outputs(5792) <= not b or a;
    layer6_outputs(5793) <= a or b;
    layer6_outputs(5794) <= b;
    layer6_outputs(5795) <= not (a xor b);
    layer6_outputs(5796) <= not a;
    layer6_outputs(5797) <= not b;
    layer6_outputs(5798) <= not b or a;
    layer6_outputs(5799) <= a and not b;
    layer6_outputs(5800) <= not (a and b);
    layer6_outputs(5801) <= a and not b;
    layer6_outputs(5802) <= not a;
    layer6_outputs(5803) <= not (a or b);
    layer6_outputs(5804) <= not (a xor b);
    layer6_outputs(5805) <= not (a xor b);
    layer6_outputs(5806) <= b and not a;
    layer6_outputs(5807) <= not b;
    layer6_outputs(5808) <= not a or b;
    layer6_outputs(5809) <= not b;
    layer6_outputs(5810) <= not a or b;
    layer6_outputs(5811) <= not b;
    layer6_outputs(5812) <= a and b;
    layer6_outputs(5813) <= not b or a;
    layer6_outputs(5814) <= '1';
    layer6_outputs(5815) <= a;
    layer6_outputs(5816) <= b and not a;
    layer6_outputs(5817) <= a xor b;
    layer6_outputs(5818) <= b;
    layer6_outputs(5819) <= not (a xor b);
    layer6_outputs(5820) <= not b;
    layer6_outputs(5821) <= not (a or b);
    layer6_outputs(5822) <= not (a and b);
    layer6_outputs(5823) <= not b;
    layer6_outputs(5824) <= a and not b;
    layer6_outputs(5825) <= b;
    layer6_outputs(5826) <= a xor b;
    layer6_outputs(5827) <= not (a or b);
    layer6_outputs(5828) <= b and not a;
    layer6_outputs(5829) <= a;
    layer6_outputs(5830) <= a and not b;
    layer6_outputs(5831) <= not (a and b);
    layer6_outputs(5832) <= a;
    layer6_outputs(5833) <= a or b;
    layer6_outputs(5834) <= a and b;
    layer6_outputs(5835) <= b and not a;
    layer6_outputs(5836) <= not (a or b);
    layer6_outputs(5837) <= a;
    layer6_outputs(5838) <= not b or a;
    layer6_outputs(5839) <= a or b;
    layer6_outputs(5840) <= not b;
    layer6_outputs(5841) <= not (a xor b);
    layer6_outputs(5842) <= not a;
    layer6_outputs(5843) <= not a;
    layer6_outputs(5844) <= not b;
    layer6_outputs(5845) <= not (a and b);
    layer6_outputs(5846) <= a and not b;
    layer6_outputs(5847) <= a;
    layer6_outputs(5848) <= '1';
    layer6_outputs(5849) <= a or b;
    layer6_outputs(5850) <= not b or a;
    layer6_outputs(5851) <= not a;
    layer6_outputs(5852) <= not b;
    layer6_outputs(5853) <= a and not b;
    layer6_outputs(5854) <= not a;
    layer6_outputs(5855) <= not (a and b);
    layer6_outputs(5856) <= not b;
    layer6_outputs(5857) <= b;
    layer6_outputs(5858) <= a;
    layer6_outputs(5859) <= b;
    layer6_outputs(5860) <= not (a and b);
    layer6_outputs(5861) <= not a or b;
    layer6_outputs(5862) <= a;
    layer6_outputs(5863) <= not (a and b);
    layer6_outputs(5864) <= not b;
    layer6_outputs(5865) <= '0';
    layer6_outputs(5866) <= not (a and b);
    layer6_outputs(5867) <= not b;
    layer6_outputs(5868) <= b;
    layer6_outputs(5869) <= not a or b;
    layer6_outputs(5870) <= b;
    layer6_outputs(5871) <= a and b;
    layer6_outputs(5872) <= a;
    layer6_outputs(5873) <= b;
    layer6_outputs(5874) <= b and not a;
    layer6_outputs(5875) <= not a;
    layer6_outputs(5876) <= a;
    layer6_outputs(5877) <= not b;
    layer6_outputs(5878) <= not (a xor b);
    layer6_outputs(5879) <= a and not b;
    layer6_outputs(5880) <= b and not a;
    layer6_outputs(5881) <= not (a or b);
    layer6_outputs(5882) <= not b or a;
    layer6_outputs(5883) <= b;
    layer6_outputs(5884) <= not a;
    layer6_outputs(5885) <= a and not b;
    layer6_outputs(5886) <= not (a and b);
    layer6_outputs(5887) <= a xor b;
    layer6_outputs(5888) <= b;
    layer6_outputs(5889) <= b and not a;
    layer6_outputs(5890) <= not (a xor b);
    layer6_outputs(5891) <= a and b;
    layer6_outputs(5892) <= a;
    layer6_outputs(5893) <= not b;
    layer6_outputs(5894) <= a or b;
    layer6_outputs(5895) <= '1';
    layer6_outputs(5896) <= not (a xor b);
    layer6_outputs(5897) <= a xor b;
    layer6_outputs(5898) <= a;
    layer6_outputs(5899) <= not b or a;
    layer6_outputs(5900) <= not b;
    layer6_outputs(5901) <= a and not b;
    layer6_outputs(5902) <= a and not b;
    layer6_outputs(5903) <= b;
    layer6_outputs(5904) <= a and b;
    layer6_outputs(5905) <= not (a xor b);
    layer6_outputs(5906) <= not (a and b);
    layer6_outputs(5907) <= b and not a;
    layer6_outputs(5908) <= a;
    layer6_outputs(5909) <= not a;
    layer6_outputs(5910) <= not (a xor b);
    layer6_outputs(5911) <= not b;
    layer6_outputs(5912) <= not (a or b);
    layer6_outputs(5913) <= not b or a;
    layer6_outputs(5914) <= not b or a;
    layer6_outputs(5915) <= a;
    layer6_outputs(5916) <= a and not b;
    layer6_outputs(5917) <= a;
    layer6_outputs(5918) <= a and not b;
    layer6_outputs(5919) <= b and not a;
    layer6_outputs(5920) <= not a or b;
    layer6_outputs(5921) <= '0';
    layer6_outputs(5922) <= not (a and b);
    layer6_outputs(5923) <= not b;
    layer6_outputs(5924) <= not a or b;
    layer6_outputs(5925) <= not (a and b);
    layer6_outputs(5926) <= b and not a;
    layer6_outputs(5927) <= b;
    layer6_outputs(5928) <= not a;
    layer6_outputs(5929) <= not (a and b);
    layer6_outputs(5930) <= b;
    layer6_outputs(5931) <= a xor b;
    layer6_outputs(5932) <= not b;
    layer6_outputs(5933) <= a or b;
    layer6_outputs(5934) <= not a;
    layer6_outputs(5935) <= a;
    layer6_outputs(5936) <= not (a and b);
    layer6_outputs(5937) <= a;
    layer6_outputs(5938) <= b;
    layer6_outputs(5939) <= not (a xor b);
    layer6_outputs(5940) <= not b or a;
    layer6_outputs(5941) <= not b;
    layer6_outputs(5942) <= not (a or b);
    layer6_outputs(5943) <= not a or b;
    layer6_outputs(5944) <= not a;
    layer6_outputs(5945) <= '1';
    layer6_outputs(5946) <= '0';
    layer6_outputs(5947) <= not (a and b);
    layer6_outputs(5948) <= a;
    layer6_outputs(5949) <= not b;
    layer6_outputs(5950) <= not a or b;
    layer6_outputs(5951) <= b and not a;
    layer6_outputs(5952) <= not b;
    layer6_outputs(5953) <= a or b;
    layer6_outputs(5954) <= a or b;
    layer6_outputs(5955) <= b;
    layer6_outputs(5956) <= a and not b;
    layer6_outputs(5957) <= b;
    layer6_outputs(5958) <= not b or a;
    layer6_outputs(5959) <= b;
    layer6_outputs(5960) <= a or b;
    layer6_outputs(5961) <= not a or b;
    layer6_outputs(5962) <= a;
    layer6_outputs(5963) <= a and b;
    layer6_outputs(5964) <= not (a xor b);
    layer6_outputs(5965) <= a or b;
    layer6_outputs(5966) <= not a or b;
    layer6_outputs(5967) <= a;
    layer6_outputs(5968) <= a;
    layer6_outputs(5969) <= a or b;
    layer6_outputs(5970) <= b;
    layer6_outputs(5971) <= not a or b;
    layer6_outputs(5972) <= b;
    layer6_outputs(5973) <= b;
    layer6_outputs(5974) <= a and b;
    layer6_outputs(5975) <= not (a or b);
    layer6_outputs(5976) <= a and not b;
    layer6_outputs(5977) <= b;
    layer6_outputs(5978) <= a or b;
    layer6_outputs(5979) <= a or b;
    layer6_outputs(5980) <= a or b;
    layer6_outputs(5981) <= not (a or b);
    layer6_outputs(5982) <= not (a or b);
    layer6_outputs(5983) <= not (a and b);
    layer6_outputs(5984) <= b and not a;
    layer6_outputs(5985) <= not (a xor b);
    layer6_outputs(5986) <= not (a or b);
    layer6_outputs(5987) <= not (a or b);
    layer6_outputs(5988) <= b;
    layer6_outputs(5989) <= not (a and b);
    layer6_outputs(5990) <= not b or a;
    layer6_outputs(5991) <= not (a and b);
    layer6_outputs(5992) <= not (a xor b);
    layer6_outputs(5993) <= b;
    layer6_outputs(5994) <= a or b;
    layer6_outputs(5995) <= not a;
    layer6_outputs(5996) <= not a or b;
    layer6_outputs(5997) <= not a;
    layer6_outputs(5998) <= a and b;
    layer6_outputs(5999) <= not b or a;
    layer6_outputs(6000) <= b and not a;
    layer6_outputs(6001) <= not (a or b);
    layer6_outputs(6002) <= a xor b;
    layer6_outputs(6003) <= a and not b;
    layer6_outputs(6004) <= not (a or b);
    layer6_outputs(6005) <= not b;
    layer6_outputs(6006) <= not b or a;
    layer6_outputs(6007) <= not (a xor b);
    layer6_outputs(6008) <= not (a and b);
    layer6_outputs(6009) <= not a or b;
    layer6_outputs(6010) <= '1';
    layer6_outputs(6011) <= b and not a;
    layer6_outputs(6012) <= not a;
    layer6_outputs(6013) <= not a;
    layer6_outputs(6014) <= a xor b;
    layer6_outputs(6015) <= a xor b;
    layer6_outputs(6016) <= not a;
    layer6_outputs(6017) <= not a;
    layer6_outputs(6018) <= not b;
    layer6_outputs(6019) <= a;
    layer6_outputs(6020) <= a and not b;
    layer6_outputs(6021) <= a and b;
    layer6_outputs(6022) <= not (a and b);
    layer6_outputs(6023) <= not b;
    layer6_outputs(6024) <= a xor b;
    layer6_outputs(6025) <= not b;
    layer6_outputs(6026) <= a and b;
    layer6_outputs(6027) <= b;
    layer6_outputs(6028) <= not b;
    layer6_outputs(6029) <= '1';
    layer6_outputs(6030) <= not (a xor b);
    layer6_outputs(6031) <= not b;
    layer6_outputs(6032) <= not a;
    layer6_outputs(6033) <= '1';
    layer6_outputs(6034) <= not b;
    layer6_outputs(6035) <= not (a and b);
    layer6_outputs(6036) <= not b or a;
    layer6_outputs(6037) <= a;
    layer6_outputs(6038) <= a and not b;
    layer6_outputs(6039) <= b;
    layer6_outputs(6040) <= '1';
    layer6_outputs(6041) <= not b or a;
    layer6_outputs(6042) <= not b or a;
    layer6_outputs(6043) <= a xor b;
    layer6_outputs(6044) <= not (a and b);
    layer6_outputs(6045) <= a xor b;
    layer6_outputs(6046) <= not (a or b);
    layer6_outputs(6047) <= not (a and b);
    layer6_outputs(6048) <= not (a and b);
    layer6_outputs(6049) <= a and b;
    layer6_outputs(6050) <= not (a xor b);
    layer6_outputs(6051) <= a xor b;
    layer6_outputs(6052) <= not b or a;
    layer6_outputs(6053) <= not a or b;
    layer6_outputs(6054) <= a or b;
    layer6_outputs(6055) <= b;
    layer6_outputs(6056) <= b;
    layer6_outputs(6057) <= not a or b;
    layer6_outputs(6058) <= '1';
    layer6_outputs(6059) <= '0';
    layer6_outputs(6060) <= a;
    layer6_outputs(6061) <= b;
    layer6_outputs(6062) <= a;
    layer6_outputs(6063) <= not b or a;
    layer6_outputs(6064) <= a and not b;
    layer6_outputs(6065) <= not a or b;
    layer6_outputs(6066) <= not b;
    layer6_outputs(6067) <= a;
    layer6_outputs(6068) <= b;
    layer6_outputs(6069) <= b;
    layer6_outputs(6070) <= a or b;
    layer6_outputs(6071) <= a xor b;
    layer6_outputs(6072) <= not (a or b);
    layer6_outputs(6073) <= b;
    layer6_outputs(6074) <= a;
    layer6_outputs(6075) <= not (a or b);
    layer6_outputs(6076) <= a or b;
    layer6_outputs(6077) <= b;
    layer6_outputs(6078) <= a and not b;
    layer6_outputs(6079) <= a or b;
    layer6_outputs(6080) <= not a or b;
    layer6_outputs(6081) <= a;
    layer6_outputs(6082) <= not a;
    layer6_outputs(6083) <= a and b;
    layer6_outputs(6084) <= not a;
    layer6_outputs(6085) <= a or b;
    layer6_outputs(6086) <= not a or b;
    layer6_outputs(6087) <= not a or b;
    layer6_outputs(6088) <= not a;
    layer6_outputs(6089) <= a or b;
    layer6_outputs(6090) <= not a;
    layer6_outputs(6091) <= a;
    layer6_outputs(6092) <= not (a xor b);
    layer6_outputs(6093) <= not b;
    layer6_outputs(6094) <= not b or a;
    layer6_outputs(6095) <= b;
    layer6_outputs(6096) <= not b;
    layer6_outputs(6097) <= b and not a;
    layer6_outputs(6098) <= b and not a;
    layer6_outputs(6099) <= a or b;
    layer6_outputs(6100) <= not a or b;
    layer6_outputs(6101) <= not a;
    layer6_outputs(6102) <= not (a or b);
    layer6_outputs(6103) <= not (a and b);
    layer6_outputs(6104) <= a and b;
    layer6_outputs(6105) <= '0';
    layer6_outputs(6106) <= a xor b;
    layer6_outputs(6107) <= a or b;
    layer6_outputs(6108) <= not a;
    layer6_outputs(6109) <= a;
    layer6_outputs(6110) <= not b or a;
    layer6_outputs(6111) <= b and not a;
    layer6_outputs(6112) <= not (a xor b);
    layer6_outputs(6113) <= '1';
    layer6_outputs(6114) <= b and not a;
    layer6_outputs(6115) <= b;
    layer6_outputs(6116) <= b and not a;
    layer6_outputs(6117) <= not a;
    layer6_outputs(6118) <= b;
    layer6_outputs(6119) <= not b or a;
    layer6_outputs(6120) <= not b;
    layer6_outputs(6121) <= a and b;
    layer6_outputs(6122) <= a and not b;
    layer6_outputs(6123) <= not a or b;
    layer6_outputs(6124) <= a or b;
    layer6_outputs(6125) <= not b;
    layer6_outputs(6126) <= not (a and b);
    layer6_outputs(6127) <= not b;
    layer6_outputs(6128) <= not a;
    layer6_outputs(6129) <= a;
    layer6_outputs(6130) <= not a or b;
    layer6_outputs(6131) <= not a;
    layer6_outputs(6132) <= a;
    layer6_outputs(6133) <= a or b;
    layer6_outputs(6134) <= not a or b;
    layer6_outputs(6135) <= b;
    layer6_outputs(6136) <= not (a xor b);
    layer6_outputs(6137) <= not b;
    layer6_outputs(6138) <= a;
    layer6_outputs(6139) <= a xor b;
    layer6_outputs(6140) <= '0';
    layer6_outputs(6141) <= not a or b;
    layer6_outputs(6142) <= not (a and b);
    layer6_outputs(6143) <= '1';
    layer6_outputs(6144) <= not (a or b);
    layer6_outputs(6145) <= a and not b;
    layer6_outputs(6146) <= b and not a;
    layer6_outputs(6147) <= a and not b;
    layer6_outputs(6148) <= not b;
    layer6_outputs(6149) <= a or b;
    layer6_outputs(6150) <= not a;
    layer6_outputs(6151) <= not a or b;
    layer6_outputs(6152) <= not b or a;
    layer6_outputs(6153) <= not (a or b);
    layer6_outputs(6154) <= a and not b;
    layer6_outputs(6155) <= a;
    layer6_outputs(6156) <= not b;
    layer6_outputs(6157) <= a and not b;
    layer6_outputs(6158) <= not b or a;
    layer6_outputs(6159) <= not (a and b);
    layer6_outputs(6160) <= not (a or b);
    layer6_outputs(6161) <= b and not a;
    layer6_outputs(6162) <= not a or b;
    layer6_outputs(6163) <= a or b;
    layer6_outputs(6164) <= '1';
    layer6_outputs(6165) <= '0';
    layer6_outputs(6166) <= not b;
    layer6_outputs(6167) <= not (a and b);
    layer6_outputs(6168) <= a;
    layer6_outputs(6169) <= a and b;
    layer6_outputs(6170) <= b;
    layer6_outputs(6171) <= not b;
    layer6_outputs(6172) <= b and not a;
    layer6_outputs(6173) <= not (a xor b);
    layer6_outputs(6174) <= b;
    layer6_outputs(6175) <= not a or b;
    layer6_outputs(6176) <= not (a xor b);
    layer6_outputs(6177) <= a and not b;
    layer6_outputs(6178) <= a and b;
    layer6_outputs(6179) <= not (a or b);
    layer6_outputs(6180) <= not b or a;
    layer6_outputs(6181) <= not a;
    layer6_outputs(6182) <= b and not a;
    layer6_outputs(6183) <= a and b;
    layer6_outputs(6184) <= not (a and b);
    layer6_outputs(6185) <= a;
    layer6_outputs(6186) <= a or b;
    layer6_outputs(6187) <= a and b;
    layer6_outputs(6188) <= not a;
    layer6_outputs(6189) <= not b or a;
    layer6_outputs(6190) <= a and not b;
    layer6_outputs(6191) <= not (a or b);
    layer6_outputs(6192) <= a or b;
    layer6_outputs(6193) <= a or b;
    layer6_outputs(6194) <= '1';
    layer6_outputs(6195) <= not (a or b);
    layer6_outputs(6196) <= '0';
    layer6_outputs(6197) <= a;
    layer6_outputs(6198) <= not b;
    layer6_outputs(6199) <= a or b;
    layer6_outputs(6200) <= b and not a;
    layer6_outputs(6201) <= a;
    layer6_outputs(6202) <= a;
    layer6_outputs(6203) <= b and not a;
    layer6_outputs(6204) <= a and b;
    layer6_outputs(6205) <= a and b;
    layer6_outputs(6206) <= not (a and b);
    layer6_outputs(6207) <= a and not b;
    layer6_outputs(6208) <= not a or b;
    layer6_outputs(6209) <= not a or b;
    layer6_outputs(6210) <= a;
    layer6_outputs(6211) <= a and not b;
    layer6_outputs(6212) <= not (a or b);
    layer6_outputs(6213) <= not a;
    layer6_outputs(6214) <= a or b;
    layer6_outputs(6215) <= b and not a;
    layer6_outputs(6216) <= not (a or b);
    layer6_outputs(6217) <= b;
    layer6_outputs(6218) <= not (a or b);
    layer6_outputs(6219) <= not b or a;
    layer6_outputs(6220) <= not a or b;
    layer6_outputs(6221) <= not (a or b);
    layer6_outputs(6222) <= not a;
    layer6_outputs(6223) <= not (a and b);
    layer6_outputs(6224) <= a and b;
    layer6_outputs(6225) <= a and not b;
    layer6_outputs(6226) <= not b;
    layer6_outputs(6227) <= not b;
    layer6_outputs(6228) <= not a;
    layer6_outputs(6229) <= not b or a;
    layer6_outputs(6230) <= not (a or b);
    layer6_outputs(6231) <= not b or a;
    layer6_outputs(6232) <= a;
    layer6_outputs(6233) <= not (a or b);
    layer6_outputs(6234) <= a or b;
    layer6_outputs(6235) <= not b;
    layer6_outputs(6236) <= not b;
    layer6_outputs(6237) <= not b;
    layer6_outputs(6238) <= not (a or b);
    layer6_outputs(6239) <= b;
    layer6_outputs(6240) <= '1';
    layer6_outputs(6241) <= a;
    layer6_outputs(6242) <= not a;
    layer6_outputs(6243) <= b;
    layer6_outputs(6244) <= a and b;
    layer6_outputs(6245) <= not a;
    layer6_outputs(6246) <= a;
    layer6_outputs(6247) <= not a;
    layer6_outputs(6248) <= b;
    layer6_outputs(6249) <= a and not b;
    layer6_outputs(6250) <= not b;
    layer6_outputs(6251) <= a or b;
    layer6_outputs(6252) <= a or b;
    layer6_outputs(6253) <= b and not a;
    layer6_outputs(6254) <= b;
    layer6_outputs(6255) <= a;
    layer6_outputs(6256) <= not a;
    layer6_outputs(6257) <= not a or b;
    layer6_outputs(6258) <= a or b;
    layer6_outputs(6259) <= b and not a;
    layer6_outputs(6260) <= not b or a;
    layer6_outputs(6261) <= b and not a;
    layer6_outputs(6262) <= not (a xor b);
    layer6_outputs(6263) <= not b;
    layer6_outputs(6264) <= a or b;
    layer6_outputs(6265) <= a and not b;
    layer6_outputs(6266) <= b;
    layer6_outputs(6267) <= b;
    layer6_outputs(6268) <= not (a xor b);
    layer6_outputs(6269) <= b;
    layer6_outputs(6270) <= not a;
    layer6_outputs(6271) <= b;
    layer6_outputs(6272) <= not b or a;
    layer6_outputs(6273) <= not (a or b);
    layer6_outputs(6274) <= b and not a;
    layer6_outputs(6275) <= not a;
    layer6_outputs(6276) <= not a;
    layer6_outputs(6277) <= a and b;
    layer6_outputs(6278) <= a and b;
    layer6_outputs(6279) <= a;
    layer6_outputs(6280) <= b and not a;
    layer6_outputs(6281) <= a and not b;
    layer6_outputs(6282) <= b;
    layer6_outputs(6283) <= b;
    layer6_outputs(6284) <= a and not b;
    layer6_outputs(6285) <= a and b;
    layer6_outputs(6286) <= a and not b;
    layer6_outputs(6287) <= a and b;
    layer6_outputs(6288) <= '1';
    layer6_outputs(6289) <= not a;
    layer6_outputs(6290) <= not b;
    layer6_outputs(6291) <= b and not a;
    layer6_outputs(6292) <= b and not a;
    layer6_outputs(6293) <= b;
    layer6_outputs(6294) <= not (a and b);
    layer6_outputs(6295) <= not b;
    layer6_outputs(6296) <= a or b;
    layer6_outputs(6297) <= not (a or b);
    layer6_outputs(6298) <= a xor b;
    layer6_outputs(6299) <= b and not a;
    layer6_outputs(6300) <= not b or a;
    layer6_outputs(6301) <= not a;
    layer6_outputs(6302) <= b;
    layer6_outputs(6303) <= a;
    layer6_outputs(6304) <= a and not b;
    layer6_outputs(6305) <= not a;
    layer6_outputs(6306) <= a or b;
    layer6_outputs(6307) <= a and not b;
    layer6_outputs(6308) <= not b;
    layer6_outputs(6309) <= not b;
    layer6_outputs(6310) <= not b or a;
    layer6_outputs(6311) <= a and b;
    layer6_outputs(6312) <= a;
    layer6_outputs(6313) <= a;
    layer6_outputs(6314) <= not b;
    layer6_outputs(6315) <= not b;
    layer6_outputs(6316) <= not a or b;
    layer6_outputs(6317) <= a;
    layer6_outputs(6318) <= not (a or b);
    layer6_outputs(6319) <= not (a and b);
    layer6_outputs(6320) <= not a;
    layer6_outputs(6321) <= b;
    layer6_outputs(6322) <= a or b;
    layer6_outputs(6323) <= a and not b;
    layer6_outputs(6324) <= not a;
    layer6_outputs(6325) <= a;
    layer6_outputs(6326) <= a and not b;
    layer6_outputs(6327) <= not a or b;
    layer6_outputs(6328) <= not a;
    layer6_outputs(6329) <= a;
    layer6_outputs(6330) <= b;
    layer6_outputs(6331) <= not b;
    layer6_outputs(6332) <= a;
    layer6_outputs(6333) <= a and b;
    layer6_outputs(6334) <= not a;
    layer6_outputs(6335) <= a or b;
    layer6_outputs(6336) <= not a;
    layer6_outputs(6337) <= not (a or b);
    layer6_outputs(6338) <= a and not b;
    layer6_outputs(6339) <= a and not b;
    layer6_outputs(6340) <= not a or b;
    layer6_outputs(6341) <= not a or b;
    layer6_outputs(6342) <= not (a or b);
    layer6_outputs(6343) <= not (a or b);
    layer6_outputs(6344) <= not b;
    layer6_outputs(6345) <= not b or a;
    layer6_outputs(6346) <= not a;
    layer6_outputs(6347) <= not (a xor b);
    layer6_outputs(6348) <= not a or b;
    layer6_outputs(6349) <= a;
    layer6_outputs(6350) <= not a;
    layer6_outputs(6351) <= b;
    layer6_outputs(6352) <= not (a or b);
    layer6_outputs(6353) <= '0';
    layer6_outputs(6354) <= a xor b;
    layer6_outputs(6355) <= not (a xor b);
    layer6_outputs(6356) <= not b;
    layer6_outputs(6357) <= a and b;
    layer6_outputs(6358) <= not b or a;
    layer6_outputs(6359) <= not b;
    layer6_outputs(6360) <= not (a xor b);
    layer6_outputs(6361) <= a or b;
    layer6_outputs(6362) <= not a or b;
    layer6_outputs(6363) <= not a or b;
    layer6_outputs(6364) <= b;
    layer6_outputs(6365) <= a;
    layer6_outputs(6366) <= not a;
    layer6_outputs(6367) <= a or b;
    layer6_outputs(6368) <= not b;
    layer6_outputs(6369) <= not a or b;
    layer6_outputs(6370) <= b;
    layer6_outputs(6371) <= not (a xor b);
    layer6_outputs(6372) <= b;
    layer6_outputs(6373) <= a and not b;
    layer6_outputs(6374) <= not a;
    layer6_outputs(6375) <= not (a and b);
    layer6_outputs(6376) <= a or b;
    layer6_outputs(6377) <= b and not a;
    layer6_outputs(6378) <= b and not a;
    layer6_outputs(6379) <= not b;
    layer6_outputs(6380) <= not a;
    layer6_outputs(6381) <= not (a or b);
    layer6_outputs(6382) <= a;
    layer6_outputs(6383) <= not (a or b);
    layer6_outputs(6384) <= not b or a;
    layer6_outputs(6385) <= a and b;
    layer6_outputs(6386) <= not (a or b);
    layer6_outputs(6387) <= not (a and b);
    layer6_outputs(6388) <= not a;
    layer6_outputs(6389) <= b and not a;
    layer6_outputs(6390) <= not b;
    layer6_outputs(6391) <= a and not b;
    layer6_outputs(6392) <= b and not a;
    layer6_outputs(6393) <= not (a or b);
    layer6_outputs(6394) <= not (a or b);
    layer6_outputs(6395) <= a and b;
    layer6_outputs(6396) <= '1';
    layer6_outputs(6397) <= not a or b;
    layer6_outputs(6398) <= not b or a;
    layer6_outputs(6399) <= a xor b;
    layer6_outputs(6400) <= b and not a;
    layer6_outputs(6401) <= not (a xor b);
    layer6_outputs(6402) <= a;
    layer6_outputs(6403) <= not (a and b);
    layer6_outputs(6404) <= not a;
    layer6_outputs(6405) <= not (a and b);
    layer6_outputs(6406) <= b and not a;
    layer6_outputs(6407) <= not (a xor b);
    layer6_outputs(6408) <= not a or b;
    layer6_outputs(6409) <= not a;
    layer6_outputs(6410) <= not a or b;
    layer6_outputs(6411) <= a;
    layer6_outputs(6412) <= b;
    layer6_outputs(6413) <= not (a or b);
    layer6_outputs(6414) <= not a;
    layer6_outputs(6415) <= b;
    layer6_outputs(6416) <= not b;
    layer6_outputs(6417) <= b;
    layer6_outputs(6418) <= not (a xor b);
    layer6_outputs(6419) <= not (a or b);
    layer6_outputs(6420) <= not (a and b);
    layer6_outputs(6421) <= not (a or b);
    layer6_outputs(6422) <= not b;
    layer6_outputs(6423) <= a;
    layer6_outputs(6424) <= not b;
    layer6_outputs(6425) <= b;
    layer6_outputs(6426) <= '1';
    layer6_outputs(6427) <= a;
    layer6_outputs(6428) <= a xor b;
    layer6_outputs(6429) <= not b;
    layer6_outputs(6430) <= not (a xor b);
    layer6_outputs(6431) <= not b;
    layer6_outputs(6432) <= not b or a;
    layer6_outputs(6433) <= a and b;
    layer6_outputs(6434) <= not a;
    layer6_outputs(6435) <= a and b;
    layer6_outputs(6436) <= not a or b;
    layer6_outputs(6437) <= not a or b;
    layer6_outputs(6438) <= not (a and b);
    layer6_outputs(6439) <= not a or b;
    layer6_outputs(6440) <= a and b;
    layer6_outputs(6441) <= a;
    layer6_outputs(6442) <= a;
    layer6_outputs(6443) <= a and not b;
    layer6_outputs(6444) <= not (a and b);
    layer6_outputs(6445) <= not (a xor b);
    layer6_outputs(6446) <= a;
    layer6_outputs(6447) <= a;
    layer6_outputs(6448) <= a and b;
    layer6_outputs(6449) <= not b or a;
    layer6_outputs(6450) <= not b;
    layer6_outputs(6451) <= a and not b;
    layer6_outputs(6452) <= not a or b;
    layer6_outputs(6453) <= not b;
    layer6_outputs(6454) <= a and b;
    layer6_outputs(6455) <= a and not b;
    layer6_outputs(6456) <= '0';
    layer6_outputs(6457) <= not b;
    layer6_outputs(6458) <= b;
    layer6_outputs(6459) <= b;
    layer6_outputs(6460) <= b and not a;
    layer6_outputs(6461) <= a;
    layer6_outputs(6462) <= b and not a;
    layer6_outputs(6463) <= a and b;
    layer6_outputs(6464) <= a or b;
    layer6_outputs(6465) <= a;
    layer6_outputs(6466) <= b and not a;
    layer6_outputs(6467) <= a;
    layer6_outputs(6468) <= a and b;
    layer6_outputs(6469) <= not (a and b);
    layer6_outputs(6470) <= not b;
    layer6_outputs(6471) <= not b or a;
    layer6_outputs(6472) <= a or b;
    layer6_outputs(6473) <= b;
    layer6_outputs(6474) <= not a;
    layer6_outputs(6475) <= not a;
    layer6_outputs(6476) <= a and not b;
    layer6_outputs(6477) <= not b;
    layer6_outputs(6478) <= a and not b;
    layer6_outputs(6479) <= not a;
    layer6_outputs(6480) <= b and not a;
    layer6_outputs(6481) <= a or b;
    layer6_outputs(6482) <= a or b;
    layer6_outputs(6483) <= '0';
    layer6_outputs(6484) <= a;
    layer6_outputs(6485) <= not b;
    layer6_outputs(6486) <= '0';
    layer6_outputs(6487) <= not a;
    layer6_outputs(6488) <= a xor b;
    layer6_outputs(6489) <= a;
    layer6_outputs(6490) <= b;
    layer6_outputs(6491) <= a xor b;
    layer6_outputs(6492) <= not (a and b);
    layer6_outputs(6493) <= not (a or b);
    layer6_outputs(6494) <= '0';
    layer6_outputs(6495) <= a and not b;
    layer6_outputs(6496) <= not (a and b);
    layer6_outputs(6497) <= b;
    layer6_outputs(6498) <= a;
    layer6_outputs(6499) <= b and not a;
    layer6_outputs(6500) <= not (a or b);
    layer6_outputs(6501) <= a and b;
    layer6_outputs(6502) <= not (a and b);
    layer6_outputs(6503) <= not b or a;
    layer6_outputs(6504) <= b and not a;
    layer6_outputs(6505) <= a and b;
    layer6_outputs(6506) <= not b;
    layer6_outputs(6507) <= '1';
    layer6_outputs(6508) <= not b;
    layer6_outputs(6509) <= not b;
    layer6_outputs(6510) <= not (a or b);
    layer6_outputs(6511) <= not a;
    layer6_outputs(6512) <= not (a and b);
    layer6_outputs(6513) <= not (a and b);
    layer6_outputs(6514) <= a and not b;
    layer6_outputs(6515) <= b and not a;
    layer6_outputs(6516) <= a and b;
    layer6_outputs(6517) <= not b;
    layer6_outputs(6518) <= a and not b;
    layer6_outputs(6519) <= not (a and b);
    layer6_outputs(6520) <= a xor b;
    layer6_outputs(6521) <= not (a and b);
    layer6_outputs(6522) <= b;
    layer6_outputs(6523) <= '1';
    layer6_outputs(6524) <= b;
    layer6_outputs(6525) <= not (a xor b);
    layer6_outputs(6526) <= not (a or b);
    layer6_outputs(6527) <= b and not a;
    layer6_outputs(6528) <= a or b;
    layer6_outputs(6529) <= b;
    layer6_outputs(6530) <= a and not b;
    layer6_outputs(6531) <= not (a and b);
    layer6_outputs(6532) <= not a;
    layer6_outputs(6533) <= a;
    layer6_outputs(6534) <= not (a or b);
    layer6_outputs(6535) <= a and b;
    layer6_outputs(6536) <= not a;
    layer6_outputs(6537) <= not (a and b);
    layer6_outputs(6538) <= b;
    layer6_outputs(6539) <= b and not a;
    layer6_outputs(6540) <= not a;
    layer6_outputs(6541) <= a and b;
    layer6_outputs(6542) <= not a;
    layer6_outputs(6543) <= a or b;
    layer6_outputs(6544) <= not a or b;
    layer6_outputs(6545) <= a and not b;
    layer6_outputs(6546) <= a;
    layer6_outputs(6547) <= a and not b;
    layer6_outputs(6548) <= a;
    layer6_outputs(6549) <= a and b;
    layer6_outputs(6550) <= not b;
    layer6_outputs(6551) <= not b or a;
    layer6_outputs(6552) <= not b or a;
    layer6_outputs(6553) <= not a;
    layer6_outputs(6554) <= b;
    layer6_outputs(6555) <= b and not a;
    layer6_outputs(6556) <= a;
    layer6_outputs(6557) <= not b;
    layer6_outputs(6558) <= a;
    layer6_outputs(6559) <= not a or b;
    layer6_outputs(6560) <= not b;
    layer6_outputs(6561) <= a;
    layer6_outputs(6562) <= a and b;
    layer6_outputs(6563) <= a and not b;
    layer6_outputs(6564) <= not a;
    layer6_outputs(6565) <= not (a and b);
    layer6_outputs(6566) <= a or b;
    layer6_outputs(6567) <= b;
    layer6_outputs(6568) <= a xor b;
    layer6_outputs(6569) <= b and not a;
    layer6_outputs(6570) <= '0';
    layer6_outputs(6571) <= not a or b;
    layer6_outputs(6572) <= a and b;
    layer6_outputs(6573) <= not b;
    layer6_outputs(6574) <= not b;
    layer6_outputs(6575) <= not b;
    layer6_outputs(6576) <= not (a xor b);
    layer6_outputs(6577) <= a;
    layer6_outputs(6578) <= a;
    layer6_outputs(6579) <= b;
    layer6_outputs(6580) <= not (a and b);
    layer6_outputs(6581) <= a xor b;
    layer6_outputs(6582) <= a xor b;
    layer6_outputs(6583) <= b;
    layer6_outputs(6584) <= a;
    layer6_outputs(6585) <= b;
    layer6_outputs(6586) <= not (a and b);
    layer6_outputs(6587) <= not (a or b);
    layer6_outputs(6588) <= '0';
    layer6_outputs(6589) <= not (a or b);
    layer6_outputs(6590) <= b;
    layer6_outputs(6591) <= a xor b;
    layer6_outputs(6592) <= b and not a;
    layer6_outputs(6593) <= b;
    layer6_outputs(6594) <= not (a and b);
    layer6_outputs(6595) <= not b;
    layer6_outputs(6596) <= not a;
    layer6_outputs(6597) <= not (a or b);
    layer6_outputs(6598) <= not (a xor b);
    layer6_outputs(6599) <= a or b;
    layer6_outputs(6600) <= '0';
    layer6_outputs(6601) <= '0';
    layer6_outputs(6602) <= '1';
    layer6_outputs(6603) <= not a or b;
    layer6_outputs(6604) <= b;
    layer6_outputs(6605) <= a and b;
    layer6_outputs(6606) <= not a or b;
    layer6_outputs(6607) <= not b or a;
    layer6_outputs(6608) <= b;
    layer6_outputs(6609) <= not (a or b);
    layer6_outputs(6610) <= a and not b;
    layer6_outputs(6611) <= not a;
    layer6_outputs(6612) <= not a;
    layer6_outputs(6613) <= a and not b;
    layer6_outputs(6614) <= not (a or b);
    layer6_outputs(6615) <= not b or a;
    layer6_outputs(6616) <= a and not b;
    layer6_outputs(6617) <= '1';
    layer6_outputs(6618) <= not a or b;
    layer6_outputs(6619) <= b;
    layer6_outputs(6620) <= not a;
    layer6_outputs(6621) <= a and not b;
    layer6_outputs(6622) <= not b or a;
    layer6_outputs(6623) <= not a or b;
    layer6_outputs(6624) <= not a;
    layer6_outputs(6625) <= b;
    layer6_outputs(6626) <= b;
    layer6_outputs(6627) <= not b;
    layer6_outputs(6628) <= not a;
    layer6_outputs(6629) <= a or b;
    layer6_outputs(6630) <= a;
    layer6_outputs(6631) <= not b or a;
    layer6_outputs(6632) <= a or b;
    layer6_outputs(6633) <= not a or b;
    layer6_outputs(6634) <= '1';
    layer6_outputs(6635) <= a or b;
    layer6_outputs(6636) <= not a;
    layer6_outputs(6637) <= a;
    layer6_outputs(6638) <= a or b;
    layer6_outputs(6639) <= a xor b;
    layer6_outputs(6640) <= a;
    layer6_outputs(6641) <= a;
    layer6_outputs(6642) <= a or b;
    layer6_outputs(6643) <= a;
    layer6_outputs(6644) <= b and not a;
    layer6_outputs(6645) <= a and b;
    layer6_outputs(6646) <= b and not a;
    layer6_outputs(6647) <= b and not a;
    layer6_outputs(6648) <= not (a xor b);
    layer6_outputs(6649) <= not (a xor b);
    layer6_outputs(6650) <= not b or a;
    layer6_outputs(6651) <= a;
    layer6_outputs(6652) <= not (a xor b);
    layer6_outputs(6653) <= not (a and b);
    layer6_outputs(6654) <= not (a xor b);
    layer6_outputs(6655) <= b and not a;
    layer6_outputs(6656) <= not b;
    layer6_outputs(6657) <= b and not a;
    layer6_outputs(6658) <= not a or b;
    layer6_outputs(6659) <= not a or b;
    layer6_outputs(6660) <= not a;
    layer6_outputs(6661) <= not b or a;
    layer6_outputs(6662) <= not b;
    layer6_outputs(6663) <= not b;
    layer6_outputs(6664) <= b;
    layer6_outputs(6665) <= not a;
    layer6_outputs(6666) <= not b or a;
    layer6_outputs(6667) <= b;
    layer6_outputs(6668) <= not (a and b);
    layer6_outputs(6669) <= '1';
    layer6_outputs(6670) <= not (a and b);
    layer6_outputs(6671) <= not (a xor b);
    layer6_outputs(6672) <= a and b;
    layer6_outputs(6673) <= a;
    layer6_outputs(6674) <= a and not b;
    layer6_outputs(6675) <= b and not a;
    layer6_outputs(6676) <= a and b;
    layer6_outputs(6677) <= b;
    layer6_outputs(6678) <= a xor b;
    layer6_outputs(6679) <= a;
    layer6_outputs(6680) <= a and b;
    layer6_outputs(6681) <= not a;
    layer6_outputs(6682) <= not (a and b);
    layer6_outputs(6683) <= not (a or b);
    layer6_outputs(6684) <= a or b;
    layer6_outputs(6685) <= not (a xor b);
    layer6_outputs(6686) <= not (a or b);
    layer6_outputs(6687) <= not a;
    layer6_outputs(6688) <= a and b;
    layer6_outputs(6689) <= a and b;
    layer6_outputs(6690) <= '1';
    layer6_outputs(6691) <= not (a and b);
    layer6_outputs(6692) <= not b;
    layer6_outputs(6693) <= not a;
    layer6_outputs(6694) <= not b or a;
    layer6_outputs(6695) <= b;
    layer6_outputs(6696) <= not a or b;
    layer6_outputs(6697) <= not a;
    layer6_outputs(6698) <= b;
    layer6_outputs(6699) <= not b or a;
    layer6_outputs(6700) <= not (a xor b);
    layer6_outputs(6701) <= not a;
    layer6_outputs(6702) <= not b;
    layer6_outputs(6703) <= a xor b;
    layer6_outputs(6704) <= not (a and b);
    layer6_outputs(6705) <= b and not a;
    layer6_outputs(6706) <= a and not b;
    layer6_outputs(6707) <= a or b;
    layer6_outputs(6708) <= not a or b;
    layer6_outputs(6709) <= not a;
    layer6_outputs(6710) <= b;
    layer6_outputs(6711) <= not b;
    layer6_outputs(6712) <= not (a or b);
    layer6_outputs(6713) <= a or b;
    layer6_outputs(6714) <= not a;
    layer6_outputs(6715) <= a or b;
    layer6_outputs(6716) <= not b;
    layer6_outputs(6717) <= a;
    layer6_outputs(6718) <= not (a and b);
    layer6_outputs(6719) <= b;
    layer6_outputs(6720) <= not a or b;
    layer6_outputs(6721) <= not (a or b);
    layer6_outputs(6722) <= not a;
    layer6_outputs(6723) <= not (a or b);
    layer6_outputs(6724) <= a and b;
    layer6_outputs(6725) <= b;
    layer6_outputs(6726) <= not b;
    layer6_outputs(6727) <= not a or b;
    layer6_outputs(6728) <= not b;
    layer6_outputs(6729) <= a and not b;
    layer6_outputs(6730) <= a;
    layer6_outputs(6731) <= a;
    layer6_outputs(6732) <= b;
    layer6_outputs(6733) <= not (a or b);
    layer6_outputs(6734) <= not (a or b);
    layer6_outputs(6735) <= not a or b;
    layer6_outputs(6736) <= a;
    layer6_outputs(6737) <= not b;
    layer6_outputs(6738) <= a;
    layer6_outputs(6739) <= a or b;
    layer6_outputs(6740) <= a and b;
    layer6_outputs(6741) <= a and not b;
    layer6_outputs(6742) <= a and not b;
    layer6_outputs(6743) <= not (a or b);
    layer6_outputs(6744) <= a;
    layer6_outputs(6745) <= not b;
    layer6_outputs(6746) <= a xor b;
    layer6_outputs(6747) <= a and not b;
    layer6_outputs(6748) <= '0';
    layer6_outputs(6749) <= not a;
    layer6_outputs(6750) <= b;
    layer6_outputs(6751) <= not b;
    layer6_outputs(6752) <= a;
    layer6_outputs(6753) <= a or b;
    layer6_outputs(6754) <= '0';
    layer6_outputs(6755) <= a;
    layer6_outputs(6756) <= a or b;
    layer6_outputs(6757) <= a xor b;
    layer6_outputs(6758) <= a xor b;
    layer6_outputs(6759) <= a;
    layer6_outputs(6760) <= not a;
    layer6_outputs(6761) <= not (a or b);
    layer6_outputs(6762) <= not b or a;
    layer6_outputs(6763) <= b;
    layer6_outputs(6764) <= not (a and b);
    layer6_outputs(6765) <= not (a and b);
    layer6_outputs(6766) <= not (a or b);
    layer6_outputs(6767) <= not a;
    layer6_outputs(6768) <= not b;
    layer6_outputs(6769) <= not a;
    layer6_outputs(6770) <= b;
    layer6_outputs(6771) <= not b or a;
    layer6_outputs(6772) <= not a or b;
    layer6_outputs(6773) <= not b or a;
    layer6_outputs(6774) <= not b;
    layer6_outputs(6775) <= not b;
    layer6_outputs(6776) <= not (a xor b);
    layer6_outputs(6777) <= a or b;
    layer6_outputs(6778) <= not a;
    layer6_outputs(6779) <= not (a or b);
    layer6_outputs(6780) <= a and not b;
    layer6_outputs(6781) <= not a;
    layer6_outputs(6782) <= not b;
    layer6_outputs(6783) <= b;
    layer6_outputs(6784) <= not b;
    layer6_outputs(6785) <= not a;
    layer6_outputs(6786) <= not (a and b);
    layer6_outputs(6787) <= not b;
    layer6_outputs(6788) <= not b or a;
    layer6_outputs(6789) <= not b;
    layer6_outputs(6790) <= not a;
    layer6_outputs(6791) <= not a;
    layer6_outputs(6792) <= a xor b;
    layer6_outputs(6793) <= not (a or b);
    layer6_outputs(6794) <= a and not b;
    layer6_outputs(6795) <= a;
    layer6_outputs(6796) <= b;
    layer6_outputs(6797) <= not b;
    layer6_outputs(6798) <= not b;
    layer6_outputs(6799) <= a and b;
    layer6_outputs(6800) <= b;
    layer6_outputs(6801) <= not a;
    layer6_outputs(6802) <= not (a or b);
    layer6_outputs(6803) <= a and b;
    layer6_outputs(6804) <= a and not b;
    layer6_outputs(6805) <= not a;
    layer6_outputs(6806) <= not b;
    layer6_outputs(6807) <= not a;
    layer6_outputs(6808) <= not b;
    layer6_outputs(6809) <= not (a and b);
    layer6_outputs(6810) <= not (a xor b);
    layer6_outputs(6811) <= a and not b;
    layer6_outputs(6812) <= b;
    layer6_outputs(6813) <= a and not b;
    layer6_outputs(6814) <= a;
    layer6_outputs(6815) <= a;
    layer6_outputs(6816) <= b and not a;
    layer6_outputs(6817) <= not (a or b);
    layer6_outputs(6818) <= not b;
    layer6_outputs(6819) <= not b;
    layer6_outputs(6820) <= a;
    layer6_outputs(6821) <= a;
    layer6_outputs(6822) <= not b;
    layer6_outputs(6823) <= not (a or b);
    layer6_outputs(6824) <= b;
    layer6_outputs(6825) <= not a;
    layer6_outputs(6826) <= not a;
    layer6_outputs(6827) <= b;
    layer6_outputs(6828) <= b;
    layer6_outputs(6829) <= a;
    layer6_outputs(6830) <= b;
    layer6_outputs(6831) <= a and not b;
    layer6_outputs(6832) <= not (a and b);
    layer6_outputs(6833) <= not a or b;
    layer6_outputs(6834) <= a and b;
    layer6_outputs(6835) <= not b;
    layer6_outputs(6836) <= a xor b;
    layer6_outputs(6837) <= a;
    layer6_outputs(6838) <= b and not a;
    layer6_outputs(6839) <= not a or b;
    layer6_outputs(6840) <= not (a xor b);
    layer6_outputs(6841) <= not a or b;
    layer6_outputs(6842) <= not a;
    layer6_outputs(6843) <= not a;
    layer6_outputs(6844) <= not b;
    layer6_outputs(6845) <= b and not a;
    layer6_outputs(6846) <= a xor b;
    layer6_outputs(6847) <= not a;
    layer6_outputs(6848) <= not b;
    layer6_outputs(6849) <= b;
    layer6_outputs(6850) <= b and not a;
    layer6_outputs(6851) <= a;
    layer6_outputs(6852) <= a and b;
    layer6_outputs(6853) <= b;
    layer6_outputs(6854) <= not b or a;
    layer6_outputs(6855) <= not (a xor b);
    layer6_outputs(6856) <= a;
    layer6_outputs(6857) <= b;
    layer6_outputs(6858) <= not a or b;
    layer6_outputs(6859) <= not (a or b);
    layer6_outputs(6860) <= a;
    layer6_outputs(6861) <= not b;
    layer6_outputs(6862) <= not a;
    layer6_outputs(6863) <= a and b;
    layer6_outputs(6864) <= a;
    layer6_outputs(6865) <= b and not a;
    layer6_outputs(6866) <= not a;
    layer6_outputs(6867) <= not a or b;
    layer6_outputs(6868) <= not (a and b);
    layer6_outputs(6869) <= not a or b;
    layer6_outputs(6870) <= a or b;
    layer6_outputs(6871) <= '0';
    layer6_outputs(6872) <= a or b;
    layer6_outputs(6873) <= a or b;
    layer6_outputs(6874) <= a and b;
    layer6_outputs(6875) <= not a;
    layer6_outputs(6876) <= not a or b;
    layer6_outputs(6877) <= b;
    layer6_outputs(6878) <= not b;
    layer6_outputs(6879) <= b and not a;
    layer6_outputs(6880) <= not (a and b);
    layer6_outputs(6881) <= b;
    layer6_outputs(6882) <= not (a or b);
    layer6_outputs(6883) <= not (a xor b);
    layer6_outputs(6884) <= not a;
    layer6_outputs(6885) <= a;
    layer6_outputs(6886) <= not b;
    layer6_outputs(6887) <= a;
    layer6_outputs(6888) <= not (a and b);
    layer6_outputs(6889) <= not a;
    layer6_outputs(6890) <= not (a or b);
    layer6_outputs(6891) <= not (a xor b);
    layer6_outputs(6892) <= a;
    layer6_outputs(6893) <= b and not a;
    layer6_outputs(6894) <= not a or b;
    layer6_outputs(6895) <= b;
    layer6_outputs(6896) <= not b;
    layer6_outputs(6897) <= not b;
    layer6_outputs(6898) <= b;
    layer6_outputs(6899) <= '0';
    layer6_outputs(6900) <= a;
    layer6_outputs(6901) <= not (a or b);
    layer6_outputs(6902) <= a or b;
    layer6_outputs(6903) <= a and b;
    layer6_outputs(6904) <= a or b;
    layer6_outputs(6905) <= b and not a;
    layer6_outputs(6906) <= a;
    layer6_outputs(6907) <= a and not b;
    layer6_outputs(6908) <= not a;
    layer6_outputs(6909) <= a and not b;
    layer6_outputs(6910) <= not (a or b);
    layer6_outputs(6911) <= a xor b;
    layer6_outputs(6912) <= a or b;
    layer6_outputs(6913) <= a xor b;
    layer6_outputs(6914) <= a;
    layer6_outputs(6915) <= a or b;
    layer6_outputs(6916) <= a xor b;
    layer6_outputs(6917) <= not b;
    layer6_outputs(6918) <= a xor b;
    layer6_outputs(6919) <= not b;
    layer6_outputs(6920) <= not b;
    layer6_outputs(6921) <= not a;
    layer6_outputs(6922) <= not b;
    layer6_outputs(6923) <= a xor b;
    layer6_outputs(6924) <= '0';
    layer6_outputs(6925) <= not a;
    layer6_outputs(6926) <= a and b;
    layer6_outputs(6927) <= a and not b;
    layer6_outputs(6928) <= not (a xor b);
    layer6_outputs(6929) <= a xor b;
    layer6_outputs(6930) <= a or b;
    layer6_outputs(6931) <= not a;
    layer6_outputs(6932) <= not b or a;
    layer6_outputs(6933) <= a;
    layer6_outputs(6934) <= b;
    layer6_outputs(6935) <= not b;
    layer6_outputs(6936) <= not b;
    layer6_outputs(6937) <= a;
    layer6_outputs(6938) <= not a;
    layer6_outputs(6939) <= not (a and b);
    layer6_outputs(6940) <= not b;
    layer6_outputs(6941) <= a;
    layer6_outputs(6942) <= not a;
    layer6_outputs(6943) <= not (a or b);
    layer6_outputs(6944) <= '0';
    layer6_outputs(6945) <= a and not b;
    layer6_outputs(6946) <= not b;
    layer6_outputs(6947) <= not (a xor b);
    layer6_outputs(6948) <= a and b;
    layer6_outputs(6949) <= not (a and b);
    layer6_outputs(6950) <= not (a or b);
    layer6_outputs(6951) <= b and not a;
    layer6_outputs(6952) <= not (a and b);
    layer6_outputs(6953) <= b;
    layer6_outputs(6954) <= b;
    layer6_outputs(6955) <= not b;
    layer6_outputs(6956) <= not b;
    layer6_outputs(6957) <= a and not b;
    layer6_outputs(6958) <= not b;
    layer6_outputs(6959) <= a or b;
    layer6_outputs(6960) <= not b;
    layer6_outputs(6961) <= not (a or b);
    layer6_outputs(6962) <= '1';
    layer6_outputs(6963) <= a and b;
    layer6_outputs(6964) <= not (a and b);
    layer6_outputs(6965) <= not b;
    layer6_outputs(6966) <= b and not a;
    layer6_outputs(6967) <= not (a or b);
    layer6_outputs(6968) <= not (a xor b);
    layer6_outputs(6969) <= not (a xor b);
    layer6_outputs(6970) <= a;
    layer6_outputs(6971) <= not b or a;
    layer6_outputs(6972) <= not a or b;
    layer6_outputs(6973) <= not b;
    layer6_outputs(6974) <= not (a xor b);
    layer6_outputs(6975) <= b and not a;
    layer6_outputs(6976) <= a and b;
    layer6_outputs(6977) <= a;
    layer6_outputs(6978) <= not b;
    layer6_outputs(6979) <= not b;
    layer6_outputs(6980) <= not b;
    layer6_outputs(6981) <= b;
    layer6_outputs(6982) <= not (a or b);
    layer6_outputs(6983) <= a or b;
    layer6_outputs(6984) <= a and not b;
    layer6_outputs(6985) <= b and not a;
    layer6_outputs(6986) <= b;
    layer6_outputs(6987) <= b;
    layer6_outputs(6988) <= b;
    layer6_outputs(6989) <= not (a or b);
    layer6_outputs(6990) <= not a;
    layer6_outputs(6991) <= not a;
    layer6_outputs(6992) <= not b;
    layer6_outputs(6993) <= not b;
    layer6_outputs(6994) <= not (a and b);
    layer6_outputs(6995) <= not (a or b);
    layer6_outputs(6996) <= not b;
    layer6_outputs(6997) <= a;
    layer6_outputs(6998) <= '0';
    layer6_outputs(6999) <= a and b;
    layer6_outputs(7000) <= not (a and b);
    layer6_outputs(7001) <= a;
    layer6_outputs(7002) <= b;
    layer6_outputs(7003) <= not b;
    layer6_outputs(7004) <= a and b;
    layer6_outputs(7005) <= a and b;
    layer6_outputs(7006) <= not (a xor b);
    layer6_outputs(7007) <= not (a xor b);
    layer6_outputs(7008) <= a;
    layer6_outputs(7009) <= b;
    layer6_outputs(7010) <= not b;
    layer6_outputs(7011) <= not b;
    layer6_outputs(7012) <= b;
    layer6_outputs(7013) <= not b or a;
    layer6_outputs(7014) <= a;
    layer6_outputs(7015) <= not a or b;
    layer6_outputs(7016) <= not (a xor b);
    layer6_outputs(7017) <= not b;
    layer6_outputs(7018) <= a xor b;
    layer6_outputs(7019) <= a;
    layer6_outputs(7020) <= not b;
    layer6_outputs(7021) <= not (a or b);
    layer6_outputs(7022) <= b;
    layer6_outputs(7023) <= not b;
    layer6_outputs(7024) <= not a;
    layer6_outputs(7025) <= a xor b;
    layer6_outputs(7026) <= a;
    layer6_outputs(7027) <= '1';
    layer6_outputs(7028) <= not b;
    layer6_outputs(7029) <= not (a xor b);
    layer6_outputs(7030) <= '0';
    layer6_outputs(7031) <= a xor b;
    layer6_outputs(7032) <= a xor b;
    layer6_outputs(7033) <= a xor b;
    layer6_outputs(7034) <= not b;
    layer6_outputs(7035) <= b;
    layer6_outputs(7036) <= a and not b;
    layer6_outputs(7037) <= b;
    layer6_outputs(7038) <= a xor b;
    layer6_outputs(7039) <= a xor b;
    layer6_outputs(7040) <= not b or a;
    layer6_outputs(7041) <= not b;
    layer6_outputs(7042) <= not b;
    layer6_outputs(7043) <= b and not a;
    layer6_outputs(7044) <= a and b;
    layer6_outputs(7045) <= '0';
    layer6_outputs(7046) <= a or b;
    layer6_outputs(7047) <= not a or b;
    layer6_outputs(7048) <= not a or b;
    layer6_outputs(7049) <= b;
    layer6_outputs(7050) <= not (a or b);
    layer6_outputs(7051) <= not a;
    layer6_outputs(7052) <= a;
    layer6_outputs(7053) <= a;
    layer6_outputs(7054) <= not a;
    layer6_outputs(7055) <= b and not a;
    layer6_outputs(7056) <= b;
    layer6_outputs(7057) <= a;
    layer6_outputs(7058) <= b;
    layer6_outputs(7059) <= a and not b;
    layer6_outputs(7060) <= a xor b;
    layer6_outputs(7061) <= b;
    layer6_outputs(7062) <= not (a xor b);
    layer6_outputs(7063) <= not a or b;
    layer6_outputs(7064) <= a;
    layer6_outputs(7065) <= not b;
    layer6_outputs(7066) <= not b;
    layer6_outputs(7067) <= '0';
    layer6_outputs(7068) <= not a or b;
    layer6_outputs(7069) <= not b or a;
    layer6_outputs(7070) <= a;
    layer6_outputs(7071) <= not b;
    layer6_outputs(7072) <= a;
    layer6_outputs(7073) <= not b;
    layer6_outputs(7074) <= not b;
    layer6_outputs(7075) <= '1';
    layer6_outputs(7076) <= not b;
    layer6_outputs(7077) <= '0';
    layer6_outputs(7078) <= not (a xor b);
    layer6_outputs(7079) <= a and not b;
    layer6_outputs(7080) <= not a or b;
    layer6_outputs(7081) <= a and not b;
    layer6_outputs(7082) <= not (a xor b);
    layer6_outputs(7083) <= b;
    layer6_outputs(7084) <= not a or b;
    layer6_outputs(7085) <= '0';
    layer6_outputs(7086) <= not (a or b);
    layer6_outputs(7087) <= not (a xor b);
    layer6_outputs(7088) <= a;
    layer6_outputs(7089) <= a;
    layer6_outputs(7090) <= b;
    layer6_outputs(7091) <= not b;
    layer6_outputs(7092) <= b;
    layer6_outputs(7093) <= a and not b;
    layer6_outputs(7094) <= a or b;
    layer6_outputs(7095) <= not b;
    layer6_outputs(7096) <= b;
    layer6_outputs(7097) <= not b;
    layer6_outputs(7098) <= a and b;
    layer6_outputs(7099) <= not a;
    layer6_outputs(7100) <= a;
    layer6_outputs(7101) <= a or b;
    layer6_outputs(7102) <= not b or a;
    layer6_outputs(7103) <= '0';
    layer6_outputs(7104) <= a and b;
    layer6_outputs(7105) <= not (a xor b);
    layer6_outputs(7106) <= b;
    layer6_outputs(7107) <= a;
    layer6_outputs(7108) <= b;
    layer6_outputs(7109) <= b;
    layer6_outputs(7110) <= not b;
    layer6_outputs(7111) <= a and b;
    layer6_outputs(7112) <= a or b;
    layer6_outputs(7113) <= a and b;
    layer6_outputs(7114) <= '0';
    layer6_outputs(7115) <= not (a or b);
    layer6_outputs(7116) <= not b or a;
    layer6_outputs(7117) <= not b;
    layer6_outputs(7118) <= b and not a;
    layer6_outputs(7119) <= b;
    layer6_outputs(7120) <= a xor b;
    layer6_outputs(7121) <= b;
    layer6_outputs(7122) <= not b or a;
    layer6_outputs(7123) <= a and b;
    layer6_outputs(7124) <= b and not a;
    layer6_outputs(7125) <= not b or a;
    layer6_outputs(7126) <= a or b;
    layer6_outputs(7127) <= a or b;
    layer6_outputs(7128) <= b;
    layer6_outputs(7129) <= a and b;
    layer6_outputs(7130) <= not (a or b);
    layer6_outputs(7131) <= '1';
    layer6_outputs(7132) <= a xor b;
    layer6_outputs(7133) <= not (a xor b);
    layer6_outputs(7134) <= not b;
    layer6_outputs(7135) <= not b;
    layer6_outputs(7136) <= not b or a;
    layer6_outputs(7137) <= a and not b;
    layer6_outputs(7138) <= a xor b;
    layer6_outputs(7139) <= b;
    layer6_outputs(7140) <= a;
    layer6_outputs(7141) <= not b or a;
    layer6_outputs(7142) <= a and not b;
    layer6_outputs(7143) <= not a;
    layer6_outputs(7144) <= not b;
    layer6_outputs(7145) <= b and not a;
    layer6_outputs(7146) <= b and not a;
    layer6_outputs(7147) <= a;
    layer6_outputs(7148) <= not (a xor b);
    layer6_outputs(7149) <= a;
    layer6_outputs(7150) <= not a or b;
    layer6_outputs(7151) <= not (a or b);
    layer6_outputs(7152) <= '0';
    layer6_outputs(7153) <= not b or a;
    layer6_outputs(7154) <= a or b;
    layer6_outputs(7155) <= a and not b;
    layer6_outputs(7156) <= not (a or b);
    layer6_outputs(7157) <= a and not b;
    layer6_outputs(7158) <= a or b;
    layer6_outputs(7159) <= not a;
    layer6_outputs(7160) <= not a or b;
    layer6_outputs(7161) <= b and not a;
    layer6_outputs(7162) <= a and b;
    layer6_outputs(7163) <= a xor b;
    layer6_outputs(7164) <= not a;
    layer6_outputs(7165) <= not (a xor b);
    layer6_outputs(7166) <= a;
    layer6_outputs(7167) <= not a;
    layer6_outputs(7168) <= a xor b;
    layer6_outputs(7169) <= b and not a;
    layer6_outputs(7170) <= not b;
    layer6_outputs(7171) <= not (a xor b);
    layer6_outputs(7172) <= a;
    layer6_outputs(7173) <= not a;
    layer6_outputs(7174) <= b;
    layer6_outputs(7175) <= b and not a;
    layer6_outputs(7176) <= a and b;
    layer6_outputs(7177) <= not a;
    layer6_outputs(7178) <= a;
    layer6_outputs(7179) <= a xor b;
    layer6_outputs(7180) <= not (a and b);
    layer6_outputs(7181) <= not (a and b);
    layer6_outputs(7182) <= not a;
    layer6_outputs(7183) <= a;
    layer6_outputs(7184) <= not a or b;
    layer6_outputs(7185) <= not (a and b);
    layer6_outputs(7186) <= not (a xor b);
    layer6_outputs(7187) <= not a;
    layer6_outputs(7188) <= b;
    layer6_outputs(7189) <= b;
    layer6_outputs(7190) <= not (a or b);
    layer6_outputs(7191) <= not (a and b);
    layer6_outputs(7192) <= b and not a;
    layer6_outputs(7193) <= not a;
    layer6_outputs(7194) <= a or b;
    layer6_outputs(7195) <= not a;
    layer6_outputs(7196) <= not b or a;
    layer6_outputs(7197) <= not b;
    layer6_outputs(7198) <= b and not a;
    layer6_outputs(7199) <= b;
    layer6_outputs(7200) <= not b;
    layer6_outputs(7201) <= a xor b;
    layer6_outputs(7202) <= a and b;
    layer6_outputs(7203) <= '0';
    layer6_outputs(7204) <= b and not a;
    layer6_outputs(7205) <= a xor b;
    layer6_outputs(7206) <= not b;
    layer6_outputs(7207) <= a xor b;
    layer6_outputs(7208) <= a;
    layer6_outputs(7209) <= not (a xor b);
    layer6_outputs(7210) <= not a;
    layer6_outputs(7211) <= not b or a;
    layer6_outputs(7212) <= b;
    layer6_outputs(7213) <= a and b;
    layer6_outputs(7214) <= a;
    layer6_outputs(7215) <= '0';
    layer6_outputs(7216) <= a or b;
    layer6_outputs(7217) <= b;
    layer6_outputs(7218) <= not (a and b);
    layer6_outputs(7219) <= a and b;
    layer6_outputs(7220) <= '0';
    layer6_outputs(7221) <= a xor b;
    layer6_outputs(7222) <= a;
    layer6_outputs(7223) <= not (a xor b);
    layer6_outputs(7224) <= not b;
    layer6_outputs(7225) <= a and not b;
    layer6_outputs(7226) <= b;
    layer6_outputs(7227) <= not a;
    layer6_outputs(7228) <= a and b;
    layer6_outputs(7229) <= b and not a;
    layer6_outputs(7230) <= b and not a;
    layer6_outputs(7231) <= not (a and b);
    layer6_outputs(7232) <= not b or a;
    layer6_outputs(7233) <= not b;
    layer6_outputs(7234) <= a and b;
    layer6_outputs(7235) <= a and b;
    layer6_outputs(7236) <= a;
    layer6_outputs(7237) <= not b or a;
    layer6_outputs(7238) <= '0';
    layer6_outputs(7239) <= not b;
    layer6_outputs(7240) <= b;
    layer6_outputs(7241) <= b and not a;
    layer6_outputs(7242) <= a or b;
    layer6_outputs(7243) <= a xor b;
    layer6_outputs(7244) <= a and b;
    layer6_outputs(7245) <= not (a or b);
    layer6_outputs(7246) <= b;
    layer6_outputs(7247) <= '1';
    layer6_outputs(7248) <= a;
    layer6_outputs(7249) <= a xor b;
    layer6_outputs(7250) <= not a;
    layer6_outputs(7251) <= not (a or b);
    layer6_outputs(7252) <= not a or b;
    layer6_outputs(7253) <= a and b;
    layer6_outputs(7254) <= not b or a;
    layer6_outputs(7255) <= not b or a;
    layer6_outputs(7256) <= b;
    layer6_outputs(7257) <= not a;
    layer6_outputs(7258) <= not b;
    layer6_outputs(7259) <= not b;
    layer6_outputs(7260) <= not a or b;
    layer6_outputs(7261) <= a;
    layer6_outputs(7262) <= b and not a;
    layer6_outputs(7263) <= b;
    layer6_outputs(7264) <= a xor b;
    layer6_outputs(7265) <= a or b;
    layer6_outputs(7266) <= '1';
    layer6_outputs(7267) <= b;
    layer6_outputs(7268) <= a and b;
    layer6_outputs(7269) <= not a;
    layer6_outputs(7270) <= a and b;
    layer6_outputs(7271) <= not (a and b);
    layer6_outputs(7272) <= not b;
    layer6_outputs(7273) <= a xor b;
    layer6_outputs(7274) <= not b or a;
    layer6_outputs(7275) <= b;
    layer6_outputs(7276) <= not (a xor b);
    layer6_outputs(7277) <= b;
    layer6_outputs(7278) <= not b;
    layer6_outputs(7279) <= '1';
    layer6_outputs(7280) <= b and not a;
    layer6_outputs(7281) <= b;
    layer6_outputs(7282) <= not a;
    layer6_outputs(7283) <= a;
    layer6_outputs(7284) <= not b;
    layer6_outputs(7285) <= a;
    layer6_outputs(7286) <= a xor b;
    layer6_outputs(7287) <= not (a and b);
    layer6_outputs(7288) <= '0';
    layer6_outputs(7289) <= b and not a;
    layer6_outputs(7290) <= not b;
    layer6_outputs(7291) <= a or b;
    layer6_outputs(7292) <= b;
    layer6_outputs(7293) <= a and b;
    layer6_outputs(7294) <= '1';
    layer6_outputs(7295) <= not a or b;
    layer6_outputs(7296) <= a;
    layer6_outputs(7297) <= not (a and b);
    layer6_outputs(7298) <= not b;
    layer6_outputs(7299) <= not a;
    layer6_outputs(7300) <= a and not b;
    layer6_outputs(7301) <= not (a xor b);
    layer6_outputs(7302) <= not b;
    layer6_outputs(7303) <= not a;
    layer6_outputs(7304) <= not b;
    layer6_outputs(7305) <= '0';
    layer6_outputs(7306) <= a or b;
    layer6_outputs(7307) <= a xor b;
    layer6_outputs(7308) <= a and not b;
    layer6_outputs(7309) <= b;
    layer6_outputs(7310) <= a;
    layer6_outputs(7311) <= not (a and b);
    layer6_outputs(7312) <= a and b;
    layer6_outputs(7313) <= not (a and b);
    layer6_outputs(7314) <= a and b;
    layer6_outputs(7315) <= not (a xor b);
    layer6_outputs(7316) <= not (a xor b);
    layer6_outputs(7317) <= a xor b;
    layer6_outputs(7318) <= not a;
    layer6_outputs(7319) <= a;
    layer6_outputs(7320) <= not a;
    layer6_outputs(7321) <= not a or b;
    layer6_outputs(7322) <= not a;
    layer6_outputs(7323) <= b and not a;
    layer6_outputs(7324) <= not b;
    layer6_outputs(7325) <= not a;
    layer6_outputs(7326) <= not a;
    layer6_outputs(7327) <= b;
    layer6_outputs(7328) <= not a;
    layer6_outputs(7329) <= a xor b;
    layer6_outputs(7330) <= a;
    layer6_outputs(7331) <= a or b;
    layer6_outputs(7332) <= a and b;
    layer6_outputs(7333) <= not a;
    layer6_outputs(7334) <= not (a xor b);
    layer6_outputs(7335) <= not b;
    layer6_outputs(7336) <= not b;
    layer6_outputs(7337) <= not (a or b);
    layer6_outputs(7338) <= '1';
    layer6_outputs(7339) <= not (a xor b);
    layer6_outputs(7340) <= b;
    layer6_outputs(7341) <= not (a or b);
    layer6_outputs(7342) <= a or b;
    layer6_outputs(7343) <= not b;
    layer6_outputs(7344) <= a;
    layer6_outputs(7345) <= a;
    layer6_outputs(7346) <= not a or b;
    layer6_outputs(7347) <= a;
    layer6_outputs(7348) <= a and b;
    layer6_outputs(7349) <= a xor b;
    layer6_outputs(7350) <= a;
    layer6_outputs(7351) <= not (a and b);
    layer6_outputs(7352) <= '0';
    layer6_outputs(7353) <= not a;
    layer6_outputs(7354) <= not b or a;
    layer6_outputs(7355) <= not b;
    layer6_outputs(7356) <= b;
    layer6_outputs(7357) <= not (a and b);
    layer6_outputs(7358) <= not b or a;
    layer6_outputs(7359) <= not (a and b);
    layer6_outputs(7360) <= '1';
    layer6_outputs(7361) <= b and not a;
    layer6_outputs(7362) <= not (a xor b);
    layer6_outputs(7363) <= not a or b;
    layer6_outputs(7364) <= '0';
    layer6_outputs(7365) <= not b;
    layer6_outputs(7366) <= b;
    layer6_outputs(7367) <= not (a xor b);
    layer6_outputs(7368) <= not a or b;
    layer6_outputs(7369) <= not b or a;
    layer6_outputs(7370) <= b and not a;
    layer6_outputs(7371) <= not b or a;
    layer6_outputs(7372) <= not a or b;
    layer6_outputs(7373) <= b;
    layer6_outputs(7374) <= '1';
    layer6_outputs(7375) <= b;
    layer6_outputs(7376) <= a;
    layer6_outputs(7377) <= b and not a;
    layer6_outputs(7378) <= not (a or b);
    layer6_outputs(7379) <= not b;
    layer6_outputs(7380) <= not a;
    layer6_outputs(7381) <= a;
    layer6_outputs(7382) <= not a;
    layer6_outputs(7383) <= not a or b;
    layer6_outputs(7384) <= a and b;
    layer6_outputs(7385) <= a and b;
    layer6_outputs(7386) <= not b or a;
    layer6_outputs(7387) <= b;
    layer6_outputs(7388) <= a and not b;
    layer6_outputs(7389) <= a xor b;
    layer6_outputs(7390) <= not a or b;
    layer6_outputs(7391) <= a xor b;
    layer6_outputs(7392) <= not a;
    layer6_outputs(7393) <= a xor b;
    layer6_outputs(7394) <= a and b;
    layer6_outputs(7395) <= '0';
    layer6_outputs(7396) <= not a or b;
    layer6_outputs(7397) <= not b;
    layer6_outputs(7398) <= not (a xor b);
    layer6_outputs(7399) <= a and not b;
    layer6_outputs(7400) <= not a;
    layer6_outputs(7401) <= b;
    layer6_outputs(7402) <= not (a and b);
    layer6_outputs(7403) <= a;
    layer6_outputs(7404) <= not a;
    layer6_outputs(7405) <= b and not a;
    layer6_outputs(7406) <= not b;
    layer6_outputs(7407) <= not a or b;
    layer6_outputs(7408) <= a and not b;
    layer6_outputs(7409) <= a and not b;
    layer6_outputs(7410) <= not (a xor b);
    layer6_outputs(7411) <= not b;
    layer6_outputs(7412) <= b;
    layer6_outputs(7413) <= not b or a;
    layer6_outputs(7414) <= a and not b;
    layer6_outputs(7415) <= b;
    layer6_outputs(7416) <= not b;
    layer6_outputs(7417) <= a xor b;
    layer6_outputs(7418) <= a and b;
    layer6_outputs(7419) <= not a;
    layer6_outputs(7420) <= not a or b;
    layer6_outputs(7421) <= b;
    layer6_outputs(7422) <= not (a and b);
    layer6_outputs(7423) <= b;
    layer6_outputs(7424) <= not b or a;
    layer6_outputs(7425) <= b;
    layer6_outputs(7426) <= b and not a;
    layer6_outputs(7427) <= a and b;
    layer6_outputs(7428) <= a or b;
    layer6_outputs(7429) <= '0';
    layer6_outputs(7430) <= b and not a;
    layer6_outputs(7431) <= not b;
    layer6_outputs(7432) <= a and b;
    layer6_outputs(7433) <= a xor b;
    layer6_outputs(7434) <= '0';
    layer6_outputs(7435) <= b;
    layer6_outputs(7436) <= not b;
    layer6_outputs(7437) <= a or b;
    layer6_outputs(7438) <= not (a or b);
    layer6_outputs(7439) <= not (a or b);
    layer6_outputs(7440) <= not (a xor b);
    layer6_outputs(7441) <= not (a or b);
    layer6_outputs(7442) <= not b;
    layer6_outputs(7443) <= a;
    layer6_outputs(7444) <= a and b;
    layer6_outputs(7445) <= not b;
    layer6_outputs(7446) <= not b;
    layer6_outputs(7447) <= not b;
    layer6_outputs(7448) <= b;
    layer6_outputs(7449) <= not a;
    layer6_outputs(7450) <= not (a xor b);
    layer6_outputs(7451) <= a;
    layer6_outputs(7452) <= not (a and b);
    layer6_outputs(7453) <= not (a or b);
    layer6_outputs(7454) <= not b;
    layer6_outputs(7455) <= not a;
    layer6_outputs(7456) <= b;
    layer6_outputs(7457) <= not a or b;
    layer6_outputs(7458) <= not (a or b);
    layer6_outputs(7459) <= not b;
    layer6_outputs(7460) <= a or b;
    layer6_outputs(7461) <= '0';
    layer6_outputs(7462) <= not a;
    layer6_outputs(7463) <= not (a or b);
    layer6_outputs(7464) <= a;
    layer6_outputs(7465) <= a and b;
    layer6_outputs(7466) <= not (a and b);
    layer6_outputs(7467) <= a and not b;
    layer6_outputs(7468) <= b and not a;
    layer6_outputs(7469) <= b and not a;
    layer6_outputs(7470) <= not (a xor b);
    layer6_outputs(7471) <= not (a and b);
    layer6_outputs(7472) <= b and not a;
    layer6_outputs(7473) <= not (a xor b);
    layer6_outputs(7474) <= a;
    layer6_outputs(7475) <= not b;
    layer6_outputs(7476) <= not b or a;
    layer6_outputs(7477) <= not a;
    layer6_outputs(7478) <= b;
    layer6_outputs(7479) <= not (a or b);
    layer6_outputs(7480) <= b and not a;
    layer6_outputs(7481) <= b;
    layer6_outputs(7482) <= b;
    layer6_outputs(7483) <= a;
    layer6_outputs(7484) <= b and not a;
    layer6_outputs(7485) <= a or b;
    layer6_outputs(7486) <= '0';
    layer6_outputs(7487) <= a or b;
    layer6_outputs(7488) <= not b;
    layer6_outputs(7489) <= b;
    layer6_outputs(7490) <= b and not a;
    layer6_outputs(7491) <= not (a or b);
    layer6_outputs(7492) <= not (a and b);
    layer6_outputs(7493) <= not (a xor b);
    layer6_outputs(7494) <= b;
    layer6_outputs(7495) <= a and b;
    layer6_outputs(7496) <= not a;
    layer6_outputs(7497) <= a or b;
    layer6_outputs(7498) <= not a;
    layer6_outputs(7499) <= not (a xor b);
    layer6_outputs(7500) <= b;
    layer6_outputs(7501) <= b;
    layer6_outputs(7502) <= not b or a;
    layer6_outputs(7503) <= a;
    layer6_outputs(7504) <= not b or a;
    layer6_outputs(7505) <= a and b;
    layer6_outputs(7506) <= '0';
    layer6_outputs(7507) <= a or b;
    layer6_outputs(7508) <= a;
    layer6_outputs(7509) <= '1';
    layer6_outputs(7510) <= not a;
    layer6_outputs(7511) <= a or b;
    layer6_outputs(7512) <= a;
    layer6_outputs(7513) <= a or b;
    layer6_outputs(7514) <= not (a or b);
    layer6_outputs(7515) <= b and not a;
    layer6_outputs(7516) <= not b or a;
    layer6_outputs(7517) <= not (a xor b);
    layer6_outputs(7518) <= not (a and b);
    layer6_outputs(7519) <= not a;
    layer6_outputs(7520) <= not (a or b);
    layer6_outputs(7521) <= not b;
    layer6_outputs(7522) <= b;
    layer6_outputs(7523) <= a xor b;
    layer6_outputs(7524) <= not a or b;
    layer6_outputs(7525) <= a xor b;
    layer6_outputs(7526) <= not a;
    layer6_outputs(7527) <= not a;
    layer6_outputs(7528) <= not (a and b);
    layer6_outputs(7529) <= not (a or b);
    layer6_outputs(7530) <= b;
    layer6_outputs(7531) <= a;
    layer6_outputs(7532) <= a;
    layer6_outputs(7533) <= b;
    layer6_outputs(7534) <= not (a xor b);
    layer6_outputs(7535) <= a or b;
    layer6_outputs(7536) <= b;
    layer6_outputs(7537) <= not b or a;
    layer6_outputs(7538) <= a or b;
    layer6_outputs(7539) <= a and not b;
    layer6_outputs(7540) <= not b;
    layer6_outputs(7541) <= not b;
    layer6_outputs(7542) <= not (a or b);
    layer6_outputs(7543) <= a xor b;
    layer6_outputs(7544) <= not b;
    layer6_outputs(7545) <= '0';
    layer6_outputs(7546) <= not a or b;
    layer6_outputs(7547) <= a and b;
    layer6_outputs(7548) <= a and b;
    layer6_outputs(7549) <= not a;
    layer6_outputs(7550) <= not a;
    layer6_outputs(7551) <= not (a xor b);
    layer6_outputs(7552) <= b and not a;
    layer6_outputs(7553) <= not (a and b);
    layer6_outputs(7554) <= a and b;
    layer6_outputs(7555) <= not a;
    layer6_outputs(7556) <= not b;
    layer6_outputs(7557) <= not b;
    layer6_outputs(7558) <= a or b;
    layer6_outputs(7559) <= a and b;
    layer6_outputs(7560) <= not b;
    layer6_outputs(7561) <= a xor b;
    layer6_outputs(7562) <= a and b;
    layer6_outputs(7563) <= not a or b;
    layer6_outputs(7564) <= b and not a;
    layer6_outputs(7565) <= a;
    layer6_outputs(7566) <= not a;
    layer6_outputs(7567) <= b;
    layer6_outputs(7568) <= a;
    layer6_outputs(7569) <= not a;
    layer6_outputs(7570) <= not b or a;
    layer6_outputs(7571) <= a or b;
    layer6_outputs(7572) <= b and not a;
    layer6_outputs(7573) <= a xor b;
    layer6_outputs(7574) <= not (a xor b);
    layer6_outputs(7575) <= not b;
    layer6_outputs(7576) <= a and b;
    layer6_outputs(7577) <= not b;
    layer6_outputs(7578) <= not b or a;
    layer6_outputs(7579) <= not a or b;
    layer6_outputs(7580) <= b and not a;
    layer6_outputs(7581) <= a or b;
    layer6_outputs(7582) <= '0';
    layer6_outputs(7583) <= not (a and b);
    layer6_outputs(7584) <= a and b;
    layer6_outputs(7585) <= not b or a;
    layer6_outputs(7586) <= a xor b;
    layer6_outputs(7587) <= a or b;
    layer6_outputs(7588) <= a or b;
    layer6_outputs(7589) <= not b or a;
    layer6_outputs(7590) <= b and not a;
    layer6_outputs(7591) <= '0';
    layer6_outputs(7592) <= not (a or b);
    layer6_outputs(7593) <= not b;
    layer6_outputs(7594) <= b and not a;
    layer6_outputs(7595) <= b and not a;
    layer6_outputs(7596) <= '1';
    layer6_outputs(7597) <= not b;
    layer6_outputs(7598) <= not b;
    layer6_outputs(7599) <= not a or b;
    layer6_outputs(7600) <= a and not b;
    layer6_outputs(7601) <= a xor b;
    layer6_outputs(7602) <= a and b;
    layer6_outputs(7603) <= b;
    layer6_outputs(7604) <= b;
    layer6_outputs(7605) <= a and not b;
    layer6_outputs(7606) <= b;
    layer6_outputs(7607) <= not b;
    layer6_outputs(7608) <= not (a and b);
    layer6_outputs(7609) <= a and b;
    layer6_outputs(7610) <= not a or b;
    layer6_outputs(7611) <= b and not a;
    layer6_outputs(7612) <= '0';
    layer6_outputs(7613) <= a xor b;
    layer6_outputs(7614) <= a and b;
    layer6_outputs(7615) <= not b;
    layer6_outputs(7616) <= b;
    layer6_outputs(7617) <= not (a and b);
    layer6_outputs(7618) <= not a or b;
    layer6_outputs(7619) <= not (a and b);
    layer6_outputs(7620) <= not b or a;
    layer6_outputs(7621) <= not (a and b);
    layer6_outputs(7622) <= a and not b;
    layer6_outputs(7623) <= a and b;
    layer6_outputs(7624) <= not (a xor b);
    layer6_outputs(7625) <= a;
    layer6_outputs(7626) <= not a or b;
    layer6_outputs(7627) <= not a;
    layer6_outputs(7628) <= a;
    layer6_outputs(7629) <= not (a and b);
    layer6_outputs(7630) <= a and not b;
    layer6_outputs(7631) <= not (a and b);
    layer6_outputs(7632) <= '0';
    layer6_outputs(7633) <= b;
    layer6_outputs(7634) <= a xor b;
    layer6_outputs(7635) <= not a;
    layer6_outputs(7636) <= a;
    layer6_outputs(7637) <= not a;
    layer6_outputs(7638) <= not (a xor b);
    layer6_outputs(7639) <= not a;
    layer6_outputs(7640) <= not b or a;
    layer6_outputs(7641) <= not b or a;
    layer6_outputs(7642) <= not a;
    layer6_outputs(7643) <= not a or b;
    layer6_outputs(7644) <= a;
    layer6_outputs(7645) <= b;
    layer6_outputs(7646) <= not b or a;
    layer6_outputs(7647) <= a xor b;
    layer6_outputs(7648) <= not (a and b);
    layer6_outputs(7649) <= not (a or b);
    layer6_outputs(7650) <= b;
    layer6_outputs(7651) <= not a;
    layer6_outputs(7652) <= a or b;
    layer6_outputs(7653) <= not (a xor b);
    layer6_outputs(7654) <= not a or b;
    layer6_outputs(7655) <= a xor b;
    layer6_outputs(7656) <= not (a xor b);
    layer6_outputs(7657) <= a xor b;
    layer6_outputs(7658) <= '0';
    layer6_outputs(7659) <= a and not b;
    layer6_outputs(7660) <= b;
    layer6_outputs(7661) <= not a or b;
    layer6_outputs(7662) <= not (a or b);
    layer6_outputs(7663) <= not a;
    layer6_outputs(7664) <= b;
    layer6_outputs(7665) <= not a or b;
    layer6_outputs(7666) <= not a;
    layer6_outputs(7667) <= a and b;
    layer6_outputs(7668) <= a xor b;
    layer6_outputs(7669) <= not b or a;
    layer6_outputs(7670) <= not (a and b);
    layer6_outputs(7671) <= not b or a;
    layer6_outputs(7672) <= not a;
    layer6_outputs(7673) <= not b;
    layer6_outputs(7674) <= a and not b;
    layer6_outputs(7675) <= a xor b;
    layer6_outputs(7676) <= a;
    layer6_outputs(7677) <= a or b;
    layer6_outputs(7678) <= not a;
    layer6_outputs(7679) <= '0';
    layer7_outputs(0) <= not a;
    layer7_outputs(1) <= not (a or b);
    layer7_outputs(2) <= a and not b;
    layer7_outputs(3) <= not (a xor b);
    layer7_outputs(4) <= not (a or b);
    layer7_outputs(5) <= a and b;
    layer7_outputs(6) <= not a;
    layer7_outputs(7) <= a;
    layer7_outputs(8) <= '0';
    layer7_outputs(9) <= a or b;
    layer7_outputs(10) <= not b;
    layer7_outputs(11) <= b;
    layer7_outputs(12) <= not a;
    layer7_outputs(13) <= not b;
    layer7_outputs(14) <= not b;
    layer7_outputs(15) <= not (a or b);
    layer7_outputs(16) <= not a;
    layer7_outputs(17) <= not a;
    layer7_outputs(18) <= a xor b;
    layer7_outputs(19) <= not b;
    layer7_outputs(20) <= b;
    layer7_outputs(21) <= b;
    layer7_outputs(22) <= not (a and b);
    layer7_outputs(23) <= a xor b;
    layer7_outputs(24) <= not a;
    layer7_outputs(25) <= not (a or b);
    layer7_outputs(26) <= not a;
    layer7_outputs(27) <= not b;
    layer7_outputs(28) <= b;
    layer7_outputs(29) <= not (a xor b);
    layer7_outputs(30) <= a or b;
    layer7_outputs(31) <= not (a or b);
    layer7_outputs(32) <= not b;
    layer7_outputs(33) <= not (a xor b);
    layer7_outputs(34) <= b;
    layer7_outputs(35) <= b;
    layer7_outputs(36) <= not b or a;
    layer7_outputs(37) <= not a;
    layer7_outputs(38) <= not (a or b);
    layer7_outputs(39) <= a and b;
    layer7_outputs(40) <= not (a and b);
    layer7_outputs(41) <= not b;
    layer7_outputs(42) <= not (a and b);
    layer7_outputs(43) <= '1';
    layer7_outputs(44) <= b;
    layer7_outputs(45) <= not a;
    layer7_outputs(46) <= not b or a;
    layer7_outputs(47) <= not b;
    layer7_outputs(48) <= not (a xor b);
    layer7_outputs(49) <= a;
    layer7_outputs(50) <= b;
    layer7_outputs(51) <= not (a and b);
    layer7_outputs(52) <= not (a and b);
    layer7_outputs(53) <= a or b;
    layer7_outputs(54) <= b;
    layer7_outputs(55) <= not b or a;
    layer7_outputs(56) <= not b or a;
    layer7_outputs(57) <= a;
    layer7_outputs(58) <= b;
    layer7_outputs(59) <= not (a or b);
    layer7_outputs(60) <= b;
    layer7_outputs(61) <= not (a xor b);
    layer7_outputs(62) <= a xor b;
    layer7_outputs(63) <= a and b;
    layer7_outputs(64) <= not (a xor b);
    layer7_outputs(65) <= not (a or b);
    layer7_outputs(66) <= not a;
    layer7_outputs(67) <= a xor b;
    layer7_outputs(68) <= b and not a;
    layer7_outputs(69) <= b;
    layer7_outputs(70) <= a and b;
    layer7_outputs(71) <= not b;
    layer7_outputs(72) <= a and b;
    layer7_outputs(73) <= b;
    layer7_outputs(74) <= b;
    layer7_outputs(75) <= b and not a;
    layer7_outputs(76) <= a;
    layer7_outputs(77) <= not a or b;
    layer7_outputs(78) <= not a;
    layer7_outputs(79) <= not a;
    layer7_outputs(80) <= a and not b;
    layer7_outputs(81) <= b;
    layer7_outputs(82) <= b and not a;
    layer7_outputs(83) <= a;
    layer7_outputs(84) <= a and not b;
    layer7_outputs(85) <= b;
    layer7_outputs(86) <= not (a or b);
    layer7_outputs(87) <= not (a xor b);
    layer7_outputs(88) <= '0';
    layer7_outputs(89) <= a;
    layer7_outputs(90) <= not b;
    layer7_outputs(91) <= not a or b;
    layer7_outputs(92) <= not (a xor b);
    layer7_outputs(93) <= not b;
    layer7_outputs(94) <= not b or a;
    layer7_outputs(95) <= not b or a;
    layer7_outputs(96) <= not b or a;
    layer7_outputs(97) <= a;
    layer7_outputs(98) <= not (a xor b);
    layer7_outputs(99) <= not b or a;
    layer7_outputs(100) <= not (a or b);
    layer7_outputs(101) <= a and b;
    layer7_outputs(102) <= a or b;
    layer7_outputs(103) <= a xor b;
    layer7_outputs(104) <= '1';
    layer7_outputs(105) <= '1';
    layer7_outputs(106) <= a and not b;
    layer7_outputs(107) <= not a;
    layer7_outputs(108) <= not (a xor b);
    layer7_outputs(109) <= not b;
    layer7_outputs(110) <= b;
    layer7_outputs(111) <= a and b;
    layer7_outputs(112) <= a and b;
    layer7_outputs(113) <= b;
    layer7_outputs(114) <= not a or b;
    layer7_outputs(115) <= not a;
    layer7_outputs(116) <= a xor b;
    layer7_outputs(117) <= a;
    layer7_outputs(118) <= not b;
    layer7_outputs(119) <= not a;
    layer7_outputs(120) <= not (a xor b);
    layer7_outputs(121) <= not (a or b);
    layer7_outputs(122) <= not a;
    layer7_outputs(123) <= a and b;
    layer7_outputs(124) <= b and not a;
    layer7_outputs(125) <= not a;
    layer7_outputs(126) <= not b;
    layer7_outputs(127) <= a or b;
    layer7_outputs(128) <= not (a and b);
    layer7_outputs(129) <= not b or a;
    layer7_outputs(130) <= b;
    layer7_outputs(131) <= a xor b;
    layer7_outputs(132) <= not a;
    layer7_outputs(133) <= not b or a;
    layer7_outputs(134) <= b and not a;
    layer7_outputs(135) <= b;
    layer7_outputs(136) <= b and not a;
    layer7_outputs(137) <= not a;
    layer7_outputs(138) <= '0';
    layer7_outputs(139) <= a and b;
    layer7_outputs(140) <= a and not b;
    layer7_outputs(141) <= a and not b;
    layer7_outputs(142) <= b and not a;
    layer7_outputs(143) <= not (a xor b);
    layer7_outputs(144) <= not (a or b);
    layer7_outputs(145) <= not b or a;
    layer7_outputs(146) <= b;
    layer7_outputs(147) <= a or b;
    layer7_outputs(148) <= a xor b;
    layer7_outputs(149) <= a;
    layer7_outputs(150) <= '0';
    layer7_outputs(151) <= not (a and b);
    layer7_outputs(152) <= a or b;
    layer7_outputs(153) <= b;
    layer7_outputs(154) <= a and b;
    layer7_outputs(155) <= not a or b;
    layer7_outputs(156) <= a;
    layer7_outputs(157) <= b and not a;
    layer7_outputs(158) <= not a;
    layer7_outputs(159) <= not b;
    layer7_outputs(160) <= a;
    layer7_outputs(161) <= a;
    layer7_outputs(162) <= not b;
    layer7_outputs(163) <= a xor b;
    layer7_outputs(164) <= a or b;
    layer7_outputs(165) <= not (a xor b);
    layer7_outputs(166) <= a and not b;
    layer7_outputs(167) <= a xor b;
    layer7_outputs(168) <= b;
    layer7_outputs(169) <= b;
    layer7_outputs(170) <= not b;
    layer7_outputs(171) <= b;
    layer7_outputs(172) <= not a or b;
    layer7_outputs(173) <= a and not b;
    layer7_outputs(174) <= not (a and b);
    layer7_outputs(175) <= a;
    layer7_outputs(176) <= not b;
    layer7_outputs(177) <= b;
    layer7_outputs(178) <= not a;
    layer7_outputs(179) <= not a;
    layer7_outputs(180) <= not b;
    layer7_outputs(181) <= b and not a;
    layer7_outputs(182) <= b and not a;
    layer7_outputs(183) <= not a or b;
    layer7_outputs(184) <= not (a and b);
    layer7_outputs(185) <= not (a xor b);
    layer7_outputs(186) <= not (a xor b);
    layer7_outputs(187) <= not a;
    layer7_outputs(188) <= a or b;
    layer7_outputs(189) <= a and b;
    layer7_outputs(190) <= not (a xor b);
    layer7_outputs(191) <= b;
    layer7_outputs(192) <= b;
    layer7_outputs(193) <= a or b;
    layer7_outputs(194) <= not b or a;
    layer7_outputs(195) <= not (a xor b);
    layer7_outputs(196) <= not a or b;
    layer7_outputs(197) <= a or b;
    layer7_outputs(198) <= not a;
    layer7_outputs(199) <= a and b;
    layer7_outputs(200) <= b;
    layer7_outputs(201) <= a;
    layer7_outputs(202) <= b;
    layer7_outputs(203) <= not b;
    layer7_outputs(204) <= not a;
    layer7_outputs(205) <= not b;
    layer7_outputs(206) <= not (a and b);
    layer7_outputs(207) <= not a or b;
    layer7_outputs(208) <= not (a and b);
    layer7_outputs(209) <= a and not b;
    layer7_outputs(210) <= not (a and b);
    layer7_outputs(211) <= not a;
    layer7_outputs(212) <= not b;
    layer7_outputs(213) <= b and not a;
    layer7_outputs(214) <= not (a xor b);
    layer7_outputs(215) <= not b;
    layer7_outputs(216) <= not (a xor b);
    layer7_outputs(217) <= not b;
    layer7_outputs(218) <= '1';
    layer7_outputs(219) <= b and not a;
    layer7_outputs(220) <= not (a xor b);
    layer7_outputs(221) <= a and b;
    layer7_outputs(222) <= a or b;
    layer7_outputs(223) <= a and not b;
    layer7_outputs(224) <= not b;
    layer7_outputs(225) <= b;
    layer7_outputs(226) <= not (a and b);
    layer7_outputs(227) <= not (a or b);
    layer7_outputs(228) <= b;
    layer7_outputs(229) <= a;
    layer7_outputs(230) <= not a;
    layer7_outputs(231) <= '0';
    layer7_outputs(232) <= b and not a;
    layer7_outputs(233) <= not a or b;
    layer7_outputs(234) <= b and not a;
    layer7_outputs(235) <= not (a and b);
    layer7_outputs(236) <= a;
    layer7_outputs(237) <= not b;
    layer7_outputs(238) <= a or b;
    layer7_outputs(239) <= not (a xor b);
    layer7_outputs(240) <= not (a and b);
    layer7_outputs(241) <= not a or b;
    layer7_outputs(242) <= not (a and b);
    layer7_outputs(243) <= a xor b;
    layer7_outputs(244) <= b;
    layer7_outputs(245) <= not b or a;
    layer7_outputs(246) <= not a or b;
    layer7_outputs(247) <= not b;
    layer7_outputs(248) <= b;
    layer7_outputs(249) <= b and not a;
    layer7_outputs(250) <= a and not b;
    layer7_outputs(251) <= a and b;
    layer7_outputs(252) <= not (a and b);
    layer7_outputs(253) <= not a or b;
    layer7_outputs(254) <= b and not a;
    layer7_outputs(255) <= not (a xor b);
    layer7_outputs(256) <= b;
    layer7_outputs(257) <= not a;
    layer7_outputs(258) <= not a or b;
    layer7_outputs(259) <= a;
    layer7_outputs(260) <= not b;
    layer7_outputs(261) <= b;
    layer7_outputs(262) <= not a or b;
    layer7_outputs(263) <= a xor b;
    layer7_outputs(264) <= not a or b;
    layer7_outputs(265) <= b;
    layer7_outputs(266) <= not a;
    layer7_outputs(267) <= not b;
    layer7_outputs(268) <= not (a xor b);
    layer7_outputs(269) <= not (a xor b);
    layer7_outputs(270) <= '0';
    layer7_outputs(271) <= not a;
    layer7_outputs(272) <= a and not b;
    layer7_outputs(273) <= a;
    layer7_outputs(274) <= not (a or b);
    layer7_outputs(275) <= not b or a;
    layer7_outputs(276) <= a;
    layer7_outputs(277) <= not b;
    layer7_outputs(278) <= b and not a;
    layer7_outputs(279) <= b and not a;
    layer7_outputs(280) <= a and b;
    layer7_outputs(281) <= a and not b;
    layer7_outputs(282) <= a or b;
    layer7_outputs(283) <= not (a xor b);
    layer7_outputs(284) <= not (a or b);
    layer7_outputs(285) <= a and b;
    layer7_outputs(286) <= not a or b;
    layer7_outputs(287) <= b and not a;
    layer7_outputs(288) <= a;
    layer7_outputs(289) <= not b or a;
    layer7_outputs(290) <= not a;
    layer7_outputs(291) <= '0';
    layer7_outputs(292) <= not a;
    layer7_outputs(293) <= not a;
    layer7_outputs(294) <= a;
    layer7_outputs(295) <= not (a xor b);
    layer7_outputs(296) <= not a;
    layer7_outputs(297) <= not (a xor b);
    layer7_outputs(298) <= not a or b;
    layer7_outputs(299) <= a xor b;
    layer7_outputs(300) <= not (a and b);
    layer7_outputs(301) <= not (a or b);
    layer7_outputs(302) <= not b;
    layer7_outputs(303) <= not b;
    layer7_outputs(304) <= b;
    layer7_outputs(305) <= b;
    layer7_outputs(306) <= a;
    layer7_outputs(307) <= not a;
    layer7_outputs(308) <= not (a xor b);
    layer7_outputs(309) <= not b;
    layer7_outputs(310) <= a;
    layer7_outputs(311) <= a and b;
    layer7_outputs(312) <= a;
    layer7_outputs(313) <= not a or b;
    layer7_outputs(314) <= not b;
    layer7_outputs(315) <= a and not b;
    layer7_outputs(316) <= not a or b;
    layer7_outputs(317) <= not b or a;
    layer7_outputs(318) <= not b;
    layer7_outputs(319) <= not a;
    layer7_outputs(320) <= not a;
    layer7_outputs(321) <= a xor b;
    layer7_outputs(322) <= '1';
    layer7_outputs(323) <= not a or b;
    layer7_outputs(324) <= a;
    layer7_outputs(325) <= not a;
    layer7_outputs(326) <= b;
    layer7_outputs(327) <= a;
    layer7_outputs(328) <= a or b;
    layer7_outputs(329) <= not b;
    layer7_outputs(330) <= not a;
    layer7_outputs(331) <= not a or b;
    layer7_outputs(332) <= a and b;
    layer7_outputs(333) <= a and not b;
    layer7_outputs(334) <= a xor b;
    layer7_outputs(335) <= not b or a;
    layer7_outputs(336) <= a xor b;
    layer7_outputs(337) <= not a or b;
    layer7_outputs(338) <= not a;
    layer7_outputs(339) <= b and not a;
    layer7_outputs(340) <= not b;
    layer7_outputs(341) <= not b or a;
    layer7_outputs(342) <= b;
    layer7_outputs(343) <= a xor b;
    layer7_outputs(344) <= not a;
    layer7_outputs(345) <= not (a or b);
    layer7_outputs(346) <= not b;
    layer7_outputs(347) <= a xor b;
    layer7_outputs(348) <= a xor b;
    layer7_outputs(349) <= not (a and b);
    layer7_outputs(350) <= a and not b;
    layer7_outputs(351) <= a and not b;
    layer7_outputs(352) <= not a;
    layer7_outputs(353) <= '0';
    layer7_outputs(354) <= not a;
    layer7_outputs(355) <= b;
    layer7_outputs(356) <= a;
    layer7_outputs(357) <= a xor b;
    layer7_outputs(358) <= b;
    layer7_outputs(359) <= not (a xor b);
    layer7_outputs(360) <= not (a xor b);
    layer7_outputs(361) <= a and b;
    layer7_outputs(362) <= not a;
    layer7_outputs(363) <= b;
    layer7_outputs(364) <= a;
    layer7_outputs(365) <= not b or a;
    layer7_outputs(366) <= b and not a;
    layer7_outputs(367) <= b;
    layer7_outputs(368) <= not b;
    layer7_outputs(369) <= not (a and b);
    layer7_outputs(370) <= not (a and b);
    layer7_outputs(371) <= a;
    layer7_outputs(372) <= not (a or b);
    layer7_outputs(373) <= not (a and b);
    layer7_outputs(374) <= not a or b;
    layer7_outputs(375) <= b;
    layer7_outputs(376) <= not (a or b);
    layer7_outputs(377) <= not (a and b);
    layer7_outputs(378) <= a or b;
    layer7_outputs(379) <= not (a xor b);
    layer7_outputs(380) <= a and not b;
    layer7_outputs(381) <= a and b;
    layer7_outputs(382) <= not (a and b);
    layer7_outputs(383) <= a xor b;
    layer7_outputs(384) <= not a;
    layer7_outputs(385) <= not a;
    layer7_outputs(386) <= '1';
    layer7_outputs(387) <= not a;
    layer7_outputs(388) <= not b;
    layer7_outputs(389) <= a;
    layer7_outputs(390) <= b and not a;
    layer7_outputs(391) <= b;
    layer7_outputs(392) <= a;
    layer7_outputs(393) <= b and not a;
    layer7_outputs(394) <= not b;
    layer7_outputs(395) <= a or b;
    layer7_outputs(396) <= not a;
    layer7_outputs(397) <= a;
    layer7_outputs(398) <= b and not a;
    layer7_outputs(399) <= not a;
    layer7_outputs(400) <= a xor b;
    layer7_outputs(401) <= a;
    layer7_outputs(402) <= not a or b;
    layer7_outputs(403) <= a and b;
    layer7_outputs(404) <= not a;
    layer7_outputs(405) <= a xor b;
    layer7_outputs(406) <= b and not a;
    layer7_outputs(407) <= a;
    layer7_outputs(408) <= not (a xor b);
    layer7_outputs(409) <= not b or a;
    layer7_outputs(410) <= a or b;
    layer7_outputs(411) <= not b;
    layer7_outputs(412) <= not (a or b);
    layer7_outputs(413) <= not a;
    layer7_outputs(414) <= not a;
    layer7_outputs(415) <= not (a xor b);
    layer7_outputs(416) <= b;
    layer7_outputs(417) <= a and b;
    layer7_outputs(418) <= b and not a;
    layer7_outputs(419) <= not b;
    layer7_outputs(420) <= b;
    layer7_outputs(421) <= b;
    layer7_outputs(422) <= a and not b;
    layer7_outputs(423) <= a xor b;
    layer7_outputs(424) <= not a;
    layer7_outputs(425) <= not b;
    layer7_outputs(426) <= b;
    layer7_outputs(427) <= a xor b;
    layer7_outputs(428) <= a xor b;
    layer7_outputs(429) <= not b;
    layer7_outputs(430) <= not b or a;
    layer7_outputs(431) <= not b or a;
    layer7_outputs(432) <= '1';
    layer7_outputs(433) <= a;
    layer7_outputs(434) <= b;
    layer7_outputs(435) <= not a;
    layer7_outputs(436) <= not b;
    layer7_outputs(437) <= a;
    layer7_outputs(438) <= b;
    layer7_outputs(439) <= a;
    layer7_outputs(440) <= a and not b;
    layer7_outputs(441) <= b;
    layer7_outputs(442) <= b;
    layer7_outputs(443) <= a xor b;
    layer7_outputs(444) <= not a;
    layer7_outputs(445) <= not (a xor b);
    layer7_outputs(446) <= a;
    layer7_outputs(447) <= not a;
    layer7_outputs(448) <= not b;
    layer7_outputs(449) <= a;
    layer7_outputs(450) <= not a;
    layer7_outputs(451) <= '1';
    layer7_outputs(452) <= not a;
    layer7_outputs(453) <= not b;
    layer7_outputs(454) <= not b;
    layer7_outputs(455) <= b;
    layer7_outputs(456) <= not (a xor b);
    layer7_outputs(457) <= a and b;
    layer7_outputs(458) <= b and not a;
    layer7_outputs(459) <= b and not a;
    layer7_outputs(460) <= '1';
    layer7_outputs(461) <= a;
    layer7_outputs(462) <= not b;
    layer7_outputs(463) <= not (a xor b);
    layer7_outputs(464) <= b;
    layer7_outputs(465) <= not b;
    layer7_outputs(466) <= not (a xor b);
    layer7_outputs(467) <= a;
    layer7_outputs(468) <= not a;
    layer7_outputs(469) <= b;
    layer7_outputs(470) <= a;
    layer7_outputs(471) <= b;
    layer7_outputs(472) <= not (a xor b);
    layer7_outputs(473) <= a;
    layer7_outputs(474) <= b;
    layer7_outputs(475) <= b and not a;
    layer7_outputs(476) <= a xor b;
    layer7_outputs(477) <= a and not b;
    layer7_outputs(478) <= a;
    layer7_outputs(479) <= a and b;
    layer7_outputs(480) <= b;
    layer7_outputs(481) <= not a;
    layer7_outputs(482) <= a;
    layer7_outputs(483) <= '0';
    layer7_outputs(484) <= not (a xor b);
    layer7_outputs(485) <= not a;
    layer7_outputs(486) <= b and not a;
    layer7_outputs(487) <= not (a or b);
    layer7_outputs(488) <= not (a and b);
    layer7_outputs(489) <= not a;
    layer7_outputs(490) <= a and b;
    layer7_outputs(491) <= a and not b;
    layer7_outputs(492) <= not b;
    layer7_outputs(493) <= b;
    layer7_outputs(494) <= a;
    layer7_outputs(495) <= not b;
    layer7_outputs(496) <= b;
    layer7_outputs(497) <= not b or a;
    layer7_outputs(498) <= not (a and b);
    layer7_outputs(499) <= b;
    layer7_outputs(500) <= b;
    layer7_outputs(501) <= b;
    layer7_outputs(502) <= a and not b;
    layer7_outputs(503) <= a;
    layer7_outputs(504) <= b and not a;
    layer7_outputs(505) <= a or b;
    layer7_outputs(506) <= not b;
    layer7_outputs(507) <= not a;
    layer7_outputs(508) <= not a;
    layer7_outputs(509) <= a and b;
    layer7_outputs(510) <= not b;
    layer7_outputs(511) <= not a;
    layer7_outputs(512) <= not b;
    layer7_outputs(513) <= a xor b;
    layer7_outputs(514) <= a;
    layer7_outputs(515) <= a;
    layer7_outputs(516) <= not a or b;
    layer7_outputs(517) <= a and not b;
    layer7_outputs(518) <= a xor b;
    layer7_outputs(519) <= not b or a;
    layer7_outputs(520) <= not (a or b);
    layer7_outputs(521) <= b;
    layer7_outputs(522) <= not a;
    layer7_outputs(523) <= not a;
    layer7_outputs(524) <= not a;
    layer7_outputs(525) <= a;
    layer7_outputs(526) <= a;
    layer7_outputs(527) <= a xor b;
    layer7_outputs(528) <= b;
    layer7_outputs(529) <= not (a and b);
    layer7_outputs(530) <= not a or b;
    layer7_outputs(531) <= a;
    layer7_outputs(532) <= not b;
    layer7_outputs(533) <= '0';
    layer7_outputs(534) <= not (a and b);
    layer7_outputs(535) <= b;
    layer7_outputs(536) <= not b;
    layer7_outputs(537) <= a;
    layer7_outputs(538) <= not a;
    layer7_outputs(539) <= not (a and b);
    layer7_outputs(540) <= a;
    layer7_outputs(541) <= a xor b;
    layer7_outputs(542) <= b and not a;
    layer7_outputs(543) <= b and not a;
    layer7_outputs(544) <= a;
    layer7_outputs(545) <= not b;
    layer7_outputs(546) <= a and b;
    layer7_outputs(547) <= a;
    layer7_outputs(548) <= not b;
    layer7_outputs(549) <= not a or b;
    layer7_outputs(550) <= b and not a;
    layer7_outputs(551) <= b and not a;
    layer7_outputs(552) <= a and not b;
    layer7_outputs(553) <= a xor b;
    layer7_outputs(554) <= a and not b;
    layer7_outputs(555) <= a and b;
    layer7_outputs(556) <= not a;
    layer7_outputs(557) <= not b or a;
    layer7_outputs(558) <= not (a or b);
    layer7_outputs(559) <= not (a or b);
    layer7_outputs(560) <= not (a and b);
    layer7_outputs(561) <= not b;
    layer7_outputs(562) <= not a or b;
    layer7_outputs(563) <= b and not a;
    layer7_outputs(564) <= not (a xor b);
    layer7_outputs(565) <= not (a xor b);
    layer7_outputs(566) <= a and not b;
    layer7_outputs(567) <= not (a xor b);
    layer7_outputs(568) <= not a or b;
    layer7_outputs(569) <= a or b;
    layer7_outputs(570) <= b;
    layer7_outputs(571) <= b;
    layer7_outputs(572) <= a and b;
    layer7_outputs(573) <= b and not a;
    layer7_outputs(574) <= not a;
    layer7_outputs(575) <= not (a and b);
    layer7_outputs(576) <= not (a or b);
    layer7_outputs(577) <= not b;
    layer7_outputs(578) <= b;
    layer7_outputs(579) <= not (a xor b);
    layer7_outputs(580) <= b and not a;
    layer7_outputs(581) <= b and not a;
    layer7_outputs(582) <= b;
    layer7_outputs(583) <= not (a or b);
    layer7_outputs(584) <= not b;
    layer7_outputs(585) <= not (a xor b);
    layer7_outputs(586) <= not (a xor b);
    layer7_outputs(587) <= b;
    layer7_outputs(588) <= not a;
    layer7_outputs(589) <= not a;
    layer7_outputs(590) <= b;
    layer7_outputs(591) <= '0';
    layer7_outputs(592) <= a xor b;
    layer7_outputs(593) <= not (a xor b);
    layer7_outputs(594) <= not b or a;
    layer7_outputs(595) <= not a;
    layer7_outputs(596) <= not (a and b);
    layer7_outputs(597) <= not a;
    layer7_outputs(598) <= not a;
    layer7_outputs(599) <= not (a or b);
    layer7_outputs(600) <= b;
    layer7_outputs(601) <= not (a xor b);
    layer7_outputs(602) <= a and b;
    layer7_outputs(603) <= not a;
    layer7_outputs(604) <= not b;
    layer7_outputs(605) <= not a;
    layer7_outputs(606) <= b;
    layer7_outputs(607) <= a and not b;
    layer7_outputs(608) <= not b or a;
    layer7_outputs(609) <= not b;
    layer7_outputs(610) <= a;
    layer7_outputs(611) <= not a;
    layer7_outputs(612) <= not b;
    layer7_outputs(613) <= not b;
    layer7_outputs(614) <= b;
    layer7_outputs(615) <= a and not b;
    layer7_outputs(616) <= not b;
    layer7_outputs(617) <= not b;
    layer7_outputs(618) <= a xor b;
    layer7_outputs(619) <= a and b;
    layer7_outputs(620) <= a or b;
    layer7_outputs(621) <= not b;
    layer7_outputs(622) <= b and not a;
    layer7_outputs(623) <= a xor b;
    layer7_outputs(624) <= not a or b;
    layer7_outputs(625) <= b and not a;
    layer7_outputs(626) <= not (a or b);
    layer7_outputs(627) <= a;
    layer7_outputs(628) <= a;
    layer7_outputs(629) <= a and b;
    layer7_outputs(630) <= a and not b;
    layer7_outputs(631) <= b and not a;
    layer7_outputs(632) <= b;
    layer7_outputs(633) <= not (a or b);
    layer7_outputs(634) <= not a;
    layer7_outputs(635) <= a and b;
    layer7_outputs(636) <= not (a and b);
    layer7_outputs(637) <= b;
    layer7_outputs(638) <= not (a or b);
    layer7_outputs(639) <= a and b;
    layer7_outputs(640) <= not (a or b);
    layer7_outputs(641) <= not (a or b);
    layer7_outputs(642) <= a;
    layer7_outputs(643) <= not b;
    layer7_outputs(644) <= a;
    layer7_outputs(645) <= b;
    layer7_outputs(646) <= not b or a;
    layer7_outputs(647) <= a;
    layer7_outputs(648) <= a;
    layer7_outputs(649) <= a and b;
    layer7_outputs(650) <= not b or a;
    layer7_outputs(651) <= '1';
    layer7_outputs(652) <= a or b;
    layer7_outputs(653) <= not a;
    layer7_outputs(654) <= not a;
    layer7_outputs(655) <= not a or b;
    layer7_outputs(656) <= not a or b;
    layer7_outputs(657) <= a and not b;
    layer7_outputs(658) <= not b;
    layer7_outputs(659) <= a or b;
    layer7_outputs(660) <= a;
    layer7_outputs(661) <= not a;
    layer7_outputs(662) <= not b;
    layer7_outputs(663) <= not (a xor b);
    layer7_outputs(664) <= not a or b;
    layer7_outputs(665) <= a and not b;
    layer7_outputs(666) <= a and b;
    layer7_outputs(667) <= a;
    layer7_outputs(668) <= not b;
    layer7_outputs(669) <= b;
    layer7_outputs(670) <= not b or a;
    layer7_outputs(671) <= a and not b;
    layer7_outputs(672) <= b;
    layer7_outputs(673) <= a xor b;
    layer7_outputs(674) <= not b;
    layer7_outputs(675) <= not (a xor b);
    layer7_outputs(676) <= a and b;
    layer7_outputs(677) <= not a;
    layer7_outputs(678) <= not a or b;
    layer7_outputs(679) <= b and not a;
    layer7_outputs(680) <= not b;
    layer7_outputs(681) <= not (a xor b);
    layer7_outputs(682) <= a and b;
    layer7_outputs(683) <= not a;
    layer7_outputs(684) <= not a;
    layer7_outputs(685) <= not a;
    layer7_outputs(686) <= not (a xor b);
    layer7_outputs(687) <= not (a xor b);
    layer7_outputs(688) <= a xor b;
    layer7_outputs(689) <= not b or a;
    layer7_outputs(690) <= not (a or b);
    layer7_outputs(691) <= a;
    layer7_outputs(692) <= '0';
    layer7_outputs(693) <= not (a xor b);
    layer7_outputs(694) <= not a;
    layer7_outputs(695) <= not a;
    layer7_outputs(696) <= b;
    layer7_outputs(697) <= a;
    layer7_outputs(698) <= not (a xor b);
    layer7_outputs(699) <= not b or a;
    layer7_outputs(700) <= a;
    layer7_outputs(701) <= not (a xor b);
    layer7_outputs(702) <= a and b;
    layer7_outputs(703) <= a xor b;
    layer7_outputs(704) <= not b;
    layer7_outputs(705) <= not b;
    layer7_outputs(706) <= b;
    layer7_outputs(707) <= a and b;
    layer7_outputs(708) <= a;
    layer7_outputs(709) <= not a;
    layer7_outputs(710) <= not a or b;
    layer7_outputs(711) <= not (a and b);
    layer7_outputs(712) <= a or b;
    layer7_outputs(713) <= b;
    layer7_outputs(714) <= not b or a;
    layer7_outputs(715) <= not (a or b);
    layer7_outputs(716) <= not b;
    layer7_outputs(717) <= a or b;
    layer7_outputs(718) <= not b;
    layer7_outputs(719) <= not a;
    layer7_outputs(720) <= b;
    layer7_outputs(721) <= not b;
    layer7_outputs(722) <= not (a or b);
    layer7_outputs(723) <= b;
    layer7_outputs(724) <= not b;
    layer7_outputs(725) <= not a;
    layer7_outputs(726) <= not b;
    layer7_outputs(727) <= a and not b;
    layer7_outputs(728) <= not (a or b);
    layer7_outputs(729) <= a or b;
    layer7_outputs(730) <= b and not a;
    layer7_outputs(731) <= not a or b;
    layer7_outputs(732) <= '0';
    layer7_outputs(733) <= not (a or b);
    layer7_outputs(734) <= '1';
    layer7_outputs(735) <= not (a and b);
    layer7_outputs(736) <= not (a or b);
    layer7_outputs(737) <= a and not b;
    layer7_outputs(738) <= a or b;
    layer7_outputs(739) <= not (a or b);
    layer7_outputs(740) <= not b or a;
    layer7_outputs(741) <= '0';
    layer7_outputs(742) <= not (a or b);
    layer7_outputs(743) <= a;
    layer7_outputs(744) <= not (a or b);
    layer7_outputs(745) <= not (a xor b);
    layer7_outputs(746) <= not b;
    layer7_outputs(747) <= not a;
    layer7_outputs(748) <= not (a or b);
    layer7_outputs(749) <= not a or b;
    layer7_outputs(750) <= not (a or b);
    layer7_outputs(751) <= a;
    layer7_outputs(752) <= a xor b;
    layer7_outputs(753) <= not a or b;
    layer7_outputs(754) <= not a;
    layer7_outputs(755) <= not (a and b);
    layer7_outputs(756) <= not a or b;
    layer7_outputs(757) <= not (a or b);
    layer7_outputs(758) <= not (a xor b);
    layer7_outputs(759) <= a;
    layer7_outputs(760) <= a and b;
    layer7_outputs(761) <= b;
    layer7_outputs(762) <= a;
    layer7_outputs(763) <= not a;
    layer7_outputs(764) <= a and b;
    layer7_outputs(765) <= b;
    layer7_outputs(766) <= a and not b;
    layer7_outputs(767) <= not b;
    layer7_outputs(768) <= b;
    layer7_outputs(769) <= a xor b;
    layer7_outputs(770) <= not a;
    layer7_outputs(771) <= not (a or b);
    layer7_outputs(772) <= not a;
    layer7_outputs(773) <= a and not b;
    layer7_outputs(774) <= a and not b;
    layer7_outputs(775) <= a;
    layer7_outputs(776) <= not (a or b);
    layer7_outputs(777) <= not (a xor b);
    layer7_outputs(778) <= not b;
    layer7_outputs(779) <= b and not a;
    layer7_outputs(780) <= not b or a;
    layer7_outputs(781) <= not b or a;
    layer7_outputs(782) <= '0';
    layer7_outputs(783) <= not b or a;
    layer7_outputs(784) <= b and not a;
    layer7_outputs(785) <= a and not b;
    layer7_outputs(786) <= not a;
    layer7_outputs(787) <= b;
    layer7_outputs(788) <= a;
    layer7_outputs(789) <= not (a or b);
    layer7_outputs(790) <= a and b;
    layer7_outputs(791) <= not (a or b);
    layer7_outputs(792) <= a;
    layer7_outputs(793) <= a or b;
    layer7_outputs(794) <= not (a and b);
    layer7_outputs(795) <= b;
    layer7_outputs(796) <= a xor b;
    layer7_outputs(797) <= a;
    layer7_outputs(798) <= b;
    layer7_outputs(799) <= not a;
    layer7_outputs(800) <= not (a or b);
    layer7_outputs(801) <= a;
    layer7_outputs(802) <= not b;
    layer7_outputs(803) <= not a;
    layer7_outputs(804) <= b;
    layer7_outputs(805) <= a xor b;
    layer7_outputs(806) <= a or b;
    layer7_outputs(807) <= not b;
    layer7_outputs(808) <= b;
    layer7_outputs(809) <= b;
    layer7_outputs(810) <= not (a xor b);
    layer7_outputs(811) <= a and not b;
    layer7_outputs(812) <= not (a xor b);
    layer7_outputs(813) <= a;
    layer7_outputs(814) <= not (a and b);
    layer7_outputs(815) <= not (a or b);
    layer7_outputs(816) <= a and not b;
    layer7_outputs(817) <= a and b;
    layer7_outputs(818) <= a and not b;
    layer7_outputs(819) <= not a;
    layer7_outputs(820) <= a;
    layer7_outputs(821) <= not (a xor b);
    layer7_outputs(822) <= not a or b;
    layer7_outputs(823) <= a and not b;
    layer7_outputs(824) <= not b;
    layer7_outputs(825) <= not b;
    layer7_outputs(826) <= a xor b;
    layer7_outputs(827) <= b and not a;
    layer7_outputs(828) <= a or b;
    layer7_outputs(829) <= a and not b;
    layer7_outputs(830) <= b;
    layer7_outputs(831) <= a and b;
    layer7_outputs(832) <= not a or b;
    layer7_outputs(833) <= a;
    layer7_outputs(834) <= a and b;
    layer7_outputs(835) <= a and not b;
    layer7_outputs(836) <= b;
    layer7_outputs(837) <= a and not b;
    layer7_outputs(838) <= '0';
    layer7_outputs(839) <= not b;
    layer7_outputs(840) <= a or b;
    layer7_outputs(841) <= not (a xor b);
    layer7_outputs(842) <= a xor b;
    layer7_outputs(843) <= not b;
    layer7_outputs(844) <= not (a and b);
    layer7_outputs(845) <= not b;
    layer7_outputs(846) <= not (a or b);
    layer7_outputs(847) <= b and not a;
    layer7_outputs(848) <= b and not a;
    layer7_outputs(849) <= '1';
    layer7_outputs(850) <= not b;
    layer7_outputs(851) <= a or b;
    layer7_outputs(852) <= not b;
    layer7_outputs(853) <= not b or a;
    layer7_outputs(854) <= a and b;
    layer7_outputs(855) <= not b;
    layer7_outputs(856) <= not (a and b);
    layer7_outputs(857) <= not (a xor b);
    layer7_outputs(858) <= not b;
    layer7_outputs(859) <= not (a or b);
    layer7_outputs(860) <= not (a or b);
    layer7_outputs(861) <= not a;
    layer7_outputs(862) <= a and not b;
    layer7_outputs(863) <= a xor b;
    layer7_outputs(864) <= b;
    layer7_outputs(865) <= a or b;
    layer7_outputs(866) <= '0';
    layer7_outputs(867) <= b and not a;
    layer7_outputs(868) <= not (a and b);
    layer7_outputs(869) <= b;
    layer7_outputs(870) <= a;
    layer7_outputs(871) <= a;
    layer7_outputs(872) <= '0';
    layer7_outputs(873) <= b and not a;
    layer7_outputs(874) <= '1';
    layer7_outputs(875) <= not a;
    layer7_outputs(876) <= not a;
    layer7_outputs(877) <= a and not b;
    layer7_outputs(878) <= not (a and b);
    layer7_outputs(879) <= not b;
    layer7_outputs(880) <= a xor b;
    layer7_outputs(881) <= not (a and b);
    layer7_outputs(882) <= a and not b;
    layer7_outputs(883) <= a or b;
    layer7_outputs(884) <= a;
    layer7_outputs(885) <= not a;
    layer7_outputs(886) <= not a;
    layer7_outputs(887) <= a xor b;
    layer7_outputs(888) <= not a;
    layer7_outputs(889) <= not b;
    layer7_outputs(890) <= not a or b;
    layer7_outputs(891) <= not (a or b);
    layer7_outputs(892) <= not a;
    layer7_outputs(893) <= not (a or b);
    layer7_outputs(894) <= a and not b;
    layer7_outputs(895) <= not (a xor b);
    layer7_outputs(896) <= b;
    layer7_outputs(897) <= not a or b;
    layer7_outputs(898) <= '1';
    layer7_outputs(899) <= not (a or b);
    layer7_outputs(900) <= b;
    layer7_outputs(901) <= a;
    layer7_outputs(902) <= not b or a;
    layer7_outputs(903) <= not b;
    layer7_outputs(904) <= not b;
    layer7_outputs(905) <= not (a or b);
    layer7_outputs(906) <= a;
    layer7_outputs(907) <= a and not b;
    layer7_outputs(908) <= not a or b;
    layer7_outputs(909) <= b;
    layer7_outputs(910) <= not (a xor b);
    layer7_outputs(911) <= a or b;
    layer7_outputs(912) <= not a;
    layer7_outputs(913) <= not b;
    layer7_outputs(914) <= not b;
    layer7_outputs(915) <= not (a and b);
    layer7_outputs(916) <= not b;
    layer7_outputs(917) <= not b;
    layer7_outputs(918) <= not (a and b);
    layer7_outputs(919) <= a xor b;
    layer7_outputs(920) <= not a;
    layer7_outputs(921) <= not a;
    layer7_outputs(922) <= b and not a;
    layer7_outputs(923) <= not b or a;
    layer7_outputs(924) <= not (a and b);
    layer7_outputs(925) <= a xor b;
    layer7_outputs(926) <= not b;
    layer7_outputs(927) <= not a or b;
    layer7_outputs(928) <= not (a xor b);
    layer7_outputs(929) <= not (a xor b);
    layer7_outputs(930) <= not (a and b);
    layer7_outputs(931) <= not (a or b);
    layer7_outputs(932) <= not a;
    layer7_outputs(933) <= a;
    layer7_outputs(934) <= not a or b;
    layer7_outputs(935) <= not (a xor b);
    layer7_outputs(936) <= not (a xor b);
    layer7_outputs(937) <= not a;
    layer7_outputs(938) <= a;
    layer7_outputs(939) <= not (a and b);
    layer7_outputs(940) <= not b;
    layer7_outputs(941) <= not (a or b);
    layer7_outputs(942) <= not (a and b);
    layer7_outputs(943) <= not b;
    layer7_outputs(944) <= a or b;
    layer7_outputs(945) <= a xor b;
    layer7_outputs(946) <= b and not a;
    layer7_outputs(947) <= a and not b;
    layer7_outputs(948) <= not (a xor b);
    layer7_outputs(949) <= not a;
    layer7_outputs(950) <= a and not b;
    layer7_outputs(951) <= not (a xor b);
    layer7_outputs(952) <= not b;
    layer7_outputs(953) <= not a or b;
    layer7_outputs(954) <= a xor b;
    layer7_outputs(955) <= not a or b;
    layer7_outputs(956) <= not a;
    layer7_outputs(957) <= a;
    layer7_outputs(958) <= not a;
    layer7_outputs(959) <= not (a and b);
    layer7_outputs(960) <= a;
    layer7_outputs(961) <= not b;
    layer7_outputs(962) <= '0';
    layer7_outputs(963) <= not (a or b);
    layer7_outputs(964) <= not b or a;
    layer7_outputs(965) <= a or b;
    layer7_outputs(966) <= a or b;
    layer7_outputs(967) <= not a;
    layer7_outputs(968) <= a;
    layer7_outputs(969) <= b and not a;
    layer7_outputs(970) <= '1';
    layer7_outputs(971) <= not a;
    layer7_outputs(972) <= not (a or b);
    layer7_outputs(973) <= a and not b;
    layer7_outputs(974) <= not (a xor b);
    layer7_outputs(975) <= b;
    layer7_outputs(976) <= not (a or b);
    layer7_outputs(977) <= not (a or b);
    layer7_outputs(978) <= not (a xor b);
    layer7_outputs(979) <= a xor b;
    layer7_outputs(980) <= a xor b;
    layer7_outputs(981) <= not b;
    layer7_outputs(982) <= '1';
    layer7_outputs(983) <= not (a and b);
    layer7_outputs(984) <= a;
    layer7_outputs(985) <= a;
    layer7_outputs(986) <= a and not b;
    layer7_outputs(987) <= a or b;
    layer7_outputs(988) <= b and not a;
    layer7_outputs(989) <= b;
    layer7_outputs(990) <= not (a and b);
    layer7_outputs(991) <= a and b;
    layer7_outputs(992) <= b;
    layer7_outputs(993) <= not (a or b);
    layer7_outputs(994) <= a;
    layer7_outputs(995) <= not a;
    layer7_outputs(996) <= not b;
    layer7_outputs(997) <= not a;
    layer7_outputs(998) <= not (a xor b);
    layer7_outputs(999) <= not a or b;
    layer7_outputs(1000) <= a or b;
    layer7_outputs(1001) <= a;
    layer7_outputs(1002) <= b;
    layer7_outputs(1003) <= a xor b;
    layer7_outputs(1004) <= b;
    layer7_outputs(1005) <= b and not a;
    layer7_outputs(1006) <= b and not a;
    layer7_outputs(1007) <= b;
    layer7_outputs(1008) <= not (a or b);
    layer7_outputs(1009) <= a;
    layer7_outputs(1010) <= not b;
    layer7_outputs(1011) <= a;
    layer7_outputs(1012) <= b;
    layer7_outputs(1013) <= not (a and b);
    layer7_outputs(1014) <= not (a or b);
    layer7_outputs(1015) <= not (a xor b);
    layer7_outputs(1016) <= b;
    layer7_outputs(1017) <= not a or b;
    layer7_outputs(1018) <= not b;
    layer7_outputs(1019) <= not b or a;
    layer7_outputs(1020) <= '1';
    layer7_outputs(1021) <= '0';
    layer7_outputs(1022) <= not a;
    layer7_outputs(1023) <= not (a or b);
    layer7_outputs(1024) <= a;
    layer7_outputs(1025) <= a;
    layer7_outputs(1026) <= not b or a;
    layer7_outputs(1027) <= not (a and b);
    layer7_outputs(1028) <= not a or b;
    layer7_outputs(1029) <= not (a or b);
    layer7_outputs(1030) <= a;
    layer7_outputs(1031) <= a;
    layer7_outputs(1032) <= a;
    layer7_outputs(1033) <= b;
    layer7_outputs(1034) <= b;
    layer7_outputs(1035) <= a and b;
    layer7_outputs(1036) <= b;
    layer7_outputs(1037) <= not b;
    layer7_outputs(1038) <= not (a or b);
    layer7_outputs(1039) <= not b;
    layer7_outputs(1040) <= b;
    layer7_outputs(1041) <= a or b;
    layer7_outputs(1042) <= not b or a;
    layer7_outputs(1043) <= not b or a;
    layer7_outputs(1044) <= a and b;
    layer7_outputs(1045) <= a and not b;
    layer7_outputs(1046) <= not (a or b);
    layer7_outputs(1047) <= a or b;
    layer7_outputs(1048) <= a or b;
    layer7_outputs(1049) <= b;
    layer7_outputs(1050) <= b;
    layer7_outputs(1051) <= not a or b;
    layer7_outputs(1052) <= not a;
    layer7_outputs(1053) <= a xor b;
    layer7_outputs(1054) <= b;
    layer7_outputs(1055) <= not (a or b);
    layer7_outputs(1056) <= not b or a;
    layer7_outputs(1057) <= not (a xor b);
    layer7_outputs(1058) <= a;
    layer7_outputs(1059) <= b;
    layer7_outputs(1060) <= a and b;
    layer7_outputs(1061) <= not a;
    layer7_outputs(1062) <= a and not b;
    layer7_outputs(1063) <= b and not a;
    layer7_outputs(1064) <= not b or a;
    layer7_outputs(1065) <= b and not a;
    layer7_outputs(1066) <= b;
    layer7_outputs(1067) <= not a or b;
    layer7_outputs(1068) <= not a;
    layer7_outputs(1069) <= not (a and b);
    layer7_outputs(1070) <= not b;
    layer7_outputs(1071) <= not b;
    layer7_outputs(1072) <= not (a and b);
    layer7_outputs(1073) <= not b;
    layer7_outputs(1074) <= b;
    layer7_outputs(1075) <= not a;
    layer7_outputs(1076) <= not b;
    layer7_outputs(1077) <= b;
    layer7_outputs(1078) <= a or b;
    layer7_outputs(1079) <= b;
    layer7_outputs(1080) <= a xor b;
    layer7_outputs(1081) <= not (a xor b);
    layer7_outputs(1082) <= not a or b;
    layer7_outputs(1083) <= not a;
    layer7_outputs(1084) <= a;
    layer7_outputs(1085) <= not (a xor b);
    layer7_outputs(1086) <= not b;
    layer7_outputs(1087) <= not b;
    layer7_outputs(1088) <= not b or a;
    layer7_outputs(1089) <= not (a xor b);
    layer7_outputs(1090) <= not (a and b);
    layer7_outputs(1091) <= a xor b;
    layer7_outputs(1092) <= b and not a;
    layer7_outputs(1093) <= not a;
    layer7_outputs(1094) <= b;
    layer7_outputs(1095) <= a and b;
    layer7_outputs(1096) <= not (a or b);
    layer7_outputs(1097) <= b and not a;
    layer7_outputs(1098) <= not b;
    layer7_outputs(1099) <= a xor b;
    layer7_outputs(1100) <= not a;
    layer7_outputs(1101) <= not b or a;
    layer7_outputs(1102) <= a and not b;
    layer7_outputs(1103) <= b and not a;
    layer7_outputs(1104) <= a;
    layer7_outputs(1105) <= not b or a;
    layer7_outputs(1106) <= b;
    layer7_outputs(1107) <= not b;
    layer7_outputs(1108) <= a;
    layer7_outputs(1109) <= b;
    layer7_outputs(1110) <= a;
    layer7_outputs(1111) <= a;
    layer7_outputs(1112) <= not a;
    layer7_outputs(1113) <= '0';
    layer7_outputs(1114) <= a or b;
    layer7_outputs(1115) <= not (a or b);
    layer7_outputs(1116) <= a and not b;
    layer7_outputs(1117) <= b and not a;
    layer7_outputs(1118) <= not b;
    layer7_outputs(1119) <= a or b;
    layer7_outputs(1120) <= a xor b;
    layer7_outputs(1121) <= a;
    layer7_outputs(1122) <= b;
    layer7_outputs(1123) <= not (a or b);
    layer7_outputs(1124) <= a xor b;
    layer7_outputs(1125) <= a and not b;
    layer7_outputs(1126) <= b;
    layer7_outputs(1127) <= b;
    layer7_outputs(1128) <= not (a and b);
    layer7_outputs(1129) <= not (a xor b);
    layer7_outputs(1130) <= a xor b;
    layer7_outputs(1131) <= not b;
    layer7_outputs(1132) <= a or b;
    layer7_outputs(1133) <= a;
    layer7_outputs(1134) <= '0';
    layer7_outputs(1135) <= not (a and b);
    layer7_outputs(1136) <= not a;
    layer7_outputs(1137) <= not a;
    layer7_outputs(1138) <= not a;
    layer7_outputs(1139) <= a;
    layer7_outputs(1140) <= not a;
    layer7_outputs(1141) <= not a or b;
    layer7_outputs(1142) <= b and not a;
    layer7_outputs(1143) <= not b or a;
    layer7_outputs(1144) <= not b;
    layer7_outputs(1145) <= not (a xor b);
    layer7_outputs(1146) <= b and not a;
    layer7_outputs(1147) <= a;
    layer7_outputs(1148) <= not b or a;
    layer7_outputs(1149) <= not a or b;
    layer7_outputs(1150) <= not b;
    layer7_outputs(1151) <= b;
    layer7_outputs(1152) <= a;
    layer7_outputs(1153) <= not (a and b);
    layer7_outputs(1154) <= not (a xor b);
    layer7_outputs(1155) <= b and not a;
    layer7_outputs(1156) <= a;
    layer7_outputs(1157) <= not a or b;
    layer7_outputs(1158) <= not b;
    layer7_outputs(1159) <= a;
    layer7_outputs(1160) <= not a or b;
    layer7_outputs(1161) <= not b;
    layer7_outputs(1162) <= a;
    layer7_outputs(1163) <= not b;
    layer7_outputs(1164) <= a;
    layer7_outputs(1165) <= not (a xor b);
    layer7_outputs(1166) <= a and b;
    layer7_outputs(1167) <= b;
    layer7_outputs(1168) <= not (a and b);
    layer7_outputs(1169) <= not b or a;
    layer7_outputs(1170) <= not b;
    layer7_outputs(1171) <= not b;
    layer7_outputs(1172) <= a xor b;
    layer7_outputs(1173) <= a xor b;
    layer7_outputs(1174) <= not a;
    layer7_outputs(1175) <= not b;
    layer7_outputs(1176) <= b;
    layer7_outputs(1177) <= not a;
    layer7_outputs(1178) <= b and not a;
    layer7_outputs(1179) <= a xor b;
    layer7_outputs(1180) <= b;
    layer7_outputs(1181) <= not a;
    layer7_outputs(1182) <= b;
    layer7_outputs(1183) <= not (a xor b);
    layer7_outputs(1184) <= a xor b;
    layer7_outputs(1185) <= not b;
    layer7_outputs(1186) <= b;
    layer7_outputs(1187) <= a;
    layer7_outputs(1188) <= b and not a;
    layer7_outputs(1189) <= not b;
    layer7_outputs(1190) <= not (a and b);
    layer7_outputs(1191) <= not (a or b);
    layer7_outputs(1192) <= a xor b;
    layer7_outputs(1193) <= a and not b;
    layer7_outputs(1194) <= not a;
    layer7_outputs(1195) <= not a;
    layer7_outputs(1196) <= a;
    layer7_outputs(1197) <= not b;
    layer7_outputs(1198) <= not (a xor b);
    layer7_outputs(1199) <= a and not b;
    layer7_outputs(1200) <= a xor b;
    layer7_outputs(1201) <= not (a xor b);
    layer7_outputs(1202) <= not (a xor b);
    layer7_outputs(1203) <= not (a xor b);
    layer7_outputs(1204) <= not b;
    layer7_outputs(1205) <= a xor b;
    layer7_outputs(1206) <= a;
    layer7_outputs(1207) <= a;
    layer7_outputs(1208) <= a xor b;
    layer7_outputs(1209) <= a and b;
    layer7_outputs(1210) <= a;
    layer7_outputs(1211) <= b;
    layer7_outputs(1212) <= a;
    layer7_outputs(1213) <= b and not a;
    layer7_outputs(1214) <= b;
    layer7_outputs(1215) <= not (a and b);
    layer7_outputs(1216) <= not (a xor b);
    layer7_outputs(1217) <= b and not a;
    layer7_outputs(1218) <= a;
    layer7_outputs(1219) <= b and not a;
    layer7_outputs(1220) <= not b;
    layer7_outputs(1221) <= not a;
    layer7_outputs(1222) <= b and not a;
    layer7_outputs(1223) <= b;
    layer7_outputs(1224) <= not a or b;
    layer7_outputs(1225) <= not b or a;
    layer7_outputs(1226) <= a xor b;
    layer7_outputs(1227) <= not b;
    layer7_outputs(1228) <= not b;
    layer7_outputs(1229) <= not a or b;
    layer7_outputs(1230) <= not (a or b);
    layer7_outputs(1231) <= not a;
    layer7_outputs(1232) <= a xor b;
    layer7_outputs(1233) <= not (a xor b);
    layer7_outputs(1234) <= '0';
    layer7_outputs(1235) <= b;
    layer7_outputs(1236) <= a;
    layer7_outputs(1237) <= b;
    layer7_outputs(1238) <= a xor b;
    layer7_outputs(1239) <= a xor b;
    layer7_outputs(1240) <= not b;
    layer7_outputs(1241) <= not a;
    layer7_outputs(1242) <= not a or b;
    layer7_outputs(1243) <= a;
    layer7_outputs(1244) <= b;
    layer7_outputs(1245) <= '0';
    layer7_outputs(1246) <= a or b;
    layer7_outputs(1247) <= not (a xor b);
    layer7_outputs(1248) <= a and not b;
    layer7_outputs(1249) <= a;
    layer7_outputs(1250) <= a or b;
    layer7_outputs(1251) <= not a or b;
    layer7_outputs(1252) <= not a;
    layer7_outputs(1253) <= not a;
    layer7_outputs(1254) <= not a;
    layer7_outputs(1255) <= a and not b;
    layer7_outputs(1256) <= not b;
    layer7_outputs(1257) <= b;
    layer7_outputs(1258) <= not (a and b);
    layer7_outputs(1259) <= not b;
    layer7_outputs(1260) <= a xor b;
    layer7_outputs(1261) <= a;
    layer7_outputs(1262) <= not b;
    layer7_outputs(1263) <= b;
    layer7_outputs(1264) <= '1';
    layer7_outputs(1265) <= not (a and b);
    layer7_outputs(1266) <= a or b;
    layer7_outputs(1267) <= a;
    layer7_outputs(1268) <= a and b;
    layer7_outputs(1269) <= not a;
    layer7_outputs(1270) <= a and b;
    layer7_outputs(1271) <= a;
    layer7_outputs(1272) <= not a;
    layer7_outputs(1273) <= a;
    layer7_outputs(1274) <= not b;
    layer7_outputs(1275) <= not b;
    layer7_outputs(1276) <= a and b;
    layer7_outputs(1277) <= not (a and b);
    layer7_outputs(1278) <= not (a xor b);
    layer7_outputs(1279) <= not b or a;
    layer7_outputs(1280) <= b;
    layer7_outputs(1281) <= not (a xor b);
    layer7_outputs(1282) <= not b;
    layer7_outputs(1283) <= b and not a;
    layer7_outputs(1284) <= a xor b;
    layer7_outputs(1285) <= a or b;
    layer7_outputs(1286) <= a and b;
    layer7_outputs(1287) <= not a;
    layer7_outputs(1288) <= a xor b;
    layer7_outputs(1289) <= a;
    layer7_outputs(1290) <= b;
    layer7_outputs(1291) <= '1';
    layer7_outputs(1292) <= a and not b;
    layer7_outputs(1293) <= not b;
    layer7_outputs(1294) <= not a;
    layer7_outputs(1295) <= a;
    layer7_outputs(1296) <= b and not a;
    layer7_outputs(1297) <= not b;
    layer7_outputs(1298) <= not a;
    layer7_outputs(1299) <= not b;
    layer7_outputs(1300) <= b and not a;
    layer7_outputs(1301) <= not (a xor b);
    layer7_outputs(1302) <= not a or b;
    layer7_outputs(1303) <= a xor b;
    layer7_outputs(1304) <= a;
    layer7_outputs(1305) <= not b;
    layer7_outputs(1306) <= a and not b;
    layer7_outputs(1307) <= not a or b;
    layer7_outputs(1308) <= not (a xor b);
    layer7_outputs(1309) <= b;
    layer7_outputs(1310) <= not b;
    layer7_outputs(1311) <= b;
    layer7_outputs(1312) <= not (a and b);
    layer7_outputs(1313) <= a;
    layer7_outputs(1314) <= not a;
    layer7_outputs(1315) <= a and b;
    layer7_outputs(1316) <= not (a xor b);
    layer7_outputs(1317) <= b and not a;
    layer7_outputs(1318) <= b and not a;
    layer7_outputs(1319) <= not a;
    layer7_outputs(1320) <= '1';
    layer7_outputs(1321) <= b;
    layer7_outputs(1322) <= not b;
    layer7_outputs(1323) <= b and not a;
    layer7_outputs(1324) <= a and not b;
    layer7_outputs(1325) <= a xor b;
    layer7_outputs(1326) <= not b;
    layer7_outputs(1327) <= not (a or b);
    layer7_outputs(1328) <= b;
    layer7_outputs(1329) <= a and not b;
    layer7_outputs(1330) <= a xor b;
    layer7_outputs(1331) <= not (a or b);
    layer7_outputs(1332) <= not b or a;
    layer7_outputs(1333) <= not b or a;
    layer7_outputs(1334) <= a and b;
    layer7_outputs(1335) <= not b;
    layer7_outputs(1336) <= not a;
    layer7_outputs(1337) <= not (a or b);
    layer7_outputs(1338) <= a;
    layer7_outputs(1339) <= not a;
    layer7_outputs(1340) <= a and b;
    layer7_outputs(1341) <= '0';
    layer7_outputs(1342) <= not b;
    layer7_outputs(1343) <= not a;
    layer7_outputs(1344) <= '0';
    layer7_outputs(1345) <= not b;
    layer7_outputs(1346) <= b and not a;
    layer7_outputs(1347) <= a and not b;
    layer7_outputs(1348) <= a and not b;
    layer7_outputs(1349) <= b;
    layer7_outputs(1350) <= not (a xor b);
    layer7_outputs(1351) <= not b or a;
    layer7_outputs(1352) <= not a or b;
    layer7_outputs(1353) <= not (a and b);
    layer7_outputs(1354) <= a;
    layer7_outputs(1355) <= not (a or b);
    layer7_outputs(1356) <= a or b;
    layer7_outputs(1357) <= not (a xor b);
    layer7_outputs(1358) <= a xor b;
    layer7_outputs(1359) <= not (a and b);
    layer7_outputs(1360) <= not (a or b);
    layer7_outputs(1361) <= b;
    layer7_outputs(1362) <= not (a and b);
    layer7_outputs(1363) <= b;
    layer7_outputs(1364) <= a or b;
    layer7_outputs(1365) <= a and not b;
    layer7_outputs(1366) <= a xor b;
    layer7_outputs(1367) <= not a;
    layer7_outputs(1368) <= a;
    layer7_outputs(1369) <= not a;
    layer7_outputs(1370) <= a xor b;
    layer7_outputs(1371) <= a xor b;
    layer7_outputs(1372) <= a;
    layer7_outputs(1373) <= not (a or b);
    layer7_outputs(1374) <= b and not a;
    layer7_outputs(1375) <= a;
    layer7_outputs(1376) <= b;
    layer7_outputs(1377) <= not b or a;
    layer7_outputs(1378) <= b and not a;
    layer7_outputs(1379) <= not (a and b);
    layer7_outputs(1380) <= not (a and b);
    layer7_outputs(1381) <= a and b;
    layer7_outputs(1382) <= b;
    layer7_outputs(1383) <= not b;
    layer7_outputs(1384) <= a and not b;
    layer7_outputs(1385) <= not a;
    layer7_outputs(1386) <= not a;
    layer7_outputs(1387) <= not a;
    layer7_outputs(1388) <= not a or b;
    layer7_outputs(1389) <= a;
    layer7_outputs(1390) <= not (a xor b);
    layer7_outputs(1391) <= a and not b;
    layer7_outputs(1392) <= a or b;
    layer7_outputs(1393) <= not b;
    layer7_outputs(1394) <= a and not b;
    layer7_outputs(1395) <= b;
    layer7_outputs(1396) <= a or b;
    layer7_outputs(1397) <= a;
    layer7_outputs(1398) <= a and b;
    layer7_outputs(1399) <= not b;
    layer7_outputs(1400) <= not b;
    layer7_outputs(1401) <= not b;
    layer7_outputs(1402) <= not (a and b);
    layer7_outputs(1403) <= not a;
    layer7_outputs(1404) <= b;
    layer7_outputs(1405) <= a and b;
    layer7_outputs(1406) <= a xor b;
    layer7_outputs(1407) <= not a;
    layer7_outputs(1408) <= not a or b;
    layer7_outputs(1409) <= a and not b;
    layer7_outputs(1410) <= a;
    layer7_outputs(1411) <= b;
    layer7_outputs(1412) <= a and b;
    layer7_outputs(1413) <= not a;
    layer7_outputs(1414) <= a and not b;
    layer7_outputs(1415) <= not b;
    layer7_outputs(1416) <= not a;
    layer7_outputs(1417) <= not a or b;
    layer7_outputs(1418) <= not a;
    layer7_outputs(1419) <= not (a and b);
    layer7_outputs(1420) <= a;
    layer7_outputs(1421) <= b;
    layer7_outputs(1422) <= b;
    layer7_outputs(1423) <= a;
    layer7_outputs(1424) <= a xor b;
    layer7_outputs(1425) <= b;
    layer7_outputs(1426) <= a;
    layer7_outputs(1427) <= a;
    layer7_outputs(1428) <= a;
    layer7_outputs(1429) <= b and not a;
    layer7_outputs(1430) <= a or b;
    layer7_outputs(1431) <= a or b;
    layer7_outputs(1432) <= not a;
    layer7_outputs(1433) <= b and not a;
    layer7_outputs(1434) <= b and not a;
    layer7_outputs(1435) <= b;
    layer7_outputs(1436) <= not b;
    layer7_outputs(1437) <= a;
    layer7_outputs(1438) <= b and not a;
    layer7_outputs(1439) <= a;
    layer7_outputs(1440) <= not (a xor b);
    layer7_outputs(1441) <= not (a xor b);
    layer7_outputs(1442) <= not (a or b);
    layer7_outputs(1443) <= a xor b;
    layer7_outputs(1444) <= not (a and b);
    layer7_outputs(1445) <= not a;
    layer7_outputs(1446) <= not (a or b);
    layer7_outputs(1447) <= a and b;
    layer7_outputs(1448) <= a or b;
    layer7_outputs(1449) <= a;
    layer7_outputs(1450) <= not b;
    layer7_outputs(1451) <= a;
    layer7_outputs(1452) <= not a;
    layer7_outputs(1453) <= not a or b;
    layer7_outputs(1454) <= b and not a;
    layer7_outputs(1455) <= a;
    layer7_outputs(1456) <= not b;
    layer7_outputs(1457) <= not b;
    layer7_outputs(1458) <= '0';
    layer7_outputs(1459) <= a and b;
    layer7_outputs(1460) <= a and b;
    layer7_outputs(1461) <= '0';
    layer7_outputs(1462) <= a xor b;
    layer7_outputs(1463) <= b;
    layer7_outputs(1464) <= a xor b;
    layer7_outputs(1465) <= not b;
    layer7_outputs(1466) <= not a or b;
    layer7_outputs(1467) <= a and b;
    layer7_outputs(1468) <= a xor b;
    layer7_outputs(1469) <= not a or b;
    layer7_outputs(1470) <= not b;
    layer7_outputs(1471) <= not b or a;
    layer7_outputs(1472) <= b;
    layer7_outputs(1473) <= not (a xor b);
    layer7_outputs(1474) <= not a;
    layer7_outputs(1475) <= a or b;
    layer7_outputs(1476) <= a;
    layer7_outputs(1477) <= a xor b;
    layer7_outputs(1478) <= not (a or b);
    layer7_outputs(1479) <= not a;
    layer7_outputs(1480) <= not b;
    layer7_outputs(1481) <= b and not a;
    layer7_outputs(1482) <= a and b;
    layer7_outputs(1483) <= not a;
    layer7_outputs(1484) <= '0';
    layer7_outputs(1485) <= not (a xor b);
    layer7_outputs(1486) <= not (a or b);
    layer7_outputs(1487) <= not a;
    layer7_outputs(1488) <= not (a or b);
    layer7_outputs(1489) <= not a or b;
    layer7_outputs(1490) <= a;
    layer7_outputs(1491) <= a xor b;
    layer7_outputs(1492) <= '0';
    layer7_outputs(1493) <= a or b;
    layer7_outputs(1494) <= '1';
    layer7_outputs(1495) <= a xor b;
    layer7_outputs(1496) <= not a;
    layer7_outputs(1497) <= not a or b;
    layer7_outputs(1498) <= a;
    layer7_outputs(1499) <= b;
    layer7_outputs(1500) <= not (a and b);
    layer7_outputs(1501) <= a or b;
    layer7_outputs(1502) <= a;
    layer7_outputs(1503) <= a;
    layer7_outputs(1504) <= '1';
    layer7_outputs(1505) <= not b or a;
    layer7_outputs(1506) <= a;
    layer7_outputs(1507) <= a or b;
    layer7_outputs(1508) <= a or b;
    layer7_outputs(1509) <= not a or b;
    layer7_outputs(1510) <= a or b;
    layer7_outputs(1511) <= a or b;
    layer7_outputs(1512) <= a;
    layer7_outputs(1513) <= a xor b;
    layer7_outputs(1514) <= a or b;
    layer7_outputs(1515) <= a;
    layer7_outputs(1516) <= not b;
    layer7_outputs(1517) <= b;
    layer7_outputs(1518) <= b;
    layer7_outputs(1519) <= a;
    layer7_outputs(1520) <= b;
    layer7_outputs(1521) <= not (a and b);
    layer7_outputs(1522) <= a and b;
    layer7_outputs(1523) <= '0';
    layer7_outputs(1524) <= a xor b;
    layer7_outputs(1525) <= b;
    layer7_outputs(1526) <= a and b;
    layer7_outputs(1527) <= not a or b;
    layer7_outputs(1528) <= not a or b;
    layer7_outputs(1529) <= not b;
    layer7_outputs(1530) <= b;
    layer7_outputs(1531) <= not (a xor b);
    layer7_outputs(1532) <= a xor b;
    layer7_outputs(1533) <= not (a xor b);
    layer7_outputs(1534) <= not a or b;
    layer7_outputs(1535) <= not (a or b);
    layer7_outputs(1536) <= a xor b;
    layer7_outputs(1537) <= not a;
    layer7_outputs(1538) <= not b;
    layer7_outputs(1539) <= not (a xor b);
    layer7_outputs(1540) <= a and not b;
    layer7_outputs(1541) <= not (a xor b);
    layer7_outputs(1542) <= a;
    layer7_outputs(1543) <= a;
    layer7_outputs(1544) <= b;
    layer7_outputs(1545) <= a xor b;
    layer7_outputs(1546) <= b;
    layer7_outputs(1547) <= a;
    layer7_outputs(1548) <= not a or b;
    layer7_outputs(1549) <= not a;
    layer7_outputs(1550) <= not b;
    layer7_outputs(1551) <= not (a and b);
    layer7_outputs(1552) <= not b;
    layer7_outputs(1553) <= not b;
    layer7_outputs(1554) <= not (a xor b);
    layer7_outputs(1555) <= not b;
    layer7_outputs(1556) <= a or b;
    layer7_outputs(1557) <= a and b;
    layer7_outputs(1558) <= not (a and b);
    layer7_outputs(1559) <= a;
    layer7_outputs(1560) <= not (a and b);
    layer7_outputs(1561) <= a or b;
    layer7_outputs(1562) <= a xor b;
    layer7_outputs(1563) <= a xor b;
    layer7_outputs(1564) <= a xor b;
    layer7_outputs(1565) <= not b;
    layer7_outputs(1566) <= not (a xor b);
    layer7_outputs(1567) <= a and not b;
    layer7_outputs(1568) <= not (a and b);
    layer7_outputs(1569) <= not a;
    layer7_outputs(1570) <= a xor b;
    layer7_outputs(1571) <= not (a xor b);
    layer7_outputs(1572) <= a xor b;
    layer7_outputs(1573) <= not (a or b);
    layer7_outputs(1574) <= a and b;
    layer7_outputs(1575) <= b;
    layer7_outputs(1576) <= a;
    layer7_outputs(1577) <= b;
    layer7_outputs(1578) <= b and not a;
    layer7_outputs(1579) <= a or b;
    layer7_outputs(1580) <= b and not a;
    layer7_outputs(1581) <= not b;
    layer7_outputs(1582) <= not b;
    layer7_outputs(1583) <= a and not b;
    layer7_outputs(1584) <= not a;
    layer7_outputs(1585) <= b;
    layer7_outputs(1586) <= not (a or b);
    layer7_outputs(1587) <= a xor b;
    layer7_outputs(1588) <= b;
    layer7_outputs(1589) <= not a;
    layer7_outputs(1590) <= not (a or b);
    layer7_outputs(1591) <= not a or b;
    layer7_outputs(1592) <= not a;
    layer7_outputs(1593) <= not b;
    layer7_outputs(1594) <= b;
    layer7_outputs(1595) <= a and b;
    layer7_outputs(1596) <= not b or a;
    layer7_outputs(1597) <= '0';
    layer7_outputs(1598) <= a and b;
    layer7_outputs(1599) <= not b or a;
    layer7_outputs(1600) <= not a;
    layer7_outputs(1601) <= b;
    layer7_outputs(1602) <= b;
    layer7_outputs(1603) <= not b;
    layer7_outputs(1604) <= a;
    layer7_outputs(1605) <= '0';
    layer7_outputs(1606) <= not (a xor b);
    layer7_outputs(1607) <= b and not a;
    layer7_outputs(1608) <= a;
    layer7_outputs(1609) <= not b;
    layer7_outputs(1610) <= '1';
    layer7_outputs(1611) <= b;
    layer7_outputs(1612) <= b;
    layer7_outputs(1613) <= a or b;
    layer7_outputs(1614) <= not b or a;
    layer7_outputs(1615) <= not a;
    layer7_outputs(1616) <= a and b;
    layer7_outputs(1617) <= a;
    layer7_outputs(1618) <= a;
    layer7_outputs(1619) <= a;
    layer7_outputs(1620) <= not b;
    layer7_outputs(1621) <= a or b;
    layer7_outputs(1622) <= not b or a;
    layer7_outputs(1623) <= b;
    layer7_outputs(1624) <= a xor b;
    layer7_outputs(1625) <= b;
    layer7_outputs(1626) <= not a or b;
    layer7_outputs(1627) <= not a;
    layer7_outputs(1628) <= a and not b;
    layer7_outputs(1629) <= not b or a;
    layer7_outputs(1630) <= a xor b;
    layer7_outputs(1631) <= a;
    layer7_outputs(1632) <= a;
    layer7_outputs(1633) <= a or b;
    layer7_outputs(1634) <= not b;
    layer7_outputs(1635) <= b;
    layer7_outputs(1636) <= not a;
    layer7_outputs(1637) <= not (a or b);
    layer7_outputs(1638) <= not (a xor b);
    layer7_outputs(1639) <= not a;
    layer7_outputs(1640) <= not b or a;
    layer7_outputs(1641) <= not a;
    layer7_outputs(1642) <= not b;
    layer7_outputs(1643) <= not b or a;
    layer7_outputs(1644) <= b;
    layer7_outputs(1645) <= not b;
    layer7_outputs(1646) <= a xor b;
    layer7_outputs(1647) <= not a;
    layer7_outputs(1648) <= not a;
    layer7_outputs(1649) <= a;
    layer7_outputs(1650) <= a xor b;
    layer7_outputs(1651) <= not b or a;
    layer7_outputs(1652) <= not (a or b);
    layer7_outputs(1653) <= a;
    layer7_outputs(1654) <= b;
    layer7_outputs(1655) <= a xor b;
    layer7_outputs(1656) <= b and not a;
    layer7_outputs(1657) <= not (a and b);
    layer7_outputs(1658) <= a and b;
    layer7_outputs(1659) <= a and not b;
    layer7_outputs(1660) <= not (a or b);
    layer7_outputs(1661) <= '1';
    layer7_outputs(1662) <= a;
    layer7_outputs(1663) <= not b;
    layer7_outputs(1664) <= a and b;
    layer7_outputs(1665) <= not (a xor b);
    layer7_outputs(1666) <= b;
    layer7_outputs(1667) <= not b or a;
    layer7_outputs(1668) <= not b or a;
    layer7_outputs(1669) <= not (a and b);
    layer7_outputs(1670) <= b;
    layer7_outputs(1671) <= not b;
    layer7_outputs(1672) <= not b or a;
    layer7_outputs(1673) <= a xor b;
    layer7_outputs(1674) <= b;
    layer7_outputs(1675) <= not b;
    layer7_outputs(1676) <= not (a or b);
    layer7_outputs(1677) <= b;
    layer7_outputs(1678) <= a and not b;
    layer7_outputs(1679) <= not a;
    layer7_outputs(1680) <= '0';
    layer7_outputs(1681) <= not a;
    layer7_outputs(1682) <= not a;
    layer7_outputs(1683) <= not (a xor b);
    layer7_outputs(1684) <= not (a and b);
    layer7_outputs(1685) <= not (a xor b);
    layer7_outputs(1686) <= not a or b;
    layer7_outputs(1687) <= not b;
    layer7_outputs(1688) <= not a;
    layer7_outputs(1689) <= not (a xor b);
    layer7_outputs(1690) <= '0';
    layer7_outputs(1691) <= b;
    layer7_outputs(1692) <= not a;
    layer7_outputs(1693) <= a and not b;
    layer7_outputs(1694) <= a or b;
    layer7_outputs(1695) <= not a or b;
    layer7_outputs(1696) <= not b or a;
    layer7_outputs(1697) <= not b or a;
    layer7_outputs(1698) <= b and not a;
    layer7_outputs(1699) <= not a or b;
    layer7_outputs(1700) <= not b;
    layer7_outputs(1701) <= a;
    layer7_outputs(1702) <= a or b;
    layer7_outputs(1703) <= not b;
    layer7_outputs(1704) <= not b or a;
    layer7_outputs(1705) <= b;
    layer7_outputs(1706) <= a;
    layer7_outputs(1707) <= a and not b;
    layer7_outputs(1708) <= not b;
    layer7_outputs(1709) <= not b;
    layer7_outputs(1710) <= a xor b;
    layer7_outputs(1711) <= a and not b;
    layer7_outputs(1712) <= not a;
    layer7_outputs(1713) <= not a or b;
    layer7_outputs(1714) <= a and not b;
    layer7_outputs(1715) <= not a or b;
    layer7_outputs(1716) <= b;
    layer7_outputs(1717) <= not (a or b);
    layer7_outputs(1718) <= a and b;
    layer7_outputs(1719) <= b;
    layer7_outputs(1720) <= not a or b;
    layer7_outputs(1721) <= b and not a;
    layer7_outputs(1722) <= not (a xor b);
    layer7_outputs(1723) <= a;
    layer7_outputs(1724) <= not (a or b);
    layer7_outputs(1725) <= not a or b;
    layer7_outputs(1726) <= not b;
    layer7_outputs(1727) <= a;
    layer7_outputs(1728) <= not a or b;
    layer7_outputs(1729) <= not (a xor b);
    layer7_outputs(1730) <= not a;
    layer7_outputs(1731) <= a or b;
    layer7_outputs(1732) <= a;
    layer7_outputs(1733) <= not b;
    layer7_outputs(1734) <= b and not a;
    layer7_outputs(1735) <= not b;
    layer7_outputs(1736) <= not a;
    layer7_outputs(1737) <= not b;
    layer7_outputs(1738) <= a;
    layer7_outputs(1739) <= not a;
    layer7_outputs(1740) <= a;
    layer7_outputs(1741) <= not a;
    layer7_outputs(1742) <= a;
    layer7_outputs(1743) <= not (a xor b);
    layer7_outputs(1744) <= not (a or b);
    layer7_outputs(1745) <= '0';
    layer7_outputs(1746) <= not (a or b);
    layer7_outputs(1747) <= a and b;
    layer7_outputs(1748) <= not a or b;
    layer7_outputs(1749) <= not (a and b);
    layer7_outputs(1750) <= a xor b;
    layer7_outputs(1751) <= b and not a;
    layer7_outputs(1752) <= a;
    layer7_outputs(1753) <= not a or b;
    layer7_outputs(1754) <= not a;
    layer7_outputs(1755) <= not b;
    layer7_outputs(1756) <= '0';
    layer7_outputs(1757) <= not a;
    layer7_outputs(1758) <= not a;
    layer7_outputs(1759) <= not a;
    layer7_outputs(1760) <= a and not b;
    layer7_outputs(1761) <= not b;
    layer7_outputs(1762) <= not a;
    layer7_outputs(1763) <= not b;
    layer7_outputs(1764) <= not (a and b);
    layer7_outputs(1765) <= a and b;
    layer7_outputs(1766) <= not (a xor b);
    layer7_outputs(1767) <= not a;
    layer7_outputs(1768) <= not b or a;
    layer7_outputs(1769) <= not a or b;
    layer7_outputs(1770) <= a or b;
    layer7_outputs(1771) <= not (a xor b);
    layer7_outputs(1772) <= not b or a;
    layer7_outputs(1773) <= not (a xor b);
    layer7_outputs(1774) <= not b;
    layer7_outputs(1775) <= not b;
    layer7_outputs(1776) <= b;
    layer7_outputs(1777) <= a xor b;
    layer7_outputs(1778) <= b;
    layer7_outputs(1779) <= not (a or b);
    layer7_outputs(1780) <= a or b;
    layer7_outputs(1781) <= b and not a;
    layer7_outputs(1782) <= not a or b;
    layer7_outputs(1783) <= b and not a;
    layer7_outputs(1784) <= a xor b;
    layer7_outputs(1785) <= not b;
    layer7_outputs(1786) <= a xor b;
    layer7_outputs(1787) <= b;
    layer7_outputs(1788) <= a;
    layer7_outputs(1789) <= not (a or b);
    layer7_outputs(1790) <= not b or a;
    layer7_outputs(1791) <= not b;
    layer7_outputs(1792) <= not a;
    layer7_outputs(1793) <= b and not a;
    layer7_outputs(1794) <= a and b;
    layer7_outputs(1795) <= not (a xor b);
    layer7_outputs(1796) <= not a or b;
    layer7_outputs(1797) <= a and b;
    layer7_outputs(1798) <= b and not a;
    layer7_outputs(1799) <= not (a xor b);
    layer7_outputs(1800) <= a;
    layer7_outputs(1801) <= b;
    layer7_outputs(1802) <= not (a or b);
    layer7_outputs(1803) <= b and not a;
    layer7_outputs(1804) <= a xor b;
    layer7_outputs(1805) <= a xor b;
    layer7_outputs(1806) <= not (a xor b);
    layer7_outputs(1807) <= not b;
    layer7_outputs(1808) <= a xor b;
    layer7_outputs(1809) <= not a or b;
    layer7_outputs(1810) <= b;
    layer7_outputs(1811) <= a and not b;
    layer7_outputs(1812) <= a;
    layer7_outputs(1813) <= not b;
    layer7_outputs(1814) <= not b or a;
    layer7_outputs(1815) <= not (a or b);
    layer7_outputs(1816) <= not b;
    layer7_outputs(1817) <= not b;
    layer7_outputs(1818) <= b and not a;
    layer7_outputs(1819) <= not b;
    layer7_outputs(1820) <= not (a or b);
    layer7_outputs(1821) <= b and not a;
    layer7_outputs(1822) <= a xor b;
    layer7_outputs(1823) <= '0';
    layer7_outputs(1824) <= not b or a;
    layer7_outputs(1825) <= a;
    layer7_outputs(1826) <= not b;
    layer7_outputs(1827) <= b;
    layer7_outputs(1828) <= not b;
    layer7_outputs(1829) <= not (a xor b);
    layer7_outputs(1830) <= not a;
    layer7_outputs(1831) <= '0';
    layer7_outputs(1832) <= not a or b;
    layer7_outputs(1833) <= not b;
    layer7_outputs(1834) <= not b or a;
    layer7_outputs(1835) <= not a or b;
    layer7_outputs(1836) <= not (a or b);
    layer7_outputs(1837) <= not b;
    layer7_outputs(1838) <= not b;
    layer7_outputs(1839) <= not b;
    layer7_outputs(1840) <= b;
    layer7_outputs(1841) <= not b or a;
    layer7_outputs(1842) <= not a or b;
    layer7_outputs(1843) <= not (a xor b);
    layer7_outputs(1844) <= b;
    layer7_outputs(1845) <= a and b;
    layer7_outputs(1846) <= not (a xor b);
    layer7_outputs(1847) <= not a;
    layer7_outputs(1848) <= a xor b;
    layer7_outputs(1849) <= a xor b;
    layer7_outputs(1850) <= not (a and b);
    layer7_outputs(1851) <= not a or b;
    layer7_outputs(1852) <= a and b;
    layer7_outputs(1853) <= not b or a;
    layer7_outputs(1854) <= b and not a;
    layer7_outputs(1855) <= b and not a;
    layer7_outputs(1856) <= not b or a;
    layer7_outputs(1857) <= a and not b;
    layer7_outputs(1858) <= b;
    layer7_outputs(1859) <= not b;
    layer7_outputs(1860) <= not b;
    layer7_outputs(1861) <= b and not a;
    layer7_outputs(1862) <= not (a xor b);
    layer7_outputs(1863) <= a and b;
    layer7_outputs(1864) <= not (a or b);
    layer7_outputs(1865) <= not (a and b);
    layer7_outputs(1866) <= b and not a;
    layer7_outputs(1867) <= b;
    layer7_outputs(1868) <= a;
    layer7_outputs(1869) <= a;
    layer7_outputs(1870) <= a and not b;
    layer7_outputs(1871) <= b;
    layer7_outputs(1872) <= a xor b;
    layer7_outputs(1873) <= not (a and b);
    layer7_outputs(1874) <= a;
    layer7_outputs(1875) <= a or b;
    layer7_outputs(1876) <= not b;
    layer7_outputs(1877) <= a;
    layer7_outputs(1878) <= a;
    layer7_outputs(1879) <= a xor b;
    layer7_outputs(1880) <= a;
    layer7_outputs(1881) <= b;
    layer7_outputs(1882) <= not b;
    layer7_outputs(1883) <= not a;
    layer7_outputs(1884) <= '1';
    layer7_outputs(1885) <= b;
    layer7_outputs(1886) <= a and b;
    layer7_outputs(1887) <= not (a and b);
    layer7_outputs(1888) <= a or b;
    layer7_outputs(1889) <= not b or a;
    layer7_outputs(1890) <= b;
    layer7_outputs(1891) <= not (a and b);
    layer7_outputs(1892) <= b;
    layer7_outputs(1893) <= not a;
    layer7_outputs(1894) <= b and not a;
    layer7_outputs(1895) <= b and not a;
    layer7_outputs(1896) <= not a;
    layer7_outputs(1897) <= not a;
    layer7_outputs(1898) <= not b;
    layer7_outputs(1899) <= not (a xor b);
    layer7_outputs(1900) <= a or b;
    layer7_outputs(1901) <= '0';
    layer7_outputs(1902) <= not a or b;
    layer7_outputs(1903) <= a and not b;
    layer7_outputs(1904) <= a and not b;
    layer7_outputs(1905) <= not b;
    layer7_outputs(1906) <= b;
    layer7_outputs(1907) <= a or b;
    layer7_outputs(1908) <= a and not b;
    layer7_outputs(1909) <= not (a xor b);
    layer7_outputs(1910) <= a xor b;
    layer7_outputs(1911) <= not (a or b);
    layer7_outputs(1912) <= not (a and b);
    layer7_outputs(1913) <= a and b;
    layer7_outputs(1914) <= a and not b;
    layer7_outputs(1915) <= not b;
    layer7_outputs(1916) <= a and not b;
    layer7_outputs(1917) <= a;
    layer7_outputs(1918) <= not (a xor b);
    layer7_outputs(1919) <= b;
    layer7_outputs(1920) <= b;
    layer7_outputs(1921) <= not (a and b);
    layer7_outputs(1922) <= not b or a;
    layer7_outputs(1923) <= a;
    layer7_outputs(1924) <= not b or a;
    layer7_outputs(1925) <= not (a and b);
    layer7_outputs(1926) <= not a;
    layer7_outputs(1927) <= not b;
    layer7_outputs(1928) <= not b or a;
    layer7_outputs(1929) <= not (a xor b);
    layer7_outputs(1930) <= not b or a;
    layer7_outputs(1931) <= a or b;
    layer7_outputs(1932) <= '0';
    layer7_outputs(1933) <= not a;
    layer7_outputs(1934) <= a;
    layer7_outputs(1935) <= not a;
    layer7_outputs(1936) <= not (a xor b);
    layer7_outputs(1937) <= not (a xor b);
    layer7_outputs(1938) <= not a;
    layer7_outputs(1939) <= b;
    layer7_outputs(1940) <= not a;
    layer7_outputs(1941) <= not (a xor b);
    layer7_outputs(1942) <= b and not a;
    layer7_outputs(1943) <= a and b;
    layer7_outputs(1944) <= a xor b;
    layer7_outputs(1945) <= not (a or b);
    layer7_outputs(1946) <= a or b;
    layer7_outputs(1947) <= b;
    layer7_outputs(1948) <= not b;
    layer7_outputs(1949) <= not b;
    layer7_outputs(1950) <= not b;
    layer7_outputs(1951) <= not b or a;
    layer7_outputs(1952) <= not (a xor b);
    layer7_outputs(1953) <= not b or a;
    layer7_outputs(1954) <= not (a or b);
    layer7_outputs(1955) <= a xor b;
    layer7_outputs(1956) <= not a;
    layer7_outputs(1957) <= not b;
    layer7_outputs(1958) <= a xor b;
    layer7_outputs(1959) <= not a or b;
    layer7_outputs(1960) <= not b or a;
    layer7_outputs(1961) <= not (a or b);
    layer7_outputs(1962) <= not a;
    layer7_outputs(1963) <= a xor b;
    layer7_outputs(1964) <= not a;
    layer7_outputs(1965) <= not b;
    layer7_outputs(1966) <= not b or a;
    layer7_outputs(1967) <= a or b;
    layer7_outputs(1968) <= b;
    layer7_outputs(1969) <= b and not a;
    layer7_outputs(1970) <= not a;
    layer7_outputs(1971) <= not (a xor b);
    layer7_outputs(1972) <= a and not b;
    layer7_outputs(1973) <= not b;
    layer7_outputs(1974) <= a;
    layer7_outputs(1975) <= b;
    layer7_outputs(1976) <= a and b;
    layer7_outputs(1977) <= not (a or b);
    layer7_outputs(1978) <= a and b;
    layer7_outputs(1979) <= a and not b;
    layer7_outputs(1980) <= not b;
    layer7_outputs(1981) <= not (a xor b);
    layer7_outputs(1982) <= not (a xor b);
    layer7_outputs(1983) <= b and not a;
    layer7_outputs(1984) <= not a;
    layer7_outputs(1985) <= a;
    layer7_outputs(1986) <= not a;
    layer7_outputs(1987) <= a and b;
    layer7_outputs(1988) <= not b;
    layer7_outputs(1989) <= not (a xor b);
    layer7_outputs(1990) <= not b or a;
    layer7_outputs(1991) <= not a or b;
    layer7_outputs(1992) <= a and not b;
    layer7_outputs(1993) <= a xor b;
    layer7_outputs(1994) <= not b or a;
    layer7_outputs(1995) <= a;
    layer7_outputs(1996) <= not (a or b);
    layer7_outputs(1997) <= b;
    layer7_outputs(1998) <= a or b;
    layer7_outputs(1999) <= a or b;
    layer7_outputs(2000) <= a or b;
    layer7_outputs(2001) <= not (a xor b);
    layer7_outputs(2002) <= a xor b;
    layer7_outputs(2003) <= b and not a;
    layer7_outputs(2004) <= not (a xor b);
    layer7_outputs(2005) <= a or b;
    layer7_outputs(2006) <= a and b;
    layer7_outputs(2007) <= not b;
    layer7_outputs(2008) <= not a or b;
    layer7_outputs(2009) <= not (a xor b);
    layer7_outputs(2010) <= a;
    layer7_outputs(2011) <= not b or a;
    layer7_outputs(2012) <= not b;
    layer7_outputs(2013) <= a;
    layer7_outputs(2014) <= a;
    layer7_outputs(2015) <= not b or a;
    layer7_outputs(2016) <= not b;
    layer7_outputs(2017) <= not (a and b);
    layer7_outputs(2018) <= a and b;
    layer7_outputs(2019) <= not (a or b);
    layer7_outputs(2020) <= not b;
    layer7_outputs(2021) <= not (a and b);
    layer7_outputs(2022) <= b;
    layer7_outputs(2023) <= b;
    layer7_outputs(2024) <= not a or b;
    layer7_outputs(2025) <= not a;
    layer7_outputs(2026) <= not a;
    layer7_outputs(2027) <= a xor b;
    layer7_outputs(2028) <= not (a xor b);
    layer7_outputs(2029) <= a;
    layer7_outputs(2030) <= a xor b;
    layer7_outputs(2031) <= a xor b;
    layer7_outputs(2032) <= not b or a;
    layer7_outputs(2033) <= b;
    layer7_outputs(2034) <= '1';
    layer7_outputs(2035) <= b;
    layer7_outputs(2036) <= a or b;
    layer7_outputs(2037) <= a;
    layer7_outputs(2038) <= a xor b;
    layer7_outputs(2039) <= not a or b;
    layer7_outputs(2040) <= a and b;
    layer7_outputs(2041) <= not (a xor b);
    layer7_outputs(2042) <= a;
    layer7_outputs(2043) <= a;
    layer7_outputs(2044) <= not a;
    layer7_outputs(2045) <= not a or b;
    layer7_outputs(2046) <= not b;
    layer7_outputs(2047) <= b;
    layer7_outputs(2048) <= not b;
    layer7_outputs(2049) <= b and not a;
    layer7_outputs(2050) <= a or b;
    layer7_outputs(2051) <= a and not b;
    layer7_outputs(2052) <= not a or b;
    layer7_outputs(2053) <= a xor b;
    layer7_outputs(2054) <= b;
    layer7_outputs(2055) <= not (a or b);
    layer7_outputs(2056) <= not a;
    layer7_outputs(2057) <= a xor b;
    layer7_outputs(2058) <= not a;
    layer7_outputs(2059) <= a;
    layer7_outputs(2060) <= not (a or b);
    layer7_outputs(2061) <= b and not a;
    layer7_outputs(2062) <= not a;
    layer7_outputs(2063) <= not b;
    layer7_outputs(2064) <= a xor b;
    layer7_outputs(2065) <= b and not a;
    layer7_outputs(2066) <= not b;
    layer7_outputs(2067) <= not (a or b);
    layer7_outputs(2068) <= not b;
    layer7_outputs(2069) <= not a;
    layer7_outputs(2070) <= not a;
    layer7_outputs(2071) <= not a or b;
    layer7_outputs(2072) <= not (a and b);
    layer7_outputs(2073) <= not (a and b);
    layer7_outputs(2074) <= a and b;
    layer7_outputs(2075) <= not b;
    layer7_outputs(2076) <= not (a xor b);
    layer7_outputs(2077) <= b;
    layer7_outputs(2078) <= a and not b;
    layer7_outputs(2079) <= b;
    layer7_outputs(2080) <= a xor b;
    layer7_outputs(2081) <= not (a xor b);
    layer7_outputs(2082) <= a xor b;
    layer7_outputs(2083) <= not a;
    layer7_outputs(2084) <= not a;
    layer7_outputs(2085) <= not b;
    layer7_outputs(2086) <= a xor b;
    layer7_outputs(2087) <= not (a or b);
    layer7_outputs(2088) <= a or b;
    layer7_outputs(2089) <= not a or b;
    layer7_outputs(2090) <= not a;
    layer7_outputs(2091) <= not b or a;
    layer7_outputs(2092) <= not a or b;
    layer7_outputs(2093) <= not a or b;
    layer7_outputs(2094) <= a or b;
    layer7_outputs(2095) <= a;
    layer7_outputs(2096) <= '0';
    layer7_outputs(2097) <= b;
    layer7_outputs(2098) <= not b;
    layer7_outputs(2099) <= not b;
    layer7_outputs(2100) <= not b;
    layer7_outputs(2101) <= a or b;
    layer7_outputs(2102) <= b and not a;
    layer7_outputs(2103) <= a and not b;
    layer7_outputs(2104) <= not a;
    layer7_outputs(2105) <= a xor b;
    layer7_outputs(2106) <= a or b;
    layer7_outputs(2107) <= not b;
    layer7_outputs(2108) <= not (a and b);
    layer7_outputs(2109) <= a;
    layer7_outputs(2110) <= not (a and b);
    layer7_outputs(2111) <= a and b;
    layer7_outputs(2112) <= a;
    layer7_outputs(2113) <= not (a xor b);
    layer7_outputs(2114) <= not b or a;
    layer7_outputs(2115) <= not (a xor b);
    layer7_outputs(2116) <= a;
    layer7_outputs(2117) <= a and b;
    layer7_outputs(2118) <= a or b;
    layer7_outputs(2119) <= a and b;
    layer7_outputs(2120) <= a xor b;
    layer7_outputs(2121) <= not a or b;
    layer7_outputs(2122) <= '0';
    layer7_outputs(2123) <= not (a or b);
    layer7_outputs(2124) <= not (a or b);
    layer7_outputs(2125) <= a;
    layer7_outputs(2126) <= b and not a;
    layer7_outputs(2127) <= a and not b;
    layer7_outputs(2128) <= not a;
    layer7_outputs(2129) <= b;
    layer7_outputs(2130) <= a or b;
    layer7_outputs(2131) <= not b or a;
    layer7_outputs(2132) <= b and not a;
    layer7_outputs(2133) <= a;
    layer7_outputs(2134) <= b;
    layer7_outputs(2135) <= not a;
    layer7_outputs(2136) <= not b;
    layer7_outputs(2137) <= not (a and b);
    layer7_outputs(2138) <= b;
    layer7_outputs(2139) <= not (a and b);
    layer7_outputs(2140) <= not (a or b);
    layer7_outputs(2141) <= b;
    layer7_outputs(2142) <= a xor b;
    layer7_outputs(2143) <= not b;
    layer7_outputs(2144) <= b and not a;
    layer7_outputs(2145) <= a;
    layer7_outputs(2146) <= a or b;
    layer7_outputs(2147) <= a and b;
    layer7_outputs(2148) <= not (a xor b);
    layer7_outputs(2149) <= a and not b;
    layer7_outputs(2150) <= b and not a;
    layer7_outputs(2151) <= a and not b;
    layer7_outputs(2152) <= a xor b;
    layer7_outputs(2153) <= b;
    layer7_outputs(2154) <= not a;
    layer7_outputs(2155) <= not b or a;
    layer7_outputs(2156) <= b;
    layer7_outputs(2157) <= b;
    layer7_outputs(2158) <= not a;
    layer7_outputs(2159) <= a;
    layer7_outputs(2160) <= a;
    layer7_outputs(2161) <= a and not b;
    layer7_outputs(2162) <= b and not a;
    layer7_outputs(2163) <= a xor b;
    layer7_outputs(2164) <= a and not b;
    layer7_outputs(2165) <= a;
    layer7_outputs(2166) <= not b or a;
    layer7_outputs(2167) <= not a;
    layer7_outputs(2168) <= not (a and b);
    layer7_outputs(2169) <= '0';
    layer7_outputs(2170) <= b;
    layer7_outputs(2171) <= a;
    layer7_outputs(2172) <= a or b;
    layer7_outputs(2173) <= b and not a;
    layer7_outputs(2174) <= not (a or b);
    layer7_outputs(2175) <= b;
    layer7_outputs(2176) <= a and not b;
    layer7_outputs(2177) <= a and b;
    layer7_outputs(2178) <= a or b;
    layer7_outputs(2179) <= b;
    layer7_outputs(2180) <= not a;
    layer7_outputs(2181) <= a or b;
    layer7_outputs(2182) <= not a;
    layer7_outputs(2183) <= not (a xor b);
    layer7_outputs(2184) <= not a or b;
    layer7_outputs(2185) <= b and not a;
    layer7_outputs(2186) <= not b;
    layer7_outputs(2187) <= not (a and b);
    layer7_outputs(2188) <= not (a and b);
    layer7_outputs(2189) <= a and not b;
    layer7_outputs(2190) <= '1';
    layer7_outputs(2191) <= b;
    layer7_outputs(2192) <= not (a and b);
    layer7_outputs(2193) <= a xor b;
    layer7_outputs(2194) <= not (a xor b);
    layer7_outputs(2195) <= b;
    layer7_outputs(2196) <= a;
    layer7_outputs(2197) <= b;
    layer7_outputs(2198) <= b;
    layer7_outputs(2199) <= b;
    layer7_outputs(2200) <= not (a or b);
    layer7_outputs(2201) <= b and not a;
    layer7_outputs(2202) <= not (a xor b);
    layer7_outputs(2203) <= not b or a;
    layer7_outputs(2204) <= a;
    layer7_outputs(2205) <= not b;
    layer7_outputs(2206) <= not b;
    layer7_outputs(2207) <= not b or a;
    layer7_outputs(2208) <= a xor b;
    layer7_outputs(2209) <= a and b;
    layer7_outputs(2210) <= b;
    layer7_outputs(2211) <= not a or b;
    layer7_outputs(2212) <= not (a and b);
    layer7_outputs(2213) <= b;
    layer7_outputs(2214) <= a;
    layer7_outputs(2215) <= not a or b;
    layer7_outputs(2216) <= not (a or b);
    layer7_outputs(2217) <= a;
    layer7_outputs(2218) <= not b;
    layer7_outputs(2219) <= '1';
    layer7_outputs(2220) <= a;
    layer7_outputs(2221) <= not a;
    layer7_outputs(2222) <= not b;
    layer7_outputs(2223) <= b;
    layer7_outputs(2224) <= not (a xor b);
    layer7_outputs(2225) <= not (a xor b);
    layer7_outputs(2226) <= b;
    layer7_outputs(2227) <= not (a xor b);
    layer7_outputs(2228) <= a xor b;
    layer7_outputs(2229) <= not b;
    layer7_outputs(2230) <= not (a and b);
    layer7_outputs(2231) <= b;
    layer7_outputs(2232) <= not (a xor b);
    layer7_outputs(2233) <= not (a xor b);
    layer7_outputs(2234) <= not (a and b);
    layer7_outputs(2235) <= not (a or b);
    layer7_outputs(2236) <= a and b;
    layer7_outputs(2237) <= a;
    layer7_outputs(2238) <= b;
    layer7_outputs(2239) <= a or b;
    layer7_outputs(2240) <= not (a xor b);
    layer7_outputs(2241) <= not (a and b);
    layer7_outputs(2242) <= not a;
    layer7_outputs(2243) <= not a or b;
    layer7_outputs(2244) <= not a or b;
    layer7_outputs(2245) <= not a;
    layer7_outputs(2246) <= not (a or b);
    layer7_outputs(2247) <= not a;
    layer7_outputs(2248) <= not b or a;
    layer7_outputs(2249) <= a xor b;
    layer7_outputs(2250) <= not b;
    layer7_outputs(2251) <= not a or b;
    layer7_outputs(2252) <= not (a and b);
    layer7_outputs(2253) <= not (a xor b);
    layer7_outputs(2254) <= not b;
    layer7_outputs(2255) <= not (a xor b);
    layer7_outputs(2256) <= a or b;
    layer7_outputs(2257) <= a and not b;
    layer7_outputs(2258) <= not (a xor b);
    layer7_outputs(2259) <= b and not a;
    layer7_outputs(2260) <= b and not a;
    layer7_outputs(2261) <= not a;
    layer7_outputs(2262) <= a xor b;
    layer7_outputs(2263) <= not b or a;
    layer7_outputs(2264) <= not a or b;
    layer7_outputs(2265) <= a and not b;
    layer7_outputs(2266) <= not a;
    layer7_outputs(2267) <= a;
    layer7_outputs(2268) <= not b or a;
    layer7_outputs(2269) <= a;
    layer7_outputs(2270) <= b;
    layer7_outputs(2271) <= not b;
    layer7_outputs(2272) <= a xor b;
    layer7_outputs(2273) <= b;
    layer7_outputs(2274) <= a and not b;
    layer7_outputs(2275) <= a and not b;
    layer7_outputs(2276) <= a and not b;
    layer7_outputs(2277) <= not (a or b);
    layer7_outputs(2278) <= a and not b;
    layer7_outputs(2279) <= a and not b;
    layer7_outputs(2280) <= '0';
    layer7_outputs(2281) <= a xor b;
    layer7_outputs(2282) <= not a or b;
    layer7_outputs(2283) <= '1';
    layer7_outputs(2284) <= not (a xor b);
    layer7_outputs(2285) <= '0';
    layer7_outputs(2286) <= a xor b;
    layer7_outputs(2287) <= b;
    layer7_outputs(2288) <= a xor b;
    layer7_outputs(2289) <= '1';
    layer7_outputs(2290) <= not a or b;
    layer7_outputs(2291) <= a;
    layer7_outputs(2292) <= b;
    layer7_outputs(2293) <= not (a and b);
    layer7_outputs(2294) <= not (a or b);
    layer7_outputs(2295) <= not b or a;
    layer7_outputs(2296) <= b;
    layer7_outputs(2297) <= not b;
    layer7_outputs(2298) <= b and not a;
    layer7_outputs(2299) <= not (a xor b);
    layer7_outputs(2300) <= not b;
    layer7_outputs(2301) <= not a;
    layer7_outputs(2302) <= not a;
    layer7_outputs(2303) <= not (a or b);
    layer7_outputs(2304) <= not a;
    layer7_outputs(2305) <= not (a xor b);
    layer7_outputs(2306) <= not a or b;
    layer7_outputs(2307) <= a and b;
    layer7_outputs(2308) <= a and b;
    layer7_outputs(2309) <= b and not a;
    layer7_outputs(2310) <= not b or a;
    layer7_outputs(2311) <= not b;
    layer7_outputs(2312) <= b and not a;
    layer7_outputs(2313) <= b;
    layer7_outputs(2314) <= not a or b;
    layer7_outputs(2315) <= a xor b;
    layer7_outputs(2316) <= not a;
    layer7_outputs(2317) <= not (a or b);
    layer7_outputs(2318) <= a xor b;
    layer7_outputs(2319) <= not a;
    layer7_outputs(2320) <= not a or b;
    layer7_outputs(2321) <= not a;
    layer7_outputs(2322) <= a or b;
    layer7_outputs(2323) <= not (a or b);
    layer7_outputs(2324) <= not a or b;
    layer7_outputs(2325) <= not (a xor b);
    layer7_outputs(2326) <= '0';
    layer7_outputs(2327) <= b;
    layer7_outputs(2328) <= a and b;
    layer7_outputs(2329) <= '0';
    layer7_outputs(2330) <= not (a and b);
    layer7_outputs(2331) <= not a;
    layer7_outputs(2332) <= not a or b;
    layer7_outputs(2333) <= not b or a;
    layer7_outputs(2334) <= b;
    layer7_outputs(2335) <= b;
    layer7_outputs(2336) <= not b or a;
    layer7_outputs(2337) <= a;
    layer7_outputs(2338) <= not (a and b);
    layer7_outputs(2339) <= a and b;
    layer7_outputs(2340) <= not (a and b);
    layer7_outputs(2341) <= a;
    layer7_outputs(2342) <= not (a xor b);
    layer7_outputs(2343) <= a and b;
    layer7_outputs(2344) <= not (a or b);
    layer7_outputs(2345) <= not a or b;
    layer7_outputs(2346) <= not a;
    layer7_outputs(2347) <= not a;
    layer7_outputs(2348) <= not a or b;
    layer7_outputs(2349) <= not b;
    layer7_outputs(2350) <= a and not b;
    layer7_outputs(2351) <= not b;
    layer7_outputs(2352) <= b and not a;
    layer7_outputs(2353) <= not (a and b);
    layer7_outputs(2354) <= a;
    layer7_outputs(2355) <= not a or b;
    layer7_outputs(2356) <= b;
    layer7_outputs(2357) <= a and not b;
    layer7_outputs(2358) <= not a;
    layer7_outputs(2359) <= a xor b;
    layer7_outputs(2360) <= not b;
    layer7_outputs(2361) <= not (a xor b);
    layer7_outputs(2362) <= a and b;
    layer7_outputs(2363) <= not b;
    layer7_outputs(2364) <= a and not b;
    layer7_outputs(2365) <= not (a or b);
    layer7_outputs(2366) <= b;
    layer7_outputs(2367) <= not a;
    layer7_outputs(2368) <= a;
    layer7_outputs(2369) <= not b;
    layer7_outputs(2370) <= not a;
    layer7_outputs(2371) <= b;
    layer7_outputs(2372) <= b;
    layer7_outputs(2373) <= not b or a;
    layer7_outputs(2374) <= not a;
    layer7_outputs(2375) <= not a;
    layer7_outputs(2376) <= not a;
    layer7_outputs(2377) <= not a or b;
    layer7_outputs(2378) <= a xor b;
    layer7_outputs(2379) <= a or b;
    layer7_outputs(2380) <= a xor b;
    layer7_outputs(2381) <= '0';
    layer7_outputs(2382) <= not b;
    layer7_outputs(2383) <= not a or b;
    layer7_outputs(2384) <= a;
    layer7_outputs(2385) <= not (a and b);
    layer7_outputs(2386) <= not a or b;
    layer7_outputs(2387) <= b;
    layer7_outputs(2388) <= not (a or b);
    layer7_outputs(2389) <= not (a and b);
    layer7_outputs(2390) <= not b;
    layer7_outputs(2391) <= not b;
    layer7_outputs(2392) <= a or b;
    layer7_outputs(2393) <= a or b;
    layer7_outputs(2394) <= a and not b;
    layer7_outputs(2395) <= not a;
    layer7_outputs(2396) <= a and not b;
    layer7_outputs(2397) <= b and not a;
    layer7_outputs(2398) <= b;
    layer7_outputs(2399) <= not b;
    layer7_outputs(2400) <= a;
    layer7_outputs(2401) <= a and b;
    layer7_outputs(2402) <= a and b;
    layer7_outputs(2403) <= not (a or b);
    layer7_outputs(2404) <= b;
    layer7_outputs(2405) <= '0';
    layer7_outputs(2406) <= a and not b;
    layer7_outputs(2407) <= a or b;
    layer7_outputs(2408) <= not (a or b);
    layer7_outputs(2409) <= not b;
    layer7_outputs(2410) <= not a;
    layer7_outputs(2411) <= not (a and b);
    layer7_outputs(2412) <= a;
    layer7_outputs(2413) <= a;
    layer7_outputs(2414) <= not b;
    layer7_outputs(2415) <= b;
    layer7_outputs(2416) <= a xor b;
    layer7_outputs(2417) <= a xor b;
    layer7_outputs(2418) <= a or b;
    layer7_outputs(2419) <= not b or a;
    layer7_outputs(2420) <= a or b;
    layer7_outputs(2421) <= a or b;
    layer7_outputs(2422) <= not a;
    layer7_outputs(2423) <= not b or a;
    layer7_outputs(2424) <= a;
    layer7_outputs(2425) <= not a;
    layer7_outputs(2426) <= b;
    layer7_outputs(2427) <= not (a and b);
    layer7_outputs(2428) <= not a or b;
    layer7_outputs(2429) <= a xor b;
    layer7_outputs(2430) <= a or b;
    layer7_outputs(2431) <= a xor b;
    layer7_outputs(2432) <= not (a and b);
    layer7_outputs(2433) <= a and not b;
    layer7_outputs(2434) <= a xor b;
    layer7_outputs(2435) <= not (a and b);
    layer7_outputs(2436) <= not b or a;
    layer7_outputs(2437) <= a and b;
    layer7_outputs(2438) <= not (a and b);
    layer7_outputs(2439) <= b;
    layer7_outputs(2440) <= b;
    layer7_outputs(2441) <= not (a xor b);
    layer7_outputs(2442) <= not a;
    layer7_outputs(2443) <= not a;
    layer7_outputs(2444) <= a or b;
    layer7_outputs(2445) <= not a;
    layer7_outputs(2446) <= b and not a;
    layer7_outputs(2447) <= a and not b;
    layer7_outputs(2448) <= a or b;
    layer7_outputs(2449) <= a xor b;
    layer7_outputs(2450) <= not a or b;
    layer7_outputs(2451) <= '0';
    layer7_outputs(2452) <= not a;
    layer7_outputs(2453) <= a and b;
    layer7_outputs(2454) <= b;
    layer7_outputs(2455) <= not b;
    layer7_outputs(2456) <= b;
    layer7_outputs(2457) <= b and not a;
    layer7_outputs(2458) <= a xor b;
    layer7_outputs(2459) <= a and b;
    layer7_outputs(2460) <= '1';
    layer7_outputs(2461) <= not (a or b);
    layer7_outputs(2462) <= b and not a;
    layer7_outputs(2463) <= a;
    layer7_outputs(2464) <= b;
    layer7_outputs(2465) <= not a or b;
    layer7_outputs(2466) <= not (a xor b);
    layer7_outputs(2467) <= not a;
    layer7_outputs(2468) <= b;
    layer7_outputs(2469) <= b and not a;
    layer7_outputs(2470) <= not a;
    layer7_outputs(2471) <= not (a xor b);
    layer7_outputs(2472) <= a;
    layer7_outputs(2473) <= not b;
    layer7_outputs(2474) <= b and not a;
    layer7_outputs(2475) <= a;
    layer7_outputs(2476) <= a and not b;
    layer7_outputs(2477) <= not b;
    layer7_outputs(2478) <= not a;
    layer7_outputs(2479) <= not a;
    layer7_outputs(2480) <= a or b;
    layer7_outputs(2481) <= a xor b;
    layer7_outputs(2482) <= b;
    layer7_outputs(2483) <= b;
    layer7_outputs(2484) <= not (a or b);
    layer7_outputs(2485) <= a;
    layer7_outputs(2486) <= a or b;
    layer7_outputs(2487) <= not b or a;
    layer7_outputs(2488) <= '0';
    layer7_outputs(2489) <= not a;
    layer7_outputs(2490) <= b;
    layer7_outputs(2491) <= a;
    layer7_outputs(2492) <= not (a and b);
    layer7_outputs(2493) <= not (a xor b);
    layer7_outputs(2494) <= a;
    layer7_outputs(2495) <= b;
    layer7_outputs(2496) <= not a;
    layer7_outputs(2497) <= not a or b;
    layer7_outputs(2498) <= not (a xor b);
    layer7_outputs(2499) <= not (a and b);
    layer7_outputs(2500) <= not b or a;
    layer7_outputs(2501) <= a and b;
    layer7_outputs(2502) <= a and b;
    layer7_outputs(2503) <= not b or a;
    layer7_outputs(2504) <= b and not a;
    layer7_outputs(2505) <= b;
    layer7_outputs(2506) <= a and b;
    layer7_outputs(2507) <= not a;
    layer7_outputs(2508) <= not a;
    layer7_outputs(2509) <= a and b;
    layer7_outputs(2510) <= a;
    layer7_outputs(2511) <= not b;
    layer7_outputs(2512) <= b;
    layer7_outputs(2513) <= b and not a;
    layer7_outputs(2514) <= a;
    layer7_outputs(2515) <= not a or b;
    layer7_outputs(2516) <= b and not a;
    layer7_outputs(2517) <= b and not a;
    layer7_outputs(2518) <= not b;
    layer7_outputs(2519) <= a;
    layer7_outputs(2520) <= a and not b;
    layer7_outputs(2521) <= b and not a;
    layer7_outputs(2522) <= b;
    layer7_outputs(2523) <= not b or a;
    layer7_outputs(2524) <= a and b;
    layer7_outputs(2525) <= a and not b;
    layer7_outputs(2526) <= a and not b;
    layer7_outputs(2527) <= b;
    layer7_outputs(2528) <= a and not b;
    layer7_outputs(2529) <= not b;
    layer7_outputs(2530) <= not a;
    layer7_outputs(2531) <= not (a or b);
    layer7_outputs(2532) <= not b;
    layer7_outputs(2533) <= a or b;
    layer7_outputs(2534) <= b;
    layer7_outputs(2535) <= '1';
    layer7_outputs(2536) <= not b;
    layer7_outputs(2537) <= a;
    layer7_outputs(2538) <= a and not b;
    layer7_outputs(2539) <= not a;
    layer7_outputs(2540) <= not a;
    layer7_outputs(2541) <= not a or b;
    layer7_outputs(2542) <= not a or b;
    layer7_outputs(2543) <= a and b;
    layer7_outputs(2544) <= a or b;
    layer7_outputs(2545) <= not (a xor b);
    layer7_outputs(2546) <= not b or a;
    layer7_outputs(2547) <= b;
    layer7_outputs(2548) <= not a;
    layer7_outputs(2549) <= not (a or b);
    layer7_outputs(2550) <= not b;
    layer7_outputs(2551) <= a or b;
    layer7_outputs(2552) <= not (a xor b);
    layer7_outputs(2553) <= a;
    layer7_outputs(2554) <= a xor b;
    layer7_outputs(2555) <= a xor b;
    layer7_outputs(2556) <= not b or a;
    layer7_outputs(2557) <= not (a xor b);
    layer7_outputs(2558) <= b and not a;
    layer7_outputs(2559) <= a;
    layer7_outputs(2560) <= a or b;
    layer7_outputs(2561) <= b;
    layer7_outputs(2562) <= b;
    layer7_outputs(2563) <= a xor b;
    layer7_outputs(2564) <= b and not a;
    layer7_outputs(2565) <= a;
    layer7_outputs(2566) <= '1';
    layer7_outputs(2567) <= not a or b;
    layer7_outputs(2568) <= not b or a;
    layer7_outputs(2569) <= a and b;
    layer7_outputs(2570) <= b;
    layer7_outputs(2571) <= b;
    layer7_outputs(2572) <= not a;
    layer7_outputs(2573) <= a xor b;
    layer7_outputs(2574) <= a or b;
    layer7_outputs(2575) <= not (a xor b);
    layer7_outputs(2576) <= not (a xor b);
    layer7_outputs(2577) <= b;
    layer7_outputs(2578) <= b and not a;
    layer7_outputs(2579) <= a and not b;
    layer7_outputs(2580) <= b;
    layer7_outputs(2581) <= a or b;
    layer7_outputs(2582) <= not (a xor b);
    layer7_outputs(2583) <= not a or b;
    layer7_outputs(2584) <= not b or a;
    layer7_outputs(2585) <= not b;
    layer7_outputs(2586) <= a or b;
    layer7_outputs(2587) <= a xor b;
    layer7_outputs(2588) <= a or b;
    layer7_outputs(2589) <= not b or a;
    layer7_outputs(2590) <= b and not a;
    layer7_outputs(2591) <= a and not b;
    layer7_outputs(2592) <= b;
    layer7_outputs(2593) <= not b;
    layer7_outputs(2594) <= not (a xor b);
    layer7_outputs(2595) <= not b;
    layer7_outputs(2596) <= not b or a;
    layer7_outputs(2597) <= a xor b;
    layer7_outputs(2598) <= not b or a;
    layer7_outputs(2599) <= a xor b;
    layer7_outputs(2600) <= not b or a;
    layer7_outputs(2601) <= not b;
    layer7_outputs(2602) <= b;
    layer7_outputs(2603) <= a;
    layer7_outputs(2604) <= a;
    layer7_outputs(2605) <= not b or a;
    layer7_outputs(2606) <= a;
    layer7_outputs(2607) <= not b or a;
    layer7_outputs(2608) <= not (a or b);
    layer7_outputs(2609) <= not b;
    layer7_outputs(2610) <= a xor b;
    layer7_outputs(2611) <= a;
    layer7_outputs(2612) <= not (a xor b);
    layer7_outputs(2613) <= b and not a;
    layer7_outputs(2614) <= '0';
    layer7_outputs(2615) <= not (a and b);
    layer7_outputs(2616) <= b;
    layer7_outputs(2617) <= a and not b;
    layer7_outputs(2618) <= a or b;
    layer7_outputs(2619) <= b;
    layer7_outputs(2620) <= '0';
    layer7_outputs(2621) <= a;
    layer7_outputs(2622) <= a xor b;
    layer7_outputs(2623) <= a or b;
    layer7_outputs(2624) <= not b or a;
    layer7_outputs(2625) <= not (a and b);
    layer7_outputs(2626) <= b and not a;
    layer7_outputs(2627) <= not b;
    layer7_outputs(2628) <= a;
    layer7_outputs(2629) <= a and b;
    layer7_outputs(2630) <= '1';
    layer7_outputs(2631) <= not (a and b);
    layer7_outputs(2632) <= not (a and b);
    layer7_outputs(2633) <= a or b;
    layer7_outputs(2634) <= not b;
    layer7_outputs(2635) <= not (a and b);
    layer7_outputs(2636) <= not b;
    layer7_outputs(2637) <= '1';
    layer7_outputs(2638) <= b and not a;
    layer7_outputs(2639) <= a and b;
    layer7_outputs(2640) <= not b;
    layer7_outputs(2641) <= not (a or b);
    layer7_outputs(2642) <= not a;
    layer7_outputs(2643) <= not b;
    layer7_outputs(2644) <= not a;
    layer7_outputs(2645) <= a and not b;
    layer7_outputs(2646) <= a;
    layer7_outputs(2647) <= a xor b;
    layer7_outputs(2648) <= a and b;
    layer7_outputs(2649) <= a xor b;
    layer7_outputs(2650) <= a or b;
    layer7_outputs(2651) <= b;
    layer7_outputs(2652) <= b and not a;
    layer7_outputs(2653) <= '0';
    layer7_outputs(2654) <= a;
    layer7_outputs(2655) <= not (a xor b);
    layer7_outputs(2656) <= b and not a;
    layer7_outputs(2657) <= not b;
    layer7_outputs(2658) <= not b;
    layer7_outputs(2659) <= not a;
    layer7_outputs(2660) <= not b or a;
    layer7_outputs(2661) <= not (a xor b);
    layer7_outputs(2662) <= not (a or b);
    layer7_outputs(2663) <= a and not b;
    layer7_outputs(2664) <= a xor b;
    layer7_outputs(2665) <= a;
    layer7_outputs(2666) <= not (a or b);
    layer7_outputs(2667) <= b;
    layer7_outputs(2668) <= b;
    layer7_outputs(2669) <= a and b;
    layer7_outputs(2670) <= a and not b;
    layer7_outputs(2671) <= not (a xor b);
    layer7_outputs(2672) <= not b;
    layer7_outputs(2673) <= not a or b;
    layer7_outputs(2674) <= not b or a;
    layer7_outputs(2675) <= a xor b;
    layer7_outputs(2676) <= not (a xor b);
    layer7_outputs(2677) <= not b or a;
    layer7_outputs(2678) <= not b;
    layer7_outputs(2679) <= not b;
    layer7_outputs(2680) <= a and b;
    layer7_outputs(2681) <= a;
    layer7_outputs(2682) <= not b or a;
    layer7_outputs(2683) <= a or b;
    layer7_outputs(2684) <= a;
    layer7_outputs(2685) <= not b;
    layer7_outputs(2686) <= not b;
    layer7_outputs(2687) <= a;
    layer7_outputs(2688) <= not (a xor b);
    layer7_outputs(2689) <= '1';
    layer7_outputs(2690) <= not b;
    layer7_outputs(2691) <= a or b;
    layer7_outputs(2692) <= a;
    layer7_outputs(2693) <= not (a or b);
    layer7_outputs(2694) <= not a or b;
    layer7_outputs(2695) <= not a or b;
    layer7_outputs(2696) <= not a;
    layer7_outputs(2697) <= not a;
    layer7_outputs(2698) <= not a;
    layer7_outputs(2699) <= not a;
    layer7_outputs(2700) <= b and not a;
    layer7_outputs(2701) <= a and not b;
    layer7_outputs(2702) <= not a;
    layer7_outputs(2703) <= b;
    layer7_outputs(2704) <= a;
    layer7_outputs(2705) <= a;
    layer7_outputs(2706) <= not b;
    layer7_outputs(2707) <= a xor b;
    layer7_outputs(2708) <= not b or a;
    layer7_outputs(2709) <= a;
    layer7_outputs(2710) <= not b or a;
    layer7_outputs(2711) <= not a;
    layer7_outputs(2712) <= not a or b;
    layer7_outputs(2713) <= b;
    layer7_outputs(2714) <= a;
    layer7_outputs(2715) <= not a;
    layer7_outputs(2716) <= not a;
    layer7_outputs(2717) <= not (a or b);
    layer7_outputs(2718) <= a;
    layer7_outputs(2719) <= not (a and b);
    layer7_outputs(2720) <= a or b;
    layer7_outputs(2721) <= a or b;
    layer7_outputs(2722) <= not a or b;
    layer7_outputs(2723) <= a or b;
    layer7_outputs(2724) <= b;
    layer7_outputs(2725) <= a xor b;
    layer7_outputs(2726) <= not b;
    layer7_outputs(2727) <= b;
    layer7_outputs(2728) <= a and b;
    layer7_outputs(2729) <= not (a xor b);
    layer7_outputs(2730) <= not (a xor b);
    layer7_outputs(2731) <= a or b;
    layer7_outputs(2732) <= a;
    layer7_outputs(2733) <= not a or b;
    layer7_outputs(2734) <= b;
    layer7_outputs(2735) <= not b;
    layer7_outputs(2736) <= not (a and b);
    layer7_outputs(2737) <= a and b;
    layer7_outputs(2738) <= not (a and b);
    layer7_outputs(2739) <= a and not b;
    layer7_outputs(2740) <= not (a xor b);
    layer7_outputs(2741) <= a xor b;
    layer7_outputs(2742) <= a;
    layer7_outputs(2743) <= b;
    layer7_outputs(2744) <= not a;
    layer7_outputs(2745) <= not a;
    layer7_outputs(2746) <= b and not a;
    layer7_outputs(2747) <= not a;
    layer7_outputs(2748) <= b;
    layer7_outputs(2749) <= not b;
    layer7_outputs(2750) <= not b or a;
    layer7_outputs(2751) <= not b;
    layer7_outputs(2752) <= a;
    layer7_outputs(2753) <= not b;
    layer7_outputs(2754) <= not b;
    layer7_outputs(2755) <= not a;
    layer7_outputs(2756) <= a xor b;
    layer7_outputs(2757) <= not a;
    layer7_outputs(2758) <= b;
    layer7_outputs(2759) <= not b;
    layer7_outputs(2760) <= not (a and b);
    layer7_outputs(2761) <= a xor b;
    layer7_outputs(2762) <= a;
    layer7_outputs(2763) <= not b;
    layer7_outputs(2764) <= not (a and b);
    layer7_outputs(2765) <= a or b;
    layer7_outputs(2766) <= not (a xor b);
    layer7_outputs(2767) <= a and b;
    layer7_outputs(2768) <= not (a or b);
    layer7_outputs(2769) <= a or b;
    layer7_outputs(2770) <= a;
    layer7_outputs(2771) <= not (a xor b);
    layer7_outputs(2772) <= not b;
    layer7_outputs(2773) <= not a;
    layer7_outputs(2774) <= not b;
    layer7_outputs(2775) <= not a or b;
    layer7_outputs(2776) <= not b or a;
    layer7_outputs(2777) <= b;
    layer7_outputs(2778) <= a and b;
    layer7_outputs(2779) <= '1';
    layer7_outputs(2780) <= not b;
    layer7_outputs(2781) <= not b or a;
    layer7_outputs(2782) <= a;
    layer7_outputs(2783) <= a and b;
    layer7_outputs(2784) <= not (a xor b);
    layer7_outputs(2785) <= b and not a;
    layer7_outputs(2786) <= b and not a;
    layer7_outputs(2787) <= a xor b;
    layer7_outputs(2788) <= not b;
    layer7_outputs(2789) <= not a;
    layer7_outputs(2790) <= not (a xor b);
    layer7_outputs(2791) <= not (a and b);
    layer7_outputs(2792) <= not a;
    layer7_outputs(2793) <= a xor b;
    layer7_outputs(2794) <= not (a or b);
    layer7_outputs(2795) <= a and not b;
    layer7_outputs(2796) <= b;
    layer7_outputs(2797) <= a and not b;
    layer7_outputs(2798) <= a or b;
    layer7_outputs(2799) <= not a;
    layer7_outputs(2800) <= not (a or b);
    layer7_outputs(2801) <= not (a and b);
    layer7_outputs(2802) <= not (a xor b);
    layer7_outputs(2803) <= a xor b;
    layer7_outputs(2804) <= a or b;
    layer7_outputs(2805) <= not (a and b);
    layer7_outputs(2806) <= not (a xor b);
    layer7_outputs(2807) <= not (a or b);
    layer7_outputs(2808) <= a and b;
    layer7_outputs(2809) <= a or b;
    layer7_outputs(2810) <= b;
    layer7_outputs(2811) <= b;
    layer7_outputs(2812) <= '1';
    layer7_outputs(2813) <= not b;
    layer7_outputs(2814) <= not (a and b);
    layer7_outputs(2815) <= not (a xor b);
    layer7_outputs(2816) <= not b or a;
    layer7_outputs(2817) <= not b or a;
    layer7_outputs(2818) <= not b;
    layer7_outputs(2819) <= not b;
    layer7_outputs(2820) <= not (a or b);
    layer7_outputs(2821) <= not a;
    layer7_outputs(2822) <= not a;
    layer7_outputs(2823) <= not (a xor b);
    layer7_outputs(2824) <= a;
    layer7_outputs(2825) <= a xor b;
    layer7_outputs(2826) <= not (a xor b);
    layer7_outputs(2827) <= not (a and b);
    layer7_outputs(2828) <= a;
    layer7_outputs(2829) <= a xor b;
    layer7_outputs(2830) <= a;
    layer7_outputs(2831) <= not a;
    layer7_outputs(2832) <= b;
    layer7_outputs(2833) <= not (a xor b);
    layer7_outputs(2834) <= not a;
    layer7_outputs(2835) <= not a or b;
    layer7_outputs(2836) <= a or b;
    layer7_outputs(2837) <= a and b;
    layer7_outputs(2838) <= a and b;
    layer7_outputs(2839) <= '0';
    layer7_outputs(2840) <= a and not b;
    layer7_outputs(2841) <= a or b;
    layer7_outputs(2842) <= a and b;
    layer7_outputs(2843) <= not a;
    layer7_outputs(2844) <= a;
    layer7_outputs(2845) <= a xor b;
    layer7_outputs(2846) <= not (a xor b);
    layer7_outputs(2847) <= b and not a;
    layer7_outputs(2848) <= b and not a;
    layer7_outputs(2849) <= not a;
    layer7_outputs(2850) <= a xor b;
    layer7_outputs(2851) <= b;
    layer7_outputs(2852) <= not a;
    layer7_outputs(2853) <= not (a and b);
    layer7_outputs(2854) <= not a;
    layer7_outputs(2855) <= b and not a;
    layer7_outputs(2856) <= not a or b;
    layer7_outputs(2857) <= not (a xor b);
    layer7_outputs(2858) <= not b or a;
    layer7_outputs(2859) <= a xor b;
    layer7_outputs(2860) <= b;
    layer7_outputs(2861) <= not (a and b);
    layer7_outputs(2862) <= not (a or b);
    layer7_outputs(2863) <= not (a and b);
    layer7_outputs(2864) <= not (a or b);
    layer7_outputs(2865) <= not b or a;
    layer7_outputs(2866) <= not (a and b);
    layer7_outputs(2867) <= not b;
    layer7_outputs(2868) <= a and not b;
    layer7_outputs(2869) <= not a;
    layer7_outputs(2870) <= not b;
    layer7_outputs(2871) <= not b;
    layer7_outputs(2872) <= not b;
    layer7_outputs(2873) <= a and b;
    layer7_outputs(2874) <= not a;
    layer7_outputs(2875) <= b and not a;
    layer7_outputs(2876) <= not (a xor b);
    layer7_outputs(2877) <= a;
    layer7_outputs(2878) <= not (a xor b);
    layer7_outputs(2879) <= a and not b;
    layer7_outputs(2880) <= b;
    layer7_outputs(2881) <= b and not a;
    layer7_outputs(2882) <= a;
    layer7_outputs(2883) <= b;
    layer7_outputs(2884) <= a;
    layer7_outputs(2885) <= a xor b;
    layer7_outputs(2886) <= not b or a;
    layer7_outputs(2887) <= not b;
    layer7_outputs(2888) <= b and not a;
    layer7_outputs(2889) <= '1';
    layer7_outputs(2890) <= not b;
    layer7_outputs(2891) <= a and b;
    layer7_outputs(2892) <= a and not b;
    layer7_outputs(2893) <= a and b;
    layer7_outputs(2894) <= not (a xor b);
    layer7_outputs(2895) <= not a;
    layer7_outputs(2896) <= a and b;
    layer7_outputs(2897) <= not (a or b);
    layer7_outputs(2898) <= '0';
    layer7_outputs(2899) <= a and not b;
    layer7_outputs(2900) <= not a;
    layer7_outputs(2901) <= b;
    layer7_outputs(2902) <= '0';
    layer7_outputs(2903) <= not (a or b);
    layer7_outputs(2904) <= a;
    layer7_outputs(2905) <= a;
    layer7_outputs(2906) <= a xor b;
    layer7_outputs(2907) <= b;
    layer7_outputs(2908) <= a;
    layer7_outputs(2909) <= a xor b;
    layer7_outputs(2910) <= b;
    layer7_outputs(2911) <= not a;
    layer7_outputs(2912) <= not a;
    layer7_outputs(2913) <= not (a xor b);
    layer7_outputs(2914) <= a or b;
    layer7_outputs(2915) <= a and b;
    layer7_outputs(2916) <= not b;
    layer7_outputs(2917) <= a and not b;
    layer7_outputs(2918) <= a;
    layer7_outputs(2919) <= a;
    layer7_outputs(2920) <= not a;
    layer7_outputs(2921) <= a;
    layer7_outputs(2922) <= not a;
    layer7_outputs(2923) <= not b;
    layer7_outputs(2924) <= a and not b;
    layer7_outputs(2925) <= not b or a;
    layer7_outputs(2926) <= not b;
    layer7_outputs(2927) <= a xor b;
    layer7_outputs(2928) <= b and not a;
    layer7_outputs(2929) <= not a;
    layer7_outputs(2930) <= not (a or b);
    layer7_outputs(2931) <= not (a xor b);
    layer7_outputs(2932) <= a;
    layer7_outputs(2933) <= not b;
    layer7_outputs(2934) <= a and not b;
    layer7_outputs(2935) <= b;
    layer7_outputs(2936) <= not b;
    layer7_outputs(2937) <= b;
    layer7_outputs(2938) <= a and not b;
    layer7_outputs(2939) <= b and not a;
    layer7_outputs(2940) <= not (a or b);
    layer7_outputs(2941) <= not a;
    layer7_outputs(2942) <= not (a and b);
    layer7_outputs(2943) <= a;
    layer7_outputs(2944) <= a;
    layer7_outputs(2945) <= a or b;
    layer7_outputs(2946) <= b and not a;
    layer7_outputs(2947) <= a and b;
    layer7_outputs(2948) <= not (a or b);
    layer7_outputs(2949) <= a;
    layer7_outputs(2950) <= b;
    layer7_outputs(2951) <= b;
    layer7_outputs(2952) <= a;
    layer7_outputs(2953) <= b;
    layer7_outputs(2954) <= not b;
    layer7_outputs(2955) <= not a or b;
    layer7_outputs(2956) <= not (a and b);
    layer7_outputs(2957) <= not b;
    layer7_outputs(2958) <= a;
    layer7_outputs(2959) <= not (a and b);
    layer7_outputs(2960) <= a and b;
    layer7_outputs(2961) <= not b;
    layer7_outputs(2962) <= b;
    layer7_outputs(2963) <= not a;
    layer7_outputs(2964) <= a;
    layer7_outputs(2965) <= not b;
    layer7_outputs(2966) <= not (a or b);
    layer7_outputs(2967) <= not b;
    layer7_outputs(2968) <= a xor b;
    layer7_outputs(2969) <= b and not a;
    layer7_outputs(2970) <= not (a or b);
    layer7_outputs(2971) <= b and not a;
    layer7_outputs(2972) <= not b;
    layer7_outputs(2973) <= b;
    layer7_outputs(2974) <= a and b;
    layer7_outputs(2975) <= a xor b;
    layer7_outputs(2976) <= not (a xor b);
    layer7_outputs(2977) <= a;
    layer7_outputs(2978) <= a and not b;
    layer7_outputs(2979) <= a;
    layer7_outputs(2980) <= b and not a;
    layer7_outputs(2981) <= not a;
    layer7_outputs(2982) <= a xor b;
    layer7_outputs(2983) <= not (a or b);
    layer7_outputs(2984) <= not a or b;
    layer7_outputs(2985) <= not b or a;
    layer7_outputs(2986) <= not a;
    layer7_outputs(2987) <= not b;
    layer7_outputs(2988) <= not b or a;
    layer7_outputs(2989) <= b;
    layer7_outputs(2990) <= not (a xor b);
    layer7_outputs(2991) <= a;
    layer7_outputs(2992) <= a and b;
    layer7_outputs(2993) <= a and not b;
    layer7_outputs(2994) <= not a;
    layer7_outputs(2995) <= not (a or b);
    layer7_outputs(2996) <= a or b;
    layer7_outputs(2997) <= a;
    layer7_outputs(2998) <= not (a and b);
    layer7_outputs(2999) <= not (a and b);
    layer7_outputs(3000) <= b;
    layer7_outputs(3001) <= a and not b;
    layer7_outputs(3002) <= not a;
    layer7_outputs(3003) <= b;
    layer7_outputs(3004) <= not (a and b);
    layer7_outputs(3005) <= a xor b;
    layer7_outputs(3006) <= not b or a;
    layer7_outputs(3007) <= not a;
    layer7_outputs(3008) <= not b;
    layer7_outputs(3009) <= not b;
    layer7_outputs(3010) <= not b;
    layer7_outputs(3011) <= a and not b;
    layer7_outputs(3012) <= not b or a;
    layer7_outputs(3013) <= not b;
    layer7_outputs(3014) <= not b or a;
    layer7_outputs(3015) <= a;
    layer7_outputs(3016) <= b;
    layer7_outputs(3017) <= not a;
    layer7_outputs(3018) <= a xor b;
    layer7_outputs(3019) <= not (a xor b);
    layer7_outputs(3020) <= not (a or b);
    layer7_outputs(3021) <= b and not a;
    layer7_outputs(3022) <= not b;
    layer7_outputs(3023) <= b;
    layer7_outputs(3024) <= a;
    layer7_outputs(3025) <= not b;
    layer7_outputs(3026) <= a and not b;
    layer7_outputs(3027) <= not a;
    layer7_outputs(3028) <= b;
    layer7_outputs(3029) <= not a;
    layer7_outputs(3030) <= a and b;
    layer7_outputs(3031) <= not b or a;
    layer7_outputs(3032) <= not b;
    layer7_outputs(3033) <= not a;
    layer7_outputs(3034) <= not (a or b);
    layer7_outputs(3035) <= a and b;
    layer7_outputs(3036) <= a and not b;
    layer7_outputs(3037) <= b;
    layer7_outputs(3038) <= a and b;
    layer7_outputs(3039) <= b and not a;
    layer7_outputs(3040) <= b;
    layer7_outputs(3041) <= not b or a;
    layer7_outputs(3042) <= a and b;
    layer7_outputs(3043) <= a and not b;
    layer7_outputs(3044) <= b;
    layer7_outputs(3045) <= not (a and b);
    layer7_outputs(3046) <= a or b;
    layer7_outputs(3047) <= not (a xor b);
    layer7_outputs(3048) <= not (a and b);
    layer7_outputs(3049) <= not a;
    layer7_outputs(3050) <= not b or a;
    layer7_outputs(3051) <= a and not b;
    layer7_outputs(3052) <= a and not b;
    layer7_outputs(3053) <= a;
    layer7_outputs(3054) <= a;
    layer7_outputs(3055) <= a xor b;
    layer7_outputs(3056) <= b;
    layer7_outputs(3057) <= not b or a;
    layer7_outputs(3058) <= a and b;
    layer7_outputs(3059) <= b;
    layer7_outputs(3060) <= b and not a;
    layer7_outputs(3061) <= a or b;
    layer7_outputs(3062) <= a and not b;
    layer7_outputs(3063) <= not (a xor b);
    layer7_outputs(3064) <= a and b;
    layer7_outputs(3065) <= not b or a;
    layer7_outputs(3066) <= a;
    layer7_outputs(3067) <= not (a and b);
    layer7_outputs(3068) <= not b;
    layer7_outputs(3069) <= a and not b;
    layer7_outputs(3070) <= a and not b;
    layer7_outputs(3071) <= not a;
    layer7_outputs(3072) <= not a or b;
    layer7_outputs(3073) <= a;
    layer7_outputs(3074) <= a xor b;
    layer7_outputs(3075) <= a and not b;
    layer7_outputs(3076) <= not (a xor b);
    layer7_outputs(3077) <= a;
    layer7_outputs(3078) <= a and not b;
    layer7_outputs(3079) <= a and b;
    layer7_outputs(3080) <= a and b;
    layer7_outputs(3081) <= b and not a;
    layer7_outputs(3082) <= a;
    layer7_outputs(3083) <= a;
    layer7_outputs(3084) <= not (a and b);
    layer7_outputs(3085) <= a;
    layer7_outputs(3086) <= not (a and b);
    layer7_outputs(3087) <= a or b;
    layer7_outputs(3088) <= a xor b;
    layer7_outputs(3089) <= not b;
    layer7_outputs(3090) <= not (a xor b);
    layer7_outputs(3091) <= b;
    layer7_outputs(3092) <= not a;
    layer7_outputs(3093) <= b and not a;
    layer7_outputs(3094) <= not (a and b);
    layer7_outputs(3095) <= not a;
    layer7_outputs(3096) <= b and not a;
    layer7_outputs(3097) <= a xor b;
    layer7_outputs(3098) <= not (a and b);
    layer7_outputs(3099) <= a;
    layer7_outputs(3100) <= not b;
    layer7_outputs(3101) <= b;
    layer7_outputs(3102) <= not b or a;
    layer7_outputs(3103) <= a xor b;
    layer7_outputs(3104) <= b and not a;
    layer7_outputs(3105) <= not b;
    layer7_outputs(3106) <= b;
    layer7_outputs(3107) <= b;
    layer7_outputs(3108) <= a;
    layer7_outputs(3109) <= not a;
    layer7_outputs(3110) <= not b;
    layer7_outputs(3111) <= not b or a;
    layer7_outputs(3112) <= b;
    layer7_outputs(3113) <= not b;
    layer7_outputs(3114) <= a and b;
    layer7_outputs(3115) <= not a;
    layer7_outputs(3116) <= not (a and b);
    layer7_outputs(3117) <= a and not b;
    layer7_outputs(3118) <= a;
    layer7_outputs(3119) <= not a;
    layer7_outputs(3120) <= b;
    layer7_outputs(3121) <= a and not b;
    layer7_outputs(3122) <= not (a xor b);
    layer7_outputs(3123) <= a or b;
    layer7_outputs(3124) <= b and not a;
    layer7_outputs(3125) <= not a;
    layer7_outputs(3126) <= a xor b;
    layer7_outputs(3127) <= not (a and b);
    layer7_outputs(3128) <= not b or a;
    layer7_outputs(3129) <= a;
    layer7_outputs(3130) <= not b or a;
    layer7_outputs(3131) <= a xor b;
    layer7_outputs(3132) <= not a;
    layer7_outputs(3133) <= a and b;
    layer7_outputs(3134) <= not a;
    layer7_outputs(3135) <= '1';
    layer7_outputs(3136) <= not (a xor b);
    layer7_outputs(3137) <= not b;
    layer7_outputs(3138) <= not a;
    layer7_outputs(3139) <= a xor b;
    layer7_outputs(3140) <= not a;
    layer7_outputs(3141) <= not (a or b);
    layer7_outputs(3142) <= a;
    layer7_outputs(3143) <= a and not b;
    layer7_outputs(3144) <= not b;
    layer7_outputs(3145) <= b and not a;
    layer7_outputs(3146) <= not a or b;
    layer7_outputs(3147) <= not b;
    layer7_outputs(3148) <= a and not b;
    layer7_outputs(3149) <= not (a and b);
    layer7_outputs(3150) <= a;
    layer7_outputs(3151) <= not (a or b);
    layer7_outputs(3152) <= not (a or b);
    layer7_outputs(3153) <= a;
    layer7_outputs(3154) <= b;
    layer7_outputs(3155) <= not (a or b);
    layer7_outputs(3156) <= not b;
    layer7_outputs(3157) <= not (a and b);
    layer7_outputs(3158) <= a and not b;
    layer7_outputs(3159) <= not (a and b);
    layer7_outputs(3160) <= b;
    layer7_outputs(3161) <= not b or a;
    layer7_outputs(3162) <= not (a and b);
    layer7_outputs(3163) <= b;
    layer7_outputs(3164) <= not a;
    layer7_outputs(3165) <= b;
    layer7_outputs(3166) <= not b;
    layer7_outputs(3167) <= not (a and b);
    layer7_outputs(3168) <= not b;
    layer7_outputs(3169) <= b and not a;
    layer7_outputs(3170) <= not a;
    layer7_outputs(3171) <= not (a or b);
    layer7_outputs(3172) <= a and not b;
    layer7_outputs(3173) <= a xor b;
    layer7_outputs(3174) <= not b;
    layer7_outputs(3175) <= not b;
    layer7_outputs(3176) <= not (a xor b);
    layer7_outputs(3177) <= a;
    layer7_outputs(3178) <= a or b;
    layer7_outputs(3179) <= a;
    layer7_outputs(3180) <= not (a and b);
    layer7_outputs(3181) <= b and not a;
    layer7_outputs(3182) <= a;
    layer7_outputs(3183) <= b;
    layer7_outputs(3184) <= a or b;
    layer7_outputs(3185) <= b;
    layer7_outputs(3186) <= not a;
    layer7_outputs(3187) <= not b or a;
    layer7_outputs(3188) <= not (a xor b);
    layer7_outputs(3189) <= b and not a;
    layer7_outputs(3190) <= not (a xor b);
    layer7_outputs(3191) <= not (a xor b);
    layer7_outputs(3192) <= not b;
    layer7_outputs(3193) <= not (a and b);
    layer7_outputs(3194) <= not (a and b);
    layer7_outputs(3195) <= not a;
    layer7_outputs(3196) <= not a;
    layer7_outputs(3197) <= b;
    layer7_outputs(3198) <= b;
    layer7_outputs(3199) <= not a;
    layer7_outputs(3200) <= not b or a;
    layer7_outputs(3201) <= not b or a;
    layer7_outputs(3202) <= not b or a;
    layer7_outputs(3203) <= '1';
    layer7_outputs(3204) <= b;
    layer7_outputs(3205) <= a xor b;
    layer7_outputs(3206) <= a or b;
    layer7_outputs(3207) <= a;
    layer7_outputs(3208) <= not b;
    layer7_outputs(3209) <= a or b;
    layer7_outputs(3210) <= b;
    layer7_outputs(3211) <= not a;
    layer7_outputs(3212) <= a;
    layer7_outputs(3213) <= a and b;
    layer7_outputs(3214) <= '1';
    layer7_outputs(3215) <= b and not a;
    layer7_outputs(3216) <= a and b;
    layer7_outputs(3217) <= a and b;
    layer7_outputs(3218) <= '1';
    layer7_outputs(3219) <= b and not a;
    layer7_outputs(3220) <= a or b;
    layer7_outputs(3221) <= not a;
    layer7_outputs(3222) <= not a;
    layer7_outputs(3223) <= b and not a;
    layer7_outputs(3224) <= a;
    layer7_outputs(3225) <= a;
    layer7_outputs(3226) <= b;
    layer7_outputs(3227) <= a and not b;
    layer7_outputs(3228) <= a;
    layer7_outputs(3229) <= not b or a;
    layer7_outputs(3230) <= '0';
    layer7_outputs(3231) <= not b;
    layer7_outputs(3232) <= not a;
    layer7_outputs(3233) <= not a or b;
    layer7_outputs(3234) <= a;
    layer7_outputs(3235) <= not b;
    layer7_outputs(3236) <= a and not b;
    layer7_outputs(3237) <= not (a and b);
    layer7_outputs(3238) <= a;
    layer7_outputs(3239) <= b;
    layer7_outputs(3240) <= b;
    layer7_outputs(3241) <= not (a and b);
    layer7_outputs(3242) <= a and not b;
    layer7_outputs(3243) <= a;
    layer7_outputs(3244) <= not (a or b);
    layer7_outputs(3245) <= b;
    layer7_outputs(3246) <= a;
    layer7_outputs(3247) <= b and not a;
    layer7_outputs(3248) <= not (a or b);
    layer7_outputs(3249) <= a or b;
    layer7_outputs(3250) <= b;
    layer7_outputs(3251) <= not a;
    layer7_outputs(3252) <= a;
    layer7_outputs(3253) <= b;
    layer7_outputs(3254) <= not b;
    layer7_outputs(3255) <= a or b;
    layer7_outputs(3256) <= not b;
    layer7_outputs(3257) <= not (a and b);
    layer7_outputs(3258) <= not b or a;
    layer7_outputs(3259) <= not a;
    layer7_outputs(3260) <= not (a and b);
    layer7_outputs(3261) <= not b;
    layer7_outputs(3262) <= not (a xor b);
    layer7_outputs(3263) <= b and not a;
    layer7_outputs(3264) <= not b or a;
    layer7_outputs(3265) <= not b or a;
    layer7_outputs(3266) <= not a;
    layer7_outputs(3267) <= not b;
    layer7_outputs(3268) <= not (a xor b);
    layer7_outputs(3269) <= a and b;
    layer7_outputs(3270) <= a xor b;
    layer7_outputs(3271) <= not (a xor b);
    layer7_outputs(3272) <= a and not b;
    layer7_outputs(3273) <= not (a or b);
    layer7_outputs(3274) <= not (a xor b);
    layer7_outputs(3275) <= a;
    layer7_outputs(3276) <= not a;
    layer7_outputs(3277) <= a;
    layer7_outputs(3278) <= b and not a;
    layer7_outputs(3279) <= a;
    layer7_outputs(3280) <= b;
    layer7_outputs(3281) <= not a;
    layer7_outputs(3282) <= b;
    layer7_outputs(3283) <= not (a xor b);
    layer7_outputs(3284) <= b;
    layer7_outputs(3285) <= not b;
    layer7_outputs(3286) <= not b;
    layer7_outputs(3287) <= a xor b;
    layer7_outputs(3288) <= not b;
    layer7_outputs(3289) <= not (a or b);
    layer7_outputs(3290) <= a and b;
    layer7_outputs(3291) <= a xor b;
    layer7_outputs(3292) <= a and not b;
    layer7_outputs(3293) <= not (a xor b);
    layer7_outputs(3294) <= a and b;
    layer7_outputs(3295) <= a xor b;
    layer7_outputs(3296) <= not (a or b);
    layer7_outputs(3297) <= b and not a;
    layer7_outputs(3298) <= not a;
    layer7_outputs(3299) <= not (a and b);
    layer7_outputs(3300) <= a and b;
    layer7_outputs(3301) <= not a;
    layer7_outputs(3302) <= a or b;
    layer7_outputs(3303) <= not b;
    layer7_outputs(3304) <= b and not a;
    layer7_outputs(3305) <= b;
    layer7_outputs(3306) <= not a or b;
    layer7_outputs(3307) <= a and not b;
    layer7_outputs(3308) <= a and b;
    layer7_outputs(3309) <= a;
    layer7_outputs(3310) <= b;
    layer7_outputs(3311) <= not b;
    layer7_outputs(3312) <= not a;
    layer7_outputs(3313) <= a xor b;
    layer7_outputs(3314) <= not a;
    layer7_outputs(3315) <= a and b;
    layer7_outputs(3316) <= not (a and b);
    layer7_outputs(3317) <= a or b;
    layer7_outputs(3318) <= b and not a;
    layer7_outputs(3319) <= not (a and b);
    layer7_outputs(3320) <= not b;
    layer7_outputs(3321) <= not (a xor b);
    layer7_outputs(3322) <= not b;
    layer7_outputs(3323) <= not (a or b);
    layer7_outputs(3324) <= a;
    layer7_outputs(3325) <= a;
    layer7_outputs(3326) <= a;
    layer7_outputs(3327) <= b and not a;
    layer7_outputs(3328) <= not (a xor b);
    layer7_outputs(3329) <= not b;
    layer7_outputs(3330) <= a xor b;
    layer7_outputs(3331) <= a and b;
    layer7_outputs(3332) <= not a or b;
    layer7_outputs(3333) <= a and not b;
    layer7_outputs(3334) <= not a or b;
    layer7_outputs(3335) <= not (a and b);
    layer7_outputs(3336) <= not b;
    layer7_outputs(3337) <= not b;
    layer7_outputs(3338) <= not a;
    layer7_outputs(3339) <= not a or b;
    layer7_outputs(3340) <= not a;
    layer7_outputs(3341) <= a xor b;
    layer7_outputs(3342) <= b;
    layer7_outputs(3343) <= not b;
    layer7_outputs(3344) <= not (a or b);
    layer7_outputs(3345) <= not a or b;
    layer7_outputs(3346) <= b;
    layer7_outputs(3347) <= not (a and b);
    layer7_outputs(3348) <= b;
    layer7_outputs(3349) <= a;
    layer7_outputs(3350) <= not a or b;
    layer7_outputs(3351) <= a and b;
    layer7_outputs(3352) <= not b or a;
    layer7_outputs(3353) <= a and b;
    layer7_outputs(3354) <= a and not b;
    layer7_outputs(3355) <= not a or b;
    layer7_outputs(3356) <= a xor b;
    layer7_outputs(3357) <= not a or b;
    layer7_outputs(3358) <= not b or a;
    layer7_outputs(3359) <= not (a xor b);
    layer7_outputs(3360) <= b;
    layer7_outputs(3361) <= a xor b;
    layer7_outputs(3362) <= '1';
    layer7_outputs(3363) <= '1';
    layer7_outputs(3364) <= b;
    layer7_outputs(3365) <= not a or b;
    layer7_outputs(3366) <= a xor b;
    layer7_outputs(3367) <= a xor b;
    layer7_outputs(3368) <= b;
    layer7_outputs(3369) <= not (a xor b);
    layer7_outputs(3370) <= a;
    layer7_outputs(3371) <= not b or a;
    layer7_outputs(3372) <= not b;
    layer7_outputs(3373) <= not b;
    layer7_outputs(3374) <= a xor b;
    layer7_outputs(3375) <= b;
    layer7_outputs(3376) <= not b;
    layer7_outputs(3377) <= not b;
    layer7_outputs(3378) <= not a or b;
    layer7_outputs(3379) <= not a;
    layer7_outputs(3380) <= b;
    layer7_outputs(3381) <= b;
    layer7_outputs(3382) <= not a;
    layer7_outputs(3383) <= not (a xor b);
    layer7_outputs(3384) <= a and b;
    layer7_outputs(3385) <= not b;
    layer7_outputs(3386) <= b;
    layer7_outputs(3387) <= a and b;
    layer7_outputs(3388) <= '0';
    layer7_outputs(3389) <= b and not a;
    layer7_outputs(3390) <= a and b;
    layer7_outputs(3391) <= a;
    layer7_outputs(3392) <= a and not b;
    layer7_outputs(3393) <= not b or a;
    layer7_outputs(3394) <= a or b;
    layer7_outputs(3395) <= a;
    layer7_outputs(3396) <= not (a or b);
    layer7_outputs(3397) <= a xor b;
    layer7_outputs(3398) <= a or b;
    layer7_outputs(3399) <= not a;
    layer7_outputs(3400) <= not a or b;
    layer7_outputs(3401) <= b;
    layer7_outputs(3402) <= not (a and b);
    layer7_outputs(3403) <= not (a xor b);
    layer7_outputs(3404) <= not a or b;
    layer7_outputs(3405) <= a and b;
    layer7_outputs(3406) <= a xor b;
    layer7_outputs(3407) <= b;
    layer7_outputs(3408) <= not a;
    layer7_outputs(3409) <= not b;
    layer7_outputs(3410) <= not (a and b);
    layer7_outputs(3411) <= a;
    layer7_outputs(3412) <= b and not a;
    layer7_outputs(3413) <= not a or b;
    layer7_outputs(3414) <= a or b;
    layer7_outputs(3415) <= a;
    layer7_outputs(3416) <= a;
    layer7_outputs(3417) <= not b or a;
    layer7_outputs(3418) <= not (a and b);
    layer7_outputs(3419) <= a;
    layer7_outputs(3420) <= not a;
    layer7_outputs(3421) <= not b;
    layer7_outputs(3422) <= not b;
    layer7_outputs(3423) <= a;
    layer7_outputs(3424) <= not a or b;
    layer7_outputs(3425) <= not a;
    layer7_outputs(3426) <= not a;
    layer7_outputs(3427) <= a xor b;
    layer7_outputs(3428) <= not b;
    layer7_outputs(3429) <= a;
    layer7_outputs(3430) <= a;
    layer7_outputs(3431) <= a xor b;
    layer7_outputs(3432) <= not b;
    layer7_outputs(3433) <= not (a and b);
    layer7_outputs(3434) <= not a;
    layer7_outputs(3435) <= b;
    layer7_outputs(3436) <= not b or a;
    layer7_outputs(3437) <= '0';
    layer7_outputs(3438) <= not (a and b);
    layer7_outputs(3439) <= not (a and b);
    layer7_outputs(3440) <= a;
    layer7_outputs(3441) <= not b or a;
    layer7_outputs(3442) <= a or b;
    layer7_outputs(3443) <= not b or a;
    layer7_outputs(3444) <= not a;
    layer7_outputs(3445) <= b and not a;
    layer7_outputs(3446) <= a;
    layer7_outputs(3447) <= a and not b;
    layer7_outputs(3448) <= b;
    layer7_outputs(3449) <= a and b;
    layer7_outputs(3450) <= not (a or b);
    layer7_outputs(3451) <= b;
    layer7_outputs(3452) <= not (a or b);
    layer7_outputs(3453) <= not a;
    layer7_outputs(3454) <= a xor b;
    layer7_outputs(3455) <= not b;
    layer7_outputs(3456) <= not (a and b);
    layer7_outputs(3457) <= not b;
    layer7_outputs(3458) <= a and b;
    layer7_outputs(3459) <= not a;
    layer7_outputs(3460) <= not a or b;
    layer7_outputs(3461) <= not b or a;
    layer7_outputs(3462) <= not a;
    layer7_outputs(3463) <= a xor b;
    layer7_outputs(3464) <= not (a or b);
    layer7_outputs(3465) <= not (a and b);
    layer7_outputs(3466) <= b;
    layer7_outputs(3467) <= b and not a;
    layer7_outputs(3468) <= a or b;
    layer7_outputs(3469) <= not b or a;
    layer7_outputs(3470) <= a;
    layer7_outputs(3471) <= a xor b;
    layer7_outputs(3472) <= not (a or b);
    layer7_outputs(3473) <= not (a or b);
    layer7_outputs(3474) <= a;
    layer7_outputs(3475) <= not a;
    layer7_outputs(3476) <= a;
    layer7_outputs(3477) <= b;
    layer7_outputs(3478) <= b;
    layer7_outputs(3479) <= a and b;
    layer7_outputs(3480) <= not b;
    layer7_outputs(3481) <= not b;
    layer7_outputs(3482) <= not a;
    layer7_outputs(3483) <= not b;
    layer7_outputs(3484) <= a xor b;
    layer7_outputs(3485) <= a and not b;
    layer7_outputs(3486) <= not a or b;
    layer7_outputs(3487) <= not (a xor b);
    layer7_outputs(3488) <= a xor b;
    layer7_outputs(3489) <= not b;
    layer7_outputs(3490) <= a and b;
    layer7_outputs(3491) <= b;
    layer7_outputs(3492) <= not b;
    layer7_outputs(3493) <= a and b;
    layer7_outputs(3494) <= a and b;
    layer7_outputs(3495) <= not (a and b);
    layer7_outputs(3496) <= not b;
    layer7_outputs(3497) <= not b;
    layer7_outputs(3498) <= not a;
    layer7_outputs(3499) <= not b;
    layer7_outputs(3500) <= a;
    layer7_outputs(3501) <= b and not a;
    layer7_outputs(3502) <= a and not b;
    layer7_outputs(3503) <= a;
    layer7_outputs(3504) <= a;
    layer7_outputs(3505) <= not (a and b);
    layer7_outputs(3506) <= not (a and b);
    layer7_outputs(3507) <= b and not a;
    layer7_outputs(3508) <= not a or b;
    layer7_outputs(3509) <= a;
    layer7_outputs(3510) <= not (a xor b);
    layer7_outputs(3511) <= a xor b;
    layer7_outputs(3512) <= not b;
    layer7_outputs(3513) <= a;
    layer7_outputs(3514) <= not b;
    layer7_outputs(3515) <= not a;
    layer7_outputs(3516) <= not b or a;
    layer7_outputs(3517) <= not b;
    layer7_outputs(3518) <= a xor b;
    layer7_outputs(3519) <= not a;
    layer7_outputs(3520) <= b;
    layer7_outputs(3521) <= not b;
    layer7_outputs(3522) <= not a;
    layer7_outputs(3523) <= not (a xor b);
    layer7_outputs(3524) <= a or b;
    layer7_outputs(3525) <= not (a and b);
    layer7_outputs(3526) <= a;
    layer7_outputs(3527) <= a or b;
    layer7_outputs(3528) <= not a;
    layer7_outputs(3529) <= not b or a;
    layer7_outputs(3530) <= not a or b;
    layer7_outputs(3531) <= a or b;
    layer7_outputs(3532) <= not b;
    layer7_outputs(3533) <= a or b;
    layer7_outputs(3534) <= b and not a;
    layer7_outputs(3535) <= not (a xor b);
    layer7_outputs(3536) <= b;
    layer7_outputs(3537) <= not (a xor b);
    layer7_outputs(3538) <= not b;
    layer7_outputs(3539) <= not a or b;
    layer7_outputs(3540) <= not (a xor b);
    layer7_outputs(3541) <= a and not b;
    layer7_outputs(3542) <= not a;
    layer7_outputs(3543) <= b;
    layer7_outputs(3544) <= not a;
    layer7_outputs(3545) <= a;
    layer7_outputs(3546) <= a or b;
    layer7_outputs(3547) <= not (a xor b);
    layer7_outputs(3548) <= not b or a;
    layer7_outputs(3549) <= not (a or b);
    layer7_outputs(3550) <= a;
    layer7_outputs(3551) <= not b;
    layer7_outputs(3552) <= not (a xor b);
    layer7_outputs(3553) <= a or b;
    layer7_outputs(3554) <= not b;
    layer7_outputs(3555) <= not a;
    layer7_outputs(3556) <= b and not a;
    layer7_outputs(3557) <= not a;
    layer7_outputs(3558) <= not a or b;
    layer7_outputs(3559) <= not a;
    layer7_outputs(3560) <= b;
    layer7_outputs(3561) <= b and not a;
    layer7_outputs(3562) <= a;
    layer7_outputs(3563) <= not (a or b);
    layer7_outputs(3564) <= not (a xor b);
    layer7_outputs(3565) <= a;
    layer7_outputs(3566) <= not a;
    layer7_outputs(3567) <= a and b;
    layer7_outputs(3568) <= not b;
    layer7_outputs(3569) <= a and not b;
    layer7_outputs(3570) <= a;
    layer7_outputs(3571) <= not b;
    layer7_outputs(3572) <= a xor b;
    layer7_outputs(3573) <= not a;
    layer7_outputs(3574) <= a and b;
    layer7_outputs(3575) <= not a or b;
    layer7_outputs(3576) <= not b;
    layer7_outputs(3577) <= not (a and b);
    layer7_outputs(3578) <= not a;
    layer7_outputs(3579) <= a or b;
    layer7_outputs(3580) <= b and not a;
    layer7_outputs(3581) <= not (a xor b);
    layer7_outputs(3582) <= not (a or b);
    layer7_outputs(3583) <= b;
    layer7_outputs(3584) <= b;
    layer7_outputs(3585) <= a xor b;
    layer7_outputs(3586) <= a and b;
    layer7_outputs(3587) <= a or b;
    layer7_outputs(3588) <= a xor b;
    layer7_outputs(3589) <= not b;
    layer7_outputs(3590) <= a;
    layer7_outputs(3591) <= not (a xor b);
    layer7_outputs(3592) <= not b;
    layer7_outputs(3593) <= a and not b;
    layer7_outputs(3594) <= not b;
    layer7_outputs(3595) <= not (a xor b);
    layer7_outputs(3596) <= not (a or b);
    layer7_outputs(3597) <= not (a xor b);
    layer7_outputs(3598) <= '1';
    layer7_outputs(3599) <= a;
    layer7_outputs(3600) <= b;
    layer7_outputs(3601) <= a or b;
    layer7_outputs(3602) <= '0';
    layer7_outputs(3603) <= a xor b;
    layer7_outputs(3604) <= not (a and b);
    layer7_outputs(3605) <= not b;
    layer7_outputs(3606) <= not a or b;
    layer7_outputs(3607) <= not (a xor b);
    layer7_outputs(3608) <= b;
    layer7_outputs(3609) <= a xor b;
    layer7_outputs(3610) <= not (a xor b);
    layer7_outputs(3611) <= a;
    layer7_outputs(3612) <= not a or b;
    layer7_outputs(3613) <= b and not a;
    layer7_outputs(3614) <= a xor b;
    layer7_outputs(3615) <= a or b;
    layer7_outputs(3616) <= a;
    layer7_outputs(3617) <= a and not b;
    layer7_outputs(3618) <= not b;
    layer7_outputs(3619) <= a and b;
    layer7_outputs(3620) <= not (a and b);
    layer7_outputs(3621) <= a and not b;
    layer7_outputs(3622) <= not a or b;
    layer7_outputs(3623) <= not a;
    layer7_outputs(3624) <= not a or b;
    layer7_outputs(3625) <= not a or b;
    layer7_outputs(3626) <= a or b;
    layer7_outputs(3627) <= not b;
    layer7_outputs(3628) <= a and not b;
    layer7_outputs(3629) <= a;
    layer7_outputs(3630) <= '1';
    layer7_outputs(3631) <= not (a and b);
    layer7_outputs(3632) <= b;
    layer7_outputs(3633) <= a and b;
    layer7_outputs(3634) <= not b or a;
    layer7_outputs(3635) <= not (a or b);
    layer7_outputs(3636) <= a and not b;
    layer7_outputs(3637) <= not a;
    layer7_outputs(3638) <= not a;
    layer7_outputs(3639) <= a or b;
    layer7_outputs(3640) <= a or b;
    layer7_outputs(3641) <= b;
    layer7_outputs(3642) <= not a;
    layer7_outputs(3643) <= a xor b;
    layer7_outputs(3644) <= not b;
    layer7_outputs(3645) <= not (a or b);
    layer7_outputs(3646) <= not b;
    layer7_outputs(3647) <= not a;
    layer7_outputs(3648) <= not (a xor b);
    layer7_outputs(3649) <= not b;
    layer7_outputs(3650) <= not (a xor b);
    layer7_outputs(3651) <= not b or a;
    layer7_outputs(3652) <= not (a or b);
    layer7_outputs(3653) <= '0';
    layer7_outputs(3654) <= a xor b;
    layer7_outputs(3655) <= a and b;
    layer7_outputs(3656) <= not b or a;
    layer7_outputs(3657) <= not (a xor b);
    layer7_outputs(3658) <= not (a or b);
    layer7_outputs(3659) <= not a or b;
    layer7_outputs(3660) <= a;
    layer7_outputs(3661) <= a;
    layer7_outputs(3662) <= not (a or b);
    layer7_outputs(3663) <= a;
    layer7_outputs(3664) <= not a;
    layer7_outputs(3665) <= not (a xor b);
    layer7_outputs(3666) <= not b or a;
    layer7_outputs(3667) <= a;
    layer7_outputs(3668) <= b;
    layer7_outputs(3669) <= a;
    layer7_outputs(3670) <= not b;
    layer7_outputs(3671) <= b and not a;
    layer7_outputs(3672) <= not (a xor b);
    layer7_outputs(3673) <= not b;
    layer7_outputs(3674) <= a;
    layer7_outputs(3675) <= a xor b;
    layer7_outputs(3676) <= b;
    layer7_outputs(3677) <= b;
    layer7_outputs(3678) <= a xor b;
    layer7_outputs(3679) <= a;
    layer7_outputs(3680) <= not (a or b);
    layer7_outputs(3681) <= a and b;
    layer7_outputs(3682) <= a;
    layer7_outputs(3683) <= not b;
    layer7_outputs(3684) <= not (a and b);
    layer7_outputs(3685) <= not (a xor b);
    layer7_outputs(3686) <= a and not b;
    layer7_outputs(3687) <= not a;
    layer7_outputs(3688) <= not (a xor b);
    layer7_outputs(3689) <= a and b;
    layer7_outputs(3690) <= not a;
    layer7_outputs(3691) <= not b or a;
    layer7_outputs(3692) <= not a;
    layer7_outputs(3693) <= b;
    layer7_outputs(3694) <= not a;
    layer7_outputs(3695) <= not (a or b);
    layer7_outputs(3696) <= '1';
    layer7_outputs(3697) <= not b;
    layer7_outputs(3698) <= a;
    layer7_outputs(3699) <= b and not a;
    layer7_outputs(3700) <= b;
    layer7_outputs(3701) <= not (a xor b);
    layer7_outputs(3702) <= a;
    layer7_outputs(3703) <= a xor b;
    layer7_outputs(3704) <= a;
    layer7_outputs(3705) <= b;
    layer7_outputs(3706) <= a or b;
    layer7_outputs(3707) <= a and b;
    layer7_outputs(3708) <= b and not a;
    layer7_outputs(3709) <= a xor b;
    layer7_outputs(3710) <= a xor b;
    layer7_outputs(3711) <= a and b;
    layer7_outputs(3712) <= '1';
    layer7_outputs(3713) <= a and b;
    layer7_outputs(3714) <= a;
    layer7_outputs(3715) <= not (a xor b);
    layer7_outputs(3716) <= a or b;
    layer7_outputs(3717) <= not a;
    layer7_outputs(3718) <= b;
    layer7_outputs(3719) <= not a or b;
    layer7_outputs(3720) <= b and not a;
    layer7_outputs(3721) <= not a or b;
    layer7_outputs(3722) <= not a;
    layer7_outputs(3723) <= not (a or b);
    layer7_outputs(3724) <= b;
    layer7_outputs(3725) <= not b;
    layer7_outputs(3726) <= a;
    layer7_outputs(3727) <= not a;
    layer7_outputs(3728) <= '1';
    layer7_outputs(3729) <= a and b;
    layer7_outputs(3730) <= not b or a;
    layer7_outputs(3731) <= b and not a;
    layer7_outputs(3732) <= a xor b;
    layer7_outputs(3733) <= not a;
    layer7_outputs(3734) <= b;
    layer7_outputs(3735) <= a and not b;
    layer7_outputs(3736) <= not b;
    layer7_outputs(3737) <= a and not b;
    layer7_outputs(3738) <= a and not b;
    layer7_outputs(3739) <= a;
    layer7_outputs(3740) <= b;
    layer7_outputs(3741) <= a and not b;
    layer7_outputs(3742) <= a or b;
    layer7_outputs(3743) <= a;
    layer7_outputs(3744) <= a;
    layer7_outputs(3745) <= b;
    layer7_outputs(3746) <= not a or b;
    layer7_outputs(3747) <= not a;
    layer7_outputs(3748) <= not a or b;
    layer7_outputs(3749) <= not b;
    layer7_outputs(3750) <= b;
    layer7_outputs(3751) <= b;
    layer7_outputs(3752) <= a xor b;
    layer7_outputs(3753) <= a or b;
    layer7_outputs(3754) <= not b;
    layer7_outputs(3755) <= a and b;
    layer7_outputs(3756) <= not a;
    layer7_outputs(3757) <= not b;
    layer7_outputs(3758) <= b;
    layer7_outputs(3759) <= not a;
    layer7_outputs(3760) <= not (a and b);
    layer7_outputs(3761) <= not (a xor b);
    layer7_outputs(3762) <= b and not a;
    layer7_outputs(3763) <= b and not a;
    layer7_outputs(3764) <= a;
    layer7_outputs(3765) <= not a;
    layer7_outputs(3766) <= not b;
    layer7_outputs(3767) <= a xor b;
    layer7_outputs(3768) <= b;
    layer7_outputs(3769) <= not a;
    layer7_outputs(3770) <= b and not a;
    layer7_outputs(3771) <= not b;
    layer7_outputs(3772) <= b;
    layer7_outputs(3773) <= not b or a;
    layer7_outputs(3774) <= a and not b;
    layer7_outputs(3775) <= a;
    layer7_outputs(3776) <= a or b;
    layer7_outputs(3777) <= not (a xor b);
    layer7_outputs(3778) <= b;
    layer7_outputs(3779) <= b;
    layer7_outputs(3780) <= a xor b;
    layer7_outputs(3781) <= not (a xor b);
    layer7_outputs(3782) <= a or b;
    layer7_outputs(3783) <= a;
    layer7_outputs(3784) <= not b or a;
    layer7_outputs(3785) <= not (a xor b);
    layer7_outputs(3786) <= a;
    layer7_outputs(3787) <= not a;
    layer7_outputs(3788) <= a xor b;
    layer7_outputs(3789) <= a and b;
    layer7_outputs(3790) <= not (a and b);
    layer7_outputs(3791) <= not b or a;
    layer7_outputs(3792) <= a and b;
    layer7_outputs(3793) <= a and b;
    layer7_outputs(3794) <= a;
    layer7_outputs(3795) <= not a;
    layer7_outputs(3796) <= not (a xor b);
    layer7_outputs(3797) <= not (a and b);
    layer7_outputs(3798) <= not b;
    layer7_outputs(3799) <= a;
    layer7_outputs(3800) <= not (a or b);
    layer7_outputs(3801) <= not a;
    layer7_outputs(3802) <= not b or a;
    layer7_outputs(3803) <= not (a and b);
    layer7_outputs(3804) <= not a;
    layer7_outputs(3805) <= not a or b;
    layer7_outputs(3806) <= not b or a;
    layer7_outputs(3807) <= a xor b;
    layer7_outputs(3808) <= not b;
    layer7_outputs(3809) <= not b or a;
    layer7_outputs(3810) <= not (a or b);
    layer7_outputs(3811) <= not a;
    layer7_outputs(3812) <= a and not b;
    layer7_outputs(3813) <= a xor b;
    layer7_outputs(3814) <= a or b;
    layer7_outputs(3815) <= a;
    layer7_outputs(3816) <= a;
    layer7_outputs(3817) <= a;
    layer7_outputs(3818) <= not b or a;
    layer7_outputs(3819) <= '1';
    layer7_outputs(3820) <= not (a xor b);
    layer7_outputs(3821) <= b;
    layer7_outputs(3822) <= a or b;
    layer7_outputs(3823) <= a or b;
    layer7_outputs(3824) <= a and b;
    layer7_outputs(3825) <= b;
    layer7_outputs(3826) <= not a or b;
    layer7_outputs(3827) <= b;
    layer7_outputs(3828) <= not b;
    layer7_outputs(3829) <= not b or a;
    layer7_outputs(3830) <= b and not a;
    layer7_outputs(3831) <= b and not a;
    layer7_outputs(3832) <= a or b;
    layer7_outputs(3833) <= not b or a;
    layer7_outputs(3834) <= a;
    layer7_outputs(3835) <= a or b;
    layer7_outputs(3836) <= not (a or b);
    layer7_outputs(3837) <= b;
    layer7_outputs(3838) <= not b;
    layer7_outputs(3839) <= not a;
    layer7_outputs(3840) <= a or b;
    layer7_outputs(3841) <= a or b;
    layer7_outputs(3842) <= not a;
    layer7_outputs(3843) <= not a;
    layer7_outputs(3844) <= not b;
    layer7_outputs(3845) <= a or b;
    layer7_outputs(3846) <= a xor b;
    layer7_outputs(3847) <= a xor b;
    layer7_outputs(3848) <= not (a and b);
    layer7_outputs(3849) <= b;
    layer7_outputs(3850) <= a xor b;
    layer7_outputs(3851) <= a or b;
    layer7_outputs(3852) <= b;
    layer7_outputs(3853) <= not a;
    layer7_outputs(3854) <= b;
    layer7_outputs(3855) <= a and b;
    layer7_outputs(3856) <= a or b;
    layer7_outputs(3857) <= not b;
    layer7_outputs(3858) <= not a or b;
    layer7_outputs(3859) <= b and not a;
    layer7_outputs(3860) <= b and not a;
    layer7_outputs(3861) <= not b or a;
    layer7_outputs(3862) <= not (a and b);
    layer7_outputs(3863) <= a and not b;
    layer7_outputs(3864) <= a xor b;
    layer7_outputs(3865) <= not b;
    layer7_outputs(3866) <= a;
    layer7_outputs(3867) <= a;
    layer7_outputs(3868) <= not b;
    layer7_outputs(3869) <= not b or a;
    layer7_outputs(3870) <= b;
    layer7_outputs(3871) <= not (a or b);
    layer7_outputs(3872) <= a or b;
    layer7_outputs(3873) <= not a;
    layer7_outputs(3874) <= not a or b;
    layer7_outputs(3875) <= not a or b;
    layer7_outputs(3876) <= b and not a;
    layer7_outputs(3877) <= '1';
    layer7_outputs(3878) <= not (a and b);
    layer7_outputs(3879) <= not (a xor b);
    layer7_outputs(3880) <= not (a xor b);
    layer7_outputs(3881) <= not (a xor b);
    layer7_outputs(3882) <= not a or b;
    layer7_outputs(3883) <= b and not a;
    layer7_outputs(3884) <= b and not a;
    layer7_outputs(3885) <= not a;
    layer7_outputs(3886) <= not a;
    layer7_outputs(3887) <= a and b;
    layer7_outputs(3888) <= not a;
    layer7_outputs(3889) <= not (a and b);
    layer7_outputs(3890) <= a and not b;
    layer7_outputs(3891) <= a or b;
    layer7_outputs(3892) <= a;
    layer7_outputs(3893) <= not a;
    layer7_outputs(3894) <= a;
    layer7_outputs(3895) <= not b;
    layer7_outputs(3896) <= not b;
    layer7_outputs(3897) <= not (a or b);
    layer7_outputs(3898) <= a and not b;
    layer7_outputs(3899) <= not a;
    layer7_outputs(3900) <= not b;
    layer7_outputs(3901) <= not b;
    layer7_outputs(3902) <= not a or b;
    layer7_outputs(3903) <= not b or a;
    layer7_outputs(3904) <= a and b;
    layer7_outputs(3905) <= a xor b;
    layer7_outputs(3906) <= a;
    layer7_outputs(3907) <= not b;
    layer7_outputs(3908) <= not a;
    layer7_outputs(3909) <= not b;
    layer7_outputs(3910) <= a xor b;
    layer7_outputs(3911) <= a xor b;
    layer7_outputs(3912) <= not a or b;
    layer7_outputs(3913) <= not a;
    layer7_outputs(3914) <= not b;
    layer7_outputs(3915) <= b;
    layer7_outputs(3916) <= b and not a;
    layer7_outputs(3917) <= a;
    layer7_outputs(3918) <= a or b;
    layer7_outputs(3919) <= not (a or b);
    layer7_outputs(3920) <= not b or a;
    layer7_outputs(3921) <= not (a xor b);
    layer7_outputs(3922) <= b;
    layer7_outputs(3923) <= a;
    layer7_outputs(3924) <= not b;
    layer7_outputs(3925) <= b and not a;
    layer7_outputs(3926) <= a xor b;
    layer7_outputs(3927) <= '1';
    layer7_outputs(3928) <= a;
    layer7_outputs(3929) <= not (a xor b);
    layer7_outputs(3930) <= a or b;
    layer7_outputs(3931) <= not a;
    layer7_outputs(3932) <= not a;
    layer7_outputs(3933) <= '0';
    layer7_outputs(3934) <= a or b;
    layer7_outputs(3935) <= not a;
    layer7_outputs(3936) <= not a;
    layer7_outputs(3937) <= not (a xor b);
    layer7_outputs(3938) <= a;
    layer7_outputs(3939) <= b;
    layer7_outputs(3940) <= not (a xor b);
    layer7_outputs(3941) <= not b;
    layer7_outputs(3942) <= b and not a;
    layer7_outputs(3943) <= not (a or b);
    layer7_outputs(3944) <= not (a or b);
    layer7_outputs(3945) <= not a;
    layer7_outputs(3946) <= not a;
    layer7_outputs(3947) <= b;
    layer7_outputs(3948) <= b;
    layer7_outputs(3949) <= b;
    layer7_outputs(3950) <= not b;
    layer7_outputs(3951) <= b;
    layer7_outputs(3952) <= b;
    layer7_outputs(3953) <= not (a and b);
    layer7_outputs(3954) <= a xor b;
    layer7_outputs(3955) <= not (a or b);
    layer7_outputs(3956) <= a or b;
    layer7_outputs(3957) <= not (a or b);
    layer7_outputs(3958) <= not b;
    layer7_outputs(3959) <= a xor b;
    layer7_outputs(3960) <= not a;
    layer7_outputs(3961) <= not b;
    layer7_outputs(3962) <= not a or b;
    layer7_outputs(3963) <= a xor b;
    layer7_outputs(3964) <= not b or a;
    layer7_outputs(3965) <= a;
    layer7_outputs(3966) <= a;
    layer7_outputs(3967) <= not b;
    layer7_outputs(3968) <= a and b;
    layer7_outputs(3969) <= a;
    layer7_outputs(3970) <= not b or a;
    layer7_outputs(3971) <= a or b;
    layer7_outputs(3972) <= not a or b;
    layer7_outputs(3973) <= a or b;
    layer7_outputs(3974) <= a;
    layer7_outputs(3975) <= not a;
    layer7_outputs(3976) <= a or b;
    layer7_outputs(3977) <= not b or a;
    layer7_outputs(3978) <= a and not b;
    layer7_outputs(3979) <= '0';
    layer7_outputs(3980) <= not b;
    layer7_outputs(3981) <= not b;
    layer7_outputs(3982) <= not b;
    layer7_outputs(3983) <= not (a and b);
    layer7_outputs(3984) <= a;
    layer7_outputs(3985) <= not b or a;
    layer7_outputs(3986) <= not a;
    layer7_outputs(3987) <= not (a or b);
    layer7_outputs(3988) <= not (a xor b);
    layer7_outputs(3989) <= not b;
    layer7_outputs(3990) <= a and b;
    layer7_outputs(3991) <= not a;
    layer7_outputs(3992) <= a;
    layer7_outputs(3993) <= not (a xor b);
    layer7_outputs(3994) <= not (a and b);
    layer7_outputs(3995) <= b and not a;
    layer7_outputs(3996) <= b;
    layer7_outputs(3997) <= a and b;
    layer7_outputs(3998) <= not b or a;
    layer7_outputs(3999) <= not b or a;
    layer7_outputs(4000) <= not (a xor b);
    layer7_outputs(4001) <= not b or a;
    layer7_outputs(4002) <= a and b;
    layer7_outputs(4003) <= b;
    layer7_outputs(4004) <= b and not a;
    layer7_outputs(4005) <= not a;
    layer7_outputs(4006) <= not b;
    layer7_outputs(4007) <= not (a and b);
    layer7_outputs(4008) <= b and not a;
    layer7_outputs(4009) <= a or b;
    layer7_outputs(4010) <= not (a or b);
    layer7_outputs(4011) <= not b;
    layer7_outputs(4012) <= not b;
    layer7_outputs(4013) <= a and not b;
    layer7_outputs(4014) <= not a;
    layer7_outputs(4015) <= not (a and b);
    layer7_outputs(4016) <= not b;
    layer7_outputs(4017) <= a;
    layer7_outputs(4018) <= not (a and b);
    layer7_outputs(4019) <= '1';
    layer7_outputs(4020) <= a and b;
    layer7_outputs(4021) <= b;
    layer7_outputs(4022) <= not b or a;
    layer7_outputs(4023) <= not b;
    layer7_outputs(4024) <= a xor b;
    layer7_outputs(4025) <= b;
    layer7_outputs(4026) <= a;
    layer7_outputs(4027) <= not b;
    layer7_outputs(4028) <= a and b;
    layer7_outputs(4029) <= not (a and b);
    layer7_outputs(4030) <= not b;
    layer7_outputs(4031) <= a xor b;
    layer7_outputs(4032) <= a;
    layer7_outputs(4033) <= b;
    layer7_outputs(4034) <= b;
    layer7_outputs(4035) <= a and b;
    layer7_outputs(4036) <= not b or a;
    layer7_outputs(4037) <= a;
    layer7_outputs(4038) <= a or b;
    layer7_outputs(4039) <= a;
    layer7_outputs(4040) <= '1';
    layer7_outputs(4041) <= not b;
    layer7_outputs(4042) <= b;
    layer7_outputs(4043) <= not (a or b);
    layer7_outputs(4044) <= not (a xor b);
    layer7_outputs(4045) <= b;
    layer7_outputs(4046) <= not b;
    layer7_outputs(4047) <= not b;
    layer7_outputs(4048) <= a xor b;
    layer7_outputs(4049) <= not (a and b);
    layer7_outputs(4050) <= not b;
    layer7_outputs(4051) <= not b or a;
    layer7_outputs(4052) <= not (a and b);
    layer7_outputs(4053) <= not (a xor b);
    layer7_outputs(4054) <= not (a xor b);
    layer7_outputs(4055) <= a or b;
    layer7_outputs(4056) <= not (a and b);
    layer7_outputs(4057) <= a;
    layer7_outputs(4058) <= not b or a;
    layer7_outputs(4059) <= not (a xor b);
    layer7_outputs(4060) <= not (a and b);
    layer7_outputs(4061) <= not a;
    layer7_outputs(4062) <= b;
    layer7_outputs(4063) <= b;
    layer7_outputs(4064) <= not b;
    layer7_outputs(4065) <= not (a and b);
    layer7_outputs(4066) <= a;
    layer7_outputs(4067) <= not a or b;
    layer7_outputs(4068) <= a xor b;
    layer7_outputs(4069) <= b and not a;
    layer7_outputs(4070) <= not a;
    layer7_outputs(4071) <= not a or b;
    layer7_outputs(4072) <= b and not a;
    layer7_outputs(4073) <= not b;
    layer7_outputs(4074) <= a xor b;
    layer7_outputs(4075) <= not a or b;
    layer7_outputs(4076) <= not b;
    layer7_outputs(4077) <= not b;
    layer7_outputs(4078) <= not a;
    layer7_outputs(4079) <= not (a or b);
    layer7_outputs(4080) <= b;
    layer7_outputs(4081) <= not b;
    layer7_outputs(4082) <= a and not b;
    layer7_outputs(4083) <= not a;
    layer7_outputs(4084) <= not b or a;
    layer7_outputs(4085) <= not (a or b);
    layer7_outputs(4086) <= not (a xor b);
    layer7_outputs(4087) <= not a;
    layer7_outputs(4088) <= b;
    layer7_outputs(4089) <= not a;
    layer7_outputs(4090) <= a;
    layer7_outputs(4091) <= not (a and b);
    layer7_outputs(4092) <= not (a or b);
    layer7_outputs(4093) <= a;
    layer7_outputs(4094) <= not b;
    layer7_outputs(4095) <= a and b;
    layer7_outputs(4096) <= a;
    layer7_outputs(4097) <= a or b;
    layer7_outputs(4098) <= b;
    layer7_outputs(4099) <= b;
    layer7_outputs(4100) <= a and b;
    layer7_outputs(4101) <= b;
    layer7_outputs(4102) <= not b or a;
    layer7_outputs(4103) <= not (a xor b);
    layer7_outputs(4104) <= not b or a;
    layer7_outputs(4105) <= b and not a;
    layer7_outputs(4106) <= b;
    layer7_outputs(4107) <= not b or a;
    layer7_outputs(4108) <= not (a and b);
    layer7_outputs(4109) <= a;
    layer7_outputs(4110) <= a or b;
    layer7_outputs(4111) <= '1';
    layer7_outputs(4112) <= b;
    layer7_outputs(4113) <= not a or b;
    layer7_outputs(4114) <= a and not b;
    layer7_outputs(4115) <= a or b;
    layer7_outputs(4116) <= a and b;
    layer7_outputs(4117) <= not b;
    layer7_outputs(4118) <= a;
    layer7_outputs(4119) <= a and b;
    layer7_outputs(4120) <= a xor b;
    layer7_outputs(4121) <= not b or a;
    layer7_outputs(4122) <= not (a and b);
    layer7_outputs(4123) <= '0';
    layer7_outputs(4124) <= b and not a;
    layer7_outputs(4125) <= a and b;
    layer7_outputs(4126) <= b and not a;
    layer7_outputs(4127) <= a and not b;
    layer7_outputs(4128) <= not a or b;
    layer7_outputs(4129) <= not b;
    layer7_outputs(4130) <= not b or a;
    layer7_outputs(4131) <= not (a xor b);
    layer7_outputs(4132) <= a xor b;
    layer7_outputs(4133) <= not (a and b);
    layer7_outputs(4134) <= not b;
    layer7_outputs(4135) <= not a;
    layer7_outputs(4136) <= not (a or b);
    layer7_outputs(4137) <= a and b;
    layer7_outputs(4138) <= a or b;
    layer7_outputs(4139) <= b and not a;
    layer7_outputs(4140) <= b;
    layer7_outputs(4141) <= a and b;
    layer7_outputs(4142) <= a xor b;
    layer7_outputs(4143) <= not (a or b);
    layer7_outputs(4144) <= not (a xor b);
    layer7_outputs(4145) <= not a or b;
    layer7_outputs(4146) <= not b or a;
    layer7_outputs(4147) <= not a or b;
    layer7_outputs(4148) <= a or b;
    layer7_outputs(4149) <= a and not b;
    layer7_outputs(4150) <= not (a and b);
    layer7_outputs(4151) <= not (a and b);
    layer7_outputs(4152) <= a;
    layer7_outputs(4153) <= '1';
    layer7_outputs(4154) <= b;
    layer7_outputs(4155) <= not b or a;
    layer7_outputs(4156) <= not b;
    layer7_outputs(4157) <= not b;
    layer7_outputs(4158) <= a xor b;
    layer7_outputs(4159) <= b;
    layer7_outputs(4160) <= not (a xor b);
    layer7_outputs(4161) <= a xor b;
    layer7_outputs(4162) <= a;
    layer7_outputs(4163) <= not b;
    layer7_outputs(4164) <= not b or a;
    layer7_outputs(4165) <= b;
    layer7_outputs(4166) <= not a;
    layer7_outputs(4167) <= not a;
    layer7_outputs(4168) <= b and not a;
    layer7_outputs(4169) <= not (a xor b);
    layer7_outputs(4170) <= not (a and b);
    layer7_outputs(4171) <= a and not b;
    layer7_outputs(4172) <= b and not a;
    layer7_outputs(4173) <= a;
    layer7_outputs(4174) <= not (a xor b);
    layer7_outputs(4175) <= not (a and b);
    layer7_outputs(4176) <= not (a or b);
    layer7_outputs(4177) <= a;
    layer7_outputs(4178) <= b;
    layer7_outputs(4179) <= a;
    layer7_outputs(4180) <= a and not b;
    layer7_outputs(4181) <= a and not b;
    layer7_outputs(4182) <= not (a and b);
    layer7_outputs(4183) <= a and b;
    layer7_outputs(4184) <= not b;
    layer7_outputs(4185) <= a;
    layer7_outputs(4186) <= not a or b;
    layer7_outputs(4187) <= not (a xor b);
    layer7_outputs(4188) <= not a or b;
    layer7_outputs(4189) <= a;
    layer7_outputs(4190) <= a and b;
    layer7_outputs(4191) <= not (a xor b);
    layer7_outputs(4192) <= not a;
    layer7_outputs(4193) <= not (a and b);
    layer7_outputs(4194) <= not (a xor b);
    layer7_outputs(4195) <= not a;
    layer7_outputs(4196) <= a;
    layer7_outputs(4197) <= a xor b;
    layer7_outputs(4198) <= a or b;
    layer7_outputs(4199) <= not b;
    layer7_outputs(4200) <= a and b;
    layer7_outputs(4201) <= not a or b;
    layer7_outputs(4202) <= a or b;
    layer7_outputs(4203) <= b;
    layer7_outputs(4204) <= not b;
    layer7_outputs(4205) <= '0';
    layer7_outputs(4206) <= '0';
    layer7_outputs(4207) <= b and not a;
    layer7_outputs(4208) <= b;
    layer7_outputs(4209) <= not b;
    layer7_outputs(4210) <= not b;
    layer7_outputs(4211) <= not b;
    layer7_outputs(4212) <= not (a and b);
    layer7_outputs(4213) <= not b;
    layer7_outputs(4214) <= not a;
    layer7_outputs(4215) <= a or b;
    layer7_outputs(4216) <= a or b;
    layer7_outputs(4217) <= not b;
    layer7_outputs(4218) <= not (a xor b);
    layer7_outputs(4219) <= a or b;
    layer7_outputs(4220) <= not (a xor b);
    layer7_outputs(4221) <= not a or b;
    layer7_outputs(4222) <= a;
    layer7_outputs(4223) <= a;
    layer7_outputs(4224) <= not a or b;
    layer7_outputs(4225) <= not (a xor b);
    layer7_outputs(4226) <= not a;
    layer7_outputs(4227) <= not a;
    layer7_outputs(4228) <= not b or a;
    layer7_outputs(4229) <= a;
    layer7_outputs(4230) <= not (a or b);
    layer7_outputs(4231) <= a or b;
    layer7_outputs(4232) <= not (a or b);
    layer7_outputs(4233) <= a or b;
    layer7_outputs(4234) <= not a;
    layer7_outputs(4235) <= a xor b;
    layer7_outputs(4236) <= not (a and b);
    layer7_outputs(4237) <= a;
    layer7_outputs(4238) <= not b;
    layer7_outputs(4239) <= a;
    layer7_outputs(4240) <= b;
    layer7_outputs(4241) <= not a;
    layer7_outputs(4242) <= a and b;
    layer7_outputs(4243) <= not (a xor b);
    layer7_outputs(4244) <= not b;
    layer7_outputs(4245) <= not (a or b);
    layer7_outputs(4246) <= not (a or b);
    layer7_outputs(4247) <= not a;
    layer7_outputs(4248) <= a;
    layer7_outputs(4249) <= not b or a;
    layer7_outputs(4250) <= a xor b;
    layer7_outputs(4251) <= a and not b;
    layer7_outputs(4252) <= not (a and b);
    layer7_outputs(4253) <= not b or a;
    layer7_outputs(4254) <= not a;
    layer7_outputs(4255) <= '0';
    layer7_outputs(4256) <= a;
    layer7_outputs(4257) <= not a;
    layer7_outputs(4258) <= not (a and b);
    layer7_outputs(4259) <= b;
    layer7_outputs(4260) <= a xor b;
    layer7_outputs(4261) <= a and b;
    layer7_outputs(4262) <= not b;
    layer7_outputs(4263) <= b and not a;
    layer7_outputs(4264) <= a;
    layer7_outputs(4265) <= a xor b;
    layer7_outputs(4266) <= b;
    layer7_outputs(4267) <= a xor b;
    layer7_outputs(4268) <= b;
    layer7_outputs(4269) <= a or b;
    layer7_outputs(4270) <= b;
    layer7_outputs(4271) <= not a;
    layer7_outputs(4272) <= not a;
    layer7_outputs(4273) <= not b;
    layer7_outputs(4274) <= not b;
    layer7_outputs(4275) <= a;
    layer7_outputs(4276) <= not b or a;
    layer7_outputs(4277) <= not (a or b);
    layer7_outputs(4278) <= not a;
    layer7_outputs(4279) <= not (a or b);
    layer7_outputs(4280) <= b;
    layer7_outputs(4281) <= b;
    layer7_outputs(4282) <= not (a or b);
    layer7_outputs(4283) <= a and not b;
    layer7_outputs(4284) <= not (a and b);
    layer7_outputs(4285) <= b;
    layer7_outputs(4286) <= not b;
    layer7_outputs(4287) <= a and b;
    layer7_outputs(4288) <= a or b;
    layer7_outputs(4289) <= not (a and b);
    layer7_outputs(4290) <= b;
    layer7_outputs(4291) <= not (a xor b);
    layer7_outputs(4292) <= a and b;
    layer7_outputs(4293) <= a;
    layer7_outputs(4294) <= not b;
    layer7_outputs(4295) <= a xor b;
    layer7_outputs(4296) <= not a;
    layer7_outputs(4297) <= not a;
    layer7_outputs(4298) <= not (a xor b);
    layer7_outputs(4299) <= not a;
    layer7_outputs(4300) <= a and b;
    layer7_outputs(4301) <= not (a xor b);
    layer7_outputs(4302) <= b and not a;
    layer7_outputs(4303) <= not a;
    layer7_outputs(4304) <= a;
    layer7_outputs(4305) <= not a;
    layer7_outputs(4306) <= not a or b;
    layer7_outputs(4307) <= a and not b;
    layer7_outputs(4308) <= b;
    layer7_outputs(4309) <= a;
    layer7_outputs(4310) <= not b;
    layer7_outputs(4311) <= b;
    layer7_outputs(4312) <= not a or b;
    layer7_outputs(4313) <= not (a xor b);
    layer7_outputs(4314) <= b and not a;
    layer7_outputs(4315) <= b and not a;
    layer7_outputs(4316) <= a;
    layer7_outputs(4317) <= a;
    layer7_outputs(4318) <= not (a xor b);
    layer7_outputs(4319) <= a and not b;
    layer7_outputs(4320) <= b and not a;
    layer7_outputs(4321) <= a or b;
    layer7_outputs(4322) <= b;
    layer7_outputs(4323) <= b and not a;
    layer7_outputs(4324) <= not b;
    layer7_outputs(4325) <= not a or b;
    layer7_outputs(4326) <= not (a and b);
    layer7_outputs(4327) <= not b;
    layer7_outputs(4328) <= not b;
    layer7_outputs(4329) <= not a or b;
    layer7_outputs(4330) <= b and not a;
    layer7_outputs(4331) <= not b;
    layer7_outputs(4332) <= not a;
    layer7_outputs(4333) <= b;
    layer7_outputs(4334) <= not b or a;
    layer7_outputs(4335) <= a;
    layer7_outputs(4336) <= b;
    layer7_outputs(4337) <= not b or a;
    layer7_outputs(4338) <= b;
    layer7_outputs(4339) <= b and not a;
    layer7_outputs(4340) <= not a or b;
    layer7_outputs(4341) <= b;
    layer7_outputs(4342) <= a or b;
    layer7_outputs(4343) <= a;
    layer7_outputs(4344) <= b and not a;
    layer7_outputs(4345) <= a or b;
    layer7_outputs(4346) <= not a;
    layer7_outputs(4347) <= not (a xor b);
    layer7_outputs(4348) <= not a;
    layer7_outputs(4349) <= not a;
    layer7_outputs(4350) <= not b;
    layer7_outputs(4351) <= not a or b;
    layer7_outputs(4352) <= not b;
    layer7_outputs(4353) <= a and not b;
    layer7_outputs(4354) <= a;
    layer7_outputs(4355) <= a xor b;
    layer7_outputs(4356) <= a and not b;
    layer7_outputs(4357) <= not (a and b);
    layer7_outputs(4358) <= b;
    layer7_outputs(4359) <= not a;
    layer7_outputs(4360) <= a and b;
    layer7_outputs(4361) <= b;
    layer7_outputs(4362) <= '1';
    layer7_outputs(4363) <= not a;
    layer7_outputs(4364) <= not (a xor b);
    layer7_outputs(4365) <= b and not a;
    layer7_outputs(4366) <= b and not a;
    layer7_outputs(4367) <= not b;
    layer7_outputs(4368) <= not b;
    layer7_outputs(4369) <= a and not b;
    layer7_outputs(4370) <= a and b;
    layer7_outputs(4371) <= not a;
    layer7_outputs(4372) <= not (a or b);
    layer7_outputs(4373) <= not a;
    layer7_outputs(4374) <= a;
    layer7_outputs(4375) <= not b or a;
    layer7_outputs(4376) <= a and b;
    layer7_outputs(4377) <= b;
    layer7_outputs(4378) <= a;
    layer7_outputs(4379) <= b;
    layer7_outputs(4380) <= not (a xor b);
    layer7_outputs(4381) <= not (a and b);
    layer7_outputs(4382) <= not b;
    layer7_outputs(4383) <= b and not a;
    layer7_outputs(4384) <= not (a and b);
    layer7_outputs(4385) <= a xor b;
    layer7_outputs(4386) <= not b or a;
    layer7_outputs(4387) <= a;
    layer7_outputs(4388) <= a xor b;
    layer7_outputs(4389) <= a xor b;
    layer7_outputs(4390) <= a or b;
    layer7_outputs(4391) <= b;
    layer7_outputs(4392) <= a;
    layer7_outputs(4393) <= a;
    layer7_outputs(4394) <= not a;
    layer7_outputs(4395) <= a xor b;
    layer7_outputs(4396) <= a xor b;
    layer7_outputs(4397) <= a;
    layer7_outputs(4398) <= a and b;
    layer7_outputs(4399) <= a and b;
    layer7_outputs(4400) <= a;
    layer7_outputs(4401) <= a;
    layer7_outputs(4402) <= not b;
    layer7_outputs(4403) <= a;
    layer7_outputs(4404) <= a and not b;
    layer7_outputs(4405) <= not a or b;
    layer7_outputs(4406) <= not b;
    layer7_outputs(4407) <= a and not b;
    layer7_outputs(4408) <= not a;
    layer7_outputs(4409) <= a;
    layer7_outputs(4410) <= not a or b;
    layer7_outputs(4411) <= a;
    layer7_outputs(4412) <= a;
    layer7_outputs(4413) <= b;
    layer7_outputs(4414) <= not (a or b);
    layer7_outputs(4415) <= not a or b;
    layer7_outputs(4416) <= not (a or b);
    layer7_outputs(4417) <= not (a xor b);
    layer7_outputs(4418) <= not b or a;
    layer7_outputs(4419) <= b;
    layer7_outputs(4420) <= a and not b;
    layer7_outputs(4421) <= not b;
    layer7_outputs(4422) <= a or b;
    layer7_outputs(4423) <= b and not a;
    layer7_outputs(4424) <= not a or b;
    layer7_outputs(4425) <= a xor b;
    layer7_outputs(4426) <= a and not b;
    layer7_outputs(4427) <= not a;
    layer7_outputs(4428) <= '0';
    layer7_outputs(4429) <= a and not b;
    layer7_outputs(4430) <= not b;
    layer7_outputs(4431) <= not (a xor b);
    layer7_outputs(4432) <= not a;
    layer7_outputs(4433) <= a xor b;
    layer7_outputs(4434) <= b;
    layer7_outputs(4435) <= a;
    layer7_outputs(4436) <= a and b;
    layer7_outputs(4437) <= b and not a;
    layer7_outputs(4438) <= not (a or b);
    layer7_outputs(4439) <= not (a xor b);
    layer7_outputs(4440) <= not a or b;
    layer7_outputs(4441) <= not a;
    layer7_outputs(4442) <= a;
    layer7_outputs(4443) <= not a;
    layer7_outputs(4444) <= a and b;
    layer7_outputs(4445) <= b;
    layer7_outputs(4446) <= b and not a;
    layer7_outputs(4447) <= a;
    layer7_outputs(4448) <= a and not b;
    layer7_outputs(4449) <= not a;
    layer7_outputs(4450) <= not a;
    layer7_outputs(4451) <= not (a xor b);
    layer7_outputs(4452) <= not a;
    layer7_outputs(4453) <= b and not a;
    layer7_outputs(4454) <= a;
    layer7_outputs(4455) <= b;
    layer7_outputs(4456) <= not a or b;
    layer7_outputs(4457) <= not a;
    layer7_outputs(4458) <= not (a xor b);
    layer7_outputs(4459) <= '0';
    layer7_outputs(4460) <= a or b;
    layer7_outputs(4461) <= a and b;
    layer7_outputs(4462) <= not b;
    layer7_outputs(4463) <= a;
    layer7_outputs(4464) <= a xor b;
    layer7_outputs(4465) <= b;
    layer7_outputs(4466) <= not a or b;
    layer7_outputs(4467) <= a and b;
    layer7_outputs(4468) <= not b;
    layer7_outputs(4469) <= not a;
    layer7_outputs(4470) <= not b;
    layer7_outputs(4471) <= not (a and b);
    layer7_outputs(4472) <= not a or b;
    layer7_outputs(4473) <= b and not a;
    layer7_outputs(4474) <= not b;
    layer7_outputs(4475) <= not b or a;
    layer7_outputs(4476) <= not b;
    layer7_outputs(4477) <= a and b;
    layer7_outputs(4478) <= not (a or b);
    layer7_outputs(4479) <= a;
    layer7_outputs(4480) <= not (a xor b);
    layer7_outputs(4481) <= a and b;
    layer7_outputs(4482) <= not a;
    layer7_outputs(4483) <= not b;
    layer7_outputs(4484) <= a xor b;
    layer7_outputs(4485) <= not a;
    layer7_outputs(4486) <= b;
    layer7_outputs(4487) <= b;
    layer7_outputs(4488) <= not b;
    layer7_outputs(4489) <= b;
    layer7_outputs(4490) <= a and b;
    layer7_outputs(4491) <= a;
    layer7_outputs(4492) <= not b;
    layer7_outputs(4493) <= b and not a;
    layer7_outputs(4494) <= not b or a;
    layer7_outputs(4495) <= a xor b;
    layer7_outputs(4496) <= not b;
    layer7_outputs(4497) <= not (a xor b);
    layer7_outputs(4498) <= a xor b;
    layer7_outputs(4499) <= a xor b;
    layer7_outputs(4500) <= not a or b;
    layer7_outputs(4501) <= not (a xor b);
    layer7_outputs(4502) <= a or b;
    layer7_outputs(4503) <= not (a xor b);
    layer7_outputs(4504) <= a xor b;
    layer7_outputs(4505) <= '0';
    layer7_outputs(4506) <= b;
    layer7_outputs(4507) <= a;
    layer7_outputs(4508) <= not (a xor b);
    layer7_outputs(4509) <= not (a or b);
    layer7_outputs(4510) <= not (a or b);
    layer7_outputs(4511) <= b;
    layer7_outputs(4512) <= a and not b;
    layer7_outputs(4513) <= not a or b;
    layer7_outputs(4514) <= b;
    layer7_outputs(4515) <= not (a and b);
    layer7_outputs(4516) <= not b;
    layer7_outputs(4517) <= not (a xor b);
    layer7_outputs(4518) <= a and not b;
    layer7_outputs(4519) <= a;
    layer7_outputs(4520) <= a;
    layer7_outputs(4521) <= not b;
    layer7_outputs(4522) <= a xor b;
    layer7_outputs(4523) <= not b;
    layer7_outputs(4524) <= a;
    layer7_outputs(4525) <= a or b;
    layer7_outputs(4526) <= not (a or b);
    layer7_outputs(4527) <= not (a xor b);
    layer7_outputs(4528) <= '1';
    layer7_outputs(4529) <= a xor b;
    layer7_outputs(4530) <= a and b;
    layer7_outputs(4531) <= a;
    layer7_outputs(4532) <= not a;
    layer7_outputs(4533) <= a;
    layer7_outputs(4534) <= b;
    layer7_outputs(4535) <= not (a or b);
    layer7_outputs(4536) <= not b or a;
    layer7_outputs(4537) <= not b;
    layer7_outputs(4538) <= b and not a;
    layer7_outputs(4539) <= a;
    layer7_outputs(4540) <= not a;
    layer7_outputs(4541) <= not b;
    layer7_outputs(4542) <= a;
    layer7_outputs(4543) <= not (a xor b);
    layer7_outputs(4544) <= a and b;
    layer7_outputs(4545) <= not b;
    layer7_outputs(4546) <= not (a and b);
    layer7_outputs(4547) <= not (a xor b);
    layer7_outputs(4548) <= not b;
    layer7_outputs(4549) <= a xor b;
    layer7_outputs(4550) <= not b or a;
    layer7_outputs(4551) <= not (a xor b);
    layer7_outputs(4552) <= b;
    layer7_outputs(4553) <= not a;
    layer7_outputs(4554) <= b;
    layer7_outputs(4555) <= a and b;
    layer7_outputs(4556) <= b;
    layer7_outputs(4557) <= not b or a;
    layer7_outputs(4558) <= a or b;
    layer7_outputs(4559) <= b and not a;
    layer7_outputs(4560) <= a xor b;
    layer7_outputs(4561) <= not (a or b);
    layer7_outputs(4562) <= b;
    layer7_outputs(4563) <= not b;
    layer7_outputs(4564) <= b and not a;
    layer7_outputs(4565) <= a xor b;
    layer7_outputs(4566) <= not (a and b);
    layer7_outputs(4567) <= a;
    layer7_outputs(4568) <= not b;
    layer7_outputs(4569) <= not a;
    layer7_outputs(4570) <= a xor b;
    layer7_outputs(4571) <= a and b;
    layer7_outputs(4572) <= not b or a;
    layer7_outputs(4573) <= not (a and b);
    layer7_outputs(4574) <= a;
    layer7_outputs(4575) <= not (a or b);
    layer7_outputs(4576) <= a or b;
    layer7_outputs(4577) <= b and not a;
    layer7_outputs(4578) <= a;
    layer7_outputs(4579) <= b;
    layer7_outputs(4580) <= not a;
    layer7_outputs(4581) <= not a;
    layer7_outputs(4582) <= not (a xor b);
    layer7_outputs(4583) <= not (a or b);
    layer7_outputs(4584) <= b;
    layer7_outputs(4585) <= a and b;
    layer7_outputs(4586) <= a xor b;
    layer7_outputs(4587) <= not (a or b);
    layer7_outputs(4588) <= a and b;
    layer7_outputs(4589) <= a xor b;
    layer7_outputs(4590) <= a and not b;
    layer7_outputs(4591) <= not b;
    layer7_outputs(4592) <= a and b;
    layer7_outputs(4593) <= b;
    layer7_outputs(4594) <= a and b;
    layer7_outputs(4595) <= a xor b;
    layer7_outputs(4596) <= not a;
    layer7_outputs(4597) <= b;
    layer7_outputs(4598) <= a and not b;
    layer7_outputs(4599) <= b;
    layer7_outputs(4600) <= a and b;
    layer7_outputs(4601) <= a and not b;
    layer7_outputs(4602) <= not b;
    layer7_outputs(4603) <= a;
    layer7_outputs(4604) <= not (a xor b);
    layer7_outputs(4605) <= a xor b;
    layer7_outputs(4606) <= not b;
    layer7_outputs(4607) <= not b;
    layer7_outputs(4608) <= not a;
    layer7_outputs(4609) <= a or b;
    layer7_outputs(4610) <= a or b;
    layer7_outputs(4611) <= not (a and b);
    layer7_outputs(4612) <= a;
    layer7_outputs(4613) <= not b;
    layer7_outputs(4614) <= a;
    layer7_outputs(4615) <= not (a xor b);
    layer7_outputs(4616) <= not (a and b);
    layer7_outputs(4617) <= a and not b;
    layer7_outputs(4618) <= not a;
    layer7_outputs(4619) <= b and not a;
    layer7_outputs(4620) <= a and b;
    layer7_outputs(4621) <= not a;
    layer7_outputs(4622) <= '0';
    layer7_outputs(4623) <= not a or b;
    layer7_outputs(4624) <= a xor b;
    layer7_outputs(4625) <= a;
    layer7_outputs(4626) <= b;
    layer7_outputs(4627) <= a and b;
    layer7_outputs(4628) <= a or b;
    layer7_outputs(4629) <= not a;
    layer7_outputs(4630) <= b;
    layer7_outputs(4631) <= not (a or b);
    layer7_outputs(4632) <= not b or a;
    layer7_outputs(4633) <= not b;
    layer7_outputs(4634) <= a;
    layer7_outputs(4635) <= b;
    layer7_outputs(4636) <= not (a xor b);
    layer7_outputs(4637) <= not b;
    layer7_outputs(4638) <= not (a xor b);
    layer7_outputs(4639) <= a xor b;
    layer7_outputs(4640) <= not (a xor b);
    layer7_outputs(4641) <= a;
    layer7_outputs(4642) <= a xor b;
    layer7_outputs(4643) <= a;
    layer7_outputs(4644) <= b and not a;
    layer7_outputs(4645) <= not a;
    layer7_outputs(4646) <= a xor b;
    layer7_outputs(4647) <= not b;
    layer7_outputs(4648) <= not (a and b);
    layer7_outputs(4649) <= not (a and b);
    layer7_outputs(4650) <= not (a and b);
    layer7_outputs(4651) <= a xor b;
    layer7_outputs(4652) <= a and b;
    layer7_outputs(4653) <= a;
    layer7_outputs(4654) <= not a;
    layer7_outputs(4655) <= not a;
    layer7_outputs(4656) <= a;
    layer7_outputs(4657) <= not (a xor b);
    layer7_outputs(4658) <= '0';
    layer7_outputs(4659) <= b;
    layer7_outputs(4660) <= a;
    layer7_outputs(4661) <= a;
    layer7_outputs(4662) <= not (a and b);
    layer7_outputs(4663) <= not b or a;
    layer7_outputs(4664) <= not a;
    layer7_outputs(4665) <= a and b;
    layer7_outputs(4666) <= not a;
    layer7_outputs(4667) <= not b or a;
    layer7_outputs(4668) <= not b;
    layer7_outputs(4669) <= not a;
    layer7_outputs(4670) <= not b or a;
    layer7_outputs(4671) <= not a;
    layer7_outputs(4672) <= a and not b;
    layer7_outputs(4673) <= not a;
    layer7_outputs(4674) <= a and not b;
    layer7_outputs(4675) <= a and b;
    layer7_outputs(4676) <= not a;
    layer7_outputs(4677) <= a xor b;
    layer7_outputs(4678) <= a xor b;
    layer7_outputs(4679) <= b;
    layer7_outputs(4680) <= a xor b;
    layer7_outputs(4681) <= not (a and b);
    layer7_outputs(4682) <= not a;
    layer7_outputs(4683) <= a;
    layer7_outputs(4684) <= a;
    layer7_outputs(4685) <= not b;
    layer7_outputs(4686) <= not a;
    layer7_outputs(4687) <= a;
    layer7_outputs(4688) <= b;
    layer7_outputs(4689) <= not b;
    layer7_outputs(4690) <= not (a and b);
    layer7_outputs(4691) <= not a;
    layer7_outputs(4692) <= not b;
    layer7_outputs(4693) <= not b or a;
    layer7_outputs(4694) <= not a or b;
    layer7_outputs(4695) <= not a or b;
    layer7_outputs(4696) <= a;
    layer7_outputs(4697) <= not (a and b);
    layer7_outputs(4698) <= a or b;
    layer7_outputs(4699) <= not a or b;
    layer7_outputs(4700) <= a or b;
    layer7_outputs(4701) <= a xor b;
    layer7_outputs(4702) <= b;
    layer7_outputs(4703) <= '1';
    layer7_outputs(4704) <= '0';
    layer7_outputs(4705) <= b and not a;
    layer7_outputs(4706) <= b;
    layer7_outputs(4707) <= b;
    layer7_outputs(4708) <= not a;
    layer7_outputs(4709) <= a xor b;
    layer7_outputs(4710) <= a or b;
    layer7_outputs(4711) <= a or b;
    layer7_outputs(4712) <= not (a xor b);
    layer7_outputs(4713) <= a and b;
    layer7_outputs(4714) <= a;
    layer7_outputs(4715) <= b;
    layer7_outputs(4716) <= b;
    layer7_outputs(4717) <= a or b;
    layer7_outputs(4718) <= a;
    layer7_outputs(4719) <= a;
    layer7_outputs(4720) <= not b or a;
    layer7_outputs(4721) <= b;
    layer7_outputs(4722) <= not b;
    layer7_outputs(4723) <= not (a and b);
    layer7_outputs(4724) <= b and not a;
    layer7_outputs(4725) <= not a;
    layer7_outputs(4726) <= a or b;
    layer7_outputs(4727) <= b;
    layer7_outputs(4728) <= b and not a;
    layer7_outputs(4729) <= not a;
    layer7_outputs(4730) <= a;
    layer7_outputs(4731) <= b and not a;
    layer7_outputs(4732) <= not (a and b);
    layer7_outputs(4733) <= a and not b;
    layer7_outputs(4734) <= a and b;
    layer7_outputs(4735) <= a xor b;
    layer7_outputs(4736) <= not (a and b);
    layer7_outputs(4737) <= not b or a;
    layer7_outputs(4738) <= b and not a;
    layer7_outputs(4739) <= not (a and b);
    layer7_outputs(4740) <= not b or a;
    layer7_outputs(4741) <= not a;
    layer7_outputs(4742) <= a and b;
    layer7_outputs(4743) <= not (a xor b);
    layer7_outputs(4744) <= not a or b;
    layer7_outputs(4745) <= a or b;
    layer7_outputs(4746) <= b and not a;
    layer7_outputs(4747) <= not b;
    layer7_outputs(4748) <= not a;
    layer7_outputs(4749) <= not (a or b);
    layer7_outputs(4750) <= not b or a;
    layer7_outputs(4751) <= a or b;
    layer7_outputs(4752) <= a xor b;
    layer7_outputs(4753) <= a xor b;
    layer7_outputs(4754) <= '1';
    layer7_outputs(4755) <= a and not b;
    layer7_outputs(4756) <= a and b;
    layer7_outputs(4757) <= not a;
    layer7_outputs(4758) <= a and b;
    layer7_outputs(4759) <= not a or b;
    layer7_outputs(4760) <= not (a or b);
    layer7_outputs(4761) <= a;
    layer7_outputs(4762) <= a;
    layer7_outputs(4763) <= not b;
    layer7_outputs(4764) <= not (a and b);
    layer7_outputs(4765) <= not (a xor b);
    layer7_outputs(4766) <= not a;
    layer7_outputs(4767) <= not b;
    layer7_outputs(4768) <= a and not b;
    layer7_outputs(4769) <= a xor b;
    layer7_outputs(4770) <= b;
    layer7_outputs(4771) <= not (a or b);
    layer7_outputs(4772) <= b;
    layer7_outputs(4773) <= b;
    layer7_outputs(4774) <= a;
    layer7_outputs(4775) <= not (a xor b);
    layer7_outputs(4776) <= not a or b;
    layer7_outputs(4777) <= not a;
    layer7_outputs(4778) <= not a;
    layer7_outputs(4779) <= a and b;
    layer7_outputs(4780) <= not a;
    layer7_outputs(4781) <= not b;
    layer7_outputs(4782) <= not b;
    layer7_outputs(4783) <= b;
    layer7_outputs(4784) <= not b or a;
    layer7_outputs(4785) <= a;
    layer7_outputs(4786) <= not a or b;
    layer7_outputs(4787) <= not a or b;
    layer7_outputs(4788) <= not a;
    layer7_outputs(4789) <= not a;
    layer7_outputs(4790) <= a xor b;
    layer7_outputs(4791) <= not a;
    layer7_outputs(4792) <= not b or a;
    layer7_outputs(4793) <= not (a xor b);
    layer7_outputs(4794) <= a and not b;
    layer7_outputs(4795) <= a xor b;
    layer7_outputs(4796) <= a and not b;
    layer7_outputs(4797) <= b;
    layer7_outputs(4798) <= '1';
    layer7_outputs(4799) <= not a;
    layer7_outputs(4800) <= not a;
    layer7_outputs(4801) <= a and not b;
    layer7_outputs(4802) <= a and b;
    layer7_outputs(4803) <= not b;
    layer7_outputs(4804) <= a xor b;
    layer7_outputs(4805) <= not (a or b);
    layer7_outputs(4806) <= not (a or b);
    layer7_outputs(4807) <= not b;
    layer7_outputs(4808) <= not b;
    layer7_outputs(4809) <= a;
    layer7_outputs(4810) <= not a or b;
    layer7_outputs(4811) <= a;
    layer7_outputs(4812) <= not (a and b);
    layer7_outputs(4813) <= not (a and b);
    layer7_outputs(4814) <= not a;
    layer7_outputs(4815) <= a;
    layer7_outputs(4816) <= a or b;
    layer7_outputs(4817) <= not b;
    layer7_outputs(4818) <= not (a xor b);
    layer7_outputs(4819) <= a;
    layer7_outputs(4820) <= a;
    layer7_outputs(4821) <= not b;
    layer7_outputs(4822) <= not b;
    layer7_outputs(4823) <= b;
    layer7_outputs(4824) <= b;
    layer7_outputs(4825) <= a and b;
    layer7_outputs(4826) <= not (a xor b);
    layer7_outputs(4827) <= not b;
    layer7_outputs(4828) <= not b;
    layer7_outputs(4829) <= not b;
    layer7_outputs(4830) <= b;
    layer7_outputs(4831) <= not a or b;
    layer7_outputs(4832) <= not (a and b);
    layer7_outputs(4833) <= a or b;
    layer7_outputs(4834) <= a;
    layer7_outputs(4835) <= a xor b;
    layer7_outputs(4836) <= a and not b;
    layer7_outputs(4837) <= not a or b;
    layer7_outputs(4838) <= not (a or b);
    layer7_outputs(4839) <= not b or a;
    layer7_outputs(4840) <= a;
    layer7_outputs(4841) <= b and not a;
    layer7_outputs(4842) <= not b;
    layer7_outputs(4843) <= not b;
    layer7_outputs(4844) <= not (a xor b);
    layer7_outputs(4845) <= a;
    layer7_outputs(4846) <= a and b;
    layer7_outputs(4847) <= '0';
    layer7_outputs(4848) <= not b;
    layer7_outputs(4849) <= not b;
    layer7_outputs(4850) <= not b;
    layer7_outputs(4851) <= a and not b;
    layer7_outputs(4852) <= not b or a;
    layer7_outputs(4853) <= not (a xor b);
    layer7_outputs(4854) <= not a or b;
    layer7_outputs(4855) <= a xor b;
    layer7_outputs(4856) <= not (a or b);
    layer7_outputs(4857) <= a;
    layer7_outputs(4858) <= not b;
    layer7_outputs(4859) <= a xor b;
    layer7_outputs(4860) <= a;
    layer7_outputs(4861) <= a;
    layer7_outputs(4862) <= '0';
    layer7_outputs(4863) <= not b;
    layer7_outputs(4864) <= a;
    layer7_outputs(4865) <= not a or b;
    layer7_outputs(4866) <= a or b;
    layer7_outputs(4867) <= not b;
    layer7_outputs(4868) <= b;
    layer7_outputs(4869) <= not b;
    layer7_outputs(4870) <= not a or b;
    layer7_outputs(4871) <= a xor b;
    layer7_outputs(4872) <= not a or b;
    layer7_outputs(4873) <= a or b;
    layer7_outputs(4874) <= not (a or b);
    layer7_outputs(4875) <= not (a xor b);
    layer7_outputs(4876) <= not a;
    layer7_outputs(4877) <= not (a xor b);
    layer7_outputs(4878) <= not a;
    layer7_outputs(4879) <= not a;
    layer7_outputs(4880) <= a xor b;
    layer7_outputs(4881) <= not b or a;
    layer7_outputs(4882) <= a and not b;
    layer7_outputs(4883) <= a xor b;
    layer7_outputs(4884) <= not b or a;
    layer7_outputs(4885) <= not b or a;
    layer7_outputs(4886) <= b;
    layer7_outputs(4887) <= a;
    layer7_outputs(4888) <= a or b;
    layer7_outputs(4889) <= not (a xor b);
    layer7_outputs(4890) <= not (a and b);
    layer7_outputs(4891) <= not a;
    layer7_outputs(4892) <= not b;
    layer7_outputs(4893) <= b and not a;
    layer7_outputs(4894) <= b and not a;
    layer7_outputs(4895) <= a and not b;
    layer7_outputs(4896) <= not (a xor b);
    layer7_outputs(4897) <= b;
    layer7_outputs(4898) <= not (a and b);
    layer7_outputs(4899) <= not b or a;
    layer7_outputs(4900) <= b;
    layer7_outputs(4901) <= a or b;
    layer7_outputs(4902) <= not (a or b);
    layer7_outputs(4903) <= b;
    layer7_outputs(4904) <= a or b;
    layer7_outputs(4905) <= a and b;
    layer7_outputs(4906) <= not a;
    layer7_outputs(4907) <= not (a or b);
    layer7_outputs(4908) <= a;
    layer7_outputs(4909) <= not (a or b);
    layer7_outputs(4910) <= a;
    layer7_outputs(4911) <= not b;
    layer7_outputs(4912) <= not (a xor b);
    layer7_outputs(4913) <= not b;
    layer7_outputs(4914) <= b;
    layer7_outputs(4915) <= a and b;
    layer7_outputs(4916) <= not (a xor b);
    layer7_outputs(4917) <= a;
    layer7_outputs(4918) <= not a;
    layer7_outputs(4919) <= a xor b;
    layer7_outputs(4920) <= not a;
    layer7_outputs(4921) <= a xor b;
    layer7_outputs(4922) <= '0';
    layer7_outputs(4923) <= a or b;
    layer7_outputs(4924) <= not (a or b);
    layer7_outputs(4925) <= not b;
    layer7_outputs(4926) <= not a or b;
    layer7_outputs(4927) <= not b;
    layer7_outputs(4928) <= a and not b;
    layer7_outputs(4929) <= not b;
    layer7_outputs(4930) <= a and not b;
    layer7_outputs(4931) <= not (a and b);
    layer7_outputs(4932) <= not (a and b);
    layer7_outputs(4933) <= not b;
    layer7_outputs(4934) <= not (a and b);
    layer7_outputs(4935) <= a and not b;
    layer7_outputs(4936) <= not b or a;
    layer7_outputs(4937) <= not b or a;
    layer7_outputs(4938) <= not (a or b);
    layer7_outputs(4939) <= not b;
    layer7_outputs(4940) <= not b;
    layer7_outputs(4941) <= b and not a;
    layer7_outputs(4942) <= b and not a;
    layer7_outputs(4943) <= not a or b;
    layer7_outputs(4944) <= not a;
    layer7_outputs(4945) <= not a;
    layer7_outputs(4946) <= not a;
    layer7_outputs(4947) <= a and not b;
    layer7_outputs(4948) <= a or b;
    layer7_outputs(4949) <= b;
    layer7_outputs(4950) <= a;
    layer7_outputs(4951) <= not a;
    layer7_outputs(4952) <= not (a or b);
    layer7_outputs(4953) <= a;
    layer7_outputs(4954) <= '0';
    layer7_outputs(4955) <= not b;
    layer7_outputs(4956) <= not a;
    layer7_outputs(4957) <= a xor b;
    layer7_outputs(4958) <= b;
    layer7_outputs(4959) <= b and not a;
    layer7_outputs(4960) <= not a;
    layer7_outputs(4961) <= not (a and b);
    layer7_outputs(4962) <= b;
    layer7_outputs(4963) <= not b or a;
    layer7_outputs(4964) <= '0';
    layer7_outputs(4965) <= not (a or b);
    layer7_outputs(4966) <= a xor b;
    layer7_outputs(4967) <= not a or b;
    layer7_outputs(4968) <= a and not b;
    layer7_outputs(4969) <= not b or a;
    layer7_outputs(4970) <= not (a and b);
    layer7_outputs(4971) <= a and not b;
    layer7_outputs(4972) <= not b;
    layer7_outputs(4973) <= a;
    layer7_outputs(4974) <= not b;
    layer7_outputs(4975) <= not b;
    layer7_outputs(4976) <= a;
    layer7_outputs(4977) <= a and b;
    layer7_outputs(4978) <= a and b;
    layer7_outputs(4979) <= not b;
    layer7_outputs(4980) <= a or b;
    layer7_outputs(4981) <= not a;
    layer7_outputs(4982) <= not b;
    layer7_outputs(4983) <= not b;
    layer7_outputs(4984) <= not b or a;
    layer7_outputs(4985) <= b;
    layer7_outputs(4986) <= not b;
    layer7_outputs(4987) <= '0';
    layer7_outputs(4988) <= not (a and b);
    layer7_outputs(4989) <= not a or b;
    layer7_outputs(4990) <= a or b;
    layer7_outputs(4991) <= '1';
    layer7_outputs(4992) <= b and not a;
    layer7_outputs(4993) <= not a or b;
    layer7_outputs(4994) <= b;
    layer7_outputs(4995) <= b and not a;
    layer7_outputs(4996) <= not a;
    layer7_outputs(4997) <= b;
    layer7_outputs(4998) <= a;
    layer7_outputs(4999) <= b and not a;
    layer7_outputs(5000) <= not a or b;
    layer7_outputs(5001) <= a;
    layer7_outputs(5002) <= a;
    layer7_outputs(5003) <= b;
    layer7_outputs(5004) <= a and b;
    layer7_outputs(5005) <= not a;
    layer7_outputs(5006) <= a and b;
    layer7_outputs(5007) <= not a or b;
    layer7_outputs(5008) <= a xor b;
    layer7_outputs(5009) <= '0';
    layer7_outputs(5010) <= not (a xor b);
    layer7_outputs(5011) <= not (a xor b);
    layer7_outputs(5012) <= not a;
    layer7_outputs(5013) <= a or b;
    layer7_outputs(5014) <= a xor b;
    layer7_outputs(5015) <= not (a xor b);
    layer7_outputs(5016) <= not (a or b);
    layer7_outputs(5017) <= not a;
    layer7_outputs(5018) <= not (a and b);
    layer7_outputs(5019) <= not a;
    layer7_outputs(5020) <= not (a and b);
    layer7_outputs(5021) <= b and not a;
    layer7_outputs(5022) <= a and not b;
    layer7_outputs(5023) <= a and not b;
    layer7_outputs(5024) <= not b or a;
    layer7_outputs(5025) <= not a;
    layer7_outputs(5026) <= not (a and b);
    layer7_outputs(5027) <= not (a xor b);
    layer7_outputs(5028) <= b;
    layer7_outputs(5029) <= not a or b;
    layer7_outputs(5030) <= not b;
    layer7_outputs(5031) <= not (a xor b);
    layer7_outputs(5032) <= a;
    layer7_outputs(5033) <= a;
    layer7_outputs(5034) <= not (a and b);
    layer7_outputs(5035) <= not a;
    layer7_outputs(5036) <= not a or b;
    layer7_outputs(5037) <= a xor b;
    layer7_outputs(5038) <= a;
    layer7_outputs(5039) <= not a;
    layer7_outputs(5040) <= not b;
    layer7_outputs(5041) <= not a;
    layer7_outputs(5042) <= a;
    layer7_outputs(5043) <= not a;
    layer7_outputs(5044) <= b;
    layer7_outputs(5045) <= a and b;
    layer7_outputs(5046) <= a;
    layer7_outputs(5047) <= not a;
    layer7_outputs(5048) <= not (a and b);
    layer7_outputs(5049) <= a or b;
    layer7_outputs(5050) <= a;
    layer7_outputs(5051) <= not a;
    layer7_outputs(5052) <= not a;
    layer7_outputs(5053) <= a;
    layer7_outputs(5054) <= a xor b;
    layer7_outputs(5055) <= not (a xor b);
    layer7_outputs(5056) <= '0';
    layer7_outputs(5057) <= not a;
    layer7_outputs(5058) <= a xor b;
    layer7_outputs(5059) <= b and not a;
    layer7_outputs(5060) <= not b;
    layer7_outputs(5061) <= not a or b;
    layer7_outputs(5062) <= not (a xor b);
    layer7_outputs(5063) <= a xor b;
    layer7_outputs(5064) <= a;
    layer7_outputs(5065) <= b;
    layer7_outputs(5066) <= not b;
    layer7_outputs(5067) <= a and not b;
    layer7_outputs(5068) <= not b or a;
    layer7_outputs(5069) <= not a;
    layer7_outputs(5070) <= a;
    layer7_outputs(5071) <= a and b;
    layer7_outputs(5072) <= a xor b;
    layer7_outputs(5073) <= not (a xor b);
    layer7_outputs(5074) <= a xor b;
    layer7_outputs(5075) <= not b;
    layer7_outputs(5076) <= a xor b;
    layer7_outputs(5077) <= b and not a;
    layer7_outputs(5078) <= a and b;
    layer7_outputs(5079) <= b and not a;
    layer7_outputs(5080) <= not b or a;
    layer7_outputs(5081) <= b;
    layer7_outputs(5082) <= not a;
    layer7_outputs(5083) <= not a or b;
    layer7_outputs(5084) <= b;
    layer7_outputs(5085) <= not a;
    layer7_outputs(5086) <= b and not a;
    layer7_outputs(5087) <= not (a or b);
    layer7_outputs(5088) <= b;
    layer7_outputs(5089) <= a;
    layer7_outputs(5090) <= b;
    layer7_outputs(5091) <= '1';
    layer7_outputs(5092) <= not b;
    layer7_outputs(5093) <= not (a xor b);
    layer7_outputs(5094) <= a and b;
    layer7_outputs(5095) <= not a;
    layer7_outputs(5096) <= '0';
    layer7_outputs(5097) <= not a;
    layer7_outputs(5098) <= a and b;
    layer7_outputs(5099) <= a xor b;
    layer7_outputs(5100) <= b;
    layer7_outputs(5101) <= a;
    layer7_outputs(5102) <= b and not a;
    layer7_outputs(5103) <= b;
    layer7_outputs(5104) <= not b;
    layer7_outputs(5105) <= not a or b;
    layer7_outputs(5106) <= b;
    layer7_outputs(5107) <= a and b;
    layer7_outputs(5108) <= a;
    layer7_outputs(5109) <= not a;
    layer7_outputs(5110) <= b and not a;
    layer7_outputs(5111) <= b;
    layer7_outputs(5112) <= '0';
    layer7_outputs(5113) <= not (a xor b);
    layer7_outputs(5114) <= a xor b;
    layer7_outputs(5115) <= not b;
    layer7_outputs(5116) <= not a;
    layer7_outputs(5117) <= a and not b;
    layer7_outputs(5118) <= not a;
    layer7_outputs(5119) <= not (a or b);
    layer7_outputs(5120) <= '1';
    layer7_outputs(5121) <= not a;
    layer7_outputs(5122) <= not (a xor b);
    layer7_outputs(5123) <= a or b;
    layer7_outputs(5124) <= not b;
    layer7_outputs(5125) <= not (a or b);
    layer7_outputs(5126) <= a;
    layer7_outputs(5127) <= not (a or b);
    layer7_outputs(5128) <= b and not a;
    layer7_outputs(5129) <= a and b;
    layer7_outputs(5130) <= a and b;
    layer7_outputs(5131) <= a;
    layer7_outputs(5132) <= not b or a;
    layer7_outputs(5133) <= not b;
    layer7_outputs(5134) <= not b;
    layer7_outputs(5135) <= a and b;
    layer7_outputs(5136) <= a;
    layer7_outputs(5137) <= a;
    layer7_outputs(5138) <= a or b;
    layer7_outputs(5139) <= a xor b;
    layer7_outputs(5140) <= a;
    layer7_outputs(5141) <= b;
    layer7_outputs(5142) <= not b or a;
    layer7_outputs(5143) <= a xor b;
    layer7_outputs(5144) <= not a;
    layer7_outputs(5145) <= b;
    layer7_outputs(5146) <= not b;
    layer7_outputs(5147) <= not b;
    layer7_outputs(5148) <= not b;
    layer7_outputs(5149) <= not b;
    layer7_outputs(5150) <= b and not a;
    layer7_outputs(5151) <= b;
    layer7_outputs(5152) <= not a;
    layer7_outputs(5153) <= '0';
    layer7_outputs(5154) <= not (a or b);
    layer7_outputs(5155) <= not (a xor b);
    layer7_outputs(5156) <= b;
    layer7_outputs(5157) <= a and not b;
    layer7_outputs(5158) <= not a;
    layer7_outputs(5159) <= a and not b;
    layer7_outputs(5160) <= b;
    layer7_outputs(5161) <= not (a and b);
    layer7_outputs(5162) <= a and b;
    layer7_outputs(5163) <= not (a and b);
    layer7_outputs(5164) <= a or b;
    layer7_outputs(5165) <= '0';
    layer7_outputs(5166) <= b and not a;
    layer7_outputs(5167) <= not (a xor b);
    layer7_outputs(5168) <= a;
    layer7_outputs(5169) <= not (a xor b);
    layer7_outputs(5170) <= a xor b;
    layer7_outputs(5171) <= a;
    layer7_outputs(5172) <= not b;
    layer7_outputs(5173) <= not a or b;
    layer7_outputs(5174) <= '0';
    layer7_outputs(5175) <= not b;
    layer7_outputs(5176) <= a;
    layer7_outputs(5177) <= a and not b;
    layer7_outputs(5178) <= a or b;
    layer7_outputs(5179) <= not b;
    layer7_outputs(5180) <= b;
    layer7_outputs(5181) <= a;
    layer7_outputs(5182) <= a xor b;
    layer7_outputs(5183) <= not (a and b);
    layer7_outputs(5184) <= not a;
    layer7_outputs(5185) <= a and b;
    layer7_outputs(5186) <= b and not a;
    layer7_outputs(5187) <= '1';
    layer7_outputs(5188) <= not b;
    layer7_outputs(5189) <= a and b;
    layer7_outputs(5190) <= not (a and b);
    layer7_outputs(5191) <= not a;
    layer7_outputs(5192) <= not (a or b);
    layer7_outputs(5193) <= not b;
    layer7_outputs(5194) <= a xor b;
    layer7_outputs(5195) <= b;
    layer7_outputs(5196) <= a;
    layer7_outputs(5197) <= not a;
    layer7_outputs(5198) <= '0';
    layer7_outputs(5199) <= b and not a;
    layer7_outputs(5200) <= a xor b;
    layer7_outputs(5201) <= b;
    layer7_outputs(5202) <= not (a and b);
    layer7_outputs(5203) <= a;
    layer7_outputs(5204) <= a xor b;
    layer7_outputs(5205) <= not (a or b);
    layer7_outputs(5206) <= not a;
    layer7_outputs(5207) <= a and not b;
    layer7_outputs(5208) <= a xor b;
    layer7_outputs(5209) <= not b;
    layer7_outputs(5210) <= a and not b;
    layer7_outputs(5211) <= a or b;
    layer7_outputs(5212) <= not a;
    layer7_outputs(5213) <= not b;
    layer7_outputs(5214) <= a xor b;
    layer7_outputs(5215) <= a or b;
    layer7_outputs(5216) <= '1';
    layer7_outputs(5217) <= a;
    layer7_outputs(5218) <= '0';
    layer7_outputs(5219) <= b;
    layer7_outputs(5220) <= not (a and b);
    layer7_outputs(5221) <= b and not a;
    layer7_outputs(5222) <= not (a and b);
    layer7_outputs(5223) <= b and not a;
    layer7_outputs(5224) <= not b;
    layer7_outputs(5225) <= not b or a;
    layer7_outputs(5226) <= not b;
    layer7_outputs(5227) <= not (a and b);
    layer7_outputs(5228) <= a and not b;
    layer7_outputs(5229) <= not a or b;
    layer7_outputs(5230) <= not a or b;
    layer7_outputs(5231) <= not (a or b);
    layer7_outputs(5232) <= b and not a;
    layer7_outputs(5233) <= a xor b;
    layer7_outputs(5234) <= not (a xor b);
    layer7_outputs(5235) <= not b;
    layer7_outputs(5236) <= not (a or b);
    layer7_outputs(5237) <= a;
    layer7_outputs(5238) <= not a;
    layer7_outputs(5239) <= b;
    layer7_outputs(5240) <= b;
    layer7_outputs(5241) <= not b;
    layer7_outputs(5242) <= not (a and b);
    layer7_outputs(5243) <= not b;
    layer7_outputs(5244) <= b;
    layer7_outputs(5245) <= a;
    layer7_outputs(5246) <= b;
    layer7_outputs(5247) <= not a;
    layer7_outputs(5248) <= not a;
    layer7_outputs(5249) <= b;
    layer7_outputs(5250) <= not (a xor b);
    layer7_outputs(5251) <= not a;
    layer7_outputs(5252) <= a and b;
    layer7_outputs(5253) <= not b;
    layer7_outputs(5254) <= not a;
    layer7_outputs(5255) <= not a or b;
    layer7_outputs(5256) <= not (a or b);
    layer7_outputs(5257) <= b and not a;
    layer7_outputs(5258) <= a and not b;
    layer7_outputs(5259) <= not a;
    layer7_outputs(5260) <= a or b;
    layer7_outputs(5261) <= not (a and b);
    layer7_outputs(5262) <= not (a xor b);
    layer7_outputs(5263) <= b;
    layer7_outputs(5264) <= a;
    layer7_outputs(5265) <= not (a xor b);
    layer7_outputs(5266) <= b;
    layer7_outputs(5267) <= a and b;
    layer7_outputs(5268) <= a xor b;
    layer7_outputs(5269) <= not (a xor b);
    layer7_outputs(5270) <= b;
    layer7_outputs(5271) <= not a;
    layer7_outputs(5272) <= not (a or b);
    layer7_outputs(5273) <= not b;
    layer7_outputs(5274) <= a;
    layer7_outputs(5275) <= b;
    layer7_outputs(5276) <= a xor b;
    layer7_outputs(5277) <= a and b;
    layer7_outputs(5278) <= not b or a;
    layer7_outputs(5279) <= not a;
    layer7_outputs(5280) <= not a;
    layer7_outputs(5281) <= not (a and b);
    layer7_outputs(5282) <= a;
    layer7_outputs(5283) <= a;
    layer7_outputs(5284) <= not (a or b);
    layer7_outputs(5285) <= b and not a;
    layer7_outputs(5286) <= b;
    layer7_outputs(5287) <= a or b;
    layer7_outputs(5288) <= a xor b;
    layer7_outputs(5289) <= a xor b;
    layer7_outputs(5290) <= not a;
    layer7_outputs(5291) <= not a;
    layer7_outputs(5292) <= not (a xor b);
    layer7_outputs(5293) <= not (a or b);
    layer7_outputs(5294) <= a;
    layer7_outputs(5295) <= a;
    layer7_outputs(5296) <= a;
    layer7_outputs(5297) <= not b or a;
    layer7_outputs(5298) <= a and not b;
    layer7_outputs(5299) <= b;
    layer7_outputs(5300) <= b;
    layer7_outputs(5301) <= b;
    layer7_outputs(5302) <= a xor b;
    layer7_outputs(5303) <= b and not a;
    layer7_outputs(5304) <= a;
    layer7_outputs(5305) <= not (a and b);
    layer7_outputs(5306) <= '0';
    layer7_outputs(5307) <= not (a or b);
    layer7_outputs(5308) <= a and b;
    layer7_outputs(5309) <= not (a xor b);
    layer7_outputs(5310) <= b and not a;
    layer7_outputs(5311) <= not (a xor b);
    layer7_outputs(5312) <= not (a or b);
    layer7_outputs(5313) <= not b;
    layer7_outputs(5314) <= a;
    layer7_outputs(5315) <= not b;
    layer7_outputs(5316) <= a or b;
    layer7_outputs(5317) <= a;
    layer7_outputs(5318) <= b and not a;
    layer7_outputs(5319) <= not b or a;
    layer7_outputs(5320) <= a;
    layer7_outputs(5321) <= a;
    layer7_outputs(5322) <= not (a or b);
    layer7_outputs(5323) <= not a;
    layer7_outputs(5324) <= '1';
    layer7_outputs(5325) <= a xor b;
    layer7_outputs(5326) <= not (a and b);
    layer7_outputs(5327) <= '1';
    layer7_outputs(5328) <= not (a or b);
    layer7_outputs(5329) <= not b;
    layer7_outputs(5330) <= a or b;
    layer7_outputs(5331) <= a;
    layer7_outputs(5332) <= not b;
    layer7_outputs(5333) <= not b;
    layer7_outputs(5334) <= not a or b;
    layer7_outputs(5335) <= b and not a;
    layer7_outputs(5336) <= a and not b;
    layer7_outputs(5337) <= a and not b;
    layer7_outputs(5338) <= a and b;
    layer7_outputs(5339) <= not a;
    layer7_outputs(5340) <= not b or a;
    layer7_outputs(5341) <= b;
    layer7_outputs(5342) <= not b;
    layer7_outputs(5343) <= not b;
    layer7_outputs(5344) <= not (a and b);
    layer7_outputs(5345) <= not b;
    layer7_outputs(5346) <= not a;
    layer7_outputs(5347) <= b;
    layer7_outputs(5348) <= b;
    layer7_outputs(5349) <= not b;
    layer7_outputs(5350) <= not b or a;
    layer7_outputs(5351) <= not (a or b);
    layer7_outputs(5352) <= not a or b;
    layer7_outputs(5353) <= a or b;
    layer7_outputs(5354) <= not (a xor b);
    layer7_outputs(5355) <= a and not b;
    layer7_outputs(5356) <= b;
    layer7_outputs(5357) <= not (a or b);
    layer7_outputs(5358) <= a and not b;
    layer7_outputs(5359) <= not b;
    layer7_outputs(5360) <= not (a and b);
    layer7_outputs(5361) <= not (a and b);
    layer7_outputs(5362) <= not a or b;
    layer7_outputs(5363) <= a;
    layer7_outputs(5364) <= not a or b;
    layer7_outputs(5365) <= not b;
    layer7_outputs(5366) <= b and not a;
    layer7_outputs(5367) <= b;
    layer7_outputs(5368) <= a;
    layer7_outputs(5369) <= a and b;
    layer7_outputs(5370) <= '1';
    layer7_outputs(5371) <= b;
    layer7_outputs(5372) <= not a;
    layer7_outputs(5373) <= a and b;
    layer7_outputs(5374) <= not (a xor b);
    layer7_outputs(5375) <= not (a or b);
    layer7_outputs(5376) <= a or b;
    layer7_outputs(5377) <= not (a and b);
    layer7_outputs(5378) <= a or b;
    layer7_outputs(5379) <= b;
    layer7_outputs(5380) <= not a;
    layer7_outputs(5381) <= not b;
    layer7_outputs(5382) <= a and b;
    layer7_outputs(5383) <= not (a xor b);
    layer7_outputs(5384) <= b;
    layer7_outputs(5385) <= '1';
    layer7_outputs(5386) <= not (a and b);
    layer7_outputs(5387) <= not b;
    layer7_outputs(5388) <= a;
    layer7_outputs(5389) <= not (a xor b);
    layer7_outputs(5390) <= a xor b;
    layer7_outputs(5391) <= a;
    layer7_outputs(5392) <= not (a xor b);
    layer7_outputs(5393) <= a and not b;
    layer7_outputs(5394) <= not (a xor b);
    layer7_outputs(5395) <= not b or a;
    layer7_outputs(5396) <= not (a xor b);
    layer7_outputs(5397) <= b;
    layer7_outputs(5398) <= b;
    layer7_outputs(5399) <= a;
    layer7_outputs(5400) <= not a or b;
    layer7_outputs(5401) <= not b;
    layer7_outputs(5402) <= a;
    layer7_outputs(5403) <= not b;
    layer7_outputs(5404) <= not a;
    layer7_outputs(5405) <= a xor b;
    layer7_outputs(5406) <= not b;
    layer7_outputs(5407) <= a;
    layer7_outputs(5408) <= not (a or b);
    layer7_outputs(5409) <= b;
    layer7_outputs(5410) <= not b;
    layer7_outputs(5411) <= a and not b;
    layer7_outputs(5412) <= not a;
    layer7_outputs(5413) <= b;
    layer7_outputs(5414) <= not b;
    layer7_outputs(5415) <= b;
    layer7_outputs(5416) <= a or b;
    layer7_outputs(5417) <= not a;
    layer7_outputs(5418) <= not (a and b);
    layer7_outputs(5419) <= not b;
    layer7_outputs(5420) <= b and not a;
    layer7_outputs(5421) <= not b or a;
    layer7_outputs(5422) <= a xor b;
    layer7_outputs(5423) <= not (a xor b);
    layer7_outputs(5424) <= a xor b;
    layer7_outputs(5425) <= a and not b;
    layer7_outputs(5426) <= not a;
    layer7_outputs(5427) <= not a or b;
    layer7_outputs(5428) <= not (a and b);
    layer7_outputs(5429) <= a and b;
    layer7_outputs(5430) <= not b;
    layer7_outputs(5431) <= not b;
    layer7_outputs(5432) <= a and b;
    layer7_outputs(5433) <= a or b;
    layer7_outputs(5434) <= not (a or b);
    layer7_outputs(5435) <= not b or a;
    layer7_outputs(5436) <= not b;
    layer7_outputs(5437) <= not (a and b);
    layer7_outputs(5438) <= not (a xor b);
    layer7_outputs(5439) <= b and not a;
    layer7_outputs(5440) <= a or b;
    layer7_outputs(5441) <= not (a and b);
    layer7_outputs(5442) <= b and not a;
    layer7_outputs(5443) <= not a or b;
    layer7_outputs(5444) <= a and b;
    layer7_outputs(5445) <= a and b;
    layer7_outputs(5446) <= not (a and b);
    layer7_outputs(5447) <= b;
    layer7_outputs(5448) <= not b or a;
    layer7_outputs(5449) <= '1';
    layer7_outputs(5450) <= not (a and b);
    layer7_outputs(5451) <= not a;
    layer7_outputs(5452) <= b;
    layer7_outputs(5453) <= not b;
    layer7_outputs(5454) <= '0';
    layer7_outputs(5455) <= a;
    layer7_outputs(5456) <= b;
    layer7_outputs(5457) <= a or b;
    layer7_outputs(5458) <= a and not b;
    layer7_outputs(5459) <= b;
    layer7_outputs(5460) <= a and not b;
    layer7_outputs(5461) <= not b;
    layer7_outputs(5462) <= not a;
    layer7_outputs(5463) <= '0';
    layer7_outputs(5464) <= not (a or b);
    layer7_outputs(5465) <= not b;
    layer7_outputs(5466) <= a;
    layer7_outputs(5467) <= b;
    layer7_outputs(5468) <= a or b;
    layer7_outputs(5469) <= not (a xor b);
    layer7_outputs(5470) <= not b;
    layer7_outputs(5471) <= not a;
    layer7_outputs(5472) <= not a or b;
    layer7_outputs(5473) <= not b;
    layer7_outputs(5474) <= a or b;
    layer7_outputs(5475) <= not (a or b);
    layer7_outputs(5476) <= b and not a;
    layer7_outputs(5477) <= b;
    layer7_outputs(5478) <= b;
    layer7_outputs(5479) <= not b;
    layer7_outputs(5480) <= not a or b;
    layer7_outputs(5481) <= not b or a;
    layer7_outputs(5482) <= not (a or b);
    layer7_outputs(5483) <= b;
    layer7_outputs(5484) <= b;
    layer7_outputs(5485) <= not (a or b);
    layer7_outputs(5486) <= not b;
    layer7_outputs(5487) <= not b;
    layer7_outputs(5488) <= a xor b;
    layer7_outputs(5489) <= a and not b;
    layer7_outputs(5490) <= not (a or b);
    layer7_outputs(5491) <= a;
    layer7_outputs(5492) <= a and not b;
    layer7_outputs(5493) <= a or b;
    layer7_outputs(5494) <= '1';
    layer7_outputs(5495) <= not b;
    layer7_outputs(5496) <= not b;
    layer7_outputs(5497) <= not b or a;
    layer7_outputs(5498) <= a or b;
    layer7_outputs(5499) <= not b;
    layer7_outputs(5500) <= a xor b;
    layer7_outputs(5501) <= a xor b;
    layer7_outputs(5502) <= a;
    layer7_outputs(5503) <= a and b;
    layer7_outputs(5504) <= not b;
    layer7_outputs(5505) <= b;
    layer7_outputs(5506) <= b;
    layer7_outputs(5507) <= not (a xor b);
    layer7_outputs(5508) <= not (a xor b);
    layer7_outputs(5509) <= not b;
    layer7_outputs(5510) <= not a;
    layer7_outputs(5511) <= a and not b;
    layer7_outputs(5512) <= a;
    layer7_outputs(5513) <= '1';
    layer7_outputs(5514) <= '0';
    layer7_outputs(5515) <= b and not a;
    layer7_outputs(5516) <= not b;
    layer7_outputs(5517) <= not b;
    layer7_outputs(5518) <= not (a xor b);
    layer7_outputs(5519) <= a or b;
    layer7_outputs(5520) <= not b or a;
    layer7_outputs(5521) <= a and b;
    layer7_outputs(5522) <= a or b;
    layer7_outputs(5523) <= a;
    layer7_outputs(5524) <= not b;
    layer7_outputs(5525) <= not (a xor b);
    layer7_outputs(5526) <= a xor b;
    layer7_outputs(5527) <= not a or b;
    layer7_outputs(5528) <= not b;
    layer7_outputs(5529) <= not (a and b);
    layer7_outputs(5530) <= not b;
    layer7_outputs(5531) <= a;
    layer7_outputs(5532) <= a and not b;
    layer7_outputs(5533) <= a or b;
    layer7_outputs(5534) <= a and b;
    layer7_outputs(5535) <= a or b;
    layer7_outputs(5536) <= not a;
    layer7_outputs(5537) <= b;
    layer7_outputs(5538) <= not b;
    layer7_outputs(5539) <= not a;
    layer7_outputs(5540) <= b;
    layer7_outputs(5541) <= not b or a;
    layer7_outputs(5542) <= not (a xor b);
    layer7_outputs(5543) <= a or b;
    layer7_outputs(5544) <= b and not a;
    layer7_outputs(5545) <= a and not b;
    layer7_outputs(5546) <= b;
    layer7_outputs(5547) <= a and b;
    layer7_outputs(5548) <= b and not a;
    layer7_outputs(5549) <= b and not a;
    layer7_outputs(5550) <= b;
    layer7_outputs(5551) <= b and not a;
    layer7_outputs(5552) <= b;
    layer7_outputs(5553) <= not (a or b);
    layer7_outputs(5554) <= a;
    layer7_outputs(5555) <= not b;
    layer7_outputs(5556) <= a;
    layer7_outputs(5557) <= a;
    layer7_outputs(5558) <= a and b;
    layer7_outputs(5559) <= '0';
    layer7_outputs(5560) <= not b or a;
    layer7_outputs(5561) <= not a;
    layer7_outputs(5562) <= not b or a;
    layer7_outputs(5563) <= not a or b;
    layer7_outputs(5564) <= b;
    layer7_outputs(5565) <= a;
    layer7_outputs(5566) <= not a;
    layer7_outputs(5567) <= a;
    layer7_outputs(5568) <= not (a xor b);
    layer7_outputs(5569) <= not (a or b);
    layer7_outputs(5570) <= a;
    layer7_outputs(5571) <= b;
    layer7_outputs(5572) <= not (a or b);
    layer7_outputs(5573) <= b and not a;
    layer7_outputs(5574) <= not b;
    layer7_outputs(5575) <= a and b;
    layer7_outputs(5576) <= not (a and b);
    layer7_outputs(5577) <= a and not b;
    layer7_outputs(5578) <= a xor b;
    layer7_outputs(5579) <= a xor b;
    layer7_outputs(5580) <= not b;
    layer7_outputs(5581) <= not a;
    layer7_outputs(5582) <= a xor b;
    layer7_outputs(5583) <= a xor b;
    layer7_outputs(5584) <= not (a xor b);
    layer7_outputs(5585) <= '1';
    layer7_outputs(5586) <= not (a or b);
    layer7_outputs(5587) <= not b;
    layer7_outputs(5588) <= not (a and b);
    layer7_outputs(5589) <= a;
    layer7_outputs(5590) <= a;
    layer7_outputs(5591) <= not b;
    layer7_outputs(5592) <= a;
    layer7_outputs(5593) <= not b or a;
    layer7_outputs(5594) <= not (a xor b);
    layer7_outputs(5595) <= not a;
    layer7_outputs(5596) <= not (a and b);
    layer7_outputs(5597) <= not a or b;
    layer7_outputs(5598) <= a and b;
    layer7_outputs(5599) <= b;
    layer7_outputs(5600) <= '0';
    layer7_outputs(5601) <= a xor b;
    layer7_outputs(5602) <= a;
    layer7_outputs(5603) <= '0';
    layer7_outputs(5604) <= not a;
    layer7_outputs(5605) <= not b or a;
    layer7_outputs(5606) <= b;
    layer7_outputs(5607) <= '1';
    layer7_outputs(5608) <= a;
    layer7_outputs(5609) <= not (a and b);
    layer7_outputs(5610) <= a or b;
    layer7_outputs(5611) <= a or b;
    layer7_outputs(5612) <= a;
    layer7_outputs(5613) <= a;
    layer7_outputs(5614) <= not (a and b);
    layer7_outputs(5615) <= not (a or b);
    layer7_outputs(5616) <= b;
    layer7_outputs(5617) <= a;
    layer7_outputs(5618) <= b and not a;
    layer7_outputs(5619) <= b;
    layer7_outputs(5620) <= not a;
    layer7_outputs(5621) <= not b;
    layer7_outputs(5622) <= not b;
    layer7_outputs(5623) <= b;
    layer7_outputs(5624) <= a;
    layer7_outputs(5625) <= '0';
    layer7_outputs(5626) <= not b or a;
    layer7_outputs(5627) <= not (a or b);
    layer7_outputs(5628) <= not b;
    layer7_outputs(5629) <= a or b;
    layer7_outputs(5630) <= not a or b;
    layer7_outputs(5631) <= not a;
    layer7_outputs(5632) <= not (a or b);
    layer7_outputs(5633) <= not (a xor b);
    layer7_outputs(5634) <= a or b;
    layer7_outputs(5635) <= not a;
    layer7_outputs(5636) <= not b or a;
    layer7_outputs(5637) <= not b;
    layer7_outputs(5638) <= a and not b;
    layer7_outputs(5639) <= a and not b;
    layer7_outputs(5640) <= a xor b;
    layer7_outputs(5641) <= a;
    layer7_outputs(5642) <= not b;
    layer7_outputs(5643) <= b;
    layer7_outputs(5644) <= not b or a;
    layer7_outputs(5645) <= a and not b;
    layer7_outputs(5646) <= not (a or b);
    layer7_outputs(5647) <= not a;
    layer7_outputs(5648) <= b;
    layer7_outputs(5649) <= a and not b;
    layer7_outputs(5650) <= not b;
    layer7_outputs(5651) <= a and not b;
    layer7_outputs(5652) <= not a or b;
    layer7_outputs(5653) <= a xor b;
    layer7_outputs(5654) <= a or b;
    layer7_outputs(5655) <= not b;
    layer7_outputs(5656) <= b and not a;
    layer7_outputs(5657) <= a;
    layer7_outputs(5658) <= not a;
    layer7_outputs(5659) <= a;
    layer7_outputs(5660) <= not (a xor b);
    layer7_outputs(5661) <= b;
    layer7_outputs(5662) <= a;
    layer7_outputs(5663) <= not (a or b);
    layer7_outputs(5664) <= not a or b;
    layer7_outputs(5665) <= '0';
    layer7_outputs(5666) <= a or b;
    layer7_outputs(5667) <= not a;
    layer7_outputs(5668) <= not a;
    layer7_outputs(5669) <= not b;
    layer7_outputs(5670) <= not (a xor b);
    layer7_outputs(5671) <= a and b;
    layer7_outputs(5672) <= not b;
    layer7_outputs(5673) <= not a;
    layer7_outputs(5674) <= b;
    layer7_outputs(5675) <= not (a or b);
    layer7_outputs(5676) <= not b;
    layer7_outputs(5677) <= not a;
    layer7_outputs(5678) <= a xor b;
    layer7_outputs(5679) <= not (a or b);
    layer7_outputs(5680) <= not a;
    layer7_outputs(5681) <= a and not b;
    layer7_outputs(5682) <= a xor b;
    layer7_outputs(5683) <= not (a and b);
    layer7_outputs(5684) <= not b;
    layer7_outputs(5685) <= b and not a;
    layer7_outputs(5686) <= a and b;
    layer7_outputs(5687) <= not (a xor b);
    layer7_outputs(5688) <= not (a xor b);
    layer7_outputs(5689) <= a;
    layer7_outputs(5690) <= a xor b;
    layer7_outputs(5691) <= not (a or b);
    layer7_outputs(5692) <= not a;
    layer7_outputs(5693) <= b and not a;
    layer7_outputs(5694) <= b;
    layer7_outputs(5695) <= not (a xor b);
    layer7_outputs(5696) <= not b;
    layer7_outputs(5697) <= not (a xor b);
    layer7_outputs(5698) <= '1';
    layer7_outputs(5699) <= b and not a;
    layer7_outputs(5700) <= b;
    layer7_outputs(5701) <= b and not a;
    layer7_outputs(5702) <= not (a and b);
    layer7_outputs(5703) <= not b;
    layer7_outputs(5704) <= not b or a;
    layer7_outputs(5705) <= not a or b;
    layer7_outputs(5706) <= a xor b;
    layer7_outputs(5707) <= b;
    layer7_outputs(5708) <= not b;
    layer7_outputs(5709) <= b and not a;
    layer7_outputs(5710) <= b;
    layer7_outputs(5711) <= b;
    layer7_outputs(5712) <= not a;
    layer7_outputs(5713) <= not b;
    layer7_outputs(5714) <= not a or b;
    layer7_outputs(5715) <= a or b;
    layer7_outputs(5716) <= a and not b;
    layer7_outputs(5717) <= not (a xor b);
    layer7_outputs(5718) <= not a;
    layer7_outputs(5719) <= not (a or b);
    layer7_outputs(5720) <= not b or a;
    layer7_outputs(5721) <= not (a or b);
    layer7_outputs(5722) <= a and not b;
    layer7_outputs(5723) <= a and b;
    layer7_outputs(5724) <= not a;
    layer7_outputs(5725) <= a;
    layer7_outputs(5726) <= not (a or b);
    layer7_outputs(5727) <= not b;
    layer7_outputs(5728) <= not a or b;
    layer7_outputs(5729) <= not a;
    layer7_outputs(5730) <= a or b;
    layer7_outputs(5731) <= not b or a;
    layer7_outputs(5732) <= a and b;
    layer7_outputs(5733) <= not (a or b);
    layer7_outputs(5734) <= b;
    layer7_outputs(5735) <= not a;
    layer7_outputs(5736) <= a and not b;
    layer7_outputs(5737) <= b and not a;
    layer7_outputs(5738) <= b;
    layer7_outputs(5739) <= not (a xor b);
    layer7_outputs(5740) <= '0';
    layer7_outputs(5741) <= not a;
    layer7_outputs(5742) <= a;
    layer7_outputs(5743) <= not (a and b);
    layer7_outputs(5744) <= not (a xor b);
    layer7_outputs(5745) <= a and b;
    layer7_outputs(5746) <= a and b;
    layer7_outputs(5747) <= not b;
    layer7_outputs(5748) <= not a;
    layer7_outputs(5749) <= a and not b;
    layer7_outputs(5750) <= not a or b;
    layer7_outputs(5751) <= not b;
    layer7_outputs(5752) <= b;
    layer7_outputs(5753) <= '1';
    layer7_outputs(5754) <= not b or a;
    layer7_outputs(5755) <= a or b;
    layer7_outputs(5756) <= not (a and b);
    layer7_outputs(5757) <= a and not b;
    layer7_outputs(5758) <= b;
    layer7_outputs(5759) <= b and not a;
    layer7_outputs(5760) <= a and not b;
    layer7_outputs(5761) <= b;
    layer7_outputs(5762) <= '1';
    layer7_outputs(5763) <= a and not b;
    layer7_outputs(5764) <= not (a xor b);
    layer7_outputs(5765) <= a;
    layer7_outputs(5766) <= a;
    layer7_outputs(5767) <= not b;
    layer7_outputs(5768) <= not (a or b);
    layer7_outputs(5769) <= not a or b;
    layer7_outputs(5770) <= b;
    layer7_outputs(5771) <= not (a or b);
    layer7_outputs(5772) <= not b or a;
    layer7_outputs(5773) <= a xor b;
    layer7_outputs(5774) <= b;
    layer7_outputs(5775) <= not (a xor b);
    layer7_outputs(5776) <= b;
    layer7_outputs(5777) <= a xor b;
    layer7_outputs(5778) <= b;
    layer7_outputs(5779) <= a and not b;
    layer7_outputs(5780) <= a;
    layer7_outputs(5781) <= b;
    layer7_outputs(5782) <= a or b;
    layer7_outputs(5783) <= a;
    layer7_outputs(5784) <= not (a or b);
    layer7_outputs(5785) <= b;
    layer7_outputs(5786) <= not b;
    layer7_outputs(5787) <= not a;
    layer7_outputs(5788) <= not (a xor b);
    layer7_outputs(5789) <= a xor b;
    layer7_outputs(5790) <= not b;
    layer7_outputs(5791) <= not b;
    layer7_outputs(5792) <= not b or a;
    layer7_outputs(5793) <= a and not b;
    layer7_outputs(5794) <= not (a and b);
    layer7_outputs(5795) <= a;
    layer7_outputs(5796) <= not b;
    layer7_outputs(5797) <= b and not a;
    layer7_outputs(5798) <= not b;
    layer7_outputs(5799) <= not b;
    layer7_outputs(5800) <= a xor b;
    layer7_outputs(5801) <= a and b;
    layer7_outputs(5802) <= not (a xor b);
    layer7_outputs(5803) <= not (a and b);
    layer7_outputs(5804) <= a xor b;
    layer7_outputs(5805) <= a and b;
    layer7_outputs(5806) <= not (a or b);
    layer7_outputs(5807) <= not a;
    layer7_outputs(5808) <= not (a and b);
    layer7_outputs(5809) <= not a;
    layer7_outputs(5810) <= not b;
    layer7_outputs(5811) <= not (a and b);
    layer7_outputs(5812) <= a xor b;
    layer7_outputs(5813) <= b;
    layer7_outputs(5814) <= b;
    layer7_outputs(5815) <= a xor b;
    layer7_outputs(5816) <= a and b;
    layer7_outputs(5817) <= not (a and b);
    layer7_outputs(5818) <= a xor b;
    layer7_outputs(5819) <= not a or b;
    layer7_outputs(5820) <= not (a or b);
    layer7_outputs(5821) <= not b or a;
    layer7_outputs(5822) <= a;
    layer7_outputs(5823) <= b;
    layer7_outputs(5824) <= not b;
    layer7_outputs(5825) <= a;
    layer7_outputs(5826) <= not a;
    layer7_outputs(5827) <= not (a and b);
    layer7_outputs(5828) <= not a or b;
    layer7_outputs(5829) <= not a;
    layer7_outputs(5830) <= a and b;
    layer7_outputs(5831) <= not (a or b);
    layer7_outputs(5832) <= a or b;
    layer7_outputs(5833) <= b;
    layer7_outputs(5834) <= not (a and b);
    layer7_outputs(5835) <= not (a xor b);
    layer7_outputs(5836) <= a and b;
    layer7_outputs(5837) <= a and b;
    layer7_outputs(5838) <= a xor b;
    layer7_outputs(5839) <= not (a and b);
    layer7_outputs(5840) <= a;
    layer7_outputs(5841) <= a or b;
    layer7_outputs(5842) <= not (a and b);
    layer7_outputs(5843) <= not a;
    layer7_outputs(5844) <= a and b;
    layer7_outputs(5845) <= not (a xor b);
    layer7_outputs(5846) <= a;
    layer7_outputs(5847) <= not b;
    layer7_outputs(5848) <= b;
    layer7_outputs(5849) <= not b or a;
    layer7_outputs(5850) <= not (a or b);
    layer7_outputs(5851) <= not (a and b);
    layer7_outputs(5852) <= a;
    layer7_outputs(5853) <= a and b;
    layer7_outputs(5854) <= not (a or b);
    layer7_outputs(5855) <= a xor b;
    layer7_outputs(5856) <= not a;
    layer7_outputs(5857) <= not (a xor b);
    layer7_outputs(5858) <= a;
    layer7_outputs(5859) <= not (a or b);
    layer7_outputs(5860) <= not b;
    layer7_outputs(5861) <= a and not b;
    layer7_outputs(5862) <= a xor b;
    layer7_outputs(5863) <= a or b;
    layer7_outputs(5864) <= b;
    layer7_outputs(5865) <= a;
    layer7_outputs(5866) <= not (a and b);
    layer7_outputs(5867) <= a;
    layer7_outputs(5868) <= not (a xor b);
    layer7_outputs(5869) <= a xor b;
    layer7_outputs(5870) <= a;
    layer7_outputs(5871) <= not (a and b);
    layer7_outputs(5872) <= not (a and b);
    layer7_outputs(5873) <= a and not b;
    layer7_outputs(5874) <= b and not a;
    layer7_outputs(5875) <= not (a or b);
    layer7_outputs(5876) <= a or b;
    layer7_outputs(5877) <= a xor b;
    layer7_outputs(5878) <= a and not b;
    layer7_outputs(5879) <= not a;
    layer7_outputs(5880) <= not a;
    layer7_outputs(5881) <= a;
    layer7_outputs(5882) <= not (a xor b);
    layer7_outputs(5883) <= '0';
    layer7_outputs(5884) <= not (a or b);
    layer7_outputs(5885) <= a;
    layer7_outputs(5886) <= '0';
    layer7_outputs(5887) <= '0';
    layer7_outputs(5888) <= not a;
    layer7_outputs(5889) <= a xor b;
    layer7_outputs(5890) <= not (a xor b);
    layer7_outputs(5891) <= not b;
    layer7_outputs(5892) <= not (a or b);
    layer7_outputs(5893) <= not (a and b);
    layer7_outputs(5894) <= b;
    layer7_outputs(5895) <= a and not b;
    layer7_outputs(5896) <= not (a xor b);
    layer7_outputs(5897) <= not (a or b);
    layer7_outputs(5898) <= not (a and b);
    layer7_outputs(5899) <= b and not a;
    layer7_outputs(5900) <= a;
    layer7_outputs(5901) <= a;
    layer7_outputs(5902) <= '1';
    layer7_outputs(5903) <= b;
    layer7_outputs(5904) <= not b;
    layer7_outputs(5905) <= b;
    layer7_outputs(5906) <= not (a and b);
    layer7_outputs(5907) <= not b;
    layer7_outputs(5908) <= a or b;
    layer7_outputs(5909) <= b;
    layer7_outputs(5910) <= b;
    layer7_outputs(5911) <= a;
    layer7_outputs(5912) <= not (a and b);
    layer7_outputs(5913) <= not (a xor b);
    layer7_outputs(5914) <= a xor b;
    layer7_outputs(5915) <= not a;
    layer7_outputs(5916) <= '1';
    layer7_outputs(5917) <= not a;
    layer7_outputs(5918) <= a;
    layer7_outputs(5919) <= a;
    layer7_outputs(5920) <= not b or a;
    layer7_outputs(5921) <= not (a xor b);
    layer7_outputs(5922) <= a;
    layer7_outputs(5923) <= not (a xor b);
    layer7_outputs(5924) <= a;
    layer7_outputs(5925) <= not a or b;
    layer7_outputs(5926) <= not a;
    layer7_outputs(5927) <= a;
    layer7_outputs(5928) <= not a;
    layer7_outputs(5929) <= not a;
    layer7_outputs(5930) <= a or b;
    layer7_outputs(5931) <= not (a xor b);
    layer7_outputs(5932) <= not a;
    layer7_outputs(5933) <= not a or b;
    layer7_outputs(5934) <= not a or b;
    layer7_outputs(5935) <= not b;
    layer7_outputs(5936) <= not a;
    layer7_outputs(5937) <= not b;
    layer7_outputs(5938) <= a and b;
    layer7_outputs(5939) <= not b or a;
    layer7_outputs(5940) <= not b;
    layer7_outputs(5941) <= not b;
    layer7_outputs(5942) <= a;
    layer7_outputs(5943) <= a;
    layer7_outputs(5944) <= a xor b;
    layer7_outputs(5945) <= b and not a;
    layer7_outputs(5946) <= a;
    layer7_outputs(5947) <= not a;
    layer7_outputs(5948) <= a;
    layer7_outputs(5949) <= a and b;
    layer7_outputs(5950) <= not (a or b);
    layer7_outputs(5951) <= a;
    layer7_outputs(5952) <= a xor b;
    layer7_outputs(5953) <= not a;
    layer7_outputs(5954) <= a;
    layer7_outputs(5955) <= not a;
    layer7_outputs(5956) <= a and not b;
    layer7_outputs(5957) <= not a;
    layer7_outputs(5958) <= not (a xor b);
    layer7_outputs(5959) <= a xor b;
    layer7_outputs(5960) <= b;
    layer7_outputs(5961) <= '1';
    layer7_outputs(5962) <= a;
    layer7_outputs(5963) <= a and not b;
    layer7_outputs(5964) <= not b;
    layer7_outputs(5965) <= a xor b;
    layer7_outputs(5966) <= a;
    layer7_outputs(5967) <= not a or b;
    layer7_outputs(5968) <= not (a xor b);
    layer7_outputs(5969) <= not b;
    layer7_outputs(5970) <= a and not b;
    layer7_outputs(5971) <= not (a and b);
    layer7_outputs(5972) <= not b;
    layer7_outputs(5973) <= not b or a;
    layer7_outputs(5974) <= a and b;
    layer7_outputs(5975) <= b;
    layer7_outputs(5976) <= not (a xor b);
    layer7_outputs(5977) <= not b or a;
    layer7_outputs(5978) <= not b;
    layer7_outputs(5979) <= not (a or b);
    layer7_outputs(5980) <= not a;
    layer7_outputs(5981) <= not (a xor b);
    layer7_outputs(5982) <= a and b;
    layer7_outputs(5983) <= not a;
    layer7_outputs(5984) <= not a;
    layer7_outputs(5985) <= not (a xor b);
    layer7_outputs(5986) <= not (a or b);
    layer7_outputs(5987) <= not b;
    layer7_outputs(5988) <= a;
    layer7_outputs(5989) <= not (a and b);
    layer7_outputs(5990) <= not a;
    layer7_outputs(5991) <= not a or b;
    layer7_outputs(5992) <= not a or b;
    layer7_outputs(5993) <= not b;
    layer7_outputs(5994) <= not b;
    layer7_outputs(5995) <= b;
    layer7_outputs(5996) <= a and not b;
    layer7_outputs(5997) <= not a;
    layer7_outputs(5998) <= a;
    layer7_outputs(5999) <= a or b;
    layer7_outputs(6000) <= not a or b;
    layer7_outputs(6001) <= not (a xor b);
    layer7_outputs(6002) <= not b;
    layer7_outputs(6003) <= a and b;
    layer7_outputs(6004) <= not a;
    layer7_outputs(6005) <= a and b;
    layer7_outputs(6006) <= not (a xor b);
    layer7_outputs(6007) <= b;
    layer7_outputs(6008) <= not a or b;
    layer7_outputs(6009) <= not (a xor b);
    layer7_outputs(6010) <= a;
    layer7_outputs(6011) <= not a;
    layer7_outputs(6012) <= not a or b;
    layer7_outputs(6013) <= not a or b;
    layer7_outputs(6014) <= not a or b;
    layer7_outputs(6015) <= not (a xor b);
    layer7_outputs(6016) <= not b or a;
    layer7_outputs(6017) <= a xor b;
    layer7_outputs(6018) <= a or b;
    layer7_outputs(6019) <= a or b;
    layer7_outputs(6020) <= not a;
    layer7_outputs(6021) <= not b;
    layer7_outputs(6022) <= a or b;
    layer7_outputs(6023) <= not a;
    layer7_outputs(6024) <= a;
    layer7_outputs(6025) <= not a or b;
    layer7_outputs(6026) <= a or b;
    layer7_outputs(6027) <= b;
    layer7_outputs(6028) <= a xor b;
    layer7_outputs(6029) <= a and b;
    layer7_outputs(6030) <= not a;
    layer7_outputs(6031) <= not a;
    layer7_outputs(6032) <= not (a and b);
    layer7_outputs(6033) <= not a or b;
    layer7_outputs(6034) <= b;
    layer7_outputs(6035) <= not a;
    layer7_outputs(6036) <= not a;
    layer7_outputs(6037) <= a or b;
    layer7_outputs(6038) <= a or b;
    layer7_outputs(6039) <= a and not b;
    layer7_outputs(6040) <= not (a and b);
    layer7_outputs(6041) <= not b or a;
    layer7_outputs(6042) <= not (a xor b);
    layer7_outputs(6043) <= b and not a;
    layer7_outputs(6044) <= not b;
    layer7_outputs(6045) <= a xor b;
    layer7_outputs(6046) <= a and not b;
    layer7_outputs(6047) <= not a;
    layer7_outputs(6048) <= not b;
    layer7_outputs(6049) <= a;
    layer7_outputs(6050) <= not b;
    layer7_outputs(6051) <= a;
    layer7_outputs(6052) <= not a;
    layer7_outputs(6053) <= a;
    layer7_outputs(6054) <= a;
    layer7_outputs(6055) <= not a;
    layer7_outputs(6056) <= not (a xor b);
    layer7_outputs(6057) <= b;
    layer7_outputs(6058) <= b and not a;
    layer7_outputs(6059) <= a or b;
    layer7_outputs(6060) <= not a;
    layer7_outputs(6061) <= not a;
    layer7_outputs(6062) <= not b;
    layer7_outputs(6063) <= a or b;
    layer7_outputs(6064) <= a xor b;
    layer7_outputs(6065) <= b;
    layer7_outputs(6066) <= a xor b;
    layer7_outputs(6067) <= not a or b;
    layer7_outputs(6068) <= a and not b;
    layer7_outputs(6069) <= not a;
    layer7_outputs(6070) <= a xor b;
    layer7_outputs(6071) <= not (a xor b);
    layer7_outputs(6072) <= a and b;
    layer7_outputs(6073) <= a;
    layer7_outputs(6074) <= a or b;
    layer7_outputs(6075) <= not b;
    layer7_outputs(6076) <= not (a xor b);
    layer7_outputs(6077) <= b;
    layer7_outputs(6078) <= a and b;
    layer7_outputs(6079) <= b;
    layer7_outputs(6080) <= not (a and b);
    layer7_outputs(6081) <= a;
    layer7_outputs(6082) <= b and not a;
    layer7_outputs(6083) <= not b;
    layer7_outputs(6084) <= not a or b;
    layer7_outputs(6085) <= b;
    layer7_outputs(6086) <= a or b;
    layer7_outputs(6087) <= a xor b;
    layer7_outputs(6088) <= a;
    layer7_outputs(6089) <= a and b;
    layer7_outputs(6090) <= b;
    layer7_outputs(6091) <= not b or a;
    layer7_outputs(6092) <= not (a and b);
    layer7_outputs(6093) <= a xor b;
    layer7_outputs(6094) <= a;
    layer7_outputs(6095) <= not (a and b);
    layer7_outputs(6096) <= not (a and b);
    layer7_outputs(6097) <= not (a xor b);
    layer7_outputs(6098) <= not b or a;
    layer7_outputs(6099) <= not b or a;
    layer7_outputs(6100) <= '1';
    layer7_outputs(6101) <= not a;
    layer7_outputs(6102) <= a and not b;
    layer7_outputs(6103) <= b;
    layer7_outputs(6104) <= not b;
    layer7_outputs(6105) <= b and not a;
    layer7_outputs(6106) <= b and not a;
    layer7_outputs(6107) <= not b;
    layer7_outputs(6108) <= b;
    layer7_outputs(6109) <= b and not a;
    layer7_outputs(6110) <= not a;
    layer7_outputs(6111) <= b;
    layer7_outputs(6112) <= not (a or b);
    layer7_outputs(6113) <= a;
    layer7_outputs(6114) <= b;
    layer7_outputs(6115) <= a;
    layer7_outputs(6116) <= a;
    layer7_outputs(6117) <= a and b;
    layer7_outputs(6118) <= not a;
    layer7_outputs(6119) <= b;
    layer7_outputs(6120) <= b;
    layer7_outputs(6121) <= a or b;
    layer7_outputs(6122) <= not b;
    layer7_outputs(6123) <= not a;
    layer7_outputs(6124) <= not b;
    layer7_outputs(6125) <= a or b;
    layer7_outputs(6126) <= not a;
    layer7_outputs(6127) <= not b;
    layer7_outputs(6128) <= a and b;
    layer7_outputs(6129) <= b;
    layer7_outputs(6130) <= b and not a;
    layer7_outputs(6131) <= not b;
    layer7_outputs(6132) <= not a;
    layer7_outputs(6133) <= b;
    layer7_outputs(6134) <= not b;
    layer7_outputs(6135) <= a and b;
    layer7_outputs(6136) <= a;
    layer7_outputs(6137) <= a xor b;
    layer7_outputs(6138) <= not b or a;
    layer7_outputs(6139) <= a and b;
    layer7_outputs(6140) <= not a;
    layer7_outputs(6141) <= b;
    layer7_outputs(6142) <= not b;
    layer7_outputs(6143) <= not a or b;
    layer7_outputs(6144) <= not a or b;
    layer7_outputs(6145) <= a and not b;
    layer7_outputs(6146) <= a and not b;
    layer7_outputs(6147) <= b;
    layer7_outputs(6148) <= not a;
    layer7_outputs(6149) <= not a or b;
    layer7_outputs(6150) <= a and not b;
    layer7_outputs(6151) <= not a or b;
    layer7_outputs(6152) <= b;
    layer7_outputs(6153) <= a and b;
    layer7_outputs(6154) <= not b or a;
    layer7_outputs(6155) <= not a;
    layer7_outputs(6156) <= not a or b;
    layer7_outputs(6157) <= not (a xor b);
    layer7_outputs(6158) <= a xor b;
    layer7_outputs(6159) <= a or b;
    layer7_outputs(6160) <= a and not b;
    layer7_outputs(6161) <= a xor b;
    layer7_outputs(6162) <= a xor b;
    layer7_outputs(6163) <= not b;
    layer7_outputs(6164) <= '1';
    layer7_outputs(6165) <= not b or a;
    layer7_outputs(6166) <= not b;
    layer7_outputs(6167) <= not (a xor b);
    layer7_outputs(6168) <= not b or a;
    layer7_outputs(6169) <= not (a or b);
    layer7_outputs(6170) <= a;
    layer7_outputs(6171) <= b;
    layer7_outputs(6172) <= not a;
    layer7_outputs(6173) <= not (a xor b);
    layer7_outputs(6174) <= a or b;
    layer7_outputs(6175) <= b;
    layer7_outputs(6176) <= not (a or b);
    layer7_outputs(6177) <= not (a xor b);
    layer7_outputs(6178) <= a xor b;
    layer7_outputs(6179) <= not b;
    layer7_outputs(6180) <= not b or a;
    layer7_outputs(6181) <= a;
    layer7_outputs(6182) <= a and b;
    layer7_outputs(6183) <= not (a and b);
    layer7_outputs(6184) <= not b;
    layer7_outputs(6185) <= a xor b;
    layer7_outputs(6186) <= a;
    layer7_outputs(6187) <= b and not a;
    layer7_outputs(6188) <= a and not b;
    layer7_outputs(6189) <= a;
    layer7_outputs(6190) <= not a;
    layer7_outputs(6191) <= not a;
    layer7_outputs(6192) <= not a;
    layer7_outputs(6193) <= not b or a;
    layer7_outputs(6194) <= a xor b;
    layer7_outputs(6195) <= not (a and b);
    layer7_outputs(6196) <= not (a or b);
    layer7_outputs(6197) <= a or b;
    layer7_outputs(6198) <= not (a and b);
    layer7_outputs(6199) <= a xor b;
    layer7_outputs(6200) <= not a;
    layer7_outputs(6201) <= a;
    layer7_outputs(6202) <= not b or a;
    layer7_outputs(6203) <= not b;
    layer7_outputs(6204) <= a and b;
    layer7_outputs(6205) <= not (a or b);
    layer7_outputs(6206) <= not b;
    layer7_outputs(6207) <= not (a or b);
    layer7_outputs(6208) <= a and b;
    layer7_outputs(6209) <= not a;
    layer7_outputs(6210) <= b and not a;
    layer7_outputs(6211) <= a and b;
    layer7_outputs(6212) <= b;
    layer7_outputs(6213) <= b;
    layer7_outputs(6214) <= a;
    layer7_outputs(6215) <= not a;
    layer7_outputs(6216) <= not (a xor b);
    layer7_outputs(6217) <= b;
    layer7_outputs(6218) <= a or b;
    layer7_outputs(6219) <= a;
    layer7_outputs(6220) <= not (a or b);
    layer7_outputs(6221) <= not b;
    layer7_outputs(6222) <= a and not b;
    layer7_outputs(6223) <= b and not a;
    layer7_outputs(6224) <= a or b;
    layer7_outputs(6225) <= a;
    layer7_outputs(6226) <= b;
    layer7_outputs(6227) <= a and not b;
    layer7_outputs(6228) <= not (a or b);
    layer7_outputs(6229) <= a or b;
    layer7_outputs(6230) <= a or b;
    layer7_outputs(6231) <= b and not a;
    layer7_outputs(6232) <= not a;
    layer7_outputs(6233) <= not a;
    layer7_outputs(6234) <= not a;
    layer7_outputs(6235) <= a;
    layer7_outputs(6236) <= not (a xor b);
    layer7_outputs(6237) <= a and not b;
    layer7_outputs(6238) <= not a;
    layer7_outputs(6239) <= a xor b;
    layer7_outputs(6240) <= not (a xor b);
    layer7_outputs(6241) <= a xor b;
    layer7_outputs(6242) <= a and b;
    layer7_outputs(6243) <= b;
    layer7_outputs(6244) <= b;
    layer7_outputs(6245) <= not (a or b);
    layer7_outputs(6246) <= a xor b;
    layer7_outputs(6247) <= b and not a;
    layer7_outputs(6248) <= a or b;
    layer7_outputs(6249) <= not (a or b);
    layer7_outputs(6250) <= a and not b;
    layer7_outputs(6251) <= not b;
    layer7_outputs(6252) <= b;
    layer7_outputs(6253) <= a;
    layer7_outputs(6254) <= a and b;
    layer7_outputs(6255) <= a xor b;
    layer7_outputs(6256) <= b;
    layer7_outputs(6257) <= '1';
    layer7_outputs(6258) <= a and not b;
    layer7_outputs(6259) <= '1';
    layer7_outputs(6260) <= not a;
    layer7_outputs(6261) <= not a;
    layer7_outputs(6262) <= not b;
    layer7_outputs(6263) <= not b;
    layer7_outputs(6264) <= a xor b;
    layer7_outputs(6265) <= not (a and b);
    layer7_outputs(6266) <= a and not b;
    layer7_outputs(6267) <= a;
    layer7_outputs(6268) <= not b;
    layer7_outputs(6269) <= not (a xor b);
    layer7_outputs(6270) <= a and not b;
    layer7_outputs(6271) <= not b;
    layer7_outputs(6272) <= b;
    layer7_outputs(6273) <= b;
    layer7_outputs(6274) <= not b;
    layer7_outputs(6275) <= b;
    layer7_outputs(6276) <= a or b;
    layer7_outputs(6277) <= a or b;
    layer7_outputs(6278) <= b;
    layer7_outputs(6279) <= not b or a;
    layer7_outputs(6280) <= a xor b;
    layer7_outputs(6281) <= not b;
    layer7_outputs(6282) <= not (a and b);
    layer7_outputs(6283) <= b and not a;
    layer7_outputs(6284) <= a;
    layer7_outputs(6285) <= b and not a;
    layer7_outputs(6286) <= a xor b;
    layer7_outputs(6287) <= not a;
    layer7_outputs(6288) <= not b;
    layer7_outputs(6289) <= a and b;
    layer7_outputs(6290) <= not (a xor b);
    layer7_outputs(6291) <= not b;
    layer7_outputs(6292) <= not a;
    layer7_outputs(6293) <= '1';
    layer7_outputs(6294) <= a;
    layer7_outputs(6295) <= a or b;
    layer7_outputs(6296) <= not a;
    layer7_outputs(6297) <= a and not b;
    layer7_outputs(6298) <= a;
    layer7_outputs(6299) <= a;
    layer7_outputs(6300) <= a and b;
    layer7_outputs(6301) <= not (a or b);
    layer7_outputs(6302) <= a or b;
    layer7_outputs(6303) <= b;
    layer7_outputs(6304) <= a and not b;
    layer7_outputs(6305) <= not a or b;
    layer7_outputs(6306) <= not (a xor b);
    layer7_outputs(6307) <= a and b;
    layer7_outputs(6308) <= not a or b;
    layer7_outputs(6309) <= b;
    layer7_outputs(6310) <= '0';
    layer7_outputs(6311) <= a;
    layer7_outputs(6312) <= b;
    layer7_outputs(6313) <= not (a and b);
    layer7_outputs(6314) <= a xor b;
    layer7_outputs(6315) <= b;
    layer7_outputs(6316) <= b;
    layer7_outputs(6317) <= not (a xor b);
    layer7_outputs(6318) <= not b;
    layer7_outputs(6319) <= not a;
    layer7_outputs(6320) <= a xor b;
    layer7_outputs(6321) <= not a;
    layer7_outputs(6322) <= b and not a;
    layer7_outputs(6323) <= a;
    layer7_outputs(6324) <= a and b;
    layer7_outputs(6325) <= b and not a;
    layer7_outputs(6326) <= not b;
    layer7_outputs(6327) <= a;
    layer7_outputs(6328) <= b;
    layer7_outputs(6329) <= a;
    layer7_outputs(6330) <= a or b;
    layer7_outputs(6331) <= a;
    layer7_outputs(6332) <= not b;
    layer7_outputs(6333) <= not (a xor b);
    layer7_outputs(6334) <= b and not a;
    layer7_outputs(6335) <= a;
    layer7_outputs(6336) <= not a;
    layer7_outputs(6337) <= a xor b;
    layer7_outputs(6338) <= not a;
    layer7_outputs(6339) <= a xor b;
    layer7_outputs(6340) <= not (a and b);
    layer7_outputs(6341) <= b;
    layer7_outputs(6342) <= a;
    layer7_outputs(6343) <= not b;
    layer7_outputs(6344) <= a or b;
    layer7_outputs(6345) <= not b;
    layer7_outputs(6346) <= not (a or b);
    layer7_outputs(6347) <= not a;
    layer7_outputs(6348) <= a and b;
    layer7_outputs(6349) <= not (a or b);
    layer7_outputs(6350) <= not a;
    layer7_outputs(6351) <= not (a and b);
    layer7_outputs(6352) <= b;
    layer7_outputs(6353) <= not (a or b);
    layer7_outputs(6354) <= not a or b;
    layer7_outputs(6355) <= '0';
    layer7_outputs(6356) <= not a;
    layer7_outputs(6357) <= not (a xor b);
    layer7_outputs(6358) <= a xor b;
    layer7_outputs(6359) <= not a;
    layer7_outputs(6360) <= not b;
    layer7_outputs(6361) <= b;
    layer7_outputs(6362) <= a;
    layer7_outputs(6363) <= not (a xor b);
    layer7_outputs(6364) <= not b;
    layer7_outputs(6365) <= not b;
    layer7_outputs(6366) <= not a or b;
    layer7_outputs(6367) <= b;
    layer7_outputs(6368) <= a and not b;
    layer7_outputs(6369) <= not a or b;
    layer7_outputs(6370) <= b;
    layer7_outputs(6371) <= not (a xor b);
    layer7_outputs(6372) <= not b;
    layer7_outputs(6373) <= b;
    layer7_outputs(6374) <= b;
    layer7_outputs(6375) <= a and b;
    layer7_outputs(6376) <= not b;
    layer7_outputs(6377) <= not a;
    layer7_outputs(6378) <= b;
    layer7_outputs(6379) <= not a;
    layer7_outputs(6380) <= not (a xor b);
    layer7_outputs(6381) <= not b;
    layer7_outputs(6382) <= b and not a;
    layer7_outputs(6383) <= a;
    layer7_outputs(6384) <= not b;
    layer7_outputs(6385) <= not b or a;
    layer7_outputs(6386) <= not a;
    layer7_outputs(6387) <= b;
    layer7_outputs(6388) <= a and b;
    layer7_outputs(6389) <= not (a xor b);
    layer7_outputs(6390) <= b;
    layer7_outputs(6391) <= not a;
    layer7_outputs(6392) <= b;
    layer7_outputs(6393) <= not a;
    layer7_outputs(6394) <= a or b;
    layer7_outputs(6395) <= not a;
    layer7_outputs(6396) <= a or b;
    layer7_outputs(6397) <= not b or a;
    layer7_outputs(6398) <= not b;
    layer7_outputs(6399) <= b;
    layer7_outputs(6400) <= b;
    layer7_outputs(6401) <= a;
    layer7_outputs(6402) <= not b;
    layer7_outputs(6403) <= not a or b;
    layer7_outputs(6404) <= not (a and b);
    layer7_outputs(6405) <= not a;
    layer7_outputs(6406) <= a and b;
    layer7_outputs(6407) <= not b or a;
    layer7_outputs(6408) <= a;
    layer7_outputs(6409) <= a;
    layer7_outputs(6410) <= not (a xor b);
    layer7_outputs(6411) <= not a;
    layer7_outputs(6412) <= a;
    layer7_outputs(6413) <= a;
    layer7_outputs(6414) <= not b;
    layer7_outputs(6415) <= '1';
    layer7_outputs(6416) <= a and not b;
    layer7_outputs(6417) <= not b;
    layer7_outputs(6418) <= not (a and b);
    layer7_outputs(6419) <= a xor b;
    layer7_outputs(6420) <= b and not a;
    layer7_outputs(6421) <= not b or a;
    layer7_outputs(6422) <= not (a and b);
    layer7_outputs(6423) <= a;
    layer7_outputs(6424) <= a or b;
    layer7_outputs(6425) <= b;
    layer7_outputs(6426) <= not a or b;
    layer7_outputs(6427) <= not (a xor b);
    layer7_outputs(6428) <= a xor b;
    layer7_outputs(6429) <= a and b;
    layer7_outputs(6430) <= a xor b;
    layer7_outputs(6431) <= not a;
    layer7_outputs(6432) <= a and not b;
    layer7_outputs(6433) <= a xor b;
    layer7_outputs(6434) <= a or b;
    layer7_outputs(6435) <= b;
    layer7_outputs(6436) <= not (a or b);
    layer7_outputs(6437) <= a and not b;
    layer7_outputs(6438) <= not (a and b);
    layer7_outputs(6439) <= '1';
    layer7_outputs(6440) <= b;
    layer7_outputs(6441) <= a or b;
    layer7_outputs(6442) <= not b;
    layer7_outputs(6443) <= not (a and b);
    layer7_outputs(6444) <= a xor b;
    layer7_outputs(6445) <= not b or a;
    layer7_outputs(6446) <= not b;
    layer7_outputs(6447) <= a xor b;
    layer7_outputs(6448) <= not (a or b);
    layer7_outputs(6449) <= not b;
    layer7_outputs(6450) <= not a or b;
    layer7_outputs(6451) <= not b;
    layer7_outputs(6452) <= not (a or b);
    layer7_outputs(6453) <= not b;
    layer7_outputs(6454) <= not b;
    layer7_outputs(6455) <= not a;
    layer7_outputs(6456) <= b;
    layer7_outputs(6457) <= a xor b;
    layer7_outputs(6458) <= a xor b;
    layer7_outputs(6459) <= not a;
    layer7_outputs(6460) <= not b;
    layer7_outputs(6461) <= a and b;
    layer7_outputs(6462) <= b;
    layer7_outputs(6463) <= not (a xor b);
    layer7_outputs(6464) <= not b or a;
    layer7_outputs(6465) <= a;
    layer7_outputs(6466) <= a xor b;
    layer7_outputs(6467) <= b;
    layer7_outputs(6468) <= not a;
    layer7_outputs(6469) <= not (a xor b);
    layer7_outputs(6470) <= not (a or b);
    layer7_outputs(6471) <= b;
    layer7_outputs(6472) <= not a or b;
    layer7_outputs(6473) <= a;
    layer7_outputs(6474) <= not a;
    layer7_outputs(6475) <= a and not b;
    layer7_outputs(6476) <= not a or b;
    layer7_outputs(6477) <= a and not b;
    layer7_outputs(6478) <= a and not b;
    layer7_outputs(6479) <= b and not a;
    layer7_outputs(6480) <= not b;
    layer7_outputs(6481) <= not a or b;
    layer7_outputs(6482) <= not a;
    layer7_outputs(6483) <= a or b;
    layer7_outputs(6484) <= b;
    layer7_outputs(6485) <= a;
    layer7_outputs(6486) <= not b;
    layer7_outputs(6487) <= '0';
    layer7_outputs(6488) <= a and b;
    layer7_outputs(6489) <= '1';
    layer7_outputs(6490) <= '0';
    layer7_outputs(6491) <= b and not a;
    layer7_outputs(6492) <= a and b;
    layer7_outputs(6493) <= b;
    layer7_outputs(6494) <= a;
    layer7_outputs(6495) <= b;
    layer7_outputs(6496) <= not (a xor b);
    layer7_outputs(6497) <= not a;
    layer7_outputs(6498) <= not a;
    layer7_outputs(6499) <= a or b;
    layer7_outputs(6500) <= not b;
    layer7_outputs(6501) <= a xor b;
    layer7_outputs(6502) <= not a;
    layer7_outputs(6503) <= a;
    layer7_outputs(6504) <= b and not a;
    layer7_outputs(6505) <= a and not b;
    layer7_outputs(6506) <= not (a and b);
    layer7_outputs(6507) <= b;
    layer7_outputs(6508) <= a and b;
    layer7_outputs(6509) <= not (a and b);
    layer7_outputs(6510) <= b;
    layer7_outputs(6511) <= a and b;
    layer7_outputs(6512) <= not b;
    layer7_outputs(6513) <= not a or b;
    layer7_outputs(6514) <= a;
    layer7_outputs(6515) <= not b;
    layer7_outputs(6516) <= a or b;
    layer7_outputs(6517) <= a or b;
    layer7_outputs(6518) <= not (a or b);
    layer7_outputs(6519) <= not a;
    layer7_outputs(6520) <= not b;
    layer7_outputs(6521) <= not a;
    layer7_outputs(6522) <= a xor b;
    layer7_outputs(6523) <= not (a and b);
    layer7_outputs(6524) <= not (a or b);
    layer7_outputs(6525) <= a;
    layer7_outputs(6526) <= not b or a;
    layer7_outputs(6527) <= b;
    layer7_outputs(6528) <= a;
    layer7_outputs(6529) <= not (a or b);
    layer7_outputs(6530) <= not a;
    layer7_outputs(6531) <= b;
    layer7_outputs(6532) <= not (a or b);
    layer7_outputs(6533) <= b;
    layer7_outputs(6534) <= not b;
    layer7_outputs(6535) <= b;
    layer7_outputs(6536) <= a and b;
    layer7_outputs(6537) <= b;
    layer7_outputs(6538) <= not b;
    layer7_outputs(6539) <= not a;
    layer7_outputs(6540) <= not (a or b);
    layer7_outputs(6541) <= b;
    layer7_outputs(6542) <= not b;
    layer7_outputs(6543) <= not b;
    layer7_outputs(6544) <= b and not a;
    layer7_outputs(6545) <= not b or a;
    layer7_outputs(6546) <= a and b;
    layer7_outputs(6547) <= '0';
    layer7_outputs(6548) <= a xor b;
    layer7_outputs(6549) <= '0';
    layer7_outputs(6550) <= '1';
    layer7_outputs(6551) <= a;
    layer7_outputs(6552) <= a;
    layer7_outputs(6553) <= a and b;
    layer7_outputs(6554) <= not (a xor b);
    layer7_outputs(6555) <= a;
    layer7_outputs(6556) <= b and not a;
    layer7_outputs(6557) <= a;
    layer7_outputs(6558) <= not b;
    layer7_outputs(6559) <= not b;
    layer7_outputs(6560) <= a and b;
    layer7_outputs(6561) <= not b or a;
    layer7_outputs(6562) <= a;
    layer7_outputs(6563) <= a xor b;
    layer7_outputs(6564) <= a;
    layer7_outputs(6565) <= not b;
    layer7_outputs(6566) <= not a or b;
    layer7_outputs(6567) <= not a;
    layer7_outputs(6568) <= not a or b;
    layer7_outputs(6569) <= not b;
    layer7_outputs(6570) <= a;
    layer7_outputs(6571) <= a xor b;
    layer7_outputs(6572) <= a or b;
    layer7_outputs(6573) <= not a;
    layer7_outputs(6574) <= a and not b;
    layer7_outputs(6575) <= not a or b;
    layer7_outputs(6576) <= a xor b;
    layer7_outputs(6577) <= not (a xor b);
    layer7_outputs(6578) <= '0';
    layer7_outputs(6579) <= not b;
    layer7_outputs(6580) <= not b or a;
    layer7_outputs(6581) <= b;
    layer7_outputs(6582) <= a;
    layer7_outputs(6583) <= not a or b;
    layer7_outputs(6584) <= not b;
    layer7_outputs(6585) <= not a;
    layer7_outputs(6586) <= not b;
    layer7_outputs(6587) <= not b;
    layer7_outputs(6588) <= not (a or b);
    layer7_outputs(6589) <= a or b;
    layer7_outputs(6590) <= not a or b;
    layer7_outputs(6591) <= not b;
    layer7_outputs(6592) <= a;
    layer7_outputs(6593) <= b;
    layer7_outputs(6594) <= not (a xor b);
    layer7_outputs(6595) <= a and not b;
    layer7_outputs(6596) <= not a or b;
    layer7_outputs(6597) <= a and b;
    layer7_outputs(6598) <= '0';
    layer7_outputs(6599) <= not a;
    layer7_outputs(6600) <= not b or a;
    layer7_outputs(6601) <= not (a or b);
    layer7_outputs(6602) <= a;
    layer7_outputs(6603) <= not a or b;
    layer7_outputs(6604) <= not b or a;
    layer7_outputs(6605) <= a and b;
    layer7_outputs(6606) <= a;
    layer7_outputs(6607) <= not (a or b);
    layer7_outputs(6608) <= b;
    layer7_outputs(6609) <= not b;
    layer7_outputs(6610) <= not a or b;
    layer7_outputs(6611) <= not b;
    layer7_outputs(6612) <= a;
    layer7_outputs(6613) <= a or b;
    layer7_outputs(6614) <= a;
    layer7_outputs(6615) <= not (a and b);
    layer7_outputs(6616) <= not (a and b);
    layer7_outputs(6617) <= not b;
    layer7_outputs(6618) <= a;
    layer7_outputs(6619) <= not a;
    layer7_outputs(6620) <= not a;
    layer7_outputs(6621) <= a xor b;
    layer7_outputs(6622) <= a or b;
    layer7_outputs(6623) <= a and not b;
    layer7_outputs(6624) <= not b;
    layer7_outputs(6625) <= not a;
    layer7_outputs(6626) <= b;
    layer7_outputs(6627) <= not a or b;
    layer7_outputs(6628) <= b;
    layer7_outputs(6629) <= not b;
    layer7_outputs(6630) <= not a;
    layer7_outputs(6631) <= not b;
    layer7_outputs(6632) <= a;
    layer7_outputs(6633) <= not a;
    layer7_outputs(6634) <= a xor b;
    layer7_outputs(6635) <= a or b;
    layer7_outputs(6636) <= b;
    layer7_outputs(6637) <= b;
    layer7_outputs(6638) <= not (a and b);
    layer7_outputs(6639) <= b and not a;
    layer7_outputs(6640) <= a and not b;
    layer7_outputs(6641) <= b;
    layer7_outputs(6642) <= not a;
    layer7_outputs(6643) <= not (a or b);
    layer7_outputs(6644) <= b;
    layer7_outputs(6645) <= a and b;
    layer7_outputs(6646) <= not (a xor b);
    layer7_outputs(6647) <= a and not b;
    layer7_outputs(6648) <= not a or b;
    layer7_outputs(6649) <= not b or a;
    layer7_outputs(6650) <= a and b;
    layer7_outputs(6651) <= b;
    layer7_outputs(6652) <= not b;
    layer7_outputs(6653) <= a;
    layer7_outputs(6654) <= a and not b;
    layer7_outputs(6655) <= not (a xor b);
    layer7_outputs(6656) <= a;
    layer7_outputs(6657) <= a and not b;
    layer7_outputs(6658) <= a;
    layer7_outputs(6659) <= a;
    layer7_outputs(6660) <= not (a or b);
    layer7_outputs(6661) <= a xor b;
    layer7_outputs(6662) <= not (a or b);
    layer7_outputs(6663) <= not a;
    layer7_outputs(6664) <= not (a xor b);
    layer7_outputs(6665) <= '0';
    layer7_outputs(6666) <= not (a xor b);
    layer7_outputs(6667) <= not (a xor b);
    layer7_outputs(6668) <= b and not a;
    layer7_outputs(6669) <= not a;
    layer7_outputs(6670) <= not a or b;
    layer7_outputs(6671) <= b;
    layer7_outputs(6672) <= a and not b;
    layer7_outputs(6673) <= not (a and b);
    layer7_outputs(6674) <= b;
    layer7_outputs(6675) <= a xor b;
    layer7_outputs(6676) <= a;
    layer7_outputs(6677) <= not b;
    layer7_outputs(6678) <= not (a xor b);
    layer7_outputs(6679) <= a;
    layer7_outputs(6680) <= not b;
    layer7_outputs(6681) <= not (a and b);
    layer7_outputs(6682) <= not (a xor b);
    layer7_outputs(6683) <= not (a xor b);
    layer7_outputs(6684) <= a xor b;
    layer7_outputs(6685) <= a and not b;
    layer7_outputs(6686) <= b;
    layer7_outputs(6687) <= a and b;
    layer7_outputs(6688) <= a and not b;
    layer7_outputs(6689) <= b;
    layer7_outputs(6690) <= a xor b;
    layer7_outputs(6691) <= not (a xor b);
    layer7_outputs(6692) <= not b;
    layer7_outputs(6693) <= not b or a;
    layer7_outputs(6694) <= not (a or b);
    layer7_outputs(6695) <= a or b;
    layer7_outputs(6696) <= not b or a;
    layer7_outputs(6697) <= a and b;
    layer7_outputs(6698) <= b;
    layer7_outputs(6699) <= not b;
    layer7_outputs(6700) <= a and not b;
    layer7_outputs(6701) <= a or b;
    layer7_outputs(6702) <= b;
    layer7_outputs(6703) <= not b;
    layer7_outputs(6704) <= a or b;
    layer7_outputs(6705) <= not b or a;
    layer7_outputs(6706) <= not b;
    layer7_outputs(6707) <= not b;
    layer7_outputs(6708) <= a and b;
    layer7_outputs(6709) <= b;
    layer7_outputs(6710) <= a;
    layer7_outputs(6711) <= a and b;
    layer7_outputs(6712) <= not a;
    layer7_outputs(6713) <= b;
    layer7_outputs(6714) <= b;
    layer7_outputs(6715) <= a;
    layer7_outputs(6716) <= b and not a;
    layer7_outputs(6717) <= not b or a;
    layer7_outputs(6718) <= not b or a;
    layer7_outputs(6719) <= not (a and b);
    layer7_outputs(6720) <= not (a and b);
    layer7_outputs(6721) <= not b;
    layer7_outputs(6722) <= b;
    layer7_outputs(6723) <= a and b;
    layer7_outputs(6724) <= not b;
    layer7_outputs(6725) <= not b;
    layer7_outputs(6726) <= not b;
    layer7_outputs(6727) <= b and not a;
    layer7_outputs(6728) <= not a or b;
    layer7_outputs(6729) <= b;
    layer7_outputs(6730) <= not a;
    layer7_outputs(6731) <= a and not b;
    layer7_outputs(6732) <= not a;
    layer7_outputs(6733) <= not b or a;
    layer7_outputs(6734) <= a;
    layer7_outputs(6735) <= not b or a;
    layer7_outputs(6736) <= not (a and b);
    layer7_outputs(6737) <= a and not b;
    layer7_outputs(6738) <= not a or b;
    layer7_outputs(6739) <= not (a or b);
    layer7_outputs(6740) <= a;
    layer7_outputs(6741) <= not a or b;
    layer7_outputs(6742) <= b and not a;
    layer7_outputs(6743) <= not (a xor b);
    layer7_outputs(6744) <= a or b;
    layer7_outputs(6745) <= a;
    layer7_outputs(6746) <= a xor b;
    layer7_outputs(6747) <= a;
    layer7_outputs(6748) <= not b or a;
    layer7_outputs(6749) <= a and b;
    layer7_outputs(6750) <= not (a and b);
    layer7_outputs(6751) <= b;
    layer7_outputs(6752) <= b;
    layer7_outputs(6753) <= not b;
    layer7_outputs(6754) <= not (a and b);
    layer7_outputs(6755) <= not a;
    layer7_outputs(6756) <= not (a xor b);
    layer7_outputs(6757) <= a and b;
    layer7_outputs(6758) <= a and b;
    layer7_outputs(6759) <= b;
    layer7_outputs(6760) <= not b or a;
    layer7_outputs(6761) <= not (a or b);
    layer7_outputs(6762) <= b;
    layer7_outputs(6763) <= not a;
    layer7_outputs(6764) <= not a or b;
    layer7_outputs(6765) <= not b or a;
    layer7_outputs(6766) <= a and not b;
    layer7_outputs(6767) <= not b;
    layer7_outputs(6768) <= a and b;
    layer7_outputs(6769) <= not (a xor b);
    layer7_outputs(6770) <= not (a and b);
    layer7_outputs(6771) <= b;
    layer7_outputs(6772) <= not a or b;
    layer7_outputs(6773) <= b;
    layer7_outputs(6774) <= a;
    layer7_outputs(6775) <= not b;
    layer7_outputs(6776) <= not b or a;
    layer7_outputs(6777) <= a;
    layer7_outputs(6778) <= b;
    layer7_outputs(6779) <= not b;
    layer7_outputs(6780) <= a;
    layer7_outputs(6781) <= not (a xor b);
    layer7_outputs(6782) <= a or b;
    layer7_outputs(6783) <= not (a and b);
    layer7_outputs(6784) <= not b;
    layer7_outputs(6785) <= not a;
    layer7_outputs(6786) <= not (a xor b);
    layer7_outputs(6787) <= a;
    layer7_outputs(6788) <= a;
    layer7_outputs(6789) <= b;
    layer7_outputs(6790) <= a or b;
    layer7_outputs(6791) <= b;
    layer7_outputs(6792) <= not a;
    layer7_outputs(6793) <= not a or b;
    layer7_outputs(6794) <= b and not a;
    layer7_outputs(6795) <= not a or b;
    layer7_outputs(6796) <= a and not b;
    layer7_outputs(6797) <= not a;
    layer7_outputs(6798) <= not b or a;
    layer7_outputs(6799) <= a;
    layer7_outputs(6800) <= a and b;
    layer7_outputs(6801) <= not b or a;
    layer7_outputs(6802) <= not (a and b);
    layer7_outputs(6803) <= not (a xor b);
    layer7_outputs(6804) <= not b;
    layer7_outputs(6805) <= not a;
    layer7_outputs(6806) <= not (a xor b);
    layer7_outputs(6807) <= a or b;
    layer7_outputs(6808) <= not a or b;
    layer7_outputs(6809) <= not b or a;
    layer7_outputs(6810) <= b;
    layer7_outputs(6811) <= not (a xor b);
    layer7_outputs(6812) <= not a;
    layer7_outputs(6813) <= not b;
    layer7_outputs(6814) <= a;
    layer7_outputs(6815) <= not (a xor b);
    layer7_outputs(6816) <= not (a and b);
    layer7_outputs(6817) <= a;
    layer7_outputs(6818) <= a xor b;
    layer7_outputs(6819) <= a or b;
    layer7_outputs(6820) <= not a;
    layer7_outputs(6821) <= a and b;
    layer7_outputs(6822) <= not a or b;
    layer7_outputs(6823) <= not a;
    layer7_outputs(6824) <= not b or a;
    layer7_outputs(6825) <= not (a xor b);
    layer7_outputs(6826) <= a;
    layer7_outputs(6827) <= b;
    layer7_outputs(6828) <= not b or a;
    layer7_outputs(6829) <= a or b;
    layer7_outputs(6830) <= not b;
    layer7_outputs(6831) <= not a or b;
    layer7_outputs(6832) <= not a;
    layer7_outputs(6833) <= a and b;
    layer7_outputs(6834) <= b;
    layer7_outputs(6835) <= not a;
    layer7_outputs(6836) <= not (a or b);
    layer7_outputs(6837) <= not a;
    layer7_outputs(6838) <= not a;
    layer7_outputs(6839) <= b;
    layer7_outputs(6840) <= not (a xor b);
    layer7_outputs(6841) <= a or b;
    layer7_outputs(6842) <= not b;
    layer7_outputs(6843) <= not (a or b);
    layer7_outputs(6844) <= a and b;
    layer7_outputs(6845) <= a and b;
    layer7_outputs(6846) <= not a;
    layer7_outputs(6847) <= not b;
    layer7_outputs(6848) <= not a;
    layer7_outputs(6849) <= not (a and b);
    layer7_outputs(6850) <= not (a xor b);
    layer7_outputs(6851) <= not (a and b);
    layer7_outputs(6852) <= b and not a;
    layer7_outputs(6853) <= a and b;
    layer7_outputs(6854) <= a xor b;
    layer7_outputs(6855) <= not a;
    layer7_outputs(6856) <= not b or a;
    layer7_outputs(6857) <= b;
    layer7_outputs(6858) <= b;
    layer7_outputs(6859) <= a;
    layer7_outputs(6860) <= not b or a;
    layer7_outputs(6861) <= not a;
    layer7_outputs(6862) <= not a;
    layer7_outputs(6863) <= a and not b;
    layer7_outputs(6864) <= not b;
    layer7_outputs(6865) <= not (a or b);
    layer7_outputs(6866) <= a;
    layer7_outputs(6867) <= b;
    layer7_outputs(6868) <= a and not b;
    layer7_outputs(6869) <= a;
    layer7_outputs(6870) <= not a;
    layer7_outputs(6871) <= not a;
    layer7_outputs(6872) <= '1';
    layer7_outputs(6873) <= not a or b;
    layer7_outputs(6874) <= a xor b;
    layer7_outputs(6875) <= b and not a;
    layer7_outputs(6876) <= not b;
    layer7_outputs(6877) <= a and b;
    layer7_outputs(6878) <= a and not b;
    layer7_outputs(6879) <= not (a or b);
    layer7_outputs(6880) <= not a;
    layer7_outputs(6881) <= a xor b;
    layer7_outputs(6882) <= b and not a;
    layer7_outputs(6883) <= a and b;
    layer7_outputs(6884) <= a or b;
    layer7_outputs(6885) <= a xor b;
    layer7_outputs(6886) <= a;
    layer7_outputs(6887) <= a;
    layer7_outputs(6888) <= not (a xor b);
    layer7_outputs(6889) <= a or b;
    layer7_outputs(6890) <= not a;
    layer7_outputs(6891) <= a and b;
    layer7_outputs(6892) <= '0';
    layer7_outputs(6893) <= a;
    layer7_outputs(6894) <= b and not a;
    layer7_outputs(6895) <= not (a and b);
    layer7_outputs(6896) <= not a;
    layer7_outputs(6897) <= a;
    layer7_outputs(6898) <= a;
    layer7_outputs(6899) <= not b;
    layer7_outputs(6900) <= b;
    layer7_outputs(6901) <= a or b;
    layer7_outputs(6902) <= not (a and b);
    layer7_outputs(6903) <= not a;
    layer7_outputs(6904) <= not b or a;
    layer7_outputs(6905) <= a and b;
    layer7_outputs(6906) <= a or b;
    layer7_outputs(6907) <= '0';
    layer7_outputs(6908) <= a and b;
    layer7_outputs(6909) <= not b;
    layer7_outputs(6910) <= b;
    layer7_outputs(6911) <= a and not b;
    layer7_outputs(6912) <= not b or a;
    layer7_outputs(6913) <= a and not b;
    layer7_outputs(6914) <= a and not b;
    layer7_outputs(6915) <= a or b;
    layer7_outputs(6916) <= not a or b;
    layer7_outputs(6917) <= a;
    layer7_outputs(6918) <= not a;
    layer7_outputs(6919) <= not a;
    layer7_outputs(6920) <= b;
    layer7_outputs(6921) <= not b or a;
    layer7_outputs(6922) <= not b or a;
    layer7_outputs(6923) <= a xor b;
    layer7_outputs(6924) <= b and not a;
    layer7_outputs(6925) <= not (a or b);
    layer7_outputs(6926) <= a and b;
    layer7_outputs(6927) <= a and b;
    layer7_outputs(6928) <= not b;
    layer7_outputs(6929) <= a and not b;
    layer7_outputs(6930) <= not a or b;
    layer7_outputs(6931) <= not (a or b);
    layer7_outputs(6932) <= '0';
    layer7_outputs(6933) <= not a or b;
    layer7_outputs(6934) <= a;
    layer7_outputs(6935) <= not (a or b);
    layer7_outputs(6936) <= not a;
    layer7_outputs(6937) <= a or b;
    layer7_outputs(6938) <= a or b;
    layer7_outputs(6939) <= not (a xor b);
    layer7_outputs(6940) <= not b;
    layer7_outputs(6941) <= not b;
    layer7_outputs(6942) <= a;
    layer7_outputs(6943) <= a xor b;
    layer7_outputs(6944) <= a;
    layer7_outputs(6945) <= not (a and b);
    layer7_outputs(6946) <= not b;
    layer7_outputs(6947) <= b and not a;
    layer7_outputs(6948) <= not b;
    layer7_outputs(6949) <= b;
    layer7_outputs(6950) <= '0';
    layer7_outputs(6951) <= '0';
    layer7_outputs(6952) <= b;
    layer7_outputs(6953) <= not b;
    layer7_outputs(6954) <= not b;
    layer7_outputs(6955) <= not (a and b);
    layer7_outputs(6956) <= a xor b;
    layer7_outputs(6957) <= not (a xor b);
    layer7_outputs(6958) <= not a or b;
    layer7_outputs(6959) <= not b;
    layer7_outputs(6960) <= a and not b;
    layer7_outputs(6961) <= not (a xor b);
    layer7_outputs(6962) <= not a;
    layer7_outputs(6963) <= a;
    layer7_outputs(6964) <= not (a or b);
    layer7_outputs(6965) <= '0';
    layer7_outputs(6966) <= not (a xor b);
    layer7_outputs(6967) <= b and not a;
    layer7_outputs(6968) <= a and b;
    layer7_outputs(6969) <= a xor b;
    layer7_outputs(6970) <= not a or b;
    layer7_outputs(6971) <= not a;
    layer7_outputs(6972) <= a and b;
    layer7_outputs(6973) <= a xor b;
    layer7_outputs(6974) <= not a;
    layer7_outputs(6975) <= not (a and b);
    layer7_outputs(6976) <= not b;
    layer7_outputs(6977) <= a or b;
    layer7_outputs(6978) <= not a or b;
    layer7_outputs(6979) <= not (a and b);
    layer7_outputs(6980) <= a;
    layer7_outputs(6981) <= not (a xor b);
    layer7_outputs(6982) <= a;
    layer7_outputs(6983) <= not a or b;
    layer7_outputs(6984) <= not b;
    layer7_outputs(6985) <= not b or a;
    layer7_outputs(6986) <= not a;
    layer7_outputs(6987) <= a and b;
    layer7_outputs(6988) <= not (a or b);
    layer7_outputs(6989) <= not (a or b);
    layer7_outputs(6990) <= not a or b;
    layer7_outputs(6991) <= a and not b;
    layer7_outputs(6992) <= not a or b;
    layer7_outputs(6993) <= not (a or b);
    layer7_outputs(6994) <= not (a or b);
    layer7_outputs(6995) <= not (a xor b);
    layer7_outputs(6996) <= not a;
    layer7_outputs(6997) <= a xor b;
    layer7_outputs(6998) <= not a or b;
    layer7_outputs(6999) <= a;
    layer7_outputs(7000) <= b;
    layer7_outputs(7001) <= a and not b;
    layer7_outputs(7002) <= not b;
    layer7_outputs(7003) <= not a or b;
    layer7_outputs(7004) <= not b or a;
    layer7_outputs(7005) <= not a;
    layer7_outputs(7006) <= b and not a;
    layer7_outputs(7007) <= a;
    layer7_outputs(7008) <= a;
    layer7_outputs(7009) <= a xor b;
    layer7_outputs(7010) <= a or b;
    layer7_outputs(7011) <= a or b;
    layer7_outputs(7012) <= a and not b;
    layer7_outputs(7013) <= not (a xor b);
    layer7_outputs(7014) <= b;
    layer7_outputs(7015) <= b;
    layer7_outputs(7016) <= a and not b;
    layer7_outputs(7017) <= not a or b;
    layer7_outputs(7018) <= not a or b;
    layer7_outputs(7019) <= a or b;
    layer7_outputs(7020) <= not b or a;
    layer7_outputs(7021) <= not a;
    layer7_outputs(7022) <= b and not a;
    layer7_outputs(7023) <= b;
    layer7_outputs(7024) <= a xor b;
    layer7_outputs(7025) <= a and not b;
    layer7_outputs(7026) <= a and not b;
    layer7_outputs(7027) <= a or b;
    layer7_outputs(7028) <= not b or a;
    layer7_outputs(7029) <= not a or b;
    layer7_outputs(7030) <= not a;
    layer7_outputs(7031) <= not b;
    layer7_outputs(7032) <= b;
    layer7_outputs(7033) <= not a;
    layer7_outputs(7034) <= not b;
    layer7_outputs(7035) <= not b;
    layer7_outputs(7036) <= not (a or b);
    layer7_outputs(7037) <= not a or b;
    layer7_outputs(7038) <= a;
    layer7_outputs(7039) <= a or b;
    layer7_outputs(7040) <= not b;
    layer7_outputs(7041) <= not b;
    layer7_outputs(7042) <= a xor b;
    layer7_outputs(7043) <= a xor b;
    layer7_outputs(7044) <= b;
    layer7_outputs(7045) <= b;
    layer7_outputs(7046) <= a;
    layer7_outputs(7047) <= not (a and b);
    layer7_outputs(7048) <= '1';
    layer7_outputs(7049) <= '1';
    layer7_outputs(7050) <= a;
    layer7_outputs(7051) <= b;
    layer7_outputs(7052) <= not a;
    layer7_outputs(7053) <= a or b;
    layer7_outputs(7054) <= b and not a;
    layer7_outputs(7055) <= not (a and b);
    layer7_outputs(7056) <= not b;
    layer7_outputs(7057) <= a xor b;
    layer7_outputs(7058) <= a;
    layer7_outputs(7059) <= a;
    layer7_outputs(7060) <= not (a and b);
    layer7_outputs(7061) <= not (a xor b);
    layer7_outputs(7062) <= not a or b;
    layer7_outputs(7063) <= a and not b;
    layer7_outputs(7064) <= not a or b;
    layer7_outputs(7065) <= '0';
    layer7_outputs(7066) <= '1';
    layer7_outputs(7067) <= a and not b;
    layer7_outputs(7068) <= a;
    layer7_outputs(7069) <= not (a xor b);
    layer7_outputs(7070) <= a xor b;
    layer7_outputs(7071) <= '0';
    layer7_outputs(7072) <= not (a xor b);
    layer7_outputs(7073) <= not (a or b);
    layer7_outputs(7074) <= b;
    layer7_outputs(7075) <= a;
    layer7_outputs(7076) <= a and not b;
    layer7_outputs(7077) <= a and b;
    layer7_outputs(7078) <= not (a and b);
    layer7_outputs(7079) <= not a or b;
    layer7_outputs(7080) <= b and not a;
    layer7_outputs(7081) <= not b;
    layer7_outputs(7082) <= b;
    layer7_outputs(7083) <= a;
    layer7_outputs(7084) <= not (a xor b);
    layer7_outputs(7085) <= not a;
    layer7_outputs(7086) <= a or b;
    layer7_outputs(7087) <= not a;
    layer7_outputs(7088) <= not b;
    layer7_outputs(7089) <= not b or a;
    layer7_outputs(7090) <= a xor b;
    layer7_outputs(7091) <= not (a xor b);
    layer7_outputs(7092) <= not a;
    layer7_outputs(7093) <= a xor b;
    layer7_outputs(7094) <= not (a and b);
    layer7_outputs(7095) <= b;
    layer7_outputs(7096) <= a;
    layer7_outputs(7097) <= a and not b;
    layer7_outputs(7098) <= '1';
    layer7_outputs(7099) <= a;
    layer7_outputs(7100) <= a;
    layer7_outputs(7101) <= b and not a;
    layer7_outputs(7102) <= not b;
    layer7_outputs(7103) <= a or b;
    layer7_outputs(7104) <= a;
    layer7_outputs(7105) <= a or b;
    layer7_outputs(7106) <= not a or b;
    layer7_outputs(7107) <= b;
    layer7_outputs(7108) <= not b;
    layer7_outputs(7109) <= a;
    layer7_outputs(7110) <= b;
    layer7_outputs(7111) <= a or b;
    layer7_outputs(7112) <= not a;
    layer7_outputs(7113) <= a;
    layer7_outputs(7114) <= not b or a;
    layer7_outputs(7115) <= not a;
    layer7_outputs(7116) <= not a;
    layer7_outputs(7117) <= not b;
    layer7_outputs(7118) <= a;
    layer7_outputs(7119) <= not a;
    layer7_outputs(7120) <= b;
    layer7_outputs(7121) <= a and not b;
    layer7_outputs(7122) <= b and not a;
    layer7_outputs(7123) <= not (a and b);
    layer7_outputs(7124) <= not a or b;
    layer7_outputs(7125) <= b and not a;
    layer7_outputs(7126) <= a;
    layer7_outputs(7127) <= a and b;
    layer7_outputs(7128) <= b;
    layer7_outputs(7129) <= not (a or b);
    layer7_outputs(7130) <= a and not b;
    layer7_outputs(7131) <= not b;
    layer7_outputs(7132) <= not (a or b);
    layer7_outputs(7133) <= a and not b;
    layer7_outputs(7134) <= not a;
    layer7_outputs(7135) <= a;
    layer7_outputs(7136) <= b;
    layer7_outputs(7137) <= not b;
    layer7_outputs(7138) <= a xor b;
    layer7_outputs(7139) <= b;
    layer7_outputs(7140) <= a and not b;
    layer7_outputs(7141) <= a and not b;
    layer7_outputs(7142) <= not b or a;
    layer7_outputs(7143) <= a xor b;
    layer7_outputs(7144) <= not (a xor b);
    layer7_outputs(7145) <= not b;
    layer7_outputs(7146) <= b and not a;
    layer7_outputs(7147) <= not (a or b);
    layer7_outputs(7148) <= a;
    layer7_outputs(7149) <= b and not a;
    layer7_outputs(7150) <= b and not a;
    layer7_outputs(7151) <= not (a and b);
    layer7_outputs(7152) <= a and not b;
    layer7_outputs(7153) <= not b;
    layer7_outputs(7154) <= a and b;
    layer7_outputs(7155) <= b and not a;
    layer7_outputs(7156) <= not (a xor b);
    layer7_outputs(7157) <= a xor b;
    layer7_outputs(7158) <= not (a or b);
    layer7_outputs(7159) <= b;
    layer7_outputs(7160) <= not (a and b);
    layer7_outputs(7161) <= a xor b;
    layer7_outputs(7162) <= a;
    layer7_outputs(7163) <= not b;
    layer7_outputs(7164) <= a;
    layer7_outputs(7165) <= not b or a;
    layer7_outputs(7166) <= a;
    layer7_outputs(7167) <= a and b;
    layer7_outputs(7168) <= b and not a;
    layer7_outputs(7169) <= b;
    layer7_outputs(7170) <= b;
    layer7_outputs(7171) <= not (a xor b);
    layer7_outputs(7172) <= a or b;
    layer7_outputs(7173) <= not a or b;
    layer7_outputs(7174) <= not (a and b);
    layer7_outputs(7175) <= not a or b;
    layer7_outputs(7176) <= b and not a;
    layer7_outputs(7177) <= a and b;
    layer7_outputs(7178) <= not a;
    layer7_outputs(7179) <= not b;
    layer7_outputs(7180) <= not b or a;
    layer7_outputs(7181) <= not (a xor b);
    layer7_outputs(7182) <= a xor b;
    layer7_outputs(7183) <= not b or a;
    layer7_outputs(7184) <= b;
    layer7_outputs(7185) <= a and b;
    layer7_outputs(7186) <= b and not a;
    layer7_outputs(7187) <= a xor b;
    layer7_outputs(7188) <= b and not a;
    layer7_outputs(7189) <= a;
    layer7_outputs(7190) <= a and not b;
    layer7_outputs(7191) <= not a;
    layer7_outputs(7192) <= '1';
    layer7_outputs(7193) <= not (a xor b);
    layer7_outputs(7194) <= a;
    layer7_outputs(7195) <= a and b;
    layer7_outputs(7196) <= not b;
    layer7_outputs(7197) <= a xor b;
    layer7_outputs(7198) <= not a;
    layer7_outputs(7199) <= a and not b;
    layer7_outputs(7200) <= a;
    layer7_outputs(7201) <= not b;
    layer7_outputs(7202) <= a or b;
    layer7_outputs(7203) <= not (a or b);
    layer7_outputs(7204) <= a or b;
    layer7_outputs(7205) <= a and b;
    layer7_outputs(7206) <= b;
    layer7_outputs(7207) <= b;
    layer7_outputs(7208) <= not (a and b);
    layer7_outputs(7209) <= a and not b;
    layer7_outputs(7210) <= a xor b;
    layer7_outputs(7211) <= a and b;
    layer7_outputs(7212) <= not a or b;
    layer7_outputs(7213) <= b;
    layer7_outputs(7214) <= '1';
    layer7_outputs(7215) <= not a;
    layer7_outputs(7216) <= a and not b;
    layer7_outputs(7217) <= not (a or b);
    layer7_outputs(7218) <= not b;
    layer7_outputs(7219) <= a;
    layer7_outputs(7220) <= a;
    layer7_outputs(7221) <= a;
    layer7_outputs(7222) <= not b;
    layer7_outputs(7223) <= not b;
    layer7_outputs(7224) <= not (a and b);
    layer7_outputs(7225) <= not a;
    layer7_outputs(7226) <= not b;
    layer7_outputs(7227) <= b and not a;
    layer7_outputs(7228) <= a;
    layer7_outputs(7229) <= not b;
    layer7_outputs(7230) <= not (a or b);
    layer7_outputs(7231) <= '1';
    layer7_outputs(7232) <= a and not b;
    layer7_outputs(7233) <= '1';
    layer7_outputs(7234) <= not b;
    layer7_outputs(7235) <= b and not a;
    layer7_outputs(7236) <= not a;
    layer7_outputs(7237) <= b and not a;
    layer7_outputs(7238) <= a and b;
    layer7_outputs(7239) <= a xor b;
    layer7_outputs(7240) <= not b or a;
    layer7_outputs(7241) <= not b;
    layer7_outputs(7242) <= not b or a;
    layer7_outputs(7243) <= not a or b;
    layer7_outputs(7244) <= a and b;
    layer7_outputs(7245) <= not b;
    layer7_outputs(7246) <= not b;
    layer7_outputs(7247) <= not (a or b);
    layer7_outputs(7248) <= a;
    layer7_outputs(7249) <= b and not a;
    layer7_outputs(7250) <= not b;
    layer7_outputs(7251) <= b;
    layer7_outputs(7252) <= b;
    layer7_outputs(7253) <= not a or b;
    layer7_outputs(7254) <= not a;
    layer7_outputs(7255) <= a xor b;
    layer7_outputs(7256) <= a and not b;
    layer7_outputs(7257) <= a;
    layer7_outputs(7258) <= b and not a;
    layer7_outputs(7259) <= b;
    layer7_outputs(7260) <= not (a or b);
    layer7_outputs(7261) <= not a;
    layer7_outputs(7262) <= b and not a;
    layer7_outputs(7263) <= not b or a;
    layer7_outputs(7264) <= b and not a;
    layer7_outputs(7265) <= b;
    layer7_outputs(7266) <= b and not a;
    layer7_outputs(7267) <= not (a and b);
    layer7_outputs(7268) <= b;
    layer7_outputs(7269) <= not (a xor b);
    layer7_outputs(7270) <= not a;
    layer7_outputs(7271) <= not (a or b);
    layer7_outputs(7272) <= a xor b;
    layer7_outputs(7273) <= a or b;
    layer7_outputs(7274) <= a xor b;
    layer7_outputs(7275) <= a xor b;
    layer7_outputs(7276) <= b;
    layer7_outputs(7277) <= not (a and b);
    layer7_outputs(7278) <= a and not b;
    layer7_outputs(7279) <= not (a xor b);
    layer7_outputs(7280) <= a;
    layer7_outputs(7281) <= a xor b;
    layer7_outputs(7282) <= not a or b;
    layer7_outputs(7283) <= b;
    layer7_outputs(7284) <= a;
    layer7_outputs(7285) <= b and not a;
    layer7_outputs(7286) <= not a;
    layer7_outputs(7287) <= b and not a;
    layer7_outputs(7288) <= a;
    layer7_outputs(7289) <= a;
    layer7_outputs(7290) <= b;
    layer7_outputs(7291) <= a xor b;
    layer7_outputs(7292) <= not b;
    layer7_outputs(7293) <= '0';
    layer7_outputs(7294) <= not a;
    layer7_outputs(7295) <= b and not a;
    layer7_outputs(7296) <= a and b;
    layer7_outputs(7297) <= not (a or b);
    layer7_outputs(7298) <= a;
    layer7_outputs(7299) <= b;
    layer7_outputs(7300) <= not (a or b);
    layer7_outputs(7301) <= a;
    layer7_outputs(7302) <= not a or b;
    layer7_outputs(7303) <= not b;
    layer7_outputs(7304) <= a;
    layer7_outputs(7305) <= a;
    layer7_outputs(7306) <= b;
    layer7_outputs(7307) <= not (a xor b);
    layer7_outputs(7308) <= not b;
    layer7_outputs(7309) <= not a;
    layer7_outputs(7310) <= not a;
    layer7_outputs(7311) <= not a or b;
    layer7_outputs(7312) <= b and not a;
    layer7_outputs(7313) <= a xor b;
    layer7_outputs(7314) <= a and not b;
    layer7_outputs(7315) <= not b;
    layer7_outputs(7316) <= not a;
    layer7_outputs(7317) <= not a;
    layer7_outputs(7318) <= b;
    layer7_outputs(7319) <= b;
    layer7_outputs(7320) <= a and b;
    layer7_outputs(7321) <= not a;
    layer7_outputs(7322) <= b;
    layer7_outputs(7323) <= not (a or b);
    layer7_outputs(7324) <= not b;
    layer7_outputs(7325) <= b and not a;
    layer7_outputs(7326) <= not (a and b);
    layer7_outputs(7327) <= not (a xor b);
    layer7_outputs(7328) <= not a;
    layer7_outputs(7329) <= not b;
    layer7_outputs(7330) <= not b;
    layer7_outputs(7331) <= b and not a;
    layer7_outputs(7332) <= not a;
    layer7_outputs(7333) <= a and not b;
    layer7_outputs(7334) <= not b;
    layer7_outputs(7335) <= not (a xor b);
    layer7_outputs(7336) <= a;
    layer7_outputs(7337) <= not (a xor b);
    layer7_outputs(7338) <= not a;
    layer7_outputs(7339) <= a or b;
    layer7_outputs(7340) <= a or b;
    layer7_outputs(7341) <= a and not b;
    layer7_outputs(7342) <= not (a xor b);
    layer7_outputs(7343) <= not a;
    layer7_outputs(7344) <= b and not a;
    layer7_outputs(7345) <= not a or b;
    layer7_outputs(7346) <= b and not a;
    layer7_outputs(7347) <= b and not a;
    layer7_outputs(7348) <= not b;
    layer7_outputs(7349) <= a xor b;
    layer7_outputs(7350) <= not b or a;
    layer7_outputs(7351) <= a and not b;
    layer7_outputs(7352) <= a and b;
    layer7_outputs(7353) <= a xor b;
    layer7_outputs(7354) <= not (a or b);
    layer7_outputs(7355) <= not b or a;
    layer7_outputs(7356) <= not b or a;
    layer7_outputs(7357) <= a and b;
    layer7_outputs(7358) <= a and b;
    layer7_outputs(7359) <= '0';
    layer7_outputs(7360) <= not (a xor b);
    layer7_outputs(7361) <= a or b;
    layer7_outputs(7362) <= a;
    layer7_outputs(7363) <= a;
    layer7_outputs(7364) <= b and not a;
    layer7_outputs(7365) <= not (a and b);
    layer7_outputs(7366) <= not a or b;
    layer7_outputs(7367) <= a and b;
    layer7_outputs(7368) <= not (a or b);
    layer7_outputs(7369) <= not a;
    layer7_outputs(7370) <= a and not b;
    layer7_outputs(7371) <= a xor b;
    layer7_outputs(7372) <= a or b;
    layer7_outputs(7373) <= a and b;
    layer7_outputs(7374) <= a;
    layer7_outputs(7375) <= '0';
    layer7_outputs(7376) <= not b;
    layer7_outputs(7377) <= a;
    layer7_outputs(7378) <= not (a or b);
    layer7_outputs(7379) <= a;
    layer7_outputs(7380) <= not b;
    layer7_outputs(7381) <= not b;
    layer7_outputs(7382) <= not a;
    layer7_outputs(7383) <= not b;
    layer7_outputs(7384) <= not (a or b);
    layer7_outputs(7385) <= a or b;
    layer7_outputs(7386) <= not b;
    layer7_outputs(7387) <= a;
    layer7_outputs(7388) <= not b;
    layer7_outputs(7389) <= b and not a;
    layer7_outputs(7390) <= a and b;
    layer7_outputs(7391) <= not (a xor b);
    layer7_outputs(7392) <= not a;
    layer7_outputs(7393) <= not (a or b);
    layer7_outputs(7394) <= not (a and b);
    layer7_outputs(7395) <= a;
    layer7_outputs(7396) <= not (a xor b);
    layer7_outputs(7397) <= not (a or b);
    layer7_outputs(7398) <= not b;
    layer7_outputs(7399) <= not (a xor b);
    layer7_outputs(7400) <= a and b;
    layer7_outputs(7401) <= a and b;
    layer7_outputs(7402) <= not (a or b);
    layer7_outputs(7403) <= not (a xor b);
    layer7_outputs(7404) <= b;
    layer7_outputs(7405) <= a xor b;
    layer7_outputs(7406) <= b and not a;
    layer7_outputs(7407) <= a or b;
    layer7_outputs(7408) <= b;
    layer7_outputs(7409) <= a and b;
    layer7_outputs(7410) <= not a;
    layer7_outputs(7411) <= a and b;
    layer7_outputs(7412) <= a xor b;
    layer7_outputs(7413) <= a and b;
    layer7_outputs(7414) <= b and not a;
    layer7_outputs(7415) <= a and b;
    layer7_outputs(7416) <= not (a or b);
    layer7_outputs(7417) <= not (a xor b);
    layer7_outputs(7418) <= not b;
    layer7_outputs(7419) <= a or b;
    layer7_outputs(7420) <= not a;
    layer7_outputs(7421) <= not b or a;
    layer7_outputs(7422) <= not a or b;
    layer7_outputs(7423) <= a xor b;
    layer7_outputs(7424) <= b;
    layer7_outputs(7425) <= a and not b;
    layer7_outputs(7426) <= not a;
    layer7_outputs(7427) <= not a or b;
    layer7_outputs(7428) <= b and not a;
    layer7_outputs(7429) <= b;
    layer7_outputs(7430) <= b;
    layer7_outputs(7431) <= a and not b;
    layer7_outputs(7432) <= a xor b;
    layer7_outputs(7433) <= not (a or b);
    layer7_outputs(7434) <= a and not b;
    layer7_outputs(7435) <= b;
    layer7_outputs(7436) <= not (a and b);
    layer7_outputs(7437) <= a and not b;
    layer7_outputs(7438) <= b and not a;
    layer7_outputs(7439) <= not (a or b);
    layer7_outputs(7440) <= not a;
    layer7_outputs(7441) <= not a or b;
    layer7_outputs(7442) <= not b or a;
    layer7_outputs(7443) <= b;
    layer7_outputs(7444) <= not (a or b);
    layer7_outputs(7445) <= a and not b;
    layer7_outputs(7446) <= not b;
    layer7_outputs(7447) <= not a or b;
    layer7_outputs(7448) <= not a;
    layer7_outputs(7449) <= not a or b;
    layer7_outputs(7450) <= not (a or b);
    layer7_outputs(7451) <= not (a or b);
    layer7_outputs(7452) <= a;
    layer7_outputs(7453) <= not b;
    layer7_outputs(7454) <= not a;
    layer7_outputs(7455) <= a or b;
    layer7_outputs(7456) <= a and not b;
    layer7_outputs(7457) <= a;
    layer7_outputs(7458) <= a;
    layer7_outputs(7459) <= b;
    layer7_outputs(7460) <= a xor b;
    layer7_outputs(7461) <= a;
    layer7_outputs(7462) <= not (a xor b);
    layer7_outputs(7463) <= not b;
    layer7_outputs(7464) <= a and b;
    layer7_outputs(7465) <= a xor b;
    layer7_outputs(7466) <= not b or a;
    layer7_outputs(7467) <= not b;
    layer7_outputs(7468) <= a;
    layer7_outputs(7469) <= not (a and b);
    layer7_outputs(7470) <= not (a and b);
    layer7_outputs(7471) <= a;
    layer7_outputs(7472) <= not a;
    layer7_outputs(7473) <= a or b;
    layer7_outputs(7474) <= a;
    layer7_outputs(7475) <= not b or a;
    layer7_outputs(7476) <= b;
    layer7_outputs(7477) <= not b or a;
    layer7_outputs(7478) <= not a;
    layer7_outputs(7479) <= '1';
    layer7_outputs(7480) <= b;
    layer7_outputs(7481) <= not b;
    layer7_outputs(7482) <= not a;
    layer7_outputs(7483) <= not a or b;
    layer7_outputs(7484) <= not (a or b);
    layer7_outputs(7485) <= a and not b;
    layer7_outputs(7486) <= a and not b;
    layer7_outputs(7487) <= not (a and b);
    layer7_outputs(7488) <= b;
    layer7_outputs(7489) <= b and not a;
    layer7_outputs(7490) <= a and b;
    layer7_outputs(7491) <= not a;
    layer7_outputs(7492) <= not b or a;
    layer7_outputs(7493) <= not b or a;
    layer7_outputs(7494) <= b;
    layer7_outputs(7495) <= a and not b;
    layer7_outputs(7496) <= not (a or b);
    layer7_outputs(7497) <= not a;
    layer7_outputs(7498) <= not b or a;
    layer7_outputs(7499) <= not a or b;
    layer7_outputs(7500) <= not a or b;
    layer7_outputs(7501) <= b and not a;
    layer7_outputs(7502) <= a or b;
    layer7_outputs(7503) <= a;
    layer7_outputs(7504) <= a or b;
    layer7_outputs(7505) <= not (a xor b);
    layer7_outputs(7506) <= a and b;
    layer7_outputs(7507) <= not a;
    layer7_outputs(7508) <= '0';
    layer7_outputs(7509) <= not (a and b);
    layer7_outputs(7510) <= a and b;
    layer7_outputs(7511) <= not a or b;
    layer7_outputs(7512) <= not b;
    layer7_outputs(7513) <= a xor b;
    layer7_outputs(7514) <= not b;
    layer7_outputs(7515) <= a and b;
    layer7_outputs(7516) <= not (a or b);
    layer7_outputs(7517) <= a or b;
    layer7_outputs(7518) <= not (a xor b);
    layer7_outputs(7519) <= not (a xor b);
    layer7_outputs(7520) <= a or b;
    layer7_outputs(7521) <= not b or a;
    layer7_outputs(7522) <= not a or b;
    layer7_outputs(7523) <= not a or b;
    layer7_outputs(7524) <= not (a and b);
    layer7_outputs(7525) <= a;
    layer7_outputs(7526) <= a xor b;
    layer7_outputs(7527) <= b;
    layer7_outputs(7528) <= not a;
    layer7_outputs(7529) <= b;
    layer7_outputs(7530) <= not a;
    layer7_outputs(7531) <= not a or b;
    layer7_outputs(7532) <= a xor b;
    layer7_outputs(7533) <= b and not a;
    layer7_outputs(7534) <= not b or a;
    layer7_outputs(7535) <= not (a xor b);
    layer7_outputs(7536) <= a and b;
    layer7_outputs(7537) <= not b;
    layer7_outputs(7538) <= not (a xor b);
    layer7_outputs(7539) <= not a or b;
    layer7_outputs(7540) <= a;
    layer7_outputs(7541) <= not a or b;
    layer7_outputs(7542) <= not b;
    layer7_outputs(7543) <= not (a and b);
    layer7_outputs(7544) <= not b or a;
    layer7_outputs(7545) <= not (a or b);
    layer7_outputs(7546) <= not a;
    layer7_outputs(7547) <= not b;
    layer7_outputs(7548) <= not (a and b);
    layer7_outputs(7549) <= b;
    layer7_outputs(7550) <= b;
    layer7_outputs(7551) <= b and not a;
    layer7_outputs(7552) <= not a;
    layer7_outputs(7553) <= not (a and b);
    layer7_outputs(7554) <= a;
    layer7_outputs(7555) <= a or b;
    layer7_outputs(7556) <= b and not a;
    layer7_outputs(7557) <= a and not b;
    layer7_outputs(7558) <= a or b;
    layer7_outputs(7559) <= not (a and b);
    layer7_outputs(7560) <= not b or a;
    layer7_outputs(7561) <= a or b;
    layer7_outputs(7562) <= a;
    layer7_outputs(7563) <= not (a xor b);
    layer7_outputs(7564) <= not a or b;
    layer7_outputs(7565) <= b;
    layer7_outputs(7566) <= not (a and b);
    layer7_outputs(7567) <= a and b;
    layer7_outputs(7568) <= not a or b;
    layer7_outputs(7569) <= not (a and b);
    layer7_outputs(7570) <= not b;
    layer7_outputs(7571) <= b;
    layer7_outputs(7572) <= not (a and b);
    layer7_outputs(7573) <= not b;
    layer7_outputs(7574) <= a xor b;
    layer7_outputs(7575) <= not (a or b);
    layer7_outputs(7576) <= not b;
    layer7_outputs(7577) <= b;
    layer7_outputs(7578) <= not b;
    layer7_outputs(7579) <= not (a and b);
    layer7_outputs(7580) <= b;
    layer7_outputs(7581) <= a xor b;
    layer7_outputs(7582) <= not (a or b);
    layer7_outputs(7583) <= not a;
    layer7_outputs(7584) <= not b or a;
    layer7_outputs(7585) <= not b or a;
    layer7_outputs(7586) <= not (a or b);
    layer7_outputs(7587) <= a xor b;
    layer7_outputs(7588) <= b;
    layer7_outputs(7589) <= not a or b;
    layer7_outputs(7590) <= not a;
    layer7_outputs(7591) <= b;
    layer7_outputs(7592) <= a xor b;
    layer7_outputs(7593) <= a or b;
    layer7_outputs(7594) <= b;
    layer7_outputs(7595) <= not b;
    layer7_outputs(7596) <= not (a xor b);
    layer7_outputs(7597) <= not (a xor b);
    layer7_outputs(7598) <= b;
    layer7_outputs(7599) <= not b;
    layer7_outputs(7600) <= not a or b;
    layer7_outputs(7601) <= not a;
    layer7_outputs(7602) <= not b;
    layer7_outputs(7603) <= a;
    layer7_outputs(7604) <= a;
    layer7_outputs(7605) <= not b;
    layer7_outputs(7606) <= a;
    layer7_outputs(7607) <= a and b;
    layer7_outputs(7608) <= not a;
    layer7_outputs(7609) <= not (a or b);
    layer7_outputs(7610) <= '1';
    layer7_outputs(7611) <= not (a and b);
    layer7_outputs(7612) <= not (a and b);
    layer7_outputs(7613) <= a xor b;
    layer7_outputs(7614) <= a or b;
    layer7_outputs(7615) <= not a or b;
    layer7_outputs(7616) <= not (a xor b);
    layer7_outputs(7617) <= not b;
    layer7_outputs(7618) <= b;
    layer7_outputs(7619) <= a and not b;
    layer7_outputs(7620) <= a or b;
    layer7_outputs(7621) <= not (a or b);
    layer7_outputs(7622) <= not a or b;
    layer7_outputs(7623) <= a or b;
    layer7_outputs(7624) <= a;
    layer7_outputs(7625) <= not (a and b);
    layer7_outputs(7626) <= a and not b;
    layer7_outputs(7627) <= a;
    layer7_outputs(7628) <= a;
    layer7_outputs(7629) <= not (a xor b);
    layer7_outputs(7630) <= not (a and b);
    layer7_outputs(7631) <= b;
    layer7_outputs(7632) <= a and not b;
    layer7_outputs(7633) <= not b or a;
    layer7_outputs(7634) <= b and not a;
    layer7_outputs(7635) <= a;
    layer7_outputs(7636) <= not (a or b);
    layer7_outputs(7637) <= not b;
    layer7_outputs(7638) <= not (a and b);
    layer7_outputs(7639) <= not a or b;
    layer7_outputs(7640) <= not (a or b);
    layer7_outputs(7641) <= not (a and b);
    layer7_outputs(7642) <= not b;
    layer7_outputs(7643) <= not (a xor b);
    layer7_outputs(7644) <= a or b;
    layer7_outputs(7645) <= not a;
    layer7_outputs(7646) <= not (a or b);
    layer7_outputs(7647) <= b;
    layer7_outputs(7648) <= '0';
    layer7_outputs(7649) <= '1';
    layer7_outputs(7650) <= b and not a;
    layer7_outputs(7651) <= a and b;
    layer7_outputs(7652) <= not (a and b);
    layer7_outputs(7653) <= '1';
    layer7_outputs(7654) <= not (a and b);
    layer7_outputs(7655) <= a xor b;
    layer7_outputs(7656) <= not a;
    layer7_outputs(7657) <= not b;
    layer7_outputs(7658) <= a or b;
    layer7_outputs(7659) <= a;
    layer7_outputs(7660) <= a or b;
    layer7_outputs(7661) <= b and not a;
    layer7_outputs(7662) <= not a or b;
    layer7_outputs(7663) <= a and b;
    layer7_outputs(7664) <= not (a xor b);
    layer7_outputs(7665) <= a and b;
    layer7_outputs(7666) <= not b;
    layer7_outputs(7667) <= a xor b;
    layer7_outputs(7668) <= b;
    layer7_outputs(7669) <= a and not b;
    layer7_outputs(7670) <= not b or a;
    layer7_outputs(7671) <= not b;
    layer7_outputs(7672) <= not b;
    layer7_outputs(7673) <= not b or a;
    layer7_outputs(7674) <= not a;
    layer7_outputs(7675) <= not a;
    layer7_outputs(7676) <= b;
    layer7_outputs(7677) <= not a or b;
    layer7_outputs(7678) <= not b;
    layer7_outputs(7679) <= not a;
    layer8_outputs(0) <= b;
    layer8_outputs(1) <= not (a xor b);
    layer8_outputs(2) <= a;
    layer8_outputs(3) <= not (a xor b);
    layer8_outputs(4) <= a;
    layer8_outputs(5) <= a and b;
    layer8_outputs(6) <= not a or b;
    layer8_outputs(7) <= not a or b;
    layer8_outputs(8) <= a;
    layer8_outputs(9) <= not (a xor b);
    layer8_outputs(10) <= a and not b;
    layer8_outputs(11) <= not b;
    layer8_outputs(12) <= not (a or b);
    layer8_outputs(13) <= a;
    layer8_outputs(14) <= b;
    layer8_outputs(15) <= not (a xor b);
    layer8_outputs(16) <= not a or b;
    layer8_outputs(17) <= not b;
    layer8_outputs(18) <= not (a xor b);
    layer8_outputs(19) <= not (a xor b);
    layer8_outputs(20) <= b and not a;
    layer8_outputs(21) <= not a;
    layer8_outputs(22) <= not b or a;
    layer8_outputs(23) <= not b;
    layer8_outputs(24) <= not a;
    layer8_outputs(25) <= a;
    layer8_outputs(26) <= not a;
    layer8_outputs(27) <= not b;
    layer8_outputs(28) <= b;
    layer8_outputs(29) <= a and b;
    layer8_outputs(30) <= not (a or b);
    layer8_outputs(31) <= not (a or b);
    layer8_outputs(32) <= not (a and b);
    layer8_outputs(33) <= not b or a;
    layer8_outputs(34) <= a and not b;
    layer8_outputs(35) <= not (a or b);
    layer8_outputs(36) <= a xor b;
    layer8_outputs(37) <= not a;
    layer8_outputs(38) <= a;
    layer8_outputs(39) <= not b or a;
    layer8_outputs(40) <= a;
    layer8_outputs(41) <= not (a or b);
    layer8_outputs(42) <= a;
    layer8_outputs(43) <= not (a xor b);
    layer8_outputs(44) <= a and not b;
    layer8_outputs(45) <= not b or a;
    layer8_outputs(46) <= not b or a;
    layer8_outputs(47) <= not b;
    layer8_outputs(48) <= not (a xor b);
    layer8_outputs(49) <= a;
    layer8_outputs(50) <= b;
    layer8_outputs(51) <= a;
    layer8_outputs(52) <= b;
    layer8_outputs(53) <= b;
    layer8_outputs(54) <= b and not a;
    layer8_outputs(55) <= b;
    layer8_outputs(56) <= not a or b;
    layer8_outputs(57) <= b;
    layer8_outputs(58) <= a;
    layer8_outputs(59) <= not (a xor b);
    layer8_outputs(60) <= a;
    layer8_outputs(61) <= not a;
    layer8_outputs(62) <= a and not b;
    layer8_outputs(63) <= a xor b;
    layer8_outputs(64) <= not (a xor b);
    layer8_outputs(65) <= a;
    layer8_outputs(66) <= a and b;
    layer8_outputs(67) <= a xor b;
    layer8_outputs(68) <= a xor b;
    layer8_outputs(69) <= a xor b;
    layer8_outputs(70) <= a;
    layer8_outputs(71) <= not a;
    layer8_outputs(72) <= not (a or b);
    layer8_outputs(73) <= not (a xor b);
    layer8_outputs(74) <= a and not b;
    layer8_outputs(75) <= a xor b;
    layer8_outputs(76) <= not b;
    layer8_outputs(77) <= b and not a;
    layer8_outputs(78) <= not a or b;
    layer8_outputs(79) <= b;
    layer8_outputs(80) <= not b;
    layer8_outputs(81) <= not a;
    layer8_outputs(82) <= not (a and b);
    layer8_outputs(83) <= b;
    layer8_outputs(84) <= not a;
    layer8_outputs(85) <= b;
    layer8_outputs(86) <= a or b;
    layer8_outputs(87) <= a and not b;
    layer8_outputs(88) <= a xor b;
    layer8_outputs(89) <= b;
    layer8_outputs(90) <= '0';
    layer8_outputs(91) <= a and b;
    layer8_outputs(92) <= not a;
    layer8_outputs(93) <= a or b;
    layer8_outputs(94) <= a xor b;
    layer8_outputs(95) <= a xor b;
    layer8_outputs(96) <= not b;
    layer8_outputs(97) <= b;
    layer8_outputs(98) <= not b;
    layer8_outputs(99) <= a xor b;
    layer8_outputs(100) <= not a;
    layer8_outputs(101) <= not a;
    layer8_outputs(102) <= not (a xor b);
    layer8_outputs(103) <= not b;
    layer8_outputs(104) <= not b;
    layer8_outputs(105) <= not a;
    layer8_outputs(106) <= not b;
    layer8_outputs(107) <= not b;
    layer8_outputs(108) <= b;
    layer8_outputs(109) <= a;
    layer8_outputs(110) <= not (a xor b);
    layer8_outputs(111) <= not (a or b);
    layer8_outputs(112) <= a;
    layer8_outputs(113) <= a and not b;
    layer8_outputs(114) <= not (a or b);
    layer8_outputs(115) <= not (a xor b);
    layer8_outputs(116) <= not (a and b);
    layer8_outputs(117) <= not (a xor b);
    layer8_outputs(118) <= a and b;
    layer8_outputs(119) <= not b;
    layer8_outputs(120) <= not (a and b);
    layer8_outputs(121) <= not b or a;
    layer8_outputs(122) <= b and not a;
    layer8_outputs(123) <= not b or a;
    layer8_outputs(124) <= not a;
    layer8_outputs(125) <= a;
    layer8_outputs(126) <= b;
    layer8_outputs(127) <= a xor b;
    layer8_outputs(128) <= a xor b;
    layer8_outputs(129) <= not a or b;
    layer8_outputs(130) <= not (a and b);
    layer8_outputs(131) <= b and not a;
    layer8_outputs(132) <= b;
    layer8_outputs(133) <= b;
    layer8_outputs(134) <= a;
    layer8_outputs(135) <= not (a and b);
    layer8_outputs(136) <= not a;
    layer8_outputs(137) <= b and not a;
    layer8_outputs(138) <= not a or b;
    layer8_outputs(139) <= a;
    layer8_outputs(140) <= a or b;
    layer8_outputs(141) <= a and b;
    layer8_outputs(142) <= not (a xor b);
    layer8_outputs(143) <= a;
    layer8_outputs(144) <= not (a or b);
    layer8_outputs(145) <= not b or a;
    layer8_outputs(146) <= b;
    layer8_outputs(147) <= b;
    layer8_outputs(148) <= a xor b;
    layer8_outputs(149) <= b;
    layer8_outputs(150) <= not (a xor b);
    layer8_outputs(151) <= not (a xor b);
    layer8_outputs(152) <= a xor b;
    layer8_outputs(153) <= not (a and b);
    layer8_outputs(154) <= a xor b;
    layer8_outputs(155) <= b;
    layer8_outputs(156) <= not (a and b);
    layer8_outputs(157) <= b and not a;
    layer8_outputs(158) <= a xor b;
    layer8_outputs(159) <= b;
    layer8_outputs(160) <= a and b;
    layer8_outputs(161) <= a;
    layer8_outputs(162) <= a xor b;
    layer8_outputs(163) <= a xor b;
    layer8_outputs(164) <= b;
    layer8_outputs(165) <= a;
    layer8_outputs(166) <= b and not a;
    layer8_outputs(167) <= a;
    layer8_outputs(168) <= b and not a;
    layer8_outputs(169) <= b;
    layer8_outputs(170) <= b;
    layer8_outputs(171) <= not a;
    layer8_outputs(172) <= a or b;
    layer8_outputs(173) <= a;
    layer8_outputs(174) <= a;
    layer8_outputs(175) <= a;
    layer8_outputs(176) <= a;
    layer8_outputs(177) <= not (a xor b);
    layer8_outputs(178) <= a xor b;
    layer8_outputs(179) <= not a;
    layer8_outputs(180) <= not (a or b);
    layer8_outputs(181) <= not a or b;
    layer8_outputs(182) <= a or b;
    layer8_outputs(183) <= b;
    layer8_outputs(184) <= '1';
    layer8_outputs(185) <= b;
    layer8_outputs(186) <= not (a and b);
    layer8_outputs(187) <= b and not a;
    layer8_outputs(188) <= b;
    layer8_outputs(189) <= not (a xor b);
    layer8_outputs(190) <= not b;
    layer8_outputs(191) <= a and not b;
    layer8_outputs(192) <= not a;
    layer8_outputs(193) <= a;
    layer8_outputs(194) <= a and not b;
    layer8_outputs(195) <= not b;
    layer8_outputs(196) <= not (a xor b);
    layer8_outputs(197) <= a and b;
    layer8_outputs(198) <= b;
    layer8_outputs(199) <= not a or b;
    layer8_outputs(200) <= not (a or b);
    layer8_outputs(201) <= a;
    layer8_outputs(202) <= not a;
    layer8_outputs(203) <= not a;
    layer8_outputs(204) <= not (a xor b);
    layer8_outputs(205) <= b and not a;
    layer8_outputs(206) <= a xor b;
    layer8_outputs(207) <= not a;
    layer8_outputs(208) <= not a;
    layer8_outputs(209) <= not b or a;
    layer8_outputs(210) <= not a;
    layer8_outputs(211) <= a;
    layer8_outputs(212) <= a xor b;
    layer8_outputs(213) <= not (a xor b);
    layer8_outputs(214) <= not a;
    layer8_outputs(215) <= not a;
    layer8_outputs(216) <= a;
    layer8_outputs(217) <= not b;
    layer8_outputs(218) <= not (a and b);
    layer8_outputs(219) <= b;
    layer8_outputs(220) <= not (a and b);
    layer8_outputs(221) <= not b or a;
    layer8_outputs(222) <= a or b;
    layer8_outputs(223) <= not (a and b);
    layer8_outputs(224) <= not (a xor b);
    layer8_outputs(225) <= not a;
    layer8_outputs(226) <= a and not b;
    layer8_outputs(227) <= a;
    layer8_outputs(228) <= not b or a;
    layer8_outputs(229) <= not (a xor b);
    layer8_outputs(230) <= b;
    layer8_outputs(231) <= not b;
    layer8_outputs(232) <= not (a or b);
    layer8_outputs(233) <= a;
    layer8_outputs(234) <= a xor b;
    layer8_outputs(235) <= not a;
    layer8_outputs(236) <= not (a xor b);
    layer8_outputs(237) <= a;
    layer8_outputs(238) <= not (a or b);
    layer8_outputs(239) <= a;
    layer8_outputs(240) <= not b;
    layer8_outputs(241) <= a and b;
    layer8_outputs(242) <= not a;
    layer8_outputs(243) <= a or b;
    layer8_outputs(244) <= not b;
    layer8_outputs(245) <= not b or a;
    layer8_outputs(246) <= b;
    layer8_outputs(247) <= not (a xor b);
    layer8_outputs(248) <= b;
    layer8_outputs(249) <= a and not b;
    layer8_outputs(250) <= b;
    layer8_outputs(251) <= b;
    layer8_outputs(252) <= not (a or b);
    layer8_outputs(253) <= a;
    layer8_outputs(254) <= not a;
    layer8_outputs(255) <= a or b;
    layer8_outputs(256) <= not (a xor b);
    layer8_outputs(257) <= not b;
    layer8_outputs(258) <= a and b;
    layer8_outputs(259) <= a;
    layer8_outputs(260) <= not a;
    layer8_outputs(261) <= a;
    layer8_outputs(262) <= a;
    layer8_outputs(263) <= b;
    layer8_outputs(264) <= not a;
    layer8_outputs(265) <= b;
    layer8_outputs(266) <= not b;
    layer8_outputs(267) <= a;
    layer8_outputs(268) <= a and not b;
    layer8_outputs(269) <= not (a or b);
    layer8_outputs(270) <= not (a xor b);
    layer8_outputs(271) <= not b;
    layer8_outputs(272) <= '1';
    layer8_outputs(273) <= b;
    layer8_outputs(274) <= a xor b;
    layer8_outputs(275) <= not b;
    layer8_outputs(276) <= a;
    layer8_outputs(277) <= not a or b;
    layer8_outputs(278) <= b;
    layer8_outputs(279) <= not (a xor b);
    layer8_outputs(280) <= not a;
    layer8_outputs(281) <= a;
    layer8_outputs(282) <= b and not a;
    layer8_outputs(283) <= b;
    layer8_outputs(284) <= not (a and b);
    layer8_outputs(285) <= b;
    layer8_outputs(286) <= not (a and b);
    layer8_outputs(287) <= not a or b;
    layer8_outputs(288) <= a;
    layer8_outputs(289) <= not (a xor b);
    layer8_outputs(290) <= a;
    layer8_outputs(291) <= a or b;
    layer8_outputs(292) <= not a;
    layer8_outputs(293) <= a xor b;
    layer8_outputs(294) <= b and not a;
    layer8_outputs(295) <= not a;
    layer8_outputs(296) <= not b or a;
    layer8_outputs(297) <= '1';
    layer8_outputs(298) <= a xor b;
    layer8_outputs(299) <= b and not a;
    layer8_outputs(300) <= b and not a;
    layer8_outputs(301) <= not b;
    layer8_outputs(302) <= a or b;
    layer8_outputs(303) <= b and not a;
    layer8_outputs(304) <= not b;
    layer8_outputs(305) <= not a or b;
    layer8_outputs(306) <= a;
    layer8_outputs(307) <= not b or a;
    layer8_outputs(308) <= not a;
    layer8_outputs(309) <= not b or a;
    layer8_outputs(310) <= a xor b;
    layer8_outputs(311) <= not a;
    layer8_outputs(312) <= not a;
    layer8_outputs(313) <= not a;
    layer8_outputs(314) <= a;
    layer8_outputs(315) <= not a or b;
    layer8_outputs(316) <= a;
    layer8_outputs(317) <= a and b;
    layer8_outputs(318) <= b and not a;
    layer8_outputs(319) <= b;
    layer8_outputs(320) <= not (a xor b);
    layer8_outputs(321) <= b;
    layer8_outputs(322) <= a;
    layer8_outputs(323) <= b and not a;
    layer8_outputs(324) <= a and not b;
    layer8_outputs(325) <= a xor b;
    layer8_outputs(326) <= a xor b;
    layer8_outputs(327) <= b;
    layer8_outputs(328) <= a xor b;
    layer8_outputs(329) <= not a;
    layer8_outputs(330) <= a xor b;
    layer8_outputs(331) <= not b;
    layer8_outputs(332) <= b and not a;
    layer8_outputs(333) <= b;
    layer8_outputs(334) <= a xor b;
    layer8_outputs(335) <= a xor b;
    layer8_outputs(336) <= a and not b;
    layer8_outputs(337) <= not (a xor b);
    layer8_outputs(338) <= a and b;
    layer8_outputs(339) <= b;
    layer8_outputs(340) <= not (a or b);
    layer8_outputs(341) <= a xor b;
    layer8_outputs(342) <= b;
    layer8_outputs(343) <= not b;
    layer8_outputs(344) <= not b or a;
    layer8_outputs(345) <= a and not b;
    layer8_outputs(346) <= not b or a;
    layer8_outputs(347) <= not (a xor b);
    layer8_outputs(348) <= b and not a;
    layer8_outputs(349) <= '1';
    layer8_outputs(350) <= a xor b;
    layer8_outputs(351) <= a or b;
    layer8_outputs(352) <= b;
    layer8_outputs(353) <= b and not a;
    layer8_outputs(354) <= not b;
    layer8_outputs(355) <= a and b;
    layer8_outputs(356) <= not (a xor b);
    layer8_outputs(357) <= b;
    layer8_outputs(358) <= a and b;
    layer8_outputs(359) <= not a;
    layer8_outputs(360) <= not (a or b);
    layer8_outputs(361) <= b and not a;
    layer8_outputs(362) <= a xor b;
    layer8_outputs(363) <= not a;
    layer8_outputs(364) <= not (a or b);
    layer8_outputs(365) <= not (a xor b);
    layer8_outputs(366) <= a xor b;
    layer8_outputs(367) <= a;
    layer8_outputs(368) <= not (a xor b);
    layer8_outputs(369) <= not (a or b);
    layer8_outputs(370) <= b;
    layer8_outputs(371) <= b;
    layer8_outputs(372) <= a;
    layer8_outputs(373) <= not (a xor b);
    layer8_outputs(374) <= a and not b;
    layer8_outputs(375) <= not b;
    layer8_outputs(376) <= b and not a;
    layer8_outputs(377) <= a xor b;
    layer8_outputs(378) <= not (a xor b);
    layer8_outputs(379) <= a or b;
    layer8_outputs(380) <= not (a xor b);
    layer8_outputs(381) <= not b;
    layer8_outputs(382) <= a or b;
    layer8_outputs(383) <= not a or b;
    layer8_outputs(384) <= not a;
    layer8_outputs(385) <= a xor b;
    layer8_outputs(386) <= b;
    layer8_outputs(387) <= a;
    layer8_outputs(388) <= a xor b;
    layer8_outputs(389) <= not (a and b);
    layer8_outputs(390) <= b;
    layer8_outputs(391) <= not b or a;
    layer8_outputs(392) <= a xor b;
    layer8_outputs(393) <= not b;
    layer8_outputs(394) <= not b;
    layer8_outputs(395) <= a;
    layer8_outputs(396) <= a xor b;
    layer8_outputs(397) <= not (a xor b);
    layer8_outputs(398) <= b;
    layer8_outputs(399) <= not b or a;
    layer8_outputs(400) <= not b or a;
    layer8_outputs(401) <= not a;
    layer8_outputs(402) <= b and not a;
    layer8_outputs(403) <= a;
    layer8_outputs(404) <= not a;
    layer8_outputs(405) <= b and not a;
    layer8_outputs(406) <= not (a and b);
    layer8_outputs(407) <= not a or b;
    layer8_outputs(408) <= a or b;
    layer8_outputs(409) <= not (a or b);
    layer8_outputs(410) <= not a or b;
    layer8_outputs(411) <= b and not a;
    layer8_outputs(412) <= b;
    layer8_outputs(413) <= b;
    layer8_outputs(414) <= a;
    layer8_outputs(415) <= a;
    layer8_outputs(416) <= a or b;
    layer8_outputs(417) <= a xor b;
    layer8_outputs(418) <= '0';
    layer8_outputs(419) <= b and not a;
    layer8_outputs(420) <= b and not a;
    layer8_outputs(421) <= a and not b;
    layer8_outputs(422) <= a xor b;
    layer8_outputs(423) <= a and not b;
    layer8_outputs(424) <= not b;
    layer8_outputs(425) <= not b;
    layer8_outputs(426) <= a and b;
    layer8_outputs(427) <= a;
    layer8_outputs(428) <= not (a xor b);
    layer8_outputs(429) <= b;
    layer8_outputs(430) <= not a or b;
    layer8_outputs(431) <= b;
    layer8_outputs(432) <= not b or a;
    layer8_outputs(433) <= not (a xor b);
    layer8_outputs(434) <= a;
    layer8_outputs(435) <= a and b;
    layer8_outputs(436) <= b and not a;
    layer8_outputs(437) <= a;
    layer8_outputs(438) <= a;
    layer8_outputs(439) <= not (a or b);
    layer8_outputs(440) <= not a;
    layer8_outputs(441) <= not (a xor b);
    layer8_outputs(442) <= not b or a;
    layer8_outputs(443) <= not a;
    layer8_outputs(444) <= a xor b;
    layer8_outputs(445) <= a;
    layer8_outputs(446) <= b;
    layer8_outputs(447) <= not (a or b);
    layer8_outputs(448) <= not a;
    layer8_outputs(449) <= not a;
    layer8_outputs(450) <= a xor b;
    layer8_outputs(451) <= not (a and b);
    layer8_outputs(452) <= not b or a;
    layer8_outputs(453) <= b;
    layer8_outputs(454) <= not b or a;
    layer8_outputs(455) <= not b;
    layer8_outputs(456) <= not (a or b);
    layer8_outputs(457) <= not a;
    layer8_outputs(458) <= not a or b;
    layer8_outputs(459) <= a xor b;
    layer8_outputs(460) <= b;
    layer8_outputs(461) <= b and not a;
    layer8_outputs(462) <= a;
    layer8_outputs(463) <= a or b;
    layer8_outputs(464) <= a and not b;
    layer8_outputs(465) <= b;
    layer8_outputs(466) <= not (a xor b);
    layer8_outputs(467) <= a xor b;
    layer8_outputs(468) <= a and not b;
    layer8_outputs(469) <= b;
    layer8_outputs(470) <= a;
    layer8_outputs(471) <= not b;
    layer8_outputs(472) <= a and not b;
    layer8_outputs(473) <= not a;
    layer8_outputs(474) <= not (a xor b);
    layer8_outputs(475) <= a and not b;
    layer8_outputs(476) <= b and not a;
    layer8_outputs(477) <= not (a or b);
    layer8_outputs(478) <= not (a and b);
    layer8_outputs(479) <= a;
    layer8_outputs(480) <= not a;
    layer8_outputs(481) <= not (a or b);
    layer8_outputs(482) <= not a;
    layer8_outputs(483) <= not (a xor b);
    layer8_outputs(484) <= not (a or b);
    layer8_outputs(485) <= not (a xor b);
    layer8_outputs(486) <= a xor b;
    layer8_outputs(487) <= not (a xor b);
    layer8_outputs(488) <= b;
    layer8_outputs(489) <= not (a xor b);
    layer8_outputs(490) <= b;
    layer8_outputs(491) <= not b;
    layer8_outputs(492) <= not (a xor b);
    layer8_outputs(493) <= not b;
    layer8_outputs(494) <= not a;
    layer8_outputs(495) <= not b;
    layer8_outputs(496) <= not a;
    layer8_outputs(497) <= b;
    layer8_outputs(498) <= a;
    layer8_outputs(499) <= b and not a;
    layer8_outputs(500) <= not a;
    layer8_outputs(501) <= not a;
    layer8_outputs(502) <= a xor b;
    layer8_outputs(503) <= not b;
    layer8_outputs(504) <= '0';
    layer8_outputs(505) <= b;
    layer8_outputs(506) <= not (a xor b);
    layer8_outputs(507) <= a;
    layer8_outputs(508) <= a;
    layer8_outputs(509) <= a and b;
    layer8_outputs(510) <= not (a xor b);
    layer8_outputs(511) <= a xor b;
    layer8_outputs(512) <= a and b;
    layer8_outputs(513) <= not (a xor b);
    layer8_outputs(514) <= a and not b;
    layer8_outputs(515) <= not a;
    layer8_outputs(516) <= not b;
    layer8_outputs(517) <= not b or a;
    layer8_outputs(518) <= a or b;
    layer8_outputs(519) <= a and not b;
    layer8_outputs(520) <= not b;
    layer8_outputs(521) <= a xor b;
    layer8_outputs(522) <= b;
    layer8_outputs(523) <= a and not b;
    layer8_outputs(524) <= not a or b;
    layer8_outputs(525) <= b;
    layer8_outputs(526) <= b;
    layer8_outputs(527) <= not (a or b);
    layer8_outputs(528) <= not (a xor b);
    layer8_outputs(529) <= not (a and b);
    layer8_outputs(530) <= not (a and b);
    layer8_outputs(531) <= b;
    layer8_outputs(532) <= not (a xor b);
    layer8_outputs(533) <= a or b;
    layer8_outputs(534) <= not (a and b);
    layer8_outputs(535) <= not b;
    layer8_outputs(536) <= b;
    layer8_outputs(537) <= not b or a;
    layer8_outputs(538) <= not a;
    layer8_outputs(539) <= a and b;
    layer8_outputs(540) <= a xor b;
    layer8_outputs(541) <= not a or b;
    layer8_outputs(542) <= b;
    layer8_outputs(543) <= a xor b;
    layer8_outputs(544) <= b;
    layer8_outputs(545) <= a xor b;
    layer8_outputs(546) <= not (a xor b);
    layer8_outputs(547) <= not a;
    layer8_outputs(548) <= not b;
    layer8_outputs(549) <= a xor b;
    layer8_outputs(550) <= a;
    layer8_outputs(551) <= a xor b;
    layer8_outputs(552) <= b and not a;
    layer8_outputs(553) <= a xor b;
    layer8_outputs(554) <= a;
    layer8_outputs(555) <= not (a xor b);
    layer8_outputs(556) <= not a or b;
    layer8_outputs(557) <= '0';
    layer8_outputs(558) <= b;
    layer8_outputs(559) <= not a or b;
    layer8_outputs(560) <= a xor b;
    layer8_outputs(561) <= not b;
    layer8_outputs(562) <= not a;
    layer8_outputs(563) <= not b;
    layer8_outputs(564) <= b;
    layer8_outputs(565) <= a and b;
    layer8_outputs(566) <= a;
    layer8_outputs(567) <= b and not a;
    layer8_outputs(568) <= a;
    layer8_outputs(569) <= a xor b;
    layer8_outputs(570) <= not b;
    layer8_outputs(571) <= b and not a;
    layer8_outputs(572) <= not b;
    layer8_outputs(573) <= a and b;
    layer8_outputs(574) <= a;
    layer8_outputs(575) <= not b;
    layer8_outputs(576) <= b;
    layer8_outputs(577) <= not a;
    layer8_outputs(578) <= not a;
    layer8_outputs(579) <= '0';
    layer8_outputs(580) <= not a;
    layer8_outputs(581) <= a or b;
    layer8_outputs(582) <= not b or a;
    layer8_outputs(583) <= not (a or b);
    layer8_outputs(584) <= not (a or b);
    layer8_outputs(585) <= not (a xor b);
    layer8_outputs(586) <= not (a xor b);
    layer8_outputs(587) <= not a;
    layer8_outputs(588) <= a xor b;
    layer8_outputs(589) <= not (a or b);
    layer8_outputs(590) <= not a;
    layer8_outputs(591) <= not a;
    layer8_outputs(592) <= b and not a;
    layer8_outputs(593) <= a;
    layer8_outputs(594) <= not a;
    layer8_outputs(595) <= b;
    layer8_outputs(596) <= not b;
    layer8_outputs(597) <= a xor b;
    layer8_outputs(598) <= not b;
    layer8_outputs(599) <= a xor b;
    layer8_outputs(600) <= not (a or b);
    layer8_outputs(601) <= not b or a;
    layer8_outputs(602) <= a and b;
    layer8_outputs(603) <= not b;
    layer8_outputs(604) <= not (a or b);
    layer8_outputs(605) <= not a;
    layer8_outputs(606) <= not b;
    layer8_outputs(607) <= not a;
    layer8_outputs(608) <= b;
    layer8_outputs(609) <= a xor b;
    layer8_outputs(610) <= a and b;
    layer8_outputs(611) <= not (a or b);
    layer8_outputs(612) <= not a;
    layer8_outputs(613) <= b;
    layer8_outputs(614) <= a and b;
    layer8_outputs(615) <= b;
    layer8_outputs(616) <= not (a and b);
    layer8_outputs(617) <= b;
    layer8_outputs(618) <= a;
    layer8_outputs(619) <= a xor b;
    layer8_outputs(620) <= not (a or b);
    layer8_outputs(621) <= not b or a;
    layer8_outputs(622) <= not b;
    layer8_outputs(623) <= not (a and b);
    layer8_outputs(624) <= not (a xor b);
    layer8_outputs(625) <= a and not b;
    layer8_outputs(626) <= not a;
    layer8_outputs(627) <= not a;
    layer8_outputs(628) <= not (a xor b);
    layer8_outputs(629) <= a or b;
    layer8_outputs(630) <= not (a and b);
    layer8_outputs(631) <= '0';
    layer8_outputs(632) <= not b;
    layer8_outputs(633) <= not (a xor b);
    layer8_outputs(634) <= a and b;
    layer8_outputs(635) <= a;
    layer8_outputs(636) <= not a or b;
    layer8_outputs(637) <= not a;
    layer8_outputs(638) <= a and not b;
    layer8_outputs(639) <= a xor b;
    layer8_outputs(640) <= not (a xor b);
    layer8_outputs(641) <= b;
    layer8_outputs(642) <= a xor b;
    layer8_outputs(643) <= not (a and b);
    layer8_outputs(644) <= b;
    layer8_outputs(645) <= b and not a;
    layer8_outputs(646) <= a;
    layer8_outputs(647) <= not b;
    layer8_outputs(648) <= not (a and b);
    layer8_outputs(649) <= not (a or b);
    layer8_outputs(650) <= a;
    layer8_outputs(651) <= not (a xor b);
    layer8_outputs(652) <= b;
    layer8_outputs(653) <= not (a xor b);
    layer8_outputs(654) <= not (a xor b);
    layer8_outputs(655) <= not (a xor b);
    layer8_outputs(656) <= not (a xor b);
    layer8_outputs(657) <= b;
    layer8_outputs(658) <= a xor b;
    layer8_outputs(659) <= not b;
    layer8_outputs(660) <= not (a and b);
    layer8_outputs(661) <= not a;
    layer8_outputs(662) <= not (a xor b);
    layer8_outputs(663) <= '1';
    layer8_outputs(664) <= b and not a;
    layer8_outputs(665) <= not a or b;
    layer8_outputs(666) <= a xor b;
    layer8_outputs(667) <= a;
    layer8_outputs(668) <= a;
    layer8_outputs(669) <= a xor b;
    layer8_outputs(670) <= not (a xor b);
    layer8_outputs(671) <= not (a and b);
    layer8_outputs(672) <= a xor b;
    layer8_outputs(673) <= a or b;
    layer8_outputs(674) <= a xor b;
    layer8_outputs(675) <= not b;
    layer8_outputs(676) <= a xor b;
    layer8_outputs(677) <= not a;
    layer8_outputs(678) <= b;
    layer8_outputs(679) <= b and not a;
    layer8_outputs(680) <= a xor b;
    layer8_outputs(681) <= a;
    layer8_outputs(682) <= b;
    layer8_outputs(683) <= a or b;
    layer8_outputs(684) <= a and b;
    layer8_outputs(685) <= b;
    layer8_outputs(686) <= not a or b;
    layer8_outputs(687) <= not b;
    layer8_outputs(688) <= b;
    layer8_outputs(689) <= b and not a;
    layer8_outputs(690) <= b;
    layer8_outputs(691) <= not a;
    layer8_outputs(692) <= '0';
    layer8_outputs(693) <= not a or b;
    layer8_outputs(694) <= not b;
    layer8_outputs(695) <= b;
    layer8_outputs(696) <= not b;
    layer8_outputs(697) <= not (a xor b);
    layer8_outputs(698) <= a;
    layer8_outputs(699) <= not (a and b);
    layer8_outputs(700) <= not b;
    layer8_outputs(701) <= not a or b;
    layer8_outputs(702) <= not b;
    layer8_outputs(703) <= not a;
    layer8_outputs(704) <= not (a and b);
    layer8_outputs(705) <= not b;
    layer8_outputs(706) <= b;
    layer8_outputs(707) <= b and not a;
    layer8_outputs(708) <= not (a or b);
    layer8_outputs(709) <= not (a xor b);
    layer8_outputs(710) <= not (a and b);
    layer8_outputs(711) <= not (a xor b);
    layer8_outputs(712) <= not a or b;
    layer8_outputs(713) <= not a;
    layer8_outputs(714) <= not (a or b);
    layer8_outputs(715) <= a xor b;
    layer8_outputs(716) <= a;
    layer8_outputs(717) <= b;
    layer8_outputs(718) <= not a;
    layer8_outputs(719) <= not b or a;
    layer8_outputs(720) <= not (a or b);
    layer8_outputs(721) <= a xor b;
    layer8_outputs(722) <= not b;
    layer8_outputs(723) <= b;
    layer8_outputs(724) <= b;
    layer8_outputs(725) <= a xor b;
    layer8_outputs(726) <= not (a and b);
    layer8_outputs(727) <= not b;
    layer8_outputs(728) <= '0';
    layer8_outputs(729) <= not b;
    layer8_outputs(730) <= not a or b;
    layer8_outputs(731) <= not a;
    layer8_outputs(732) <= b;
    layer8_outputs(733) <= not b;
    layer8_outputs(734) <= b;
    layer8_outputs(735) <= b and not a;
    layer8_outputs(736) <= a xor b;
    layer8_outputs(737) <= not b or a;
    layer8_outputs(738) <= a;
    layer8_outputs(739) <= a and b;
    layer8_outputs(740) <= a xor b;
    layer8_outputs(741) <= a or b;
    layer8_outputs(742) <= not a;
    layer8_outputs(743) <= b and not a;
    layer8_outputs(744) <= a;
    layer8_outputs(745) <= b;
    layer8_outputs(746) <= a;
    layer8_outputs(747) <= a xor b;
    layer8_outputs(748) <= not (a xor b);
    layer8_outputs(749) <= a and b;
    layer8_outputs(750) <= a and b;
    layer8_outputs(751) <= not b;
    layer8_outputs(752) <= not b or a;
    layer8_outputs(753) <= a;
    layer8_outputs(754) <= not a;
    layer8_outputs(755) <= a or b;
    layer8_outputs(756) <= not b;
    layer8_outputs(757) <= a;
    layer8_outputs(758) <= a xor b;
    layer8_outputs(759) <= a and not b;
    layer8_outputs(760) <= a;
    layer8_outputs(761) <= not (a or b);
    layer8_outputs(762) <= b and not a;
    layer8_outputs(763) <= a;
    layer8_outputs(764) <= '1';
    layer8_outputs(765) <= not (a xor b);
    layer8_outputs(766) <= not a;
    layer8_outputs(767) <= not (a and b);
    layer8_outputs(768) <= not a;
    layer8_outputs(769) <= b;
    layer8_outputs(770) <= b and not a;
    layer8_outputs(771) <= a;
    layer8_outputs(772) <= not a;
    layer8_outputs(773) <= b;
    layer8_outputs(774) <= a xor b;
    layer8_outputs(775) <= a or b;
    layer8_outputs(776) <= not a;
    layer8_outputs(777) <= a xor b;
    layer8_outputs(778) <= '0';
    layer8_outputs(779) <= a and not b;
    layer8_outputs(780) <= a and b;
    layer8_outputs(781) <= not (a xor b);
    layer8_outputs(782) <= a xor b;
    layer8_outputs(783) <= not b;
    layer8_outputs(784) <= not b;
    layer8_outputs(785) <= a;
    layer8_outputs(786) <= a;
    layer8_outputs(787) <= not b;
    layer8_outputs(788) <= not a;
    layer8_outputs(789) <= a or b;
    layer8_outputs(790) <= a;
    layer8_outputs(791) <= b;
    layer8_outputs(792) <= a or b;
    layer8_outputs(793) <= not (a xor b);
    layer8_outputs(794) <= a;
    layer8_outputs(795) <= a xor b;
    layer8_outputs(796) <= a xor b;
    layer8_outputs(797) <= not (a or b);
    layer8_outputs(798) <= b and not a;
    layer8_outputs(799) <= a or b;
    layer8_outputs(800) <= b;
    layer8_outputs(801) <= not a or b;
    layer8_outputs(802) <= not (a and b);
    layer8_outputs(803) <= a and b;
    layer8_outputs(804) <= not b or a;
    layer8_outputs(805) <= a and not b;
    layer8_outputs(806) <= b and not a;
    layer8_outputs(807) <= '0';
    layer8_outputs(808) <= a and not b;
    layer8_outputs(809) <= b and not a;
    layer8_outputs(810) <= not a or b;
    layer8_outputs(811) <= not b;
    layer8_outputs(812) <= a and b;
    layer8_outputs(813) <= a and b;
    layer8_outputs(814) <= a;
    layer8_outputs(815) <= a xor b;
    layer8_outputs(816) <= a and not b;
    layer8_outputs(817) <= not a;
    layer8_outputs(818) <= not (a or b);
    layer8_outputs(819) <= not b;
    layer8_outputs(820) <= b and not a;
    layer8_outputs(821) <= a or b;
    layer8_outputs(822) <= a xor b;
    layer8_outputs(823) <= '0';
    layer8_outputs(824) <= not b;
    layer8_outputs(825) <= not a;
    layer8_outputs(826) <= a;
    layer8_outputs(827) <= b and not a;
    layer8_outputs(828) <= b;
    layer8_outputs(829) <= a;
    layer8_outputs(830) <= not b;
    layer8_outputs(831) <= b and not a;
    layer8_outputs(832) <= b;
    layer8_outputs(833) <= not b;
    layer8_outputs(834) <= a;
    layer8_outputs(835) <= not (a xor b);
    layer8_outputs(836) <= b and not a;
    layer8_outputs(837) <= a and b;
    layer8_outputs(838) <= not b or a;
    layer8_outputs(839) <= a;
    layer8_outputs(840) <= a;
    layer8_outputs(841) <= not a or b;
    layer8_outputs(842) <= a;
    layer8_outputs(843) <= b;
    layer8_outputs(844) <= a and not b;
    layer8_outputs(845) <= a xor b;
    layer8_outputs(846) <= a and not b;
    layer8_outputs(847) <= b and not a;
    layer8_outputs(848) <= not (a or b);
    layer8_outputs(849) <= not b or a;
    layer8_outputs(850) <= a xor b;
    layer8_outputs(851) <= a xor b;
    layer8_outputs(852) <= not a or b;
    layer8_outputs(853) <= a xor b;
    layer8_outputs(854) <= a and not b;
    layer8_outputs(855) <= not (a xor b);
    layer8_outputs(856) <= a and not b;
    layer8_outputs(857) <= not b;
    layer8_outputs(858) <= not a;
    layer8_outputs(859) <= a;
    layer8_outputs(860) <= a;
    layer8_outputs(861) <= a;
    layer8_outputs(862) <= not (a xor b);
    layer8_outputs(863) <= not a;
    layer8_outputs(864) <= a and not b;
    layer8_outputs(865) <= a or b;
    layer8_outputs(866) <= not (a or b);
    layer8_outputs(867) <= not b;
    layer8_outputs(868) <= not b;
    layer8_outputs(869) <= a and not b;
    layer8_outputs(870) <= b and not a;
    layer8_outputs(871) <= a xor b;
    layer8_outputs(872) <= not a or b;
    layer8_outputs(873) <= not b;
    layer8_outputs(874) <= not b or a;
    layer8_outputs(875) <= b and not a;
    layer8_outputs(876) <= a xor b;
    layer8_outputs(877) <= a or b;
    layer8_outputs(878) <= not b or a;
    layer8_outputs(879) <= '0';
    layer8_outputs(880) <= not a;
    layer8_outputs(881) <= a xor b;
    layer8_outputs(882) <= a xor b;
    layer8_outputs(883) <= a and not b;
    layer8_outputs(884) <= a or b;
    layer8_outputs(885) <= a xor b;
    layer8_outputs(886) <= not a;
    layer8_outputs(887) <= not b or a;
    layer8_outputs(888) <= not b;
    layer8_outputs(889) <= not (a xor b);
    layer8_outputs(890) <= not a;
    layer8_outputs(891) <= not b;
    layer8_outputs(892) <= '1';
    layer8_outputs(893) <= a and b;
    layer8_outputs(894) <= not b;
    layer8_outputs(895) <= not (a and b);
    layer8_outputs(896) <= not a;
    layer8_outputs(897) <= b and not a;
    layer8_outputs(898) <= a xor b;
    layer8_outputs(899) <= a;
    layer8_outputs(900) <= a and b;
    layer8_outputs(901) <= '1';
    layer8_outputs(902) <= not a;
    layer8_outputs(903) <= not (a and b);
    layer8_outputs(904) <= not a or b;
    layer8_outputs(905) <= not b;
    layer8_outputs(906) <= not a or b;
    layer8_outputs(907) <= a xor b;
    layer8_outputs(908) <= not b;
    layer8_outputs(909) <= not (a and b);
    layer8_outputs(910) <= not (a or b);
    layer8_outputs(911) <= not a;
    layer8_outputs(912) <= a xor b;
    layer8_outputs(913) <= a;
    layer8_outputs(914) <= a;
    layer8_outputs(915) <= a or b;
    layer8_outputs(916) <= not a;
    layer8_outputs(917) <= not (a xor b);
    layer8_outputs(918) <= b;
    layer8_outputs(919) <= b and not a;
    layer8_outputs(920) <= a;
    layer8_outputs(921) <= b and not a;
    layer8_outputs(922) <= not a;
    layer8_outputs(923) <= not b;
    layer8_outputs(924) <= b;
    layer8_outputs(925) <= not a;
    layer8_outputs(926) <= b;
    layer8_outputs(927) <= not b or a;
    layer8_outputs(928) <= b and not a;
    layer8_outputs(929) <= b;
    layer8_outputs(930) <= not a or b;
    layer8_outputs(931) <= a xor b;
    layer8_outputs(932) <= not a;
    layer8_outputs(933) <= a;
    layer8_outputs(934) <= a xor b;
    layer8_outputs(935) <= a xor b;
    layer8_outputs(936) <= not b;
    layer8_outputs(937) <= a;
    layer8_outputs(938) <= not b;
    layer8_outputs(939) <= not b;
    layer8_outputs(940) <= a xor b;
    layer8_outputs(941) <= a xor b;
    layer8_outputs(942) <= not (a and b);
    layer8_outputs(943) <= a or b;
    layer8_outputs(944) <= not a or b;
    layer8_outputs(945) <= not b;
    layer8_outputs(946) <= not a;
    layer8_outputs(947) <= not b;
    layer8_outputs(948) <= b;
    layer8_outputs(949) <= a and b;
    layer8_outputs(950) <= not (a xor b);
    layer8_outputs(951) <= not a;
    layer8_outputs(952) <= not b;
    layer8_outputs(953) <= not b;
    layer8_outputs(954) <= a xor b;
    layer8_outputs(955) <= not b or a;
    layer8_outputs(956) <= not (a and b);
    layer8_outputs(957) <= not (a xor b);
    layer8_outputs(958) <= not (a xor b);
    layer8_outputs(959) <= a;
    layer8_outputs(960) <= b;
    layer8_outputs(961) <= not b or a;
    layer8_outputs(962) <= not (a xor b);
    layer8_outputs(963) <= a and not b;
    layer8_outputs(964) <= a xor b;
    layer8_outputs(965) <= not (a and b);
    layer8_outputs(966) <= a xor b;
    layer8_outputs(967) <= not a;
    layer8_outputs(968) <= not b;
    layer8_outputs(969) <= not b;
    layer8_outputs(970) <= not a;
    layer8_outputs(971) <= b and not a;
    layer8_outputs(972) <= a;
    layer8_outputs(973) <= a;
    layer8_outputs(974) <= not b or a;
    layer8_outputs(975) <= not a;
    layer8_outputs(976) <= not (a xor b);
    layer8_outputs(977) <= b;
    layer8_outputs(978) <= a xor b;
    layer8_outputs(979) <= b;
    layer8_outputs(980) <= not (a xor b);
    layer8_outputs(981) <= b;
    layer8_outputs(982) <= a xor b;
    layer8_outputs(983) <= a xor b;
    layer8_outputs(984) <= a;
    layer8_outputs(985) <= not (a or b);
    layer8_outputs(986) <= b and not a;
    layer8_outputs(987) <= not a or b;
    layer8_outputs(988) <= not (a or b);
    layer8_outputs(989) <= not a or b;
    layer8_outputs(990) <= b;
    layer8_outputs(991) <= not (a or b);
    layer8_outputs(992) <= not b;
    layer8_outputs(993) <= b;
    layer8_outputs(994) <= a xor b;
    layer8_outputs(995) <= a and not b;
    layer8_outputs(996) <= not a;
    layer8_outputs(997) <= a and not b;
    layer8_outputs(998) <= b;
    layer8_outputs(999) <= not a;
    layer8_outputs(1000) <= not a;
    layer8_outputs(1001) <= not (a and b);
    layer8_outputs(1002) <= b and not a;
    layer8_outputs(1003) <= a;
    layer8_outputs(1004) <= b;
    layer8_outputs(1005) <= a;
    layer8_outputs(1006) <= a xor b;
    layer8_outputs(1007) <= not (a xor b);
    layer8_outputs(1008) <= b;
    layer8_outputs(1009) <= not a;
    layer8_outputs(1010) <= not b or a;
    layer8_outputs(1011) <= b;
    layer8_outputs(1012) <= a xor b;
    layer8_outputs(1013) <= b and not a;
    layer8_outputs(1014) <= b;
    layer8_outputs(1015) <= '1';
    layer8_outputs(1016) <= not b;
    layer8_outputs(1017) <= not a or b;
    layer8_outputs(1018) <= a xor b;
    layer8_outputs(1019) <= not b;
    layer8_outputs(1020) <= not (a or b);
    layer8_outputs(1021) <= not b;
    layer8_outputs(1022) <= b;
    layer8_outputs(1023) <= not (a and b);
    layer8_outputs(1024) <= not a;
    layer8_outputs(1025) <= a;
    layer8_outputs(1026) <= not b;
    layer8_outputs(1027) <= not a;
    layer8_outputs(1028) <= b;
    layer8_outputs(1029) <= b;
    layer8_outputs(1030) <= a;
    layer8_outputs(1031) <= a xor b;
    layer8_outputs(1032) <= a;
    layer8_outputs(1033) <= not (a and b);
    layer8_outputs(1034) <= b;
    layer8_outputs(1035) <= not (a or b);
    layer8_outputs(1036) <= not b;
    layer8_outputs(1037) <= not a;
    layer8_outputs(1038) <= not (a xor b);
    layer8_outputs(1039) <= not (a or b);
    layer8_outputs(1040) <= b;
    layer8_outputs(1041) <= not b or a;
    layer8_outputs(1042) <= a and b;
    layer8_outputs(1043) <= a xor b;
    layer8_outputs(1044) <= a;
    layer8_outputs(1045) <= b;
    layer8_outputs(1046) <= not b;
    layer8_outputs(1047) <= not (a xor b);
    layer8_outputs(1048) <= b;
    layer8_outputs(1049) <= not b;
    layer8_outputs(1050) <= a;
    layer8_outputs(1051) <= a and b;
    layer8_outputs(1052) <= not (a xor b);
    layer8_outputs(1053) <= a and b;
    layer8_outputs(1054) <= not a;
    layer8_outputs(1055) <= not (a and b);
    layer8_outputs(1056) <= a and b;
    layer8_outputs(1057) <= not (a xor b);
    layer8_outputs(1058) <= a and b;
    layer8_outputs(1059) <= not b;
    layer8_outputs(1060) <= not b;
    layer8_outputs(1061) <= not (a xor b);
    layer8_outputs(1062) <= not (a or b);
    layer8_outputs(1063) <= a;
    layer8_outputs(1064) <= a xor b;
    layer8_outputs(1065) <= not a or b;
    layer8_outputs(1066) <= not (a xor b);
    layer8_outputs(1067) <= a and b;
    layer8_outputs(1068) <= a and b;
    layer8_outputs(1069) <= not (a or b);
    layer8_outputs(1070) <= b;
    layer8_outputs(1071) <= a;
    layer8_outputs(1072) <= not b;
    layer8_outputs(1073) <= a or b;
    layer8_outputs(1074) <= a;
    layer8_outputs(1075) <= a and not b;
    layer8_outputs(1076) <= b;
    layer8_outputs(1077) <= not b;
    layer8_outputs(1078) <= a or b;
    layer8_outputs(1079) <= a;
    layer8_outputs(1080) <= not a or b;
    layer8_outputs(1081) <= not b;
    layer8_outputs(1082) <= not b or a;
    layer8_outputs(1083) <= not a;
    layer8_outputs(1084) <= not b;
    layer8_outputs(1085) <= not b;
    layer8_outputs(1086) <= b;
    layer8_outputs(1087) <= not b;
    layer8_outputs(1088) <= not b;
    layer8_outputs(1089) <= not b;
    layer8_outputs(1090) <= not a;
    layer8_outputs(1091) <= a and b;
    layer8_outputs(1092) <= not b;
    layer8_outputs(1093) <= not (a or b);
    layer8_outputs(1094) <= not (a xor b);
    layer8_outputs(1095) <= not a;
    layer8_outputs(1096) <= b;
    layer8_outputs(1097) <= not b or a;
    layer8_outputs(1098) <= a and not b;
    layer8_outputs(1099) <= not (a xor b);
    layer8_outputs(1100) <= b and not a;
    layer8_outputs(1101) <= not (a xor b);
    layer8_outputs(1102) <= not b or a;
    layer8_outputs(1103) <= not (a and b);
    layer8_outputs(1104) <= a xor b;
    layer8_outputs(1105) <= not (a xor b);
    layer8_outputs(1106) <= b and not a;
    layer8_outputs(1107) <= b;
    layer8_outputs(1108) <= not (a or b);
    layer8_outputs(1109) <= a and b;
    layer8_outputs(1110) <= a and not b;
    layer8_outputs(1111) <= not a or b;
    layer8_outputs(1112) <= a;
    layer8_outputs(1113) <= not a;
    layer8_outputs(1114) <= not (a or b);
    layer8_outputs(1115) <= not a;
    layer8_outputs(1116) <= not b or a;
    layer8_outputs(1117) <= a xor b;
    layer8_outputs(1118) <= not (a xor b);
    layer8_outputs(1119) <= a or b;
    layer8_outputs(1120) <= not a;
    layer8_outputs(1121) <= a or b;
    layer8_outputs(1122) <= not a;
    layer8_outputs(1123) <= a xor b;
    layer8_outputs(1124) <= not (a or b);
    layer8_outputs(1125) <= not (a xor b);
    layer8_outputs(1126) <= b and not a;
    layer8_outputs(1127) <= a xor b;
    layer8_outputs(1128) <= not b;
    layer8_outputs(1129) <= a xor b;
    layer8_outputs(1130) <= not a;
    layer8_outputs(1131) <= not b;
    layer8_outputs(1132) <= a xor b;
    layer8_outputs(1133) <= b;
    layer8_outputs(1134) <= a;
    layer8_outputs(1135) <= a;
    layer8_outputs(1136) <= b;
    layer8_outputs(1137) <= a and b;
    layer8_outputs(1138) <= not (a and b);
    layer8_outputs(1139) <= not a or b;
    layer8_outputs(1140) <= not (a and b);
    layer8_outputs(1141) <= not a;
    layer8_outputs(1142) <= not a;
    layer8_outputs(1143) <= a and not b;
    layer8_outputs(1144) <= a;
    layer8_outputs(1145) <= not a or b;
    layer8_outputs(1146) <= a;
    layer8_outputs(1147) <= a and not b;
    layer8_outputs(1148) <= not (a or b);
    layer8_outputs(1149) <= a and not b;
    layer8_outputs(1150) <= not a;
    layer8_outputs(1151) <= a xor b;
    layer8_outputs(1152) <= a xor b;
    layer8_outputs(1153) <= not a;
    layer8_outputs(1154) <= a xor b;
    layer8_outputs(1155) <= a xor b;
    layer8_outputs(1156) <= not a or b;
    layer8_outputs(1157) <= not a;
    layer8_outputs(1158) <= a or b;
    layer8_outputs(1159) <= b;
    layer8_outputs(1160) <= not (a xor b);
    layer8_outputs(1161) <= not b or a;
    layer8_outputs(1162) <= a;
    layer8_outputs(1163) <= a xor b;
    layer8_outputs(1164) <= a;
    layer8_outputs(1165) <= a xor b;
    layer8_outputs(1166) <= a;
    layer8_outputs(1167) <= not a or b;
    layer8_outputs(1168) <= not b;
    layer8_outputs(1169) <= b and not a;
    layer8_outputs(1170) <= not (a xor b);
    layer8_outputs(1171) <= a and b;
    layer8_outputs(1172) <= not (a xor b);
    layer8_outputs(1173) <= a;
    layer8_outputs(1174) <= '1';
    layer8_outputs(1175) <= a and not b;
    layer8_outputs(1176) <= a and b;
    layer8_outputs(1177) <= not b;
    layer8_outputs(1178) <= not b;
    layer8_outputs(1179) <= not a or b;
    layer8_outputs(1180) <= b;
    layer8_outputs(1181) <= b;
    layer8_outputs(1182) <= not a;
    layer8_outputs(1183) <= '1';
    layer8_outputs(1184) <= not (a and b);
    layer8_outputs(1185) <= not a or b;
    layer8_outputs(1186) <= not (a and b);
    layer8_outputs(1187) <= not a or b;
    layer8_outputs(1188) <= not (a xor b);
    layer8_outputs(1189) <= b and not a;
    layer8_outputs(1190) <= a or b;
    layer8_outputs(1191) <= a;
    layer8_outputs(1192) <= a or b;
    layer8_outputs(1193) <= not (a xor b);
    layer8_outputs(1194) <= a and not b;
    layer8_outputs(1195) <= b;
    layer8_outputs(1196) <= not a or b;
    layer8_outputs(1197) <= not a;
    layer8_outputs(1198) <= not a;
    layer8_outputs(1199) <= not a;
    layer8_outputs(1200) <= not (a xor b);
    layer8_outputs(1201) <= a;
    layer8_outputs(1202) <= not a;
    layer8_outputs(1203) <= not b;
    layer8_outputs(1204) <= a;
    layer8_outputs(1205) <= b;
    layer8_outputs(1206) <= not (a xor b);
    layer8_outputs(1207) <= not (a xor b);
    layer8_outputs(1208) <= not a or b;
    layer8_outputs(1209) <= not (a xor b);
    layer8_outputs(1210) <= not a;
    layer8_outputs(1211) <= a xor b;
    layer8_outputs(1212) <= not b;
    layer8_outputs(1213) <= not b;
    layer8_outputs(1214) <= a;
    layer8_outputs(1215) <= b;
    layer8_outputs(1216) <= not (a xor b);
    layer8_outputs(1217) <= not a;
    layer8_outputs(1218) <= not b or a;
    layer8_outputs(1219) <= not a or b;
    layer8_outputs(1220) <= not (a xor b);
    layer8_outputs(1221) <= '1';
    layer8_outputs(1222) <= a xor b;
    layer8_outputs(1223) <= not (a or b);
    layer8_outputs(1224) <= a xor b;
    layer8_outputs(1225) <= not a or b;
    layer8_outputs(1226) <= not b;
    layer8_outputs(1227) <= a xor b;
    layer8_outputs(1228) <= not b;
    layer8_outputs(1229) <= a and b;
    layer8_outputs(1230) <= not (a or b);
    layer8_outputs(1231) <= a xor b;
    layer8_outputs(1232) <= b;
    layer8_outputs(1233) <= not a;
    layer8_outputs(1234) <= not a;
    layer8_outputs(1235) <= not (a and b);
    layer8_outputs(1236) <= not (a xor b);
    layer8_outputs(1237) <= not b;
    layer8_outputs(1238) <= not (a or b);
    layer8_outputs(1239) <= not (a and b);
    layer8_outputs(1240) <= a xor b;
    layer8_outputs(1241) <= not a or b;
    layer8_outputs(1242) <= b;
    layer8_outputs(1243) <= not b;
    layer8_outputs(1244) <= a and not b;
    layer8_outputs(1245) <= not a;
    layer8_outputs(1246) <= a xor b;
    layer8_outputs(1247) <= b;
    layer8_outputs(1248) <= not (a xor b);
    layer8_outputs(1249) <= a and not b;
    layer8_outputs(1250) <= a and not b;
    layer8_outputs(1251) <= b;
    layer8_outputs(1252) <= b and not a;
    layer8_outputs(1253) <= a or b;
    layer8_outputs(1254) <= a and b;
    layer8_outputs(1255) <= a and b;
    layer8_outputs(1256) <= a or b;
    layer8_outputs(1257) <= a and b;
    layer8_outputs(1258) <= not b;
    layer8_outputs(1259) <= not a;
    layer8_outputs(1260) <= a;
    layer8_outputs(1261) <= a or b;
    layer8_outputs(1262) <= not b;
    layer8_outputs(1263) <= not a;
    layer8_outputs(1264) <= not b;
    layer8_outputs(1265) <= b;
    layer8_outputs(1266) <= a xor b;
    layer8_outputs(1267) <= not b or a;
    layer8_outputs(1268) <= a xor b;
    layer8_outputs(1269) <= a;
    layer8_outputs(1270) <= a;
    layer8_outputs(1271) <= not a;
    layer8_outputs(1272) <= not a or b;
    layer8_outputs(1273) <= a;
    layer8_outputs(1274) <= a xor b;
    layer8_outputs(1275) <= a and not b;
    layer8_outputs(1276) <= a;
    layer8_outputs(1277) <= a xor b;
    layer8_outputs(1278) <= not a;
    layer8_outputs(1279) <= b;
    layer8_outputs(1280) <= not (a and b);
    layer8_outputs(1281) <= not b;
    layer8_outputs(1282) <= b;
    layer8_outputs(1283) <= not (a xor b);
    layer8_outputs(1284) <= a or b;
    layer8_outputs(1285) <= not (a or b);
    layer8_outputs(1286) <= b;
    layer8_outputs(1287) <= a;
    layer8_outputs(1288) <= a;
    layer8_outputs(1289) <= a;
    layer8_outputs(1290) <= not b;
    layer8_outputs(1291) <= not a;
    layer8_outputs(1292) <= a or b;
    layer8_outputs(1293) <= a xor b;
    layer8_outputs(1294) <= not a;
    layer8_outputs(1295) <= a;
    layer8_outputs(1296) <= a and b;
    layer8_outputs(1297) <= a and b;
    layer8_outputs(1298) <= b;
    layer8_outputs(1299) <= a xor b;
    layer8_outputs(1300) <= not (a xor b);
    layer8_outputs(1301) <= b and not a;
    layer8_outputs(1302) <= not a;
    layer8_outputs(1303) <= not b;
    layer8_outputs(1304) <= b;
    layer8_outputs(1305) <= not (a or b);
    layer8_outputs(1306) <= a or b;
    layer8_outputs(1307) <= b and not a;
    layer8_outputs(1308) <= not a;
    layer8_outputs(1309) <= not a;
    layer8_outputs(1310) <= b and not a;
    layer8_outputs(1311) <= a and b;
    layer8_outputs(1312) <= not (a xor b);
    layer8_outputs(1313) <= a and not b;
    layer8_outputs(1314) <= not (a xor b);
    layer8_outputs(1315) <= a xor b;
    layer8_outputs(1316) <= b and not a;
    layer8_outputs(1317) <= not (a xor b);
    layer8_outputs(1318) <= a;
    layer8_outputs(1319) <= a or b;
    layer8_outputs(1320) <= b and not a;
    layer8_outputs(1321) <= not a;
    layer8_outputs(1322) <= not a or b;
    layer8_outputs(1323) <= not b;
    layer8_outputs(1324) <= not (a and b);
    layer8_outputs(1325) <= b and not a;
    layer8_outputs(1326) <= not a;
    layer8_outputs(1327) <= a xor b;
    layer8_outputs(1328) <= not (a or b);
    layer8_outputs(1329) <= a and not b;
    layer8_outputs(1330) <= not b;
    layer8_outputs(1331) <= b;
    layer8_outputs(1332) <= a or b;
    layer8_outputs(1333) <= not a;
    layer8_outputs(1334) <= not (a xor b);
    layer8_outputs(1335) <= a xor b;
    layer8_outputs(1336) <= not (a xor b);
    layer8_outputs(1337) <= not (a and b);
    layer8_outputs(1338) <= not a or b;
    layer8_outputs(1339) <= not a;
    layer8_outputs(1340) <= a;
    layer8_outputs(1341) <= not a or b;
    layer8_outputs(1342) <= a xor b;
    layer8_outputs(1343) <= not (a xor b);
    layer8_outputs(1344) <= a;
    layer8_outputs(1345) <= a;
    layer8_outputs(1346) <= not a;
    layer8_outputs(1347) <= a;
    layer8_outputs(1348) <= a or b;
    layer8_outputs(1349) <= a xor b;
    layer8_outputs(1350) <= not (a xor b);
    layer8_outputs(1351) <= a xor b;
    layer8_outputs(1352) <= a or b;
    layer8_outputs(1353) <= not b or a;
    layer8_outputs(1354) <= not b;
    layer8_outputs(1355) <= not (a or b);
    layer8_outputs(1356) <= a and not b;
    layer8_outputs(1357) <= not b or a;
    layer8_outputs(1358) <= not b;
    layer8_outputs(1359) <= a or b;
    layer8_outputs(1360) <= a and b;
    layer8_outputs(1361) <= not b;
    layer8_outputs(1362) <= not b;
    layer8_outputs(1363) <= b and not a;
    layer8_outputs(1364) <= a xor b;
    layer8_outputs(1365) <= a xor b;
    layer8_outputs(1366) <= not b;
    layer8_outputs(1367) <= not b;
    layer8_outputs(1368) <= '1';
    layer8_outputs(1369) <= not a;
    layer8_outputs(1370) <= a;
    layer8_outputs(1371) <= not a or b;
    layer8_outputs(1372) <= not a;
    layer8_outputs(1373) <= not a or b;
    layer8_outputs(1374) <= not b;
    layer8_outputs(1375) <= a and b;
    layer8_outputs(1376) <= not b;
    layer8_outputs(1377) <= not b;
    layer8_outputs(1378) <= b;
    layer8_outputs(1379) <= not b;
    layer8_outputs(1380) <= not a;
    layer8_outputs(1381) <= not a;
    layer8_outputs(1382) <= not b;
    layer8_outputs(1383) <= a;
    layer8_outputs(1384) <= b;
    layer8_outputs(1385) <= b;
    layer8_outputs(1386) <= not (a or b);
    layer8_outputs(1387) <= b and not a;
    layer8_outputs(1388) <= not a or b;
    layer8_outputs(1389) <= not (a xor b);
    layer8_outputs(1390) <= not (a or b);
    layer8_outputs(1391) <= '0';
    layer8_outputs(1392) <= b;
    layer8_outputs(1393) <= b and not a;
    layer8_outputs(1394) <= not (a and b);
    layer8_outputs(1395) <= not a;
    layer8_outputs(1396) <= a or b;
    layer8_outputs(1397) <= a;
    layer8_outputs(1398) <= a;
    layer8_outputs(1399) <= a;
    layer8_outputs(1400) <= b;
    layer8_outputs(1401) <= a;
    layer8_outputs(1402) <= b;
    layer8_outputs(1403) <= not a;
    layer8_outputs(1404) <= a and not b;
    layer8_outputs(1405) <= not b;
    layer8_outputs(1406) <= a and not b;
    layer8_outputs(1407) <= a and not b;
    layer8_outputs(1408) <= not (a xor b);
    layer8_outputs(1409) <= not b;
    layer8_outputs(1410) <= '1';
    layer8_outputs(1411) <= not a;
    layer8_outputs(1412) <= not (a and b);
    layer8_outputs(1413) <= not (a and b);
    layer8_outputs(1414) <= not a or b;
    layer8_outputs(1415) <= not a or b;
    layer8_outputs(1416) <= not a;
    layer8_outputs(1417) <= a and not b;
    layer8_outputs(1418) <= not b;
    layer8_outputs(1419) <= a xor b;
    layer8_outputs(1420) <= a;
    layer8_outputs(1421) <= b;
    layer8_outputs(1422) <= a or b;
    layer8_outputs(1423) <= a;
    layer8_outputs(1424) <= not b or a;
    layer8_outputs(1425) <= not (a xor b);
    layer8_outputs(1426) <= b;
    layer8_outputs(1427) <= not a;
    layer8_outputs(1428) <= b;
    layer8_outputs(1429) <= not a or b;
    layer8_outputs(1430) <= not b;
    layer8_outputs(1431) <= not a;
    layer8_outputs(1432) <= a or b;
    layer8_outputs(1433) <= a xor b;
    layer8_outputs(1434) <= a or b;
    layer8_outputs(1435) <= a and not b;
    layer8_outputs(1436) <= not a or b;
    layer8_outputs(1437) <= not a;
    layer8_outputs(1438) <= a;
    layer8_outputs(1439) <= not a or b;
    layer8_outputs(1440) <= not a;
    layer8_outputs(1441) <= a xor b;
    layer8_outputs(1442) <= a xor b;
    layer8_outputs(1443) <= not (a or b);
    layer8_outputs(1444) <= a;
    layer8_outputs(1445) <= not (a xor b);
    layer8_outputs(1446) <= a;
    layer8_outputs(1447) <= a xor b;
    layer8_outputs(1448) <= not b;
    layer8_outputs(1449) <= a xor b;
    layer8_outputs(1450) <= b;
    layer8_outputs(1451) <= not (a xor b);
    layer8_outputs(1452) <= a;
    layer8_outputs(1453) <= '0';
    layer8_outputs(1454) <= a;
    layer8_outputs(1455) <= not (a and b);
    layer8_outputs(1456) <= b and not a;
    layer8_outputs(1457) <= b;
    layer8_outputs(1458) <= b;
    layer8_outputs(1459) <= not b;
    layer8_outputs(1460) <= not b;
    layer8_outputs(1461) <= a;
    layer8_outputs(1462) <= b and not a;
    layer8_outputs(1463) <= a xor b;
    layer8_outputs(1464) <= a;
    layer8_outputs(1465) <= not (a xor b);
    layer8_outputs(1466) <= not b;
    layer8_outputs(1467) <= a;
    layer8_outputs(1468) <= a or b;
    layer8_outputs(1469) <= b;
    layer8_outputs(1470) <= a and not b;
    layer8_outputs(1471) <= not (a and b);
    layer8_outputs(1472) <= not a;
    layer8_outputs(1473) <= not b;
    layer8_outputs(1474) <= b and not a;
    layer8_outputs(1475) <= b;
    layer8_outputs(1476) <= a;
    layer8_outputs(1477) <= a and b;
    layer8_outputs(1478) <= not a;
    layer8_outputs(1479) <= not b;
    layer8_outputs(1480) <= b;
    layer8_outputs(1481) <= not (a or b);
    layer8_outputs(1482) <= a xor b;
    layer8_outputs(1483) <= not b;
    layer8_outputs(1484) <= not (a or b);
    layer8_outputs(1485) <= a xor b;
    layer8_outputs(1486) <= not (a or b);
    layer8_outputs(1487) <= not (a xor b);
    layer8_outputs(1488) <= not a;
    layer8_outputs(1489) <= a and b;
    layer8_outputs(1490) <= a;
    layer8_outputs(1491) <= a xor b;
    layer8_outputs(1492) <= a xor b;
    layer8_outputs(1493) <= not (a xor b);
    layer8_outputs(1494) <= not a;
    layer8_outputs(1495) <= b and not a;
    layer8_outputs(1496) <= not a;
    layer8_outputs(1497) <= not a or b;
    layer8_outputs(1498) <= a and not b;
    layer8_outputs(1499) <= b and not a;
    layer8_outputs(1500) <= a;
    layer8_outputs(1501) <= not (a or b);
    layer8_outputs(1502) <= a or b;
    layer8_outputs(1503) <= not b;
    layer8_outputs(1504) <= a xor b;
    layer8_outputs(1505) <= a;
    layer8_outputs(1506) <= b;
    layer8_outputs(1507) <= not (a and b);
    layer8_outputs(1508) <= not (a xor b);
    layer8_outputs(1509) <= not a or b;
    layer8_outputs(1510) <= not b;
    layer8_outputs(1511) <= a and b;
    layer8_outputs(1512) <= not a;
    layer8_outputs(1513) <= not (a and b);
    layer8_outputs(1514) <= a or b;
    layer8_outputs(1515) <= a xor b;
    layer8_outputs(1516) <= not a;
    layer8_outputs(1517) <= not b or a;
    layer8_outputs(1518) <= not (a xor b);
    layer8_outputs(1519) <= a and not b;
    layer8_outputs(1520) <= not (a xor b);
    layer8_outputs(1521) <= a xor b;
    layer8_outputs(1522) <= not (a or b);
    layer8_outputs(1523) <= a;
    layer8_outputs(1524) <= not (a xor b);
    layer8_outputs(1525) <= not (a or b);
    layer8_outputs(1526) <= a;
    layer8_outputs(1527) <= a xor b;
    layer8_outputs(1528) <= not b or a;
    layer8_outputs(1529) <= not (a and b);
    layer8_outputs(1530) <= b and not a;
    layer8_outputs(1531) <= b;
    layer8_outputs(1532) <= not (a or b);
    layer8_outputs(1533) <= a and not b;
    layer8_outputs(1534) <= not (a xor b);
    layer8_outputs(1535) <= not b;
    layer8_outputs(1536) <= not a;
    layer8_outputs(1537) <= b;
    layer8_outputs(1538) <= a or b;
    layer8_outputs(1539) <= not (a or b);
    layer8_outputs(1540) <= not b;
    layer8_outputs(1541) <= not (a and b);
    layer8_outputs(1542) <= not a;
    layer8_outputs(1543) <= not b or a;
    layer8_outputs(1544) <= not (a xor b);
    layer8_outputs(1545) <= not b;
    layer8_outputs(1546) <= not (a xor b);
    layer8_outputs(1547) <= not (a xor b);
    layer8_outputs(1548) <= b;
    layer8_outputs(1549) <= a;
    layer8_outputs(1550) <= not b;
    layer8_outputs(1551) <= not b;
    layer8_outputs(1552) <= not a;
    layer8_outputs(1553) <= not a;
    layer8_outputs(1554) <= b;
    layer8_outputs(1555) <= b;
    layer8_outputs(1556) <= not (a or b);
    layer8_outputs(1557) <= a xor b;
    layer8_outputs(1558) <= a and b;
    layer8_outputs(1559) <= not a or b;
    layer8_outputs(1560) <= '0';
    layer8_outputs(1561) <= not (a xor b);
    layer8_outputs(1562) <= not a;
    layer8_outputs(1563) <= not a or b;
    layer8_outputs(1564) <= a;
    layer8_outputs(1565) <= not b or a;
    layer8_outputs(1566) <= not (a xor b);
    layer8_outputs(1567) <= not a or b;
    layer8_outputs(1568) <= b;
    layer8_outputs(1569) <= not (a xor b);
    layer8_outputs(1570) <= not a;
    layer8_outputs(1571) <= '1';
    layer8_outputs(1572) <= not (a or b);
    layer8_outputs(1573) <= not a;
    layer8_outputs(1574) <= not b;
    layer8_outputs(1575) <= a or b;
    layer8_outputs(1576) <= not (a and b);
    layer8_outputs(1577) <= a;
    layer8_outputs(1578) <= not a;
    layer8_outputs(1579) <= not b;
    layer8_outputs(1580) <= not (a and b);
    layer8_outputs(1581) <= not b or a;
    layer8_outputs(1582) <= a and not b;
    layer8_outputs(1583) <= b and not a;
    layer8_outputs(1584) <= a;
    layer8_outputs(1585) <= not b;
    layer8_outputs(1586) <= a or b;
    layer8_outputs(1587) <= not (a and b);
    layer8_outputs(1588) <= not a or b;
    layer8_outputs(1589) <= a or b;
    layer8_outputs(1590) <= not (a xor b);
    layer8_outputs(1591) <= a and b;
    layer8_outputs(1592) <= a and b;
    layer8_outputs(1593) <= a or b;
    layer8_outputs(1594) <= a and b;
    layer8_outputs(1595) <= not a;
    layer8_outputs(1596) <= a;
    layer8_outputs(1597) <= not a;
    layer8_outputs(1598) <= a xor b;
    layer8_outputs(1599) <= not b;
    layer8_outputs(1600) <= not (a or b);
    layer8_outputs(1601) <= not a;
    layer8_outputs(1602) <= not (a and b);
    layer8_outputs(1603) <= not a;
    layer8_outputs(1604) <= not a or b;
    layer8_outputs(1605) <= not (a or b);
    layer8_outputs(1606) <= not a or b;
    layer8_outputs(1607) <= b and not a;
    layer8_outputs(1608) <= not a or b;
    layer8_outputs(1609) <= b and not a;
    layer8_outputs(1610) <= a xor b;
    layer8_outputs(1611) <= not (a xor b);
    layer8_outputs(1612) <= not a;
    layer8_outputs(1613) <= not b;
    layer8_outputs(1614) <= a xor b;
    layer8_outputs(1615) <= a and not b;
    layer8_outputs(1616) <= not b or a;
    layer8_outputs(1617) <= a;
    layer8_outputs(1618) <= a;
    layer8_outputs(1619) <= a and b;
    layer8_outputs(1620) <= not b;
    layer8_outputs(1621) <= not a;
    layer8_outputs(1622) <= a and b;
    layer8_outputs(1623) <= a xor b;
    layer8_outputs(1624) <= b;
    layer8_outputs(1625) <= b;
    layer8_outputs(1626) <= b and not a;
    layer8_outputs(1627) <= not (a xor b);
    layer8_outputs(1628) <= not (a or b);
    layer8_outputs(1629) <= not (a or b);
    layer8_outputs(1630) <= not (a or b);
    layer8_outputs(1631) <= not a;
    layer8_outputs(1632) <= a xor b;
    layer8_outputs(1633) <= a or b;
    layer8_outputs(1634) <= not b;
    layer8_outputs(1635) <= b;
    layer8_outputs(1636) <= a;
    layer8_outputs(1637) <= a or b;
    layer8_outputs(1638) <= not (a and b);
    layer8_outputs(1639) <= a;
    layer8_outputs(1640) <= a;
    layer8_outputs(1641) <= a;
    layer8_outputs(1642) <= not a or b;
    layer8_outputs(1643) <= b;
    layer8_outputs(1644) <= not (a and b);
    layer8_outputs(1645) <= a;
    layer8_outputs(1646) <= a and not b;
    layer8_outputs(1647) <= not a or b;
    layer8_outputs(1648) <= a and not b;
    layer8_outputs(1649) <= a and b;
    layer8_outputs(1650) <= b;
    layer8_outputs(1651) <= a xor b;
    layer8_outputs(1652) <= a;
    layer8_outputs(1653) <= a or b;
    layer8_outputs(1654) <= a xor b;
    layer8_outputs(1655) <= a xor b;
    layer8_outputs(1656) <= b;
    layer8_outputs(1657) <= a;
    layer8_outputs(1658) <= a or b;
    layer8_outputs(1659) <= a or b;
    layer8_outputs(1660) <= not (a and b);
    layer8_outputs(1661) <= not (a xor b);
    layer8_outputs(1662) <= b;
    layer8_outputs(1663) <= not (a xor b);
    layer8_outputs(1664) <= a and b;
    layer8_outputs(1665) <= not a;
    layer8_outputs(1666) <= not (a xor b);
    layer8_outputs(1667) <= a and not b;
    layer8_outputs(1668) <= b;
    layer8_outputs(1669) <= not b;
    layer8_outputs(1670) <= not b;
    layer8_outputs(1671) <= not a;
    layer8_outputs(1672) <= not b or a;
    layer8_outputs(1673) <= not b or a;
    layer8_outputs(1674) <= not a;
    layer8_outputs(1675) <= a;
    layer8_outputs(1676) <= not a or b;
    layer8_outputs(1677) <= not b;
    layer8_outputs(1678) <= not a;
    layer8_outputs(1679) <= not (a xor b);
    layer8_outputs(1680) <= b;
    layer8_outputs(1681) <= a;
    layer8_outputs(1682) <= a and not b;
    layer8_outputs(1683) <= b and not a;
    layer8_outputs(1684) <= not a;
    layer8_outputs(1685) <= not (a and b);
    layer8_outputs(1686) <= not (a xor b);
    layer8_outputs(1687) <= not a;
    layer8_outputs(1688) <= a;
    layer8_outputs(1689) <= not (a xor b);
    layer8_outputs(1690) <= not a;
    layer8_outputs(1691) <= b;
    layer8_outputs(1692) <= a and not b;
    layer8_outputs(1693) <= a and b;
    layer8_outputs(1694) <= b;
    layer8_outputs(1695) <= a or b;
    layer8_outputs(1696) <= not b or a;
    layer8_outputs(1697) <= b;
    layer8_outputs(1698) <= b;
    layer8_outputs(1699) <= not b;
    layer8_outputs(1700) <= b and not a;
    layer8_outputs(1701) <= not (a or b);
    layer8_outputs(1702) <= a and b;
    layer8_outputs(1703) <= not a;
    layer8_outputs(1704) <= a;
    layer8_outputs(1705) <= not a or b;
    layer8_outputs(1706) <= a xor b;
    layer8_outputs(1707) <= a;
    layer8_outputs(1708) <= a xor b;
    layer8_outputs(1709) <= b and not a;
    layer8_outputs(1710) <= a or b;
    layer8_outputs(1711) <= a and b;
    layer8_outputs(1712) <= not (a and b);
    layer8_outputs(1713) <= not b;
    layer8_outputs(1714) <= a;
    layer8_outputs(1715) <= not b;
    layer8_outputs(1716) <= a xor b;
    layer8_outputs(1717) <= not a or b;
    layer8_outputs(1718) <= not (a xor b);
    layer8_outputs(1719) <= not a;
    layer8_outputs(1720) <= not (a or b);
    layer8_outputs(1721) <= not a;
    layer8_outputs(1722) <= a xor b;
    layer8_outputs(1723) <= not (a and b);
    layer8_outputs(1724) <= b;
    layer8_outputs(1725) <= not b or a;
    layer8_outputs(1726) <= a;
    layer8_outputs(1727) <= a xor b;
    layer8_outputs(1728) <= b;
    layer8_outputs(1729) <= b;
    layer8_outputs(1730) <= not (a xor b);
    layer8_outputs(1731) <= not a;
    layer8_outputs(1732) <= b and not a;
    layer8_outputs(1733) <= a or b;
    layer8_outputs(1734) <= not (a xor b);
    layer8_outputs(1735) <= not (a xor b);
    layer8_outputs(1736) <= not a;
    layer8_outputs(1737) <= not a;
    layer8_outputs(1738) <= not a;
    layer8_outputs(1739) <= not b or a;
    layer8_outputs(1740) <= a;
    layer8_outputs(1741) <= a and b;
    layer8_outputs(1742) <= a;
    layer8_outputs(1743) <= not (a and b);
    layer8_outputs(1744) <= not a or b;
    layer8_outputs(1745) <= not a;
    layer8_outputs(1746) <= not b;
    layer8_outputs(1747) <= a xor b;
    layer8_outputs(1748) <= a and b;
    layer8_outputs(1749) <= '0';
    layer8_outputs(1750) <= b;
    layer8_outputs(1751) <= b;
    layer8_outputs(1752) <= not b;
    layer8_outputs(1753) <= not a or b;
    layer8_outputs(1754) <= not (a and b);
    layer8_outputs(1755) <= not b;
    layer8_outputs(1756) <= not a;
    layer8_outputs(1757) <= not b;
    layer8_outputs(1758) <= not b or a;
    layer8_outputs(1759) <= not a;
    layer8_outputs(1760) <= not (a xor b);
    layer8_outputs(1761) <= a and not b;
    layer8_outputs(1762) <= not (a or b);
    layer8_outputs(1763) <= a or b;
    layer8_outputs(1764) <= not a;
    layer8_outputs(1765) <= a xor b;
    layer8_outputs(1766) <= a and not b;
    layer8_outputs(1767) <= not a;
    layer8_outputs(1768) <= b;
    layer8_outputs(1769) <= b;
    layer8_outputs(1770) <= b;
    layer8_outputs(1771) <= a xor b;
    layer8_outputs(1772) <= not a;
    layer8_outputs(1773) <= not (a xor b);
    layer8_outputs(1774) <= b and not a;
    layer8_outputs(1775) <= not b or a;
    layer8_outputs(1776) <= not b or a;
    layer8_outputs(1777) <= not a;
    layer8_outputs(1778) <= not (a xor b);
    layer8_outputs(1779) <= a and b;
    layer8_outputs(1780) <= not b;
    layer8_outputs(1781) <= not a or b;
    layer8_outputs(1782) <= a;
    layer8_outputs(1783) <= b and not a;
    layer8_outputs(1784) <= b;
    layer8_outputs(1785) <= not b;
    layer8_outputs(1786) <= not a;
    layer8_outputs(1787) <= b;
    layer8_outputs(1788) <= b;
    layer8_outputs(1789) <= b;
    layer8_outputs(1790) <= a;
    layer8_outputs(1791) <= a;
    layer8_outputs(1792) <= a and not b;
    layer8_outputs(1793) <= not a;
    layer8_outputs(1794) <= a;
    layer8_outputs(1795) <= b and not a;
    layer8_outputs(1796) <= not b;
    layer8_outputs(1797) <= a;
    layer8_outputs(1798) <= b;
    layer8_outputs(1799) <= a and b;
    layer8_outputs(1800) <= not (a and b);
    layer8_outputs(1801) <= a xor b;
    layer8_outputs(1802) <= a or b;
    layer8_outputs(1803) <= not (a or b);
    layer8_outputs(1804) <= a xor b;
    layer8_outputs(1805) <= not a or b;
    layer8_outputs(1806) <= not (a xor b);
    layer8_outputs(1807) <= a and b;
    layer8_outputs(1808) <= not (a xor b);
    layer8_outputs(1809) <= a xor b;
    layer8_outputs(1810) <= not b;
    layer8_outputs(1811) <= a and b;
    layer8_outputs(1812) <= not a;
    layer8_outputs(1813) <= not b;
    layer8_outputs(1814) <= a and not b;
    layer8_outputs(1815) <= not b;
    layer8_outputs(1816) <= a or b;
    layer8_outputs(1817) <= not (a xor b);
    layer8_outputs(1818) <= a xor b;
    layer8_outputs(1819) <= b;
    layer8_outputs(1820) <= a;
    layer8_outputs(1821) <= not a or b;
    layer8_outputs(1822) <= not (a xor b);
    layer8_outputs(1823) <= b and not a;
    layer8_outputs(1824) <= not a;
    layer8_outputs(1825) <= a xor b;
    layer8_outputs(1826) <= a xor b;
    layer8_outputs(1827) <= not (a xor b);
    layer8_outputs(1828) <= a;
    layer8_outputs(1829) <= not (a or b);
    layer8_outputs(1830) <= a and not b;
    layer8_outputs(1831) <= b and not a;
    layer8_outputs(1832) <= not b;
    layer8_outputs(1833) <= not b;
    layer8_outputs(1834) <= a;
    layer8_outputs(1835) <= not a or b;
    layer8_outputs(1836) <= a and b;
    layer8_outputs(1837) <= not b;
    layer8_outputs(1838) <= not a;
    layer8_outputs(1839) <= a xor b;
    layer8_outputs(1840) <= b;
    layer8_outputs(1841) <= a;
    layer8_outputs(1842) <= a xor b;
    layer8_outputs(1843) <= a xor b;
    layer8_outputs(1844) <= a;
    layer8_outputs(1845) <= not b;
    layer8_outputs(1846) <= a xor b;
    layer8_outputs(1847) <= not a;
    layer8_outputs(1848) <= a xor b;
    layer8_outputs(1849) <= not b;
    layer8_outputs(1850) <= not b;
    layer8_outputs(1851) <= b;
    layer8_outputs(1852) <= not a;
    layer8_outputs(1853) <= not (a xor b);
    layer8_outputs(1854) <= a xor b;
    layer8_outputs(1855) <= not a;
    layer8_outputs(1856) <= a and not b;
    layer8_outputs(1857) <= not (a xor b);
    layer8_outputs(1858) <= not a;
    layer8_outputs(1859) <= not (a xor b);
    layer8_outputs(1860) <= not b;
    layer8_outputs(1861) <= not b;
    layer8_outputs(1862) <= not (a xor b);
    layer8_outputs(1863) <= '0';
    layer8_outputs(1864) <= a and not b;
    layer8_outputs(1865) <= not b;
    layer8_outputs(1866) <= '1';
    layer8_outputs(1867) <= not b or a;
    layer8_outputs(1868) <= not (a xor b);
    layer8_outputs(1869) <= not a or b;
    layer8_outputs(1870) <= b and not a;
    layer8_outputs(1871) <= not (a or b);
    layer8_outputs(1872) <= b;
    layer8_outputs(1873) <= not (a xor b);
    layer8_outputs(1874) <= not (a and b);
    layer8_outputs(1875) <= not (a xor b);
    layer8_outputs(1876) <= not a or b;
    layer8_outputs(1877) <= a or b;
    layer8_outputs(1878) <= a;
    layer8_outputs(1879) <= a;
    layer8_outputs(1880) <= not a;
    layer8_outputs(1881) <= not a;
    layer8_outputs(1882) <= not a;
    layer8_outputs(1883) <= not (a xor b);
    layer8_outputs(1884) <= b;
    layer8_outputs(1885) <= not a;
    layer8_outputs(1886) <= b;
    layer8_outputs(1887) <= a;
    layer8_outputs(1888) <= not (a or b);
    layer8_outputs(1889) <= a or b;
    layer8_outputs(1890) <= not a;
    layer8_outputs(1891) <= a xor b;
    layer8_outputs(1892) <= not a;
    layer8_outputs(1893) <= a;
    layer8_outputs(1894) <= not b;
    layer8_outputs(1895) <= a xor b;
    layer8_outputs(1896) <= not a;
    layer8_outputs(1897) <= b;
    layer8_outputs(1898) <= a and b;
    layer8_outputs(1899) <= not (a and b);
    layer8_outputs(1900) <= not a;
    layer8_outputs(1901) <= a;
    layer8_outputs(1902) <= not b;
    layer8_outputs(1903) <= a;
    layer8_outputs(1904) <= not a;
    layer8_outputs(1905) <= a or b;
    layer8_outputs(1906) <= not (a and b);
    layer8_outputs(1907) <= not b;
    layer8_outputs(1908) <= a and b;
    layer8_outputs(1909) <= not a;
    layer8_outputs(1910) <= not (a xor b);
    layer8_outputs(1911) <= a xor b;
    layer8_outputs(1912) <= a;
    layer8_outputs(1913) <= a or b;
    layer8_outputs(1914) <= b and not a;
    layer8_outputs(1915) <= not b;
    layer8_outputs(1916) <= b;
    layer8_outputs(1917) <= not (a xor b);
    layer8_outputs(1918) <= not b;
    layer8_outputs(1919) <= a;
    layer8_outputs(1920) <= not (a or b);
    layer8_outputs(1921) <= not (a xor b);
    layer8_outputs(1922) <= not b;
    layer8_outputs(1923) <= a and not b;
    layer8_outputs(1924) <= not b;
    layer8_outputs(1925) <= a;
    layer8_outputs(1926) <= a or b;
    layer8_outputs(1927) <= not b;
    layer8_outputs(1928) <= b;
    layer8_outputs(1929) <= not a;
    layer8_outputs(1930) <= a and b;
    layer8_outputs(1931) <= not (a and b);
    layer8_outputs(1932) <= not b;
    layer8_outputs(1933) <= a;
    layer8_outputs(1934) <= not a;
    layer8_outputs(1935) <= a or b;
    layer8_outputs(1936) <= not b or a;
    layer8_outputs(1937) <= b;
    layer8_outputs(1938) <= not (a or b);
    layer8_outputs(1939) <= not b or a;
    layer8_outputs(1940) <= not a;
    layer8_outputs(1941) <= a xor b;
    layer8_outputs(1942) <= not a;
    layer8_outputs(1943) <= a xor b;
    layer8_outputs(1944) <= a or b;
    layer8_outputs(1945) <= not (a and b);
    layer8_outputs(1946) <= a xor b;
    layer8_outputs(1947) <= b;
    layer8_outputs(1948) <= not b or a;
    layer8_outputs(1949) <= '0';
    layer8_outputs(1950) <= not a;
    layer8_outputs(1951) <= not b;
    layer8_outputs(1952) <= not b;
    layer8_outputs(1953) <= not a;
    layer8_outputs(1954) <= a and not b;
    layer8_outputs(1955) <= a and b;
    layer8_outputs(1956) <= not b;
    layer8_outputs(1957) <= b;
    layer8_outputs(1958) <= not a or b;
    layer8_outputs(1959) <= a;
    layer8_outputs(1960) <= a xor b;
    layer8_outputs(1961) <= b and not a;
    layer8_outputs(1962) <= b and not a;
    layer8_outputs(1963) <= not a;
    layer8_outputs(1964) <= a and not b;
    layer8_outputs(1965) <= a and b;
    layer8_outputs(1966) <= a and b;
    layer8_outputs(1967) <= b;
    layer8_outputs(1968) <= a xor b;
    layer8_outputs(1969) <= b;
    layer8_outputs(1970) <= a xor b;
    layer8_outputs(1971) <= a and not b;
    layer8_outputs(1972) <= a or b;
    layer8_outputs(1973) <= not (a xor b);
    layer8_outputs(1974) <= not a;
    layer8_outputs(1975) <= not b;
    layer8_outputs(1976) <= not (a or b);
    layer8_outputs(1977) <= not (a or b);
    layer8_outputs(1978) <= b;
    layer8_outputs(1979) <= not a;
    layer8_outputs(1980) <= a xor b;
    layer8_outputs(1981) <= a;
    layer8_outputs(1982) <= not (a or b);
    layer8_outputs(1983) <= b;
    layer8_outputs(1984) <= not (a and b);
    layer8_outputs(1985) <= b and not a;
    layer8_outputs(1986) <= not b;
    layer8_outputs(1987) <= not b;
    layer8_outputs(1988) <= not (a or b);
    layer8_outputs(1989) <= b;
    layer8_outputs(1990) <= b and not a;
    layer8_outputs(1991) <= not (a and b);
    layer8_outputs(1992) <= a or b;
    layer8_outputs(1993) <= a xor b;
    layer8_outputs(1994) <= not a;
    layer8_outputs(1995) <= not (a and b);
    layer8_outputs(1996) <= a and not b;
    layer8_outputs(1997) <= not (a and b);
    layer8_outputs(1998) <= not (a xor b);
    layer8_outputs(1999) <= b;
    layer8_outputs(2000) <= a;
    layer8_outputs(2001) <= a;
    layer8_outputs(2002) <= a;
    layer8_outputs(2003) <= not a;
    layer8_outputs(2004) <= a and not b;
    layer8_outputs(2005) <= not b;
    layer8_outputs(2006) <= not b;
    layer8_outputs(2007) <= a and not b;
    layer8_outputs(2008) <= not (a xor b);
    layer8_outputs(2009) <= not a;
    layer8_outputs(2010) <= a;
    layer8_outputs(2011) <= not (a xor b);
    layer8_outputs(2012) <= not a;
    layer8_outputs(2013) <= a or b;
    layer8_outputs(2014) <= a xor b;
    layer8_outputs(2015) <= b;
    layer8_outputs(2016) <= not (a and b);
    layer8_outputs(2017) <= a;
    layer8_outputs(2018) <= not (a xor b);
    layer8_outputs(2019) <= a;
    layer8_outputs(2020) <= a or b;
    layer8_outputs(2021) <= a xor b;
    layer8_outputs(2022) <= b;
    layer8_outputs(2023) <= a;
    layer8_outputs(2024) <= not a;
    layer8_outputs(2025) <= not (a or b);
    layer8_outputs(2026) <= b and not a;
    layer8_outputs(2027) <= b;
    layer8_outputs(2028) <= not b;
    layer8_outputs(2029) <= not b;
    layer8_outputs(2030) <= b;
    layer8_outputs(2031) <= not (a xor b);
    layer8_outputs(2032) <= not (a and b);
    layer8_outputs(2033) <= b;
    layer8_outputs(2034) <= b and not a;
    layer8_outputs(2035) <= b;
    layer8_outputs(2036) <= not (a xor b);
    layer8_outputs(2037) <= a xor b;
    layer8_outputs(2038) <= a or b;
    layer8_outputs(2039) <= not a;
    layer8_outputs(2040) <= not (a xor b);
    layer8_outputs(2041) <= not b or a;
    layer8_outputs(2042) <= a;
    layer8_outputs(2043) <= not (a and b);
    layer8_outputs(2044) <= not a;
    layer8_outputs(2045) <= not a or b;
    layer8_outputs(2046) <= b and not a;
    layer8_outputs(2047) <= not b;
    layer8_outputs(2048) <= b;
    layer8_outputs(2049) <= a or b;
    layer8_outputs(2050) <= b;
    layer8_outputs(2051) <= a;
    layer8_outputs(2052) <= not a;
    layer8_outputs(2053) <= not a or b;
    layer8_outputs(2054) <= not a or b;
    layer8_outputs(2055) <= not (a or b);
    layer8_outputs(2056) <= not a or b;
    layer8_outputs(2057) <= not a;
    layer8_outputs(2058) <= not (a or b);
    layer8_outputs(2059) <= '0';
    layer8_outputs(2060) <= not a;
    layer8_outputs(2061) <= a;
    layer8_outputs(2062) <= b;
    layer8_outputs(2063) <= not (a xor b);
    layer8_outputs(2064) <= not b or a;
    layer8_outputs(2065) <= a xor b;
    layer8_outputs(2066) <= a;
    layer8_outputs(2067) <= not a or b;
    layer8_outputs(2068) <= a;
    layer8_outputs(2069) <= b;
    layer8_outputs(2070) <= a or b;
    layer8_outputs(2071) <= a;
    layer8_outputs(2072) <= a or b;
    layer8_outputs(2073) <= b;
    layer8_outputs(2074) <= not (a or b);
    layer8_outputs(2075) <= not (a xor b);
    layer8_outputs(2076) <= a xor b;
    layer8_outputs(2077) <= not b;
    layer8_outputs(2078) <= a and b;
    layer8_outputs(2079) <= not (a or b);
    layer8_outputs(2080) <= b and not a;
    layer8_outputs(2081) <= not b;
    layer8_outputs(2082) <= not (a xor b);
    layer8_outputs(2083) <= not b;
    layer8_outputs(2084) <= b;
    layer8_outputs(2085) <= b;
    layer8_outputs(2086) <= not (a xor b);
    layer8_outputs(2087) <= a;
    layer8_outputs(2088) <= b and not a;
    layer8_outputs(2089) <= a;
    layer8_outputs(2090) <= b;
    layer8_outputs(2091) <= b;
    layer8_outputs(2092) <= not (a xor b);
    layer8_outputs(2093) <= a or b;
    layer8_outputs(2094) <= not (a xor b);
    layer8_outputs(2095) <= not (a xor b);
    layer8_outputs(2096) <= a;
    layer8_outputs(2097) <= a and not b;
    layer8_outputs(2098) <= not a or b;
    layer8_outputs(2099) <= a and b;
    layer8_outputs(2100) <= not (a or b);
    layer8_outputs(2101) <= a and not b;
    layer8_outputs(2102) <= not b;
    layer8_outputs(2103) <= a and b;
    layer8_outputs(2104) <= not (a xor b);
    layer8_outputs(2105) <= not b;
    layer8_outputs(2106) <= a;
    layer8_outputs(2107) <= not b;
    layer8_outputs(2108) <= a and b;
    layer8_outputs(2109) <= not (a xor b);
    layer8_outputs(2110) <= not b;
    layer8_outputs(2111) <= b and not a;
    layer8_outputs(2112) <= a;
    layer8_outputs(2113) <= a xor b;
    layer8_outputs(2114) <= a and not b;
    layer8_outputs(2115) <= not a;
    layer8_outputs(2116) <= b;
    layer8_outputs(2117) <= not (a or b);
    layer8_outputs(2118) <= not (a xor b);
    layer8_outputs(2119) <= not (a xor b);
    layer8_outputs(2120) <= not b or a;
    layer8_outputs(2121) <= a;
    layer8_outputs(2122) <= not b;
    layer8_outputs(2123) <= not b or a;
    layer8_outputs(2124) <= not a;
    layer8_outputs(2125) <= not b;
    layer8_outputs(2126) <= not a;
    layer8_outputs(2127) <= not (a xor b);
    layer8_outputs(2128) <= not a or b;
    layer8_outputs(2129) <= not (a xor b);
    layer8_outputs(2130) <= not (a xor b);
    layer8_outputs(2131) <= a and not b;
    layer8_outputs(2132) <= not (a xor b);
    layer8_outputs(2133) <= not (a and b);
    layer8_outputs(2134) <= b;
    layer8_outputs(2135) <= a and b;
    layer8_outputs(2136) <= not b or a;
    layer8_outputs(2137) <= '0';
    layer8_outputs(2138) <= not (a and b);
    layer8_outputs(2139) <= a and not b;
    layer8_outputs(2140) <= a xor b;
    layer8_outputs(2141) <= not b;
    layer8_outputs(2142) <= b and not a;
    layer8_outputs(2143) <= not (a xor b);
    layer8_outputs(2144) <= b;
    layer8_outputs(2145) <= '1';
    layer8_outputs(2146) <= not b or a;
    layer8_outputs(2147) <= not a or b;
    layer8_outputs(2148) <= a xor b;
    layer8_outputs(2149) <= a or b;
    layer8_outputs(2150) <= a;
    layer8_outputs(2151) <= not (a or b);
    layer8_outputs(2152) <= a and b;
    layer8_outputs(2153) <= a;
    layer8_outputs(2154) <= a xor b;
    layer8_outputs(2155) <= not a or b;
    layer8_outputs(2156) <= a and not b;
    layer8_outputs(2157) <= a or b;
    layer8_outputs(2158) <= a or b;
    layer8_outputs(2159) <= not (a and b);
    layer8_outputs(2160) <= a or b;
    layer8_outputs(2161) <= b;
    layer8_outputs(2162) <= not a;
    layer8_outputs(2163) <= not (a and b);
    layer8_outputs(2164) <= not a;
    layer8_outputs(2165) <= a;
    layer8_outputs(2166) <= a and b;
    layer8_outputs(2167) <= not (a or b);
    layer8_outputs(2168) <= b;
    layer8_outputs(2169) <= a;
    layer8_outputs(2170) <= b and not a;
    layer8_outputs(2171) <= a and not b;
    layer8_outputs(2172) <= '1';
    layer8_outputs(2173) <= a;
    layer8_outputs(2174) <= not (a xor b);
    layer8_outputs(2175) <= a;
    layer8_outputs(2176) <= b and not a;
    layer8_outputs(2177) <= b;
    layer8_outputs(2178) <= b and not a;
    layer8_outputs(2179) <= not (a xor b);
    layer8_outputs(2180) <= not (a and b);
    layer8_outputs(2181) <= not b;
    layer8_outputs(2182) <= a;
    layer8_outputs(2183) <= not b;
    layer8_outputs(2184) <= not (a or b);
    layer8_outputs(2185) <= not (a or b);
    layer8_outputs(2186) <= not (a or b);
    layer8_outputs(2187) <= not b;
    layer8_outputs(2188) <= b and not a;
    layer8_outputs(2189) <= a and not b;
    layer8_outputs(2190) <= '0';
    layer8_outputs(2191) <= not b or a;
    layer8_outputs(2192) <= not (a xor b);
    layer8_outputs(2193) <= not (a and b);
    layer8_outputs(2194) <= not (a xor b);
    layer8_outputs(2195) <= not b;
    layer8_outputs(2196) <= not a;
    layer8_outputs(2197) <= b;
    layer8_outputs(2198) <= a and not b;
    layer8_outputs(2199) <= not (a xor b);
    layer8_outputs(2200) <= b;
    layer8_outputs(2201) <= not (a or b);
    layer8_outputs(2202) <= a;
    layer8_outputs(2203) <= b;
    layer8_outputs(2204) <= a;
    layer8_outputs(2205) <= not a;
    layer8_outputs(2206) <= not a;
    layer8_outputs(2207) <= not (a xor b);
    layer8_outputs(2208) <= not a;
    layer8_outputs(2209) <= a;
    layer8_outputs(2210) <= not a;
    layer8_outputs(2211) <= not b or a;
    layer8_outputs(2212) <= not a or b;
    layer8_outputs(2213) <= not (a xor b);
    layer8_outputs(2214) <= b;
    layer8_outputs(2215) <= not b;
    layer8_outputs(2216) <= b;
    layer8_outputs(2217) <= not a;
    layer8_outputs(2218) <= b;
    layer8_outputs(2219) <= a;
    layer8_outputs(2220) <= not (a xor b);
    layer8_outputs(2221) <= a and b;
    layer8_outputs(2222) <= a xor b;
    layer8_outputs(2223) <= b and not a;
    layer8_outputs(2224) <= b;
    layer8_outputs(2225) <= a xor b;
    layer8_outputs(2226) <= not (a and b);
    layer8_outputs(2227) <= a;
    layer8_outputs(2228) <= not b;
    layer8_outputs(2229) <= not (a xor b);
    layer8_outputs(2230) <= a xor b;
    layer8_outputs(2231) <= a xor b;
    layer8_outputs(2232) <= a xor b;
    layer8_outputs(2233) <= a xor b;
    layer8_outputs(2234) <= not (a and b);
    layer8_outputs(2235) <= not (a xor b);
    layer8_outputs(2236) <= a and not b;
    layer8_outputs(2237) <= a;
    layer8_outputs(2238) <= a;
    layer8_outputs(2239) <= a and b;
    layer8_outputs(2240) <= a;
    layer8_outputs(2241) <= not b;
    layer8_outputs(2242) <= b;
    layer8_outputs(2243) <= a xor b;
    layer8_outputs(2244) <= a;
    layer8_outputs(2245) <= a or b;
    layer8_outputs(2246) <= a and b;
    layer8_outputs(2247) <= b;
    layer8_outputs(2248) <= b;
    layer8_outputs(2249) <= b and not a;
    layer8_outputs(2250) <= not b or a;
    layer8_outputs(2251) <= not b;
    layer8_outputs(2252) <= a and b;
    layer8_outputs(2253) <= not (a xor b);
    layer8_outputs(2254) <= not b or a;
    layer8_outputs(2255) <= a or b;
    layer8_outputs(2256) <= a;
    layer8_outputs(2257) <= not (a or b);
    layer8_outputs(2258) <= b;
    layer8_outputs(2259) <= a;
    layer8_outputs(2260) <= b;
    layer8_outputs(2261) <= not b;
    layer8_outputs(2262) <= not (a xor b);
    layer8_outputs(2263) <= b and not a;
    layer8_outputs(2264) <= not a;
    layer8_outputs(2265) <= not (a or b);
    layer8_outputs(2266) <= not b;
    layer8_outputs(2267) <= a;
    layer8_outputs(2268) <= b and not a;
    layer8_outputs(2269) <= b;
    layer8_outputs(2270) <= not (a xor b);
    layer8_outputs(2271) <= a;
    layer8_outputs(2272) <= not (a or b);
    layer8_outputs(2273) <= not b or a;
    layer8_outputs(2274) <= a xor b;
    layer8_outputs(2275) <= a;
    layer8_outputs(2276) <= not b or a;
    layer8_outputs(2277) <= not (a and b);
    layer8_outputs(2278) <= a;
    layer8_outputs(2279) <= b;
    layer8_outputs(2280) <= not a;
    layer8_outputs(2281) <= a;
    layer8_outputs(2282) <= a and b;
    layer8_outputs(2283) <= a or b;
    layer8_outputs(2284) <= a and not b;
    layer8_outputs(2285) <= b and not a;
    layer8_outputs(2286) <= b;
    layer8_outputs(2287) <= not (a xor b);
    layer8_outputs(2288) <= a;
    layer8_outputs(2289) <= '0';
    layer8_outputs(2290) <= a;
    layer8_outputs(2291) <= not (a xor b);
    layer8_outputs(2292) <= not (a xor b);
    layer8_outputs(2293) <= b and not a;
    layer8_outputs(2294) <= b;
    layer8_outputs(2295) <= a;
    layer8_outputs(2296) <= not (a xor b);
    layer8_outputs(2297) <= not (a xor b);
    layer8_outputs(2298) <= a;
    layer8_outputs(2299) <= not (a xor b);
    layer8_outputs(2300) <= not b;
    layer8_outputs(2301) <= a;
    layer8_outputs(2302) <= a or b;
    layer8_outputs(2303) <= a;
    layer8_outputs(2304) <= a xor b;
    layer8_outputs(2305) <= a;
    layer8_outputs(2306) <= b;
    layer8_outputs(2307) <= a xor b;
    layer8_outputs(2308) <= a xor b;
    layer8_outputs(2309) <= a;
    layer8_outputs(2310) <= a xor b;
    layer8_outputs(2311) <= not a;
    layer8_outputs(2312) <= b;
    layer8_outputs(2313) <= a;
    layer8_outputs(2314) <= not b;
    layer8_outputs(2315) <= a or b;
    layer8_outputs(2316) <= not a;
    layer8_outputs(2317) <= not b;
    layer8_outputs(2318) <= a or b;
    layer8_outputs(2319) <= not a or b;
    layer8_outputs(2320) <= not b;
    layer8_outputs(2321) <= not (a or b);
    layer8_outputs(2322) <= b;
    layer8_outputs(2323) <= a xor b;
    layer8_outputs(2324) <= b;
    layer8_outputs(2325) <= a;
    layer8_outputs(2326) <= not (a or b);
    layer8_outputs(2327) <= a or b;
    layer8_outputs(2328) <= a;
    layer8_outputs(2329) <= a xor b;
    layer8_outputs(2330) <= not a or b;
    layer8_outputs(2331) <= not (a xor b);
    layer8_outputs(2332) <= not (a xor b);
    layer8_outputs(2333) <= b;
    layer8_outputs(2334) <= a and b;
    layer8_outputs(2335) <= not b;
    layer8_outputs(2336) <= not (a and b);
    layer8_outputs(2337) <= not (a and b);
    layer8_outputs(2338) <= a and b;
    layer8_outputs(2339) <= a xor b;
    layer8_outputs(2340) <= a and not b;
    layer8_outputs(2341) <= not b;
    layer8_outputs(2342) <= not a or b;
    layer8_outputs(2343) <= not (a xor b);
    layer8_outputs(2344) <= a and b;
    layer8_outputs(2345) <= not b;
    layer8_outputs(2346) <= not a;
    layer8_outputs(2347) <= not a;
    layer8_outputs(2348) <= not (a and b);
    layer8_outputs(2349) <= not b or a;
    layer8_outputs(2350) <= b;
    layer8_outputs(2351) <= not (a or b);
    layer8_outputs(2352) <= not b or a;
    layer8_outputs(2353) <= a;
    layer8_outputs(2354) <= b;
    layer8_outputs(2355) <= a and not b;
    layer8_outputs(2356) <= not b;
    layer8_outputs(2357) <= not (a and b);
    layer8_outputs(2358) <= not a;
    layer8_outputs(2359) <= not a;
    layer8_outputs(2360) <= not a;
    layer8_outputs(2361) <= not a;
    layer8_outputs(2362) <= a xor b;
    layer8_outputs(2363) <= b and not a;
    layer8_outputs(2364) <= not b;
    layer8_outputs(2365) <= not b;
    layer8_outputs(2366) <= not (a or b);
    layer8_outputs(2367) <= not (a and b);
    layer8_outputs(2368) <= not (a xor b);
    layer8_outputs(2369) <= a;
    layer8_outputs(2370) <= a;
    layer8_outputs(2371) <= a and not b;
    layer8_outputs(2372) <= b;
    layer8_outputs(2373) <= not (a and b);
    layer8_outputs(2374) <= not a or b;
    layer8_outputs(2375) <= not (a and b);
    layer8_outputs(2376) <= not (a or b);
    layer8_outputs(2377) <= a;
    layer8_outputs(2378) <= not (a xor b);
    layer8_outputs(2379) <= not (a xor b);
    layer8_outputs(2380) <= b;
    layer8_outputs(2381) <= not b;
    layer8_outputs(2382) <= not (a xor b);
    layer8_outputs(2383) <= not (a xor b);
    layer8_outputs(2384) <= '1';
    layer8_outputs(2385) <= a and not b;
    layer8_outputs(2386) <= not (a xor b);
    layer8_outputs(2387) <= b and not a;
    layer8_outputs(2388) <= a xor b;
    layer8_outputs(2389) <= not a;
    layer8_outputs(2390) <= a xor b;
    layer8_outputs(2391) <= not (a and b);
    layer8_outputs(2392) <= not b;
    layer8_outputs(2393) <= a and not b;
    layer8_outputs(2394) <= not a or b;
    layer8_outputs(2395) <= not (a xor b);
    layer8_outputs(2396) <= a and b;
    layer8_outputs(2397) <= b;
    layer8_outputs(2398) <= not (a and b);
    layer8_outputs(2399) <= a;
    layer8_outputs(2400) <= b;
    layer8_outputs(2401) <= not (a or b);
    layer8_outputs(2402) <= '1';
    layer8_outputs(2403) <= not a or b;
    layer8_outputs(2404) <= not a or b;
    layer8_outputs(2405) <= a;
    layer8_outputs(2406) <= a xor b;
    layer8_outputs(2407) <= b;
    layer8_outputs(2408) <= a and b;
    layer8_outputs(2409) <= not a;
    layer8_outputs(2410) <= not (a xor b);
    layer8_outputs(2411) <= not a;
    layer8_outputs(2412) <= a xor b;
    layer8_outputs(2413) <= a and not b;
    layer8_outputs(2414) <= not a;
    layer8_outputs(2415) <= a;
    layer8_outputs(2416) <= a;
    layer8_outputs(2417) <= not (a xor b);
    layer8_outputs(2418) <= not (a xor b);
    layer8_outputs(2419) <= not (a and b);
    layer8_outputs(2420) <= not b;
    layer8_outputs(2421) <= not a or b;
    layer8_outputs(2422) <= a xor b;
    layer8_outputs(2423) <= not (a or b);
    layer8_outputs(2424) <= not (a xor b);
    layer8_outputs(2425) <= a xor b;
    layer8_outputs(2426) <= b;
    layer8_outputs(2427) <= a;
    layer8_outputs(2428) <= a xor b;
    layer8_outputs(2429) <= a and not b;
    layer8_outputs(2430) <= b;
    layer8_outputs(2431) <= not (a xor b);
    layer8_outputs(2432) <= b and not a;
    layer8_outputs(2433) <= not (a xor b);
    layer8_outputs(2434) <= a and b;
    layer8_outputs(2435) <= not b;
    layer8_outputs(2436) <= not b or a;
    layer8_outputs(2437) <= not (a or b);
    layer8_outputs(2438) <= a;
    layer8_outputs(2439) <= a xor b;
    layer8_outputs(2440) <= a or b;
    layer8_outputs(2441) <= '1';
    layer8_outputs(2442) <= a and not b;
    layer8_outputs(2443) <= not b;
    layer8_outputs(2444) <= not (a xor b);
    layer8_outputs(2445) <= not (a xor b);
    layer8_outputs(2446) <= not b;
    layer8_outputs(2447) <= not (a and b);
    layer8_outputs(2448) <= not a or b;
    layer8_outputs(2449) <= not (a and b);
    layer8_outputs(2450) <= b and not a;
    layer8_outputs(2451) <= not (a xor b);
    layer8_outputs(2452) <= b and not a;
    layer8_outputs(2453) <= a or b;
    layer8_outputs(2454) <= a;
    layer8_outputs(2455) <= b and not a;
    layer8_outputs(2456) <= not (a and b);
    layer8_outputs(2457) <= not (a xor b);
    layer8_outputs(2458) <= a xor b;
    layer8_outputs(2459) <= b;
    layer8_outputs(2460) <= a xor b;
    layer8_outputs(2461) <= not b or a;
    layer8_outputs(2462) <= a;
    layer8_outputs(2463) <= a xor b;
    layer8_outputs(2464) <= not (a xor b);
    layer8_outputs(2465) <= b and not a;
    layer8_outputs(2466) <= not (a xor b);
    layer8_outputs(2467) <= '1';
    layer8_outputs(2468) <= a;
    layer8_outputs(2469) <= not a;
    layer8_outputs(2470) <= not b or a;
    layer8_outputs(2471) <= a xor b;
    layer8_outputs(2472) <= not a;
    layer8_outputs(2473) <= a xor b;
    layer8_outputs(2474) <= a;
    layer8_outputs(2475) <= a xor b;
    layer8_outputs(2476) <= a xor b;
    layer8_outputs(2477) <= not (a xor b);
    layer8_outputs(2478) <= not a;
    layer8_outputs(2479) <= a;
    layer8_outputs(2480) <= a xor b;
    layer8_outputs(2481) <= b;
    layer8_outputs(2482) <= a xor b;
    layer8_outputs(2483) <= not b;
    layer8_outputs(2484) <= b;
    layer8_outputs(2485) <= a;
    layer8_outputs(2486) <= a xor b;
    layer8_outputs(2487) <= b;
    layer8_outputs(2488) <= a and b;
    layer8_outputs(2489) <= a xor b;
    layer8_outputs(2490) <= not a;
    layer8_outputs(2491) <= a and not b;
    layer8_outputs(2492) <= a and b;
    layer8_outputs(2493) <= a xor b;
    layer8_outputs(2494) <= a and b;
    layer8_outputs(2495) <= b;
    layer8_outputs(2496) <= b;
    layer8_outputs(2497) <= not a;
    layer8_outputs(2498) <= a or b;
    layer8_outputs(2499) <= not b;
    layer8_outputs(2500) <= a xor b;
    layer8_outputs(2501) <= a and not b;
    layer8_outputs(2502) <= not (a xor b);
    layer8_outputs(2503) <= not b;
    layer8_outputs(2504) <= not b;
    layer8_outputs(2505) <= not b;
    layer8_outputs(2506) <= not a;
    layer8_outputs(2507) <= a;
    layer8_outputs(2508) <= not b;
    layer8_outputs(2509) <= a;
    layer8_outputs(2510) <= not b;
    layer8_outputs(2511) <= b and not a;
    layer8_outputs(2512) <= not b;
    layer8_outputs(2513) <= not b;
    layer8_outputs(2514) <= a and b;
    layer8_outputs(2515) <= not b or a;
    layer8_outputs(2516) <= not b or a;
    layer8_outputs(2517) <= not a;
    layer8_outputs(2518) <= a or b;
    layer8_outputs(2519) <= b;
    layer8_outputs(2520) <= not b or a;
    layer8_outputs(2521) <= b and not a;
    layer8_outputs(2522) <= b;
    layer8_outputs(2523) <= a and b;
    layer8_outputs(2524) <= not a or b;
    layer8_outputs(2525) <= a xor b;
    layer8_outputs(2526) <= not a;
    layer8_outputs(2527) <= b and not a;
    layer8_outputs(2528) <= not (a xor b);
    layer8_outputs(2529) <= a and not b;
    layer8_outputs(2530) <= b;
    layer8_outputs(2531) <= not (a and b);
    layer8_outputs(2532) <= not a;
    layer8_outputs(2533) <= not b;
    layer8_outputs(2534) <= not (a xor b);
    layer8_outputs(2535) <= a and b;
    layer8_outputs(2536) <= a or b;
    layer8_outputs(2537) <= a xor b;
    layer8_outputs(2538) <= '0';
    layer8_outputs(2539) <= a;
    layer8_outputs(2540) <= not b;
    layer8_outputs(2541) <= not (a xor b);
    layer8_outputs(2542) <= b;
    layer8_outputs(2543) <= a xor b;
    layer8_outputs(2544) <= a and not b;
    layer8_outputs(2545) <= not (a xor b);
    layer8_outputs(2546) <= a and not b;
    layer8_outputs(2547) <= not b;
    layer8_outputs(2548) <= a and b;
    layer8_outputs(2549) <= a and not b;
    layer8_outputs(2550) <= a xor b;
    layer8_outputs(2551) <= not a or b;
    layer8_outputs(2552) <= b;
    layer8_outputs(2553) <= not (a xor b);
    layer8_outputs(2554) <= b;
    layer8_outputs(2555) <= not (a xor b);
    layer8_outputs(2556) <= not b;
    layer8_outputs(2557) <= not b or a;
    layer8_outputs(2558) <= not a;
    layer8_outputs(2559) <= not (a xor b);
    layer8_outputs(2560) <= not b;
    layer8_outputs(2561) <= b and not a;
    layer8_outputs(2562) <= b;
    layer8_outputs(2563) <= b and not a;
    layer8_outputs(2564) <= b and not a;
    layer8_outputs(2565) <= not b;
    layer8_outputs(2566) <= b;
    layer8_outputs(2567) <= a;
    layer8_outputs(2568) <= not b or a;
    layer8_outputs(2569) <= not b or a;
    layer8_outputs(2570) <= a or b;
    layer8_outputs(2571) <= not a;
    layer8_outputs(2572) <= b;
    layer8_outputs(2573) <= not (a and b);
    layer8_outputs(2574) <= b;
    layer8_outputs(2575) <= a xor b;
    layer8_outputs(2576) <= a;
    layer8_outputs(2577) <= not b or a;
    layer8_outputs(2578) <= b;
    layer8_outputs(2579) <= a xor b;
    layer8_outputs(2580) <= not (a xor b);
    layer8_outputs(2581) <= not (a xor b);
    layer8_outputs(2582) <= not (a or b);
    layer8_outputs(2583) <= not a;
    layer8_outputs(2584) <= a and not b;
    layer8_outputs(2585) <= b;
    layer8_outputs(2586) <= not (a xor b);
    layer8_outputs(2587) <= not (a or b);
    layer8_outputs(2588) <= a xor b;
    layer8_outputs(2589) <= a;
    layer8_outputs(2590) <= not (a xor b);
    layer8_outputs(2591) <= not (a or b);
    layer8_outputs(2592) <= not (a and b);
    layer8_outputs(2593) <= a;
    layer8_outputs(2594) <= a and not b;
    layer8_outputs(2595) <= a;
    layer8_outputs(2596) <= not b;
    layer8_outputs(2597) <= not (a and b);
    layer8_outputs(2598) <= not b;
    layer8_outputs(2599) <= not (a and b);
    layer8_outputs(2600) <= a;
    layer8_outputs(2601) <= b;
    layer8_outputs(2602) <= a;
    layer8_outputs(2603) <= not a;
    layer8_outputs(2604) <= not (a and b);
    layer8_outputs(2605) <= not b;
    layer8_outputs(2606) <= a xor b;
    layer8_outputs(2607) <= not (a xor b);
    layer8_outputs(2608) <= a and not b;
    layer8_outputs(2609) <= not (a and b);
    layer8_outputs(2610) <= b and not a;
    layer8_outputs(2611) <= not b;
    layer8_outputs(2612) <= not a;
    layer8_outputs(2613) <= b and not a;
    layer8_outputs(2614) <= not (a or b);
    layer8_outputs(2615) <= a xor b;
    layer8_outputs(2616) <= a and b;
    layer8_outputs(2617) <= not a;
    layer8_outputs(2618) <= b;
    layer8_outputs(2619) <= not b;
    layer8_outputs(2620) <= not b;
    layer8_outputs(2621) <= not b;
    layer8_outputs(2622) <= b;
    layer8_outputs(2623) <= a;
    layer8_outputs(2624) <= a and b;
    layer8_outputs(2625) <= '1';
    layer8_outputs(2626) <= not a;
    layer8_outputs(2627) <= a or b;
    layer8_outputs(2628) <= not b;
    layer8_outputs(2629) <= b;
    layer8_outputs(2630) <= a;
    layer8_outputs(2631) <= not b;
    layer8_outputs(2632) <= '1';
    layer8_outputs(2633) <= b and not a;
    layer8_outputs(2634) <= a xor b;
    layer8_outputs(2635) <= not b;
    layer8_outputs(2636) <= a xor b;
    layer8_outputs(2637) <= b and not a;
    layer8_outputs(2638) <= not b or a;
    layer8_outputs(2639) <= not b;
    layer8_outputs(2640) <= not b;
    layer8_outputs(2641) <= a xor b;
    layer8_outputs(2642) <= not (a xor b);
    layer8_outputs(2643) <= not a;
    layer8_outputs(2644) <= a xor b;
    layer8_outputs(2645) <= not b;
    layer8_outputs(2646) <= not a;
    layer8_outputs(2647) <= not (a xor b);
    layer8_outputs(2648) <= a;
    layer8_outputs(2649) <= a or b;
    layer8_outputs(2650) <= a xor b;
    layer8_outputs(2651) <= a and b;
    layer8_outputs(2652) <= not (a xor b);
    layer8_outputs(2653) <= a and b;
    layer8_outputs(2654) <= not (a xor b);
    layer8_outputs(2655) <= a;
    layer8_outputs(2656) <= not (a and b);
    layer8_outputs(2657) <= not (a or b);
    layer8_outputs(2658) <= not b;
    layer8_outputs(2659) <= not b;
    layer8_outputs(2660) <= b;
    layer8_outputs(2661) <= not (a xor b);
    layer8_outputs(2662) <= a and b;
    layer8_outputs(2663) <= not b;
    layer8_outputs(2664) <= not b;
    layer8_outputs(2665) <= a xor b;
    layer8_outputs(2666) <= not (a xor b);
    layer8_outputs(2667) <= not (a and b);
    layer8_outputs(2668) <= not a;
    layer8_outputs(2669) <= b;
    layer8_outputs(2670) <= a xor b;
    layer8_outputs(2671) <= not b or a;
    layer8_outputs(2672) <= not (a or b);
    layer8_outputs(2673) <= b;
    layer8_outputs(2674) <= not b;
    layer8_outputs(2675) <= a;
    layer8_outputs(2676) <= a;
    layer8_outputs(2677) <= not a or b;
    layer8_outputs(2678) <= a;
    layer8_outputs(2679) <= not b;
    layer8_outputs(2680) <= a or b;
    layer8_outputs(2681) <= b;
    layer8_outputs(2682) <= a xor b;
    layer8_outputs(2683) <= a xor b;
    layer8_outputs(2684) <= b and not a;
    layer8_outputs(2685) <= not a or b;
    layer8_outputs(2686) <= not a;
    layer8_outputs(2687) <= a;
    layer8_outputs(2688) <= not (a and b);
    layer8_outputs(2689) <= not (a xor b);
    layer8_outputs(2690) <= a and b;
    layer8_outputs(2691) <= a;
    layer8_outputs(2692) <= not b;
    layer8_outputs(2693) <= b;
    layer8_outputs(2694) <= not b;
    layer8_outputs(2695) <= a and not b;
    layer8_outputs(2696) <= not b;
    layer8_outputs(2697) <= a or b;
    layer8_outputs(2698) <= not a;
    layer8_outputs(2699) <= not b or a;
    layer8_outputs(2700) <= a and b;
    layer8_outputs(2701) <= a xor b;
    layer8_outputs(2702) <= not b;
    layer8_outputs(2703) <= not a;
    layer8_outputs(2704) <= a and not b;
    layer8_outputs(2705) <= not (a xor b);
    layer8_outputs(2706) <= b and not a;
    layer8_outputs(2707) <= a and not b;
    layer8_outputs(2708) <= a;
    layer8_outputs(2709) <= not a;
    layer8_outputs(2710) <= not b or a;
    layer8_outputs(2711) <= b;
    layer8_outputs(2712) <= a;
    layer8_outputs(2713) <= a xor b;
    layer8_outputs(2714) <= not a or b;
    layer8_outputs(2715) <= not a or b;
    layer8_outputs(2716) <= a;
    layer8_outputs(2717) <= a;
    layer8_outputs(2718) <= not a or b;
    layer8_outputs(2719) <= a;
    layer8_outputs(2720) <= a xor b;
    layer8_outputs(2721) <= a;
    layer8_outputs(2722) <= a;
    layer8_outputs(2723) <= a xor b;
    layer8_outputs(2724) <= b;
    layer8_outputs(2725) <= not b;
    layer8_outputs(2726) <= not a;
    layer8_outputs(2727) <= a and b;
    layer8_outputs(2728) <= not b;
    layer8_outputs(2729) <= not a or b;
    layer8_outputs(2730) <= not b;
    layer8_outputs(2731) <= not b;
    layer8_outputs(2732) <= b and not a;
    layer8_outputs(2733) <= not (a xor b);
    layer8_outputs(2734) <= a and b;
    layer8_outputs(2735) <= b and not a;
    layer8_outputs(2736) <= not a;
    layer8_outputs(2737) <= '1';
    layer8_outputs(2738) <= a;
    layer8_outputs(2739) <= a and not b;
    layer8_outputs(2740) <= not a or b;
    layer8_outputs(2741) <= b;
    layer8_outputs(2742) <= a;
    layer8_outputs(2743) <= b;
    layer8_outputs(2744) <= a;
    layer8_outputs(2745) <= not b;
    layer8_outputs(2746) <= a or b;
    layer8_outputs(2747) <= b;
    layer8_outputs(2748) <= b;
    layer8_outputs(2749) <= a xor b;
    layer8_outputs(2750) <= not a;
    layer8_outputs(2751) <= b and not a;
    layer8_outputs(2752) <= not b;
    layer8_outputs(2753) <= not b or a;
    layer8_outputs(2754) <= a;
    layer8_outputs(2755) <= not b or a;
    layer8_outputs(2756) <= not a;
    layer8_outputs(2757) <= not a;
    layer8_outputs(2758) <= not a;
    layer8_outputs(2759) <= not a or b;
    layer8_outputs(2760) <= b;
    layer8_outputs(2761) <= a;
    layer8_outputs(2762) <= not a;
    layer8_outputs(2763) <= not a;
    layer8_outputs(2764) <= not a;
    layer8_outputs(2765) <= not (a and b);
    layer8_outputs(2766) <= not a;
    layer8_outputs(2767) <= b;
    layer8_outputs(2768) <= not b;
    layer8_outputs(2769) <= '0';
    layer8_outputs(2770) <= b and not a;
    layer8_outputs(2771) <= not (a or b);
    layer8_outputs(2772) <= not a;
    layer8_outputs(2773) <= a xor b;
    layer8_outputs(2774) <= not b or a;
    layer8_outputs(2775) <= a;
    layer8_outputs(2776) <= not a;
    layer8_outputs(2777) <= a or b;
    layer8_outputs(2778) <= not b or a;
    layer8_outputs(2779) <= not (a xor b);
    layer8_outputs(2780) <= not (a or b);
    layer8_outputs(2781) <= not b;
    layer8_outputs(2782) <= not b;
    layer8_outputs(2783) <= not a;
    layer8_outputs(2784) <= not b;
    layer8_outputs(2785) <= not b;
    layer8_outputs(2786) <= a or b;
    layer8_outputs(2787) <= b;
    layer8_outputs(2788) <= not (a xor b);
    layer8_outputs(2789) <= not b or a;
    layer8_outputs(2790) <= not (a xor b);
    layer8_outputs(2791) <= a or b;
    layer8_outputs(2792) <= a and b;
    layer8_outputs(2793) <= a;
    layer8_outputs(2794) <= not (a xor b);
    layer8_outputs(2795) <= not b;
    layer8_outputs(2796) <= a;
    layer8_outputs(2797) <= a or b;
    layer8_outputs(2798) <= a and not b;
    layer8_outputs(2799) <= not b or a;
    layer8_outputs(2800) <= not (a xor b);
    layer8_outputs(2801) <= a xor b;
    layer8_outputs(2802) <= a or b;
    layer8_outputs(2803) <= b;
    layer8_outputs(2804) <= not a or b;
    layer8_outputs(2805) <= not b;
    layer8_outputs(2806) <= not a or b;
    layer8_outputs(2807) <= not (a xor b);
    layer8_outputs(2808) <= a;
    layer8_outputs(2809) <= not a or b;
    layer8_outputs(2810) <= not (a xor b);
    layer8_outputs(2811) <= a or b;
    layer8_outputs(2812) <= b;
    layer8_outputs(2813) <= a and b;
    layer8_outputs(2814) <= not (a or b);
    layer8_outputs(2815) <= b and not a;
    layer8_outputs(2816) <= a;
    layer8_outputs(2817) <= b;
    layer8_outputs(2818) <= not b;
    layer8_outputs(2819) <= not (a or b);
    layer8_outputs(2820) <= a xor b;
    layer8_outputs(2821) <= not a;
    layer8_outputs(2822) <= not a;
    layer8_outputs(2823) <= not (a xor b);
    layer8_outputs(2824) <= not (a and b);
    layer8_outputs(2825) <= not (a and b);
    layer8_outputs(2826) <= not a;
    layer8_outputs(2827) <= a or b;
    layer8_outputs(2828) <= not (a xor b);
    layer8_outputs(2829) <= b and not a;
    layer8_outputs(2830) <= b;
    layer8_outputs(2831) <= not (a xor b);
    layer8_outputs(2832) <= not a;
    layer8_outputs(2833) <= not (a and b);
    layer8_outputs(2834) <= not (a or b);
    layer8_outputs(2835) <= a and not b;
    layer8_outputs(2836) <= a or b;
    layer8_outputs(2837) <= a;
    layer8_outputs(2838) <= b;
    layer8_outputs(2839) <= not (a xor b);
    layer8_outputs(2840) <= a and not b;
    layer8_outputs(2841) <= b and not a;
    layer8_outputs(2842) <= not b;
    layer8_outputs(2843) <= not b;
    layer8_outputs(2844) <= a or b;
    layer8_outputs(2845) <= not (a xor b);
    layer8_outputs(2846) <= a xor b;
    layer8_outputs(2847) <= b;
    layer8_outputs(2848) <= not b;
    layer8_outputs(2849) <= a or b;
    layer8_outputs(2850) <= b;
    layer8_outputs(2851) <= a;
    layer8_outputs(2852) <= b;
    layer8_outputs(2853) <= not (a xor b);
    layer8_outputs(2854) <= not a;
    layer8_outputs(2855) <= b and not a;
    layer8_outputs(2856) <= not (a or b);
    layer8_outputs(2857) <= not (a and b);
    layer8_outputs(2858) <= not (a or b);
    layer8_outputs(2859) <= a;
    layer8_outputs(2860) <= not (a or b);
    layer8_outputs(2861) <= not (a xor b);
    layer8_outputs(2862) <= not a;
    layer8_outputs(2863) <= not b;
    layer8_outputs(2864) <= '0';
    layer8_outputs(2865) <= a;
    layer8_outputs(2866) <= b and not a;
    layer8_outputs(2867) <= b;
    layer8_outputs(2868) <= not (a or b);
    layer8_outputs(2869) <= b;
    layer8_outputs(2870) <= a or b;
    layer8_outputs(2871) <= a and not b;
    layer8_outputs(2872) <= not a;
    layer8_outputs(2873) <= not (a or b);
    layer8_outputs(2874) <= not (a xor b);
    layer8_outputs(2875) <= a and b;
    layer8_outputs(2876) <= a or b;
    layer8_outputs(2877) <= not a;
    layer8_outputs(2878) <= a or b;
    layer8_outputs(2879) <= a;
    layer8_outputs(2880) <= not a;
    layer8_outputs(2881) <= b;
    layer8_outputs(2882) <= not (a xor b);
    layer8_outputs(2883) <= a;
    layer8_outputs(2884) <= a and b;
    layer8_outputs(2885) <= not (a xor b);
    layer8_outputs(2886) <= not (a and b);
    layer8_outputs(2887) <= a and b;
    layer8_outputs(2888) <= b;
    layer8_outputs(2889) <= not b;
    layer8_outputs(2890) <= a or b;
    layer8_outputs(2891) <= b;
    layer8_outputs(2892) <= not b;
    layer8_outputs(2893) <= a;
    layer8_outputs(2894) <= b;
    layer8_outputs(2895) <= b;
    layer8_outputs(2896) <= a;
    layer8_outputs(2897) <= a or b;
    layer8_outputs(2898) <= a;
    layer8_outputs(2899) <= a;
    layer8_outputs(2900) <= a xor b;
    layer8_outputs(2901) <= a or b;
    layer8_outputs(2902) <= a;
    layer8_outputs(2903) <= a or b;
    layer8_outputs(2904) <= a or b;
    layer8_outputs(2905) <= a and not b;
    layer8_outputs(2906) <= not (a and b);
    layer8_outputs(2907) <= b and not a;
    layer8_outputs(2908) <= b and not a;
    layer8_outputs(2909) <= a or b;
    layer8_outputs(2910) <= b and not a;
    layer8_outputs(2911) <= a xor b;
    layer8_outputs(2912) <= a and not b;
    layer8_outputs(2913) <= not b or a;
    layer8_outputs(2914) <= a and b;
    layer8_outputs(2915) <= not a;
    layer8_outputs(2916) <= not (a and b);
    layer8_outputs(2917) <= not b or a;
    layer8_outputs(2918) <= not b or a;
    layer8_outputs(2919) <= a and b;
    layer8_outputs(2920) <= not b or a;
    layer8_outputs(2921) <= a or b;
    layer8_outputs(2922) <= b and not a;
    layer8_outputs(2923) <= not (a and b);
    layer8_outputs(2924) <= a and not b;
    layer8_outputs(2925) <= not b or a;
    layer8_outputs(2926) <= a xor b;
    layer8_outputs(2927) <= not a;
    layer8_outputs(2928) <= a;
    layer8_outputs(2929) <= b;
    layer8_outputs(2930) <= not (a xor b);
    layer8_outputs(2931) <= not b or a;
    layer8_outputs(2932) <= a or b;
    layer8_outputs(2933) <= a and not b;
    layer8_outputs(2934) <= a;
    layer8_outputs(2935) <= a;
    layer8_outputs(2936) <= not b;
    layer8_outputs(2937) <= not a;
    layer8_outputs(2938) <= not b;
    layer8_outputs(2939) <= b;
    layer8_outputs(2940) <= a;
    layer8_outputs(2941) <= a;
    layer8_outputs(2942) <= a xor b;
    layer8_outputs(2943) <= a;
    layer8_outputs(2944) <= b and not a;
    layer8_outputs(2945) <= a;
    layer8_outputs(2946) <= b;
    layer8_outputs(2947) <= not b;
    layer8_outputs(2948) <= not b or a;
    layer8_outputs(2949) <= not a;
    layer8_outputs(2950) <= not a;
    layer8_outputs(2951) <= a xor b;
    layer8_outputs(2952) <= a;
    layer8_outputs(2953) <= not b;
    layer8_outputs(2954) <= not b or a;
    layer8_outputs(2955) <= b;
    layer8_outputs(2956) <= a;
    layer8_outputs(2957) <= a;
    layer8_outputs(2958) <= a;
    layer8_outputs(2959) <= b;
    layer8_outputs(2960) <= a;
    layer8_outputs(2961) <= not (a or b);
    layer8_outputs(2962) <= not b or a;
    layer8_outputs(2963) <= not (a or b);
    layer8_outputs(2964) <= not b;
    layer8_outputs(2965) <= not (a and b);
    layer8_outputs(2966) <= not b;
    layer8_outputs(2967) <= b;
    layer8_outputs(2968) <= not b;
    layer8_outputs(2969) <= b;
    layer8_outputs(2970) <= not a or b;
    layer8_outputs(2971) <= not b;
    layer8_outputs(2972) <= not (a or b);
    layer8_outputs(2973) <= not a;
    layer8_outputs(2974) <= not b or a;
    layer8_outputs(2975) <= not b;
    layer8_outputs(2976) <= a;
    layer8_outputs(2977) <= not b or a;
    layer8_outputs(2978) <= not b;
    layer8_outputs(2979) <= not a;
    layer8_outputs(2980) <= not (a xor b);
    layer8_outputs(2981) <= not b or a;
    layer8_outputs(2982) <= a;
    layer8_outputs(2983) <= not b;
    layer8_outputs(2984) <= b;
    layer8_outputs(2985) <= a xor b;
    layer8_outputs(2986) <= a;
    layer8_outputs(2987) <= a and b;
    layer8_outputs(2988) <= a;
    layer8_outputs(2989) <= a;
    layer8_outputs(2990) <= b;
    layer8_outputs(2991) <= a;
    layer8_outputs(2992) <= not (a xor b);
    layer8_outputs(2993) <= not a;
    layer8_outputs(2994) <= not b;
    layer8_outputs(2995) <= a xor b;
    layer8_outputs(2996) <= b;
    layer8_outputs(2997) <= not b;
    layer8_outputs(2998) <= not a or b;
    layer8_outputs(2999) <= not a or b;
    layer8_outputs(3000) <= a and not b;
    layer8_outputs(3001) <= b;
    layer8_outputs(3002) <= b;
    layer8_outputs(3003) <= b;
    layer8_outputs(3004) <= a xor b;
    layer8_outputs(3005) <= b;
    layer8_outputs(3006) <= a xor b;
    layer8_outputs(3007) <= b;
    layer8_outputs(3008) <= not (a xor b);
    layer8_outputs(3009) <= not a;
    layer8_outputs(3010) <= a xor b;
    layer8_outputs(3011) <= a xor b;
    layer8_outputs(3012) <= not b;
    layer8_outputs(3013) <= a;
    layer8_outputs(3014) <= b and not a;
    layer8_outputs(3015) <= b;
    layer8_outputs(3016) <= not b or a;
    layer8_outputs(3017) <= not b or a;
    layer8_outputs(3018) <= not (a and b);
    layer8_outputs(3019) <= not (a and b);
    layer8_outputs(3020) <= a;
    layer8_outputs(3021) <= not (a xor b);
    layer8_outputs(3022) <= not b;
    layer8_outputs(3023) <= not b;
    layer8_outputs(3024) <= '1';
    layer8_outputs(3025) <= not (a or b);
    layer8_outputs(3026) <= not a;
    layer8_outputs(3027) <= b;
    layer8_outputs(3028) <= a or b;
    layer8_outputs(3029) <= not (a and b);
    layer8_outputs(3030) <= not (a xor b);
    layer8_outputs(3031) <= a;
    layer8_outputs(3032) <= a and b;
    layer8_outputs(3033) <= b and not a;
    layer8_outputs(3034) <= b;
    layer8_outputs(3035) <= a and b;
    layer8_outputs(3036) <= not b;
    layer8_outputs(3037) <= not a;
    layer8_outputs(3038) <= a xor b;
    layer8_outputs(3039) <= a xor b;
    layer8_outputs(3040) <= not a or b;
    layer8_outputs(3041) <= a xor b;
    layer8_outputs(3042) <= a;
    layer8_outputs(3043) <= a;
    layer8_outputs(3044) <= a;
    layer8_outputs(3045) <= not b;
    layer8_outputs(3046) <= a;
    layer8_outputs(3047) <= a;
    layer8_outputs(3048) <= b;
    layer8_outputs(3049) <= a xor b;
    layer8_outputs(3050) <= not (a or b);
    layer8_outputs(3051) <= not a;
    layer8_outputs(3052) <= not b;
    layer8_outputs(3053) <= not b;
    layer8_outputs(3054) <= b and not a;
    layer8_outputs(3055) <= not a;
    layer8_outputs(3056) <= '1';
    layer8_outputs(3057) <= not b;
    layer8_outputs(3058) <= a or b;
    layer8_outputs(3059) <= not (a or b);
    layer8_outputs(3060) <= a and b;
    layer8_outputs(3061) <= not a or b;
    layer8_outputs(3062) <= a xor b;
    layer8_outputs(3063) <= not a;
    layer8_outputs(3064) <= b;
    layer8_outputs(3065) <= a;
    layer8_outputs(3066) <= not a;
    layer8_outputs(3067) <= a or b;
    layer8_outputs(3068) <= not (a and b);
    layer8_outputs(3069) <= b;
    layer8_outputs(3070) <= a;
    layer8_outputs(3071) <= not (a and b);
    layer8_outputs(3072) <= not (a and b);
    layer8_outputs(3073) <= a xor b;
    layer8_outputs(3074) <= not (a or b);
    layer8_outputs(3075) <= not b or a;
    layer8_outputs(3076) <= not (a xor b);
    layer8_outputs(3077) <= not (a and b);
    layer8_outputs(3078) <= not a or b;
    layer8_outputs(3079) <= b and not a;
    layer8_outputs(3080) <= not (a xor b);
    layer8_outputs(3081) <= not a or b;
    layer8_outputs(3082) <= not b;
    layer8_outputs(3083) <= not (a xor b);
    layer8_outputs(3084) <= a xor b;
    layer8_outputs(3085) <= a or b;
    layer8_outputs(3086) <= not a;
    layer8_outputs(3087) <= a xor b;
    layer8_outputs(3088) <= b;
    layer8_outputs(3089) <= not (a or b);
    layer8_outputs(3090) <= a;
    layer8_outputs(3091) <= '1';
    layer8_outputs(3092) <= not a;
    layer8_outputs(3093) <= a;
    layer8_outputs(3094) <= a;
    layer8_outputs(3095) <= a and not b;
    layer8_outputs(3096) <= not b;
    layer8_outputs(3097) <= not (a or b);
    layer8_outputs(3098) <= not (a xor b);
    layer8_outputs(3099) <= a;
    layer8_outputs(3100) <= not b or a;
    layer8_outputs(3101) <= a and b;
    layer8_outputs(3102) <= b;
    layer8_outputs(3103) <= not (a xor b);
    layer8_outputs(3104) <= not (a xor b);
    layer8_outputs(3105) <= not (a and b);
    layer8_outputs(3106) <= not (a or b);
    layer8_outputs(3107) <= not a or b;
    layer8_outputs(3108) <= a and b;
    layer8_outputs(3109) <= a xor b;
    layer8_outputs(3110) <= not a;
    layer8_outputs(3111) <= a xor b;
    layer8_outputs(3112) <= not a or b;
    layer8_outputs(3113) <= not a;
    layer8_outputs(3114) <= not (a and b);
    layer8_outputs(3115) <= not (a xor b);
    layer8_outputs(3116) <= not b or a;
    layer8_outputs(3117) <= not (a and b);
    layer8_outputs(3118) <= b;
    layer8_outputs(3119) <= not b;
    layer8_outputs(3120) <= a and not b;
    layer8_outputs(3121) <= not b or a;
    layer8_outputs(3122) <= not (a xor b);
    layer8_outputs(3123) <= not (a xor b);
    layer8_outputs(3124) <= not (a or b);
    layer8_outputs(3125) <= not (a or b);
    layer8_outputs(3126) <= not a;
    layer8_outputs(3127) <= a and not b;
    layer8_outputs(3128) <= not (a and b);
    layer8_outputs(3129) <= not b;
    layer8_outputs(3130) <= b and not a;
    layer8_outputs(3131) <= not (a or b);
    layer8_outputs(3132) <= a;
    layer8_outputs(3133) <= not b;
    layer8_outputs(3134) <= not (a xor b);
    layer8_outputs(3135) <= not (a or b);
    layer8_outputs(3136) <= not b;
    layer8_outputs(3137) <= not a;
    layer8_outputs(3138) <= not (a xor b);
    layer8_outputs(3139) <= b and not a;
    layer8_outputs(3140) <= not b;
    layer8_outputs(3141) <= not (a xor b);
    layer8_outputs(3142) <= not b;
    layer8_outputs(3143) <= a;
    layer8_outputs(3144) <= a and not b;
    layer8_outputs(3145) <= a;
    layer8_outputs(3146) <= not a;
    layer8_outputs(3147) <= not b;
    layer8_outputs(3148) <= not (a and b);
    layer8_outputs(3149) <= a and not b;
    layer8_outputs(3150) <= not b;
    layer8_outputs(3151) <= b and not a;
    layer8_outputs(3152) <= '0';
    layer8_outputs(3153) <= not (a or b);
    layer8_outputs(3154) <= a;
    layer8_outputs(3155) <= not (a or b);
    layer8_outputs(3156) <= not b;
    layer8_outputs(3157) <= a xor b;
    layer8_outputs(3158) <= not b or a;
    layer8_outputs(3159) <= not b;
    layer8_outputs(3160) <= not (a xor b);
    layer8_outputs(3161) <= b;
    layer8_outputs(3162) <= a xor b;
    layer8_outputs(3163) <= not (a xor b);
    layer8_outputs(3164) <= not a;
    layer8_outputs(3165) <= a xor b;
    layer8_outputs(3166) <= a xor b;
    layer8_outputs(3167) <= a and b;
    layer8_outputs(3168) <= a;
    layer8_outputs(3169) <= a;
    layer8_outputs(3170) <= b and not a;
    layer8_outputs(3171) <= a xor b;
    layer8_outputs(3172) <= not a or b;
    layer8_outputs(3173) <= not b or a;
    layer8_outputs(3174) <= not b;
    layer8_outputs(3175) <= a and not b;
    layer8_outputs(3176) <= not (a xor b);
    layer8_outputs(3177) <= not a or b;
    layer8_outputs(3178) <= a and not b;
    layer8_outputs(3179) <= a;
    layer8_outputs(3180) <= b;
    layer8_outputs(3181) <= not a;
    layer8_outputs(3182) <= '1';
    layer8_outputs(3183) <= b;
    layer8_outputs(3184) <= not b;
    layer8_outputs(3185) <= a and not b;
    layer8_outputs(3186) <= not b or a;
    layer8_outputs(3187) <= a xor b;
    layer8_outputs(3188) <= b;
    layer8_outputs(3189) <= not (a xor b);
    layer8_outputs(3190) <= not (a or b);
    layer8_outputs(3191) <= b;
    layer8_outputs(3192) <= a or b;
    layer8_outputs(3193) <= a xor b;
    layer8_outputs(3194) <= not a or b;
    layer8_outputs(3195) <= not (a xor b);
    layer8_outputs(3196) <= b;
    layer8_outputs(3197) <= a;
    layer8_outputs(3198) <= not (a xor b);
    layer8_outputs(3199) <= b;
    layer8_outputs(3200) <= not b;
    layer8_outputs(3201) <= not a;
    layer8_outputs(3202) <= a xor b;
    layer8_outputs(3203) <= a;
    layer8_outputs(3204) <= a and not b;
    layer8_outputs(3205) <= not a;
    layer8_outputs(3206) <= not a;
    layer8_outputs(3207) <= not a or b;
    layer8_outputs(3208) <= not (a xor b);
    layer8_outputs(3209) <= a or b;
    layer8_outputs(3210) <= not b;
    layer8_outputs(3211) <= not a;
    layer8_outputs(3212) <= not (a xor b);
    layer8_outputs(3213) <= a;
    layer8_outputs(3214) <= b;
    layer8_outputs(3215) <= '0';
    layer8_outputs(3216) <= not a or b;
    layer8_outputs(3217) <= not (a and b);
    layer8_outputs(3218) <= not (a and b);
    layer8_outputs(3219) <= a xor b;
    layer8_outputs(3220) <= not b or a;
    layer8_outputs(3221) <= a xor b;
    layer8_outputs(3222) <= not (a and b);
    layer8_outputs(3223) <= a;
    layer8_outputs(3224) <= not a;
    layer8_outputs(3225) <= not a;
    layer8_outputs(3226) <= not a or b;
    layer8_outputs(3227) <= b;
    layer8_outputs(3228) <= a xor b;
    layer8_outputs(3229) <= not (a xor b);
    layer8_outputs(3230) <= a xor b;
    layer8_outputs(3231) <= a;
    layer8_outputs(3232) <= a;
    layer8_outputs(3233) <= b;
    layer8_outputs(3234) <= a;
    layer8_outputs(3235) <= not a;
    layer8_outputs(3236) <= not (a xor b);
    layer8_outputs(3237) <= not a;
    layer8_outputs(3238) <= not b;
    layer8_outputs(3239) <= not b;
    layer8_outputs(3240) <= a;
    layer8_outputs(3241) <= '0';
    layer8_outputs(3242) <= b;
    layer8_outputs(3243) <= a;
    layer8_outputs(3244) <= a and b;
    layer8_outputs(3245) <= a xor b;
    layer8_outputs(3246) <= not b or a;
    layer8_outputs(3247) <= a and not b;
    layer8_outputs(3248) <= a;
    layer8_outputs(3249) <= not (a or b);
    layer8_outputs(3250) <= not a;
    layer8_outputs(3251) <= a and b;
    layer8_outputs(3252) <= b and not a;
    layer8_outputs(3253) <= b;
    layer8_outputs(3254) <= a and not b;
    layer8_outputs(3255) <= '0';
    layer8_outputs(3256) <= not a;
    layer8_outputs(3257) <= not b;
    layer8_outputs(3258) <= a and b;
    layer8_outputs(3259) <= b;
    layer8_outputs(3260) <= a xor b;
    layer8_outputs(3261) <= not b;
    layer8_outputs(3262) <= '1';
    layer8_outputs(3263) <= a and b;
    layer8_outputs(3264) <= not b or a;
    layer8_outputs(3265) <= not b;
    layer8_outputs(3266) <= not (a and b);
    layer8_outputs(3267) <= a and b;
    layer8_outputs(3268) <= not (a xor b);
    layer8_outputs(3269) <= not (a and b);
    layer8_outputs(3270) <= not a;
    layer8_outputs(3271) <= a xor b;
    layer8_outputs(3272) <= a and not b;
    layer8_outputs(3273) <= a;
    layer8_outputs(3274) <= a xor b;
    layer8_outputs(3275) <= not (a or b);
    layer8_outputs(3276) <= not b or a;
    layer8_outputs(3277) <= not a;
    layer8_outputs(3278) <= a xor b;
    layer8_outputs(3279) <= not (a xor b);
    layer8_outputs(3280) <= not (a xor b);
    layer8_outputs(3281) <= a or b;
    layer8_outputs(3282) <= a;
    layer8_outputs(3283) <= b;
    layer8_outputs(3284) <= b;
    layer8_outputs(3285) <= a xor b;
    layer8_outputs(3286) <= a and b;
    layer8_outputs(3287) <= not a;
    layer8_outputs(3288) <= not a;
    layer8_outputs(3289) <= a or b;
    layer8_outputs(3290) <= a or b;
    layer8_outputs(3291) <= not (a xor b);
    layer8_outputs(3292) <= a xor b;
    layer8_outputs(3293) <= not (a and b);
    layer8_outputs(3294) <= not (a and b);
    layer8_outputs(3295) <= not a;
    layer8_outputs(3296) <= a and b;
    layer8_outputs(3297) <= b and not a;
    layer8_outputs(3298) <= not (a and b);
    layer8_outputs(3299) <= a xor b;
    layer8_outputs(3300) <= a;
    layer8_outputs(3301) <= not (a xor b);
    layer8_outputs(3302) <= not (a or b);
    layer8_outputs(3303) <= a xor b;
    layer8_outputs(3304) <= not a;
    layer8_outputs(3305) <= a or b;
    layer8_outputs(3306) <= not a;
    layer8_outputs(3307) <= not (a xor b);
    layer8_outputs(3308) <= not (a and b);
    layer8_outputs(3309) <= not b or a;
    layer8_outputs(3310) <= b and not a;
    layer8_outputs(3311) <= a xor b;
    layer8_outputs(3312) <= a;
    layer8_outputs(3313) <= a xor b;
    layer8_outputs(3314) <= not b;
    layer8_outputs(3315) <= a xor b;
    layer8_outputs(3316) <= a and b;
    layer8_outputs(3317) <= not a;
    layer8_outputs(3318) <= b and not a;
    layer8_outputs(3319) <= b and not a;
    layer8_outputs(3320) <= not (a and b);
    layer8_outputs(3321) <= b;
    layer8_outputs(3322) <= not b or a;
    layer8_outputs(3323) <= not a;
    layer8_outputs(3324) <= not (a xor b);
    layer8_outputs(3325) <= a;
    layer8_outputs(3326) <= b and not a;
    layer8_outputs(3327) <= a;
    layer8_outputs(3328) <= not a;
    layer8_outputs(3329) <= b;
    layer8_outputs(3330) <= not (a or b);
    layer8_outputs(3331) <= a;
    layer8_outputs(3332) <= not (a and b);
    layer8_outputs(3333) <= b;
    layer8_outputs(3334) <= b;
    layer8_outputs(3335) <= a and b;
    layer8_outputs(3336) <= not a;
    layer8_outputs(3337) <= not (a or b);
    layer8_outputs(3338) <= a and b;
    layer8_outputs(3339) <= not (a xor b);
    layer8_outputs(3340) <= not (a or b);
    layer8_outputs(3341) <= b and not a;
    layer8_outputs(3342) <= not (a and b);
    layer8_outputs(3343) <= a;
    layer8_outputs(3344) <= not b or a;
    layer8_outputs(3345) <= a;
    layer8_outputs(3346) <= not b or a;
    layer8_outputs(3347) <= not b or a;
    layer8_outputs(3348) <= a and not b;
    layer8_outputs(3349) <= b and not a;
    layer8_outputs(3350) <= b;
    layer8_outputs(3351) <= b;
    layer8_outputs(3352) <= a;
    layer8_outputs(3353) <= a xor b;
    layer8_outputs(3354) <= b;
    layer8_outputs(3355) <= b;
    layer8_outputs(3356) <= b;
    layer8_outputs(3357) <= not b;
    layer8_outputs(3358) <= b and not a;
    layer8_outputs(3359) <= a xor b;
    layer8_outputs(3360) <= not (a xor b);
    layer8_outputs(3361) <= a;
    layer8_outputs(3362) <= not (a xor b);
    layer8_outputs(3363) <= not a;
    layer8_outputs(3364) <= not a;
    layer8_outputs(3365) <= b and not a;
    layer8_outputs(3366) <= not b;
    layer8_outputs(3367) <= not a;
    layer8_outputs(3368) <= b;
    layer8_outputs(3369) <= not b;
    layer8_outputs(3370) <= b;
    layer8_outputs(3371) <= a;
    layer8_outputs(3372) <= not (a and b);
    layer8_outputs(3373) <= a;
    layer8_outputs(3374) <= not b or a;
    layer8_outputs(3375) <= b;
    layer8_outputs(3376) <= a;
    layer8_outputs(3377) <= not b;
    layer8_outputs(3378) <= b;
    layer8_outputs(3379) <= b and not a;
    layer8_outputs(3380) <= a or b;
    layer8_outputs(3381) <= not (a and b);
    layer8_outputs(3382) <= a and b;
    layer8_outputs(3383) <= not a or b;
    layer8_outputs(3384) <= not (a or b);
    layer8_outputs(3385) <= not (a xor b);
    layer8_outputs(3386) <= not a;
    layer8_outputs(3387) <= not b or a;
    layer8_outputs(3388) <= a and not b;
    layer8_outputs(3389) <= b;
    layer8_outputs(3390) <= b;
    layer8_outputs(3391) <= not a;
    layer8_outputs(3392) <= not b;
    layer8_outputs(3393) <= a xor b;
    layer8_outputs(3394) <= not b or a;
    layer8_outputs(3395) <= not (a and b);
    layer8_outputs(3396) <= not a or b;
    layer8_outputs(3397) <= not (a xor b);
    layer8_outputs(3398) <= not a;
    layer8_outputs(3399) <= not a;
    layer8_outputs(3400) <= not a or b;
    layer8_outputs(3401) <= a xor b;
    layer8_outputs(3402) <= '1';
    layer8_outputs(3403) <= not a;
    layer8_outputs(3404) <= not a;
    layer8_outputs(3405) <= not b;
    layer8_outputs(3406) <= not a or b;
    layer8_outputs(3407) <= a and not b;
    layer8_outputs(3408) <= not a;
    layer8_outputs(3409) <= not a;
    layer8_outputs(3410) <= a and b;
    layer8_outputs(3411) <= not b;
    layer8_outputs(3412) <= b;
    layer8_outputs(3413) <= a or b;
    layer8_outputs(3414) <= not a;
    layer8_outputs(3415) <= not a;
    layer8_outputs(3416) <= not b;
    layer8_outputs(3417) <= a and not b;
    layer8_outputs(3418) <= b and not a;
    layer8_outputs(3419) <= not b;
    layer8_outputs(3420) <= b;
    layer8_outputs(3421) <= b;
    layer8_outputs(3422) <= a xor b;
    layer8_outputs(3423) <= not (a and b);
    layer8_outputs(3424) <= a;
    layer8_outputs(3425) <= a xor b;
    layer8_outputs(3426) <= a;
    layer8_outputs(3427) <= a or b;
    layer8_outputs(3428) <= not b;
    layer8_outputs(3429) <= a;
    layer8_outputs(3430) <= a;
    layer8_outputs(3431) <= a or b;
    layer8_outputs(3432) <= not (a and b);
    layer8_outputs(3433) <= a and not b;
    layer8_outputs(3434) <= not a;
    layer8_outputs(3435) <= a;
    layer8_outputs(3436) <= not b or a;
    layer8_outputs(3437) <= a;
    layer8_outputs(3438) <= not a;
    layer8_outputs(3439) <= not b or a;
    layer8_outputs(3440) <= not a;
    layer8_outputs(3441) <= a;
    layer8_outputs(3442) <= b;
    layer8_outputs(3443) <= not a or b;
    layer8_outputs(3444) <= b and not a;
    layer8_outputs(3445) <= a and not b;
    layer8_outputs(3446) <= a and b;
    layer8_outputs(3447) <= not (a xor b);
    layer8_outputs(3448) <= not b;
    layer8_outputs(3449) <= a and b;
    layer8_outputs(3450) <= a xor b;
    layer8_outputs(3451) <= not (a xor b);
    layer8_outputs(3452) <= not (a xor b);
    layer8_outputs(3453) <= not a;
    layer8_outputs(3454) <= not b;
    layer8_outputs(3455) <= a;
    layer8_outputs(3456) <= not a or b;
    layer8_outputs(3457) <= not (a or b);
    layer8_outputs(3458) <= a or b;
    layer8_outputs(3459) <= a or b;
    layer8_outputs(3460) <= not (a xor b);
    layer8_outputs(3461) <= not a;
    layer8_outputs(3462) <= not a or b;
    layer8_outputs(3463) <= b and not a;
    layer8_outputs(3464) <= not (a xor b);
    layer8_outputs(3465) <= not b or a;
    layer8_outputs(3466) <= a or b;
    layer8_outputs(3467) <= not (a xor b);
    layer8_outputs(3468) <= a and b;
    layer8_outputs(3469) <= not (a and b);
    layer8_outputs(3470) <= a or b;
    layer8_outputs(3471) <= a;
    layer8_outputs(3472) <= '1';
    layer8_outputs(3473) <= not b;
    layer8_outputs(3474) <= not a or b;
    layer8_outputs(3475) <= not b;
    layer8_outputs(3476) <= not a or b;
    layer8_outputs(3477) <= a xor b;
    layer8_outputs(3478) <= not a;
    layer8_outputs(3479) <= not a;
    layer8_outputs(3480) <= not b;
    layer8_outputs(3481) <= not (a xor b);
    layer8_outputs(3482) <= not a or b;
    layer8_outputs(3483) <= not b or a;
    layer8_outputs(3484) <= not (a xor b);
    layer8_outputs(3485) <= not b or a;
    layer8_outputs(3486) <= not (a and b);
    layer8_outputs(3487) <= not b;
    layer8_outputs(3488) <= not a or b;
    layer8_outputs(3489) <= b and not a;
    layer8_outputs(3490) <= a xor b;
    layer8_outputs(3491) <= a xor b;
    layer8_outputs(3492) <= a xor b;
    layer8_outputs(3493) <= a;
    layer8_outputs(3494) <= a or b;
    layer8_outputs(3495) <= a;
    layer8_outputs(3496) <= not a or b;
    layer8_outputs(3497) <= not (a and b);
    layer8_outputs(3498) <= not (a xor b);
    layer8_outputs(3499) <= not a;
    layer8_outputs(3500) <= not b;
    layer8_outputs(3501) <= b;
    layer8_outputs(3502) <= not a;
    layer8_outputs(3503) <= b;
    layer8_outputs(3504) <= not (a xor b);
    layer8_outputs(3505) <= a xor b;
    layer8_outputs(3506) <= not b;
    layer8_outputs(3507) <= a xor b;
    layer8_outputs(3508) <= not a;
    layer8_outputs(3509) <= not (a xor b);
    layer8_outputs(3510) <= b;
    layer8_outputs(3511) <= not a;
    layer8_outputs(3512) <= a;
    layer8_outputs(3513) <= not (a and b);
    layer8_outputs(3514) <= a;
    layer8_outputs(3515) <= b;
    layer8_outputs(3516) <= not a;
    layer8_outputs(3517) <= not a;
    layer8_outputs(3518) <= not (a xor b);
    layer8_outputs(3519) <= not (a or b);
    layer8_outputs(3520) <= not b or a;
    layer8_outputs(3521) <= not (a and b);
    layer8_outputs(3522) <= b;
    layer8_outputs(3523) <= a xor b;
    layer8_outputs(3524) <= not (a xor b);
    layer8_outputs(3525) <= a xor b;
    layer8_outputs(3526) <= a;
    layer8_outputs(3527) <= not b;
    layer8_outputs(3528) <= not a;
    layer8_outputs(3529) <= a;
    layer8_outputs(3530) <= a;
    layer8_outputs(3531) <= a or b;
    layer8_outputs(3532) <= not a;
    layer8_outputs(3533) <= a and not b;
    layer8_outputs(3534) <= a xor b;
    layer8_outputs(3535) <= a or b;
    layer8_outputs(3536) <= a;
    layer8_outputs(3537) <= not (a or b);
    layer8_outputs(3538) <= a and b;
    layer8_outputs(3539) <= not (a xor b);
    layer8_outputs(3540) <= b;
    layer8_outputs(3541) <= not (a xor b);
    layer8_outputs(3542) <= b and not a;
    layer8_outputs(3543) <= not (a or b);
    layer8_outputs(3544) <= b;
    layer8_outputs(3545) <= not a;
    layer8_outputs(3546) <= b and not a;
    layer8_outputs(3547) <= not (a xor b);
    layer8_outputs(3548) <= not (a xor b);
    layer8_outputs(3549) <= a and not b;
    layer8_outputs(3550) <= a xor b;
    layer8_outputs(3551) <= a and b;
    layer8_outputs(3552) <= a;
    layer8_outputs(3553) <= not (a xor b);
    layer8_outputs(3554) <= a;
    layer8_outputs(3555) <= b and not a;
    layer8_outputs(3556) <= a xor b;
    layer8_outputs(3557) <= a;
    layer8_outputs(3558) <= not a;
    layer8_outputs(3559) <= b;
    layer8_outputs(3560) <= not a or b;
    layer8_outputs(3561) <= not a;
    layer8_outputs(3562) <= b and not a;
    layer8_outputs(3563) <= a;
    layer8_outputs(3564) <= not (a or b);
    layer8_outputs(3565) <= not (a or b);
    layer8_outputs(3566) <= b;
    layer8_outputs(3567) <= not a;
    layer8_outputs(3568) <= not b;
    layer8_outputs(3569) <= not b;
    layer8_outputs(3570) <= b;
    layer8_outputs(3571) <= a;
    layer8_outputs(3572) <= a or b;
    layer8_outputs(3573) <= a and not b;
    layer8_outputs(3574) <= a and b;
    layer8_outputs(3575) <= not (a or b);
    layer8_outputs(3576) <= a xor b;
    layer8_outputs(3577) <= b and not a;
    layer8_outputs(3578) <= not a;
    layer8_outputs(3579) <= not a or b;
    layer8_outputs(3580) <= not a or b;
    layer8_outputs(3581) <= a and b;
    layer8_outputs(3582) <= a and b;
    layer8_outputs(3583) <= b;
    layer8_outputs(3584) <= a xor b;
    layer8_outputs(3585) <= b;
    layer8_outputs(3586) <= b;
    layer8_outputs(3587) <= a;
    layer8_outputs(3588) <= not (a or b);
    layer8_outputs(3589) <= b and not a;
    layer8_outputs(3590) <= b;
    layer8_outputs(3591) <= not b;
    layer8_outputs(3592) <= a and b;
    layer8_outputs(3593) <= a or b;
    layer8_outputs(3594) <= not (a and b);
    layer8_outputs(3595) <= b and not a;
    layer8_outputs(3596) <= a or b;
    layer8_outputs(3597) <= not b;
    layer8_outputs(3598) <= not b or a;
    layer8_outputs(3599) <= a xor b;
    layer8_outputs(3600) <= not (a and b);
    layer8_outputs(3601) <= not (a xor b);
    layer8_outputs(3602) <= not a;
    layer8_outputs(3603) <= not (a xor b);
    layer8_outputs(3604) <= a xor b;
    layer8_outputs(3605) <= b;
    layer8_outputs(3606) <= not b;
    layer8_outputs(3607) <= a xor b;
    layer8_outputs(3608) <= a and b;
    layer8_outputs(3609) <= not b;
    layer8_outputs(3610) <= not a;
    layer8_outputs(3611) <= not b;
    layer8_outputs(3612) <= not (a xor b);
    layer8_outputs(3613) <= not b;
    layer8_outputs(3614) <= a xor b;
    layer8_outputs(3615) <= b;
    layer8_outputs(3616) <= not b;
    layer8_outputs(3617) <= not (a or b);
    layer8_outputs(3618) <= not b;
    layer8_outputs(3619) <= a xor b;
    layer8_outputs(3620) <= not a or b;
    layer8_outputs(3621) <= b and not a;
    layer8_outputs(3622) <= not (a xor b);
    layer8_outputs(3623) <= a;
    layer8_outputs(3624) <= not (a and b);
    layer8_outputs(3625) <= not (a xor b);
    layer8_outputs(3626) <= a or b;
    layer8_outputs(3627) <= a xor b;
    layer8_outputs(3628) <= a xor b;
    layer8_outputs(3629) <= not (a xor b);
    layer8_outputs(3630) <= a;
    layer8_outputs(3631) <= not (a and b);
    layer8_outputs(3632) <= not a;
    layer8_outputs(3633) <= a and b;
    layer8_outputs(3634) <= b;
    layer8_outputs(3635) <= b and not a;
    layer8_outputs(3636) <= not (a xor b);
    layer8_outputs(3637) <= not b;
    layer8_outputs(3638) <= not (a and b);
    layer8_outputs(3639) <= not b;
    layer8_outputs(3640) <= not a;
    layer8_outputs(3641) <= not b;
    layer8_outputs(3642) <= not a;
    layer8_outputs(3643) <= not (a xor b);
    layer8_outputs(3644) <= not b;
    layer8_outputs(3645) <= a;
    layer8_outputs(3646) <= not a;
    layer8_outputs(3647) <= not (a or b);
    layer8_outputs(3648) <= a;
    layer8_outputs(3649) <= b and not a;
    layer8_outputs(3650) <= not b;
    layer8_outputs(3651) <= b and not a;
    layer8_outputs(3652) <= a and not b;
    layer8_outputs(3653) <= not (a and b);
    layer8_outputs(3654) <= not b;
    layer8_outputs(3655) <= a and not b;
    layer8_outputs(3656) <= a xor b;
    layer8_outputs(3657) <= not (a or b);
    layer8_outputs(3658) <= b;
    layer8_outputs(3659) <= b;
    layer8_outputs(3660) <= a;
    layer8_outputs(3661) <= not a;
    layer8_outputs(3662) <= not a or b;
    layer8_outputs(3663) <= not a;
    layer8_outputs(3664) <= not b or a;
    layer8_outputs(3665) <= not b or a;
    layer8_outputs(3666) <= not (a or b);
    layer8_outputs(3667) <= not (a xor b);
    layer8_outputs(3668) <= not (a xor b);
    layer8_outputs(3669) <= not b;
    layer8_outputs(3670) <= not (a xor b);
    layer8_outputs(3671) <= a;
    layer8_outputs(3672) <= a xor b;
    layer8_outputs(3673) <= a;
    layer8_outputs(3674) <= not (a and b);
    layer8_outputs(3675) <= not b;
    layer8_outputs(3676) <= not a;
    layer8_outputs(3677) <= not (a and b);
    layer8_outputs(3678) <= a xor b;
    layer8_outputs(3679) <= not a;
    layer8_outputs(3680) <= not b or a;
    layer8_outputs(3681) <= b;
    layer8_outputs(3682) <= a;
    layer8_outputs(3683) <= a;
    layer8_outputs(3684) <= not b;
    layer8_outputs(3685) <= not b;
    layer8_outputs(3686) <= a xor b;
    layer8_outputs(3687) <= a xor b;
    layer8_outputs(3688) <= a;
    layer8_outputs(3689) <= not (a and b);
    layer8_outputs(3690) <= not (a or b);
    layer8_outputs(3691) <= not a or b;
    layer8_outputs(3692) <= not (a xor b);
    layer8_outputs(3693) <= not (a xor b);
    layer8_outputs(3694) <= a xor b;
    layer8_outputs(3695) <= not b;
    layer8_outputs(3696) <= b;
    layer8_outputs(3697) <= b;
    layer8_outputs(3698) <= b;
    layer8_outputs(3699) <= not b;
    layer8_outputs(3700) <= a xor b;
    layer8_outputs(3701) <= not b;
    layer8_outputs(3702) <= not a;
    layer8_outputs(3703) <= not b;
    layer8_outputs(3704) <= not (a xor b);
    layer8_outputs(3705) <= not (a and b);
    layer8_outputs(3706) <= not a;
    layer8_outputs(3707) <= a xor b;
    layer8_outputs(3708) <= not b;
    layer8_outputs(3709) <= not b;
    layer8_outputs(3710) <= not b;
    layer8_outputs(3711) <= '0';
    layer8_outputs(3712) <= not b;
    layer8_outputs(3713) <= not b;
    layer8_outputs(3714) <= a;
    layer8_outputs(3715) <= b and not a;
    layer8_outputs(3716) <= a and not b;
    layer8_outputs(3717) <= a xor b;
    layer8_outputs(3718) <= a;
    layer8_outputs(3719) <= a xor b;
    layer8_outputs(3720) <= not (a xor b);
    layer8_outputs(3721) <= a and not b;
    layer8_outputs(3722) <= not b;
    layer8_outputs(3723) <= b;
    layer8_outputs(3724) <= a;
    layer8_outputs(3725) <= a or b;
    layer8_outputs(3726) <= not b;
    layer8_outputs(3727) <= not b;
    layer8_outputs(3728) <= b;
    layer8_outputs(3729) <= a and not b;
    layer8_outputs(3730) <= b;
    layer8_outputs(3731) <= not a or b;
    layer8_outputs(3732) <= not b;
    layer8_outputs(3733) <= b and not a;
    layer8_outputs(3734) <= a and b;
    layer8_outputs(3735) <= a;
    layer8_outputs(3736) <= a and b;
    layer8_outputs(3737) <= not (a or b);
    layer8_outputs(3738) <= not (a xor b);
    layer8_outputs(3739) <= not a;
    layer8_outputs(3740) <= a;
    layer8_outputs(3741) <= a and not b;
    layer8_outputs(3742) <= not (a and b);
    layer8_outputs(3743) <= a xor b;
    layer8_outputs(3744) <= not (a xor b);
    layer8_outputs(3745) <= a and not b;
    layer8_outputs(3746) <= a xor b;
    layer8_outputs(3747) <= b;
    layer8_outputs(3748) <= b and not a;
    layer8_outputs(3749) <= not b or a;
    layer8_outputs(3750) <= a xor b;
    layer8_outputs(3751) <= not (a xor b);
    layer8_outputs(3752) <= b;
    layer8_outputs(3753) <= not b;
    layer8_outputs(3754) <= a xor b;
    layer8_outputs(3755) <= not (a xor b);
    layer8_outputs(3756) <= not (a or b);
    layer8_outputs(3757) <= a and not b;
    layer8_outputs(3758) <= a;
    layer8_outputs(3759) <= not (a xor b);
    layer8_outputs(3760) <= not (a or b);
    layer8_outputs(3761) <= a or b;
    layer8_outputs(3762) <= not a;
    layer8_outputs(3763) <= not (a xor b);
    layer8_outputs(3764) <= b and not a;
    layer8_outputs(3765) <= not a;
    layer8_outputs(3766) <= a xor b;
    layer8_outputs(3767) <= not a;
    layer8_outputs(3768) <= not b;
    layer8_outputs(3769) <= a;
    layer8_outputs(3770) <= not a or b;
    layer8_outputs(3771) <= b and not a;
    layer8_outputs(3772) <= not b;
    layer8_outputs(3773) <= b;
    layer8_outputs(3774) <= not a;
    layer8_outputs(3775) <= not a or b;
    layer8_outputs(3776) <= not (a or b);
    layer8_outputs(3777) <= not b;
    layer8_outputs(3778) <= not (a or b);
    layer8_outputs(3779) <= not b;
    layer8_outputs(3780) <= a and not b;
    layer8_outputs(3781) <= a and b;
    layer8_outputs(3782) <= a or b;
    layer8_outputs(3783) <= not (a and b);
    layer8_outputs(3784) <= not (a xor b);
    layer8_outputs(3785) <= not (a or b);
    layer8_outputs(3786) <= a xor b;
    layer8_outputs(3787) <= not (a xor b);
    layer8_outputs(3788) <= b;
    layer8_outputs(3789) <= not b;
    layer8_outputs(3790) <= not b;
    layer8_outputs(3791) <= not a;
    layer8_outputs(3792) <= a;
    layer8_outputs(3793) <= not a;
    layer8_outputs(3794) <= not a;
    layer8_outputs(3795) <= a or b;
    layer8_outputs(3796) <= not b or a;
    layer8_outputs(3797) <= a xor b;
    layer8_outputs(3798) <= not b;
    layer8_outputs(3799) <= a xor b;
    layer8_outputs(3800) <= not a;
    layer8_outputs(3801) <= a xor b;
    layer8_outputs(3802) <= a;
    layer8_outputs(3803) <= a;
    layer8_outputs(3804) <= a and not b;
    layer8_outputs(3805) <= b;
    layer8_outputs(3806) <= b;
    layer8_outputs(3807) <= not b;
    layer8_outputs(3808) <= a xor b;
    layer8_outputs(3809) <= not b;
    layer8_outputs(3810) <= not a or b;
    layer8_outputs(3811) <= not a;
    layer8_outputs(3812) <= not (a xor b);
    layer8_outputs(3813) <= not (a and b);
    layer8_outputs(3814) <= not b or a;
    layer8_outputs(3815) <= b;
    layer8_outputs(3816) <= not a;
    layer8_outputs(3817) <= not a;
    layer8_outputs(3818) <= b;
    layer8_outputs(3819) <= not b or a;
    layer8_outputs(3820) <= a;
    layer8_outputs(3821) <= a;
    layer8_outputs(3822) <= b and not a;
    layer8_outputs(3823) <= not a;
    layer8_outputs(3824) <= not (a xor b);
    layer8_outputs(3825) <= a;
    layer8_outputs(3826) <= a or b;
    layer8_outputs(3827) <= a xor b;
    layer8_outputs(3828) <= not (a and b);
    layer8_outputs(3829) <= not (a xor b);
    layer8_outputs(3830) <= a and not b;
    layer8_outputs(3831) <= not (a or b);
    layer8_outputs(3832) <= a;
    layer8_outputs(3833) <= b and not a;
    layer8_outputs(3834) <= a and b;
    layer8_outputs(3835) <= not b or a;
    layer8_outputs(3836) <= b;
    layer8_outputs(3837) <= not b;
    layer8_outputs(3838) <= a xor b;
    layer8_outputs(3839) <= not a or b;
    layer8_outputs(3840) <= a and not b;
    layer8_outputs(3841) <= not b or a;
    layer8_outputs(3842) <= '0';
    layer8_outputs(3843) <= a;
    layer8_outputs(3844) <= not (a xor b);
    layer8_outputs(3845) <= a xor b;
    layer8_outputs(3846) <= not a;
    layer8_outputs(3847) <= not a;
    layer8_outputs(3848) <= b;
    layer8_outputs(3849) <= b and not a;
    layer8_outputs(3850) <= not b;
    layer8_outputs(3851) <= not b;
    layer8_outputs(3852) <= a;
    layer8_outputs(3853) <= not (a xor b);
    layer8_outputs(3854) <= not a;
    layer8_outputs(3855) <= a;
    layer8_outputs(3856) <= not a;
    layer8_outputs(3857) <= b;
    layer8_outputs(3858) <= a;
    layer8_outputs(3859) <= b and not a;
    layer8_outputs(3860) <= not a;
    layer8_outputs(3861) <= not (a and b);
    layer8_outputs(3862) <= not a or b;
    layer8_outputs(3863) <= a and b;
    layer8_outputs(3864) <= a;
    layer8_outputs(3865) <= not (a xor b);
    layer8_outputs(3866) <= a and not b;
    layer8_outputs(3867) <= not a;
    layer8_outputs(3868) <= not (a xor b);
    layer8_outputs(3869) <= a;
    layer8_outputs(3870) <= b;
    layer8_outputs(3871) <= a;
    layer8_outputs(3872) <= b;
    layer8_outputs(3873) <= not b;
    layer8_outputs(3874) <= a;
    layer8_outputs(3875) <= not (a xor b);
    layer8_outputs(3876) <= a;
    layer8_outputs(3877) <= not (a xor b);
    layer8_outputs(3878) <= not (a xor b);
    layer8_outputs(3879) <= not (a xor b);
    layer8_outputs(3880) <= not a;
    layer8_outputs(3881) <= a and not b;
    layer8_outputs(3882) <= not b;
    layer8_outputs(3883) <= not b;
    layer8_outputs(3884) <= a xor b;
    layer8_outputs(3885) <= b;
    layer8_outputs(3886) <= not (a and b);
    layer8_outputs(3887) <= b;
    layer8_outputs(3888) <= b;
    layer8_outputs(3889) <= a or b;
    layer8_outputs(3890) <= not b;
    layer8_outputs(3891) <= a xor b;
    layer8_outputs(3892) <= not b or a;
    layer8_outputs(3893) <= b;
    layer8_outputs(3894) <= a xor b;
    layer8_outputs(3895) <= not a or b;
    layer8_outputs(3896) <= not (a and b);
    layer8_outputs(3897) <= not a;
    layer8_outputs(3898) <= not a or b;
    layer8_outputs(3899) <= not b;
    layer8_outputs(3900) <= not b;
    layer8_outputs(3901) <= a xor b;
    layer8_outputs(3902) <= a xor b;
    layer8_outputs(3903) <= not b or a;
    layer8_outputs(3904) <= not (a and b);
    layer8_outputs(3905) <= not a or b;
    layer8_outputs(3906) <= not (a xor b);
    layer8_outputs(3907) <= not (a or b);
    layer8_outputs(3908) <= not (a xor b);
    layer8_outputs(3909) <= b;
    layer8_outputs(3910) <= a;
    layer8_outputs(3911) <= a and not b;
    layer8_outputs(3912) <= a;
    layer8_outputs(3913) <= a;
    layer8_outputs(3914) <= not (a or b);
    layer8_outputs(3915) <= a;
    layer8_outputs(3916) <= a xor b;
    layer8_outputs(3917) <= b;
    layer8_outputs(3918) <= a and b;
    layer8_outputs(3919) <= a and b;
    layer8_outputs(3920) <= not (a xor b);
    layer8_outputs(3921) <= b;
    layer8_outputs(3922) <= a and b;
    layer8_outputs(3923) <= not b;
    layer8_outputs(3924) <= not (a and b);
    layer8_outputs(3925) <= not (a and b);
    layer8_outputs(3926) <= a xor b;
    layer8_outputs(3927) <= not b;
    layer8_outputs(3928) <= b and not a;
    layer8_outputs(3929) <= a;
    layer8_outputs(3930) <= a and b;
    layer8_outputs(3931) <= not b or a;
    layer8_outputs(3932) <= a;
    layer8_outputs(3933) <= not (a or b);
    layer8_outputs(3934) <= a;
    layer8_outputs(3935) <= not a;
    layer8_outputs(3936) <= a and not b;
    layer8_outputs(3937) <= a;
    layer8_outputs(3938) <= not b;
    layer8_outputs(3939) <= not (a and b);
    layer8_outputs(3940) <= a;
    layer8_outputs(3941) <= b;
    layer8_outputs(3942) <= not b or a;
    layer8_outputs(3943) <= a and b;
    layer8_outputs(3944) <= not a;
    layer8_outputs(3945) <= not a;
    layer8_outputs(3946) <= not b or a;
    layer8_outputs(3947) <= a xor b;
    layer8_outputs(3948) <= a xor b;
    layer8_outputs(3949) <= not (a xor b);
    layer8_outputs(3950) <= not b or a;
    layer8_outputs(3951) <= b and not a;
    layer8_outputs(3952) <= a or b;
    layer8_outputs(3953) <= not b;
    layer8_outputs(3954) <= b;
    layer8_outputs(3955) <= not b or a;
    layer8_outputs(3956) <= a xor b;
    layer8_outputs(3957) <= not a;
    layer8_outputs(3958) <= a and b;
    layer8_outputs(3959) <= a or b;
    layer8_outputs(3960) <= not (a or b);
    layer8_outputs(3961) <= not b;
    layer8_outputs(3962) <= not (a xor b);
    layer8_outputs(3963) <= not b;
    layer8_outputs(3964) <= b;
    layer8_outputs(3965) <= a;
    layer8_outputs(3966) <= not (a xor b);
    layer8_outputs(3967) <= not (a and b);
    layer8_outputs(3968) <= not b;
    layer8_outputs(3969) <= not b;
    layer8_outputs(3970) <= a xor b;
    layer8_outputs(3971) <= a xor b;
    layer8_outputs(3972) <= not (a xor b);
    layer8_outputs(3973) <= a and not b;
    layer8_outputs(3974) <= a and b;
    layer8_outputs(3975) <= not a;
    layer8_outputs(3976) <= not (a or b);
    layer8_outputs(3977) <= not (a xor b);
    layer8_outputs(3978) <= a xor b;
    layer8_outputs(3979) <= a;
    layer8_outputs(3980) <= not (a or b);
    layer8_outputs(3981) <= a or b;
    layer8_outputs(3982) <= not b;
    layer8_outputs(3983) <= a xor b;
    layer8_outputs(3984) <= a xor b;
    layer8_outputs(3985) <= a and b;
    layer8_outputs(3986) <= a xor b;
    layer8_outputs(3987) <= not b or a;
    layer8_outputs(3988) <= not (a and b);
    layer8_outputs(3989) <= a;
    layer8_outputs(3990) <= a and b;
    layer8_outputs(3991) <= not b or a;
    layer8_outputs(3992) <= not b;
    layer8_outputs(3993) <= b and not a;
    layer8_outputs(3994) <= a;
    layer8_outputs(3995) <= b;
    layer8_outputs(3996) <= not (a xor b);
    layer8_outputs(3997) <= a and b;
    layer8_outputs(3998) <= a xor b;
    layer8_outputs(3999) <= not b or a;
    layer8_outputs(4000) <= a xor b;
    layer8_outputs(4001) <= not b;
    layer8_outputs(4002) <= a;
    layer8_outputs(4003) <= a;
    layer8_outputs(4004) <= not (a xor b);
    layer8_outputs(4005) <= b and not a;
    layer8_outputs(4006) <= not (a and b);
    layer8_outputs(4007) <= not (a xor b);
    layer8_outputs(4008) <= not b;
    layer8_outputs(4009) <= not a;
    layer8_outputs(4010) <= a and not b;
    layer8_outputs(4011) <= not (a xor b);
    layer8_outputs(4012) <= not b;
    layer8_outputs(4013) <= not (a xor b);
    layer8_outputs(4014) <= b;
    layer8_outputs(4015) <= not (a xor b);
    layer8_outputs(4016) <= not a;
    layer8_outputs(4017) <= a;
    layer8_outputs(4018) <= b;
    layer8_outputs(4019) <= a;
    layer8_outputs(4020) <= b;
    layer8_outputs(4021) <= not a or b;
    layer8_outputs(4022) <= not (a and b);
    layer8_outputs(4023) <= not a or b;
    layer8_outputs(4024) <= b;
    layer8_outputs(4025) <= not (a xor b);
    layer8_outputs(4026) <= a xor b;
    layer8_outputs(4027) <= b;
    layer8_outputs(4028) <= not (a xor b);
    layer8_outputs(4029) <= not a;
    layer8_outputs(4030) <= a;
    layer8_outputs(4031) <= a xor b;
    layer8_outputs(4032) <= a xor b;
    layer8_outputs(4033) <= a or b;
    layer8_outputs(4034) <= a xor b;
    layer8_outputs(4035) <= a;
    layer8_outputs(4036) <= not (a or b);
    layer8_outputs(4037) <= b;
    layer8_outputs(4038) <= b;
    layer8_outputs(4039) <= not a;
    layer8_outputs(4040) <= a;
    layer8_outputs(4041) <= not (a xor b);
    layer8_outputs(4042) <= not (a xor b);
    layer8_outputs(4043) <= a;
    layer8_outputs(4044) <= a or b;
    layer8_outputs(4045) <= not (a xor b);
    layer8_outputs(4046) <= not b or a;
    layer8_outputs(4047) <= not a or b;
    layer8_outputs(4048) <= a xor b;
    layer8_outputs(4049) <= not a;
    layer8_outputs(4050) <= not a or b;
    layer8_outputs(4051) <= b;
    layer8_outputs(4052) <= not a;
    layer8_outputs(4053) <= b;
    layer8_outputs(4054) <= not b or a;
    layer8_outputs(4055) <= not a;
    layer8_outputs(4056) <= a or b;
    layer8_outputs(4057) <= not a or b;
    layer8_outputs(4058) <= not b or a;
    layer8_outputs(4059) <= b;
    layer8_outputs(4060) <= a xor b;
    layer8_outputs(4061) <= b;
    layer8_outputs(4062) <= a xor b;
    layer8_outputs(4063) <= b;
    layer8_outputs(4064) <= a;
    layer8_outputs(4065) <= not a or b;
    layer8_outputs(4066) <= not b;
    layer8_outputs(4067) <= a and b;
    layer8_outputs(4068) <= a xor b;
    layer8_outputs(4069) <= a or b;
    layer8_outputs(4070) <= a and not b;
    layer8_outputs(4071) <= a and b;
    layer8_outputs(4072) <= not (a and b);
    layer8_outputs(4073) <= not (a or b);
    layer8_outputs(4074) <= a;
    layer8_outputs(4075) <= a or b;
    layer8_outputs(4076) <= not a;
    layer8_outputs(4077) <= not b;
    layer8_outputs(4078) <= not (a xor b);
    layer8_outputs(4079) <= a or b;
    layer8_outputs(4080) <= a;
    layer8_outputs(4081) <= a xor b;
    layer8_outputs(4082) <= not b;
    layer8_outputs(4083) <= b;
    layer8_outputs(4084) <= not (a xor b);
    layer8_outputs(4085) <= not a;
    layer8_outputs(4086) <= a xor b;
    layer8_outputs(4087) <= not (a and b);
    layer8_outputs(4088) <= not (a xor b);
    layer8_outputs(4089) <= a and not b;
    layer8_outputs(4090) <= not a;
    layer8_outputs(4091) <= not (a xor b);
    layer8_outputs(4092) <= not (a xor b);
    layer8_outputs(4093) <= not b or a;
    layer8_outputs(4094) <= not a;
    layer8_outputs(4095) <= not a;
    layer8_outputs(4096) <= a and not b;
    layer8_outputs(4097) <= a or b;
    layer8_outputs(4098) <= not (a xor b);
    layer8_outputs(4099) <= not b;
    layer8_outputs(4100) <= not a or b;
    layer8_outputs(4101) <= a xor b;
    layer8_outputs(4102) <= a xor b;
    layer8_outputs(4103) <= b and not a;
    layer8_outputs(4104) <= not (a xor b);
    layer8_outputs(4105) <= a and b;
    layer8_outputs(4106) <= b and not a;
    layer8_outputs(4107) <= a xor b;
    layer8_outputs(4108) <= a xor b;
    layer8_outputs(4109) <= b and not a;
    layer8_outputs(4110) <= not (a and b);
    layer8_outputs(4111) <= not (a or b);
    layer8_outputs(4112) <= a and not b;
    layer8_outputs(4113) <= a or b;
    layer8_outputs(4114) <= not (a xor b);
    layer8_outputs(4115) <= b;
    layer8_outputs(4116) <= a xor b;
    layer8_outputs(4117) <= a xor b;
    layer8_outputs(4118) <= a and b;
    layer8_outputs(4119) <= not (a or b);
    layer8_outputs(4120) <= a;
    layer8_outputs(4121) <= a and not b;
    layer8_outputs(4122) <= not a;
    layer8_outputs(4123) <= not (a and b);
    layer8_outputs(4124) <= not a;
    layer8_outputs(4125) <= not a;
    layer8_outputs(4126) <= '0';
    layer8_outputs(4127) <= a;
    layer8_outputs(4128) <= b;
    layer8_outputs(4129) <= not (a and b);
    layer8_outputs(4130) <= a;
    layer8_outputs(4131) <= a or b;
    layer8_outputs(4132) <= not b;
    layer8_outputs(4133) <= a xor b;
    layer8_outputs(4134) <= a and not b;
    layer8_outputs(4135) <= not (a xor b);
    layer8_outputs(4136) <= a;
    layer8_outputs(4137) <= not b or a;
    layer8_outputs(4138) <= a xor b;
    layer8_outputs(4139) <= a xor b;
    layer8_outputs(4140) <= not (a xor b);
    layer8_outputs(4141) <= not (a xor b);
    layer8_outputs(4142) <= a;
    layer8_outputs(4143) <= not (a xor b);
    layer8_outputs(4144) <= not (a or b);
    layer8_outputs(4145) <= a;
    layer8_outputs(4146) <= not a or b;
    layer8_outputs(4147) <= a or b;
    layer8_outputs(4148) <= not a;
    layer8_outputs(4149) <= b and not a;
    layer8_outputs(4150) <= a and not b;
    layer8_outputs(4151) <= b and not a;
    layer8_outputs(4152) <= not (a xor b);
    layer8_outputs(4153) <= a;
    layer8_outputs(4154) <= not b;
    layer8_outputs(4155) <= not a;
    layer8_outputs(4156) <= not a;
    layer8_outputs(4157) <= a xor b;
    layer8_outputs(4158) <= a xor b;
    layer8_outputs(4159) <= a;
    layer8_outputs(4160) <= a or b;
    layer8_outputs(4161) <= not a;
    layer8_outputs(4162) <= b and not a;
    layer8_outputs(4163) <= not b or a;
    layer8_outputs(4164) <= a and not b;
    layer8_outputs(4165) <= a xor b;
    layer8_outputs(4166) <= a;
    layer8_outputs(4167) <= a xor b;
    layer8_outputs(4168) <= not b;
    layer8_outputs(4169) <= b and not a;
    layer8_outputs(4170) <= not b;
    layer8_outputs(4171) <= a and not b;
    layer8_outputs(4172) <= not a;
    layer8_outputs(4173) <= not (a xor b);
    layer8_outputs(4174) <= not a;
    layer8_outputs(4175) <= not b;
    layer8_outputs(4176) <= not a;
    layer8_outputs(4177) <= not (a and b);
    layer8_outputs(4178) <= b;
    layer8_outputs(4179) <= not b or a;
    layer8_outputs(4180) <= a and b;
    layer8_outputs(4181) <= b;
    layer8_outputs(4182) <= a and b;
    layer8_outputs(4183) <= b;
    layer8_outputs(4184) <= b;
    layer8_outputs(4185) <= not b;
    layer8_outputs(4186) <= a xor b;
    layer8_outputs(4187) <= a;
    layer8_outputs(4188) <= a and b;
    layer8_outputs(4189) <= a;
    layer8_outputs(4190) <= not (a and b);
    layer8_outputs(4191) <= not (a xor b);
    layer8_outputs(4192) <= a and b;
    layer8_outputs(4193) <= not (a or b);
    layer8_outputs(4194) <= a or b;
    layer8_outputs(4195) <= '1';
    layer8_outputs(4196) <= not a or b;
    layer8_outputs(4197) <= not (a xor b);
    layer8_outputs(4198) <= '0';
    layer8_outputs(4199) <= a xor b;
    layer8_outputs(4200) <= not (a or b);
    layer8_outputs(4201) <= b;
    layer8_outputs(4202) <= not b;
    layer8_outputs(4203) <= a xor b;
    layer8_outputs(4204) <= not (a and b);
    layer8_outputs(4205) <= a or b;
    layer8_outputs(4206) <= not (a or b);
    layer8_outputs(4207) <= b;
    layer8_outputs(4208) <= not b;
    layer8_outputs(4209) <= not (a xor b);
    layer8_outputs(4210) <= a or b;
    layer8_outputs(4211) <= not (a xor b);
    layer8_outputs(4212) <= not b;
    layer8_outputs(4213) <= not b;
    layer8_outputs(4214) <= b;
    layer8_outputs(4215) <= b;
    layer8_outputs(4216) <= not a;
    layer8_outputs(4217) <= not (a xor b);
    layer8_outputs(4218) <= b;
    layer8_outputs(4219) <= not (a or b);
    layer8_outputs(4220) <= b and not a;
    layer8_outputs(4221) <= not a;
    layer8_outputs(4222) <= not b;
    layer8_outputs(4223) <= b;
    layer8_outputs(4224) <= a or b;
    layer8_outputs(4225) <= '0';
    layer8_outputs(4226) <= a;
    layer8_outputs(4227) <= a xor b;
    layer8_outputs(4228) <= a;
    layer8_outputs(4229) <= a and not b;
    layer8_outputs(4230) <= not a;
    layer8_outputs(4231) <= b;
    layer8_outputs(4232) <= a xor b;
    layer8_outputs(4233) <= a xor b;
    layer8_outputs(4234) <= '1';
    layer8_outputs(4235) <= b and not a;
    layer8_outputs(4236) <= not a or b;
    layer8_outputs(4237) <= not a;
    layer8_outputs(4238) <= a;
    layer8_outputs(4239) <= b and not a;
    layer8_outputs(4240) <= a;
    layer8_outputs(4241) <= a xor b;
    layer8_outputs(4242) <= not (a or b);
    layer8_outputs(4243) <= b;
    layer8_outputs(4244) <= a;
    layer8_outputs(4245) <= not a;
    layer8_outputs(4246) <= a;
    layer8_outputs(4247) <= a;
    layer8_outputs(4248) <= not b or a;
    layer8_outputs(4249) <= not (a xor b);
    layer8_outputs(4250) <= a;
    layer8_outputs(4251) <= not b or a;
    layer8_outputs(4252) <= a;
    layer8_outputs(4253) <= not a;
    layer8_outputs(4254) <= not (a or b);
    layer8_outputs(4255) <= not b;
    layer8_outputs(4256) <= a or b;
    layer8_outputs(4257) <= not (a xor b);
    layer8_outputs(4258) <= not b;
    layer8_outputs(4259) <= b;
    layer8_outputs(4260) <= not (a xor b);
    layer8_outputs(4261) <= not b;
    layer8_outputs(4262) <= not a;
    layer8_outputs(4263) <= a and b;
    layer8_outputs(4264) <= a and b;
    layer8_outputs(4265) <= a xor b;
    layer8_outputs(4266) <= not a or b;
    layer8_outputs(4267) <= a and not b;
    layer8_outputs(4268) <= a and b;
    layer8_outputs(4269) <= b;
    layer8_outputs(4270) <= not b or a;
    layer8_outputs(4271) <= b and not a;
    layer8_outputs(4272) <= not b;
    layer8_outputs(4273) <= not b or a;
    layer8_outputs(4274) <= a and not b;
    layer8_outputs(4275) <= a;
    layer8_outputs(4276) <= b;
    layer8_outputs(4277) <= not b or a;
    layer8_outputs(4278) <= not a;
    layer8_outputs(4279) <= not b;
    layer8_outputs(4280) <= not b;
    layer8_outputs(4281) <= not (a xor b);
    layer8_outputs(4282) <= a;
    layer8_outputs(4283) <= a xor b;
    layer8_outputs(4284) <= a or b;
    layer8_outputs(4285) <= a and not b;
    layer8_outputs(4286) <= not b;
    layer8_outputs(4287) <= not b;
    layer8_outputs(4288) <= not (a xor b);
    layer8_outputs(4289) <= b;
    layer8_outputs(4290) <= a or b;
    layer8_outputs(4291) <= b;
    layer8_outputs(4292) <= not a;
    layer8_outputs(4293) <= b;
    layer8_outputs(4294) <= a and b;
    layer8_outputs(4295) <= b;
    layer8_outputs(4296) <= a xor b;
    layer8_outputs(4297) <= b and not a;
    layer8_outputs(4298) <= not b;
    layer8_outputs(4299) <= not a;
    layer8_outputs(4300) <= b;
    layer8_outputs(4301) <= not a;
    layer8_outputs(4302) <= not (a xor b);
    layer8_outputs(4303) <= not (a xor b);
    layer8_outputs(4304) <= a;
    layer8_outputs(4305) <= not (a xor b);
    layer8_outputs(4306) <= not b or a;
    layer8_outputs(4307) <= a;
    layer8_outputs(4308) <= not a;
    layer8_outputs(4309) <= b;
    layer8_outputs(4310) <= not b;
    layer8_outputs(4311) <= not (a xor b);
    layer8_outputs(4312) <= b;
    layer8_outputs(4313) <= a xor b;
    layer8_outputs(4314) <= a xor b;
    layer8_outputs(4315) <= b and not a;
    layer8_outputs(4316) <= a;
    layer8_outputs(4317) <= a;
    layer8_outputs(4318) <= b and not a;
    layer8_outputs(4319) <= a xor b;
    layer8_outputs(4320) <= a xor b;
    layer8_outputs(4321) <= not a;
    layer8_outputs(4322) <= b;
    layer8_outputs(4323) <= not (a xor b);
    layer8_outputs(4324) <= not b or a;
    layer8_outputs(4325) <= a or b;
    layer8_outputs(4326) <= a;
    layer8_outputs(4327) <= not (a xor b);
    layer8_outputs(4328) <= b;
    layer8_outputs(4329) <= not a;
    layer8_outputs(4330) <= b;
    layer8_outputs(4331) <= not (a or b);
    layer8_outputs(4332) <= not b;
    layer8_outputs(4333) <= a;
    layer8_outputs(4334) <= not (a or b);
    layer8_outputs(4335) <= b;
    layer8_outputs(4336) <= not a;
    layer8_outputs(4337) <= not (a xor b);
    layer8_outputs(4338) <= a and not b;
    layer8_outputs(4339) <= not b;
    layer8_outputs(4340) <= not a;
    layer8_outputs(4341) <= b;
    layer8_outputs(4342) <= not (a xor b);
    layer8_outputs(4343) <= b;
    layer8_outputs(4344) <= not b;
    layer8_outputs(4345) <= a xor b;
    layer8_outputs(4346) <= not a;
    layer8_outputs(4347) <= a;
    layer8_outputs(4348) <= not (a xor b);
    layer8_outputs(4349) <= not a;
    layer8_outputs(4350) <= a and not b;
    layer8_outputs(4351) <= not a;
    layer8_outputs(4352) <= not b;
    layer8_outputs(4353) <= a and not b;
    layer8_outputs(4354) <= not a;
    layer8_outputs(4355) <= a;
    layer8_outputs(4356) <= not b;
    layer8_outputs(4357) <= not a or b;
    layer8_outputs(4358) <= a;
    layer8_outputs(4359) <= not b;
    layer8_outputs(4360) <= not (a xor b);
    layer8_outputs(4361) <= a and not b;
    layer8_outputs(4362) <= a xor b;
    layer8_outputs(4363) <= a xor b;
    layer8_outputs(4364) <= not a;
    layer8_outputs(4365) <= not (a xor b);
    layer8_outputs(4366) <= not (a xor b);
    layer8_outputs(4367) <= a or b;
    layer8_outputs(4368) <= not b;
    layer8_outputs(4369) <= not b;
    layer8_outputs(4370) <= a;
    layer8_outputs(4371) <= b;
    layer8_outputs(4372) <= b;
    layer8_outputs(4373) <= not a;
    layer8_outputs(4374) <= a or b;
    layer8_outputs(4375) <= not b;
    layer8_outputs(4376) <= a xor b;
    layer8_outputs(4377) <= a;
    layer8_outputs(4378) <= b and not a;
    layer8_outputs(4379) <= not (a and b);
    layer8_outputs(4380) <= not (a and b);
    layer8_outputs(4381) <= not a or b;
    layer8_outputs(4382) <= not b;
    layer8_outputs(4383) <= not (a and b);
    layer8_outputs(4384) <= not a;
    layer8_outputs(4385) <= not b;
    layer8_outputs(4386) <= a;
    layer8_outputs(4387) <= not b;
    layer8_outputs(4388) <= b;
    layer8_outputs(4389) <= not b;
    layer8_outputs(4390) <= a;
    layer8_outputs(4391) <= b and not a;
    layer8_outputs(4392) <= a;
    layer8_outputs(4393) <= a xor b;
    layer8_outputs(4394) <= a or b;
    layer8_outputs(4395) <= b;
    layer8_outputs(4396) <= a;
    layer8_outputs(4397) <= not (a xor b);
    layer8_outputs(4398) <= not b or a;
    layer8_outputs(4399) <= not b or a;
    layer8_outputs(4400) <= a and b;
    layer8_outputs(4401) <= not b;
    layer8_outputs(4402) <= a;
    layer8_outputs(4403) <= not a or b;
    layer8_outputs(4404) <= a and not b;
    layer8_outputs(4405) <= not (a or b);
    layer8_outputs(4406) <= not b;
    layer8_outputs(4407) <= not a;
    layer8_outputs(4408) <= not b or a;
    layer8_outputs(4409) <= not a;
    layer8_outputs(4410) <= a;
    layer8_outputs(4411) <= not (a xor b);
    layer8_outputs(4412) <= b and not a;
    layer8_outputs(4413) <= not (a or b);
    layer8_outputs(4414) <= b;
    layer8_outputs(4415) <= a and b;
    layer8_outputs(4416) <= not b or a;
    layer8_outputs(4417) <= a xor b;
    layer8_outputs(4418) <= a or b;
    layer8_outputs(4419) <= not a;
    layer8_outputs(4420) <= a or b;
    layer8_outputs(4421) <= b and not a;
    layer8_outputs(4422) <= not (a or b);
    layer8_outputs(4423) <= '0';
    layer8_outputs(4424) <= not b or a;
    layer8_outputs(4425) <= not b or a;
    layer8_outputs(4426) <= not (a and b);
    layer8_outputs(4427) <= not b;
    layer8_outputs(4428) <= not b;
    layer8_outputs(4429) <= a;
    layer8_outputs(4430) <= not a;
    layer8_outputs(4431) <= a and b;
    layer8_outputs(4432) <= a;
    layer8_outputs(4433) <= a;
    layer8_outputs(4434) <= not (a and b);
    layer8_outputs(4435) <= '1';
    layer8_outputs(4436) <= b;
    layer8_outputs(4437) <= not a;
    layer8_outputs(4438) <= not a;
    layer8_outputs(4439) <= not (a and b);
    layer8_outputs(4440) <= not b or a;
    layer8_outputs(4441) <= a or b;
    layer8_outputs(4442) <= b;
    layer8_outputs(4443) <= a;
    layer8_outputs(4444) <= not (a xor b);
    layer8_outputs(4445) <= a xor b;
    layer8_outputs(4446) <= a xor b;
    layer8_outputs(4447) <= '0';
    layer8_outputs(4448) <= a xor b;
    layer8_outputs(4449) <= a xor b;
    layer8_outputs(4450) <= not (a or b);
    layer8_outputs(4451) <= not b or a;
    layer8_outputs(4452) <= a and b;
    layer8_outputs(4453) <= not b;
    layer8_outputs(4454) <= a and b;
    layer8_outputs(4455) <= b and not a;
    layer8_outputs(4456) <= '0';
    layer8_outputs(4457) <= not b;
    layer8_outputs(4458) <= not b;
    layer8_outputs(4459) <= b;
    layer8_outputs(4460) <= a or b;
    layer8_outputs(4461) <= not a;
    layer8_outputs(4462) <= not (a xor b);
    layer8_outputs(4463) <= not a or b;
    layer8_outputs(4464) <= not b;
    layer8_outputs(4465) <= not a;
    layer8_outputs(4466) <= b and not a;
    layer8_outputs(4467) <= b and not a;
    layer8_outputs(4468) <= not (a xor b);
    layer8_outputs(4469) <= a xor b;
    layer8_outputs(4470) <= not (a xor b);
    layer8_outputs(4471) <= a;
    layer8_outputs(4472) <= a and not b;
    layer8_outputs(4473) <= a or b;
    layer8_outputs(4474) <= not b;
    layer8_outputs(4475) <= not (a and b);
    layer8_outputs(4476) <= a;
    layer8_outputs(4477) <= not b;
    layer8_outputs(4478) <= not (a or b);
    layer8_outputs(4479) <= not a or b;
    layer8_outputs(4480) <= not a;
    layer8_outputs(4481) <= a;
    layer8_outputs(4482) <= a or b;
    layer8_outputs(4483) <= not b;
    layer8_outputs(4484) <= not (a xor b);
    layer8_outputs(4485) <= a or b;
    layer8_outputs(4486) <= a;
    layer8_outputs(4487) <= a or b;
    layer8_outputs(4488) <= b;
    layer8_outputs(4489) <= not (a xor b);
    layer8_outputs(4490) <= not b;
    layer8_outputs(4491) <= not a;
    layer8_outputs(4492) <= not (a xor b);
    layer8_outputs(4493) <= a;
    layer8_outputs(4494) <= '0';
    layer8_outputs(4495) <= a xor b;
    layer8_outputs(4496) <= a and b;
    layer8_outputs(4497) <= not (a xor b);
    layer8_outputs(4498) <= a xor b;
    layer8_outputs(4499) <= not a;
    layer8_outputs(4500) <= not a or b;
    layer8_outputs(4501) <= a and not b;
    layer8_outputs(4502) <= not (a xor b);
    layer8_outputs(4503) <= a or b;
    layer8_outputs(4504) <= b;
    layer8_outputs(4505) <= a;
    layer8_outputs(4506) <= a and not b;
    layer8_outputs(4507) <= not a or b;
    layer8_outputs(4508) <= a xor b;
    layer8_outputs(4509) <= not (a xor b);
    layer8_outputs(4510) <= a or b;
    layer8_outputs(4511) <= b and not a;
    layer8_outputs(4512) <= b;
    layer8_outputs(4513) <= a and not b;
    layer8_outputs(4514) <= a and b;
    layer8_outputs(4515) <= a or b;
    layer8_outputs(4516) <= not (a xor b);
    layer8_outputs(4517) <= a xor b;
    layer8_outputs(4518) <= not (a and b);
    layer8_outputs(4519) <= b;
    layer8_outputs(4520) <= a xor b;
    layer8_outputs(4521) <= not a;
    layer8_outputs(4522) <= a xor b;
    layer8_outputs(4523) <= b and not a;
    layer8_outputs(4524) <= a and not b;
    layer8_outputs(4525) <= a;
    layer8_outputs(4526) <= a xor b;
    layer8_outputs(4527) <= a and not b;
    layer8_outputs(4528) <= a and b;
    layer8_outputs(4529) <= not (a xor b);
    layer8_outputs(4530) <= b;
    layer8_outputs(4531) <= a;
    layer8_outputs(4532) <= not (a xor b);
    layer8_outputs(4533) <= not (a xor b);
    layer8_outputs(4534) <= not b or a;
    layer8_outputs(4535) <= a xor b;
    layer8_outputs(4536) <= a xor b;
    layer8_outputs(4537) <= a and b;
    layer8_outputs(4538) <= not (a xor b);
    layer8_outputs(4539) <= a;
    layer8_outputs(4540) <= a or b;
    layer8_outputs(4541) <= a;
    layer8_outputs(4542) <= b;
    layer8_outputs(4543) <= not (a xor b);
    layer8_outputs(4544) <= not a;
    layer8_outputs(4545) <= not b;
    layer8_outputs(4546) <= not (a xor b);
    layer8_outputs(4547) <= not (a and b);
    layer8_outputs(4548) <= not a;
    layer8_outputs(4549) <= not b;
    layer8_outputs(4550) <= not a;
    layer8_outputs(4551) <= b;
    layer8_outputs(4552) <= b;
    layer8_outputs(4553) <= not (a and b);
    layer8_outputs(4554) <= b;
    layer8_outputs(4555) <= not a;
    layer8_outputs(4556) <= not (a and b);
    layer8_outputs(4557) <= a xor b;
    layer8_outputs(4558) <= b;
    layer8_outputs(4559) <= '1';
    layer8_outputs(4560) <= a and b;
    layer8_outputs(4561) <= a and b;
    layer8_outputs(4562) <= not a or b;
    layer8_outputs(4563) <= not (a or b);
    layer8_outputs(4564) <= not b;
    layer8_outputs(4565) <= not (a xor b);
    layer8_outputs(4566) <= a or b;
    layer8_outputs(4567) <= b;
    layer8_outputs(4568) <= '0';
    layer8_outputs(4569) <= a and not b;
    layer8_outputs(4570) <= not (a xor b);
    layer8_outputs(4571) <= a or b;
    layer8_outputs(4572) <= not b;
    layer8_outputs(4573) <= a and b;
    layer8_outputs(4574) <= b and not a;
    layer8_outputs(4575) <= not a;
    layer8_outputs(4576) <= b;
    layer8_outputs(4577) <= a xor b;
    layer8_outputs(4578) <= a and b;
    layer8_outputs(4579) <= a xor b;
    layer8_outputs(4580) <= not (a xor b);
    layer8_outputs(4581) <= b;
    layer8_outputs(4582) <= not a;
    layer8_outputs(4583) <= not b or a;
    layer8_outputs(4584) <= b;
    layer8_outputs(4585) <= not b;
    layer8_outputs(4586) <= not a;
    layer8_outputs(4587) <= not a;
    layer8_outputs(4588) <= not (a xor b);
    layer8_outputs(4589) <= not a or b;
    layer8_outputs(4590) <= not (a or b);
    layer8_outputs(4591) <= not a or b;
    layer8_outputs(4592) <= b and not a;
    layer8_outputs(4593) <= '1';
    layer8_outputs(4594) <= a and b;
    layer8_outputs(4595) <= a;
    layer8_outputs(4596) <= b;
    layer8_outputs(4597) <= a;
    layer8_outputs(4598) <= a xor b;
    layer8_outputs(4599) <= not (a xor b);
    layer8_outputs(4600) <= a and not b;
    layer8_outputs(4601) <= '0';
    layer8_outputs(4602) <= not (a xor b);
    layer8_outputs(4603) <= not (a or b);
    layer8_outputs(4604) <= not a;
    layer8_outputs(4605) <= a;
    layer8_outputs(4606) <= not b;
    layer8_outputs(4607) <= not b;
    layer8_outputs(4608) <= a xor b;
    layer8_outputs(4609) <= not a;
    layer8_outputs(4610) <= not a or b;
    layer8_outputs(4611) <= a xor b;
    layer8_outputs(4612) <= not (a xor b);
    layer8_outputs(4613) <= not (a and b);
    layer8_outputs(4614) <= not (a xor b);
    layer8_outputs(4615) <= not (a and b);
    layer8_outputs(4616) <= not (a xor b);
    layer8_outputs(4617) <= b;
    layer8_outputs(4618) <= not (a or b);
    layer8_outputs(4619) <= a and b;
    layer8_outputs(4620) <= a or b;
    layer8_outputs(4621) <= a or b;
    layer8_outputs(4622) <= a or b;
    layer8_outputs(4623) <= not (a and b);
    layer8_outputs(4624) <= not a;
    layer8_outputs(4625) <= not b or a;
    layer8_outputs(4626) <= a or b;
    layer8_outputs(4627) <= not (a and b);
    layer8_outputs(4628) <= b;
    layer8_outputs(4629) <= not b or a;
    layer8_outputs(4630) <= a;
    layer8_outputs(4631) <= b;
    layer8_outputs(4632) <= not b;
    layer8_outputs(4633) <= not b;
    layer8_outputs(4634) <= not a;
    layer8_outputs(4635) <= b;
    layer8_outputs(4636) <= b;
    layer8_outputs(4637) <= not (a or b);
    layer8_outputs(4638) <= a;
    layer8_outputs(4639) <= not (a and b);
    layer8_outputs(4640) <= not a;
    layer8_outputs(4641) <= not (a and b);
    layer8_outputs(4642) <= not a;
    layer8_outputs(4643) <= not a or b;
    layer8_outputs(4644) <= b;
    layer8_outputs(4645) <= a xor b;
    layer8_outputs(4646) <= b and not a;
    layer8_outputs(4647) <= not b;
    layer8_outputs(4648) <= not a or b;
    layer8_outputs(4649) <= b;
    layer8_outputs(4650) <= a;
    layer8_outputs(4651) <= not b;
    layer8_outputs(4652) <= a xor b;
    layer8_outputs(4653) <= not (a and b);
    layer8_outputs(4654) <= a and not b;
    layer8_outputs(4655) <= a xor b;
    layer8_outputs(4656) <= not b;
    layer8_outputs(4657) <= b;
    layer8_outputs(4658) <= not b or a;
    layer8_outputs(4659) <= a and b;
    layer8_outputs(4660) <= not (a xor b);
    layer8_outputs(4661) <= a;
    layer8_outputs(4662) <= a;
    layer8_outputs(4663) <= not a or b;
    layer8_outputs(4664) <= not (a or b);
    layer8_outputs(4665) <= b and not a;
    layer8_outputs(4666) <= a and b;
    layer8_outputs(4667) <= a and b;
    layer8_outputs(4668) <= not a;
    layer8_outputs(4669) <= a;
    layer8_outputs(4670) <= a;
    layer8_outputs(4671) <= not b;
    layer8_outputs(4672) <= a or b;
    layer8_outputs(4673) <= not (a or b);
    layer8_outputs(4674) <= a;
    layer8_outputs(4675) <= not (a or b);
    layer8_outputs(4676) <= a and not b;
    layer8_outputs(4677) <= not (a or b);
    layer8_outputs(4678) <= a xor b;
    layer8_outputs(4679) <= a and not b;
    layer8_outputs(4680) <= a and b;
    layer8_outputs(4681) <= not b or a;
    layer8_outputs(4682) <= not b;
    layer8_outputs(4683) <= a;
    layer8_outputs(4684) <= a and b;
    layer8_outputs(4685) <= a or b;
    layer8_outputs(4686) <= not a;
    layer8_outputs(4687) <= not (a and b);
    layer8_outputs(4688) <= a and b;
    layer8_outputs(4689) <= a and b;
    layer8_outputs(4690) <= b;
    layer8_outputs(4691) <= not (a or b);
    layer8_outputs(4692) <= b and not a;
    layer8_outputs(4693) <= b;
    layer8_outputs(4694) <= not a;
    layer8_outputs(4695) <= b;
    layer8_outputs(4696) <= not b or a;
    layer8_outputs(4697) <= not b;
    layer8_outputs(4698) <= not a;
    layer8_outputs(4699) <= not b;
    layer8_outputs(4700) <= a and b;
    layer8_outputs(4701) <= not a;
    layer8_outputs(4702) <= a;
    layer8_outputs(4703) <= b;
    layer8_outputs(4704) <= not a;
    layer8_outputs(4705) <= a or b;
    layer8_outputs(4706) <= b;
    layer8_outputs(4707) <= '1';
    layer8_outputs(4708) <= b and not a;
    layer8_outputs(4709) <= a xor b;
    layer8_outputs(4710) <= b;
    layer8_outputs(4711) <= a xor b;
    layer8_outputs(4712) <= not (a or b);
    layer8_outputs(4713) <= not (a xor b);
    layer8_outputs(4714) <= not a;
    layer8_outputs(4715) <= a xor b;
    layer8_outputs(4716) <= a or b;
    layer8_outputs(4717) <= not a;
    layer8_outputs(4718) <= a;
    layer8_outputs(4719) <= not (a xor b);
    layer8_outputs(4720) <= not b or a;
    layer8_outputs(4721) <= not (a xor b);
    layer8_outputs(4722) <= b and not a;
    layer8_outputs(4723) <= not (a xor b);
    layer8_outputs(4724) <= b;
    layer8_outputs(4725) <= not a;
    layer8_outputs(4726) <= not a or b;
    layer8_outputs(4727) <= b;
    layer8_outputs(4728) <= not a;
    layer8_outputs(4729) <= a or b;
    layer8_outputs(4730) <= b;
    layer8_outputs(4731) <= a or b;
    layer8_outputs(4732) <= b and not a;
    layer8_outputs(4733) <= not (a or b);
    layer8_outputs(4734) <= b;
    layer8_outputs(4735) <= a and b;
    layer8_outputs(4736) <= not a or b;
    layer8_outputs(4737) <= not a;
    layer8_outputs(4738) <= a or b;
    layer8_outputs(4739) <= not (a xor b);
    layer8_outputs(4740) <= a or b;
    layer8_outputs(4741) <= not b;
    layer8_outputs(4742) <= a and b;
    layer8_outputs(4743) <= b;
    layer8_outputs(4744) <= not (a or b);
    layer8_outputs(4745) <= not b;
    layer8_outputs(4746) <= not a or b;
    layer8_outputs(4747) <= not b;
    layer8_outputs(4748) <= a or b;
    layer8_outputs(4749) <= not (a xor b);
    layer8_outputs(4750) <= not a;
    layer8_outputs(4751) <= not b;
    layer8_outputs(4752) <= not a or b;
    layer8_outputs(4753) <= not a;
    layer8_outputs(4754) <= not a;
    layer8_outputs(4755) <= not b;
    layer8_outputs(4756) <= not b;
    layer8_outputs(4757) <= not (a and b);
    layer8_outputs(4758) <= not (a xor b);
    layer8_outputs(4759) <= not b;
    layer8_outputs(4760) <= b and not a;
    layer8_outputs(4761) <= not b;
    layer8_outputs(4762) <= not (a and b);
    layer8_outputs(4763) <= not a;
    layer8_outputs(4764) <= not (a or b);
    layer8_outputs(4765) <= a xor b;
    layer8_outputs(4766) <= a and b;
    layer8_outputs(4767) <= b;
    layer8_outputs(4768) <= not a;
    layer8_outputs(4769) <= not b;
    layer8_outputs(4770) <= b;
    layer8_outputs(4771) <= not a;
    layer8_outputs(4772) <= not b or a;
    layer8_outputs(4773) <= a and b;
    layer8_outputs(4774) <= a xor b;
    layer8_outputs(4775) <= not a;
    layer8_outputs(4776) <= b and not a;
    layer8_outputs(4777) <= a and not b;
    layer8_outputs(4778) <= b and not a;
    layer8_outputs(4779) <= a and not b;
    layer8_outputs(4780) <= not (a xor b);
    layer8_outputs(4781) <= not (a xor b);
    layer8_outputs(4782) <= not (a xor b);
    layer8_outputs(4783) <= b and not a;
    layer8_outputs(4784) <= b and not a;
    layer8_outputs(4785) <= a;
    layer8_outputs(4786) <= not (a xor b);
    layer8_outputs(4787) <= not (a and b);
    layer8_outputs(4788) <= not a;
    layer8_outputs(4789) <= not a;
    layer8_outputs(4790) <= not (a xor b);
    layer8_outputs(4791) <= a xor b;
    layer8_outputs(4792) <= a xor b;
    layer8_outputs(4793) <= b;
    layer8_outputs(4794) <= a or b;
    layer8_outputs(4795) <= not a;
    layer8_outputs(4796) <= a and not b;
    layer8_outputs(4797) <= not b;
    layer8_outputs(4798) <= b;
    layer8_outputs(4799) <= a xor b;
    layer8_outputs(4800) <= not a;
    layer8_outputs(4801) <= not b;
    layer8_outputs(4802) <= a;
    layer8_outputs(4803) <= not a;
    layer8_outputs(4804) <= a or b;
    layer8_outputs(4805) <= not a or b;
    layer8_outputs(4806) <= not (a xor b);
    layer8_outputs(4807) <= a xor b;
    layer8_outputs(4808) <= not b or a;
    layer8_outputs(4809) <= a and b;
    layer8_outputs(4810) <= a;
    layer8_outputs(4811) <= not (a xor b);
    layer8_outputs(4812) <= not b;
    layer8_outputs(4813) <= not (a xor b);
    layer8_outputs(4814) <= not a or b;
    layer8_outputs(4815) <= b and not a;
    layer8_outputs(4816) <= a or b;
    layer8_outputs(4817) <= a;
    layer8_outputs(4818) <= a;
    layer8_outputs(4819) <= not a;
    layer8_outputs(4820) <= a and b;
    layer8_outputs(4821) <= not b;
    layer8_outputs(4822) <= a xor b;
    layer8_outputs(4823) <= not b;
    layer8_outputs(4824) <= not a;
    layer8_outputs(4825) <= b;
    layer8_outputs(4826) <= not a;
    layer8_outputs(4827) <= not b;
    layer8_outputs(4828) <= not (a and b);
    layer8_outputs(4829) <= b;
    layer8_outputs(4830) <= not a;
    layer8_outputs(4831) <= a xor b;
    layer8_outputs(4832) <= a and not b;
    layer8_outputs(4833) <= b;
    layer8_outputs(4834) <= b;
    layer8_outputs(4835) <= not (a xor b);
    layer8_outputs(4836) <= b;
    layer8_outputs(4837) <= a and not b;
    layer8_outputs(4838) <= not b;
    layer8_outputs(4839) <= not b;
    layer8_outputs(4840) <= not a or b;
    layer8_outputs(4841) <= a xor b;
    layer8_outputs(4842) <= not a or b;
    layer8_outputs(4843) <= not b or a;
    layer8_outputs(4844) <= not b;
    layer8_outputs(4845) <= a and not b;
    layer8_outputs(4846) <= not (a xor b);
    layer8_outputs(4847) <= not a or b;
    layer8_outputs(4848) <= not b or a;
    layer8_outputs(4849) <= b and not a;
    layer8_outputs(4850) <= not b;
    layer8_outputs(4851) <= a xor b;
    layer8_outputs(4852) <= not a;
    layer8_outputs(4853) <= a and not b;
    layer8_outputs(4854) <= b and not a;
    layer8_outputs(4855) <= not a;
    layer8_outputs(4856) <= not (a or b);
    layer8_outputs(4857) <= a or b;
    layer8_outputs(4858) <= a and not b;
    layer8_outputs(4859) <= b;
    layer8_outputs(4860) <= b;
    layer8_outputs(4861) <= not (a or b);
    layer8_outputs(4862) <= a;
    layer8_outputs(4863) <= not b;
    layer8_outputs(4864) <= b;
    layer8_outputs(4865) <= not (a or b);
    layer8_outputs(4866) <= not b;
    layer8_outputs(4867) <= a;
    layer8_outputs(4868) <= not a or b;
    layer8_outputs(4869) <= '1';
    layer8_outputs(4870) <= not (a xor b);
    layer8_outputs(4871) <= a;
    layer8_outputs(4872) <= not a or b;
    layer8_outputs(4873) <= b and not a;
    layer8_outputs(4874) <= not a or b;
    layer8_outputs(4875) <= not b;
    layer8_outputs(4876) <= a;
    layer8_outputs(4877) <= a xor b;
    layer8_outputs(4878) <= not a;
    layer8_outputs(4879) <= a or b;
    layer8_outputs(4880) <= a;
    layer8_outputs(4881) <= not (a or b);
    layer8_outputs(4882) <= not (a xor b);
    layer8_outputs(4883) <= a or b;
    layer8_outputs(4884) <= b and not a;
    layer8_outputs(4885) <= a and not b;
    layer8_outputs(4886) <= b;
    layer8_outputs(4887) <= '0';
    layer8_outputs(4888) <= not b or a;
    layer8_outputs(4889) <= b;
    layer8_outputs(4890) <= not b;
    layer8_outputs(4891) <= not b;
    layer8_outputs(4892) <= not b or a;
    layer8_outputs(4893) <= not (a or b);
    layer8_outputs(4894) <= b and not a;
    layer8_outputs(4895) <= not a;
    layer8_outputs(4896) <= not a;
    layer8_outputs(4897) <= not (a and b);
    layer8_outputs(4898) <= a;
    layer8_outputs(4899) <= not (a or b);
    layer8_outputs(4900) <= not b;
    layer8_outputs(4901) <= b;
    layer8_outputs(4902) <= a xor b;
    layer8_outputs(4903) <= not b;
    layer8_outputs(4904) <= b and not a;
    layer8_outputs(4905) <= a or b;
    layer8_outputs(4906) <= a and b;
    layer8_outputs(4907) <= b;
    layer8_outputs(4908) <= a;
    layer8_outputs(4909) <= b;
    layer8_outputs(4910) <= not (a xor b);
    layer8_outputs(4911) <= not b;
    layer8_outputs(4912) <= not b;
    layer8_outputs(4913) <= not a or b;
    layer8_outputs(4914) <= a xor b;
    layer8_outputs(4915) <= b;
    layer8_outputs(4916) <= not b or a;
    layer8_outputs(4917) <= a and not b;
    layer8_outputs(4918) <= not (a or b);
    layer8_outputs(4919) <= not b or a;
    layer8_outputs(4920) <= a;
    layer8_outputs(4921) <= b and not a;
    layer8_outputs(4922) <= b;
    layer8_outputs(4923) <= a xor b;
    layer8_outputs(4924) <= b;
    layer8_outputs(4925) <= a and not b;
    layer8_outputs(4926) <= a;
    layer8_outputs(4927) <= a;
    layer8_outputs(4928) <= not (a and b);
    layer8_outputs(4929) <= a;
    layer8_outputs(4930) <= b;
    layer8_outputs(4931) <= not a;
    layer8_outputs(4932) <= not (a xor b);
    layer8_outputs(4933) <= a xor b;
    layer8_outputs(4934) <= not a or b;
    layer8_outputs(4935) <= not a;
    layer8_outputs(4936) <= not (a or b);
    layer8_outputs(4937) <= not b;
    layer8_outputs(4938) <= not a;
    layer8_outputs(4939) <= not b;
    layer8_outputs(4940) <= not b;
    layer8_outputs(4941) <= not a or b;
    layer8_outputs(4942) <= a xor b;
    layer8_outputs(4943) <= a;
    layer8_outputs(4944) <= not b;
    layer8_outputs(4945) <= not a;
    layer8_outputs(4946) <= a xor b;
    layer8_outputs(4947) <= a;
    layer8_outputs(4948) <= a xor b;
    layer8_outputs(4949) <= b;
    layer8_outputs(4950) <= a;
    layer8_outputs(4951) <= a or b;
    layer8_outputs(4952) <= not b;
    layer8_outputs(4953) <= not (a or b);
    layer8_outputs(4954) <= a xor b;
    layer8_outputs(4955) <= a;
    layer8_outputs(4956) <= not b or a;
    layer8_outputs(4957) <= b;
    layer8_outputs(4958) <= a or b;
    layer8_outputs(4959) <= a xor b;
    layer8_outputs(4960) <= not a or b;
    layer8_outputs(4961) <= b;
    layer8_outputs(4962) <= not a;
    layer8_outputs(4963) <= not b or a;
    layer8_outputs(4964) <= not a or b;
    layer8_outputs(4965) <= not (a xor b);
    layer8_outputs(4966) <= not (a xor b);
    layer8_outputs(4967) <= b;
    layer8_outputs(4968) <= a;
    layer8_outputs(4969) <= not a;
    layer8_outputs(4970) <= not (a xor b);
    layer8_outputs(4971) <= a or b;
    layer8_outputs(4972) <= not a;
    layer8_outputs(4973) <= not b;
    layer8_outputs(4974) <= a xor b;
    layer8_outputs(4975) <= b;
    layer8_outputs(4976) <= not b;
    layer8_outputs(4977) <= b;
    layer8_outputs(4978) <= not a;
    layer8_outputs(4979) <= not b;
    layer8_outputs(4980) <= not b;
    layer8_outputs(4981) <= a and not b;
    layer8_outputs(4982) <= not b or a;
    layer8_outputs(4983) <= not (a or b);
    layer8_outputs(4984) <= not b;
    layer8_outputs(4985) <= b and not a;
    layer8_outputs(4986) <= b;
    layer8_outputs(4987) <= a and not b;
    layer8_outputs(4988) <= not a or b;
    layer8_outputs(4989) <= a or b;
    layer8_outputs(4990) <= not a or b;
    layer8_outputs(4991) <= b and not a;
    layer8_outputs(4992) <= a and b;
    layer8_outputs(4993) <= not a or b;
    layer8_outputs(4994) <= a;
    layer8_outputs(4995) <= a or b;
    layer8_outputs(4996) <= not a or b;
    layer8_outputs(4997) <= not a or b;
    layer8_outputs(4998) <= not a;
    layer8_outputs(4999) <= a;
    layer8_outputs(5000) <= not b;
    layer8_outputs(5001) <= not a;
    layer8_outputs(5002) <= not a;
    layer8_outputs(5003) <= a;
    layer8_outputs(5004) <= a;
    layer8_outputs(5005) <= not a or b;
    layer8_outputs(5006) <= b;
    layer8_outputs(5007) <= not a;
    layer8_outputs(5008) <= not a or b;
    layer8_outputs(5009) <= a and not b;
    layer8_outputs(5010) <= a and b;
    layer8_outputs(5011) <= not a;
    layer8_outputs(5012) <= not (a or b);
    layer8_outputs(5013) <= a or b;
    layer8_outputs(5014) <= not (a xor b);
    layer8_outputs(5015) <= a xor b;
    layer8_outputs(5016) <= a;
    layer8_outputs(5017) <= a;
    layer8_outputs(5018) <= a and not b;
    layer8_outputs(5019) <= a xor b;
    layer8_outputs(5020) <= not (a or b);
    layer8_outputs(5021) <= a xor b;
    layer8_outputs(5022) <= a xor b;
    layer8_outputs(5023) <= a xor b;
    layer8_outputs(5024) <= a xor b;
    layer8_outputs(5025) <= a and not b;
    layer8_outputs(5026) <= a and b;
    layer8_outputs(5027) <= '0';
    layer8_outputs(5028) <= not b;
    layer8_outputs(5029) <= not (a xor b);
    layer8_outputs(5030) <= not (a xor b);
    layer8_outputs(5031) <= not a;
    layer8_outputs(5032) <= a;
    layer8_outputs(5033) <= b and not a;
    layer8_outputs(5034) <= not a;
    layer8_outputs(5035) <= not (a or b);
    layer8_outputs(5036) <= a;
    layer8_outputs(5037) <= not (a and b);
    layer8_outputs(5038) <= b;
    layer8_outputs(5039) <= not b or a;
    layer8_outputs(5040) <= not (a xor b);
    layer8_outputs(5041) <= a or b;
    layer8_outputs(5042) <= b and not a;
    layer8_outputs(5043) <= a and b;
    layer8_outputs(5044) <= a and b;
    layer8_outputs(5045) <= not a;
    layer8_outputs(5046) <= a xor b;
    layer8_outputs(5047) <= not (a or b);
    layer8_outputs(5048) <= not a;
    layer8_outputs(5049) <= a or b;
    layer8_outputs(5050) <= b;
    layer8_outputs(5051) <= b;
    layer8_outputs(5052) <= not b;
    layer8_outputs(5053) <= not (a xor b);
    layer8_outputs(5054) <= a;
    layer8_outputs(5055) <= b;
    layer8_outputs(5056) <= b;
    layer8_outputs(5057) <= not (a and b);
    layer8_outputs(5058) <= not (a xor b);
    layer8_outputs(5059) <= a and b;
    layer8_outputs(5060) <= not (a xor b);
    layer8_outputs(5061) <= a and not b;
    layer8_outputs(5062) <= not (a or b);
    layer8_outputs(5063) <= a xor b;
    layer8_outputs(5064) <= a xor b;
    layer8_outputs(5065) <= not a or b;
    layer8_outputs(5066) <= b;
    layer8_outputs(5067) <= not a;
    layer8_outputs(5068) <= not (a xor b);
    layer8_outputs(5069) <= a;
    layer8_outputs(5070) <= b;
    layer8_outputs(5071) <= not a;
    layer8_outputs(5072) <= not (a xor b);
    layer8_outputs(5073) <= a xor b;
    layer8_outputs(5074) <= not (a xor b);
    layer8_outputs(5075) <= a xor b;
    layer8_outputs(5076) <= not b;
    layer8_outputs(5077) <= a and b;
    layer8_outputs(5078) <= not b;
    layer8_outputs(5079) <= not b or a;
    layer8_outputs(5080) <= not (a and b);
    layer8_outputs(5081) <= a xor b;
    layer8_outputs(5082) <= a xor b;
    layer8_outputs(5083) <= not a;
    layer8_outputs(5084) <= a or b;
    layer8_outputs(5085) <= b;
    layer8_outputs(5086) <= not (a or b);
    layer8_outputs(5087) <= not (a xor b);
    layer8_outputs(5088) <= a xor b;
    layer8_outputs(5089) <= not b or a;
    layer8_outputs(5090) <= a and not b;
    layer8_outputs(5091) <= a xor b;
    layer8_outputs(5092) <= not a;
    layer8_outputs(5093) <= a;
    layer8_outputs(5094) <= a;
    layer8_outputs(5095) <= a and b;
    layer8_outputs(5096) <= a or b;
    layer8_outputs(5097) <= not (a xor b);
    layer8_outputs(5098) <= b;
    layer8_outputs(5099) <= b and not a;
    layer8_outputs(5100) <= a or b;
    layer8_outputs(5101) <= b and not a;
    layer8_outputs(5102) <= not b;
    layer8_outputs(5103) <= b;
    layer8_outputs(5104) <= b and not a;
    layer8_outputs(5105) <= not (a xor b);
    layer8_outputs(5106) <= a xor b;
    layer8_outputs(5107) <= not (a xor b);
    layer8_outputs(5108) <= a or b;
    layer8_outputs(5109) <= a or b;
    layer8_outputs(5110) <= a xor b;
    layer8_outputs(5111) <= a and not b;
    layer8_outputs(5112) <= b;
    layer8_outputs(5113) <= b;
    layer8_outputs(5114) <= b and not a;
    layer8_outputs(5115) <= b and not a;
    layer8_outputs(5116) <= not a;
    layer8_outputs(5117) <= a;
    layer8_outputs(5118) <= b;
    layer8_outputs(5119) <= not (a or b);
    layer8_outputs(5120) <= not a;
    layer8_outputs(5121) <= not (a or b);
    layer8_outputs(5122) <= not a;
    layer8_outputs(5123) <= not (a or b);
    layer8_outputs(5124) <= a;
    layer8_outputs(5125) <= not (a or b);
    layer8_outputs(5126) <= not (a xor b);
    layer8_outputs(5127) <= a xor b;
    layer8_outputs(5128) <= not a;
    layer8_outputs(5129) <= not (a xor b);
    layer8_outputs(5130) <= a and not b;
    layer8_outputs(5131) <= a xor b;
    layer8_outputs(5132) <= b;
    layer8_outputs(5133) <= a;
    layer8_outputs(5134) <= '1';
    layer8_outputs(5135) <= not b;
    layer8_outputs(5136) <= a xor b;
    layer8_outputs(5137) <= a xor b;
    layer8_outputs(5138) <= a;
    layer8_outputs(5139) <= not (a xor b);
    layer8_outputs(5140) <= not b;
    layer8_outputs(5141) <= not a;
    layer8_outputs(5142) <= a;
    layer8_outputs(5143) <= a xor b;
    layer8_outputs(5144) <= a;
    layer8_outputs(5145) <= a xor b;
    layer8_outputs(5146) <= a;
    layer8_outputs(5147) <= not (a or b);
    layer8_outputs(5148) <= a;
    layer8_outputs(5149) <= b;
    layer8_outputs(5150) <= a or b;
    layer8_outputs(5151) <= not (a xor b);
    layer8_outputs(5152) <= b;
    layer8_outputs(5153) <= b;
    layer8_outputs(5154) <= not b or a;
    layer8_outputs(5155) <= b and not a;
    layer8_outputs(5156) <= a xor b;
    layer8_outputs(5157) <= not (a xor b);
    layer8_outputs(5158) <= a;
    layer8_outputs(5159) <= b;
    layer8_outputs(5160) <= not (a or b);
    layer8_outputs(5161) <= not (a xor b);
    layer8_outputs(5162) <= a;
    layer8_outputs(5163) <= not a;
    layer8_outputs(5164) <= a xor b;
    layer8_outputs(5165) <= '1';
    layer8_outputs(5166) <= not a;
    layer8_outputs(5167) <= a xor b;
    layer8_outputs(5168) <= b and not a;
    layer8_outputs(5169) <= not a;
    layer8_outputs(5170) <= not a or b;
    layer8_outputs(5171) <= not (a and b);
    layer8_outputs(5172) <= not a;
    layer8_outputs(5173) <= not a or b;
    layer8_outputs(5174) <= not (a or b);
    layer8_outputs(5175) <= a;
    layer8_outputs(5176) <= b;
    layer8_outputs(5177) <= b;
    layer8_outputs(5178) <= a xor b;
    layer8_outputs(5179) <= b and not a;
    layer8_outputs(5180) <= not (a and b);
    layer8_outputs(5181) <= not (a or b);
    layer8_outputs(5182) <= not b;
    layer8_outputs(5183) <= a and not b;
    layer8_outputs(5184) <= not a or b;
    layer8_outputs(5185) <= '0';
    layer8_outputs(5186) <= not (a xor b);
    layer8_outputs(5187) <= a xor b;
    layer8_outputs(5188) <= a xor b;
    layer8_outputs(5189) <= b;
    layer8_outputs(5190) <= a;
    layer8_outputs(5191) <= a;
    layer8_outputs(5192) <= not (a xor b);
    layer8_outputs(5193) <= not (a and b);
    layer8_outputs(5194) <= not (a or b);
    layer8_outputs(5195) <= not a;
    layer8_outputs(5196) <= a and b;
    layer8_outputs(5197) <= a xor b;
    layer8_outputs(5198) <= b and not a;
    layer8_outputs(5199) <= not a;
    layer8_outputs(5200) <= not (a xor b);
    layer8_outputs(5201) <= a;
    layer8_outputs(5202) <= b and not a;
    layer8_outputs(5203) <= not a;
    layer8_outputs(5204) <= b;
    layer8_outputs(5205) <= a xor b;
    layer8_outputs(5206) <= a and not b;
    layer8_outputs(5207) <= not a;
    layer8_outputs(5208) <= a xor b;
    layer8_outputs(5209) <= a and b;
    layer8_outputs(5210) <= a;
    layer8_outputs(5211) <= a;
    layer8_outputs(5212) <= a or b;
    layer8_outputs(5213) <= b;
    layer8_outputs(5214) <= not (a xor b);
    layer8_outputs(5215) <= b;
    layer8_outputs(5216) <= a;
    layer8_outputs(5217) <= not b;
    layer8_outputs(5218) <= b and not a;
    layer8_outputs(5219) <= not a;
    layer8_outputs(5220) <= not b or a;
    layer8_outputs(5221) <= b;
    layer8_outputs(5222) <= b;
    layer8_outputs(5223) <= not (a xor b);
    layer8_outputs(5224) <= not (a or b);
    layer8_outputs(5225) <= not a;
    layer8_outputs(5226) <= not a;
    layer8_outputs(5227) <= a and b;
    layer8_outputs(5228) <= not (a or b);
    layer8_outputs(5229) <= b;
    layer8_outputs(5230) <= b;
    layer8_outputs(5231) <= b and not a;
    layer8_outputs(5232) <= not (a xor b);
    layer8_outputs(5233) <= not b;
    layer8_outputs(5234) <= a or b;
    layer8_outputs(5235) <= not a;
    layer8_outputs(5236) <= a and not b;
    layer8_outputs(5237) <= not b or a;
    layer8_outputs(5238) <= a or b;
    layer8_outputs(5239) <= a and b;
    layer8_outputs(5240) <= a or b;
    layer8_outputs(5241) <= a;
    layer8_outputs(5242) <= not a;
    layer8_outputs(5243) <= not b;
    layer8_outputs(5244) <= a and not b;
    layer8_outputs(5245) <= a and b;
    layer8_outputs(5246) <= not a;
    layer8_outputs(5247) <= a;
    layer8_outputs(5248) <= not a;
    layer8_outputs(5249) <= not b;
    layer8_outputs(5250) <= not b;
    layer8_outputs(5251) <= a or b;
    layer8_outputs(5252) <= not (a xor b);
    layer8_outputs(5253) <= not a;
    layer8_outputs(5254) <= b;
    layer8_outputs(5255) <= a or b;
    layer8_outputs(5256) <= not a or b;
    layer8_outputs(5257) <= b;
    layer8_outputs(5258) <= not a;
    layer8_outputs(5259) <= b and not a;
    layer8_outputs(5260) <= not a;
    layer8_outputs(5261) <= a xor b;
    layer8_outputs(5262) <= not a;
    layer8_outputs(5263) <= not b or a;
    layer8_outputs(5264) <= b;
    layer8_outputs(5265) <= not b;
    layer8_outputs(5266) <= a;
    layer8_outputs(5267) <= not a;
    layer8_outputs(5268) <= b;
    layer8_outputs(5269) <= not a or b;
    layer8_outputs(5270) <= a xor b;
    layer8_outputs(5271) <= not (a xor b);
    layer8_outputs(5272) <= a;
    layer8_outputs(5273) <= b;
    layer8_outputs(5274) <= not (a or b);
    layer8_outputs(5275) <= a or b;
    layer8_outputs(5276) <= a xor b;
    layer8_outputs(5277) <= b;
    layer8_outputs(5278) <= not b;
    layer8_outputs(5279) <= not (a xor b);
    layer8_outputs(5280) <= '1';
    layer8_outputs(5281) <= a xor b;
    layer8_outputs(5282) <= a;
    layer8_outputs(5283) <= not (a or b);
    layer8_outputs(5284) <= a xor b;
    layer8_outputs(5285) <= not (a or b);
    layer8_outputs(5286) <= not b or a;
    layer8_outputs(5287) <= not b or a;
    layer8_outputs(5288) <= not a or b;
    layer8_outputs(5289) <= b;
    layer8_outputs(5290) <= not b;
    layer8_outputs(5291) <= a;
    layer8_outputs(5292) <= not a or b;
    layer8_outputs(5293) <= a and not b;
    layer8_outputs(5294) <= a or b;
    layer8_outputs(5295) <= not a;
    layer8_outputs(5296) <= a;
    layer8_outputs(5297) <= not (a xor b);
    layer8_outputs(5298) <= a xor b;
    layer8_outputs(5299) <= not (a xor b);
    layer8_outputs(5300) <= not (a or b);
    layer8_outputs(5301) <= b and not a;
    layer8_outputs(5302) <= a xor b;
    layer8_outputs(5303) <= a and b;
    layer8_outputs(5304) <= not (a xor b);
    layer8_outputs(5305) <= not (a and b);
    layer8_outputs(5306) <= not a;
    layer8_outputs(5307) <= not (a xor b);
    layer8_outputs(5308) <= a and not b;
    layer8_outputs(5309) <= b;
    layer8_outputs(5310) <= a or b;
    layer8_outputs(5311) <= not a;
    layer8_outputs(5312) <= a and b;
    layer8_outputs(5313) <= '0';
    layer8_outputs(5314) <= not a;
    layer8_outputs(5315) <= not a;
    layer8_outputs(5316) <= not b;
    layer8_outputs(5317) <= not (a and b);
    layer8_outputs(5318) <= b;
    layer8_outputs(5319) <= a or b;
    layer8_outputs(5320) <= not (a and b);
    layer8_outputs(5321) <= b and not a;
    layer8_outputs(5322) <= a;
    layer8_outputs(5323) <= b;
    layer8_outputs(5324) <= not a;
    layer8_outputs(5325) <= not a;
    layer8_outputs(5326) <= not a;
    layer8_outputs(5327) <= not b;
    layer8_outputs(5328) <= a;
    layer8_outputs(5329) <= b and not a;
    layer8_outputs(5330) <= not b;
    layer8_outputs(5331) <= b and not a;
    layer8_outputs(5332) <= b;
    layer8_outputs(5333) <= a xor b;
    layer8_outputs(5334) <= not a;
    layer8_outputs(5335) <= not b;
    layer8_outputs(5336) <= a xor b;
    layer8_outputs(5337) <= a and not b;
    layer8_outputs(5338) <= a and not b;
    layer8_outputs(5339) <= b;
    layer8_outputs(5340) <= not a or b;
    layer8_outputs(5341) <= a xor b;
    layer8_outputs(5342) <= not (a or b);
    layer8_outputs(5343) <= not b;
    layer8_outputs(5344) <= a and b;
    layer8_outputs(5345) <= not a;
    layer8_outputs(5346) <= b and not a;
    layer8_outputs(5347) <= not b;
    layer8_outputs(5348) <= a and b;
    layer8_outputs(5349) <= not (a and b);
    layer8_outputs(5350) <= not b;
    layer8_outputs(5351) <= a xor b;
    layer8_outputs(5352) <= b;
    layer8_outputs(5353) <= a and b;
    layer8_outputs(5354) <= a and not b;
    layer8_outputs(5355) <= a xor b;
    layer8_outputs(5356) <= b;
    layer8_outputs(5357) <= b;
    layer8_outputs(5358) <= not b;
    layer8_outputs(5359) <= a and b;
    layer8_outputs(5360) <= not a;
    layer8_outputs(5361) <= not a;
    layer8_outputs(5362) <= not (a and b);
    layer8_outputs(5363) <= not a;
    layer8_outputs(5364) <= not (a xor b);
    layer8_outputs(5365) <= not (a xor b);
    layer8_outputs(5366) <= a xor b;
    layer8_outputs(5367) <= a;
    layer8_outputs(5368) <= not a;
    layer8_outputs(5369) <= not a or b;
    layer8_outputs(5370) <= a;
    layer8_outputs(5371) <= not (a and b);
    layer8_outputs(5372) <= not b or a;
    layer8_outputs(5373) <= not (a xor b);
    layer8_outputs(5374) <= b;
    layer8_outputs(5375) <= not (a or b);
    layer8_outputs(5376) <= not (a xor b);
    layer8_outputs(5377) <= not a;
    layer8_outputs(5378) <= a and b;
    layer8_outputs(5379) <= not a;
    layer8_outputs(5380) <= a;
    layer8_outputs(5381) <= a xor b;
    layer8_outputs(5382) <= b;
    layer8_outputs(5383) <= not (a and b);
    layer8_outputs(5384) <= not (a or b);
    layer8_outputs(5385) <= not b;
    layer8_outputs(5386) <= not a;
    layer8_outputs(5387) <= not a;
    layer8_outputs(5388) <= a;
    layer8_outputs(5389) <= not b;
    layer8_outputs(5390) <= a and b;
    layer8_outputs(5391) <= a or b;
    layer8_outputs(5392) <= not a;
    layer8_outputs(5393) <= b;
    layer8_outputs(5394) <= not (a or b);
    layer8_outputs(5395) <= not b;
    layer8_outputs(5396) <= not b or a;
    layer8_outputs(5397) <= not (a xor b);
    layer8_outputs(5398) <= b;
    layer8_outputs(5399) <= not b;
    layer8_outputs(5400) <= b;
    layer8_outputs(5401) <= not b;
    layer8_outputs(5402) <= a xor b;
    layer8_outputs(5403) <= not a;
    layer8_outputs(5404) <= a;
    layer8_outputs(5405) <= not a;
    layer8_outputs(5406) <= not a or b;
    layer8_outputs(5407) <= a xor b;
    layer8_outputs(5408) <= a;
    layer8_outputs(5409) <= not a;
    layer8_outputs(5410) <= a xor b;
    layer8_outputs(5411) <= not (a and b);
    layer8_outputs(5412) <= a;
    layer8_outputs(5413) <= not b;
    layer8_outputs(5414) <= a xor b;
    layer8_outputs(5415) <= not b or a;
    layer8_outputs(5416) <= not b;
    layer8_outputs(5417) <= not (a xor b);
    layer8_outputs(5418) <= a and b;
    layer8_outputs(5419) <= a xor b;
    layer8_outputs(5420) <= not (a and b);
    layer8_outputs(5421) <= not a or b;
    layer8_outputs(5422) <= not (a or b);
    layer8_outputs(5423) <= not b;
    layer8_outputs(5424) <= a or b;
    layer8_outputs(5425) <= a xor b;
    layer8_outputs(5426) <= not a;
    layer8_outputs(5427) <= a and b;
    layer8_outputs(5428) <= a and b;
    layer8_outputs(5429) <= a and b;
    layer8_outputs(5430) <= a and b;
    layer8_outputs(5431) <= not (a and b);
    layer8_outputs(5432) <= b;
    layer8_outputs(5433) <= not (a or b);
    layer8_outputs(5434) <= not (a or b);
    layer8_outputs(5435) <= a xor b;
    layer8_outputs(5436) <= b;
    layer8_outputs(5437) <= a and b;
    layer8_outputs(5438) <= not a or b;
    layer8_outputs(5439) <= b and not a;
    layer8_outputs(5440) <= a;
    layer8_outputs(5441) <= not a or b;
    layer8_outputs(5442) <= b;
    layer8_outputs(5443) <= not a or b;
    layer8_outputs(5444) <= not (a xor b);
    layer8_outputs(5445) <= not b;
    layer8_outputs(5446) <= a and not b;
    layer8_outputs(5447) <= not b;
    layer8_outputs(5448) <= a or b;
    layer8_outputs(5449) <= not a;
    layer8_outputs(5450) <= not (a xor b);
    layer8_outputs(5451) <= a;
    layer8_outputs(5452) <= not b;
    layer8_outputs(5453) <= not (a xor b);
    layer8_outputs(5454) <= not (a xor b);
    layer8_outputs(5455) <= not a;
    layer8_outputs(5456) <= a;
    layer8_outputs(5457) <= b;
    layer8_outputs(5458) <= not b;
    layer8_outputs(5459) <= a;
    layer8_outputs(5460) <= not a;
    layer8_outputs(5461) <= a xor b;
    layer8_outputs(5462) <= not a or b;
    layer8_outputs(5463) <= not (a xor b);
    layer8_outputs(5464) <= b;
    layer8_outputs(5465) <= b;
    layer8_outputs(5466) <= '0';
    layer8_outputs(5467) <= not a;
    layer8_outputs(5468) <= b;
    layer8_outputs(5469) <= a or b;
    layer8_outputs(5470) <= b and not a;
    layer8_outputs(5471) <= not b or a;
    layer8_outputs(5472) <= b and not a;
    layer8_outputs(5473) <= not b;
    layer8_outputs(5474) <= not a;
    layer8_outputs(5475) <= not (a xor b);
    layer8_outputs(5476) <= not a;
    layer8_outputs(5477) <= not b;
    layer8_outputs(5478) <= a;
    layer8_outputs(5479) <= not a;
    layer8_outputs(5480) <= not a;
    layer8_outputs(5481) <= '0';
    layer8_outputs(5482) <= not b;
    layer8_outputs(5483) <= a;
    layer8_outputs(5484) <= not (a xor b);
    layer8_outputs(5485) <= not b;
    layer8_outputs(5486) <= not a;
    layer8_outputs(5487) <= a xor b;
    layer8_outputs(5488) <= not a or b;
    layer8_outputs(5489) <= a;
    layer8_outputs(5490) <= a and b;
    layer8_outputs(5491) <= not (a xor b);
    layer8_outputs(5492) <= not b;
    layer8_outputs(5493) <= not (a or b);
    layer8_outputs(5494) <= not (a xor b);
    layer8_outputs(5495) <= b;
    layer8_outputs(5496) <= a xor b;
    layer8_outputs(5497) <= not a;
    layer8_outputs(5498) <= a or b;
    layer8_outputs(5499) <= b;
    layer8_outputs(5500) <= not a;
    layer8_outputs(5501) <= a;
    layer8_outputs(5502) <= a;
    layer8_outputs(5503) <= not (a xor b);
    layer8_outputs(5504) <= not b;
    layer8_outputs(5505) <= not a;
    layer8_outputs(5506) <= a or b;
    layer8_outputs(5507) <= not (a xor b);
    layer8_outputs(5508) <= b;
    layer8_outputs(5509) <= not b;
    layer8_outputs(5510) <= '0';
    layer8_outputs(5511) <= a;
    layer8_outputs(5512) <= not a;
    layer8_outputs(5513) <= a;
    layer8_outputs(5514) <= not a;
    layer8_outputs(5515) <= not a or b;
    layer8_outputs(5516) <= not (a xor b);
    layer8_outputs(5517) <= not b or a;
    layer8_outputs(5518) <= a or b;
    layer8_outputs(5519) <= not a;
    layer8_outputs(5520) <= not b or a;
    layer8_outputs(5521) <= not (a xor b);
    layer8_outputs(5522) <= not (a xor b);
    layer8_outputs(5523) <= a or b;
    layer8_outputs(5524) <= not b;
    layer8_outputs(5525) <= not (a and b);
    layer8_outputs(5526) <= not (a xor b);
    layer8_outputs(5527) <= b;
    layer8_outputs(5528) <= a;
    layer8_outputs(5529) <= b;
    layer8_outputs(5530) <= not a;
    layer8_outputs(5531) <= not a;
    layer8_outputs(5532) <= a;
    layer8_outputs(5533) <= a and b;
    layer8_outputs(5534) <= not (a xor b);
    layer8_outputs(5535) <= a xor b;
    layer8_outputs(5536) <= a xor b;
    layer8_outputs(5537) <= a;
    layer8_outputs(5538) <= not (a xor b);
    layer8_outputs(5539) <= not a or b;
    layer8_outputs(5540) <= a xor b;
    layer8_outputs(5541) <= not b;
    layer8_outputs(5542) <= not (a or b);
    layer8_outputs(5543) <= not a;
    layer8_outputs(5544) <= not b;
    layer8_outputs(5545) <= b;
    layer8_outputs(5546) <= b;
    layer8_outputs(5547) <= a xor b;
    layer8_outputs(5548) <= a and b;
    layer8_outputs(5549) <= a;
    layer8_outputs(5550) <= not a;
    layer8_outputs(5551) <= not b;
    layer8_outputs(5552) <= a and not b;
    layer8_outputs(5553) <= b;
    layer8_outputs(5554) <= not (a or b);
    layer8_outputs(5555) <= not b;
    layer8_outputs(5556) <= a;
    layer8_outputs(5557) <= not (a and b);
    layer8_outputs(5558) <= not a or b;
    layer8_outputs(5559) <= b;
    layer8_outputs(5560) <= not (a xor b);
    layer8_outputs(5561) <= b;
    layer8_outputs(5562) <= not a;
    layer8_outputs(5563) <= not (a and b);
    layer8_outputs(5564) <= not (a and b);
    layer8_outputs(5565) <= b and not a;
    layer8_outputs(5566) <= not b or a;
    layer8_outputs(5567) <= not b;
    layer8_outputs(5568) <= a and not b;
    layer8_outputs(5569) <= not a;
    layer8_outputs(5570) <= not (a and b);
    layer8_outputs(5571) <= not (a xor b);
    layer8_outputs(5572) <= not (a and b);
    layer8_outputs(5573) <= not b or a;
    layer8_outputs(5574) <= a;
    layer8_outputs(5575) <= not a;
    layer8_outputs(5576) <= not (a xor b);
    layer8_outputs(5577) <= not a;
    layer8_outputs(5578) <= not a;
    layer8_outputs(5579) <= not (a and b);
    layer8_outputs(5580) <= a and b;
    layer8_outputs(5581) <= not (a xor b);
    layer8_outputs(5582) <= not b;
    layer8_outputs(5583) <= a;
    layer8_outputs(5584) <= a and b;
    layer8_outputs(5585) <= a xor b;
    layer8_outputs(5586) <= not (a xor b);
    layer8_outputs(5587) <= a;
    layer8_outputs(5588) <= not b;
    layer8_outputs(5589) <= a xor b;
    layer8_outputs(5590) <= a xor b;
    layer8_outputs(5591) <= not b;
    layer8_outputs(5592) <= not b;
    layer8_outputs(5593) <= a or b;
    layer8_outputs(5594) <= a;
    layer8_outputs(5595) <= a xor b;
    layer8_outputs(5596) <= b and not a;
    layer8_outputs(5597) <= b and not a;
    layer8_outputs(5598) <= a and not b;
    layer8_outputs(5599) <= not b or a;
    layer8_outputs(5600) <= not (a xor b);
    layer8_outputs(5601) <= a xor b;
    layer8_outputs(5602) <= a;
    layer8_outputs(5603) <= not (a xor b);
    layer8_outputs(5604) <= b and not a;
    layer8_outputs(5605) <= a xor b;
    layer8_outputs(5606) <= a;
    layer8_outputs(5607) <= not b or a;
    layer8_outputs(5608) <= b and not a;
    layer8_outputs(5609) <= a and b;
    layer8_outputs(5610) <= a;
    layer8_outputs(5611) <= a xor b;
    layer8_outputs(5612) <= b;
    layer8_outputs(5613) <= a or b;
    layer8_outputs(5614) <= not (a and b);
    layer8_outputs(5615) <= a and not b;
    layer8_outputs(5616) <= not a;
    layer8_outputs(5617) <= b;
    layer8_outputs(5618) <= a xor b;
    layer8_outputs(5619) <= not b;
    layer8_outputs(5620) <= not (a xor b);
    layer8_outputs(5621) <= not b or a;
    layer8_outputs(5622) <= b;
    layer8_outputs(5623) <= not (a xor b);
    layer8_outputs(5624) <= a and b;
    layer8_outputs(5625) <= not (a or b);
    layer8_outputs(5626) <= not (a or b);
    layer8_outputs(5627) <= not b;
    layer8_outputs(5628) <= b;
    layer8_outputs(5629) <= a and not b;
    layer8_outputs(5630) <= b and not a;
    layer8_outputs(5631) <= b;
    layer8_outputs(5632) <= not a;
    layer8_outputs(5633) <= not a;
    layer8_outputs(5634) <= b and not a;
    layer8_outputs(5635) <= a;
    layer8_outputs(5636) <= not b;
    layer8_outputs(5637) <= not (a xor b);
    layer8_outputs(5638) <= not a;
    layer8_outputs(5639) <= not a;
    layer8_outputs(5640) <= not b;
    layer8_outputs(5641) <= a or b;
    layer8_outputs(5642) <= a;
    layer8_outputs(5643) <= a or b;
    layer8_outputs(5644) <= not b or a;
    layer8_outputs(5645) <= not a or b;
    layer8_outputs(5646) <= not (a xor b);
    layer8_outputs(5647) <= a and b;
    layer8_outputs(5648) <= not a;
    layer8_outputs(5649) <= not a;
    layer8_outputs(5650) <= not b;
    layer8_outputs(5651) <= b and not a;
    layer8_outputs(5652) <= not (a and b);
    layer8_outputs(5653) <= b;
    layer8_outputs(5654) <= not b or a;
    layer8_outputs(5655) <= not a;
    layer8_outputs(5656) <= b;
    layer8_outputs(5657) <= not b or a;
    layer8_outputs(5658) <= a xor b;
    layer8_outputs(5659) <= a;
    layer8_outputs(5660) <= not a;
    layer8_outputs(5661) <= b;
    layer8_outputs(5662) <= a;
    layer8_outputs(5663) <= b;
    layer8_outputs(5664) <= a xor b;
    layer8_outputs(5665) <= a xor b;
    layer8_outputs(5666) <= not a or b;
    layer8_outputs(5667) <= b;
    layer8_outputs(5668) <= not b or a;
    layer8_outputs(5669) <= a xor b;
    layer8_outputs(5670) <= not a;
    layer8_outputs(5671) <= not a or b;
    layer8_outputs(5672) <= b and not a;
    layer8_outputs(5673) <= not (a xor b);
    layer8_outputs(5674) <= not b;
    layer8_outputs(5675) <= b;
    layer8_outputs(5676) <= not (a xor b);
    layer8_outputs(5677) <= b;
    layer8_outputs(5678) <= not (a or b);
    layer8_outputs(5679) <= a and not b;
    layer8_outputs(5680) <= a or b;
    layer8_outputs(5681) <= not (a or b);
    layer8_outputs(5682) <= not a;
    layer8_outputs(5683) <= a;
    layer8_outputs(5684) <= not a;
    layer8_outputs(5685) <= not a;
    layer8_outputs(5686) <= a xor b;
    layer8_outputs(5687) <= not b;
    layer8_outputs(5688) <= not (a xor b);
    layer8_outputs(5689) <= b;
    layer8_outputs(5690) <= a or b;
    layer8_outputs(5691) <= a and not b;
    layer8_outputs(5692) <= a and not b;
    layer8_outputs(5693) <= not a or b;
    layer8_outputs(5694) <= a and not b;
    layer8_outputs(5695) <= not (a xor b);
    layer8_outputs(5696) <= not (a xor b);
    layer8_outputs(5697) <= '1';
    layer8_outputs(5698) <= not b;
    layer8_outputs(5699) <= b;
    layer8_outputs(5700) <= not b;
    layer8_outputs(5701) <= a;
    layer8_outputs(5702) <= b;
    layer8_outputs(5703) <= a xor b;
    layer8_outputs(5704) <= not b;
    layer8_outputs(5705) <= b;
    layer8_outputs(5706) <= a and b;
    layer8_outputs(5707) <= not (a or b);
    layer8_outputs(5708) <= not a;
    layer8_outputs(5709) <= not b;
    layer8_outputs(5710) <= a or b;
    layer8_outputs(5711) <= a;
    layer8_outputs(5712) <= b;
    layer8_outputs(5713) <= not (a and b);
    layer8_outputs(5714) <= not (a or b);
    layer8_outputs(5715) <= b;
    layer8_outputs(5716) <= not (a xor b);
    layer8_outputs(5717) <= a;
    layer8_outputs(5718) <= a and not b;
    layer8_outputs(5719) <= not b;
    layer8_outputs(5720) <= not a;
    layer8_outputs(5721) <= a xor b;
    layer8_outputs(5722) <= a and b;
    layer8_outputs(5723) <= not b or a;
    layer8_outputs(5724) <= a;
    layer8_outputs(5725) <= not (a or b);
    layer8_outputs(5726) <= not b;
    layer8_outputs(5727) <= b and not a;
    layer8_outputs(5728) <= a;
    layer8_outputs(5729) <= not b;
    layer8_outputs(5730) <= a and b;
    layer8_outputs(5731) <= not (a xor b);
    layer8_outputs(5732) <= not a or b;
    layer8_outputs(5733) <= not b;
    layer8_outputs(5734) <= not b or a;
    layer8_outputs(5735) <= a xor b;
    layer8_outputs(5736) <= a xor b;
    layer8_outputs(5737) <= not (a xor b);
    layer8_outputs(5738) <= not a;
    layer8_outputs(5739) <= b;
    layer8_outputs(5740) <= a or b;
    layer8_outputs(5741) <= not b;
    layer8_outputs(5742) <= b;
    layer8_outputs(5743) <= not (a or b);
    layer8_outputs(5744) <= a or b;
    layer8_outputs(5745) <= b and not a;
    layer8_outputs(5746) <= not b or a;
    layer8_outputs(5747) <= not b;
    layer8_outputs(5748) <= not a;
    layer8_outputs(5749) <= not b or a;
    layer8_outputs(5750) <= not a;
    layer8_outputs(5751) <= a and not b;
    layer8_outputs(5752) <= not b;
    layer8_outputs(5753) <= not (a and b);
    layer8_outputs(5754) <= a;
    layer8_outputs(5755) <= not b;
    layer8_outputs(5756) <= not a;
    layer8_outputs(5757) <= a and not b;
    layer8_outputs(5758) <= not b;
    layer8_outputs(5759) <= not (a xor b);
    layer8_outputs(5760) <= a;
    layer8_outputs(5761) <= b and not a;
    layer8_outputs(5762) <= not b;
    layer8_outputs(5763) <= not b;
    layer8_outputs(5764) <= a and b;
    layer8_outputs(5765) <= b;
    layer8_outputs(5766) <= a and b;
    layer8_outputs(5767) <= not a or b;
    layer8_outputs(5768) <= b;
    layer8_outputs(5769) <= b;
    layer8_outputs(5770) <= b and not a;
    layer8_outputs(5771) <= a xor b;
    layer8_outputs(5772) <= not a;
    layer8_outputs(5773) <= not (a xor b);
    layer8_outputs(5774) <= a and b;
    layer8_outputs(5775) <= a;
    layer8_outputs(5776) <= not b;
    layer8_outputs(5777) <= b and not a;
    layer8_outputs(5778) <= not b;
    layer8_outputs(5779) <= not (a xor b);
    layer8_outputs(5780) <= not b;
    layer8_outputs(5781) <= not a;
    layer8_outputs(5782) <= a and b;
    layer8_outputs(5783) <= a;
    layer8_outputs(5784) <= not b;
    layer8_outputs(5785) <= not a;
    layer8_outputs(5786) <= a;
    layer8_outputs(5787) <= not a or b;
    layer8_outputs(5788) <= not (a or b);
    layer8_outputs(5789) <= a xor b;
    layer8_outputs(5790) <= not (a or b);
    layer8_outputs(5791) <= not (a or b);
    layer8_outputs(5792) <= not a;
    layer8_outputs(5793) <= not a;
    layer8_outputs(5794) <= b and not a;
    layer8_outputs(5795) <= a;
    layer8_outputs(5796) <= a;
    layer8_outputs(5797) <= a;
    layer8_outputs(5798) <= not a or b;
    layer8_outputs(5799) <= not b;
    layer8_outputs(5800) <= not (a xor b);
    layer8_outputs(5801) <= not (a xor b);
    layer8_outputs(5802) <= a;
    layer8_outputs(5803) <= a;
    layer8_outputs(5804) <= b;
    layer8_outputs(5805) <= a xor b;
    layer8_outputs(5806) <= a xor b;
    layer8_outputs(5807) <= b;
    layer8_outputs(5808) <= not a;
    layer8_outputs(5809) <= not (a xor b);
    layer8_outputs(5810) <= not b;
    layer8_outputs(5811) <= not (a xor b);
    layer8_outputs(5812) <= not (a and b);
    layer8_outputs(5813) <= not a;
    layer8_outputs(5814) <= not a;
    layer8_outputs(5815) <= not a;
    layer8_outputs(5816) <= a;
    layer8_outputs(5817) <= a xor b;
    layer8_outputs(5818) <= not a;
    layer8_outputs(5819) <= a xor b;
    layer8_outputs(5820) <= not b;
    layer8_outputs(5821) <= not a or b;
    layer8_outputs(5822) <= not a or b;
    layer8_outputs(5823) <= a or b;
    layer8_outputs(5824) <= not a;
    layer8_outputs(5825) <= '0';
    layer8_outputs(5826) <= a or b;
    layer8_outputs(5827) <= not a;
    layer8_outputs(5828) <= a;
    layer8_outputs(5829) <= not b;
    layer8_outputs(5830) <= a xor b;
    layer8_outputs(5831) <= b;
    layer8_outputs(5832) <= not b or a;
    layer8_outputs(5833) <= a;
    layer8_outputs(5834) <= a xor b;
    layer8_outputs(5835) <= a and b;
    layer8_outputs(5836) <= not (a and b);
    layer8_outputs(5837) <= not a or b;
    layer8_outputs(5838) <= a;
    layer8_outputs(5839) <= b;
    layer8_outputs(5840) <= b;
    layer8_outputs(5841) <= a and not b;
    layer8_outputs(5842) <= not (a or b);
    layer8_outputs(5843) <= b;
    layer8_outputs(5844) <= not b or a;
    layer8_outputs(5845) <= a or b;
    layer8_outputs(5846) <= not b or a;
    layer8_outputs(5847) <= a;
    layer8_outputs(5848) <= a xor b;
    layer8_outputs(5849) <= a xor b;
    layer8_outputs(5850) <= b;
    layer8_outputs(5851) <= a;
    layer8_outputs(5852) <= a or b;
    layer8_outputs(5853) <= not b;
    layer8_outputs(5854) <= not b;
    layer8_outputs(5855) <= a;
    layer8_outputs(5856) <= b and not a;
    layer8_outputs(5857) <= a;
    layer8_outputs(5858) <= a;
    layer8_outputs(5859) <= not (a xor b);
    layer8_outputs(5860) <= a or b;
    layer8_outputs(5861) <= b;
    layer8_outputs(5862) <= a;
    layer8_outputs(5863) <= a or b;
    layer8_outputs(5864) <= a xor b;
    layer8_outputs(5865) <= a xor b;
    layer8_outputs(5866) <= a;
    layer8_outputs(5867) <= not (a or b);
    layer8_outputs(5868) <= not (a xor b);
    layer8_outputs(5869) <= a and not b;
    layer8_outputs(5870) <= not b;
    layer8_outputs(5871) <= not a;
    layer8_outputs(5872) <= a or b;
    layer8_outputs(5873) <= a;
    layer8_outputs(5874) <= not (a xor b);
    layer8_outputs(5875) <= not (a or b);
    layer8_outputs(5876) <= not a;
    layer8_outputs(5877) <= a or b;
    layer8_outputs(5878) <= b and not a;
    layer8_outputs(5879) <= a xor b;
    layer8_outputs(5880) <= not a;
    layer8_outputs(5881) <= not (a xor b);
    layer8_outputs(5882) <= not (a and b);
    layer8_outputs(5883) <= not b or a;
    layer8_outputs(5884) <= not a;
    layer8_outputs(5885) <= not a or b;
    layer8_outputs(5886) <= b and not a;
    layer8_outputs(5887) <= b;
    layer8_outputs(5888) <= not a or b;
    layer8_outputs(5889) <= not (a xor b);
    layer8_outputs(5890) <= not (a or b);
    layer8_outputs(5891) <= not (a xor b);
    layer8_outputs(5892) <= a or b;
    layer8_outputs(5893) <= not a;
    layer8_outputs(5894) <= not (a and b);
    layer8_outputs(5895) <= a and not b;
    layer8_outputs(5896) <= not (a and b);
    layer8_outputs(5897) <= not a;
    layer8_outputs(5898) <= not b or a;
    layer8_outputs(5899) <= not a;
    layer8_outputs(5900) <= a or b;
    layer8_outputs(5901) <= a or b;
    layer8_outputs(5902) <= not a;
    layer8_outputs(5903) <= a;
    layer8_outputs(5904) <= not (a xor b);
    layer8_outputs(5905) <= b;
    layer8_outputs(5906) <= not (a or b);
    layer8_outputs(5907) <= not (a and b);
    layer8_outputs(5908) <= not b or a;
    layer8_outputs(5909) <= b;
    layer8_outputs(5910) <= not a;
    layer8_outputs(5911) <= not (a or b);
    layer8_outputs(5912) <= a and not b;
    layer8_outputs(5913) <= a or b;
    layer8_outputs(5914) <= a;
    layer8_outputs(5915) <= not a;
    layer8_outputs(5916) <= a or b;
    layer8_outputs(5917) <= not a;
    layer8_outputs(5918) <= a and not b;
    layer8_outputs(5919) <= not (a xor b);
    layer8_outputs(5920) <= not b or a;
    layer8_outputs(5921) <= a;
    layer8_outputs(5922) <= not a;
    layer8_outputs(5923) <= not a;
    layer8_outputs(5924) <= not a;
    layer8_outputs(5925) <= not b;
    layer8_outputs(5926) <= not (a xor b);
    layer8_outputs(5927) <= not (a xor b);
    layer8_outputs(5928) <= not a;
    layer8_outputs(5929) <= not a;
    layer8_outputs(5930) <= not b;
    layer8_outputs(5931) <= not (a xor b);
    layer8_outputs(5932) <= not (a or b);
    layer8_outputs(5933) <= b;
    layer8_outputs(5934) <= not b or a;
    layer8_outputs(5935) <= b;
    layer8_outputs(5936) <= '0';
    layer8_outputs(5937) <= a xor b;
    layer8_outputs(5938) <= not a or b;
    layer8_outputs(5939) <= not (a or b);
    layer8_outputs(5940) <= not b or a;
    layer8_outputs(5941) <= b and not a;
    layer8_outputs(5942) <= b;
    layer8_outputs(5943) <= not a;
    layer8_outputs(5944) <= not (a xor b);
    layer8_outputs(5945) <= a xor b;
    layer8_outputs(5946) <= a and not b;
    layer8_outputs(5947) <= not a;
    layer8_outputs(5948) <= not b;
    layer8_outputs(5949) <= a and b;
    layer8_outputs(5950) <= not b;
    layer8_outputs(5951) <= not a;
    layer8_outputs(5952) <= a;
    layer8_outputs(5953) <= not b or a;
    layer8_outputs(5954) <= b and not a;
    layer8_outputs(5955) <= a or b;
    layer8_outputs(5956) <= b;
    layer8_outputs(5957) <= not b;
    layer8_outputs(5958) <= b;
    layer8_outputs(5959) <= a xor b;
    layer8_outputs(5960) <= not b;
    layer8_outputs(5961) <= a xor b;
    layer8_outputs(5962) <= a;
    layer8_outputs(5963) <= b and not a;
    layer8_outputs(5964) <= not (a xor b);
    layer8_outputs(5965) <= a xor b;
    layer8_outputs(5966) <= not b;
    layer8_outputs(5967) <= a xor b;
    layer8_outputs(5968) <= not (a or b);
    layer8_outputs(5969) <= b;
    layer8_outputs(5970) <= not (a xor b);
    layer8_outputs(5971) <= a;
    layer8_outputs(5972) <= a or b;
    layer8_outputs(5973) <= not (a and b);
    layer8_outputs(5974) <= a xor b;
    layer8_outputs(5975) <= not a or b;
    layer8_outputs(5976) <= a or b;
    layer8_outputs(5977) <= a and not b;
    layer8_outputs(5978) <= b;
    layer8_outputs(5979) <= not b;
    layer8_outputs(5980) <= not (a xor b);
    layer8_outputs(5981) <= not a;
    layer8_outputs(5982) <= not a;
    layer8_outputs(5983) <= b;
    layer8_outputs(5984) <= not b;
    layer8_outputs(5985) <= a and b;
    layer8_outputs(5986) <= not (a xor b);
    layer8_outputs(5987) <= not b;
    layer8_outputs(5988) <= not a;
    layer8_outputs(5989) <= not b;
    layer8_outputs(5990) <= a;
    layer8_outputs(5991) <= a;
    layer8_outputs(5992) <= not a;
    layer8_outputs(5993) <= not a;
    layer8_outputs(5994) <= not b or a;
    layer8_outputs(5995) <= not (a or b);
    layer8_outputs(5996) <= a and not b;
    layer8_outputs(5997) <= not (a xor b);
    layer8_outputs(5998) <= not (a or b);
    layer8_outputs(5999) <= '1';
    layer8_outputs(6000) <= a xor b;
    layer8_outputs(6001) <= b and not a;
    layer8_outputs(6002) <= not b or a;
    layer8_outputs(6003) <= a and not b;
    layer8_outputs(6004) <= b and not a;
    layer8_outputs(6005) <= not a;
    layer8_outputs(6006) <= a;
    layer8_outputs(6007) <= a xor b;
    layer8_outputs(6008) <= not (a and b);
    layer8_outputs(6009) <= not b or a;
    layer8_outputs(6010) <= a and b;
    layer8_outputs(6011) <= a xor b;
    layer8_outputs(6012) <= not (a xor b);
    layer8_outputs(6013) <= b;
    layer8_outputs(6014) <= not a;
    layer8_outputs(6015) <= not b or a;
    layer8_outputs(6016) <= not b;
    layer8_outputs(6017) <= a and not b;
    layer8_outputs(6018) <= not a;
    layer8_outputs(6019) <= b;
    layer8_outputs(6020) <= not a;
    layer8_outputs(6021) <= not b;
    layer8_outputs(6022) <= a;
    layer8_outputs(6023) <= not (a xor b);
    layer8_outputs(6024) <= not a;
    layer8_outputs(6025) <= not a;
    layer8_outputs(6026) <= not b;
    layer8_outputs(6027) <= a xor b;
    layer8_outputs(6028) <= not b;
    layer8_outputs(6029) <= a xor b;
    layer8_outputs(6030) <= a and not b;
    layer8_outputs(6031) <= not a or b;
    layer8_outputs(6032) <= not (a or b);
    layer8_outputs(6033) <= b;
    layer8_outputs(6034) <= not a;
    layer8_outputs(6035) <= not b;
    layer8_outputs(6036) <= a and not b;
    layer8_outputs(6037) <= b;
    layer8_outputs(6038) <= not a;
    layer8_outputs(6039) <= not (a and b);
    layer8_outputs(6040) <= b;
    layer8_outputs(6041) <= not a;
    layer8_outputs(6042) <= not a;
    layer8_outputs(6043) <= b;
    layer8_outputs(6044) <= not (a or b);
    layer8_outputs(6045) <= a;
    layer8_outputs(6046) <= not b;
    layer8_outputs(6047) <= a and b;
    layer8_outputs(6048) <= not a or b;
    layer8_outputs(6049) <= not a or b;
    layer8_outputs(6050) <= a xor b;
    layer8_outputs(6051) <= a and not b;
    layer8_outputs(6052) <= a or b;
    layer8_outputs(6053) <= a xor b;
    layer8_outputs(6054) <= not b;
    layer8_outputs(6055) <= not (a xor b);
    layer8_outputs(6056) <= a and b;
    layer8_outputs(6057) <= not b or a;
    layer8_outputs(6058) <= b;
    layer8_outputs(6059) <= not (a xor b);
    layer8_outputs(6060) <= a xor b;
    layer8_outputs(6061) <= not a;
    layer8_outputs(6062) <= not b;
    layer8_outputs(6063) <= not b;
    layer8_outputs(6064) <= not a;
    layer8_outputs(6065) <= b;
    layer8_outputs(6066) <= not b;
    layer8_outputs(6067) <= a and not b;
    layer8_outputs(6068) <= not (a xor b);
    layer8_outputs(6069) <= a;
    layer8_outputs(6070) <= not (a xor b);
    layer8_outputs(6071) <= b;
    layer8_outputs(6072) <= not b;
    layer8_outputs(6073) <= a and b;
    layer8_outputs(6074) <= a or b;
    layer8_outputs(6075) <= not a;
    layer8_outputs(6076) <= a xor b;
    layer8_outputs(6077) <= not a;
    layer8_outputs(6078) <= b;
    layer8_outputs(6079) <= not (a xor b);
    layer8_outputs(6080) <= a;
    layer8_outputs(6081) <= not (a xor b);
    layer8_outputs(6082) <= a;
    layer8_outputs(6083) <= a or b;
    layer8_outputs(6084) <= not a;
    layer8_outputs(6085) <= a;
    layer8_outputs(6086) <= not (a and b);
    layer8_outputs(6087) <= not (a xor b);
    layer8_outputs(6088) <= not (a and b);
    layer8_outputs(6089) <= a xor b;
    layer8_outputs(6090) <= a;
    layer8_outputs(6091) <= not (a xor b);
    layer8_outputs(6092) <= not a;
    layer8_outputs(6093) <= not (a xor b);
    layer8_outputs(6094) <= not a;
    layer8_outputs(6095) <= a xor b;
    layer8_outputs(6096) <= not a;
    layer8_outputs(6097) <= not a or b;
    layer8_outputs(6098) <= not b;
    layer8_outputs(6099) <= a and not b;
    layer8_outputs(6100) <= not (a xor b);
    layer8_outputs(6101) <= a;
    layer8_outputs(6102) <= a or b;
    layer8_outputs(6103) <= a or b;
    layer8_outputs(6104) <= not b;
    layer8_outputs(6105) <= b;
    layer8_outputs(6106) <= not a or b;
    layer8_outputs(6107) <= not (a and b);
    layer8_outputs(6108) <= not (a and b);
    layer8_outputs(6109) <= not (a xor b);
    layer8_outputs(6110) <= not (a xor b);
    layer8_outputs(6111) <= not (a or b);
    layer8_outputs(6112) <= not a;
    layer8_outputs(6113) <= b;
    layer8_outputs(6114) <= b;
    layer8_outputs(6115) <= not (a xor b);
    layer8_outputs(6116) <= a and not b;
    layer8_outputs(6117) <= not b;
    layer8_outputs(6118) <= not (a and b);
    layer8_outputs(6119) <= not b;
    layer8_outputs(6120) <= a;
    layer8_outputs(6121) <= not (a xor b);
    layer8_outputs(6122) <= not a;
    layer8_outputs(6123) <= a xor b;
    layer8_outputs(6124) <= a or b;
    layer8_outputs(6125) <= not (a or b);
    layer8_outputs(6126) <= a xor b;
    layer8_outputs(6127) <= a xor b;
    layer8_outputs(6128) <= not (a or b);
    layer8_outputs(6129) <= not (a xor b);
    layer8_outputs(6130) <= a xor b;
    layer8_outputs(6131) <= not (a and b);
    layer8_outputs(6132) <= not (a and b);
    layer8_outputs(6133) <= not (a and b);
    layer8_outputs(6134) <= a;
    layer8_outputs(6135) <= a and b;
    layer8_outputs(6136) <= not a;
    layer8_outputs(6137) <= not a;
    layer8_outputs(6138) <= not (a and b);
    layer8_outputs(6139) <= not a;
    layer8_outputs(6140) <= not a;
    layer8_outputs(6141) <= b and not a;
    layer8_outputs(6142) <= not (a xor b);
    layer8_outputs(6143) <= a and b;
    layer8_outputs(6144) <= a xor b;
    layer8_outputs(6145) <= not b;
    layer8_outputs(6146) <= a xor b;
    layer8_outputs(6147) <= a xor b;
    layer8_outputs(6148) <= not a;
    layer8_outputs(6149) <= a and b;
    layer8_outputs(6150) <= a xor b;
    layer8_outputs(6151) <= not (a and b);
    layer8_outputs(6152) <= not (a xor b);
    layer8_outputs(6153) <= not b;
    layer8_outputs(6154) <= not a or b;
    layer8_outputs(6155) <= a xor b;
    layer8_outputs(6156) <= b;
    layer8_outputs(6157) <= a xor b;
    layer8_outputs(6158) <= b and not a;
    layer8_outputs(6159) <= not (a or b);
    layer8_outputs(6160) <= a xor b;
    layer8_outputs(6161) <= a xor b;
    layer8_outputs(6162) <= b;
    layer8_outputs(6163) <= not (a xor b);
    layer8_outputs(6164) <= a xor b;
    layer8_outputs(6165) <= a or b;
    layer8_outputs(6166) <= b and not a;
    layer8_outputs(6167) <= a or b;
    layer8_outputs(6168) <= not (a and b);
    layer8_outputs(6169) <= a;
    layer8_outputs(6170) <= b and not a;
    layer8_outputs(6171) <= not a;
    layer8_outputs(6172) <= not a or b;
    layer8_outputs(6173) <= a xor b;
    layer8_outputs(6174) <= a and not b;
    layer8_outputs(6175) <= not b or a;
    layer8_outputs(6176) <= b;
    layer8_outputs(6177) <= a xor b;
    layer8_outputs(6178) <= b;
    layer8_outputs(6179) <= not b;
    layer8_outputs(6180) <= a xor b;
    layer8_outputs(6181) <= a and b;
    layer8_outputs(6182) <= b;
    layer8_outputs(6183) <= not b or a;
    layer8_outputs(6184) <= not b;
    layer8_outputs(6185) <= not a or b;
    layer8_outputs(6186) <= b;
    layer8_outputs(6187) <= a or b;
    layer8_outputs(6188) <= not b;
    layer8_outputs(6189) <= a and not b;
    layer8_outputs(6190) <= not a;
    layer8_outputs(6191) <= b;
    layer8_outputs(6192) <= not (a or b);
    layer8_outputs(6193) <= not (a or b);
    layer8_outputs(6194) <= not a;
    layer8_outputs(6195) <= b;
    layer8_outputs(6196) <= b and not a;
    layer8_outputs(6197) <= not a;
    layer8_outputs(6198) <= not b;
    layer8_outputs(6199) <= a and b;
    layer8_outputs(6200) <= b and not a;
    layer8_outputs(6201) <= b;
    layer8_outputs(6202) <= not b or a;
    layer8_outputs(6203) <= not b;
    layer8_outputs(6204) <= not b;
    layer8_outputs(6205) <= a or b;
    layer8_outputs(6206) <= not (a xor b);
    layer8_outputs(6207) <= b;
    layer8_outputs(6208) <= not b;
    layer8_outputs(6209) <= b and not a;
    layer8_outputs(6210) <= not a or b;
    layer8_outputs(6211) <= a xor b;
    layer8_outputs(6212) <= not b;
    layer8_outputs(6213) <= a;
    layer8_outputs(6214) <= not b;
    layer8_outputs(6215) <= not b;
    layer8_outputs(6216) <= a xor b;
    layer8_outputs(6217) <= a xor b;
    layer8_outputs(6218) <= not (a or b);
    layer8_outputs(6219) <= a or b;
    layer8_outputs(6220) <= a and b;
    layer8_outputs(6221) <= a and b;
    layer8_outputs(6222) <= not a;
    layer8_outputs(6223) <= not (a xor b);
    layer8_outputs(6224) <= not a or b;
    layer8_outputs(6225) <= '0';
    layer8_outputs(6226) <= not (a or b);
    layer8_outputs(6227) <= not b;
    layer8_outputs(6228) <= not b;
    layer8_outputs(6229) <= b;
    layer8_outputs(6230) <= a and not b;
    layer8_outputs(6231) <= a;
    layer8_outputs(6232) <= not a;
    layer8_outputs(6233) <= b;
    layer8_outputs(6234) <= a and b;
    layer8_outputs(6235) <= not (a or b);
    layer8_outputs(6236) <= b;
    layer8_outputs(6237) <= not b;
    layer8_outputs(6238) <= not (a and b);
    layer8_outputs(6239) <= not b;
    layer8_outputs(6240) <= not (a xor b);
    layer8_outputs(6241) <= not a;
    layer8_outputs(6242) <= not a;
    layer8_outputs(6243) <= a;
    layer8_outputs(6244) <= b;
    layer8_outputs(6245) <= not (a or b);
    layer8_outputs(6246) <= b;
    layer8_outputs(6247) <= not a or b;
    layer8_outputs(6248) <= not (a xor b);
    layer8_outputs(6249) <= a;
    layer8_outputs(6250) <= b;
    layer8_outputs(6251) <= not a or b;
    layer8_outputs(6252) <= not b or a;
    layer8_outputs(6253) <= not (a and b);
    layer8_outputs(6254) <= b;
    layer8_outputs(6255) <= not a or b;
    layer8_outputs(6256) <= a;
    layer8_outputs(6257) <= a;
    layer8_outputs(6258) <= not b or a;
    layer8_outputs(6259) <= not b;
    layer8_outputs(6260) <= not (a xor b);
    layer8_outputs(6261) <= a and b;
    layer8_outputs(6262) <= b and not a;
    layer8_outputs(6263) <= a;
    layer8_outputs(6264) <= not a;
    layer8_outputs(6265) <= not (a and b);
    layer8_outputs(6266) <= not (a or b);
    layer8_outputs(6267) <= not a;
    layer8_outputs(6268) <= not b;
    layer8_outputs(6269) <= a and b;
    layer8_outputs(6270) <= a or b;
    layer8_outputs(6271) <= b and not a;
    layer8_outputs(6272) <= a xor b;
    layer8_outputs(6273) <= not b or a;
    layer8_outputs(6274) <= not a or b;
    layer8_outputs(6275) <= a and not b;
    layer8_outputs(6276) <= b and not a;
    layer8_outputs(6277) <= b;
    layer8_outputs(6278) <= a;
    layer8_outputs(6279) <= a xor b;
    layer8_outputs(6280) <= a xor b;
    layer8_outputs(6281) <= b;
    layer8_outputs(6282) <= not b or a;
    layer8_outputs(6283) <= not b;
    layer8_outputs(6284) <= not b;
    layer8_outputs(6285) <= b;
    layer8_outputs(6286) <= not (a xor b);
    layer8_outputs(6287) <= a or b;
    layer8_outputs(6288) <= a or b;
    layer8_outputs(6289) <= not (a or b);
    layer8_outputs(6290) <= not (a xor b);
    layer8_outputs(6291) <= '0';
    layer8_outputs(6292) <= not b;
    layer8_outputs(6293) <= a and b;
    layer8_outputs(6294) <= not (a xor b);
    layer8_outputs(6295) <= a;
    layer8_outputs(6296) <= not b or a;
    layer8_outputs(6297) <= not b or a;
    layer8_outputs(6298) <= not b or a;
    layer8_outputs(6299) <= not a or b;
    layer8_outputs(6300) <= a xor b;
    layer8_outputs(6301) <= a and not b;
    layer8_outputs(6302) <= not (a and b);
    layer8_outputs(6303) <= not a or b;
    layer8_outputs(6304) <= a and not b;
    layer8_outputs(6305) <= b;
    layer8_outputs(6306) <= not (a or b);
    layer8_outputs(6307) <= a and not b;
    layer8_outputs(6308) <= not (a and b);
    layer8_outputs(6309) <= not b;
    layer8_outputs(6310) <= a;
    layer8_outputs(6311) <= not a;
    layer8_outputs(6312) <= b and not a;
    layer8_outputs(6313) <= not b;
    layer8_outputs(6314) <= b;
    layer8_outputs(6315) <= a and b;
    layer8_outputs(6316) <= not (a xor b);
    layer8_outputs(6317) <= not (a xor b);
    layer8_outputs(6318) <= b;
    layer8_outputs(6319) <= a;
    layer8_outputs(6320) <= not (a xor b);
    layer8_outputs(6321) <= a xor b;
    layer8_outputs(6322) <= b and not a;
    layer8_outputs(6323) <= b;
    layer8_outputs(6324) <= not b;
    layer8_outputs(6325) <= not b;
    layer8_outputs(6326) <= a;
    layer8_outputs(6327) <= not a;
    layer8_outputs(6328) <= a and not b;
    layer8_outputs(6329) <= not a;
    layer8_outputs(6330) <= not (a and b);
    layer8_outputs(6331) <= b;
    layer8_outputs(6332) <= b;
    layer8_outputs(6333) <= not b;
    layer8_outputs(6334) <= a or b;
    layer8_outputs(6335) <= b and not a;
    layer8_outputs(6336) <= a and not b;
    layer8_outputs(6337) <= not (a or b);
    layer8_outputs(6338) <= a and b;
    layer8_outputs(6339) <= a or b;
    layer8_outputs(6340) <= not (a or b);
    layer8_outputs(6341) <= not b or a;
    layer8_outputs(6342) <= not b;
    layer8_outputs(6343) <= b and not a;
    layer8_outputs(6344) <= not (a or b);
    layer8_outputs(6345) <= a xor b;
    layer8_outputs(6346) <= b and not a;
    layer8_outputs(6347) <= b;
    layer8_outputs(6348) <= a xor b;
    layer8_outputs(6349) <= not b;
    layer8_outputs(6350) <= not b;
    layer8_outputs(6351) <= not a;
    layer8_outputs(6352) <= b;
    layer8_outputs(6353) <= a;
    layer8_outputs(6354) <= b;
    layer8_outputs(6355) <= not (a xor b);
    layer8_outputs(6356) <= not (a and b);
    layer8_outputs(6357) <= a and b;
    layer8_outputs(6358) <= not (a and b);
    layer8_outputs(6359) <= not b;
    layer8_outputs(6360) <= not (a xor b);
    layer8_outputs(6361) <= not b;
    layer8_outputs(6362) <= not (a xor b);
    layer8_outputs(6363) <= not b;
    layer8_outputs(6364) <= a;
    layer8_outputs(6365) <= not (a xor b);
    layer8_outputs(6366) <= not (a xor b);
    layer8_outputs(6367) <= not (a xor b);
    layer8_outputs(6368) <= not a;
    layer8_outputs(6369) <= b;
    layer8_outputs(6370) <= b;
    layer8_outputs(6371) <= not (a xor b);
    layer8_outputs(6372) <= not a or b;
    layer8_outputs(6373) <= not (a or b);
    layer8_outputs(6374) <= a xor b;
    layer8_outputs(6375) <= not b;
    layer8_outputs(6376) <= a xor b;
    layer8_outputs(6377) <= a xor b;
    layer8_outputs(6378) <= not a;
    layer8_outputs(6379) <= not a;
    layer8_outputs(6380) <= not a;
    layer8_outputs(6381) <= not a;
    layer8_outputs(6382) <= not a or b;
    layer8_outputs(6383) <= a xor b;
    layer8_outputs(6384) <= b and not a;
    layer8_outputs(6385) <= not b;
    layer8_outputs(6386) <= a xor b;
    layer8_outputs(6387) <= a and not b;
    layer8_outputs(6388) <= not a;
    layer8_outputs(6389) <= a or b;
    layer8_outputs(6390) <= a;
    layer8_outputs(6391) <= not (a xor b);
    layer8_outputs(6392) <= a;
    layer8_outputs(6393) <= a;
    layer8_outputs(6394) <= not a;
    layer8_outputs(6395) <= a;
    layer8_outputs(6396) <= a;
    layer8_outputs(6397) <= not b;
    layer8_outputs(6398) <= b;
    layer8_outputs(6399) <= not (a or b);
    layer8_outputs(6400) <= not a;
    layer8_outputs(6401) <= a;
    layer8_outputs(6402) <= a and not b;
    layer8_outputs(6403) <= a xor b;
    layer8_outputs(6404) <= a;
    layer8_outputs(6405) <= not a;
    layer8_outputs(6406) <= a;
    layer8_outputs(6407) <= not (a xor b);
    layer8_outputs(6408) <= not (a xor b);
    layer8_outputs(6409) <= not (a and b);
    layer8_outputs(6410) <= b and not a;
    layer8_outputs(6411) <= not b;
    layer8_outputs(6412) <= not a;
    layer8_outputs(6413) <= not (a xor b);
    layer8_outputs(6414) <= not b;
    layer8_outputs(6415) <= a and not b;
    layer8_outputs(6416) <= b and not a;
    layer8_outputs(6417) <= b;
    layer8_outputs(6418) <= b;
    layer8_outputs(6419) <= not (a xor b);
    layer8_outputs(6420) <= b;
    layer8_outputs(6421) <= a;
    layer8_outputs(6422) <= b;
    layer8_outputs(6423) <= not b;
    layer8_outputs(6424) <= b;
    layer8_outputs(6425) <= not (a and b);
    layer8_outputs(6426) <= b;
    layer8_outputs(6427) <= a;
    layer8_outputs(6428) <= not b or a;
    layer8_outputs(6429) <= b and not a;
    layer8_outputs(6430) <= not b;
    layer8_outputs(6431) <= a or b;
    layer8_outputs(6432) <= not b;
    layer8_outputs(6433) <= not b;
    layer8_outputs(6434) <= b;
    layer8_outputs(6435) <= a and b;
    layer8_outputs(6436) <= a;
    layer8_outputs(6437) <= a or b;
    layer8_outputs(6438) <= not b;
    layer8_outputs(6439) <= not (a or b);
    layer8_outputs(6440) <= a and b;
    layer8_outputs(6441) <= not (a and b);
    layer8_outputs(6442) <= a;
    layer8_outputs(6443) <= not b;
    layer8_outputs(6444) <= not b;
    layer8_outputs(6445) <= not a or b;
    layer8_outputs(6446) <= b;
    layer8_outputs(6447) <= a;
    layer8_outputs(6448) <= a and b;
    layer8_outputs(6449) <= b and not a;
    layer8_outputs(6450) <= a;
    layer8_outputs(6451) <= not (a or b);
    layer8_outputs(6452) <= not a;
    layer8_outputs(6453) <= b and not a;
    layer8_outputs(6454) <= not (a xor b);
    layer8_outputs(6455) <= a;
    layer8_outputs(6456) <= not a or b;
    layer8_outputs(6457) <= b and not a;
    layer8_outputs(6458) <= not a;
    layer8_outputs(6459) <= not b;
    layer8_outputs(6460) <= not (a and b);
    layer8_outputs(6461) <= a or b;
    layer8_outputs(6462) <= not (a xor b);
    layer8_outputs(6463) <= a and not b;
    layer8_outputs(6464) <= a;
    layer8_outputs(6465) <= b;
    layer8_outputs(6466) <= not b;
    layer8_outputs(6467) <= a and b;
    layer8_outputs(6468) <= not a;
    layer8_outputs(6469) <= not (a and b);
    layer8_outputs(6470) <= b;
    layer8_outputs(6471) <= a and b;
    layer8_outputs(6472) <= a or b;
    layer8_outputs(6473) <= not a;
    layer8_outputs(6474) <= a or b;
    layer8_outputs(6475) <= not a;
    layer8_outputs(6476) <= b and not a;
    layer8_outputs(6477) <= not (a xor b);
    layer8_outputs(6478) <= a;
    layer8_outputs(6479) <= a;
    layer8_outputs(6480) <= not (a and b);
    layer8_outputs(6481) <= not a or b;
    layer8_outputs(6482) <= not b;
    layer8_outputs(6483) <= b and not a;
    layer8_outputs(6484) <= not (a xor b);
    layer8_outputs(6485) <= not b;
    layer8_outputs(6486) <= a;
    layer8_outputs(6487) <= not (a xor b);
    layer8_outputs(6488) <= a and b;
    layer8_outputs(6489) <= b;
    layer8_outputs(6490) <= a;
    layer8_outputs(6491) <= a and b;
    layer8_outputs(6492) <= a xor b;
    layer8_outputs(6493) <= not (a or b);
    layer8_outputs(6494) <= not (a or b);
    layer8_outputs(6495) <= a and not b;
    layer8_outputs(6496) <= not b;
    layer8_outputs(6497) <= a xor b;
    layer8_outputs(6498) <= a and not b;
    layer8_outputs(6499) <= not (a xor b);
    layer8_outputs(6500) <= b and not a;
    layer8_outputs(6501) <= a and b;
    layer8_outputs(6502) <= not a;
    layer8_outputs(6503) <= not b;
    layer8_outputs(6504) <= not (a xor b);
    layer8_outputs(6505) <= a or b;
    layer8_outputs(6506) <= a and b;
    layer8_outputs(6507) <= a xor b;
    layer8_outputs(6508) <= not a;
    layer8_outputs(6509) <= not b;
    layer8_outputs(6510) <= not a;
    layer8_outputs(6511) <= not b or a;
    layer8_outputs(6512) <= a xor b;
    layer8_outputs(6513) <= not b;
    layer8_outputs(6514) <= not a;
    layer8_outputs(6515) <= not (a xor b);
    layer8_outputs(6516) <= not a;
    layer8_outputs(6517) <= not (a and b);
    layer8_outputs(6518) <= b;
    layer8_outputs(6519) <= a or b;
    layer8_outputs(6520) <= not b;
    layer8_outputs(6521) <= a;
    layer8_outputs(6522) <= not (a and b);
    layer8_outputs(6523) <= not b or a;
    layer8_outputs(6524) <= a;
    layer8_outputs(6525) <= a and b;
    layer8_outputs(6526) <= not b;
    layer8_outputs(6527) <= not (a or b);
    layer8_outputs(6528) <= '0';
    layer8_outputs(6529) <= not (a xor b);
    layer8_outputs(6530) <= not b;
    layer8_outputs(6531) <= not a or b;
    layer8_outputs(6532) <= b and not a;
    layer8_outputs(6533) <= b;
    layer8_outputs(6534) <= not (a and b);
    layer8_outputs(6535) <= a xor b;
    layer8_outputs(6536) <= not b or a;
    layer8_outputs(6537) <= not a;
    layer8_outputs(6538) <= a xor b;
    layer8_outputs(6539) <= not b or a;
    layer8_outputs(6540) <= a;
    layer8_outputs(6541) <= not (a xor b);
    layer8_outputs(6542) <= not (a xor b);
    layer8_outputs(6543) <= not b;
    layer8_outputs(6544) <= not b;
    layer8_outputs(6545) <= b;
    layer8_outputs(6546) <= not a;
    layer8_outputs(6547) <= not b or a;
    layer8_outputs(6548) <= not b;
    layer8_outputs(6549) <= not b or a;
    layer8_outputs(6550) <= a or b;
    layer8_outputs(6551) <= not (a or b);
    layer8_outputs(6552) <= not a;
    layer8_outputs(6553) <= a and b;
    layer8_outputs(6554) <= a and b;
    layer8_outputs(6555) <= not (a and b);
    layer8_outputs(6556) <= not a;
    layer8_outputs(6557) <= a;
    layer8_outputs(6558) <= b and not a;
    layer8_outputs(6559) <= not b;
    layer8_outputs(6560) <= not b;
    layer8_outputs(6561) <= not a;
    layer8_outputs(6562) <= b;
    layer8_outputs(6563) <= not (a or b);
    layer8_outputs(6564) <= a xor b;
    layer8_outputs(6565) <= a and b;
    layer8_outputs(6566) <= not a;
    layer8_outputs(6567) <= not (a xor b);
    layer8_outputs(6568) <= not b;
    layer8_outputs(6569) <= a or b;
    layer8_outputs(6570) <= not a or b;
    layer8_outputs(6571) <= not (a or b);
    layer8_outputs(6572) <= not b or a;
    layer8_outputs(6573) <= not (a xor b);
    layer8_outputs(6574) <= not (a xor b);
    layer8_outputs(6575) <= not b or a;
    layer8_outputs(6576) <= b and not a;
    layer8_outputs(6577) <= a;
    layer8_outputs(6578) <= not b;
    layer8_outputs(6579) <= a and b;
    layer8_outputs(6580) <= a and not b;
    layer8_outputs(6581) <= not b;
    layer8_outputs(6582) <= not a;
    layer8_outputs(6583) <= not (a xor b);
    layer8_outputs(6584) <= a and b;
    layer8_outputs(6585) <= b;
    layer8_outputs(6586) <= b and not a;
    layer8_outputs(6587) <= not b;
    layer8_outputs(6588) <= not (a xor b);
    layer8_outputs(6589) <= not b;
    layer8_outputs(6590) <= not a;
    layer8_outputs(6591) <= not a;
    layer8_outputs(6592) <= a xor b;
    layer8_outputs(6593) <= not a;
    layer8_outputs(6594) <= not b;
    layer8_outputs(6595) <= not b;
    layer8_outputs(6596) <= b;
    layer8_outputs(6597) <= not (a or b);
    layer8_outputs(6598) <= a and b;
    layer8_outputs(6599) <= not (a xor b);
    layer8_outputs(6600) <= not b;
    layer8_outputs(6601) <= b and not a;
    layer8_outputs(6602) <= b;
    layer8_outputs(6603) <= not a or b;
    layer8_outputs(6604) <= a;
    layer8_outputs(6605) <= a xor b;
    layer8_outputs(6606) <= a xor b;
    layer8_outputs(6607) <= a xor b;
    layer8_outputs(6608) <= a and b;
    layer8_outputs(6609) <= a;
    layer8_outputs(6610) <= not a;
    layer8_outputs(6611) <= not b;
    layer8_outputs(6612) <= not (a or b);
    layer8_outputs(6613) <= a;
    layer8_outputs(6614) <= a or b;
    layer8_outputs(6615) <= not (a xor b);
    layer8_outputs(6616) <= a or b;
    layer8_outputs(6617) <= b;
    layer8_outputs(6618) <= a xor b;
    layer8_outputs(6619) <= not (a xor b);
    layer8_outputs(6620) <= not b;
    layer8_outputs(6621) <= a or b;
    layer8_outputs(6622) <= a xor b;
    layer8_outputs(6623) <= not a or b;
    layer8_outputs(6624) <= b;
    layer8_outputs(6625) <= not b;
    layer8_outputs(6626) <= not a;
    layer8_outputs(6627) <= not b;
    layer8_outputs(6628) <= b;
    layer8_outputs(6629) <= a;
    layer8_outputs(6630) <= not (a xor b);
    layer8_outputs(6631) <= b;
    layer8_outputs(6632) <= b;
    layer8_outputs(6633) <= not b;
    layer8_outputs(6634) <= not a or b;
    layer8_outputs(6635) <= not a;
    layer8_outputs(6636) <= a and not b;
    layer8_outputs(6637) <= not a or b;
    layer8_outputs(6638) <= not a;
    layer8_outputs(6639) <= b and not a;
    layer8_outputs(6640) <= not b;
    layer8_outputs(6641) <= not (a xor b);
    layer8_outputs(6642) <= b;
    layer8_outputs(6643) <= not (a xor b);
    layer8_outputs(6644) <= b;
    layer8_outputs(6645) <= a and not b;
    layer8_outputs(6646) <= b;
    layer8_outputs(6647) <= not (a and b);
    layer8_outputs(6648) <= a xor b;
    layer8_outputs(6649) <= not b;
    layer8_outputs(6650) <= a or b;
    layer8_outputs(6651) <= not a or b;
    layer8_outputs(6652) <= a and b;
    layer8_outputs(6653) <= not b;
    layer8_outputs(6654) <= not b or a;
    layer8_outputs(6655) <= not b or a;
    layer8_outputs(6656) <= not (a or b);
    layer8_outputs(6657) <= a xor b;
    layer8_outputs(6658) <= a and b;
    layer8_outputs(6659) <= not b or a;
    layer8_outputs(6660) <= not b;
    layer8_outputs(6661) <= not a;
    layer8_outputs(6662) <= not b or a;
    layer8_outputs(6663) <= a xor b;
    layer8_outputs(6664) <= a and b;
    layer8_outputs(6665) <= b and not a;
    layer8_outputs(6666) <= a xor b;
    layer8_outputs(6667) <= not (a xor b);
    layer8_outputs(6668) <= not a;
    layer8_outputs(6669) <= b and not a;
    layer8_outputs(6670) <= not (a xor b);
    layer8_outputs(6671) <= a;
    layer8_outputs(6672) <= b;
    layer8_outputs(6673) <= not a or b;
    layer8_outputs(6674) <= not b or a;
    layer8_outputs(6675) <= b;
    layer8_outputs(6676) <= not (a or b);
    layer8_outputs(6677) <= a;
    layer8_outputs(6678) <= a;
    layer8_outputs(6679) <= a and b;
    layer8_outputs(6680) <= '1';
    layer8_outputs(6681) <= not (a or b);
    layer8_outputs(6682) <= a;
    layer8_outputs(6683) <= a;
    layer8_outputs(6684) <= not (a or b);
    layer8_outputs(6685) <= not a;
    layer8_outputs(6686) <= b;
    layer8_outputs(6687) <= not a or b;
    layer8_outputs(6688) <= not a;
    layer8_outputs(6689) <= a and not b;
    layer8_outputs(6690) <= a xor b;
    layer8_outputs(6691) <= not (a or b);
    layer8_outputs(6692) <= b;
    layer8_outputs(6693) <= not b;
    layer8_outputs(6694) <= a xor b;
    layer8_outputs(6695) <= not a or b;
    layer8_outputs(6696) <= not a;
    layer8_outputs(6697) <= not b;
    layer8_outputs(6698) <= not b;
    layer8_outputs(6699) <= a xor b;
    layer8_outputs(6700) <= b;
    layer8_outputs(6701) <= not a;
    layer8_outputs(6702) <= b;
    layer8_outputs(6703) <= not a;
    layer8_outputs(6704) <= a xor b;
    layer8_outputs(6705) <= a;
    layer8_outputs(6706) <= not b or a;
    layer8_outputs(6707) <= not (a and b);
    layer8_outputs(6708) <= not a;
    layer8_outputs(6709) <= a and not b;
    layer8_outputs(6710) <= not a or b;
    layer8_outputs(6711) <= a;
    layer8_outputs(6712) <= a or b;
    layer8_outputs(6713) <= not (a or b);
    layer8_outputs(6714) <= a and b;
    layer8_outputs(6715) <= a or b;
    layer8_outputs(6716) <= not b or a;
    layer8_outputs(6717) <= a;
    layer8_outputs(6718) <= not (a xor b);
    layer8_outputs(6719) <= b and not a;
    layer8_outputs(6720) <= not (a xor b);
    layer8_outputs(6721) <= not b or a;
    layer8_outputs(6722) <= b;
    layer8_outputs(6723) <= not (a xor b);
    layer8_outputs(6724) <= not a;
    layer8_outputs(6725) <= not (a xor b);
    layer8_outputs(6726) <= b;
    layer8_outputs(6727) <= a;
    layer8_outputs(6728) <= a;
    layer8_outputs(6729) <= a xor b;
    layer8_outputs(6730) <= not b;
    layer8_outputs(6731) <= a xor b;
    layer8_outputs(6732) <= b and not a;
    layer8_outputs(6733) <= not (a xor b);
    layer8_outputs(6734) <= not b;
    layer8_outputs(6735) <= not (a xor b);
    layer8_outputs(6736) <= not a;
    layer8_outputs(6737) <= not (a xor b);
    layer8_outputs(6738) <= not (a xor b);
    layer8_outputs(6739) <= not (a or b);
    layer8_outputs(6740) <= not (a or b);
    layer8_outputs(6741) <= not (a and b);
    layer8_outputs(6742) <= not (a xor b);
    layer8_outputs(6743) <= a and not b;
    layer8_outputs(6744) <= not (a xor b);
    layer8_outputs(6745) <= a;
    layer8_outputs(6746) <= a and b;
    layer8_outputs(6747) <= a and not b;
    layer8_outputs(6748) <= not (a and b);
    layer8_outputs(6749) <= not b;
    layer8_outputs(6750) <= not a;
    layer8_outputs(6751) <= not b or a;
    layer8_outputs(6752) <= not a;
    layer8_outputs(6753) <= not b;
    layer8_outputs(6754) <= '0';
    layer8_outputs(6755) <= a xor b;
    layer8_outputs(6756) <= not b or a;
    layer8_outputs(6757) <= not (a and b);
    layer8_outputs(6758) <= a;
    layer8_outputs(6759) <= not b;
    layer8_outputs(6760) <= not a;
    layer8_outputs(6761) <= a and b;
    layer8_outputs(6762) <= b;
    layer8_outputs(6763) <= not b;
    layer8_outputs(6764) <= a or b;
    layer8_outputs(6765) <= not a or b;
    layer8_outputs(6766) <= not b;
    layer8_outputs(6767) <= a;
    layer8_outputs(6768) <= a xor b;
    layer8_outputs(6769) <= a;
    layer8_outputs(6770) <= b and not a;
    layer8_outputs(6771) <= a and b;
    layer8_outputs(6772) <= not a or b;
    layer8_outputs(6773) <= not a or b;
    layer8_outputs(6774) <= not a;
    layer8_outputs(6775) <= not a;
    layer8_outputs(6776) <= not b;
    layer8_outputs(6777) <= not (a and b);
    layer8_outputs(6778) <= not b;
    layer8_outputs(6779) <= not a;
    layer8_outputs(6780) <= a and not b;
    layer8_outputs(6781) <= b;
    layer8_outputs(6782) <= not a or b;
    layer8_outputs(6783) <= a;
    layer8_outputs(6784) <= b;
    layer8_outputs(6785) <= a or b;
    layer8_outputs(6786) <= not (a xor b);
    layer8_outputs(6787) <= not b;
    layer8_outputs(6788) <= '1';
    layer8_outputs(6789) <= a xor b;
    layer8_outputs(6790) <= not b;
    layer8_outputs(6791) <= a xor b;
    layer8_outputs(6792) <= not b;
    layer8_outputs(6793) <= not a or b;
    layer8_outputs(6794) <= not (a or b);
    layer8_outputs(6795) <= b;
    layer8_outputs(6796) <= a and b;
    layer8_outputs(6797) <= not (a xor b);
    layer8_outputs(6798) <= b and not a;
    layer8_outputs(6799) <= not a;
    layer8_outputs(6800) <= not b or a;
    layer8_outputs(6801) <= not a or b;
    layer8_outputs(6802) <= a;
    layer8_outputs(6803) <= a;
    layer8_outputs(6804) <= not a;
    layer8_outputs(6805) <= a or b;
    layer8_outputs(6806) <= a and b;
    layer8_outputs(6807) <= not a;
    layer8_outputs(6808) <= b;
    layer8_outputs(6809) <= not a or b;
    layer8_outputs(6810) <= a;
    layer8_outputs(6811) <= not b or a;
    layer8_outputs(6812) <= b;
    layer8_outputs(6813) <= b;
    layer8_outputs(6814) <= a and not b;
    layer8_outputs(6815) <= a xor b;
    layer8_outputs(6816) <= not a;
    layer8_outputs(6817) <= a;
    layer8_outputs(6818) <= b;
    layer8_outputs(6819) <= not a or b;
    layer8_outputs(6820) <= a or b;
    layer8_outputs(6821) <= not a;
    layer8_outputs(6822) <= not (a and b);
    layer8_outputs(6823) <= a and not b;
    layer8_outputs(6824) <= not (a xor b);
    layer8_outputs(6825) <= not b;
    layer8_outputs(6826) <= not b or a;
    layer8_outputs(6827) <= not a;
    layer8_outputs(6828) <= '0';
    layer8_outputs(6829) <= not (a xor b);
    layer8_outputs(6830) <= not (a xor b);
    layer8_outputs(6831) <= not a;
    layer8_outputs(6832) <= not (a or b);
    layer8_outputs(6833) <= not a or b;
    layer8_outputs(6834) <= b and not a;
    layer8_outputs(6835) <= not b or a;
    layer8_outputs(6836) <= a and b;
    layer8_outputs(6837) <= not (a xor b);
    layer8_outputs(6838) <= b;
    layer8_outputs(6839) <= a and not b;
    layer8_outputs(6840) <= b;
    layer8_outputs(6841) <= not b or a;
    layer8_outputs(6842) <= not a or b;
    layer8_outputs(6843) <= a;
    layer8_outputs(6844) <= b;
    layer8_outputs(6845) <= b;
    layer8_outputs(6846) <= a;
    layer8_outputs(6847) <= not b;
    layer8_outputs(6848) <= not b;
    layer8_outputs(6849) <= not a;
    layer8_outputs(6850) <= not a;
    layer8_outputs(6851) <= b and not a;
    layer8_outputs(6852) <= a;
    layer8_outputs(6853) <= not a or b;
    layer8_outputs(6854) <= not a;
    layer8_outputs(6855) <= not (a or b);
    layer8_outputs(6856) <= not (a xor b);
    layer8_outputs(6857) <= not a;
    layer8_outputs(6858) <= not a;
    layer8_outputs(6859) <= b;
    layer8_outputs(6860) <= not b;
    layer8_outputs(6861) <= not b;
    layer8_outputs(6862) <= b;
    layer8_outputs(6863) <= a;
    layer8_outputs(6864) <= not (a xor b);
    layer8_outputs(6865) <= a and not b;
    layer8_outputs(6866) <= not a;
    layer8_outputs(6867) <= a xor b;
    layer8_outputs(6868) <= not a;
    layer8_outputs(6869) <= b and not a;
    layer8_outputs(6870) <= not (a xor b);
    layer8_outputs(6871) <= a xor b;
    layer8_outputs(6872) <= not (a xor b);
    layer8_outputs(6873) <= not a;
    layer8_outputs(6874) <= not a or b;
    layer8_outputs(6875) <= a;
    layer8_outputs(6876) <= a;
    layer8_outputs(6877) <= a and not b;
    layer8_outputs(6878) <= not a or b;
    layer8_outputs(6879) <= not b;
    layer8_outputs(6880) <= not (a xor b);
    layer8_outputs(6881) <= b;
    layer8_outputs(6882) <= not a;
    layer8_outputs(6883) <= a;
    layer8_outputs(6884) <= b;
    layer8_outputs(6885) <= a;
    layer8_outputs(6886) <= not (a or b);
    layer8_outputs(6887) <= not b;
    layer8_outputs(6888) <= a xor b;
    layer8_outputs(6889) <= not b;
    layer8_outputs(6890) <= not b;
    layer8_outputs(6891) <= b and not a;
    layer8_outputs(6892) <= not (a xor b);
    layer8_outputs(6893) <= not (a or b);
    layer8_outputs(6894) <= not (a xor b);
    layer8_outputs(6895) <= not (a xor b);
    layer8_outputs(6896) <= a and not b;
    layer8_outputs(6897) <= b;
    layer8_outputs(6898) <= not (a and b);
    layer8_outputs(6899) <= not (a or b);
    layer8_outputs(6900) <= not (a and b);
    layer8_outputs(6901) <= not b;
    layer8_outputs(6902) <= a;
    layer8_outputs(6903) <= b;
    layer8_outputs(6904) <= a and b;
    layer8_outputs(6905) <= a or b;
    layer8_outputs(6906) <= b;
    layer8_outputs(6907) <= not a;
    layer8_outputs(6908) <= not (a xor b);
    layer8_outputs(6909) <= not a;
    layer8_outputs(6910) <= a;
    layer8_outputs(6911) <= a;
    layer8_outputs(6912) <= not (a xor b);
    layer8_outputs(6913) <= not (a xor b);
    layer8_outputs(6914) <= a;
    layer8_outputs(6915) <= not (a xor b);
    layer8_outputs(6916) <= b and not a;
    layer8_outputs(6917) <= a xor b;
    layer8_outputs(6918) <= not a;
    layer8_outputs(6919) <= b;
    layer8_outputs(6920) <= not b;
    layer8_outputs(6921) <= not (a and b);
    layer8_outputs(6922) <= not b;
    layer8_outputs(6923) <= a xor b;
    layer8_outputs(6924) <= not (a xor b);
    layer8_outputs(6925) <= a and not b;
    layer8_outputs(6926) <= not b;
    layer8_outputs(6927) <= a and not b;
    layer8_outputs(6928) <= b;
    layer8_outputs(6929) <= not b;
    layer8_outputs(6930) <= a and b;
    layer8_outputs(6931) <= not (a xor b);
    layer8_outputs(6932) <= not b or a;
    layer8_outputs(6933) <= a or b;
    layer8_outputs(6934) <= not a;
    layer8_outputs(6935) <= not (a xor b);
    layer8_outputs(6936) <= a;
    layer8_outputs(6937) <= a or b;
    layer8_outputs(6938) <= not (a or b);
    layer8_outputs(6939) <= not b;
    layer8_outputs(6940) <= b;
    layer8_outputs(6941) <= not (a xor b);
    layer8_outputs(6942) <= not a;
    layer8_outputs(6943) <= not b;
    layer8_outputs(6944) <= a or b;
    layer8_outputs(6945) <= a or b;
    layer8_outputs(6946) <= not b;
    layer8_outputs(6947) <= a and b;
    layer8_outputs(6948) <= not (a xor b);
    layer8_outputs(6949) <= not (a xor b);
    layer8_outputs(6950) <= not b;
    layer8_outputs(6951) <= a;
    layer8_outputs(6952) <= not a or b;
    layer8_outputs(6953) <= a and not b;
    layer8_outputs(6954) <= a or b;
    layer8_outputs(6955) <= a;
    layer8_outputs(6956) <= not a;
    layer8_outputs(6957) <= b;
    layer8_outputs(6958) <= b;
    layer8_outputs(6959) <= not a;
    layer8_outputs(6960) <= a;
    layer8_outputs(6961) <= not a or b;
    layer8_outputs(6962) <= not (a xor b);
    layer8_outputs(6963) <= not b;
    layer8_outputs(6964) <= '1';
    layer8_outputs(6965) <= not a;
    layer8_outputs(6966) <= a;
    layer8_outputs(6967) <= a;
    layer8_outputs(6968) <= a or b;
    layer8_outputs(6969) <= a xor b;
    layer8_outputs(6970) <= a;
    layer8_outputs(6971) <= not a or b;
    layer8_outputs(6972) <= not b or a;
    layer8_outputs(6973) <= not a;
    layer8_outputs(6974) <= not a or b;
    layer8_outputs(6975) <= b;
    layer8_outputs(6976) <= not a or b;
    layer8_outputs(6977) <= not a or b;
    layer8_outputs(6978) <= a and b;
    layer8_outputs(6979) <= not (a and b);
    layer8_outputs(6980) <= b;
    layer8_outputs(6981) <= b and not a;
    layer8_outputs(6982) <= not b;
    layer8_outputs(6983) <= not a;
    layer8_outputs(6984) <= a or b;
    layer8_outputs(6985) <= a xor b;
    layer8_outputs(6986) <= not (a xor b);
    layer8_outputs(6987) <= b;
    layer8_outputs(6988) <= not b;
    layer8_outputs(6989) <= not b;
    layer8_outputs(6990) <= not (a xor b);
    layer8_outputs(6991) <= a and b;
    layer8_outputs(6992) <= a xor b;
    layer8_outputs(6993) <= not a;
    layer8_outputs(6994) <= a and b;
    layer8_outputs(6995) <= a and b;
    layer8_outputs(6996) <= not a;
    layer8_outputs(6997) <= a and not b;
    layer8_outputs(6998) <= a and not b;
    layer8_outputs(6999) <= a and b;
    layer8_outputs(7000) <= not (a and b);
    layer8_outputs(7001) <= a and b;
    layer8_outputs(7002) <= a and not b;
    layer8_outputs(7003) <= a;
    layer8_outputs(7004) <= not a;
    layer8_outputs(7005) <= not b;
    layer8_outputs(7006) <= a or b;
    layer8_outputs(7007) <= a;
    layer8_outputs(7008) <= a xor b;
    layer8_outputs(7009) <= not a;
    layer8_outputs(7010) <= not a or b;
    layer8_outputs(7011) <= a or b;
    layer8_outputs(7012) <= not a;
    layer8_outputs(7013) <= not a;
    layer8_outputs(7014) <= a and not b;
    layer8_outputs(7015) <= not (a and b);
    layer8_outputs(7016) <= not a;
    layer8_outputs(7017) <= a xor b;
    layer8_outputs(7018) <= b;
    layer8_outputs(7019) <= a;
    layer8_outputs(7020) <= b;
    layer8_outputs(7021) <= not a;
    layer8_outputs(7022) <= not a;
    layer8_outputs(7023) <= not (a or b);
    layer8_outputs(7024) <= a and b;
    layer8_outputs(7025) <= not b;
    layer8_outputs(7026) <= not (a xor b);
    layer8_outputs(7027) <= a and not b;
    layer8_outputs(7028) <= not (a xor b);
    layer8_outputs(7029) <= not b or a;
    layer8_outputs(7030) <= a;
    layer8_outputs(7031) <= a;
    layer8_outputs(7032) <= a;
    layer8_outputs(7033) <= a xor b;
    layer8_outputs(7034) <= a or b;
    layer8_outputs(7035) <= not (a and b);
    layer8_outputs(7036) <= not (a xor b);
    layer8_outputs(7037) <= a;
    layer8_outputs(7038) <= a;
    layer8_outputs(7039) <= b and not a;
    layer8_outputs(7040) <= not (a xor b);
    layer8_outputs(7041) <= not b;
    layer8_outputs(7042) <= a and not b;
    layer8_outputs(7043) <= not (a xor b);
    layer8_outputs(7044) <= a xor b;
    layer8_outputs(7045) <= a xor b;
    layer8_outputs(7046) <= not (a xor b);
    layer8_outputs(7047) <= not (a and b);
    layer8_outputs(7048) <= b;
    layer8_outputs(7049) <= not (a xor b);
    layer8_outputs(7050) <= a and not b;
    layer8_outputs(7051) <= a xor b;
    layer8_outputs(7052) <= not a or b;
    layer8_outputs(7053) <= not a or b;
    layer8_outputs(7054) <= not (a or b);
    layer8_outputs(7055) <= not (a and b);
    layer8_outputs(7056) <= not b or a;
    layer8_outputs(7057) <= b;
    layer8_outputs(7058) <= b and not a;
    layer8_outputs(7059) <= not a or b;
    layer8_outputs(7060) <= not (a xor b);
    layer8_outputs(7061) <= a and not b;
    layer8_outputs(7062) <= not b;
    layer8_outputs(7063) <= not (a xor b);
    layer8_outputs(7064) <= a;
    layer8_outputs(7065) <= a xor b;
    layer8_outputs(7066) <= b;
    layer8_outputs(7067) <= '1';
    layer8_outputs(7068) <= a and b;
    layer8_outputs(7069) <= not b;
    layer8_outputs(7070) <= a xor b;
    layer8_outputs(7071) <= a or b;
    layer8_outputs(7072) <= a or b;
    layer8_outputs(7073) <= not a;
    layer8_outputs(7074) <= not b;
    layer8_outputs(7075) <= '1';
    layer8_outputs(7076) <= not b;
    layer8_outputs(7077) <= b;
    layer8_outputs(7078) <= b;
    layer8_outputs(7079) <= not a;
    layer8_outputs(7080) <= b;
    layer8_outputs(7081) <= a;
    layer8_outputs(7082) <= not a;
    layer8_outputs(7083) <= not b;
    layer8_outputs(7084) <= a;
    layer8_outputs(7085) <= b and not a;
    layer8_outputs(7086) <= a;
    layer8_outputs(7087) <= not (a xor b);
    layer8_outputs(7088) <= b and not a;
    layer8_outputs(7089) <= a and b;
    layer8_outputs(7090) <= not b;
    layer8_outputs(7091) <= not b or a;
    layer8_outputs(7092) <= a and not b;
    layer8_outputs(7093) <= not b;
    layer8_outputs(7094) <= not a;
    layer8_outputs(7095) <= not (a xor b);
    layer8_outputs(7096) <= not b or a;
    layer8_outputs(7097) <= b and not a;
    layer8_outputs(7098) <= not b or a;
    layer8_outputs(7099) <= not (a xor b);
    layer8_outputs(7100) <= b;
    layer8_outputs(7101) <= b;
    layer8_outputs(7102) <= a or b;
    layer8_outputs(7103) <= a;
    layer8_outputs(7104) <= not a;
    layer8_outputs(7105) <= b and not a;
    layer8_outputs(7106) <= not (a and b);
    layer8_outputs(7107) <= b;
    layer8_outputs(7108) <= b and not a;
    layer8_outputs(7109) <= b;
    layer8_outputs(7110) <= a and not b;
    layer8_outputs(7111) <= not (a xor b);
    layer8_outputs(7112) <= not b;
    layer8_outputs(7113) <= not (a xor b);
    layer8_outputs(7114) <= a;
    layer8_outputs(7115) <= not a or b;
    layer8_outputs(7116) <= not (a xor b);
    layer8_outputs(7117) <= a xor b;
    layer8_outputs(7118) <= not (a xor b);
    layer8_outputs(7119) <= not b;
    layer8_outputs(7120) <= not a;
    layer8_outputs(7121) <= a xor b;
    layer8_outputs(7122) <= a;
    layer8_outputs(7123) <= a and b;
    layer8_outputs(7124) <= a and b;
    layer8_outputs(7125) <= a xor b;
    layer8_outputs(7126) <= not b;
    layer8_outputs(7127) <= not (a xor b);
    layer8_outputs(7128) <= b;
    layer8_outputs(7129) <= not a;
    layer8_outputs(7130) <= not (a xor b);
    layer8_outputs(7131) <= not (a and b);
    layer8_outputs(7132) <= a and not b;
    layer8_outputs(7133) <= b;
    layer8_outputs(7134) <= a;
    layer8_outputs(7135) <= not b;
    layer8_outputs(7136) <= not b or a;
    layer8_outputs(7137) <= not b;
    layer8_outputs(7138) <= a or b;
    layer8_outputs(7139) <= not (a or b);
    layer8_outputs(7140) <= a;
    layer8_outputs(7141) <= not a or b;
    layer8_outputs(7142) <= not a or b;
    layer8_outputs(7143) <= b and not a;
    layer8_outputs(7144) <= a or b;
    layer8_outputs(7145) <= a or b;
    layer8_outputs(7146) <= '0';
    layer8_outputs(7147) <= not a or b;
    layer8_outputs(7148) <= b;
    layer8_outputs(7149) <= not (a or b);
    layer8_outputs(7150) <= a or b;
    layer8_outputs(7151) <= b;
    layer8_outputs(7152) <= a;
    layer8_outputs(7153) <= a;
    layer8_outputs(7154) <= not b or a;
    layer8_outputs(7155) <= not b;
    layer8_outputs(7156) <= a and not b;
    layer8_outputs(7157) <= not a or b;
    layer8_outputs(7158) <= a xor b;
    layer8_outputs(7159) <= not (a and b);
    layer8_outputs(7160) <= a or b;
    layer8_outputs(7161) <= not a;
    layer8_outputs(7162) <= not b or a;
    layer8_outputs(7163) <= not a or b;
    layer8_outputs(7164) <= a xor b;
    layer8_outputs(7165) <= a xor b;
    layer8_outputs(7166) <= not b;
    layer8_outputs(7167) <= a xor b;
    layer8_outputs(7168) <= not b;
    layer8_outputs(7169) <= not (a or b);
    layer8_outputs(7170) <= not b or a;
    layer8_outputs(7171) <= not a;
    layer8_outputs(7172) <= a and b;
    layer8_outputs(7173) <= a and not b;
    layer8_outputs(7174) <= not (a or b);
    layer8_outputs(7175) <= not b or a;
    layer8_outputs(7176) <= not (a xor b);
    layer8_outputs(7177) <= not (a or b);
    layer8_outputs(7178) <= not (a xor b);
    layer8_outputs(7179) <= not b;
    layer8_outputs(7180) <= a or b;
    layer8_outputs(7181) <= a and not b;
    layer8_outputs(7182) <= not a;
    layer8_outputs(7183) <= not a;
    layer8_outputs(7184) <= not (a and b);
    layer8_outputs(7185) <= b and not a;
    layer8_outputs(7186) <= b;
    layer8_outputs(7187) <= a xor b;
    layer8_outputs(7188) <= not (a and b);
    layer8_outputs(7189) <= not b or a;
    layer8_outputs(7190) <= b;
    layer8_outputs(7191) <= not (a and b);
    layer8_outputs(7192) <= not a or b;
    layer8_outputs(7193) <= not (a xor b);
    layer8_outputs(7194) <= not a;
    layer8_outputs(7195) <= a and b;
    layer8_outputs(7196) <= b;
    layer8_outputs(7197) <= '0';
    layer8_outputs(7198) <= not b;
    layer8_outputs(7199) <= a;
    layer8_outputs(7200) <= not a or b;
    layer8_outputs(7201) <= not a;
    layer8_outputs(7202) <= a and b;
    layer8_outputs(7203) <= a and b;
    layer8_outputs(7204) <= not a;
    layer8_outputs(7205) <= a;
    layer8_outputs(7206) <= a xor b;
    layer8_outputs(7207) <= not (a and b);
    layer8_outputs(7208) <= a xor b;
    layer8_outputs(7209) <= a and not b;
    layer8_outputs(7210) <= a;
    layer8_outputs(7211) <= b;
    layer8_outputs(7212) <= not a;
    layer8_outputs(7213) <= a xor b;
    layer8_outputs(7214) <= not b;
    layer8_outputs(7215) <= a;
    layer8_outputs(7216) <= a xor b;
    layer8_outputs(7217) <= not (a xor b);
    layer8_outputs(7218) <= a xor b;
    layer8_outputs(7219) <= b;
    layer8_outputs(7220) <= b;
    layer8_outputs(7221) <= a;
    layer8_outputs(7222) <= b and not a;
    layer8_outputs(7223) <= a or b;
    layer8_outputs(7224) <= not b;
    layer8_outputs(7225) <= b;
    layer8_outputs(7226) <= not (a and b);
    layer8_outputs(7227) <= a;
    layer8_outputs(7228) <= not b;
    layer8_outputs(7229) <= not (a xor b);
    layer8_outputs(7230) <= not (a xor b);
    layer8_outputs(7231) <= a xor b;
    layer8_outputs(7232) <= not (a and b);
    layer8_outputs(7233) <= not a;
    layer8_outputs(7234) <= not (a and b);
    layer8_outputs(7235) <= not a;
    layer8_outputs(7236) <= a xor b;
    layer8_outputs(7237) <= a or b;
    layer8_outputs(7238) <= not a;
    layer8_outputs(7239) <= b;
    layer8_outputs(7240) <= not a or b;
    layer8_outputs(7241) <= not (a and b);
    layer8_outputs(7242) <= not a;
    layer8_outputs(7243) <= '0';
    layer8_outputs(7244) <= not (a xor b);
    layer8_outputs(7245) <= a or b;
    layer8_outputs(7246) <= not b or a;
    layer8_outputs(7247) <= not (a xor b);
    layer8_outputs(7248) <= not (a xor b);
    layer8_outputs(7249) <= not b or a;
    layer8_outputs(7250) <= not (a and b);
    layer8_outputs(7251) <= not (a or b);
    layer8_outputs(7252) <= not (a or b);
    layer8_outputs(7253) <= not a;
    layer8_outputs(7254) <= not a;
    layer8_outputs(7255) <= not a;
    layer8_outputs(7256) <= a;
    layer8_outputs(7257) <= a and b;
    layer8_outputs(7258) <= a and b;
    layer8_outputs(7259) <= not (a or b);
    layer8_outputs(7260) <= a xor b;
    layer8_outputs(7261) <= b;
    layer8_outputs(7262) <= a xor b;
    layer8_outputs(7263) <= not a;
    layer8_outputs(7264) <= not a;
    layer8_outputs(7265) <= b;
    layer8_outputs(7266) <= not (a and b);
    layer8_outputs(7267) <= not a;
    layer8_outputs(7268) <= a and b;
    layer8_outputs(7269) <= not (a xor b);
    layer8_outputs(7270) <= not (a xor b);
    layer8_outputs(7271) <= not a;
    layer8_outputs(7272) <= not a;
    layer8_outputs(7273) <= a xor b;
    layer8_outputs(7274) <= a or b;
    layer8_outputs(7275) <= a and not b;
    layer8_outputs(7276) <= not a or b;
    layer8_outputs(7277) <= a;
    layer8_outputs(7278) <= not b;
    layer8_outputs(7279) <= not a or b;
    layer8_outputs(7280) <= not b or a;
    layer8_outputs(7281) <= not (a or b);
    layer8_outputs(7282) <= not a;
    layer8_outputs(7283) <= not (a or b);
    layer8_outputs(7284) <= not a;
    layer8_outputs(7285) <= not b;
    layer8_outputs(7286) <= a;
    layer8_outputs(7287) <= not (a or b);
    layer8_outputs(7288) <= not a;
    layer8_outputs(7289) <= not b;
    layer8_outputs(7290) <= not (a xor b);
    layer8_outputs(7291) <= not (a xor b);
    layer8_outputs(7292) <= b;
    layer8_outputs(7293) <= a xor b;
    layer8_outputs(7294) <= not b or a;
    layer8_outputs(7295) <= not (a or b);
    layer8_outputs(7296) <= not (a and b);
    layer8_outputs(7297) <= not (a xor b);
    layer8_outputs(7298) <= a xor b;
    layer8_outputs(7299) <= not (a or b);
    layer8_outputs(7300) <= not b or a;
    layer8_outputs(7301) <= not b;
    layer8_outputs(7302) <= not (a xor b);
    layer8_outputs(7303) <= not a or b;
    layer8_outputs(7304) <= not (a xor b);
    layer8_outputs(7305) <= not b;
    layer8_outputs(7306) <= not a;
    layer8_outputs(7307) <= not (a and b);
    layer8_outputs(7308) <= a xor b;
    layer8_outputs(7309) <= not a;
    layer8_outputs(7310) <= a and not b;
    layer8_outputs(7311) <= not a;
    layer8_outputs(7312) <= not b;
    layer8_outputs(7313) <= not (a or b);
    layer8_outputs(7314) <= not a;
    layer8_outputs(7315) <= not b or a;
    layer8_outputs(7316) <= b;
    layer8_outputs(7317) <= b and not a;
    layer8_outputs(7318) <= not b;
    layer8_outputs(7319) <= not b;
    layer8_outputs(7320) <= not (a or b);
    layer8_outputs(7321) <= a and not b;
    layer8_outputs(7322) <= not a;
    layer8_outputs(7323) <= not a;
    layer8_outputs(7324) <= b;
    layer8_outputs(7325) <= a and b;
    layer8_outputs(7326) <= not (a xor b);
    layer8_outputs(7327) <= a;
    layer8_outputs(7328) <= not b;
    layer8_outputs(7329) <= not b;
    layer8_outputs(7330) <= not (a or b);
    layer8_outputs(7331) <= not b;
    layer8_outputs(7332) <= a or b;
    layer8_outputs(7333) <= not a or b;
    layer8_outputs(7334) <= not b or a;
    layer8_outputs(7335) <= a and not b;
    layer8_outputs(7336) <= a and b;
    layer8_outputs(7337) <= not a or b;
    layer8_outputs(7338) <= '1';
    layer8_outputs(7339) <= not a;
    layer8_outputs(7340) <= not b;
    layer8_outputs(7341) <= a xor b;
    layer8_outputs(7342) <= b;
    layer8_outputs(7343) <= not (a and b);
    layer8_outputs(7344) <= not b;
    layer8_outputs(7345) <= not (a xor b);
    layer8_outputs(7346) <= a and not b;
    layer8_outputs(7347) <= b;
    layer8_outputs(7348) <= b;
    layer8_outputs(7349) <= a;
    layer8_outputs(7350) <= not (a xor b);
    layer8_outputs(7351) <= not b;
    layer8_outputs(7352) <= not (a xor b);
    layer8_outputs(7353) <= a;
    layer8_outputs(7354) <= not b;
    layer8_outputs(7355) <= a xor b;
    layer8_outputs(7356) <= a xor b;
    layer8_outputs(7357) <= not a or b;
    layer8_outputs(7358) <= not b;
    layer8_outputs(7359) <= not a or b;
    layer8_outputs(7360) <= not (a xor b);
    layer8_outputs(7361) <= not b;
    layer8_outputs(7362) <= not b or a;
    layer8_outputs(7363) <= not (a or b);
    layer8_outputs(7364) <= a;
    layer8_outputs(7365) <= a xor b;
    layer8_outputs(7366) <= b;
    layer8_outputs(7367) <= not a or b;
    layer8_outputs(7368) <= b;
    layer8_outputs(7369) <= not b or a;
    layer8_outputs(7370) <= not (a xor b);
    layer8_outputs(7371) <= b;
    layer8_outputs(7372) <= not a or b;
    layer8_outputs(7373) <= not b;
    layer8_outputs(7374) <= not (a xor b);
    layer8_outputs(7375) <= b;
    layer8_outputs(7376) <= not (a and b);
    layer8_outputs(7377) <= not (a xor b);
    layer8_outputs(7378) <= b;
    layer8_outputs(7379) <= not a;
    layer8_outputs(7380) <= b;
    layer8_outputs(7381) <= not b or a;
    layer8_outputs(7382) <= a;
    layer8_outputs(7383) <= a or b;
    layer8_outputs(7384) <= not (a xor b);
    layer8_outputs(7385) <= not b or a;
    layer8_outputs(7386) <= b;
    layer8_outputs(7387) <= a or b;
    layer8_outputs(7388) <= a or b;
    layer8_outputs(7389) <= a or b;
    layer8_outputs(7390) <= '0';
    layer8_outputs(7391) <= a and not b;
    layer8_outputs(7392) <= not a or b;
    layer8_outputs(7393) <= not a;
    layer8_outputs(7394) <= b;
    layer8_outputs(7395) <= '0';
    layer8_outputs(7396) <= not b;
    layer8_outputs(7397) <= b and not a;
    layer8_outputs(7398) <= b;
    layer8_outputs(7399) <= not (a xor b);
    layer8_outputs(7400) <= a and b;
    layer8_outputs(7401) <= b and not a;
    layer8_outputs(7402) <= b and not a;
    layer8_outputs(7403) <= not a;
    layer8_outputs(7404) <= a and not b;
    layer8_outputs(7405) <= a and b;
    layer8_outputs(7406) <= b and not a;
    layer8_outputs(7407) <= b;
    layer8_outputs(7408) <= not a;
    layer8_outputs(7409) <= b and not a;
    layer8_outputs(7410) <= not b;
    layer8_outputs(7411) <= not b;
    layer8_outputs(7412) <= not (a xor b);
    layer8_outputs(7413) <= not b or a;
    layer8_outputs(7414) <= b;
    layer8_outputs(7415) <= not b or a;
    layer8_outputs(7416) <= not a;
    layer8_outputs(7417) <= not (a and b);
    layer8_outputs(7418) <= a xor b;
    layer8_outputs(7419) <= a;
    layer8_outputs(7420) <= a or b;
    layer8_outputs(7421) <= not a;
    layer8_outputs(7422) <= b;
    layer8_outputs(7423) <= not a;
    layer8_outputs(7424) <= not b;
    layer8_outputs(7425) <= not b;
    layer8_outputs(7426) <= a and not b;
    layer8_outputs(7427) <= not (a xor b);
    layer8_outputs(7428) <= not b;
    layer8_outputs(7429) <= not b;
    layer8_outputs(7430) <= not b;
    layer8_outputs(7431) <= a;
    layer8_outputs(7432) <= not (a xor b);
    layer8_outputs(7433) <= a xor b;
    layer8_outputs(7434) <= not (a xor b);
    layer8_outputs(7435) <= not b;
    layer8_outputs(7436) <= b;
    layer8_outputs(7437) <= b;
    layer8_outputs(7438) <= not (a xor b);
    layer8_outputs(7439) <= a and not b;
    layer8_outputs(7440) <= a xor b;
    layer8_outputs(7441) <= a xor b;
    layer8_outputs(7442) <= b;
    layer8_outputs(7443) <= a and b;
    layer8_outputs(7444) <= a;
    layer8_outputs(7445) <= not (a and b);
    layer8_outputs(7446) <= not b;
    layer8_outputs(7447) <= b;
    layer8_outputs(7448) <= a and not b;
    layer8_outputs(7449) <= not (a xor b);
    layer8_outputs(7450) <= not b or a;
    layer8_outputs(7451) <= a;
    layer8_outputs(7452) <= b;
    layer8_outputs(7453) <= not b;
    layer8_outputs(7454) <= b;
    layer8_outputs(7455) <= not a;
    layer8_outputs(7456) <= b;
    layer8_outputs(7457) <= not (a and b);
    layer8_outputs(7458) <= b and not a;
    layer8_outputs(7459) <= a;
    layer8_outputs(7460) <= a;
    layer8_outputs(7461) <= a;
    layer8_outputs(7462) <= not (a and b);
    layer8_outputs(7463) <= a xor b;
    layer8_outputs(7464) <= a or b;
    layer8_outputs(7465) <= a;
    layer8_outputs(7466) <= not a;
    layer8_outputs(7467) <= '1';
    layer8_outputs(7468) <= b and not a;
    layer8_outputs(7469) <= a and not b;
    layer8_outputs(7470) <= not (a or b);
    layer8_outputs(7471) <= not a;
    layer8_outputs(7472) <= a and b;
    layer8_outputs(7473) <= a xor b;
    layer8_outputs(7474) <= a and not b;
    layer8_outputs(7475) <= a or b;
    layer8_outputs(7476) <= not (a xor b);
    layer8_outputs(7477) <= not a or b;
    layer8_outputs(7478) <= not (a xor b);
    layer8_outputs(7479) <= not b;
    layer8_outputs(7480) <= not a;
    layer8_outputs(7481) <= not b or a;
    layer8_outputs(7482) <= not (a and b);
    layer8_outputs(7483) <= not a;
    layer8_outputs(7484) <= not a;
    layer8_outputs(7485) <= a xor b;
    layer8_outputs(7486) <= not (a or b);
    layer8_outputs(7487) <= not b or a;
    layer8_outputs(7488) <= not a or b;
    layer8_outputs(7489) <= not (a and b);
    layer8_outputs(7490) <= a;
    layer8_outputs(7491) <= not a;
    layer8_outputs(7492) <= not a;
    layer8_outputs(7493) <= not a;
    layer8_outputs(7494) <= a or b;
    layer8_outputs(7495) <= a xor b;
    layer8_outputs(7496) <= a xor b;
    layer8_outputs(7497) <= not a;
    layer8_outputs(7498) <= not b or a;
    layer8_outputs(7499) <= b;
    layer8_outputs(7500) <= not a;
    layer8_outputs(7501) <= not a;
    layer8_outputs(7502) <= not (a xor b);
    layer8_outputs(7503) <= not a or b;
    layer8_outputs(7504) <= not b;
    layer8_outputs(7505) <= not (a xor b);
    layer8_outputs(7506) <= not (a xor b);
    layer8_outputs(7507) <= a;
    layer8_outputs(7508) <= not a;
    layer8_outputs(7509) <= a;
    layer8_outputs(7510) <= not (a xor b);
    layer8_outputs(7511) <= b and not a;
    layer8_outputs(7512) <= not (a xor b);
    layer8_outputs(7513) <= b;
    layer8_outputs(7514) <= not b or a;
    layer8_outputs(7515) <= not a or b;
    layer8_outputs(7516) <= not (a xor b);
    layer8_outputs(7517) <= not (a xor b);
    layer8_outputs(7518) <= not a or b;
    layer8_outputs(7519) <= a or b;
    layer8_outputs(7520) <= a;
    layer8_outputs(7521) <= not a or b;
    layer8_outputs(7522) <= not b or a;
    layer8_outputs(7523) <= not b;
    layer8_outputs(7524) <= a xor b;
    layer8_outputs(7525) <= b;
    layer8_outputs(7526) <= not b or a;
    layer8_outputs(7527) <= b;
    layer8_outputs(7528) <= not (a or b);
    layer8_outputs(7529) <= a and b;
    layer8_outputs(7530) <= not a;
    layer8_outputs(7531) <= not b;
    layer8_outputs(7532) <= a xor b;
    layer8_outputs(7533) <= not (a or b);
    layer8_outputs(7534) <= a;
    layer8_outputs(7535) <= not (a xor b);
    layer8_outputs(7536) <= a xor b;
    layer8_outputs(7537) <= a xor b;
    layer8_outputs(7538) <= not a or b;
    layer8_outputs(7539) <= not a;
    layer8_outputs(7540) <= not a;
    layer8_outputs(7541) <= a or b;
    layer8_outputs(7542) <= not a;
    layer8_outputs(7543) <= not a;
    layer8_outputs(7544) <= not a;
    layer8_outputs(7545) <= not (a xor b);
    layer8_outputs(7546) <= b;
    layer8_outputs(7547) <= not (a and b);
    layer8_outputs(7548) <= not b;
    layer8_outputs(7549) <= not (a xor b);
    layer8_outputs(7550) <= not a or b;
    layer8_outputs(7551) <= not b;
    layer8_outputs(7552) <= a or b;
    layer8_outputs(7553) <= not a;
    layer8_outputs(7554) <= a;
    layer8_outputs(7555) <= not (a and b);
    layer8_outputs(7556) <= b;
    layer8_outputs(7557) <= not a;
    layer8_outputs(7558) <= a;
    layer8_outputs(7559) <= a or b;
    layer8_outputs(7560) <= not a;
    layer8_outputs(7561) <= not (a xor b);
    layer8_outputs(7562) <= not (a and b);
    layer8_outputs(7563) <= a;
    layer8_outputs(7564) <= a xor b;
    layer8_outputs(7565) <= not a or b;
    layer8_outputs(7566) <= b;
    layer8_outputs(7567) <= b;
    layer8_outputs(7568) <= a xor b;
    layer8_outputs(7569) <= not b;
    layer8_outputs(7570) <= not (a xor b);
    layer8_outputs(7571) <= not b or a;
    layer8_outputs(7572) <= '1';
    layer8_outputs(7573) <= a and not b;
    layer8_outputs(7574) <= not (a xor b);
    layer8_outputs(7575) <= not (a xor b);
    layer8_outputs(7576) <= not a or b;
    layer8_outputs(7577) <= b;
    layer8_outputs(7578) <= not (a and b);
    layer8_outputs(7579) <= not a;
    layer8_outputs(7580) <= not b;
    layer8_outputs(7581) <= a xor b;
    layer8_outputs(7582) <= a and not b;
    layer8_outputs(7583) <= a and not b;
    layer8_outputs(7584) <= not a;
    layer8_outputs(7585) <= a xor b;
    layer8_outputs(7586) <= not b;
    layer8_outputs(7587) <= '0';
    layer8_outputs(7588) <= a xor b;
    layer8_outputs(7589) <= '0';
    layer8_outputs(7590) <= a and not b;
    layer8_outputs(7591) <= not (a xor b);
    layer8_outputs(7592) <= not a;
    layer8_outputs(7593) <= b and not a;
    layer8_outputs(7594) <= b;
    layer8_outputs(7595) <= not a;
    layer8_outputs(7596) <= not b;
    layer8_outputs(7597) <= not b;
    layer8_outputs(7598) <= a and b;
    layer8_outputs(7599) <= not a or b;
    layer8_outputs(7600) <= a xor b;
    layer8_outputs(7601) <= not b;
    layer8_outputs(7602) <= not b;
    layer8_outputs(7603) <= not (a xor b);
    layer8_outputs(7604) <= not (a xor b);
    layer8_outputs(7605) <= a;
    layer8_outputs(7606) <= not (a or b);
    layer8_outputs(7607) <= not b or a;
    layer8_outputs(7608) <= b;
    layer8_outputs(7609) <= not a or b;
    layer8_outputs(7610) <= not a or b;
    layer8_outputs(7611) <= not b;
    layer8_outputs(7612) <= b;
    layer8_outputs(7613) <= not a;
    layer8_outputs(7614) <= not (a and b);
    layer8_outputs(7615) <= '1';
    layer8_outputs(7616) <= a and b;
    layer8_outputs(7617) <= not b or a;
    layer8_outputs(7618) <= not b;
    layer8_outputs(7619) <= not b or a;
    layer8_outputs(7620) <= not (a and b);
    layer8_outputs(7621) <= a;
    layer8_outputs(7622) <= not a;
    layer8_outputs(7623) <= a and not b;
    layer8_outputs(7624) <= b;
    layer8_outputs(7625) <= b and not a;
    layer8_outputs(7626) <= '1';
    layer8_outputs(7627) <= not a;
    layer8_outputs(7628) <= a xor b;
    layer8_outputs(7629) <= a;
    layer8_outputs(7630) <= not (a or b);
    layer8_outputs(7631) <= not (a or b);
    layer8_outputs(7632) <= b and not a;
    layer8_outputs(7633) <= not a;
    layer8_outputs(7634) <= a;
    layer8_outputs(7635) <= a xor b;
    layer8_outputs(7636) <= a xor b;
    layer8_outputs(7637) <= not b;
    layer8_outputs(7638) <= not a;
    layer8_outputs(7639) <= a;
    layer8_outputs(7640) <= b;
    layer8_outputs(7641) <= not (a xor b);
    layer8_outputs(7642) <= not b or a;
    layer8_outputs(7643) <= not (a or b);
    layer8_outputs(7644) <= a xor b;
    layer8_outputs(7645) <= not (a xor b);
    layer8_outputs(7646) <= not b or a;
    layer8_outputs(7647) <= not a;
    layer8_outputs(7648) <= not b;
    layer8_outputs(7649) <= b;
    layer8_outputs(7650) <= a and not b;
    layer8_outputs(7651) <= not (a xor b);
    layer8_outputs(7652) <= not a or b;
    layer8_outputs(7653) <= b and not a;
    layer8_outputs(7654) <= a or b;
    layer8_outputs(7655) <= not (a and b);
    layer8_outputs(7656) <= a or b;
    layer8_outputs(7657) <= a and not b;
    layer8_outputs(7658) <= not b;
    layer8_outputs(7659) <= a xor b;
    layer8_outputs(7660) <= a and not b;
    layer8_outputs(7661) <= not b;
    layer8_outputs(7662) <= b;
    layer8_outputs(7663) <= not (a xor b);
    layer8_outputs(7664) <= not (a and b);
    layer8_outputs(7665) <= not a;
    layer8_outputs(7666) <= a and not b;
    layer8_outputs(7667) <= a;
    layer8_outputs(7668) <= b and not a;
    layer8_outputs(7669) <= not a;
    layer8_outputs(7670) <= not b;
    layer8_outputs(7671) <= a and b;
    layer8_outputs(7672) <= a or b;
    layer8_outputs(7673) <= b;
    layer8_outputs(7674) <= a;
    layer8_outputs(7675) <= a;
    layer8_outputs(7676) <= not b;
    layer8_outputs(7677) <= not a;
    layer8_outputs(7678) <= not (a or b);
    layer8_outputs(7679) <= b;
    outputs(0) <= b;
    outputs(1) <= a xor b;
    outputs(2) <= not b;
    outputs(3) <= b;
    outputs(4) <= a xor b;
    outputs(5) <= not (a xor b);
    outputs(6) <= not (a xor b);
    outputs(7) <= a xor b;
    outputs(8) <= a;
    outputs(9) <= a xor b;
    outputs(10) <= not a;
    outputs(11) <= b;
    outputs(12) <= b;
    outputs(13) <= not b;
    outputs(14) <= not (a xor b);
    outputs(15) <= b and not a;
    outputs(16) <= a and b;
    outputs(17) <= not (a or b);
    outputs(18) <= b;
    outputs(19) <= a;
    outputs(20) <= a;
    outputs(21) <= a xor b;
    outputs(22) <= not a;
    outputs(23) <= a xor b;
    outputs(24) <= a and b;
    outputs(25) <= b and not a;
    outputs(26) <= a;
    outputs(27) <= a xor b;
    outputs(28) <= b and not a;
    outputs(29) <= not a;
    outputs(30) <= a;
    outputs(31) <= not (a xor b);
    outputs(32) <= a xor b;
    outputs(33) <= a;
    outputs(34) <= not (a or b);
    outputs(35) <= not a;
    outputs(36) <= not (a xor b);
    outputs(37) <= a xor b;
    outputs(38) <= not (a xor b);
    outputs(39) <= b;
    outputs(40) <= b;
    outputs(41) <= a;
    outputs(42) <= not (a or b);
    outputs(43) <= b;
    outputs(44) <= b;
    outputs(45) <= not (a xor b);
    outputs(46) <= b;
    outputs(47) <= a xor b;
    outputs(48) <= not b;
    outputs(49) <= b;
    outputs(50) <= not b;
    outputs(51) <= a and b;
    outputs(52) <= a and b;
    outputs(53) <= not (a xor b);
    outputs(54) <= not (a xor b);
    outputs(55) <= a xor b;
    outputs(56) <= not (a and b);
    outputs(57) <= not (a xor b);
    outputs(58) <= not b or a;
    outputs(59) <= not (a xor b);
    outputs(60) <= a xor b;
    outputs(61) <= not a;
    outputs(62) <= not (a or b);
    outputs(63) <= b;
    outputs(64) <= not b;
    outputs(65) <= a;
    outputs(66) <= a;
    outputs(67) <= not (a or b);
    outputs(68) <= not b;
    outputs(69) <= not a or b;
    outputs(70) <= not b;
    outputs(71) <= a and not b;
    outputs(72) <= not (a or b);
    outputs(73) <= not b or a;
    outputs(74) <= not (a xor b);
    outputs(75) <= b;
    outputs(76) <= a and b;
    outputs(77) <= not b;
    outputs(78) <= a;
    outputs(79) <= a xor b;
    outputs(80) <= a and not b;
    outputs(81) <= a;
    outputs(82) <= not a;
    outputs(83) <= a xor b;
    outputs(84) <= b;
    outputs(85) <= a and b;
    outputs(86) <= not (a or b);
    outputs(87) <= a xor b;
    outputs(88) <= not (a or b);
    outputs(89) <= not a;
    outputs(90) <= a;
    outputs(91) <= not b;
    outputs(92) <= a and b;
    outputs(93) <= a;
    outputs(94) <= a xor b;
    outputs(95) <= a;
    outputs(96) <= b;
    outputs(97) <= a and b;
    outputs(98) <= not a;
    outputs(99) <= not (a xor b);
    outputs(100) <= not b or a;
    outputs(101) <= b;
    outputs(102) <= a and not b;
    outputs(103) <= b;
    outputs(104) <= not a;
    outputs(105) <= a and not b;
    outputs(106) <= b;
    outputs(107) <= a xor b;
    outputs(108) <= a xor b;
    outputs(109) <= not b;
    outputs(110) <= not (a or b);
    outputs(111) <= not a or b;
    outputs(112) <= not b;
    outputs(113) <= not (a xor b);
    outputs(114) <= not (a xor b);
    outputs(115) <= a xor b;
    outputs(116) <= not (a xor b);
    outputs(117) <= b and not a;
    outputs(118) <= b and not a;
    outputs(119) <= not a;
    outputs(120) <= b;
    outputs(121) <= a xor b;
    outputs(122) <= not a;
    outputs(123) <= not a;
    outputs(124) <= a;
    outputs(125) <= b and not a;
    outputs(126) <= not (a xor b);
    outputs(127) <= a xor b;
    outputs(128) <= not (a xor b);
    outputs(129) <= a;
    outputs(130) <= a xor b;
    outputs(131) <= a xor b;
    outputs(132) <= b;
    outputs(133) <= not b;
    outputs(134) <= a;
    outputs(135) <= a xor b;
    outputs(136) <= a;
    outputs(137) <= not b;
    outputs(138) <= not (a xor b);
    outputs(139) <= not b;
    outputs(140) <= not a;
    outputs(141) <= not b;
    outputs(142) <= not b;
    outputs(143) <= a and not b;
    outputs(144) <= not b;
    outputs(145) <= a and b;
    outputs(146) <= not a;
    outputs(147) <= b;
    outputs(148) <= a and not b;
    outputs(149) <= not a;
    outputs(150) <= a xor b;
    outputs(151) <= a and b;
    outputs(152) <= a and b;
    outputs(153) <= b;
    outputs(154) <= not (a or b);
    outputs(155) <= b and not a;
    outputs(156) <= a;
    outputs(157) <= not (a and b);
    outputs(158) <= not (a or b);
    outputs(159) <= b;
    outputs(160) <= not a;
    outputs(161) <= not a;
    outputs(162) <= b;
    outputs(163) <= a and not b;
    outputs(164) <= b;
    outputs(165) <= not (a xor b);
    outputs(166) <= not (a or b);
    outputs(167) <= a xor b;
    outputs(168) <= not b;
    outputs(169) <= b;
    outputs(170) <= a;
    outputs(171) <= not b;
    outputs(172) <= a and b;
    outputs(173) <= a and b;
    outputs(174) <= not b or a;
    outputs(175) <= a or b;
    outputs(176) <= not a;
    outputs(177) <= not a;
    outputs(178) <= not (a xor b);
    outputs(179) <= a;
    outputs(180) <= a;
    outputs(181) <= a xor b;
    outputs(182) <= a xor b;
    outputs(183) <= b and not a;
    outputs(184) <= not a;
    outputs(185) <= a and b;
    outputs(186) <= b;
    outputs(187) <= not (a xor b);
    outputs(188) <= b and not a;
    outputs(189) <= a xor b;
    outputs(190) <= a;
    outputs(191) <= not (a xor b);
    outputs(192) <= a and not b;
    outputs(193) <= not (a or b);
    outputs(194) <= b;
    outputs(195) <= b and not a;
    outputs(196) <= a xor b;
    outputs(197) <= not (a or b);
    outputs(198) <= b;
    outputs(199) <= not (a and b);
    outputs(200) <= not (a or b);
    outputs(201) <= b;
    outputs(202) <= a and b;
    outputs(203) <= a;
    outputs(204) <= not a;
    outputs(205) <= not (a or b);
    outputs(206) <= not a;
    outputs(207) <= not (a or b);
    outputs(208) <= not a;
    outputs(209) <= not b;
    outputs(210) <= not b or a;
    outputs(211) <= not a;
    outputs(212) <= b;
    outputs(213) <= not (a or b);
    outputs(214) <= a and b;
    outputs(215) <= not (a or b);
    outputs(216) <= b;
    outputs(217) <= not a;
    outputs(218) <= not b;
    outputs(219) <= a xor b;
    outputs(220) <= a and b;
    outputs(221) <= not a;
    outputs(222) <= not b or a;
    outputs(223) <= a;
    outputs(224) <= a;
    outputs(225) <= a xor b;
    outputs(226) <= not b;
    outputs(227) <= b;
    outputs(228) <= not (a and b);
    outputs(229) <= a;
    outputs(230) <= b;
    outputs(231) <= not a;
    outputs(232) <= b;
    outputs(233) <= a xor b;
    outputs(234) <= a;
    outputs(235) <= a and not b;
    outputs(236) <= b;
    outputs(237) <= not (a xor b);
    outputs(238) <= not (a or b);
    outputs(239) <= not a;
    outputs(240) <= a;
    outputs(241) <= a and b;
    outputs(242) <= a;
    outputs(243) <= not (a or b);
    outputs(244) <= a or b;
    outputs(245) <= a xor b;
    outputs(246) <= not a;
    outputs(247) <= b;
    outputs(248) <= not a;
    outputs(249) <= not a;
    outputs(250) <= a;
    outputs(251) <= a and b;
    outputs(252) <= not (a xor b);
    outputs(253) <= a xor b;
    outputs(254) <= not a;
    outputs(255) <= not b;
    outputs(256) <= not b;
    outputs(257) <= a;
    outputs(258) <= not (a xor b);
    outputs(259) <= not a;
    outputs(260) <= b;
    outputs(261) <= not a;
    outputs(262) <= a;
    outputs(263) <= not (a xor b);
    outputs(264) <= a xor b;
    outputs(265) <= not b;
    outputs(266) <= not (a or b);
    outputs(267) <= a xor b;
    outputs(268) <= a xor b;
    outputs(269) <= a and b;
    outputs(270) <= a xor b;
    outputs(271) <= a xor b;
    outputs(272) <= a;
    outputs(273) <= b and not a;
    outputs(274) <= a and not b;
    outputs(275) <= a or b;
    outputs(276) <= not a;
    outputs(277) <= b;
    outputs(278) <= not (a and b);
    outputs(279) <= not a;
    outputs(280) <= a or b;
    outputs(281) <= not (a xor b);
    outputs(282) <= b and not a;
    outputs(283) <= not (a or b);
    outputs(284) <= a and b;
    outputs(285) <= a;
    outputs(286) <= b;
    outputs(287) <= not b;
    outputs(288) <= a;
    outputs(289) <= b and not a;
    outputs(290) <= not b;
    outputs(291) <= not (a or b);
    outputs(292) <= b;
    outputs(293) <= a and not b;
    outputs(294) <= not b;
    outputs(295) <= b;
    outputs(296) <= b;
    outputs(297) <= not (a and b);
    outputs(298) <= a and b;
    outputs(299) <= b;
    outputs(300) <= not (a or b);
    outputs(301) <= b;
    outputs(302) <= b and not a;
    outputs(303) <= a and b;
    outputs(304) <= not b;
    outputs(305) <= not b;
    outputs(306) <= b;
    outputs(307) <= not b;
    outputs(308) <= a xor b;
    outputs(309) <= not a;
    outputs(310) <= not b;
    outputs(311) <= not (a xor b);
    outputs(312) <= a and b;
    outputs(313) <= not a or b;
    outputs(314) <= not (a or b);
    outputs(315) <= b and not a;
    outputs(316) <= a xor b;
    outputs(317) <= not b;
    outputs(318) <= b;
    outputs(319) <= a xor b;
    outputs(320) <= b;
    outputs(321) <= not (a xor b);
    outputs(322) <= not (a xor b);
    outputs(323) <= not (a or b);
    outputs(324) <= not (a xor b);
    outputs(325) <= a xor b;
    outputs(326) <= not a;
    outputs(327) <= not b;
    outputs(328) <= b;
    outputs(329) <= a;
    outputs(330) <= b;
    outputs(331) <= a xor b;
    outputs(332) <= a and b;
    outputs(333) <= a;
    outputs(334) <= b;
    outputs(335) <= not b;
    outputs(336) <= a or b;
    outputs(337) <= not b or a;
    outputs(338) <= a;
    outputs(339) <= a xor b;
    outputs(340) <= a xor b;
    outputs(341) <= not (a xor b);
    outputs(342) <= not a;
    outputs(343) <= not a;
    outputs(344) <= not a;
    outputs(345) <= a and b;
    outputs(346) <= not (a and b);
    outputs(347) <= not a;
    outputs(348) <= not a;
    outputs(349) <= a;
    outputs(350) <= a xor b;
    outputs(351) <= not (a xor b);
    outputs(352) <= a;
    outputs(353) <= b and not a;
    outputs(354) <= b;
    outputs(355) <= b;
    outputs(356) <= a or b;
    outputs(357) <= not (a xor b);
    outputs(358) <= b and not a;
    outputs(359) <= a;
    outputs(360) <= b and not a;
    outputs(361) <= b and not a;
    outputs(362) <= not b;
    outputs(363) <= not a;
    outputs(364) <= a and b;
    outputs(365) <= a;
    outputs(366) <= not a;
    outputs(367) <= a xor b;
    outputs(368) <= not (a xor b);
    outputs(369) <= not (a xor b);
    outputs(370) <= not b;
    outputs(371) <= a xor b;
    outputs(372) <= not b;
    outputs(373) <= a and b;
    outputs(374) <= a xor b;
    outputs(375) <= a or b;
    outputs(376) <= a and not b;
    outputs(377) <= a;
    outputs(378) <= not (a or b);
    outputs(379) <= not a;
    outputs(380) <= a xor b;
    outputs(381) <= a xor b;
    outputs(382) <= not (a or b);
    outputs(383) <= not b;
    outputs(384) <= b and not a;
    outputs(385) <= not (a xor b);
    outputs(386) <= not b or a;
    outputs(387) <= not a or b;
    outputs(388) <= b;
    outputs(389) <= not a;
    outputs(390) <= a and b;
    outputs(391) <= not a or b;
    outputs(392) <= b;
    outputs(393) <= a;
    outputs(394) <= b;
    outputs(395) <= b;
    outputs(396) <= a;
    outputs(397) <= b;
    outputs(398) <= a;
    outputs(399) <= not (a or b);
    outputs(400) <= not a;
    outputs(401) <= not b;
    outputs(402) <= a xor b;
    outputs(403) <= a;
    outputs(404) <= a;
    outputs(405) <= not a;
    outputs(406) <= a;
    outputs(407) <= not a;
    outputs(408) <= a;
    outputs(409) <= not (a xor b);
    outputs(410) <= not (a or b);
    outputs(411) <= not a;
    outputs(412) <= not b;
    outputs(413) <= b;
    outputs(414) <= not a;
    outputs(415) <= a xor b;
    outputs(416) <= b;
    outputs(417) <= a and not b;
    outputs(418) <= not (a and b);
    outputs(419) <= not a;
    outputs(420) <= a;
    outputs(421) <= not (a or b);
    outputs(422) <= not (a and b);
    outputs(423) <= not b;
    outputs(424) <= a;
    outputs(425) <= not (a xor b);
    outputs(426) <= not a;
    outputs(427) <= not b;
    outputs(428) <= a xor b;
    outputs(429) <= a;
    outputs(430) <= not b;
    outputs(431) <= a xor b;
    outputs(432) <= a xor b;
    outputs(433) <= not b;
    outputs(434) <= b;
    outputs(435) <= not b;
    outputs(436) <= a and not b;
    outputs(437) <= not (a xor b);
    outputs(438) <= not (a xor b);
    outputs(439) <= a;
    outputs(440) <= not (a or b);
    outputs(441) <= b;
    outputs(442) <= not b;
    outputs(443) <= a xor b;
    outputs(444) <= a xor b;
    outputs(445) <= a and b;
    outputs(446) <= a xor b;
    outputs(447) <= not (a or b);
    outputs(448) <= not a or b;
    outputs(449) <= not a;
    outputs(450) <= a;
    outputs(451) <= not (a xor b);
    outputs(452) <= a xor b;
    outputs(453) <= not b;
    outputs(454) <= not a;
    outputs(455) <= b;
    outputs(456) <= not b;
    outputs(457) <= not a;
    outputs(458) <= a;
    outputs(459) <= a;
    outputs(460) <= not a;
    outputs(461) <= a and b;
    outputs(462) <= not (a xor b);
    outputs(463) <= a;
    outputs(464) <= a and not b;
    outputs(465) <= not (a xor b);
    outputs(466) <= b and not a;
    outputs(467) <= not a or b;
    outputs(468) <= not a;
    outputs(469) <= b;
    outputs(470) <= a and b;
    outputs(471) <= not (a or b);
    outputs(472) <= not a;
    outputs(473) <= a and b;
    outputs(474) <= not a;
    outputs(475) <= a;
    outputs(476) <= not a;
    outputs(477) <= a;
    outputs(478) <= not (a and b);
    outputs(479) <= a xor b;
    outputs(480) <= b and not a;
    outputs(481) <= b;
    outputs(482) <= a and b;
    outputs(483) <= a and not b;
    outputs(484) <= a;
    outputs(485) <= a;
    outputs(486) <= not b;
    outputs(487) <= a xor b;
    outputs(488) <= not (a xor b);
    outputs(489) <= a or b;
    outputs(490) <= not (a and b);
    outputs(491) <= not a;
    outputs(492) <= a;
    outputs(493) <= not b;
    outputs(494) <= b;
    outputs(495) <= b and not a;
    outputs(496) <= b;
    outputs(497) <= a;
    outputs(498) <= a;
    outputs(499) <= a and b;
    outputs(500) <= not a;
    outputs(501) <= not (a xor b);
    outputs(502) <= b;
    outputs(503) <= not (a or b);
    outputs(504) <= a xor b;
    outputs(505) <= not a;
    outputs(506) <= a xor b;
    outputs(507) <= not (a or b);
    outputs(508) <= a and not b;
    outputs(509) <= not a;
    outputs(510) <= b and not a;
    outputs(511) <= not (a xor b);
    outputs(512) <= a and b;
    outputs(513) <= not (a or b);
    outputs(514) <= a;
    outputs(515) <= b;
    outputs(516) <= a and not b;
    outputs(517) <= not b;
    outputs(518) <= a;
    outputs(519) <= b;
    outputs(520) <= b;
    outputs(521) <= not (a xor b);
    outputs(522) <= b and not a;
    outputs(523) <= not a;
    outputs(524) <= not (a or b);
    outputs(525) <= a;
    outputs(526) <= b;
    outputs(527) <= not b;
    outputs(528) <= not (a and b);
    outputs(529) <= not b;
    outputs(530) <= a and b;
    outputs(531) <= not a;
    outputs(532) <= not b;
    outputs(533) <= a and b;
    outputs(534) <= a;
    outputs(535) <= not b;
    outputs(536) <= not (a xor b);
    outputs(537) <= a and b;
    outputs(538) <= a;
    outputs(539) <= not a;
    outputs(540) <= not (a or b);
    outputs(541) <= not a;
    outputs(542) <= not a;
    outputs(543) <= a and not b;
    outputs(544) <= not (a xor b);
    outputs(545) <= a;
    outputs(546) <= not b;
    outputs(547) <= a and b;
    outputs(548) <= not (a or b);
    outputs(549) <= not (a xor b);
    outputs(550) <= not b;
    outputs(551) <= a;
    outputs(552) <= not (a or b);
    outputs(553) <= not b;
    outputs(554) <= a and not b;
    outputs(555) <= not a;
    outputs(556) <= not a;
    outputs(557) <= not a;
    outputs(558) <= a xor b;
    outputs(559) <= a xor b;
    outputs(560) <= a;
    outputs(561) <= not b;
    outputs(562) <= not b;
    outputs(563) <= a xor b;
    outputs(564) <= a;
    outputs(565) <= b;
    outputs(566) <= b;
    outputs(567) <= b;
    outputs(568) <= a;
    outputs(569) <= b;
    outputs(570) <= b;
    outputs(571) <= a and b;
    outputs(572) <= a xor b;
    outputs(573) <= not (a xor b);
    outputs(574) <= a xor b;
    outputs(575) <= a;
    outputs(576) <= a xor b;
    outputs(577) <= a;
    outputs(578) <= not (a xor b);
    outputs(579) <= a xor b;
    outputs(580) <= not b or a;
    outputs(581) <= not a;
    outputs(582) <= a xor b;
    outputs(583) <= a;
    outputs(584) <= a xor b;
    outputs(585) <= not a;
    outputs(586) <= a;
    outputs(587) <= a or b;
    outputs(588) <= not (a or b);
    outputs(589) <= a and not b;
    outputs(590) <= not a;
    outputs(591) <= not b;
    outputs(592) <= b;
    outputs(593) <= a;
    outputs(594) <= a;
    outputs(595) <= a xor b;
    outputs(596) <= not b;
    outputs(597) <= a and b;
    outputs(598) <= not b;
    outputs(599) <= not (a xor b);
    outputs(600) <= a;
    outputs(601) <= not b;
    outputs(602) <= not b;
    outputs(603) <= a xor b;
    outputs(604) <= b;
    outputs(605) <= not (a and b);
    outputs(606) <= a;
    outputs(607) <= a xor b;
    outputs(608) <= not (a or b);
    outputs(609) <= a and b;
    outputs(610) <= not a;
    outputs(611) <= b and not a;
    outputs(612) <= a xor b;
    outputs(613) <= b;
    outputs(614) <= not (a or b);
    outputs(615) <= b;
    outputs(616) <= not b;
    outputs(617) <= not (a xor b);
    outputs(618) <= not (a and b);
    outputs(619) <= not a;
    outputs(620) <= a and not b;
    outputs(621) <= a;
    outputs(622) <= a and not b;
    outputs(623) <= a and b;
    outputs(624) <= not (a xor b);
    outputs(625) <= a;
    outputs(626) <= not a;
    outputs(627) <= b;
    outputs(628) <= b;
    outputs(629) <= a;
    outputs(630) <= b;
    outputs(631) <= b;
    outputs(632) <= b;
    outputs(633) <= not (a xor b);
    outputs(634) <= b;
    outputs(635) <= not (a xor b);
    outputs(636) <= not (a or b);
    outputs(637) <= not (a xor b);
    outputs(638) <= not b;
    outputs(639) <= not a;
    outputs(640) <= not a;
    outputs(641) <= not (a xor b);
    outputs(642) <= not (a xor b);
    outputs(643) <= b and not a;
    outputs(644) <= a or b;
    outputs(645) <= a or b;
    outputs(646) <= b and not a;
    outputs(647) <= a and not b;
    outputs(648) <= b and not a;
    outputs(649) <= b;
    outputs(650) <= a and not b;
    outputs(651) <= not (a xor b);
    outputs(652) <= not b;
    outputs(653) <= not (a xor b);
    outputs(654) <= not (a xor b);
    outputs(655) <= a and b;
    outputs(656) <= not (a and b);
    outputs(657) <= b and not a;
    outputs(658) <= not a;
    outputs(659) <= not (a xor b);
    outputs(660) <= b and not a;
    outputs(661) <= a xor b;
    outputs(662) <= a or b;
    outputs(663) <= a xor b;
    outputs(664) <= a and not b;
    outputs(665) <= not (a xor b);
    outputs(666) <= a xor b;
    outputs(667) <= a and not b;
    outputs(668) <= a;
    outputs(669) <= not b;
    outputs(670) <= not b;
    outputs(671) <= a;
    outputs(672) <= a xor b;
    outputs(673) <= not a;
    outputs(674) <= not a;
    outputs(675) <= b;
    outputs(676) <= not (a xor b);
    outputs(677) <= b;
    outputs(678) <= a and b;
    outputs(679) <= not a;
    outputs(680) <= a and not b;
    outputs(681) <= a;
    outputs(682) <= not (a and b);
    outputs(683) <= not b or a;
    outputs(684) <= not a;
    outputs(685) <= not a or b;
    outputs(686) <= a xor b;
    outputs(687) <= not a;
    outputs(688) <= a;
    outputs(689) <= b and not a;
    outputs(690) <= b;
    outputs(691) <= not a;
    outputs(692) <= a xor b;
    outputs(693) <= b;
    outputs(694) <= a;
    outputs(695) <= not (a xor b);
    outputs(696) <= a xor b;
    outputs(697) <= b;
    outputs(698) <= not b;
    outputs(699) <= not b;
    outputs(700) <= a;
    outputs(701) <= not a;
    outputs(702) <= a and b;
    outputs(703) <= a xor b;
    outputs(704) <= b and not a;
    outputs(705) <= b;
    outputs(706) <= not a or b;
    outputs(707) <= a;
    outputs(708) <= not (a xor b);
    outputs(709) <= a and b;
    outputs(710) <= not a;
    outputs(711) <= a and b;
    outputs(712) <= not a;
    outputs(713) <= not (a or b);
    outputs(714) <= a and not b;
    outputs(715) <= not (a xor b);
    outputs(716) <= not b;
    outputs(717) <= a and b;
    outputs(718) <= not (a or b);
    outputs(719) <= not (a xor b);
    outputs(720) <= not b;
    outputs(721) <= b;
    outputs(722) <= not b;
    outputs(723) <= b and not a;
    outputs(724) <= a;
    outputs(725) <= a;
    outputs(726) <= not b;
    outputs(727) <= a;
    outputs(728) <= a;
    outputs(729) <= a xor b;
    outputs(730) <= a and b;
    outputs(731) <= not (a xor b);
    outputs(732) <= not a or b;
    outputs(733) <= a xor b;
    outputs(734) <= not (a or b);
    outputs(735) <= not (a xor b);
    outputs(736) <= not (a xor b);
    outputs(737) <= not (a xor b);
    outputs(738) <= not b;
    outputs(739) <= not (a xor b);
    outputs(740) <= not a;
    outputs(741) <= not a;
    outputs(742) <= a and not b;
    outputs(743) <= not a;
    outputs(744) <= a and b;
    outputs(745) <= a;
    outputs(746) <= b;
    outputs(747) <= b;
    outputs(748) <= a and b;
    outputs(749) <= a xor b;
    outputs(750) <= not (a xor b);
    outputs(751) <= b and not a;
    outputs(752) <= a;
    outputs(753) <= b and not a;
    outputs(754) <= not a;
    outputs(755) <= not (a xor b);
    outputs(756) <= not (a or b);
    outputs(757) <= a xor b;
    outputs(758) <= a;
    outputs(759) <= not a;
    outputs(760) <= a xor b;
    outputs(761) <= b and not a;
    outputs(762) <= b and not a;
    outputs(763) <= not a;
    outputs(764) <= a xor b;
    outputs(765) <= a;
    outputs(766) <= not b;
    outputs(767) <= not (a xor b);
    outputs(768) <= not b;
    outputs(769) <= not a;
    outputs(770) <= a and b;
    outputs(771) <= a;
    outputs(772) <= a and not b;
    outputs(773) <= a xor b;
    outputs(774) <= not a;
    outputs(775) <= b;
    outputs(776) <= b;
    outputs(777) <= not (a xor b);
    outputs(778) <= not b;
    outputs(779) <= not a;
    outputs(780) <= a and not b;
    outputs(781) <= a;
    outputs(782) <= a xor b;
    outputs(783) <= not (a xor b);
    outputs(784) <= not b;
    outputs(785) <= not (a xor b);
    outputs(786) <= not b;
    outputs(787) <= a and not b;
    outputs(788) <= a;
    outputs(789) <= b and not a;
    outputs(790) <= '0';
    outputs(791) <= a and not b;
    outputs(792) <= a and b;
    outputs(793) <= a and b;
    outputs(794) <= not b;
    outputs(795) <= b;
    outputs(796) <= a and b;
    outputs(797) <= not (a or b);
    outputs(798) <= a and b;
    outputs(799) <= b;
    outputs(800) <= a xor b;
    outputs(801) <= b;
    outputs(802) <= a and b;
    outputs(803) <= a;
    outputs(804) <= a and not b;
    outputs(805) <= not a;
    outputs(806) <= not a;
    outputs(807) <= not (a or b);
    outputs(808) <= not (a xor b);
    outputs(809) <= a xor b;
    outputs(810) <= not (a xor b);
    outputs(811) <= b and not a;
    outputs(812) <= not a;
    outputs(813) <= not b;
    outputs(814) <= b;
    outputs(815) <= not (a xor b);
    outputs(816) <= a and not b;
    outputs(817) <= not (a xor b);
    outputs(818) <= not a;
    outputs(819) <= b and not a;
    outputs(820) <= a and b;
    outputs(821) <= not b;
    outputs(822) <= not (a xor b);
    outputs(823) <= a;
    outputs(824) <= a;
    outputs(825) <= b;
    outputs(826) <= a xor b;
    outputs(827) <= a and not b;
    outputs(828) <= a xor b;
    outputs(829) <= a;
    outputs(830) <= a;
    outputs(831) <= not a;
    outputs(832) <= not (a xor b);
    outputs(833) <= not (a xor b);
    outputs(834) <= a and not b;
    outputs(835) <= not b;
    outputs(836) <= a;
    outputs(837) <= a xor b;
    outputs(838) <= not b;
    outputs(839) <= not b or a;
    outputs(840) <= not a;
    outputs(841) <= a and not b;
    outputs(842) <= b and not a;
    outputs(843) <= not (a and b);
    outputs(844) <= a xor b;
    outputs(845) <= a and b;
    outputs(846) <= not b;
    outputs(847) <= not a;
    outputs(848) <= b;
    outputs(849) <= not (a xor b);
    outputs(850) <= b;
    outputs(851) <= a xor b;
    outputs(852) <= b;
    outputs(853) <= a and b;
    outputs(854) <= a;
    outputs(855) <= b;
    outputs(856) <= b;
    outputs(857) <= b;
    outputs(858) <= not (a or b);
    outputs(859) <= b;
    outputs(860) <= not (a xor b);
    outputs(861) <= a;
    outputs(862) <= not b or a;
    outputs(863) <= not b;
    outputs(864) <= a;
    outputs(865) <= not (a or b);
    outputs(866) <= not (a xor b);
    outputs(867) <= b and not a;
    outputs(868) <= b;
    outputs(869) <= a and not b;
    outputs(870) <= b and not a;
    outputs(871) <= not a;
    outputs(872) <= a;
    outputs(873) <= b and not a;
    outputs(874) <= a and b;
    outputs(875) <= not (a xor b);
    outputs(876) <= not a;
    outputs(877) <= a and b;
    outputs(878) <= a and not b;
    outputs(879) <= not (a xor b);
    outputs(880) <= b and not a;
    outputs(881) <= a;
    outputs(882) <= a;
    outputs(883) <= not (a or b);
    outputs(884) <= not a or b;
    outputs(885) <= a and b;
    outputs(886) <= not (a xor b);
    outputs(887) <= a;
    outputs(888) <= not a;
    outputs(889) <= b and not a;
    outputs(890) <= not a;
    outputs(891) <= b;
    outputs(892) <= b and not a;
    outputs(893) <= not a;
    outputs(894) <= not b;
    outputs(895) <= a;
    outputs(896) <= not b or a;
    outputs(897) <= a and not b;
    outputs(898) <= a xor b;
    outputs(899) <= b;
    outputs(900) <= not (a xor b);
    outputs(901) <= not (a xor b);
    outputs(902) <= not a;
    outputs(903) <= b and not a;
    outputs(904) <= not b;
    outputs(905) <= a and b;
    outputs(906) <= a xor b;
    outputs(907) <= b;
    outputs(908) <= b and not a;
    outputs(909) <= b;
    outputs(910) <= a and not b;
    outputs(911) <= a and not b;
    outputs(912) <= a xor b;
    outputs(913) <= a xor b;
    outputs(914) <= a or b;
    outputs(915) <= a xor b;
    outputs(916) <= not b or a;
    outputs(917) <= not (a xor b);
    outputs(918) <= not (a or b);
    outputs(919) <= a and b;
    outputs(920) <= b;
    outputs(921) <= not b;
    outputs(922) <= not (a xor b);
    outputs(923) <= not (a xor b);
    outputs(924) <= a;
    outputs(925) <= b;
    outputs(926) <= a and b;
    outputs(927) <= not a;
    outputs(928) <= b;
    outputs(929) <= not (a or b);
    outputs(930) <= a and b;
    outputs(931) <= not a;
    outputs(932) <= a and b;
    outputs(933) <= not (a xor b);
    outputs(934) <= b;
    outputs(935) <= b and not a;
    outputs(936) <= a;
    outputs(937) <= a xor b;
    outputs(938) <= b and not a;
    outputs(939) <= a;
    outputs(940) <= a xor b;
    outputs(941) <= not (a xor b);
    outputs(942) <= b;
    outputs(943) <= a xor b;
    outputs(944) <= not (a or b);
    outputs(945) <= not a;
    outputs(946) <= not (a or b);
    outputs(947) <= not b;
    outputs(948) <= a;
    outputs(949) <= a and not b;
    outputs(950) <= a xor b;
    outputs(951) <= not (a or b);
    outputs(952) <= not a;
    outputs(953) <= not (a or b);
    outputs(954) <= b and not a;
    outputs(955) <= not (a xor b);
    outputs(956) <= b and not a;
    outputs(957) <= not (a or b);
    outputs(958) <= not (a or b);
    outputs(959) <= not b;
    outputs(960) <= a;
    outputs(961) <= b;
    outputs(962) <= not (a xor b);
    outputs(963) <= not a;
    outputs(964) <= a;
    outputs(965) <= not b;
    outputs(966) <= a and not b;
    outputs(967) <= a and not b;
    outputs(968) <= b;
    outputs(969) <= a;
    outputs(970) <= not (a xor b);
    outputs(971) <= not a;
    outputs(972) <= not (a or b);
    outputs(973) <= a and b;
    outputs(974) <= not a;
    outputs(975) <= a;
    outputs(976) <= a and not b;
    outputs(977) <= not (a or b);
    outputs(978) <= a;
    outputs(979) <= not (a or b);
    outputs(980) <= b and not a;
    outputs(981) <= not a;
    outputs(982) <= b;
    outputs(983) <= not (a or b);
    outputs(984) <= a xor b;
    outputs(985) <= a and b;
    outputs(986) <= a xor b;
    outputs(987) <= a xor b;
    outputs(988) <= a xor b;
    outputs(989) <= a;
    outputs(990) <= not (a or b);
    outputs(991) <= not b;
    outputs(992) <= b and not a;
    outputs(993) <= a;
    outputs(994) <= a xor b;
    outputs(995) <= b;
    outputs(996) <= b and not a;
    outputs(997) <= b;
    outputs(998) <= not b;
    outputs(999) <= a;
    outputs(1000) <= a;
    outputs(1001) <= not (a xor b);
    outputs(1002) <= not b;
    outputs(1003) <= a;
    outputs(1004) <= not (a or b);
    outputs(1005) <= not a;
    outputs(1006) <= b;
    outputs(1007) <= not (a xor b);
    outputs(1008) <= not (a xor b);
    outputs(1009) <= b and not a;
    outputs(1010) <= not (a xor b);
    outputs(1011) <= a and not b;
    outputs(1012) <= b and not a;
    outputs(1013) <= a and b;
    outputs(1014) <= not (a or b);
    outputs(1015) <= b and not a;
    outputs(1016) <= a and not b;
    outputs(1017) <= b;
    outputs(1018) <= not (a xor b);
    outputs(1019) <= a and b;
    outputs(1020) <= not b;
    outputs(1021) <= b;
    outputs(1022) <= a and not b;
    outputs(1023) <= a xor b;
    outputs(1024) <= not (a xor b);
    outputs(1025) <= b;
    outputs(1026) <= a;
    outputs(1027) <= b;
    outputs(1028) <= not (a or b);
    outputs(1029) <= not (a xor b);
    outputs(1030) <= not b;
    outputs(1031) <= a xor b;
    outputs(1032) <= not a;
    outputs(1033) <= a;
    outputs(1034) <= a and b;
    outputs(1035) <= not a;
    outputs(1036) <= a xor b;
    outputs(1037) <= not (a xor b);
    outputs(1038) <= a and b;
    outputs(1039) <= b and not a;
    outputs(1040) <= b;
    outputs(1041) <= a;
    outputs(1042) <= a and b;
    outputs(1043) <= a xor b;
    outputs(1044) <= not b;
    outputs(1045) <= not (a xor b);
    outputs(1046) <= not a;
    outputs(1047) <= a and b;
    outputs(1048) <= a xor b;
    outputs(1049) <= not b;
    outputs(1050) <= b and not a;
    outputs(1051) <= not (a xor b);
    outputs(1052) <= a;
    outputs(1053) <= not (a xor b);
    outputs(1054) <= not a or b;
    outputs(1055) <= not (a xor b);
    outputs(1056) <= a;
    outputs(1057) <= b and not a;
    outputs(1058) <= not (a xor b);
    outputs(1059) <= not a;
    outputs(1060) <= not b;
    outputs(1061) <= b and not a;
    outputs(1062) <= a and b;
    outputs(1063) <= a xor b;
    outputs(1064) <= a or b;
    outputs(1065) <= not (a xor b);
    outputs(1066) <= a;
    outputs(1067) <= not (a or b);
    outputs(1068) <= not a;
    outputs(1069) <= not (a xor b);
    outputs(1070) <= not b;
    outputs(1071) <= not b;
    outputs(1072) <= not b;
    outputs(1073) <= a;
    outputs(1074) <= not a;
    outputs(1075) <= not b;
    outputs(1076) <= a and not b;
    outputs(1077) <= not b or a;
    outputs(1078) <= not (a xor b);
    outputs(1079) <= not a or b;
    outputs(1080) <= a and not b;
    outputs(1081) <= not b;
    outputs(1082) <= a;
    outputs(1083) <= a xor b;
    outputs(1084) <= not a;
    outputs(1085) <= not (a xor b);
    outputs(1086) <= b;
    outputs(1087) <= a xor b;
    outputs(1088) <= not b;
    outputs(1089) <= not a or b;
    outputs(1090) <= a and not b;
    outputs(1091) <= a;
    outputs(1092) <= not (a xor b);
    outputs(1093) <= b;
    outputs(1094) <= a;
    outputs(1095) <= not (a xor b);
    outputs(1096) <= not (a or b);
    outputs(1097) <= not (a or b);
    outputs(1098) <= b and not a;
    outputs(1099) <= not b or a;
    outputs(1100) <= not (a or b);
    outputs(1101) <= a and b;
    outputs(1102) <= a;
    outputs(1103) <= not b or a;
    outputs(1104) <= not (a or b);
    outputs(1105) <= not a;
    outputs(1106) <= not b;
    outputs(1107) <= b;
    outputs(1108) <= not a;
    outputs(1109) <= a;
    outputs(1110) <= a;
    outputs(1111) <= b;
    outputs(1112) <= a and not b;
    outputs(1113) <= a;
    outputs(1114) <= not a;
    outputs(1115) <= not (a or b);
    outputs(1116) <= not (a xor b);
    outputs(1117) <= a xor b;
    outputs(1118) <= '0';
    outputs(1119) <= not b;
    outputs(1120) <= a;
    outputs(1121) <= a and b;
    outputs(1122) <= a;
    outputs(1123) <= not b;
    outputs(1124) <= a and not b;
    outputs(1125) <= a and not b;
    outputs(1126) <= not a;
    outputs(1127) <= b and not a;
    outputs(1128) <= a and b;
    outputs(1129) <= not (a or b);
    outputs(1130) <= b and not a;
    outputs(1131) <= not (a or b);
    outputs(1132) <= not (a xor b);
    outputs(1133) <= a and b;
    outputs(1134) <= a and not b;
    outputs(1135) <= b;
    outputs(1136) <= not a;
    outputs(1137) <= not (a xor b);
    outputs(1138) <= a and b;
    outputs(1139) <= a and b;
    outputs(1140) <= a xor b;
    outputs(1141) <= not b;
    outputs(1142) <= not a;
    outputs(1143) <= not (a xor b);
    outputs(1144) <= b;
    outputs(1145) <= a and b;
    outputs(1146) <= not (a or b);
    outputs(1147) <= a and not b;
    outputs(1148) <= not (a or b);
    outputs(1149) <= a xor b;
    outputs(1150) <= a and not b;
    outputs(1151) <= b;
    outputs(1152) <= a xor b;
    outputs(1153) <= a xor b;
    outputs(1154) <= a xor b;
    outputs(1155) <= a and not b;
    outputs(1156) <= not a or b;
    outputs(1157) <= not a;
    outputs(1158) <= b;
    outputs(1159) <= b;
    outputs(1160) <= not a;
    outputs(1161) <= a and b;
    outputs(1162) <= not (a or b);
    outputs(1163) <= not (a xor b);
    outputs(1164) <= a and not b;
    outputs(1165) <= not a or b;
    outputs(1166) <= not a;
    outputs(1167) <= not b;
    outputs(1168) <= a and not b;
    outputs(1169) <= a and not b;
    outputs(1170) <= not a;
    outputs(1171) <= b;
    outputs(1172) <= b;
    outputs(1173) <= b;
    outputs(1174) <= b;
    outputs(1175) <= not b;
    outputs(1176) <= a xor b;
    outputs(1177) <= b and not a;
    outputs(1178) <= a and not b;
    outputs(1179) <= not (a or b);
    outputs(1180) <= not (a xor b);
    outputs(1181) <= a and not b;
    outputs(1182) <= not b;
    outputs(1183) <= b;
    outputs(1184) <= b;
    outputs(1185) <= a and not b;
    outputs(1186) <= not (a or b);
    outputs(1187) <= b;
    outputs(1188) <= not a;
    outputs(1189) <= a and b;
    outputs(1190) <= not b;
    outputs(1191) <= not a;
    outputs(1192) <= b;
    outputs(1193) <= not (a or b);
    outputs(1194) <= a xor b;
    outputs(1195) <= a xor b;
    outputs(1196) <= a and not b;
    outputs(1197) <= b;
    outputs(1198) <= a xor b;
    outputs(1199) <= b and not a;
    outputs(1200) <= a and not b;
    outputs(1201) <= not (a xor b);
    outputs(1202) <= not (a or b);
    outputs(1203) <= not (a xor b);
    outputs(1204) <= b and not a;
    outputs(1205) <= a and b;
    outputs(1206) <= not (a xor b);
    outputs(1207) <= a and b;
    outputs(1208) <= b and not a;
    outputs(1209) <= a and b;
    outputs(1210) <= not a or b;
    outputs(1211) <= not b;
    outputs(1212) <= a;
    outputs(1213) <= b;
    outputs(1214) <= not a;
    outputs(1215) <= not (a or b);
    outputs(1216) <= a and b;
    outputs(1217) <= a xor b;
    outputs(1218) <= not (a xor b);
    outputs(1219) <= not (a or b);
    outputs(1220) <= not (a xor b);
    outputs(1221) <= a xor b;
    outputs(1222) <= b;
    outputs(1223) <= not (a and b);
    outputs(1224) <= not b;
    outputs(1225) <= a and not b;
    outputs(1226) <= not a;
    outputs(1227) <= not a;
    outputs(1228) <= a xor b;
    outputs(1229) <= '0';
    outputs(1230) <= not (a or b);
    outputs(1231) <= not (a xor b);
    outputs(1232) <= not (a or b);
    outputs(1233) <= a xor b;
    outputs(1234) <= b;
    outputs(1235) <= not b;
    outputs(1236) <= a and not b;
    outputs(1237) <= not b;
    outputs(1238) <= not (a or b);
    outputs(1239) <= a and not b;
    outputs(1240) <= a and b;
    outputs(1241) <= not (a xor b);
    outputs(1242) <= b and not a;
    outputs(1243) <= b and not a;
    outputs(1244) <= b and not a;
    outputs(1245) <= a xor b;
    outputs(1246) <= a xor b;
    outputs(1247) <= a;
    outputs(1248) <= b and not a;
    outputs(1249) <= a;
    outputs(1250) <= b;
    outputs(1251) <= not b;
    outputs(1252) <= b and not a;
    outputs(1253) <= not (a and b);
    outputs(1254) <= b;
    outputs(1255) <= not a;
    outputs(1256) <= a xor b;
    outputs(1257) <= b and not a;
    outputs(1258) <= b;
    outputs(1259) <= b;
    outputs(1260) <= not b or a;
    outputs(1261) <= not b;
    outputs(1262) <= a xor b;
    outputs(1263) <= not (a xor b);
    outputs(1264) <= b and not a;
    outputs(1265) <= not b;
    outputs(1266) <= not (a or b);
    outputs(1267) <= not (a xor b);
    outputs(1268) <= not (a xor b);
    outputs(1269) <= a and not b;
    outputs(1270) <= not (a xor b);
    outputs(1271) <= not (a and b);
    outputs(1272) <= b and not a;
    outputs(1273) <= not (a xor b);
    outputs(1274) <= not (a and b);
    outputs(1275) <= not (a or b);
    outputs(1276) <= not (a or b);
    outputs(1277) <= not (a or b);
    outputs(1278) <= not (a or b);
    outputs(1279) <= a and not b;
    outputs(1280) <= b;
    outputs(1281) <= a and b;
    outputs(1282) <= a and not b;
    outputs(1283) <= a xor b;
    outputs(1284) <= a;
    outputs(1285) <= a;
    outputs(1286) <= a;
    outputs(1287) <= b;
    outputs(1288) <= b and not a;
    outputs(1289) <= a;
    outputs(1290) <= not b;
    outputs(1291) <= not (a xor b);
    outputs(1292) <= a xor b;
    outputs(1293) <= a and not b;
    outputs(1294) <= b and not a;
    outputs(1295) <= not (a xor b);
    outputs(1296) <= b;
    outputs(1297) <= not b;
    outputs(1298) <= not (a or b);
    outputs(1299) <= a;
    outputs(1300) <= not b;
    outputs(1301) <= a and b;
    outputs(1302) <= not (a xor b);
    outputs(1303) <= b and not a;
    outputs(1304) <= b;
    outputs(1305) <= not (a xor b);
    outputs(1306) <= not (a xor b);
    outputs(1307) <= not a;
    outputs(1308) <= not (a xor b);
    outputs(1309) <= not b;
    outputs(1310) <= not b;
    outputs(1311) <= not (a xor b);
    outputs(1312) <= not (a or b);
    outputs(1313) <= a xor b;
    outputs(1314) <= not (a xor b);
    outputs(1315) <= not a;
    outputs(1316) <= not a;
    outputs(1317) <= not (a or b);
    outputs(1318) <= b;
    outputs(1319) <= not (a or b);
    outputs(1320) <= a xor b;
    outputs(1321) <= not a;
    outputs(1322) <= a xor b;
    outputs(1323) <= b and not a;
    outputs(1324) <= not b;
    outputs(1325) <= not (a xor b);
    outputs(1326) <= not a;
    outputs(1327) <= b;
    outputs(1328) <= a;
    outputs(1329) <= a;
    outputs(1330) <= not a;
    outputs(1331) <= not (a or b);
    outputs(1332) <= a xor b;
    outputs(1333) <= a and not b;
    outputs(1334) <= a xor b;
    outputs(1335) <= not a;
    outputs(1336) <= not (a or b);
    outputs(1337) <= b;
    outputs(1338) <= a and b;
    outputs(1339) <= a and b;
    outputs(1340) <= a xor b;
    outputs(1341) <= a;
    outputs(1342) <= a and not b;
    outputs(1343) <= not b;
    outputs(1344) <= a xor b;
    outputs(1345) <= b;
    outputs(1346) <= not b;
    outputs(1347) <= a and b;
    outputs(1348) <= a or b;
    outputs(1349) <= not (a or b);
    outputs(1350) <= a xor b;
    outputs(1351) <= not b;
    outputs(1352) <= a and b;
    outputs(1353) <= not (a xor b);
    outputs(1354) <= not b;
    outputs(1355) <= not b;
    outputs(1356) <= b;
    outputs(1357) <= not (a xor b);
    outputs(1358) <= a and b;
    outputs(1359) <= not (a xor b);
    outputs(1360) <= not b;
    outputs(1361) <= a xor b;
    outputs(1362) <= b and not a;
    outputs(1363) <= not (a or b);
    outputs(1364) <= b and not a;
    outputs(1365) <= a;
    outputs(1366) <= not b;
    outputs(1367) <= not b;
    outputs(1368) <= a;
    outputs(1369) <= a and not b;
    outputs(1370) <= a and not b;
    outputs(1371) <= not a;
    outputs(1372) <= a;
    outputs(1373) <= b;
    outputs(1374) <= a and not b;
    outputs(1375) <= not (a or b);
    outputs(1376) <= not b;
    outputs(1377) <= b;
    outputs(1378) <= b;
    outputs(1379) <= a and not b;
    outputs(1380) <= a xor b;
    outputs(1381) <= a xor b;
    outputs(1382) <= b;
    outputs(1383) <= not (a xor b);
    outputs(1384) <= not b;
    outputs(1385) <= a and b;
    outputs(1386) <= not a;
    outputs(1387) <= a;
    outputs(1388) <= a and not b;
    outputs(1389) <= not (a or b);
    outputs(1390) <= not a;
    outputs(1391) <= not (a xor b);
    outputs(1392) <= a;
    outputs(1393) <= a and not b;
    outputs(1394) <= not b;
    outputs(1395) <= b and not a;
    outputs(1396) <= b;
    outputs(1397) <= a xor b;
    outputs(1398) <= b;
    outputs(1399) <= a and b;
    outputs(1400) <= a xor b;
    outputs(1401) <= a and b;
    outputs(1402) <= not (a or b);
    outputs(1403) <= a and b;
    outputs(1404) <= not a;
    outputs(1405) <= a and b;
    outputs(1406) <= not b or a;
    outputs(1407) <= a;
    outputs(1408) <= a and not b;
    outputs(1409) <= a xor b;
    outputs(1410) <= a xor b;
    outputs(1411) <= a and not b;
    outputs(1412) <= '0';
    outputs(1413) <= not (a or b);
    outputs(1414) <= not (a xor b);
    outputs(1415) <= not (a xor b);
    outputs(1416) <= not a or b;
    outputs(1417) <= not a;
    outputs(1418) <= not (a xor b);
    outputs(1419) <= a;
    outputs(1420) <= not a;
    outputs(1421) <= b;
    outputs(1422) <= not (a xor b);
    outputs(1423) <= a;
    outputs(1424) <= a and b;
    outputs(1425) <= a and not b;
    outputs(1426) <= not (a xor b);
    outputs(1427) <= a and not b;
    outputs(1428) <= a and b;
    outputs(1429) <= not a;
    outputs(1430) <= a and b;
    outputs(1431) <= a and not b;
    outputs(1432) <= a xor b;
    outputs(1433) <= a;
    outputs(1434) <= not (a xor b);
    outputs(1435) <= b;
    outputs(1436) <= b;
    outputs(1437) <= a xor b;
    outputs(1438) <= a and not b;
    outputs(1439) <= a;
    outputs(1440) <= a xor b;
    outputs(1441) <= b;
    outputs(1442) <= not (a or b);
    outputs(1443) <= a and not b;
    outputs(1444) <= a and b;
    outputs(1445) <= not a;
    outputs(1446) <= b and not a;
    outputs(1447) <= not b;
    outputs(1448) <= not (a or b);
    outputs(1449) <= a xor b;
    outputs(1450) <= b;
    outputs(1451) <= a and not b;
    outputs(1452) <= a or b;
    outputs(1453) <= not b;
    outputs(1454) <= a xor b;
    outputs(1455) <= not (a or b);
    outputs(1456) <= not a or b;
    outputs(1457) <= not a;
    outputs(1458) <= not (a or b);
    outputs(1459) <= a xor b;
    outputs(1460) <= a xor b;
    outputs(1461) <= not (a xor b);
    outputs(1462) <= not b;
    outputs(1463) <= b;
    outputs(1464) <= not (a or b);
    outputs(1465) <= '0';
    outputs(1466) <= not a or b;
    outputs(1467) <= b and not a;
    outputs(1468) <= b and not a;
    outputs(1469) <= a xor b;
    outputs(1470) <= not (a and b);
    outputs(1471) <= not (a xor b);
    outputs(1472) <= a xor b;
    outputs(1473) <= a and not b;
    outputs(1474) <= a and b;
    outputs(1475) <= a and not b;
    outputs(1476) <= a and b;
    outputs(1477) <= not (a or b);
    outputs(1478) <= b;
    outputs(1479) <= b and not a;
    outputs(1480) <= b and not a;
    outputs(1481) <= b;
    outputs(1482) <= a;
    outputs(1483) <= b;
    outputs(1484) <= b and not a;
    outputs(1485) <= b and not a;
    outputs(1486) <= b;
    outputs(1487) <= not (a or b);
    outputs(1488) <= not (a or b);
    outputs(1489) <= not (a xor b);
    outputs(1490) <= a and b;
    outputs(1491) <= not (a xor b);
    outputs(1492) <= b;
    outputs(1493) <= b;
    outputs(1494) <= not (a xor b);
    outputs(1495) <= b and not a;
    outputs(1496) <= b;
    outputs(1497) <= b and not a;
    outputs(1498) <= a;
    outputs(1499) <= a and not b;
    outputs(1500) <= a;
    outputs(1501) <= a and not b;
    outputs(1502) <= b;
    outputs(1503) <= not (a and b);
    outputs(1504) <= not (a or b);
    outputs(1505) <= a;
    outputs(1506) <= b and not a;
    outputs(1507) <= a and b;
    outputs(1508) <= b;
    outputs(1509) <= not (a or b);
    outputs(1510) <= a and not b;
    outputs(1511) <= not (a xor b);
    outputs(1512) <= a xor b;
    outputs(1513) <= a and not b;
    outputs(1514) <= not (a and b);
    outputs(1515) <= a;
    outputs(1516) <= a and b;
    outputs(1517) <= a and not b;
    outputs(1518) <= not (a or b);
    outputs(1519) <= not b or a;
    outputs(1520) <= a and b;
    outputs(1521) <= b and not a;
    outputs(1522) <= not b;
    outputs(1523) <= b;
    outputs(1524) <= not (a xor b);
    outputs(1525) <= b and not a;
    outputs(1526) <= a;
    outputs(1527) <= not a;
    outputs(1528) <= a xor b;
    outputs(1529) <= not b;
    outputs(1530) <= b and not a;
    outputs(1531) <= a and not b;
    outputs(1532) <= a and not b;
    outputs(1533) <= not a;
    outputs(1534) <= a and not b;
    outputs(1535) <= not b;
    outputs(1536) <= not a;
    outputs(1537) <= a and b;
    outputs(1538) <= not (a xor b);
    outputs(1539) <= a and not b;
    outputs(1540) <= b;
    outputs(1541) <= not a;
    outputs(1542) <= a;
    outputs(1543) <= b;
    outputs(1544) <= not (a or b);
    outputs(1545) <= a;
    outputs(1546) <= not a;
    outputs(1547) <= not a;
    outputs(1548) <= not (a xor b);
    outputs(1549) <= a;
    outputs(1550) <= a;
    outputs(1551) <= not (a xor b);
    outputs(1552) <= not a;
    outputs(1553) <= b;
    outputs(1554) <= not a;
    outputs(1555) <= not b;
    outputs(1556) <= not (a xor b);
    outputs(1557) <= a xor b;
    outputs(1558) <= not (a and b);
    outputs(1559) <= not a;
    outputs(1560) <= a or b;
    outputs(1561) <= not b;
    outputs(1562) <= not b;
    outputs(1563) <= a xor b;
    outputs(1564) <= not a;
    outputs(1565) <= a xor b;
    outputs(1566) <= a;
    outputs(1567) <= not (a xor b);
    outputs(1568) <= not (a xor b);
    outputs(1569) <= a;
    outputs(1570) <= not (a xor b);
    outputs(1571) <= a;
    outputs(1572) <= not (a xor b);
    outputs(1573) <= b and not a;
    outputs(1574) <= not a;
    outputs(1575) <= b;
    outputs(1576) <= b;
    outputs(1577) <= not (a xor b);
    outputs(1578) <= not (a or b);
    outputs(1579) <= not (a or b);
    outputs(1580) <= a xor b;
    outputs(1581) <= not a;
    outputs(1582) <= a;
    outputs(1583) <= a and b;
    outputs(1584) <= b;
    outputs(1585) <= not b;
    outputs(1586) <= not (a xor b);
    outputs(1587) <= a xor b;
    outputs(1588) <= a and b;
    outputs(1589) <= a xor b;
    outputs(1590) <= not (a or b);
    outputs(1591) <= b;
    outputs(1592) <= not (a xor b);
    outputs(1593) <= b;
    outputs(1594) <= a;
    outputs(1595) <= not (a xor b);
    outputs(1596) <= b;
    outputs(1597) <= not a;
    outputs(1598) <= not a;
    outputs(1599) <= a xor b;
    outputs(1600) <= not b or a;
    outputs(1601) <= a;
    outputs(1602) <= not (a or b);
    outputs(1603) <= not (a xor b);
    outputs(1604) <= not (a xor b);
    outputs(1605) <= b and not a;
    outputs(1606) <= b;
    outputs(1607) <= not b;
    outputs(1608) <= a xor b;
    outputs(1609) <= a;
    outputs(1610) <= not (a or b);
    outputs(1611) <= b and not a;
    outputs(1612) <= a xor b;
    outputs(1613) <= b;
    outputs(1614) <= a;
    outputs(1615) <= a and b;
    outputs(1616) <= b;
    outputs(1617) <= not b;
    outputs(1618) <= not b;
    outputs(1619) <= a or b;
    outputs(1620) <= b;
    outputs(1621) <= a;
    outputs(1622) <= a and not b;
    outputs(1623) <= a xor b;
    outputs(1624) <= a xor b;
    outputs(1625) <= not (a xor b);
    outputs(1626) <= a;
    outputs(1627) <= not b;
    outputs(1628) <= not (a xor b);
    outputs(1629) <= not a;
    outputs(1630) <= b;
    outputs(1631) <= not b;
    outputs(1632) <= a or b;
    outputs(1633) <= not (a xor b);
    outputs(1634) <= not a;
    outputs(1635) <= not b or a;
    outputs(1636) <= not b;
    outputs(1637) <= not (a xor b);
    outputs(1638) <= a xor b;
    outputs(1639) <= not (a xor b);
    outputs(1640) <= not a;
    outputs(1641) <= not a;
    outputs(1642) <= not b or a;
    outputs(1643) <= a xor b;
    outputs(1644) <= a and b;
    outputs(1645) <= a xor b;
    outputs(1646) <= a xor b;
    outputs(1647) <= a xor b;
    outputs(1648) <= not b;
    outputs(1649) <= not b;
    outputs(1650) <= a and not b;
    outputs(1651) <= not a;
    outputs(1652) <= not (a xor b);
    outputs(1653) <= a xor b;
    outputs(1654) <= not a;
    outputs(1655) <= b and not a;
    outputs(1656) <= a;
    outputs(1657) <= a xor b;
    outputs(1658) <= b;
    outputs(1659) <= a xor b;
    outputs(1660) <= not b;
    outputs(1661) <= not (a and b);
    outputs(1662) <= b;
    outputs(1663) <= b;
    outputs(1664) <= a;
    outputs(1665) <= not b or a;
    outputs(1666) <= a;
    outputs(1667) <= not (a xor b);
    outputs(1668) <= not (a and b);
    outputs(1669) <= not a;
    outputs(1670) <= a;
    outputs(1671) <= not a;
    outputs(1672) <= a or b;
    outputs(1673) <= not a;
    outputs(1674) <= a and not b;
    outputs(1675) <= not a;
    outputs(1676) <= not a;
    outputs(1677) <= a xor b;
    outputs(1678) <= a xor b;
    outputs(1679) <= not (a xor b);
    outputs(1680) <= a xor b;
    outputs(1681) <= not (a xor b);
    outputs(1682) <= a;
    outputs(1683) <= not a;
    outputs(1684) <= a;
    outputs(1685) <= not (a or b);
    outputs(1686) <= b;
    outputs(1687) <= b;
    outputs(1688) <= not a;
    outputs(1689) <= a;
    outputs(1690) <= not a;
    outputs(1691) <= not b or a;
    outputs(1692) <= b;
    outputs(1693) <= a or b;
    outputs(1694) <= a;
    outputs(1695) <= b;
    outputs(1696) <= a and not b;
    outputs(1697) <= not a;
    outputs(1698) <= not b;
    outputs(1699) <= not (a xor b);
    outputs(1700) <= not (a and b);
    outputs(1701) <= a and b;
    outputs(1702) <= not (a xor b);
    outputs(1703) <= a xor b;
    outputs(1704) <= a and not b;
    outputs(1705) <= not (a or b);
    outputs(1706) <= not a;
    outputs(1707) <= not b;
    outputs(1708) <= not a;
    outputs(1709) <= not a;
    outputs(1710) <= not (a xor b);
    outputs(1711) <= not a;
    outputs(1712) <= a or b;
    outputs(1713) <= not b;
    outputs(1714) <= b;
    outputs(1715) <= b;
    outputs(1716) <= a or b;
    outputs(1717) <= not b;
    outputs(1718) <= a;
    outputs(1719) <= not a;
    outputs(1720) <= a;
    outputs(1721) <= a xor b;
    outputs(1722) <= not a or b;
    outputs(1723) <= b;
    outputs(1724) <= not (a or b);
    outputs(1725) <= not (a and b);
    outputs(1726) <= not (a xor b);
    outputs(1727) <= not (a or b);
    outputs(1728) <= b;
    outputs(1729) <= not a;
    outputs(1730) <= not b;
    outputs(1731) <= a;
    outputs(1732) <= a or b;
    outputs(1733) <= not (a xor b);
    outputs(1734) <= a and not b;
    outputs(1735) <= a;
    outputs(1736) <= a xor b;
    outputs(1737) <= a xor b;
    outputs(1738) <= not (a or b);
    outputs(1739) <= not a;
    outputs(1740) <= a;
    outputs(1741) <= not a;
    outputs(1742) <= not (a xor b);
    outputs(1743) <= '0';
    outputs(1744) <= a xor b;
    outputs(1745) <= not (a and b);
    outputs(1746) <= not b;
    outputs(1747) <= a or b;
    outputs(1748) <= a;
    outputs(1749) <= not (a xor b);
    outputs(1750) <= a xor b;
    outputs(1751) <= not a;
    outputs(1752) <= a;
    outputs(1753) <= a;
    outputs(1754) <= not a or b;
    outputs(1755) <= a;
    outputs(1756) <= not a;
    outputs(1757) <= a xor b;
    outputs(1758) <= b and not a;
    outputs(1759) <= b;
    outputs(1760) <= a xor b;
    outputs(1761) <= not b;
    outputs(1762) <= not (a xor b);
    outputs(1763) <= a and not b;
    outputs(1764) <= b;
    outputs(1765) <= a xor b;
    outputs(1766) <= a xor b;
    outputs(1767) <= not b;
    outputs(1768) <= not b;
    outputs(1769) <= not a;
    outputs(1770) <= a and not b;
    outputs(1771) <= a or b;
    outputs(1772) <= not b;
    outputs(1773) <= not (a xor b);
    outputs(1774) <= b and not a;
    outputs(1775) <= b;
    outputs(1776) <= a xor b;
    outputs(1777) <= a xor b;
    outputs(1778) <= a xor b;
    outputs(1779) <= a xor b;
    outputs(1780) <= not a;
    outputs(1781) <= not (a or b);
    outputs(1782) <= not a;
    outputs(1783) <= not (a or b);
    outputs(1784) <= a;
    outputs(1785) <= not (a xor b);
    outputs(1786) <= a and not b;
    outputs(1787) <= a;
    outputs(1788) <= a and b;
    outputs(1789) <= a xor b;
    outputs(1790) <= b;
    outputs(1791) <= not b;
    outputs(1792) <= not b or a;
    outputs(1793) <= a or b;
    outputs(1794) <= not (a xor b);
    outputs(1795) <= a and not b;
    outputs(1796) <= not a;
    outputs(1797) <= a;
    outputs(1798) <= a xor b;
    outputs(1799) <= a and b;
    outputs(1800) <= a xor b;
    outputs(1801) <= a;
    outputs(1802) <= not (a xor b);
    outputs(1803) <= a and b;
    outputs(1804) <= a and b;
    outputs(1805) <= b and not a;
    outputs(1806) <= a;
    outputs(1807) <= not (a xor b);
    outputs(1808) <= a;
    outputs(1809) <= a or b;
    outputs(1810) <= not (a xor b);
    outputs(1811) <= b;
    outputs(1812) <= not b or a;
    outputs(1813) <= not b or a;
    outputs(1814) <= not a or b;
    outputs(1815) <= a or b;
    outputs(1816) <= a xor b;
    outputs(1817) <= a xor b;
    outputs(1818) <= a or b;
    outputs(1819) <= not b;
    outputs(1820) <= not b;
    outputs(1821) <= a;
    outputs(1822) <= a;
    outputs(1823) <= not b;
    outputs(1824) <= not a;
    outputs(1825) <= a xor b;
    outputs(1826) <= a;
    outputs(1827) <= not a;
    outputs(1828) <= a xor b;
    outputs(1829) <= not b;
    outputs(1830) <= a xor b;
    outputs(1831) <= a xor b;
    outputs(1832) <= a;
    outputs(1833) <= not a;
    outputs(1834) <= not (a xor b);
    outputs(1835) <= not a or b;
    outputs(1836) <= a or b;
    outputs(1837) <= not (a xor b);
    outputs(1838) <= b and not a;
    outputs(1839) <= not (a xor b);
    outputs(1840) <= not a;
    outputs(1841) <= b;
    outputs(1842) <= a xor b;
    outputs(1843) <= a xor b;
    outputs(1844) <= not (a xor b);
    outputs(1845) <= not (a xor b);
    outputs(1846) <= a;
    outputs(1847) <= a and not b;
    outputs(1848) <= not b or a;
    outputs(1849) <= b;
    outputs(1850) <= a xor b;
    outputs(1851) <= not a;
    outputs(1852) <= a xor b;
    outputs(1853) <= a;
    outputs(1854) <= not b or a;
    outputs(1855) <= not b;
    outputs(1856) <= not (a or b);
    outputs(1857) <= b;
    outputs(1858) <= a xor b;
    outputs(1859) <= not b;
    outputs(1860) <= b and not a;
    outputs(1861) <= a and b;
    outputs(1862) <= b and not a;
    outputs(1863) <= a and not b;
    outputs(1864) <= not b;
    outputs(1865) <= not b;
    outputs(1866) <= a xor b;
    outputs(1867) <= b;
    outputs(1868) <= a xor b;
    outputs(1869) <= a;
    outputs(1870) <= not b;
    outputs(1871) <= a;
    outputs(1872) <= b and not a;
    outputs(1873) <= not a;
    outputs(1874) <= not a;
    outputs(1875) <= not b;
    outputs(1876) <= b;
    outputs(1877) <= b;
    outputs(1878) <= not (a and b);
    outputs(1879) <= not b;
    outputs(1880) <= b;
    outputs(1881) <= not b;
    outputs(1882) <= not (a xor b);
    outputs(1883) <= a;
    outputs(1884) <= a xor b;
    outputs(1885) <= not a;
    outputs(1886) <= b;
    outputs(1887) <= not a;
    outputs(1888) <= b;
    outputs(1889) <= not (a xor b);
    outputs(1890) <= b;
    outputs(1891) <= not (a xor b);
    outputs(1892) <= a xor b;
    outputs(1893) <= not a;
    outputs(1894) <= a xor b;
    outputs(1895) <= not b;
    outputs(1896) <= not (a xor b);
    outputs(1897) <= not a;
    outputs(1898) <= a xor b;
    outputs(1899) <= not (a xor b);
    outputs(1900) <= b;
    outputs(1901) <= a and not b;
    outputs(1902) <= b;
    outputs(1903) <= not (a or b);
    outputs(1904) <= not (a xor b);
    outputs(1905) <= not b;
    outputs(1906) <= not b;
    outputs(1907) <= not (a xor b);
    outputs(1908) <= not b or a;
    outputs(1909) <= b;
    outputs(1910) <= a or b;
    outputs(1911) <= a xor b;
    outputs(1912) <= b;
    outputs(1913) <= b and not a;
    outputs(1914) <= a or b;
    outputs(1915) <= not a or b;
    outputs(1916) <= not b;
    outputs(1917) <= a or b;
    outputs(1918) <= a;
    outputs(1919) <= not b;
    outputs(1920) <= b and not a;
    outputs(1921) <= not b;
    outputs(1922) <= not a;
    outputs(1923) <= a and not b;
    outputs(1924) <= not a;
    outputs(1925) <= b;
    outputs(1926) <= not b;
    outputs(1927) <= not (a xor b);
    outputs(1928) <= a;
    outputs(1929) <= not (a or b);
    outputs(1930) <= a;
    outputs(1931) <= a and not b;
    outputs(1932) <= a xor b;
    outputs(1933) <= b and not a;
    outputs(1934) <= a and b;
    outputs(1935) <= a and not b;
    outputs(1936) <= not b or a;
    outputs(1937) <= b;
    outputs(1938) <= b;
    outputs(1939) <= not b or a;
    outputs(1940) <= a;
    outputs(1941) <= not a or b;
    outputs(1942) <= b;
    outputs(1943) <= not b;
    outputs(1944) <= not a or b;
    outputs(1945) <= b;
    outputs(1946) <= a and not b;
    outputs(1947) <= a xor b;
    outputs(1948) <= not a;
    outputs(1949) <= b;
    outputs(1950) <= not a;
    outputs(1951) <= a and not b;
    outputs(1952) <= b;
    outputs(1953) <= a;
    outputs(1954) <= not b;
    outputs(1955) <= b;
    outputs(1956) <= not b;
    outputs(1957) <= a;
    outputs(1958) <= not (a and b);
    outputs(1959) <= not a;
    outputs(1960) <= not a;
    outputs(1961) <= not b;
    outputs(1962) <= not a;
    outputs(1963) <= a xor b;
    outputs(1964) <= b and not a;
    outputs(1965) <= not (a xor b);
    outputs(1966) <= a;
    outputs(1967) <= b;
    outputs(1968) <= a xor b;
    outputs(1969) <= b;
    outputs(1970) <= a;
    outputs(1971) <= not a;
    outputs(1972) <= not (a or b);
    outputs(1973) <= not b;
    outputs(1974) <= not a;
    outputs(1975) <= not b;
    outputs(1976) <= not a;
    outputs(1977) <= not (a xor b);
    outputs(1978) <= not (a or b);
    outputs(1979) <= not b;
    outputs(1980) <= a;
    outputs(1981) <= not b or a;
    outputs(1982) <= not (a or b);
    outputs(1983) <= a;
    outputs(1984) <= a xor b;
    outputs(1985) <= a xor b;
    outputs(1986) <= not a or b;
    outputs(1987) <= a and not b;
    outputs(1988) <= a;
    outputs(1989) <= not (a xor b);
    outputs(1990) <= a;
    outputs(1991) <= not (a xor b);
    outputs(1992) <= a and b;
    outputs(1993) <= b;
    outputs(1994) <= b;
    outputs(1995) <= a or b;
    outputs(1996) <= not (a xor b);
    outputs(1997) <= not b;
    outputs(1998) <= a xor b;
    outputs(1999) <= a xor b;
    outputs(2000) <= not a;
    outputs(2001) <= not (a xor b);
    outputs(2002) <= not (a xor b);
    outputs(2003) <= a and b;
    outputs(2004) <= a xor b;
    outputs(2005) <= a xor b;
    outputs(2006) <= b;
    outputs(2007) <= not b;
    outputs(2008) <= not (a and b);
    outputs(2009) <= b;
    outputs(2010) <= b and not a;
    outputs(2011) <= not (a or b);
    outputs(2012) <= a or b;
    outputs(2013) <= a and not b;
    outputs(2014) <= a;
    outputs(2015) <= a xor b;
    outputs(2016) <= b and not a;
    outputs(2017) <= not (a or b);
    outputs(2018) <= not (a or b);
    outputs(2019) <= not a;
    outputs(2020) <= b;
    outputs(2021) <= not a;
    outputs(2022) <= not (a xor b);
    outputs(2023) <= not (a or b);
    outputs(2024) <= not (a xor b);
    outputs(2025) <= not (a or b);
    outputs(2026) <= not (a xor b);
    outputs(2027) <= not b;
    outputs(2028) <= b;
    outputs(2029) <= a and not b;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= not (a and b);
    outputs(2032) <= not a;
    outputs(2033) <= a and not b;
    outputs(2034) <= not (a and b);
    outputs(2035) <= not a;
    outputs(2036) <= a and b;
    outputs(2037) <= a xor b;
    outputs(2038) <= a xor b;
    outputs(2039) <= not a;
    outputs(2040) <= not (a xor b);
    outputs(2041) <= a xor b;
    outputs(2042) <= a and b;
    outputs(2043) <= b and not a;
    outputs(2044) <= b and not a;
    outputs(2045) <= not a;
    outputs(2046) <= not a;
    outputs(2047) <= not (a and b);
    outputs(2048) <= a xor b;
    outputs(2049) <= a and b;
    outputs(2050) <= b and not a;
    outputs(2051) <= not a;
    outputs(2052) <= not (a or b);
    outputs(2053) <= b and not a;
    outputs(2054) <= not (a xor b);
    outputs(2055) <= not b or a;
    outputs(2056) <= a xor b;
    outputs(2057) <= a or b;
    outputs(2058) <= not (a xor b);
    outputs(2059) <= not (a or b);
    outputs(2060) <= not a;
    outputs(2061) <= not b;
    outputs(2062) <= not a;
    outputs(2063) <= not a;
    outputs(2064) <= not b;
    outputs(2065) <= a;
    outputs(2066) <= not (a or b);
    outputs(2067) <= a or b;
    outputs(2068) <= not (a or b);
    outputs(2069) <= a;
    outputs(2070) <= not b;
    outputs(2071) <= b;
    outputs(2072) <= not b;
    outputs(2073) <= a xor b;
    outputs(2074) <= a;
    outputs(2075) <= not a or b;
    outputs(2076) <= not (a and b);
    outputs(2077) <= not b;
    outputs(2078) <= a xor b;
    outputs(2079) <= a xor b;
    outputs(2080) <= not b;
    outputs(2081) <= b;
    outputs(2082) <= not b;
    outputs(2083) <= a;
    outputs(2084) <= b;
    outputs(2085) <= a;
    outputs(2086) <= b;
    outputs(2087) <= not b or a;
    outputs(2088) <= not (a or b);
    outputs(2089) <= a and not b;
    outputs(2090) <= not b;
    outputs(2091) <= not a;
    outputs(2092) <= b and not a;
    outputs(2093) <= not (a xor b);
    outputs(2094) <= not (a or b);
    outputs(2095) <= a and b;
    outputs(2096) <= a;
    outputs(2097) <= b;
    outputs(2098) <= a and not b;
    outputs(2099) <= not b;
    outputs(2100) <= not a;
    outputs(2101) <= a and not b;
    outputs(2102) <= a xor b;
    outputs(2103) <= a xor b;
    outputs(2104) <= a xor b;
    outputs(2105) <= not (a or b);
    outputs(2106) <= not (a or b);
    outputs(2107) <= not (a xor b);
    outputs(2108) <= b;
    outputs(2109) <= not b;
    outputs(2110) <= a and not b;
    outputs(2111) <= b;
    outputs(2112) <= a and b;
    outputs(2113) <= a xor b;
    outputs(2114) <= not (a xor b);
    outputs(2115) <= not (a or b);
    outputs(2116) <= a and not b;
    outputs(2117) <= b;
    outputs(2118) <= a xor b;
    outputs(2119) <= not (a xor b);
    outputs(2120) <= a xor b;
    outputs(2121) <= not b;
    outputs(2122) <= not (a xor b);
    outputs(2123) <= b;
    outputs(2124) <= not (a xor b);
    outputs(2125) <= not (a or b);
    outputs(2126) <= a;
    outputs(2127) <= a;
    outputs(2128) <= a xor b;
    outputs(2129) <= not b;
    outputs(2130) <= not a;
    outputs(2131) <= b and not a;
    outputs(2132) <= a and not b;
    outputs(2133) <= b;
    outputs(2134) <= not a;
    outputs(2135) <= not a;
    outputs(2136) <= b;
    outputs(2137) <= not (a xor b);
    outputs(2138) <= b and not a;
    outputs(2139) <= a xor b;
    outputs(2140) <= not a;
    outputs(2141) <= a;
    outputs(2142) <= not b;
    outputs(2143) <= b;
    outputs(2144) <= not (a or b);
    outputs(2145) <= a and b;
    outputs(2146) <= b;
    outputs(2147) <= a;
    outputs(2148) <= b;
    outputs(2149) <= not (a and b);
    outputs(2150) <= not a;
    outputs(2151) <= a xor b;
    outputs(2152) <= a xor b;
    outputs(2153) <= a;
    outputs(2154) <= a and not b;
    outputs(2155) <= a or b;
    outputs(2156) <= not (a xor b);
    outputs(2157) <= b and not a;
    outputs(2158) <= not (a or b);
    outputs(2159) <= b;
    outputs(2160) <= a;
    outputs(2161) <= not a;
    outputs(2162) <= a;
    outputs(2163) <= b;
    outputs(2164) <= a or b;
    outputs(2165) <= not a or b;
    outputs(2166) <= a xor b;
    outputs(2167) <= not a;
    outputs(2168) <= not b or a;
    outputs(2169) <= b;
    outputs(2170) <= a and not b;
    outputs(2171) <= b;
    outputs(2172) <= not b or a;
    outputs(2173) <= not (a xor b);
    outputs(2174) <= a and not b;
    outputs(2175) <= a and b;
    outputs(2176) <= a xor b;
    outputs(2177) <= a xor b;
    outputs(2178) <= a;
    outputs(2179) <= a xor b;
    outputs(2180) <= not b;
    outputs(2181) <= not a;
    outputs(2182) <= a;
    outputs(2183) <= b;
    outputs(2184) <= a;
    outputs(2185) <= not (a xor b);
    outputs(2186) <= not (a xor b);
    outputs(2187) <= a;
    outputs(2188) <= a or b;
    outputs(2189) <= a xor b;
    outputs(2190) <= b;
    outputs(2191) <= a;
    outputs(2192) <= a;
    outputs(2193) <= not (a xor b);
    outputs(2194) <= b and not a;
    outputs(2195) <= not b;
    outputs(2196) <= not b;
    outputs(2197) <= not (a xor b);
    outputs(2198) <= b;
    outputs(2199) <= a;
    outputs(2200) <= not (a xor b);
    outputs(2201) <= not a or b;
    outputs(2202) <= a xor b;
    outputs(2203) <= a;
    outputs(2204) <= not (a xor b);
    outputs(2205) <= b;
    outputs(2206) <= not b;
    outputs(2207) <= not a;
    outputs(2208) <= not b;
    outputs(2209) <= not (a xor b);
    outputs(2210) <= not b;
    outputs(2211) <= not (a xor b);
    outputs(2212) <= not b;
    outputs(2213) <= not (a xor b);
    outputs(2214) <= b;
    outputs(2215) <= a and b;
    outputs(2216) <= not b;
    outputs(2217) <= not (a xor b);
    outputs(2218) <= a;
    outputs(2219) <= b;
    outputs(2220) <= a xor b;
    outputs(2221) <= a;
    outputs(2222) <= a;
    outputs(2223) <= not b;
    outputs(2224) <= b and not a;
    outputs(2225) <= not b or a;
    outputs(2226) <= b;
    outputs(2227) <= a xor b;
    outputs(2228) <= a and not b;
    outputs(2229) <= not (a xor b);
    outputs(2230) <= a;
    outputs(2231) <= a;
    outputs(2232) <= a xor b;
    outputs(2233) <= a or b;
    outputs(2234) <= b;
    outputs(2235) <= not (a and b);
    outputs(2236) <= a xor b;
    outputs(2237) <= not (a xor b);
    outputs(2238) <= not (a xor b);
    outputs(2239) <= b;
    outputs(2240) <= not a;
    outputs(2241) <= not b;
    outputs(2242) <= a xor b;
    outputs(2243) <= a;
    outputs(2244) <= b and not a;
    outputs(2245) <= not b;
    outputs(2246) <= a and b;
    outputs(2247) <= not b or a;
    outputs(2248) <= a xor b;
    outputs(2249) <= not a or b;
    outputs(2250) <= b;
    outputs(2251) <= b;
    outputs(2252) <= not (a xor b);
    outputs(2253) <= a and not b;
    outputs(2254) <= b;
    outputs(2255) <= not (a xor b);
    outputs(2256) <= a;
    outputs(2257) <= not (a or b);
    outputs(2258) <= b;
    outputs(2259) <= b;
    outputs(2260) <= not a;
    outputs(2261) <= a xor b;
    outputs(2262) <= not (a xor b);
    outputs(2263) <= not b;
    outputs(2264) <= not (a xor b);
    outputs(2265) <= not a;
    outputs(2266) <= a;
    outputs(2267) <= not (a or b);
    outputs(2268) <= not a;
    outputs(2269) <= not (a xor b);
    outputs(2270) <= not a;
    outputs(2271) <= not (a xor b);
    outputs(2272) <= not (a xor b);
    outputs(2273) <= not b;
    outputs(2274) <= not b;
    outputs(2275) <= a;
    outputs(2276) <= a;
    outputs(2277) <= not (a xor b);
    outputs(2278) <= a xor b;
    outputs(2279) <= a xor b;
    outputs(2280) <= a and not b;
    outputs(2281) <= b;
    outputs(2282) <= a;
    outputs(2283) <= a xor b;
    outputs(2284) <= a or b;
    outputs(2285) <= a xor b;
    outputs(2286) <= not b;
    outputs(2287) <= not b;
    outputs(2288) <= b and not a;
    outputs(2289) <= not b;
    outputs(2290) <= not a or b;
    outputs(2291) <= not (a or b);
    outputs(2292) <= a or b;
    outputs(2293) <= not a;
    outputs(2294) <= not a;
    outputs(2295) <= b and not a;
    outputs(2296) <= a xor b;
    outputs(2297) <= not (a xor b);
    outputs(2298) <= not (a xor b);
    outputs(2299) <= not (a xor b);
    outputs(2300) <= a or b;
    outputs(2301) <= a xor b;
    outputs(2302) <= b;
    outputs(2303) <= not (a xor b);
    outputs(2304) <= not b;
    outputs(2305) <= a and not b;
    outputs(2306) <= not (a xor b);
    outputs(2307) <= not (a xor b);
    outputs(2308) <= not (a xor b);
    outputs(2309) <= not b;
    outputs(2310) <= b;
    outputs(2311) <= a or b;
    outputs(2312) <= not b;
    outputs(2313) <= a xor b;
    outputs(2314) <= a;
    outputs(2315) <= a and not b;
    outputs(2316) <= a or b;
    outputs(2317) <= b;
    outputs(2318) <= b and not a;
    outputs(2319) <= b;
    outputs(2320) <= not b;
    outputs(2321) <= not a;
    outputs(2322) <= b;
    outputs(2323) <= b;
    outputs(2324) <= not b or a;
    outputs(2325) <= b;
    outputs(2326) <= a;
    outputs(2327) <= a;
    outputs(2328) <= a;
    outputs(2329) <= a xor b;
    outputs(2330) <= a and not b;
    outputs(2331) <= a and not b;
    outputs(2332) <= a or b;
    outputs(2333) <= a;
    outputs(2334) <= a xor b;
    outputs(2335) <= not (a or b);
    outputs(2336) <= not a;
    outputs(2337) <= not b;
    outputs(2338) <= not (a xor b);
    outputs(2339) <= a xor b;
    outputs(2340) <= not b or a;
    outputs(2341) <= b;
    outputs(2342) <= not (a xor b);
    outputs(2343) <= a;
    outputs(2344) <= not (a xor b);
    outputs(2345) <= a and b;
    outputs(2346) <= a and not b;
    outputs(2347) <= not (a xor b);
    outputs(2348) <= a and b;
    outputs(2349) <= not a;
    outputs(2350) <= a and not b;
    outputs(2351) <= a and not b;
    outputs(2352) <= not (a xor b);
    outputs(2353) <= not (a or b);
    outputs(2354) <= a;
    outputs(2355) <= a xor b;
    outputs(2356) <= not (a xor b);
    outputs(2357) <= b;
    outputs(2358) <= not b or a;
    outputs(2359) <= not (a xor b);
    outputs(2360) <= not (a xor b);
    outputs(2361) <= a and not b;
    outputs(2362) <= a or b;
    outputs(2363) <= not b;
    outputs(2364) <= not b;
    outputs(2365) <= a;
    outputs(2366) <= not (a or b);
    outputs(2367) <= not (a xor b);
    outputs(2368) <= b and not a;
    outputs(2369) <= b and not a;
    outputs(2370) <= not (a and b);
    outputs(2371) <= not a;
    outputs(2372) <= a and b;
    outputs(2373) <= not (a xor b);
    outputs(2374) <= b;
    outputs(2375) <= not (a xor b);
    outputs(2376) <= b;
    outputs(2377) <= not (a xor b);
    outputs(2378) <= a;
    outputs(2379) <= not (a xor b);
    outputs(2380) <= not (a or b);
    outputs(2381) <= b;
    outputs(2382) <= b;
    outputs(2383) <= b;
    outputs(2384) <= b;
    outputs(2385) <= a xor b;
    outputs(2386) <= a xor b;
    outputs(2387) <= a and b;
    outputs(2388) <= not (a or b);
    outputs(2389) <= not (a xor b);
    outputs(2390) <= not (a xor b);
    outputs(2391) <= a xor b;
    outputs(2392) <= not (a xor b);
    outputs(2393) <= not a;
    outputs(2394) <= b;
    outputs(2395) <= not a;
    outputs(2396) <= b;
    outputs(2397) <= a;
    outputs(2398) <= b;
    outputs(2399) <= b;
    outputs(2400) <= b;
    outputs(2401) <= not (a or b);
    outputs(2402) <= a and b;
    outputs(2403) <= a and not b;
    outputs(2404) <= not (a xor b);
    outputs(2405) <= not (a and b);
    outputs(2406) <= not (a or b);
    outputs(2407) <= not (a and b);
    outputs(2408) <= not b;
    outputs(2409) <= a or b;
    outputs(2410) <= not (a xor b);
    outputs(2411) <= a;
    outputs(2412) <= a and b;
    outputs(2413) <= a xor b;
    outputs(2414) <= not a;
    outputs(2415) <= a;
    outputs(2416) <= not (a xor b);
    outputs(2417) <= a xor b;
    outputs(2418) <= a;
    outputs(2419) <= b and not a;
    outputs(2420) <= a xor b;
    outputs(2421) <= a xor b;
    outputs(2422) <= a xor b;
    outputs(2423) <= b;
    outputs(2424) <= not (a and b);
    outputs(2425) <= not (a xor b);
    outputs(2426) <= a and not b;
    outputs(2427) <= not a;
    outputs(2428) <= not a;
    outputs(2429) <= a xor b;
    outputs(2430) <= not b;
    outputs(2431) <= a;
    outputs(2432) <= a;
    outputs(2433) <= b;
    outputs(2434) <= b;
    outputs(2435) <= not b;
    outputs(2436) <= not a;
    outputs(2437) <= not (a or b);
    outputs(2438) <= not (a xor b);
    outputs(2439) <= not a;
    outputs(2440) <= a;
    outputs(2441) <= not (a and b);
    outputs(2442) <= not (a or b);
    outputs(2443) <= not (a xor b);
    outputs(2444) <= b and not a;
    outputs(2445) <= not b;
    outputs(2446) <= not a;
    outputs(2447) <= b and not a;
    outputs(2448) <= a;
    outputs(2449) <= not b;
    outputs(2450) <= a and b;
    outputs(2451) <= b and not a;
    outputs(2452) <= b;
    outputs(2453) <= b;
    outputs(2454) <= b;
    outputs(2455) <= a or b;
    outputs(2456) <= a xor b;
    outputs(2457) <= not b;
    outputs(2458) <= a;
    outputs(2459) <= not a;
    outputs(2460) <= not (a xor b);
    outputs(2461) <= a or b;
    outputs(2462) <= not b;
    outputs(2463) <= a xor b;
    outputs(2464) <= not a;
    outputs(2465) <= a xor b;
    outputs(2466) <= a;
    outputs(2467) <= not (a xor b);
    outputs(2468) <= b;
    outputs(2469) <= not (a and b);
    outputs(2470) <= not a;
    outputs(2471) <= a;
    outputs(2472) <= b and not a;
    outputs(2473) <= not b;
    outputs(2474) <= a and b;
    outputs(2475) <= a;
    outputs(2476) <= not (a xor b);
    outputs(2477) <= not b;
    outputs(2478) <= not (a xor b);
    outputs(2479) <= b and not a;
    outputs(2480) <= not (a xor b);
    outputs(2481) <= a xor b;
    outputs(2482) <= a;
    outputs(2483) <= a;
    outputs(2484) <= not (a xor b);
    outputs(2485) <= not (a xor b);
    outputs(2486) <= not (a xor b);
    outputs(2487) <= a or b;
    outputs(2488) <= not a;
    outputs(2489) <= b;
    outputs(2490) <= not (a or b);
    outputs(2491) <= not (a xor b);
    outputs(2492) <= a;
    outputs(2493) <= not (a xor b);
    outputs(2494) <= not a or b;
    outputs(2495) <= not (a xor b);
    outputs(2496) <= not a;
    outputs(2497) <= not (a and b);
    outputs(2498) <= not (a or b);
    outputs(2499) <= not a;
    outputs(2500) <= b;
    outputs(2501) <= not b;
    outputs(2502) <= not a;
    outputs(2503) <= a;
    outputs(2504) <= b;
    outputs(2505) <= a xor b;
    outputs(2506) <= a or b;
    outputs(2507) <= b;
    outputs(2508) <= not (a or b);
    outputs(2509) <= b;
    outputs(2510) <= b;
    outputs(2511) <= not b;
    outputs(2512) <= a xor b;
    outputs(2513) <= not (a xor b);
    outputs(2514) <= not (a xor b);
    outputs(2515) <= a;
    outputs(2516) <= not a or b;
    outputs(2517) <= a xor b;
    outputs(2518) <= a xor b;
    outputs(2519) <= not b;
    outputs(2520) <= not b;
    outputs(2521) <= not b;
    outputs(2522) <= b;
    outputs(2523) <= b;
    outputs(2524) <= a xor b;
    outputs(2525) <= b;
    outputs(2526) <= not a;
    outputs(2527) <= not (a xor b);
    outputs(2528) <= a;
    outputs(2529) <= not b;
    outputs(2530) <= b and not a;
    outputs(2531) <= a and not b;
    outputs(2532) <= a and b;
    outputs(2533) <= not b;
    outputs(2534) <= not (a xor b);
    outputs(2535) <= not b;
    outputs(2536) <= a xor b;
    outputs(2537) <= a or b;
    outputs(2538) <= a;
    outputs(2539) <= a;
    outputs(2540) <= b;
    outputs(2541) <= a and b;
    outputs(2542) <= not (a and b);
    outputs(2543) <= not b;
    outputs(2544) <= not (a xor b);
    outputs(2545) <= a xor b;
    outputs(2546) <= a xor b;
    outputs(2547) <= a or b;
    outputs(2548) <= not (a xor b);
    outputs(2549) <= a;
    outputs(2550) <= not b;
    outputs(2551) <= b;
    outputs(2552) <= a xor b;
    outputs(2553) <= not (a or b);
    outputs(2554) <= not b or a;
    outputs(2555) <= a xor b;
    outputs(2556) <= not (a and b);
    outputs(2557) <= not b;
    outputs(2558) <= not a or b;
    outputs(2559) <= a;
    outputs(2560) <= not (a xor b);
    outputs(2561) <= not (a and b);
    outputs(2562) <= not (a or b);
    outputs(2563) <= a and not b;
    outputs(2564) <= not a;
    outputs(2565) <= not (a xor b);
    outputs(2566) <= a and b;
    outputs(2567) <= b and not a;
    outputs(2568) <= not b;
    outputs(2569) <= not (a xor b);
    outputs(2570) <= a xor b;
    outputs(2571) <= b;
    outputs(2572) <= a and b;
    outputs(2573) <= not a;
    outputs(2574) <= b and not a;
    outputs(2575) <= not a;
    outputs(2576) <= not a;
    outputs(2577) <= not a;
    outputs(2578) <= not (a xor b);
    outputs(2579) <= not a;
    outputs(2580) <= not b;
    outputs(2581) <= not (a xor b);
    outputs(2582) <= not a;
    outputs(2583) <= a;
    outputs(2584) <= a xor b;
    outputs(2585) <= not (a and b);
    outputs(2586) <= not (a xor b);
    outputs(2587) <= not b;
    outputs(2588) <= not (a xor b);
    outputs(2589) <= a;
    outputs(2590) <= b;
    outputs(2591) <= not (a or b);
    outputs(2592) <= not (a xor b);
    outputs(2593) <= b;
    outputs(2594) <= a xor b;
    outputs(2595) <= not a;
    outputs(2596) <= a;
    outputs(2597) <= b and not a;
    outputs(2598) <= not b or a;
    outputs(2599) <= not b;
    outputs(2600) <= a;
    outputs(2601) <= not a or b;
    outputs(2602) <= a xor b;
    outputs(2603) <= not b or a;
    outputs(2604) <= not (a and b);
    outputs(2605) <= a xor b;
    outputs(2606) <= not (a xor b);
    outputs(2607) <= not a;
    outputs(2608) <= a xor b;
    outputs(2609) <= a xor b;
    outputs(2610) <= not (a xor b);
    outputs(2611) <= not b;
    outputs(2612) <= not (a xor b);
    outputs(2613) <= a or b;
    outputs(2614) <= not a;
    outputs(2615) <= a and not b;
    outputs(2616) <= not b;
    outputs(2617) <= not (a xor b);
    outputs(2618) <= not a or b;
    outputs(2619) <= b;
    outputs(2620) <= not (a or b);
    outputs(2621) <= not (a xor b);
    outputs(2622) <= not a;
    outputs(2623) <= a xor b;
    outputs(2624) <= a;
    outputs(2625) <= b;
    outputs(2626) <= a xor b;
    outputs(2627) <= not b;
    outputs(2628) <= not a;
    outputs(2629) <= b;
    outputs(2630) <= a and b;
    outputs(2631) <= not (a xor b);
    outputs(2632) <= not (a xor b);
    outputs(2633) <= a;
    outputs(2634) <= not (a xor b);
    outputs(2635) <= b;
    outputs(2636) <= b and not a;
    outputs(2637) <= a and b;
    outputs(2638) <= a;
    outputs(2639) <= a and not b;
    outputs(2640) <= a and not b;
    outputs(2641) <= not (a or b);
    outputs(2642) <= a;
    outputs(2643) <= not (a and b);
    outputs(2644) <= a xor b;
    outputs(2645) <= a xor b;
    outputs(2646) <= a xor b;
    outputs(2647) <= not b;
    outputs(2648) <= a xor b;
    outputs(2649) <= b;
    outputs(2650) <= a or b;
    outputs(2651) <= a or b;
    outputs(2652) <= a and not b;
    outputs(2653) <= a;
    outputs(2654) <= not (a xor b);
    outputs(2655) <= not (a xor b);
    outputs(2656) <= not b;
    outputs(2657) <= b;
    outputs(2658) <= a xor b;
    outputs(2659) <= a xor b;
    outputs(2660) <= not b;
    outputs(2661) <= not b;
    outputs(2662) <= not a;
    outputs(2663) <= a;
    outputs(2664) <= b and not a;
    outputs(2665) <= not b;
    outputs(2666) <= not (a xor b);
    outputs(2667) <= not (a xor b);
    outputs(2668) <= not b;
    outputs(2669) <= not (a or b);
    outputs(2670) <= b and not a;
    outputs(2671) <= not (a xor b);
    outputs(2672) <= a and b;
    outputs(2673) <= not (a or b);
    outputs(2674) <= b;
    outputs(2675) <= not (a xor b);
    outputs(2676) <= not a;
    outputs(2677) <= a;
    outputs(2678) <= b;
    outputs(2679) <= a xor b;
    outputs(2680) <= a;
    outputs(2681) <= a;
    outputs(2682) <= a and not b;
    outputs(2683) <= b;
    outputs(2684) <= not b or a;
    outputs(2685) <= not (a xor b);
    outputs(2686) <= a xor b;
    outputs(2687) <= a and b;
    outputs(2688) <= not (a and b);
    outputs(2689) <= not b;
    outputs(2690) <= not (a xor b);
    outputs(2691) <= not a;
    outputs(2692) <= not b;
    outputs(2693) <= not a;
    outputs(2694) <= a or b;
    outputs(2695) <= not (a and b);
    outputs(2696) <= b;
    outputs(2697) <= a or b;
    outputs(2698) <= not b;
    outputs(2699) <= a xor b;
    outputs(2700) <= a;
    outputs(2701) <= not (a xor b);
    outputs(2702) <= a xor b;
    outputs(2703) <= not a;
    outputs(2704) <= not (a xor b);
    outputs(2705) <= not (a or b);
    outputs(2706) <= not (a or b);
    outputs(2707) <= not a;
    outputs(2708) <= a;
    outputs(2709) <= b;
    outputs(2710) <= a xor b;
    outputs(2711) <= b;
    outputs(2712) <= b and not a;
    outputs(2713) <= a xor b;
    outputs(2714) <= not b;
    outputs(2715) <= not a;
    outputs(2716) <= a and b;
    outputs(2717) <= a and not b;
    outputs(2718) <= b;
    outputs(2719) <= b;
    outputs(2720) <= not a;
    outputs(2721) <= a xor b;
    outputs(2722) <= a;
    outputs(2723) <= a or b;
    outputs(2724) <= a xor b;
    outputs(2725) <= a and not b;
    outputs(2726) <= not b or a;
    outputs(2727) <= a or b;
    outputs(2728) <= a;
    outputs(2729) <= a xor b;
    outputs(2730) <= not b;
    outputs(2731) <= not b;
    outputs(2732) <= not b;
    outputs(2733) <= not a;
    outputs(2734) <= b;
    outputs(2735) <= a;
    outputs(2736) <= not a;
    outputs(2737) <= b and not a;
    outputs(2738) <= not (a xor b);
    outputs(2739) <= b and not a;
    outputs(2740) <= a xor b;
    outputs(2741) <= a xor b;
    outputs(2742) <= not b;
    outputs(2743) <= a or b;
    outputs(2744) <= b and not a;
    outputs(2745) <= not a;
    outputs(2746) <= b;
    outputs(2747) <= b and not a;
    outputs(2748) <= not b;
    outputs(2749) <= not a;
    outputs(2750) <= not (a xor b);
    outputs(2751) <= not b;
    outputs(2752) <= a;
    outputs(2753) <= a;
    outputs(2754) <= not b;
    outputs(2755) <= not a;
    outputs(2756) <= not (a xor b);
    outputs(2757) <= a;
    outputs(2758) <= a;
    outputs(2759) <= a xor b;
    outputs(2760) <= b and not a;
    outputs(2761) <= not (a xor b);
    outputs(2762) <= not a or b;
    outputs(2763) <= a or b;
    outputs(2764) <= b;
    outputs(2765) <= a and b;
    outputs(2766) <= b;
    outputs(2767) <= not (a or b);
    outputs(2768) <= not a;
    outputs(2769) <= not b;
    outputs(2770) <= not a;
    outputs(2771) <= a or b;
    outputs(2772) <= a and not b;
    outputs(2773) <= not (a or b);
    outputs(2774) <= not b;
    outputs(2775) <= not a;
    outputs(2776) <= not (a xor b);
    outputs(2777) <= not (a xor b);
    outputs(2778) <= b and not a;
    outputs(2779) <= not b;
    outputs(2780) <= not (a xor b);
    outputs(2781) <= not a;
    outputs(2782) <= b and not a;
    outputs(2783) <= not (a and b);
    outputs(2784) <= a xor b;
    outputs(2785) <= not b;
    outputs(2786) <= b and not a;
    outputs(2787) <= a;
    outputs(2788) <= a;
    outputs(2789) <= not a;
    outputs(2790) <= not b;
    outputs(2791) <= a xor b;
    outputs(2792) <= a or b;
    outputs(2793) <= a xor b;
    outputs(2794) <= a xor b;
    outputs(2795) <= a and not b;
    outputs(2796) <= b;
    outputs(2797) <= not b;
    outputs(2798) <= not a;
    outputs(2799) <= a;
    outputs(2800) <= a xor b;
    outputs(2801) <= a xor b;
    outputs(2802) <= not b;
    outputs(2803) <= a;
    outputs(2804) <= a;
    outputs(2805) <= a or b;
    outputs(2806) <= not (a xor b);
    outputs(2807) <= not (a or b);
    outputs(2808) <= b;
    outputs(2809) <= not (a xor b);
    outputs(2810) <= a xor b;
    outputs(2811) <= a;
    outputs(2812) <= a and not b;
    outputs(2813) <= b;
    outputs(2814) <= a xor b;
    outputs(2815) <= a xor b;
    outputs(2816) <= not b;
    outputs(2817) <= a and b;
    outputs(2818) <= not (a or b);
    outputs(2819) <= b;
    outputs(2820) <= not a;
    outputs(2821) <= not a or b;
    outputs(2822) <= not a;
    outputs(2823) <= a;
    outputs(2824) <= b and not a;
    outputs(2825) <= not (a and b);
    outputs(2826) <= not b;
    outputs(2827) <= a;
    outputs(2828) <= a xor b;
    outputs(2829) <= a;
    outputs(2830) <= not (a or b);
    outputs(2831) <= not (a xor b);
    outputs(2832) <= a xor b;
    outputs(2833) <= b;
    outputs(2834) <= a xor b;
    outputs(2835) <= not (a and b);
    outputs(2836) <= a and not b;
    outputs(2837) <= a xor b;
    outputs(2838) <= a and b;
    outputs(2839) <= a xor b;
    outputs(2840) <= a xor b;
    outputs(2841) <= not (a xor b);
    outputs(2842) <= not a;
    outputs(2843) <= a xor b;
    outputs(2844) <= a xor b;
    outputs(2845) <= b and not a;
    outputs(2846) <= b;
    outputs(2847) <= not b;
    outputs(2848) <= b and not a;
    outputs(2849) <= not (a or b);
    outputs(2850) <= not b;
    outputs(2851) <= b;
    outputs(2852) <= b;
    outputs(2853) <= not (a xor b);
    outputs(2854) <= b;
    outputs(2855) <= not b;
    outputs(2856) <= not (a xor b);
    outputs(2857) <= b;
    outputs(2858) <= a;
    outputs(2859) <= not a;
    outputs(2860) <= not a;
    outputs(2861) <= not (a xor b);
    outputs(2862) <= b;
    outputs(2863) <= not b;
    outputs(2864) <= a xor b;
    outputs(2865) <= not a;
    outputs(2866) <= not b;
    outputs(2867) <= b and not a;
    outputs(2868) <= not (a xor b);
    outputs(2869) <= not b;
    outputs(2870) <= not a;
    outputs(2871) <= not b or a;
    outputs(2872) <= not b;
    outputs(2873) <= not (a xor b);
    outputs(2874) <= not (a or b);
    outputs(2875) <= not b;
    outputs(2876) <= a xor b;
    outputs(2877) <= b;
    outputs(2878) <= not b or a;
    outputs(2879) <= not b;
    outputs(2880) <= a;
    outputs(2881) <= not (a xor b);
    outputs(2882) <= not (a xor b);
    outputs(2883) <= not b or a;
    outputs(2884) <= not a;
    outputs(2885) <= a and not b;
    outputs(2886) <= a;
    outputs(2887) <= b and not a;
    outputs(2888) <= a and not b;
    outputs(2889) <= not b;
    outputs(2890) <= a;
    outputs(2891) <= a and b;
    outputs(2892) <= a xor b;
    outputs(2893) <= a xor b;
    outputs(2894) <= not (a or b);
    outputs(2895) <= not a;
    outputs(2896) <= a;
    outputs(2897) <= not a or b;
    outputs(2898) <= a and b;
    outputs(2899) <= not a;
    outputs(2900) <= not (a and b);
    outputs(2901) <= b;
    outputs(2902) <= not (a xor b);
    outputs(2903) <= not a;
    outputs(2904) <= not (a or b);
    outputs(2905) <= a xor b;
    outputs(2906) <= not (a and b);
    outputs(2907) <= a;
    outputs(2908) <= not (a and b);
    outputs(2909) <= b and not a;
    outputs(2910) <= a and b;
    outputs(2911) <= not b or a;
    outputs(2912) <= not (a xor b);
    outputs(2913) <= not a;
    outputs(2914) <= not b;
    outputs(2915) <= a;
    outputs(2916) <= not (a or b);
    outputs(2917) <= a and b;
    outputs(2918) <= not (a or b);
    outputs(2919) <= a xor b;
    outputs(2920) <= not (a xor b);
    outputs(2921) <= a xor b;
    outputs(2922) <= b and not a;
    outputs(2923) <= a and not b;
    outputs(2924) <= b;
    outputs(2925) <= a xor b;
    outputs(2926) <= b;
    outputs(2927) <= a and not b;
    outputs(2928) <= not a;
    outputs(2929) <= not (a xor b);
    outputs(2930) <= a and not b;
    outputs(2931) <= not b;
    outputs(2932) <= a;
    outputs(2933) <= not (a or b);
    outputs(2934) <= a xor b;
    outputs(2935) <= not b;
    outputs(2936) <= a xor b;
    outputs(2937) <= a;
    outputs(2938) <= b;
    outputs(2939) <= a;
    outputs(2940) <= not b;
    outputs(2941) <= not b;
    outputs(2942) <= not (a and b);
    outputs(2943) <= not b;
    outputs(2944) <= a xor b;
    outputs(2945) <= not (a or b);
    outputs(2946) <= not (a xor b);
    outputs(2947) <= b;
    outputs(2948) <= a xor b;
    outputs(2949) <= b;
    outputs(2950) <= not (a xor b);
    outputs(2951) <= not (a or b);
    outputs(2952) <= a;
    outputs(2953) <= a;
    outputs(2954) <= not b;
    outputs(2955) <= not (a xor b);
    outputs(2956) <= not (a xor b);
    outputs(2957) <= not (a or b);
    outputs(2958) <= b;
    outputs(2959) <= not (a xor b);
    outputs(2960) <= b;
    outputs(2961) <= a;
    outputs(2962) <= not a or b;
    outputs(2963) <= b;
    outputs(2964) <= not (a or b);
    outputs(2965) <= not (a xor b);
    outputs(2966) <= a;
    outputs(2967) <= not a;
    outputs(2968) <= not a;
    outputs(2969) <= a or b;
    outputs(2970) <= not (a xor b);
    outputs(2971) <= a xor b;
    outputs(2972) <= a xor b;
    outputs(2973) <= b;
    outputs(2974) <= a xor b;
    outputs(2975) <= a xor b;
    outputs(2976) <= not (a xor b);
    outputs(2977) <= a xor b;
    outputs(2978) <= not (a and b);
    outputs(2979) <= b;
    outputs(2980) <= a xor b;
    outputs(2981) <= b and not a;
    outputs(2982) <= a xor b;
    outputs(2983) <= b;
    outputs(2984) <= not (a xor b);
    outputs(2985) <= not (a and b);
    outputs(2986) <= not (a and b);
    outputs(2987) <= a;
    outputs(2988) <= b;
    outputs(2989) <= not b;
    outputs(2990) <= not a;
    outputs(2991) <= a;
    outputs(2992) <= b;
    outputs(2993) <= a and b;
    outputs(2994) <= a and not b;
    outputs(2995) <= b and not a;
    outputs(2996) <= not (a xor b);
    outputs(2997) <= not a or b;
    outputs(2998) <= not a;
    outputs(2999) <= not a;
    outputs(3000) <= b;
    outputs(3001) <= a;
    outputs(3002) <= a;
    outputs(3003) <= not b;
    outputs(3004) <= a;
    outputs(3005) <= not b;
    outputs(3006) <= not (a or b);
    outputs(3007) <= not (a xor b);
    outputs(3008) <= a;
    outputs(3009) <= not (a xor b);
    outputs(3010) <= not b;
    outputs(3011) <= not a;
    outputs(3012) <= a xor b;
    outputs(3013) <= a xor b;
    outputs(3014) <= not b;
    outputs(3015) <= not (a xor b);
    outputs(3016) <= a;
    outputs(3017) <= a;
    outputs(3018) <= not b;
    outputs(3019) <= not a;
    outputs(3020) <= a xor b;
    outputs(3021) <= a;
    outputs(3022) <= a;
    outputs(3023) <= a xor b;
    outputs(3024) <= a;
    outputs(3025) <= not a;
    outputs(3026) <= a;
    outputs(3027) <= not a;
    outputs(3028) <= b and not a;
    outputs(3029) <= not a or b;
    outputs(3030) <= b;
    outputs(3031) <= not (a or b);
    outputs(3032) <= not a;
    outputs(3033) <= not a;
    outputs(3034) <= a;
    outputs(3035) <= a xor b;
    outputs(3036) <= a;
    outputs(3037) <= not (a xor b);
    outputs(3038) <= not b or a;
    outputs(3039) <= a xor b;
    outputs(3040) <= b and not a;
    outputs(3041) <= b;
    outputs(3042) <= not b;
    outputs(3043) <= a and not b;
    outputs(3044) <= a xor b;
    outputs(3045) <= a xor b;
    outputs(3046) <= b;
    outputs(3047) <= a and b;
    outputs(3048) <= a xor b;
    outputs(3049) <= a;
    outputs(3050) <= not (a xor b);
    outputs(3051) <= b and not a;
    outputs(3052) <= not a;
    outputs(3053) <= a xor b;
    outputs(3054) <= not (a xor b);
    outputs(3055) <= not (a xor b);
    outputs(3056) <= a;
    outputs(3057) <= a or b;
    outputs(3058) <= a xor b;
    outputs(3059) <= a;
    outputs(3060) <= b and not a;
    outputs(3061) <= a and b;
    outputs(3062) <= not a;
    outputs(3063) <= not b or a;
    outputs(3064) <= b and not a;
    outputs(3065) <= not (a xor b);
    outputs(3066) <= not b;
    outputs(3067) <= a xor b;
    outputs(3068) <= a xor b;
    outputs(3069) <= not b;
    outputs(3070) <= b;
    outputs(3071) <= not b;
    outputs(3072) <= not (a xor b);
    outputs(3073) <= not b;
    outputs(3074) <= a;
    outputs(3075) <= not (a and b);
    outputs(3076) <= a;
    outputs(3077) <= not b or a;
    outputs(3078) <= not b;
    outputs(3079) <= not (a or b);
    outputs(3080) <= not b;
    outputs(3081) <= not a;
    outputs(3082) <= a and b;
    outputs(3083) <= not (a xor b);
    outputs(3084) <= a;
    outputs(3085) <= not (a and b);
    outputs(3086) <= not b;
    outputs(3087) <= a and not b;
    outputs(3088) <= a and b;
    outputs(3089) <= not b or a;
    outputs(3090) <= a xor b;
    outputs(3091) <= not (a xor b);
    outputs(3092) <= not b;
    outputs(3093) <= b;
    outputs(3094) <= b and not a;
    outputs(3095) <= not a;
    outputs(3096) <= a;
    outputs(3097) <= a xor b;
    outputs(3098) <= a or b;
    outputs(3099) <= not a or b;
    outputs(3100) <= not a;
    outputs(3101) <= not a;
    outputs(3102) <= a xor b;
    outputs(3103) <= not (a xor b);
    outputs(3104) <= not a or b;
    outputs(3105) <= a and b;
    outputs(3106) <= b and not a;
    outputs(3107) <= b;
    outputs(3108) <= not a;
    outputs(3109) <= not (a xor b);
    outputs(3110) <= a;
    outputs(3111) <= a;
    outputs(3112) <= not a;
    outputs(3113) <= a xor b;
    outputs(3114) <= not b;
    outputs(3115) <= not (a xor b);
    outputs(3116) <= a xor b;
    outputs(3117) <= not (a xor b);
    outputs(3118) <= not b;
    outputs(3119) <= a;
    outputs(3120) <= b;
    outputs(3121) <= not (a and b);
    outputs(3122) <= not b;
    outputs(3123) <= not (a xor b);
    outputs(3124) <= not b;
    outputs(3125) <= b and not a;
    outputs(3126) <= a and b;
    outputs(3127) <= not (a xor b);
    outputs(3128) <= a and not b;
    outputs(3129) <= not a;
    outputs(3130) <= a xor b;
    outputs(3131) <= not (a and b);
    outputs(3132) <= not (a xor b);
    outputs(3133) <= not b;
    outputs(3134) <= a and not b;
    outputs(3135) <= a and b;
    outputs(3136) <= b;
    outputs(3137) <= not b;
    outputs(3138) <= not (a xor b);
    outputs(3139) <= not b;
    outputs(3140) <= not (a xor b);
    outputs(3141) <= a xor b;
    outputs(3142) <= not a;
    outputs(3143) <= not b;
    outputs(3144) <= a;
    outputs(3145) <= a xor b;
    outputs(3146) <= not a;
    outputs(3147) <= not b;
    outputs(3148) <= not b;
    outputs(3149) <= b;
    outputs(3150) <= a;
    outputs(3151) <= not (a or b);
    outputs(3152) <= a and not b;
    outputs(3153) <= b;
    outputs(3154) <= b;
    outputs(3155) <= a xor b;
    outputs(3156) <= not a;
    outputs(3157) <= a xor b;
    outputs(3158) <= not b;
    outputs(3159) <= a and b;
    outputs(3160) <= b;
    outputs(3161) <= not b or a;
    outputs(3162) <= not a;
    outputs(3163) <= not a or b;
    outputs(3164) <= b;
    outputs(3165) <= not (a or b);
    outputs(3166) <= b;
    outputs(3167) <= not (a xor b);
    outputs(3168) <= not b;
    outputs(3169) <= not (a xor b);
    outputs(3170) <= b and not a;
    outputs(3171) <= b;
    outputs(3172) <= not a or b;
    outputs(3173) <= a xor b;
    outputs(3174) <= a xor b;
    outputs(3175) <= a or b;
    outputs(3176) <= not (a xor b);
    outputs(3177) <= not (a and b);
    outputs(3178) <= a;
    outputs(3179) <= not b;
    outputs(3180) <= not (a xor b);
    outputs(3181) <= not (a or b);
    outputs(3182) <= a xor b;
    outputs(3183) <= b;
    outputs(3184) <= not a;
    outputs(3185) <= not a;
    outputs(3186) <= not a;
    outputs(3187) <= b and not a;
    outputs(3188) <= not b;
    outputs(3189) <= not (a xor b);
    outputs(3190) <= not a;
    outputs(3191) <= not b or a;
    outputs(3192) <= a;
    outputs(3193) <= not (a and b);
    outputs(3194) <= a;
    outputs(3195) <= a xor b;
    outputs(3196) <= not a;
    outputs(3197) <= not (a xor b);
    outputs(3198) <= not (a xor b);
    outputs(3199) <= a;
    outputs(3200) <= b and not a;
    outputs(3201) <= a;
    outputs(3202) <= a xor b;
    outputs(3203) <= a and not b;
    outputs(3204) <= a;
    outputs(3205) <= not a;
    outputs(3206) <= not (a or b);
    outputs(3207) <= a;
    outputs(3208) <= not (a xor b);
    outputs(3209) <= not b;
    outputs(3210) <= not (a xor b);
    outputs(3211) <= not b or a;
    outputs(3212) <= not (a xor b);
    outputs(3213) <= not b or a;
    outputs(3214) <= not a;
    outputs(3215) <= a xor b;
    outputs(3216) <= not b;
    outputs(3217) <= not b;
    outputs(3218) <= not b;
    outputs(3219) <= a;
    outputs(3220) <= a;
    outputs(3221) <= a xor b;
    outputs(3222) <= a;
    outputs(3223) <= a;
    outputs(3224) <= b;
    outputs(3225) <= not (a and b);
    outputs(3226) <= a and b;
    outputs(3227) <= not (a xor b);
    outputs(3228) <= a or b;
    outputs(3229) <= a xor b;
    outputs(3230) <= b;
    outputs(3231) <= not (a xor b);
    outputs(3232) <= not a;
    outputs(3233) <= a xor b;
    outputs(3234) <= not (a xor b);
    outputs(3235) <= not (a xor b);
    outputs(3236) <= not (a xor b);
    outputs(3237) <= not b;
    outputs(3238) <= not (a or b);
    outputs(3239) <= b and not a;
    outputs(3240) <= not (a xor b);
    outputs(3241) <= not a;
    outputs(3242) <= a xor b;
    outputs(3243) <= not (a xor b);
    outputs(3244) <= not (a and b);
    outputs(3245) <= a or b;
    outputs(3246) <= a;
    outputs(3247) <= b;
    outputs(3248) <= b and not a;
    outputs(3249) <= a xor b;
    outputs(3250) <= b;
    outputs(3251) <= not (a xor b);
    outputs(3252) <= a;
    outputs(3253) <= a xor b;
    outputs(3254) <= not a;
    outputs(3255) <= not a;
    outputs(3256) <= a;
    outputs(3257) <= a and b;
    outputs(3258) <= not a;
    outputs(3259) <= not b;
    outputs(3260) <= a;
    outputs(3261) <= not a or b;
    outputs(3262) <= a xor b;
    outputs(3263) <= not (a or b);
    outputs(3264) <= b;
    outputs(3265) <= a and not b;
    outputs(3266) <= not a;
    outputs(3267) <= not a;
    outputs(3268) <= b and not a;
    outputs(3269) <= not a;
    outputs(3270) <= b;
    outputs(3271) <= a and not b;
    outputs(3272) <= b;
    outputs(3273) <= not b;
    outputs(3274) <= a and not b;
    outputs(3275) <= a or b;
    outputs(3276) <= a and b;
    outputs(3277) <= a;
    outputs(3278) <= not a or b;
    outputs(3279) <= b and not a;
    outputs(3280) <= a xor b;
    outputs(3281) <= not a;
    outputs(3282) <= not (a xor b);
    outputs(3283) <= a;
    outputs(3284) <= b and not a;
    outputs(3285) <= a;
    outputs(3286) <= a and not b;
    outputs(3287) <= not a;
    outputs(3288) <= not b;
    outputs(3289) <= a or b;
    outputs(3290) <= b and not a;
    outputs(3291) <= b and not a;
    outputs(3292) <= not (a xor b);
    outputs(3293) <= not b;
    outputs(3294) <= a;
    outputs(3295) <= b;
    outputs(3296) <= a and b;
    outputs(3297) <= b;
    outputs(3298) <= not (a xor b);
    outputs(3299) <= not b;
    outputs(3300) <= a;
    outputs(3301) <= a xor b;
    outputs(3302) <= a xor b;
    outputs(3303) <= not (a xor b);
    outputs(3304) <= not (a xor b);
    outputs(3305) <= a;
    outputs(3306) <= b;
    outputs(3307) <= b;
    outputs(3308) <= not b;
    outputs(3309) <= not (a xor b);
    outputs(3310) <= b;
    outputs(3311) <= b;
    outputs(3312) <= not b or a;
    outputs(3313) <= a;
    outputs(3314) <= not (a or b);
    outputs(3315) <= not (a or b);
    outputs(3316) <= not b;
    outputs(3317) <= a;
    outputs(3318) <= not (a and b);
    outputs(3319) <= not b;
    outputs(3320) <= b;
    outputs(3321) <= not b;
    outputs(3322) <= not b or a;
    outputs(3323) <= not b;
    outputs(3324) <= b;
    outputs(3325) <= not b;
    outputs(3326) <= not (a or b);
    outputs(3327) <= not a;
    outputs(3328) <= a and not b;
    outputs(3329) <= not (a xor b);
    outputs(3330) <= not (a and b);
    outputs(3331) <= not (a or b);
    outputs(3332) <= not (a or b);
    outputs(3333) <= not (a xor b);
    outputs(3334) <= a;
    outputs(3335) <= not a;
    outputs(3336) <= a and not b;
    outputs(3337) <= not a;
    outputs(3338) <= not a or b;
    outputs(3339) <= not a;
    outputs(3340) <= not a;
    outputs(3341) <= a;
    outputs(3342) <= b;
    outputs(3343) <= not a;
    outputs(3344) <= a xor b;
    outputs(3345) <= not (a xor b);
    outputs(3346) <= not b;
    outputs(3347) <= not (a xor b);
    outputs(3348) <= a and b;
    outputs(3349) <= a xor b;
    outputs(3350) <= a;
    outputs(3351) <= not (a and b);
    outputs(3352) <= not a;
    outputs(3353) <= b;
    outputs(3354) <= b;
    outputs(3355) <= not b;
    outputs(3356) <= not (a or b);
    outputs(3357) <= a and b;
    outputs(3358) <= a and not b;
    outputs(3359) <= not a;
    outputs(3360) <= b;
    outputs(3361) <= not a or b;
    outputs(3362) <= a and b;
    outputs(3363) <= not (a xor b);
    outputs(3364) <= a;
    outputs(3365) <= a;
    outputs(3366) <= not (a xor b);
    outputs(3367) <= a xor b;
    outputs(3368) <= a xor b;
    outputs(3369) <= b;
    outputs(3370) <= not (a or b);
    outputs(3371) <= not (a xor b);
    outputs(3372) <= not b or a;
    outputs(3373) <= not b;
    outputs(3374) <= a and b;
    outputs(3375) <= not (a xor b);
    outputs(3376) <= not b;
    outputs(3377) <= a;
    outputs(3378) <= b;
    outputs(3379) <= not b;
    outputs(3380) <= b;
    outputs(3381) <= not b;
    outputs(3382) <= a;
    outputs(3383) <= not a;
    outputs(3384) <= a;
    outputs(3385) <= a and not b;
    outputs(3386) <= a xor b;
    outputs(3387) <= b;
    outputs(3388) <= not b;
    outputs(3389) <= a or b;
    outputs(3390) <= a;
    outputs(3391) <= not b;
    outputs(3392) <= a and not b;
    outputs(3393) <= a xor b;
    outputs(3394) <= a;
    outputs(3395) <= a and b;
    outputs(3396) <= not (a xor b);
    outputs(3397) <= not b;
    outputs(3398) <= not a;
    outputs(3399) <= a;
    outputs(3400) <= not a;
    outputs(3401) <= not a;
    outputs(3402) <= not b;
    outputs(3403) <= not a;
    outputs(3404) <= a xor b;
    outputs(3405) <= not a or b;
    outputs(3406) <= not b;
    outputs(3407) <= b;
    outputs(3408) <= a;
    outputs(3409) <= a;
    outputs(3410) <= a xor b;
    outputs(3411) <= not b;
    outputs(3412) <= not b;
    outputs(3413) <= not (a xor b);
    outputs(3414) <= not (a and b);
    outputs(3415) <= a and not b;
    outputs(3416) <= a and b;
    outputs(3417) <= not a;
    outputs(3418) <= not (a or b);
    outputs(3419) <= not b;
    outputs(3420) <= a xor b;
    outputs(3421) <= not (a xor b);
    outputs(3422) <= a;
    outputs(3423) <= a;
    outputs(3424) <= not (a xor b);
    outputs(3425) <= not a;
    outputs(3426) <= a;
    outputs(3427) <= a and not b;
    outputs(3428) <= not b;
    outputs(3429) <= a;
    outputs(3430) <= b;
    outputs(3431) <= not (a xor b);
    outputs(3432) <= a and b;
    outputs(3433) <= b;
    outputs(3434) <= a;
    outputs(3435) <= not (a xor b);
    outputs(3436) <= not (a xor b);
    outputs(3437) <= a;
    outputs(3438) <= not a;
    outputs(3439) <= a xor b;
    outputs(3440) <= a xor b;
    outputs(3441) <= b;
    outputs(3442) <= a xor b;
    outputs(3443) <= not (a and b);
    outputs(3444) <= a or b;
    outputs(3445) <= not b;
    outputs(3446) <= not (a xor b);
    outputs(3447) <= not b;
    outputs(3448) <= not (a xor b);
    outputs(3449) <= a;
    outputs(3450) <= not b;
    outputs(3451) <= b;
    outputs(3452) <= not b;
    outputs(3453) <= not (a xor b);
    outputs(3454) <= a and not b;
    outputs(3455) <= not (a or b);
    outputs(3456) <= a;
    outputs(3457) <= not b or a;
    outputs(3458) <= not b;
    outputs(3459) <= not a;
    outputs(3460) <= a and b;
    outputs(3461) <= not b;
    outputs(3462) <= not a;
    outputs(3463) <= not (a xor b);
    outputs(3464) <= a;
    outputs(3465) <= a;
    outputs(3466) <= not b or a;
    outputs(3467) <= a;
    outputs(3468) <= b;
    outputs(3469) <= not b;
    outputs(3470) <= not b;
    outputs(3471) <= a xor b;
    outputs(3472) <= a;
    outputs(3473) <= a and b;
    outputs(3474) <= a xor b;
    outputs(3475) <= not a;
    outputs(3476) <= not b;
    outputs(3477) <= b;
    outputs(3478) <= a and not b;
    outputs(3479) <= a xor b;
    outputs(3480) <= b;
    outputs(3481) <= not a;
    outputs(3482) <= not a;
    outputs(3483) <= not (a or b);
    outputs(3484) <= a xor b;
    outputs(3485) <= not (a xor b);
    outputs(3486) <= a and b;
    outputs(3487) <= not b;
    outputs(3488) <= not (a xor b);
    outputs(3489) <= a and b;
    outputs(3490) <= not (a xor b);
    outputs(3491) <= not a;
    outputs(3492) <= a and b;
    outputs(3493) <= a xor b;
    outputs(3494) <= not b or a;
    outputs(3495) <= a and not b;
    outputs(3496) <= a or b;
    outputs(3497) <= not b;
    outputs(3498) <= not a;
    outputs(3499) <= not (a xor b);
    outputs(3500) <= a;
    outputs(3501) <= not (a xor b);
    outputs(3502) <= b;
    outputs(3503) <= a and b;
    outputs(3504) <= a;
    outputs(3505) <= not b;
    outputs(3506) <= not b;
    outputs(3507) <= a xor b;
    outputs(3508) <= not a or b;
    outputs(3509) <= not a;
    outputs(3510) <= not (a xor b);
    outputs(3511) <= not b;
    outputs(3512) <= not (a or b);
    outputs(3513) <= not (a or b);
    outputs(3514) <= a;
    outputs(3515) <= a xor b;
    outputs(3516) <= not b;
    outputs(3517) <= b;
    outputs(3518) <= not (a or b);
    outputs(3519) <= not b;
    outputs(3520) <= not (a xor b);
    outputs(3521) <= a;
    outputs(3522) <= a and not b;
    outputs(3523) <= not (a or b);
    outputs(3524) <= not a;
    outputs(3525) <= a and not b;
    outputs(3526) <= not a;
    outputs(3527) <= not a;
    outputs(3528) <= a;
    outputs(3529) <= not (a xor b);
    outputs(3530) <= b and not a;
    outputs(3531) <= not (a xor b);
    outputs(3532) <= a or b;
    outputs(3533) <= not (a xor b);
    outputs(3534) <= not a or b;
    outputs(3535) <= not (a or b);
    outputs(3536) <= b;
    outputs(3537) <= not (a or b);
    outputs(3538) <= b and not a;
    outputs(3539) <= a;
    outputs(3540) <= not (a and b);
    outputs(3541) <= a xor b;
    outputs(3542) <= not (a xor b);
    outputs(3543) <= not a;
    outputs(3544) <= not (a or b);
    outputs(3545) <= not (a xor b);
    outputs(3546) <= a;
    outputs(3547) <= not (a or b);
    outputs(3548) <= b;
    outputs(3549) <= not (a or b);
    outputs(3550) <= not b;
    outputs(3551) <= a;
    outputs(3552) <= not a;
    outputs(3553) <= not (a xor b);
    outputs(3554) <= b and not a;
    outputs(3555) <= a;
    outputs(3556) <= not (a xor b);
    outputs(3557) <= not b or a;
    outputs(3558) <= not (a or b);
    outputs(3559) <= b;
    outputs(3560) <= a xor b;
    outputs(3561) <= not b;
    outputs(3562) <= a xor b;
    outputs(3563) <= not (a or b);
    outputs(3564) <= not a;
    outputs(3565) <= not a;
    outputs(3566) <= not b;
    outputs(3567) <= not (a xor b);
    outputs(3568) <= not a;
    outputs(3569) <= a;
    outputs(3570) <= a and b;
    outputs(3571) <= a xor b;
    outputs(3572) <= b;
    outputs(3573) <= b;
    outputs(3574) <= not b;
    outputs(3575) <= not b or a;
    outputs(3576) <= not (a xor b);
    outputs(3577) <= not a;
    outputs(3578) <= not a;
    outputs(3579) <= not a;
    outputs(3580) <= b;
    outputs(3581) <= not (a or b);
    outputs(3582) <= a xor b;
    outputs(3583) <= b;
    outputs(3584) <= b;
    outputs(3585) <= a or b;
    outputs(3586) <= not a;
    outputs(3587) <= a xor b;
    outputs(3588) <= a xor b;
    outputs(3589) <= not (a xor b);
    outputs(3590) <= a and not b;
    outputs(3591) <= not b;
    outputs(3592) <= a and b;
    outputs(3593) <= not b or a;
    outputs(3594) <= not a;
    outputs(3595) <= not a or b;
    outputs(3596) <= not a;
    outputs(3597) <= a;
    outputs(3598) <= not a;
    outputs(3599) <= not b;
    outputs(3600) <= b and not a;
    outputs(3601) <= not (a or b);
    outputs(3602) <= not (a xor b);
    outputs(3603) <= a and not b;
    outputs(3604) <= b and not a;
    outputs(3605) <= not b;
    outputs(3606) <= not a;
    outputs(3607) <= a xor b;
    outputs(3608) <= b;
    outputs(3609) <= not b;
    outputs(3610) <= a;
    outputs(3611) <= not a;
    outputs(3612) <= not (a xor b);
    outputs(3613) <= not a;
    outputs(3614) <= not (a xor b);
    outputs(3615) <= not b;
    outputs(3616) <= b and not a;
    outputs(3617) <= not (a xor b);
    outputs(3618) <= not a;
    outputs(3619) <= not (a and b);
    outputs(3620) <= not (a xor b);
    outputs(3621) <= not b or a;
    outputs(3622) <= not a or b;
    outputs(3623) <= a xor b;
    outputs(3624) <= not a;
    outputs(3625) <= b and not a;
    outputs(3626) <= b and not a;
    outputs(3627) <= not (a xor b);
    outputs(3628) <= a;
    outputs(3629) <= not b;
    outputs(3630) <= b and not a;
    outputs(3631) <= a and b;
    outputs(3632) <= not (a xor b);
    outputs(3633) <= b and not a;
    outputs(3634) <= not a;
    outputs(3635) <= not (a or b);
    outputs(3636) <= not (a and b);
    outputs(3637) <= not a;
    outputs(3638) <= not b;
    outputs(3639) <= a or b;
    outputs(3640) <= a and not b;
    outputs(3641) <= not (a or b);
    outputs(3642) <= not (a xor b);
    outputs(3643) <= not a;
    outputs(3644) <= b and not a;
    outputs(3645) <= b;
    outputs(3646) <= not (a xor b);
    outputs(3647) <= not b;
    outputs(3648) <= a xor b;
    outputs(3649) <= not a;
    outputs(3650) <= not a;
    outputs(3651) <= not (a or b);
    outputs(3652) <= not a;
    outputs(3653) <= b;
    outputs(3654) <= not (a xor b);
    outputs(3655) <= a and not b;
    outputs(3656) <= not a;
    outputs(3657) <= a;
    outputs(3658) <= a and not b;
    outputs(3659) <= a xor b;
    outputs(3660) <= not a;
    outputs(3661) <= a;
    outputs(3662) <= not b;
    outputs(3663) <= not (a xor b);
    outputs(3664) <= not a;
    outputs(3665) <= not b or a;
    outputs(3666) <= a;
    outputs(3667) <= not b;
    outputs(3668) <= a and b;
    outputs(3669) <= not b;
    outputs(3670) <= a;
    outputs(3671) <= b;
    outputs(3672) <= not a;
    outputs(3673) <= not b;
    outputs(3674) <= b;
    outputs(3675) <= a;
    outputs(3676) <= a or b;
    outputs(3677) <= b and not a;
    outputs(3678) <= not b;
    outputs(3679) <= b;
    outputs(3680) <= not (a or b);
    outputs(3681) <= a;
    outputs(3682) <= b;
    outputs(3683) <= a;
    outputs(3684) <= not a;
    outputs(3685) <= a or b;
    outputs(3686) <= not b;
    outputs(3687) <= a;
    outputs(3688) <= a;
    outputs(3689) <= a or b;
    outputs(3690) <= not (a xor b);
    outputs(3691) <= b and not a;
    outputs(3692) <= a and not b;
    outputs(3693) <= b;
    outputs(3694) <= not (a xor b);
    outputs(3695) <= b;
    outputs(3696) <= a and not b;
    outputs(3697) <= not (a xor b);
    outputs(3698) <= not a or b;
    outputs(3699) <= a;
    outputs(3700) <= b;
    outputs(3701) <= a and b;
    outputs(3702) <= not a;
    outputs(3703) <= not (a xor b);
    outputs(3704) <= not a;
    outputs(3705) <= not a;
    outputs(3706) <= not a;
    outputs(3707) <= a and not b;
    outputs(3708) <= b;
    outputs(3709) <= a or b;
    outputs(3710) <= not a;
    outputs(3711) <= not (a xor b);
    outputs(3712) <= not (a xor b);
    outputs(3713) <= not (a xor b);
    outputs(3714) <= not b;
    outputs(3715) <= b;
    outputs(3716) <= b;
    outputs(3717) <= b;
    outputs(3718) <= not (a xor b);
    outputs(3719) <= a;
    outputs(3720) <= a;
    outputs(3721) <= b;
    outputs(3722) <= b;
    outputs(3723) <= a;
    outputs(3724) <= a and b;
    outputs(3725) <= not (a or b);
    outputs(3726) <= a;
    outputs(3727) <= not (a xor b);
    outputs(3728) <= not a;
    outputs(3729) <= a;
    outputs(3730) <= b and not a;
    outputs(3731) <= a;
    outputs(3732) <= not b;
    outputs(3733) <= a xor b;
    outputs(3734) <= a;
    outputs(3735) <= a or b;
    outputs(3736) <= not (a xor b);
    outputs(3737) <= a and b;
    outputs(3738) <= a;
    outputs(3739) <= a or b;
    outputs(3740) <= not (a xor b);
    outputs(3741) <= a;
    outputs(3742) <= b;
    outputs(3743) <= not b;
    outputs(3744) <= b and not a;
    outputs(3745) <= not b;
    outputs(3746) <= a;
    outputs(3747) <= a;
    outputs(3748) <= not (a or b);
    outputs(3749) <= not a;
    outputs(3750) <= a and not b;
    outputs(3751) <= not a or b;
    outputs(3752) <= not (a xor b);
    outputs(3753) <= not (a and b);
    outputs(3754) <= not (a or b);
    outputs(3755) <= b;
    outputs(3756) <= a xor b;
    outputs(3757) <= not (a xor b);
    outputs(3758) <= not (a or b);
    outputs(3759) <= a;
    outputs(3760) <= not (a xor b);
    outputs(3761) <= a xor b;
    outputs(3762) <= not (a or b);
    outputs(3763) <= not a;
    outputs(3764) <= not b;
    outputs(3765) <= not a or b;
    outputs(3766) <= b;
    outputs(3767) <= a and not b;
    outputs(3768) <= not b;
    outputs(3769) <= not a;
    outputs(3770) <= not (a or b);
    outputs(3771) <= not b;
    outputs(3772) <= b;
    outputs(3773) <= not a;
    outputs(3774) <= not (a xor b);
    outputs(3775) <= not b;
    outputs(3776) <= a and b;
    outputs(3777) <= not a;
    outputs(3778) <= not (a xor b);
    outputs(3779) <= not b;
    outputs(3780) <= a xor b;
    outputs(3781) <= not (a xor b);
    outputs(3782) <= b;
    outputs(3783) <= not (a and b);
    outputs(3784) <= not b;
    outputs(3785) <= b;
    outputs(3786) <= b;
    outputs(3787) <= a and not b;
    outputs(3788) <= a and b;
    outputs(3789) <= a xor b;
    outputs(3790) <= b and not a;
    outputs(3791) <= not a;
    outputs(3792) <= a;
    outputs(3793) <= a xor b;
    outputs(3794) <= b;
    outputs(3795) <= a xor b;
    outputs(3796) <= b and not a;
    outputs(3797) <= not (a xor b);
    outputs(3798) <= not (a xor b);
    outputs(3799) <= b;
    outputs(3800) <= not (a or b);
    outputs(3801) <= not (a xor b);
    outputs(3802) <= a or b;
    outputs(3803) <= b;
    outputs(3804) <= a xor b;
    outputs(3805) <= b;
    outputs(3806) <= a and not b;
    outputs(3807) <= a and not b;
    outputs(3808) <= a xor b;
    outputs(3809) <= a xor b;
    outputs(3810) <= not a;
    outputs(3811) <= a;
    outputs(3812) <= a or b;
    outputs(3813) <= b;
    outputs(3814) <= a;
    outputs(3815) <= not (a or b);
    outputs(3816) <= not b;
    outputs(3817) <= not a;
    outputs(3818) <= b and not a;
    outputs(3819) <= not a;
    outputs(3820) <= a;
    outputs(3821) <= b;
    outputs(3822) <= a;
    outputs(3823) <= a xor b;
    outputs(3824) <= b;
    outputs(3825) <= b and not a;
    outputs(3826) <= a;
    outputs(3827) <= a xor b;
    outputs(3828) <= not a;
    outputs(3829) <= a xor b;
    outputs(3830) <= not b;
    outputs(3831) <= not (a and b);
    outputs(3832) <= a;
    outputs(3833) <= a;
    outputs(3834) <= a and not b;
    outputs(3835) <= b and not a;
    outputs(3836) <= not b;
    outputs(3837) <= not a;
    outputs(3838) <= not b;
    outputs(3839) <= b;
    outputs(3840) <= a;
    outputs(3841) <= a;
    outputs(3842) <= not (a xor b);
    outputs(3843) <= not a;
    outputs(3844) <= not b;
    outputs(3845) <= not a;
    outputs(3846) <= a xor b;
    outputs(3847) <= not (a xor b);
    outputs(3848) <= a xor b;
    outputs(3849) <= not (a xor b);
    outputs(3850) <= not (a xor b);
    outputs(3851) <= a xor b;
    outputs(3852) <= not a;
    outputs(3853) <= not b;
    outputs(3854) <= a xor b;
    outputs(3855) <= a and b;
    outputs(3856) <= not b;
    outputs(3857) <= not b;
    outputs(3858) <= not (a and b);
    outputs(3859) <= not a;
    outputs(3860) <= not (a xor b);
    outputs(3861) <= not (a xor b);
    outputs(3862) <= not b;
    outputs(3863) <= not a;
    outputs(3864) <= a;
    outputs(3865) <= a xor b;
    outputs(3866) <= not b or a;
    outputs(3867) <= a;
    outputs(3868) <= a and b;
    outputs(3869) <= not b or a;
    outputs(3870) <= b;
    outputs(3871) <= a xor b;
    outputs(3872) <= a xor b;
    outputs(3873) <= a xor b;
    outputs(3874) <= not (a or b);
    outputs(3875) <= not a;
    outputs(3876) <= a xor b;
    outputs(3877) <= a or b;
    outputs(3878) <= not b;
    outputs(3879) <= not b;
    outputs(3880) <= not b;
    outputs(3881) <= a and not b;
    outputs(3882) <= a;
    outputs(3883) <= not (a xor b);
    outputs(3884) <= b and not a;
    outputs(3885) <= not a;
    outputs(3886) <= a xor b;
    outputs(3887) <= not (a and b);
    outputs(3888) <= a and not b;
    outputs(3889) <= not b;
    outputs(3890) <= not a;
    outputs(3891) <= not (a and b);
    outputs(3892) <= a;
    outputs(3893) <= not a;
    outputs(3894) <= not b or a;
    outputs(3895) <= a;
    outputs(3896) <= b and not a;
    outputs(3897) <= a xor b;
    outputs(3898) <= a xor b;
    outputs(3899) <= b and not a;
    outputs(3900) <= not (a xor b);
    outputs(3901) <= not (a and b);
    outputs(3902) <= not a;
    outputs(3903) <= a xor b;
    outputs(3904) <= a and not b;
    outputs(3905) <= a;
    outputs(3906) <= not b;
    outputs(3907) <= a xor b;
    outputs(3908) <= b and not a;
    outputs(3909) <= a;
    outputs(3910) <= not b;
    outputs(3911) <= a or b;
    outputs(3912) <= not (a xor b);
    outputs(3913) <= not a;
    outputs(3914) <= b;
    outputs(3915) <= a;
    outputs(3916) <= not a;
    outputs(3917) <= not b;
    outputs(3918) <= not (a xor b);
    outputs(3919) <= not (a xor b);
    outputs(3920) <= a or b;
    outputs(3921) <= b and not a;
    outputs(3922) <= not a or b;
    outputs(3923) <= b;
    outputs(3924) <= not a;
    outputs(3925) <= not (a xor b);
    outputs(3926) <= b;
    outputs(3927) <= a;
    outputs(3928) <= not b;
    outputs(3929) <= b;
    outputs(3930) <= not (a xor b);
    outputs(3931) <= not (a xor b);
    outputs(3932) <= a xor b;
    outputs(3933) <= b;
    outputs(3934) <= b;
    outputs(3935) <= a xor b;
    outputs(3936) <= not a or b;
    outputs(3937) <= a xor b;
    outputs(3938) <= not a;
    outputs(3939) <= b;
    outputs(3940) <= not b or a;
    outputs(3941) <= a;
    outputs(3942) <= not (a or b);
    outputs(3943) <= b;
    outputs(3944) <= not b;
    outputs(3945) <= not b;
    outputs(3946) <= a or b;
    outputs(3947) <= a xor b;
    outputs(3948) <= not (a xor b);
    outputs(3949) <= a xor b;
    outputs(3950) <= a xor b;
    outputs(3951) <= a xor b;
    outputs(3952) <= not (a xor b);
    outputs(3953) <= b;
    outputs(3954) <= a or b;
    outputs(3955) <= not b;
    outputs(3956) <= b;
    outputs(3957) <= not (a xor b);
    outputs(3958) <= not (a xor b);
    outputs(3959) <= b;
    outputs(3960) <= a and not b;
    outputs(3961) <= a or b;
    outputs(3962) <= not (a and b);
    outputs(3963) <= not a;
    outputs(3964) <= a xor b;
    outputs(3965) <= a;
    outputs(3966) <= not a;
    outputs(3967) <= not b;
    outputs(3968) <= not b or a;
    outputs(3969) <= a xor b;
    outputs(3970) <= not b;
    outputs(3971) <= a xor b;
    outputs(3972) <= a and not b;
    outputs(3973) <= not (a or b);
    outputs(3974) <= a;
    outputs(3975) <= not a or b;
    outputs(3976) <= not b;
    outputs(3977) <= b;
    outputs(3978) <= b;
    outputs(3979) <= a and b;
    outputs(3980) <= not b;
    outputs(3981) <= a and not b;
    outputs(3982) <= not b;
    outputs(3983) <= a xor b;
    outputs(3984) <= not a or b;
    outputs(3985) <= b;
    outputs(3986) <= a xor b;
    outputs(3987) <= a;
    outputs(3988) <= a;
    outputs(3989) <= a xor b;
    outputs(3990) <= b and not a;
    outputs(3991) <= not a;
    outputs(3992) <= not b;
    outputs(3993) <= a xor b;
    outputs(3994) <= a xor b;
    outputs(3995) <= not b or a;
    outputs(3996) <= a;
    outputs(3997) <= not a;
    outputs(3998) <= not (a xor b);
    outputs(3999) <= not (a or b);
    outputs(4000) <= not b;
    outputs(4001) <= a xor b;
    outputs(4002) <= b;
    outputs(4003) <= not a;
    outputs(4004) <= a;
    outputs(4005) <= a;
    outputs(4006) <= a and not b;
    outputs(4007) <= not (a and b);
    outputs(4008) <= not (a or b);
    outputs(4009) <= not a or b;
    outputs(4010) <= not (a and b);
    outputs(4011) <= a and b;
    outputs(4012) <= not (a xor b);
    outputs(4013) <= not a;
    outputs(4014) <= b;
    outputs(4015) <= not a;
    outputs(4016) <= a and b;
    outputs(4017) <= a;
    outputs(4018) <= a xor b;
    outputs(4019) <= b and not a;
    outputs(4020) <= b;
    outputs(4021) <= a or b;
    outputs(4022) <= not b;
    outputs(4023) <= not (a or b);
    outputs(4024) <= a;
    outputs(4025) <= not a;
    outputs(4026) <= a;
    outputs(4027) <= a xor b;
    outputs(4028) <= not (a or b);
    outputs(4029) <= not (a xor b);
    outputs(4030) <= b;
    outputs(4031) <= not b;
    outputs(4032) <= not (a xor b);
    outputs(4033) <= not (a xor b);
    outputs(4034) <= a xor b;
    outputs(4035) <= a xor b;
    outputs(4036) <= b;
    outputs(4037) <= b and not a;
    outputs(4038) <= b;
    outputs(4039) <= not (a xor b);
    outputs(4040) <= a xor b;
    outputs(4041) <= a;
    outputs(4042) <= a xor b;
    outputs(4043) <= not b;
    outputs(4044) <= not (a xor b);
    outputs(4045) <= not b;
    outputs(4046) <= not (a xor b);
    outputs(4047) <= a and b;
    outputs(4048) <= a xor b;
    outputs(4049) <= a;
    outputs(4050) <= not a or b;
    outputs(4051) <= b;
    outputs(4052) <= not (a xor b);
    outputs(4053) <= not b;
    outputs(4054) <= not (a xor b);
    outputs(4055) <= a;
    outputs(4056) <= a;
    outputs(4057) <= not a;
    outputs(4058) <= not a;
    outputs(4059) <= a;
    outputs(4060) <= not b or a;
    outputs(4061) <= b and not a;
    outputs(4062) <= not b;
    outputs(4063) <= not b;
    outputs(4064) <= not b;
    outputs(4065) <= a xor b;
    outputs(4066) <= not a;
    outputs(4067) <= not b;
    outputs(4068) <= not (a xor b);
    outputs(4069) <= not (a or b);
    outputs(4070) <= not a or b;
    outputs(4071) <= not (a xor b);
    outputs(4072) <= a xor b;
    outputs(4073) <= a and b;
    outputs(4074) <= a and b;
    outputs(4075) <= not (a xor b);
    outputs(4076) <= b;
    outputs(4077) <= not a;
    outputs(4078) <= not (a xor b);
    outputs(4079) <= not (a xor b);
    outputs(4080) <= a;
    outputs(4081) <= not a;
    outputs(4082) <= a and b;
    outputs(4083) <= a xor b;
    outputs(4084) <= a xor b;
    outputs(4085) <= a xor b;
    outputs(4086) <= a;
    outputs(4087) <= a xor b;
    outputs(4088) <= a and not b;
    outputs(4089) <= not b;
    outputs(4090) <= a xor b;
    outputs(4091) <= not (a xor b);
    outputs(4092) <= a and not b;
    outputs(4093) <= a;
    outputs(4094) <= a;
    outputs(4095) <= b;
    outputs(4096) <= not (a xor b);
    outputs(4097) <= not (a xor b);
    outputs(4098) <= not b;
    outputs(4099) <= b;
    outputs(4100) <= b and not a;
    outputs(4101) <= not (a xor b);
    outputs(4102) <= not b;
    outputs(4103) <= not a;
    outputs(4104) <= b;
    outputs(4105) <= b and not a;
    outputs(4106) <= a xor b;
    outputs(4107) <= not a;
    outputs(4108) <= not b;
    outputs(4109) <= not (a xor b);
    outputs(4110) <= not (a or b);
    outputs(4111) <= not a;
    outputs(4112) <= not (a xor b);
    outputs(4113) <= b;
    outputs(4114) <= a;
    outputs(4115) <= not (a xor b);
    outputs(4116) <= a and not b;
    outputs(4117) <= a and not b;
    outputs(4118) <= not b;
    outputs(4119) <= a or b;
    outputs(4120) <= a xor b;
    outputs(4121) <= not (a or b);
    outputs(4122) <= b;
    outputs(4123) <= not b;
    outputs(4124) <= a xor b;
    outputs(4125) <= b;
    outputs(4126) <= not b or a;
    outputs(4127) <= a xor b;
    outputs(4128) <= not (a xor b);
    outputs(4129) <= a xor b;
    outputs(4130) <= not (a and b);
    outputs(4131) <= a or b;
    outputs(4132) <= b and not a;
    outputs(4133) <= not b or a;
    outputs(4134) <= a or b;
    outputs(4135) <= b and not a;
    outputs(4136) <= a or b;
    outputs(4137) <= a xor b;
    outputs(4138) <= a and not b;
    outputs(4139) <= a xor b;
    outputs(4140) <= not a;
    outputs(4141) <= a;
    outputs(4142) <= not a;
    outputs(4143) <= not (a xor b);
    outputs(4144) <= a and b;
    outputs(4145) <= not (a xor b);
    outputs(4146) <= a or b;
    outputs(4147) <= not b;
    outputs(4148) <= not (a xor b);
    outputs(4149) <= a xor b;
    outputs(4150) <= a xor b;
    outputs(4151) <= a and not b;
    outputs(4152) <= not b;
    outputs(4153) <= not b;
    outputs(4154) <= not (a xor b);
    outputs(4155) <= a;
    outputs(4156) <= not a;
    outputs(4157) <= a xor b;
    outputs(4158) <= not a;
    outputs(4159) <= a or b;
    outputs(4160) <= not a;
    outputs(4161) <= a xor b;
    outputs(4162) <= not (a xor b);
    outputs(4163) <= not (a xor b);
    outputs(4164) <= a and b;
    outputs(4165) <= a;
    outputs(4166) <= not a or b;
    outputs(4167) <= a and not b;
    outputs(4168) <= a xor b;
    outputs(4169) <= a and b;
    outputs(4170) <= b;
    outputs(4171) <= not (a xor b);
    outputs(4172) <= b;
    outputs(4173) <= b;
    outputs(4174) <= b;
    outputs(4175) <= a xor b;
    outputs(4176) <= a xor b;
    outputs(4177) <= b;
    outputs(4178) <= b;
    outputs(4179) <= a xor b;
    outputs(4180) <= not (a and b);
    outputs(4181) <= a xor b;
    outputs(4182) <= not a or b;
    outputs(4183) <= not a;
    outputs(4184) <= a;
    outputs(4185) <= b;
    outputs(4186) <= not (a xor b);
    outputs(4187) <= a;
    outputs(4188) <= not b;
    outputs(4189) <= not a;
    outputs(4190) <= not b;
    outputs(4191) <= a xor b;
    outputs(4192) <= a xor b;
    outputs(4193) <= b;
    outputs(4194) <= not a;
    outputs(4195) <= a and b;
    outputs(4196) <= not (a xor b);
    outputs(4197) <= not b;
    outputs(4198) <= b;
    outputs(4199) <= b;
    outputs(4200) <= not b;
    outputs(4201) <= not b;
    outputs(4202) <= b and not a;
    outputs(4203) <= not (a xor b);
    outputs(4204) <= not b;
    outputs(4205) <= not a;
    outputs(4206) <= b;
    outputs(4207) <= b and not a;
    outputs(4208) <= a;
    outputs(4209) <= a;
    outputs(4210) <= not (a or b);
    outputs(4211) <= a;
    outputs(4212) <= not a or b;
    outputs(4213) <= not (a xor b);
    outputs(4214) <= not b or a;
    outputs(4215) <= not (a xor b);
    outputs(4216) <= not b;
    outputs(4217) <= not b;
    outputs(4218) <= a xor b;
    outputs(4219) <= a;
    outputs(4220) <= not (a xor b);
    outputs(4221) <= a xor b;
    outputs(4222) <= not (a or b);
    outputs(4223) <= a;
    outputs(4224) <= a or b;
    outputs(4225) <= not (a xor b);
    outputs(4226) <= not (a xor b);
    outputs(4227) <= not (a xor b);
    outputs(4228) <= not a;
    outputs(4229) <= b and not a;
    outputs(4230) <= b;
    outputs(4231) <= not a;
    outputs(4232) <= not (a xor b);
    outputs(4233) <= a xor b;
    outputs(4234) <= not (a xor b);
    outputs(4235) <= b;
    outputs(4236) <= b;
    outputs(4237) <= a;
    outputs(4238) <= not (a xor b);
    outputs(4239) <= a xor b;
    outputs(4240) <= not a;
    outputs(4241) <= not a;
    outputs(4242) <= not (a xor b);
    outputs(4243) <= not a;
    outputs(4244) <= not (a xor b);
    outputs(4245) <= not a or b;
    outputs(4246) <= not b;
    outputs(4247) <= not a;
    outputs(4248) <= not a;
    outputs(4249) <= not a;
    outputs(4250) <= not a or b;
    outputs(4251) <= a and not b;
    outputs(4252) <= not (a xor b);
    outputs(4253) <= not (a xor b);
    outputs(4254) <= not (a xor b);
    outputs(4255) <= a or b;
    outputs(4256) <= not a or b;
    outputs(4257) <= not (a or b);
    outputs(4258) <= a and not b;
    outputs(4259) <= not (a xor b);
    outputs(4260) <= a;
    outputs(4261) <= not (a xor b);
    outputs(4262) <= b;
    outputs(4263) <= not a;
    outputs(4264) <= b;
    outputs(4265) <= a or b;
    outputs(4266) <= not a;
    outputs(4267) <= not (a xor b);
    outputs(4268) <= not b or a;
    outputs(4269) <= not a;
    outputs(4270) <= not b;
    outputs(4271) <= b and not a;
    outputs(4272) <= b;
    outputs(4273) <= a or b;
    outputs(4274) <= b;
    outputs(4275) <= a and b;
    outputs(4276) <= a;
    outputs(4277) <= not (a xor b);
    outputs(4278) <= not b;
    outputs(4279) <= a xor b;
    outputs(4280) <= not b;
    outputs(4281) <= not (a xor b);
    outputs(4282) <= a;
    outputs(4283) <= a xor b;
    outputs(4284) <= not (a xor b);
    outputs(4285) <= not a or b;
    outputs(4286) <= not (a xor b);
    outputs(4287) <= a xor b;
    outputs(4288) <= a xor b;
    outputs(4289) <= a or b;
    outputs(4290) <= not (a or b);
    outputs(4291) <= a xor b;
    outputs(4292) <= a;
    outputs(4293) <= a xor b;
    outputs(4294) <= not (a or b);
    outputs(4295) <= a and b;
    outputs(4296) <= b;
    outputs(4297) <= not b;
    outputs(4298) <= a xor b;
    outputs(4299) <= not b or a;
    outputs(4300) <= not (a xor b);
    outputs(4301) <= not (a and b);
    outputs(4302) <= not (a xor b);
    outputs(4303) <= not a;
    outputs(4304) <= a;
    outputs(4305) <= not b;
    outputs(4306) <= b;
    outputs(4307) <= a and b;
    outputs(4308) <= a xor b;
    outputs(4309) <= not b;
    outputs(4310) <= not (a xor b);
    outputs(4311) <= b and not a;
    outputs(4312) <= not (a xor b);
    outputs(4313) <= a or b;
    outputs(4314) <= not b;
    outputs(4315) <= not (a xor b);
    outputs(4316) <= not b;
    outputs(4317) <= not a;
    outputs(4318) <= not (a xor b);
    outputs(4319) <= a xor b;
    outputs(4320) <= not b;
    outputs(4321) <= not b;
    outputs(4322) <= not b;
    outputs(4323) <= a and not b;
    outputs(4324) <= b;
    outputs(4325) <= a or b;
    outputs(4326) <= not (a xor b);
    outputs(4327) <= a or b;
    outputs(4328) <= a;
    outputs(4329) <= a or b;
    outputs(4330) <= a;
    outputs(4331) <= a and not b;
    outputs(4332) <= not (a xor b);
    outputs(4333) <= b;
    outputs(4334) <= a;
    outputs(4335) <= a xor b;
    outputs(4336) <= not (a xor b);
    outputs(4337) <= not (a xor b);
    outputs(4338) <= a xor b;
    outputs(4339) <= a and not b;
    outputs(4340) <= not (a xor b);
    outputs(4341) <= a and b;
    outputs(4342) <= a xor b;
    outputs(4343) <= a xor b;
    outputs(4344) <= not (a and b);
    outputs(4345) <= a xor b;
    outputs(4346) <= not (a or b);
    outputs(4347) <= a;
    outputs(4348) <= not a;
    outputs(4349) <= b;
    outputs(4350) <= not (a or b);
    outputs(4351) <= a;
    outputs(4352) <= not (a or b);
    outputs(4353) <= a xor b;
    outputs(4354) <= a xor b;
    outputs(4355) <= not b;
    outputs(4356) <= a;
    outputs(4357) <= a;
    outputs(4358) <= b;
    outputs(4359) <= not (a xor b);
    outputs(4360) <= not (a or b);
    outputs(4361) <= not b;
    outputs(4362) <= not (a xor b);
    outputs(4363) <= not (a xor b);
    outputs(4364) <= b and not a;
    outputs(4365) <= a xor b;
    outputs(4366) <= a;
    outputs(4367) <= not (a or b);
    outputs(4368) <= b;
    outputs(4369) <= not (a xor b);
    outputs(4370) <= a;
    outputs(4371) <= a and b;
    outputs(4372) <= not (a xor b);
    outputs(4373) <= not b;
    outputs(4374) <= a or b;
    outputs(4375) <= not b or a;
    outputs(4376) <= not a;
    outputs(4377) <= not a or b;
    outputs(4378) <= b;
    outputs(4379) <= b;
    outputs(4380) <= a xor b;
    outputs(4381) <= not a;
    outputs(4382) <= not (a and b);
    outputs(4383) <= a xor b;
    outputs(4384) <= b and not a;
    outputs(4385) <= a;
    outputs(4386) <= a and b;
    outputs(4387) <= a;
    outputs(4388) <= a and not b;
    outputs(4389) <= b and not a;
    outputs(4390) <= not b;
    outputs(4391) <= a;
    outputs(4392) <= not (a xor b);
    outputs(4393) <= not (a xor b);
    outputs(4394) <= not (a xor b);
    outputs(4395) <= not a;
    outputs(4396) <= a;
    outputs(4397) <= a xor b;
    outputs(4398) <= a and b;
    outputs(4399) <= not b;
    outputs(4400) <= not (a xor b);
    outputs(4401) <= not b or a;
    outputs(4402) <= not (a and b);
    outputs(4403) <= a;
    outputs(4404) <= not b;
    outputs(4405) <= not a;
    outputs(4406) <= not a;
    outputs(4407) <= b and not a;
    outputs(4408) <= not (a xor b);
    outputs(4409) <= not (a and b);
    outputs(4410) <= a xor b;
    outputs(4411) <= not b;
    outputs(4412) <= not b;
    outputs(4413) <= a;
    outputs(4414) <= not a or b;
    outputs(4415) <= a or b;
    outputs(4416) <= a xor b;
    outputs(4417) <= a xor b;
    outputs(4418) <= a;
    outputs(4419) <= a;
    outputs(4420) <= a xor b;
    outputs(4421) <= a xor b;
    outputs(4422) <= not a;
    outputs(4423) <= b;
    outputs(4424) <= a xor b;
    outputs(4425) <= a and b;
    outputs(4426) <= not (a xor b);
    outputs(4427) <= not (a xor b);
    outputs(4428) <= a;
    outputs(4429) <= b;
    outputs(4430) <= a xor b;
    outputs(4431) <= not b or a;
    outputs(4432) <= a and b;
    outputs(4433) <= a and b;
    outputs(4434) <= not (a or b);
    outputs(4435) <= not b;
    outputs(4436) <= b;
    outputs(4437) <= a xor b;
    outputs(4438) <= a;
    outputs(4439) <= not b or a;
    outputs(4440) <= b;
    outputs(4441) <= not (a xor b);
    outputs(4442) <= a;
    outputs(4443) <= not b;
    outputs(4444) <= not a or b;
    outputs(4445) <= b and not a;
    outputs(4446) <= a xor b;
    outputs(4447) <= not a;
    outputs(4448) <= a and b;
    outputs(4449) <= not a or b;
    outputs(4450) <= a or b;
    outputs(4451) <= not b;
    outputs(4452) <= a xor b;
    outputs(4453) <= b;
    outputs(4454) <= not (a xor b);
    outputs(4455) <= not a;
    outputs(4456) <= a xor b;
    outputs(4457) <= a xor b;
    outputs(4458) <= not b;
    outputs(4459) <= not a;
    outputs(4460) <= not b;
    outputs(4461) <= not b or a;
    outputs(4462) <= not (a and b);
    outputs(4463) <= a and b;
    outputs(4464) <= a or b;
    outputs(4465) <= b;
    outputs(4466) <= not b;
    outputs(4467) <= not b;
    outputs(4468) <= a xor b;
    outputs(4469) <= b;
    outputs(4470) <= not (a xor b);
    outputs(4471) <= not b;
    outputs(4472) <= not (a xor b);
    outputs(4473) <= a and b;
    outputs(4474) <= b;
    outputs(4475) <= a xor b;
    outputs(4476) <= not (a xor b);
    outputs(4477) <= not b;
    outputs(4478) <= a and b;
    outputs(4479) <= not a;
    outputs(4480) <= not a or b;
    outputs(4481) <= b;
    outputs(4482) <= not b;
    outputs(4483) <= not b;
    outputs(4484) <= not a;
    outputs(4485) <= not a;
    outputs(4486) <= not (a xor b);
    outputs(4487) <= a and b;
    outputs(4488) <= not b or a;
    outputs(4489) <= a xor b;
    outputs(4490) <= not b;
    outputs(4491) <= not b;
    outputs(4492) <= a xor b;
    outputs(4493) <= b;
    outputs(4494) <= not a;
    outputs(4495) <= a and b;
    outputs(4496) <= a;
    outputs(4497) <= b;
    outputs(4498) <= a xor b;
    outputs(4499) <= a;
    outputs(4500) <= a xor b;
    outputs(4501) <= not (a or b);
    outputs(4502) <= not b;
    outputs(4503) <= not (a xor b);
    outputs(4504) <= not b;
    outputs(4505) <= not a;
    outputs(4506) <= not (a xor b);
    outputs(4507) <= not b or a;
    outputs(4508) <= not (a or b);
    outputs(4509) <= a xor b;
    outputs(4510) <= a xor b;
    outputs(4511) <= not a or b;
    outputs(4512) <= a;
    outputs(4513) <= b;
    outputs(4514) <= a;
    outputs(4515) <= not (a and b);
    outputs(4516) <= not b;
    outputs(4517) <= not (a or b);
    outputs(4518) <= not a or b;
    outputs(4519) <= not (a xor b);
    outputs(4520) <= a xor b;
    outputs(4521) <= not (a xor b);
    outputs(4522) <= not b or a;
    outputs(4523) <= not (a xor b);
    outputs(4524) <= b and not a;
    outputs(4525) <= a or b;
    outputs(4526) <= a;
    outputs(4527) <= a xor b;
    outputs(4528) <= not (a or b);
    outputs(4529) <= a xor b;
    outputs(4530) <= not (a xor b);
    outputs(4531) <= not b or a;
    outputs(4532) <= not b;
    outputs(4533) <= not b;
    outputs(4534) <= not b or a;
    outputs(4535) <= a and not b;
    outputs(4536) <= a and not b;
    outputs(4537) <= b;
    outputs(4538) <= b;
    outputs(4539) <= not b;
    outputs(4540) <= not b;
    outputs(4541) <= a and not b;
    outputs(4542) <= not (a xor b);
    outputs(4543) <= not a;
    outputs(4544) <= b;
    outputs(4545) <= not b or a;
    outputs(4546) <= not b or a;
    outputs(4547) <= a and not b;
    outputs(4548) <= b;
    outputs(4549) <= not a;
    outputs(4550) <= not (a and b);
    outputs(4551) <= b and not a;
    outputs(4552) <= a;
    outputs(4553) <= not a;
    outputs(4554) <= not b;
    outputs(4555) <= a xor b;
    outputs(4556) <= a and not b;
    outputs(4557) <= not a;
    outputs(4558) <= not (a or b);
    outputs(4559) <= b;
    outputs(4560) <= b;
    outputs(4561) <= not b;
    outputs(4562) <= a and b;
    outputs(4563) <= a and b;
    outputs(4564) <= not b;
    outputs(4565) <= not a or b;
    outputs(4566) <= not a or b;
    outputs(4567) <= a xor b;
    outputs(4568) <= a;
    outputs(4569) <= a;
    outputs(4570) <= a;
    outputs(4571) <= not a;
    outputs(4572) <= b and not a;
    outputs(4573) <= not (a and b);
    outputs(4574) <= a xor b;
    outputs(4575) <= not (a or b);
    outputs(4576) <= a;
    outputs(4577) <= a;
    outputs(4578) <= b and not a;
    outputs(4579) <= a and not b;
    outputs(4580) <= not (a or b);
    outputs(4581) <= a xor b;
    outputs(4582) <= a xor b;
    outputs(4583) <= b;
    outputs(4584) <= not (a xor b);
    outputs(4585) <= b;
    outputs(4586) <= a and b;
    outputs(4587) <= not a;
    outputs(4588) <= not b;
    outputs(4589) <= not b;
    outputs(4590) <= b and not a;
    outputs(4591) <= not (a or b);
    outputs(4592) <= not (a xor b);
    outputs(4593) <= a xor b;
    outputs(4594) <= a and not b;
    outputs(4595) <= not (a xor b);
    outputs(4596) <= not (a xor b);
    outputs(4597) <= not b;
    outputs(4598) <= b;
    outputs(4599) <= a xor b;
    outputs(4600) <= not (a xor b);
    outputs(4601) <= a;
    outputs(4602) <= not a or b;
    outputs(4603) <= not a or b;
    outputs(4604) <= b;
    outputs(4605) <= not b;
    outputs(4606) <= a;
    outputs(4607) <= not b;
    outputs(4608) <= a;
    outputs(4609) <= a xor b;
    outputs(4610) <= not b;
    outputs(4611) <= not (a xor b);
    outputs(4612) <= not a;
    outputs(4613) <= a and b;
    outputs(4614) <= not b;
    outputs(4615) <= b;
    outputs(4616) <= not a;
    outputs(4617) <= a;
    outputs(4618) <= not a;
    outputs(4619) <= not b;
    outputs(4620) <= not b;
    outputs(4621) <= not (a and b);
    outputs(4622) <= not a or b;
    outputs(4623) <= not (a xor b);
    outputs(4624) <= not b;
    outputs(4625) <= not a;
    outputs(4626) <= a xor b;
    outputs(4627) <= not b;
    outputs(4628) <= a;
    outputs(4629) <= a;
    outputs(4630) <= not a or b;
    outputs(4631) <= b;
    outputs(4632) <= a;
    outputs(4633) <= a;
    outputs(4634) <= a or b;
    outputs(4635) <= not (a and b);
    outputs(4636) <= a;
    outputs(4637) <= not (a xor b);
    outputs(4638) <= not a;
    outputs(4639) <= not b or a;
    outputs(4640) <= not a;
    outputs(4641) <= not b;
    outputs(4642) <= not b or a;
    outputs(4643) <= not (a xor b);
    outputs(4644) <= b;
    outputs(4645) <= not a;
    outputs(4646) <= not b;
    outputs(4647) <= a;
    outputs(4648) <= b;
    outputs(4649) <= not (a xor b);
    outputs(4650) <= a and not b;
    outputs(4651) <= a xor b;
    outputs(4652) <= a xor b;
    outputs(4653) <= not b;
    outputs(4654) <= not a;
    outputs(4655) <= not a;
    outputs(4656) <= a xor b;
    outputs(4657) <= not a;
    outputs(4658) <= b;
    outputs(4659) <= not a;
    outputs(4660) <= a;
    outputs(4661) <= not b;
    outputs(4662) <= not b;
    outputs(4663) <= b;
    outputs(4664) <= a xor b;
    outputs(4665) <= a xor b;
    outputs(4666) <= not b or a;
    outputs(4667) <= a xor b;
    outputs(4668) <= not a or b;
    outputs(4669) <= b;
    outputs(4670) <= b;
    outputs(4671) <= a and b;
    outputs(4672) <= not (a xor b);
    outputs(4673) <= a and b;
    outputs(4674) <= a;
    outputs(4675) <= b;
    outputs(4676) <= not b;
    outputs(4677) <= a xor b;
    outputs(4678) <= a xor b;
    outputs(4679) <= a xor b;
    outputs(4680) <= a xor b;
    outputs(4681) <= not b;
    outputs(4682) <= b;
    outputs(4683) <= a;
    outputs(4684) <= not b;
    outputs(4685) <= a xor b;
    outputs(4686) <= a xor b;
    outputs(4687) <= not b;
    outputs(4688) <= not (a xor b);
    outputs(4689) <= a;
    outputs(4690) <= not (a xor b);
    outputs(4691) <= a;
    outputs(4692) <= not a;
    outputs(4693) <= not (a xor b);
    outputs(4694) <= a and not b;
    outputs(4695) <= b and not a;
    outputs(4696) <= a;
    outputs(4697) <= not (a xor b);
    outputs(4698) <= not b or a;
    outputs(4699) <= a xor b;
    outputs(4700) <= b;
    outputs(4701) <= a or b;
    outputs(4702) <= not a;
    outputs(4703) <= a xor b;
    outputs(4704) <= b;
    outputs(4705) <= a and b;
    outputs(4706) <= b and not a;
    outputs(4707) <= a xor b;
    outputs(4708) <= a;
    outputs(4709) <= b;
    outputs(4710) <= a xor b;
    outputs(4711) <= a xor b;
    outputs(4712) <= not (a xor b);
    outputs(4713) <= not (a xor b);
    outputs(4714) <= not (a xor b);
    outputs(4715) <= a xor b;
    outputs(4716) <= not (a or b);
    outputs(4717) <= not (a xor b);
    outputs(4718) <= b;
    outputs(4719) <= not (a xor b);
    outputs(4720) <= a xor b;
    outputs(4721) <= not b or a;
    outputs(4722) <= not b;
    outputs(4723) <= a xor b;
    outputs(4724) <= a;
    outputs(4725) <= a xor b;
    outputs(4726) <= not b;
    outputs(4727) <= not b;
    outputs(4728) <= a;
    outputs(4729) <= a;
    outputs(4730) <= a;
    outputs(4731) <= not b;
    outputs(4732) <= a;
    outputs(4733) <= a;
    outputs(4734) <= not (a xor b);
    outputs(4735) <= a and b;
    outputs(4736) <= a xor b;
    outputs(4737) <= a and not b;
    outputs(4738) <= a or b;
    outputs(4739) <= a;
    outputs(4740) <= b;
    outputs(4741) <= b and not a;
    outputs(4742) <= not (a xor b);
    outputs(4743) <= a;
    outputs(4744) <= not b;
    outputs(4745) <= a and b;
    outputs(4746) <= b;
    outputs(4747) <= a;
    outputs(4748) <= not (a xor b);
    outputs(4749) <= b;
    outputs(4750) <= not a;
    outputs(4751) <= not a;
    outputs(4752) <= not (a xor b);
    outputs(4753) <= a xor b;
    outputs(4754) <= not (a xor b);
    outputs(4755) <= b;
    outputs(4756) <= a or b;
    outputs(4757) <= a xor b;
    outputs(4758) <= not (a xor b);
    outputs(4759) <= not b;
    outputs(4760) <= not a;
    outputs(4761) <= not b;
    outputs(4762) <= not (a or b);
    outputs(4763) <= a;
    outputs(4764) <= not b;
    outputs(4765) <= not (a xor b);
    outputs(4766) <= not b;
    outputs(4767) <= not (a xor b);
    outputs(4768) <= a;
    outputs(4769) <= a;
    outputs(4770) <= not (a xor b);
    outputs(4771) <= not a;
    outputs(4772) <= a xor b;
    outputs(4773) <= b;
    outputs(4774) <= not (a xor b);
    outputs(4775) <= b and not a;
    outputs(4776) <= b;
    outputs(4777) <= a;
    outputs(4778) <= not (a xor b);
    outputs(4779) <= not (a xor b);
    outputs(4780) <= b and not a;
    outputs(4781) <= a and b;
    outputs(4782) <= not (a or b);
    outputs(4783) <= b;
    outputs(4784) <= not a;
    outputs(4785) <= a xor b;
    outputs(4786) <= a;
    outputs(4787) <= b;
    outputs(4788) <= a or b;
    outputs(4789) <= a;
    outputs(4790) <= b;
    outputs(4791) <= not (a xor b);
    outputs(4792) <= not a;
    outputs(4793) <= a;
    outputs(4794) <= not a;
    outputs(4795) <= not b;
    outputs(4796) <= a or b;
    outputs(4797) <= not b;
    outputs(4798) <= not b;
    outputs(4799) <= b and not a;
    outputs(4800) <= a;
    outputs(4801) <= a;
    outputs(4802) <= a xor b;
    outputs(4803) <= a and b;
    outputs(4804) <= a xor b;
    outputs(4805) <= b;
    outputs(4806) <= b;
    outputs(4807) <= a;
    outputs(4808) <= a and b;
    outputs(4809) <= b;
    outputs(4810) <= a xor b;
    outputs(4811) <= not a;
    outputs(4812) <= a xor b;
    outputs(4813) <= not a;
    outputs(4814) <= not (a xor b);
    outputs(4815) <= a xor b;
    outputs(4816) <= a and not b;
    outputs(4817) <= not a;
    outputs(4818) <= not (a xor b);
    outputs(4819) <= a xor b;
    outputs(4820) <= not (a and b);
    outputs(4821) <= b;
    outputs(4822) <= a;
    outputs(4823) <= b;
    outputs(4824) <= not a;
    outputs(4825) <= not (a xor b);
    outputs(4826) <= a xor b;
    outputs(4827) <= not b;
    outputs(4828) <= a xor b;
    outputs(4829) <= not (a xor b);
    outputs(4830) <= b and not a;
    outputs(4831) <= not (a xor b);
    outputs(4832) <= a and not b;
    outputs(4833) <= not a;
    outputs(4834) <= not b;
    outputs(4835) <= not a;
    outputs(4836) <= not a;
    outputs(4837) <= not (a xor b);
    outputs(4838) <= not (a xor b);
    outputs(4839) <= not (a xor b);
    outputs(4840) <= a and not b;
    outputs(4841) <= not b;
    outputs(4842) <= not a;
    outputs(4843) <= a xor b;
    outputs(4844) <= not a or b;
    outputs(4845) <= not b;
    outputs(4846) <= not a;
    outputs(4847) <= not a;
    outputs(4848) <= not b;
    outputs(4849) <= not b or a;
    outputs(4850) <= not b;
    outputs(4851) <= not (a xor b);
    outputs(4852) <= not (a xor b);
    outputs(4853) <= b;
    outputs(4854) <= a;
    outputs(4855) <= not b or a;
    outputs(4856) <= not (a xor b);
    outputs(4857) <= a xor b;
    outputs(4858) <= a;
    outputs(4859) <= not (a xor b);
    outputs(4860) <= a xor b;
    outputs(4861) <= a or b;
    outputs(4862) <= b;
    outputs(4863) <= a;
    outputs(4864) <= a;
    outputs(4865) <= not (a or b);
    outputs(4866) <= not b;
    outputs(4867) <= not (a xor b);
    outputs(4868) <= not b;
    outputs(4869) <= not (a xor b);
    outputs(4870) <= not (a or b);
    outputs(4871) <= a and not b;
    outputs(4872) <= a;
    outputs(4873) <= not (a xor b);
    outputs(4874) <= a xor b;
    outputs(4875) <= b and not a;
    outputs(4876) <= not (a xor b);
    outputs(4877) <= a xor b;
    outputs(4878) <= not (a xor b);
    outputs(4879) <= a;
    outputs(4880) <= not a;
    outputs(4881) <= b and not a;
    outputs(4882) <= not a or b;
    outputs(4883) <= not (a xor b);
    outputs(4884) <= not a or b;
    outputs(4885) <= b;
    outputs(4886) <= b;
    outputs(4887) <= not (a xor b);
    outputs(4888) <= b and not a;
    outputs(4889) <= b and not a;
    outputs(4890) <= a;
    outputs(4891) <= not b;
    outputs(4892) <= b;
    outputs(4893) <= not (a xor b);
    outputs(4894) <= a xor b;
    outputs(4895) <= a xor b;
    outputs(4896) <= a;
    outputs(4897) <= not b;
    outputs(4898) <= not a;
    outputs(4899) <= b;
    outputs(4900) <= a;
    outputs(4901) <= a xor b;
    outputs(4902) <= a;
    outputs(4903) <= a and not b;
    outputs(4904) <= a;
    outputs(4905) <= not (a xor b);
    outputs(4906) <= a;
    outputs(4907) <= not (a xor b);
    outputs(4908) <= b;
    outputs(4909) <= a;
    outputs(4910) <= not a;
    outputs(4911) <= not (a xor b);
    outputs(4912) <= not (a xor b);
    outputs(4913) <= not b or a;
    outputs(4914) <= not (a xor b);
    outputs(4915) <= not a;
    outputs(4916) <= not (a or b);
    outputs(4917) <= a xor b;
    outputs(4918) <= not (a xor b);
    outputs(4919) <= b;
    outputs(4920) <= b and not a;
    outputs(4921) <= b;
    outputs(4922) <= a and b;
    outputs(4923) <= b;
    outputs(4924) <= not a;
    outputs(4925) <= not (a or b);
    outputs(4926) <= a xor b;
    outputs(4927) <= b;
    outputs(4928) <= not b;
    outputs(4929) <= not (a xor b);
    outputs(4930) <= a xor b;
    outputs(4931) <= not (a xor b);
    outputs(4932) <= not b;
    outputs(4933) <= b;
    outputs(4934) <= b;
    outputs(4935) <= not (a xor b);
    outputs(4936) <= not b;
    outputs(4937) <= a and not b;
    outputs(4938) <= not b;
    outputs(4939) <= a;
    outputs(4940) <= b;
    outputs(4941) <= a;
    outputs(4942) <= not b or a;
    outputs(4943) <= b;
    outputs(4944) <= not b;
    outputs(4945) <= not (a xor b);
    outputs(4946) <= not b;
    outputs(4947) <= a and b;
    outputs(4948) <= not b;
    outputs(4949) <= not (a and b);
    outputs(4950) <= not a;
    outputs(4951) <= not (a xor b);
    outputs(4952) <= b;
    outputs(4953) <= not (a xor b);
    outputs(4954) <= not (a xor b);
    outputs(4955) <= a and b;
    outputs(4956) <= not (a and b);
    outputs(4957) <= a xor b;
    outputs(4958) <= not (a and b);
    outputs(4959) <= a xor b;
    outputs(4960) <= not b;
    outputs(4961) <= not a;
    outputs(4962) <= a and b;
    outputs(4963) <= not (a or b);
    outputs(4964) <= a xor b;
    outputs(4965) <= not (a xor b);
    outputs(4966) <= a;
    outputs(4967) <= b;
    outputs(4968) <= a;
    outputs(4969) <= not a;
    outputs(4970) <= b;
    outputs(4971) <= not b;
    outputs(4972) <= a;
    outputs(4973) <= not (a xor b);
    outputs(4974) <= not a or b;
    outputs(4975) <= not b;
    outputs(4976) <= not b;
    outputs(4977) <= a;
    outputs(4978) <= a xor b;
    outputs(4979) <= not (a xor b);
    outputs(4980) <= not (a xor b);
    outputs(4981) <= b;
    outputs(4982) <= not a;
    outputs(4983) <= a xor b;
    outputs(4984) <= not a;
    outputs(4985) <= not (a xor b);
    outputs(4986) <= not (a or b);
    outputs(4987) <= not a;
    outputs(4988) <= not a;
    outputs(4989) <= a;
    outputs(4990) <= not (a or b);
    outputs(4991) <= not b;
    outputs(4992) <= not (a xor b);
    outputs(4993) <= not a;
    outputs(4994) <= a and b;
    outputs(4995) <= b;
    outputs(4996) <= not b;
    outputs(4997) <= a xor b;
    outputs(4998) <= a and b;
    outputs(4999) <= a xor b;
    outputs(5000) <= a;
    outputs(5001) <= not a;
    outputs(5002) <= not b;
    outputs(5003) <= b;
    outputs(5004) <= not (a and b);
    outputs(5005) <= not a;
    outputs(5006) <= not a or b;
    outputs(5007) <= not a or b;
    outputs(5008) <= a;
    outputs(5009) <= a or b;
    outputs(5010) <= not a;
    outputs(5011) <= a xor b;
    outputs(5012) <= b;
    outputs(5013) <= not (a xor b);
    outputs(5014) <= b and not a;
    outputs(5015) <= not (a and b);
    outputs(5016) <= not a;
    outputs(5017) <= a and b;
    outputs(5018) <= not a or b;
    outputs(5019) <= a;
    outputs(5020) <= not b;
    outputs(5021) <= not b;
    outputs(5022) <= a xor b;
    outputs(5023) <= a and b;
    outputs(5024) <= b;
    outputs(5025) <= a xor b;
    outputs(5026) <= not (a xor b);
    outputs(5027) <= not b;
    outputs(5028) <= not b;
    outputs(5029) <= b;
    outputs(5030) <= not (a xor b);
    outputs(5031) <= not b;
    outputs(5032) <= a xor b;
    outputs(5033) <= not b;
    outputs(5034) <= not (a or b);
    outputs(5035) <= not (a and b);
    outputs(5036) <= not b;
    outputs(5037) <= a or b;
    outputs(5038) <= not b;
    outputs(5039) <= not (a xor b);
    outputs(5040) <= not a;
    outputs(5041) <= a;
    outputs(5042) <= not (a xor b);
    outputs(5043) <= not (a xor b);
    outputs(5044) <= a and b;
    outputs(5045) <= a xor b;
    outputs(5046) <= not a;
    outputs(5047) <= not (a xor b);
    outputs(5048) <= a;
    outputs(5049) <= not b;
    outputs(5050) <= a xor b;
    outputs(5051) <= not b;
    outputs(5052) <= b;
    outputs(5053) <= a xor b;
    outputs(5054) <= not a;
    outputs(5055) <= a;
    outputs(5056) <= b;
    outputs(5057) <= a;
    outputs(5058) <= not b or a;
    outputs(5059) <= not (a or b);
    outputs(5060) <= a;
    outputs(5061) <= not a or b;
    outputs(5062) <= not a;
    outputs(5063) <= a xor b;
    outputs(5064) <= b and not a;
    outputs(5065) <= b and not a;
    outputs(5066) <= b;
    outputs(5067) <= not (a xor b);
    outputs(5068) <= not (a or b);
    outputs(5069) <= a xor b;
    outputs(5070) <= not a;
    outputs(5071) <= not (a or b);
    outputs(5072) <= a and not b;
    outputs(5073) <= not (a and b);
    outputs(5074) <= not b or a;
    outputs(5075) <= not (a and b);
    outputs(5076) <= a xor b;
    outputs(5077) <= not a;
    outputs(5078) <= b;
    outputs(5079) <= a;
    outputs(5080) <= b;
    outputs(5081) <= b;
    outputs(5082) <= not b;
    outputs(5083) <= not (a xor b);
    outputs(5084) <= not (a and b);
    outputs(5085) <= a and not b;
    outputs(5086) <= not b or a;
    outputs(5087) <= not (a xor b);
    outputs(5088) <= b;
    outputs(5089) <= not a;
    outputs(5090) <= not b;
    outputs(5091) <= not b or a;
    outputs(5092) <= a and b;
    outputs(5093) <= not a;
    outputs(5094) <= a;
    outputs(5095) <= not (a xor b);
    outputs(5096) <= a;
    outputs(5097) <= not (a xor b);
    outputs(5098) <= not a or b;
    outputs(5099) <= a;
    outputs(5100) <= not (a xor b);
    outputs(5101) <= not a or b;
    outputs(5102) <= not (a or b);
    outputs(5103) <= b;
    outputs(5104) <= a;
    outputs(5105) <= not a;
    outputs(5106) <= a xor b;
    outputs(5107) <= not (a and b);
    outputs(5108) <= not a;
    outputs(5109) <= a and not b;
    outputs(5110) <= not b;
    outputs(5111) <= b;
    outputs(5112) <= b;
    outputs(5113) <= a xor b;
    outputs(5114) <= not (a xor b);
    outputs(5115) <= a;
    outputs(5116) <= not a;
    outputs(5117) <= not a;
    outputs(5118) <= not (a xor b);
    outputs(5119) <= a xor b;
    outputs(5120) <= not b or a;
    outputs(5121) <= not (a and b);
    outputs(5122) <= not (a xor b);
    outputs(5123) <= not (a or b);
    outputs(5124) <= b;
    outputs(5125) <= not b;
    outputs(5126) <= b;
    outputs(5127) <= not a;
    outputs(5128) <= not (a xor b);
    outputs(5129) <= a xor b;
    outputs(5130) <= not b or a;
    outputs(5131) <= a xor b;
    outputs(5132) <= a xor b;
    outputs(5133) <= a;
    outputs(5134) <= a;
    outputs(5135) <= not (a xor b);
    outputs(5136) <= a and b;
    outputs(5137) <= not (a and b);
    outputs(5138) <= a xor b;
    outputs(5139) <= a xor b;
    outputs(5140) <= not b;
    outputs(5141) <= a xor b;
    outputs(5142) <= a xor b;
    outputs(5143) <= b and not a;
    outputs(5144) <= not (a xor b);
    outputs(5145) <= a xor b;
    outputs(5146) <= not b;
    outputs(5147) <= a xor b;
    outputs(5148) <= not a;
    outputs(5149) <= not a;
    outputs(5150) <= not a;
    outputs(5151) <= not a;
    outputs(5152) <= a xor b;
    outputs(5153) <= b and not a;
    outputs(5154) <= not (a xor b);
    outputs(5155) <= not (a xor b);
    outputs(5156) <= b;
    outputs(5157) <= not (a or b);
    outputs(5158) <= not b;
    outputs(5159) <= not (a xor b);
    outputs(5160) <= a or b;
    outputs(5161) <= not a;
    outputs(5162) <= a or b;
    outputs(5163) <= b;
    outputs(5164) <= not b;
    outputs(5165) <= a and b;
    outputs(5166) <= not b;
    outputs(5167) <= a xor b;
    outputs(5168) <= a and not b;
    outputs(5169) <= not (a xor b);
    outputs(5170) <= not b;
    outputs(5171) <= a;
    outputs(5172) <= a;
    outputs(5173) <= not (a or b);
    outputs(5174) <= not a or b;
    outputs(5175) <= not (a or b);
    outputs(5176) <= a xor b;
    outputs(5177) <= not (a or b);
    outputs(5178) <= a and not b;
    outputs(5179) <= a;
    outputs(5180) <= a;
    outputs(5181) <= a xor b;
    outputs(5182) <= not (a and b);
    outputs(5183) <= not (a and b);
    outputs(5184) <= not a;
    outputs(5185) <= b and not a;
    outputs(5186) <= not (a or b);
    outputs(5187) <= a;
    outputs(5188) <= a xor b;
    outputs(5189) <= not a;
    outputs(5190) <= not a;
    outputs(5191) <= not b;
    outputs(5192) <= a xor b;
    outputs(5193) <= not b;
    outputs(5194) <= a;
    outputs(5195) <= a;
    outputs(5196) <= not (a or b);
    outputs(5197) <= b and not a;
    outputs(5198) <= a;
    outputs(5199) <= not b;
    outputs(5200) <= not a or b;
    outputs(5201) <= a;
    outputs(5202) <= not (a or b);
    outputs(5203) <= not (a xor b);
    outputs(5204) <= a and not b;
    outputs(5205) <= a xor b;
    outputs(5206) <= a;
    outputs(5207) <= not (a xor b);
    outputs(5208) <= a and b;
    outputs(5209) <= not b or a;
    outputs(5210) <= not b;
    outputs(5211) <= not b;
    outputs(5212) <= a and b;
    outputs(5213) <= not a;
    outputs(5214) <= a;
    outputs(5215) <= not b or a;
    outputs(5216) <= b;
    outputs(5217) <= not b;
    outputs(5218) <= a xor b;
    outputs(5219) <= not b;
    outputs(5220) <= a xor b;
    outputs(5221) <= not b;
    outputs(5222) <= not b;
    outputs(5223) <= b;
    outputs(5224) <= not a;
    outputs(5225) <= not (a xor b);
    outputs(5226) <= not (a xor b);
    outputs(5227) <= b;
    outputs(5228) <= a;
    outputs(5229) <= not b;
    outputs(5230) <= not b;
    outputs(5231) <= not a;
    outputs(5232) <= b;
    outputs(5233) <= a and b;
    outputs(5234) <= not (a xor b);
    outputs(5235) <= not b or a;
    outputs(5236) <= a;
    outputs(5237) <= a;
    outputs(5238) <= not a;
    outputs(5239) <= not a;
    outputs(5240) <= not b;
    outputs(5241) <= not (a xor b);
    outputs(5242) <= b;
    outputs(5243) <= a xor b;
    outputs(5244) <= not a;
    outputs(5245) <= not a;
    outputs(5246) <= not a;
    outputs(5247) <= not a;
    outputs(5248) <= a;
    outputs(5249) <= b;
    outputs(5250) <= not (a xor b);
    outputs(5251) <= not (a xor b);
    outputs(5252) <= not b;
    outputs(5253) <= not a;
    outputs(5254) <= a and b;
    outputs(5255) <= not (a and b);
    outputs(5256) <= b;
    outputs(5257) <= a xor b;
    outputs(5258) <= a;
    outputs(5259) <= a xor b;
    outputs(5260) <= not (a xor b);
    outputs(5261) <= not a or b;
    outputs(5262) <= not (a and b);
    outputs(5263) <= a;
    outputs(5264) <= not a;
    outputs(5265) <= a and not b;
    outputs(5266) <= not b or a;
    outputs(5267) <= a and not b;
    outputs(5268) <= not a;
    outputs(5269) <= not a;
    outputs(5270) <= not (a or b);
    outputs(5271) <= a;
    outputs(5272) <= a and not b;
    outputs(5273) <= not b;
    outputs(5274) <= not a;
    outputs(5275) <= a xor b;
    outputs(5276) <= a xor b;
    outputs(5277) <= not (a xor b);
    outputs(5278) <= not b;
    outputs(5279) <= not (a xor b);
    outputs(5280) <= b;
    outputs(5281) <= a and not b;
    outputs(5282) <= not b;
    outputs(5283) <= a xor b;
    outputs(5284) <= not (a xor b);
    outputs(5285) <= not (a xor b);
    outputs(5286) <= a xor b;
    outputs(5287) <= not (a xor b);
    outputs(5288) <= a xor b;
    outputs(5289) <= not a;
    outputs(5290) <= not b or a;
    outputs(5291) <= a;
    outputs(5292) <= a xor b;
    outputs(5293) <= not (a xor b);
    outputs(5294) <= not a;
    outputs(5295) <= not (a xor b);
    outputs(5296) <= not b;
    outputs(5297) <= not b;
    outputs(5298) <= not (a xor b);
    outputs(5299) <= not a;
    outputs(5300) <= a or b;
    outputs(5301) <= not (a xor b);
    outputs(5302) <= a xor b;
    outputs(5303) <= a;
    outputs(5304) <= not (a xor b);
    outputs(5305) <= a xor b;
    outputs(5306) <= not (a xor b);
    outputs(5307) <= b;
    outputs(5308) <= a xor b;
    outputs(5309) <= b;
    outputs(5310) <= a and b;
    outputs(5311) <= not (a xor b);
    outputs(5312) <= not b;
    outputs(5313) <= not a or b;
    outputs(5314) <= b;
    outputs(5315) <= not a;
    outputs(5316) <= a;
    outputs(5317) <= not a or b;
    outputs(5318) <= not a;
    outputs(5319) <= not b;
    outputs(5320) <= not a;
    outputs(5321) <= b;
    outputs(5322) <= b;
    outputs(5323) <= a xor b;
    outputs(5324) <= b;
    outputs(5325) <= a and not b;
    outputs(5326) <= not (a and b);
    outputs(5327) <= not (a xor b);
    outputs(5328) <= not b;
    outputs(5329) <= a;
    outputs(5330) <= not (a or b);
    outputs(5331) <= a;
    outputs(5332) <= not b or a;
    outputs(5333) <= not (a and b);
    outputs(5334) <= b;
    outputs(5335) <= not (a xor b);
    outputs(5336) <= not b;
    outputs(5337) <= a;
    outputs(5338) <= a and not b;
    outputs(5339) <= b and not a;
    outputs(5340) <= a and b;
    outputs(5341) <= a xor b;
    outputs(5342) <= not b;
    outputs(5343) <= a xor b;
    outputs(5344) <= a and b;
    outputs(5345) <= not (a xor b);
    outputs(5346) <= a xor b;
    outputs(5347) <= not a;
    outputs(5348) <= not (a xor b);
    outputs(5349) <= not (a xor b);
    outputs(5350) <= not b or a;
    outputs(5351) <= not a;
    outputs(5352) <= not b;
    outputs(5353) <= not b;
    outputs(5354) <= a xor b;
    outputs(5355) <= not (a or b);
    outputs(5356) <= b;
    outputs(5357) <= a xor b;
    outputs(5358) <= not b or a;
    outputs(5359) <= b;
    outputs(5360) <= not (a or b);
    outputs(5361) <= not a;
    outputs(5362) <= a or b;
    outputs(5363) <= not b;
    outputs(5364) <= a xor b;
    outputs(5365) <= not a or b;
    outputs(5366) <= not a;
    outputs(5367) <= not (a xor b);
    outputs(5368) <= not a;
    outputs(5369) <= a xor b;
    outputs(5370) <= a xor b;
    outputs(5371) <= a and b;
    outputs(5372) <= a xor b;
    outputs(5373) <= a;
    outputs(5374) <= a xor b;
    outputs(5375) <= not (a xor b);
    outputs(5376) <= a;
    outputs(5377) <= not b or a;
    outputs(5378) <= not b or a;
    outputs(5379) <= b;
    outputs(5380) <= b and not a;
    outputs(5381) <= b;
    outputs(5382) <= not a;
    outputs(5383) <= not (a or b);
    outputs(5384) <= b and not a;
    outputs(5385) <= a and not b;
    outputs(5386) <= not (a xor b);
    outputs(5387) <= b;
    outputs(5388) <= a and not b;
    outputs(5389) <= not (a xor b);
    outputs(5390) <= not (a xor b);
    outputs(5391) <= b;
    outputs(5392) <= not (a xor b);
    outputs(5393) <= a;
    outputs(5394) <= b;
    outputs(5395) <= a and not b;
    outputs(5396) <= a;
    outputs(5397) <= a xor b;
    outputs(5398) <= not a;
    outputs(5399) <= not (a or b);
    outputs(5400) <= a xor b;
    outputs(5401) <= b;
    outputs(5402) <= not b;
    outputs(5403) <= a xor b;
    outputs(5404) <= not (a xor b);
    outputs(5405) <= a and b;
    outputs(5406) <= b and not a;
    outputs(5407) <= not (a xor b);
    outputs(5408) <= a and not b;
    outputs(5409) <= b and not a;
    outputs(5410) <= not a or b;
    outputs(5411) <= not b;
    outputs(5412) <= a;
    outputs(5413) <= b and not a;
    outputs(5414) <= a xor b;
    outputs(5415) <= not a;
    outputs(5416) <= not (a and b);
    outputs(5417) <= b and not a;
    outputs(5418) <= a xor b;
    outputs(5419) <= b and not a;
    outputs(5420) <= not (a and b);
    outputs(5421) <= a xor b;
    outputs(5422) <= a and b;
    outputs(5423) <= a and not b;
    outputs(5424) <= a;
    outputs(5425) <= b;
    outputs(5426) <= b;
    outputs(5427) <= b;
    outputs(5428) <= b and not a;
    outputs(5429) <= a and not b;
    outputs(5430) <= a;
    outputs(5431) <= not a;
    outputs(5432) <= not (a xor b);
    outputs(5433) <= not a;
    outputs(5434) <= a and b;
    outputs(5435) <= not a;
    outputs(5436) <= not b;
    outputs(5437) <= not b or a;
    outputs(5438) <= not b or a;
    outputs(5439) <= not b;
    outputs(5440) <= a and not b;
    outputs(5441) <= a xor b;
    outputs(5442) <= not (a xor b);
    outputs(5443) <= a;
    outputs(5444) <= not (a xor b);
    outputs(5445) <= not (a or b);
    outputs(5446) <= not (a or b);
    outputs(5447) <= b and not a;
    outputs(5448) <= not a;
    outputs(5449) <= a xor b;
    outputs(5450) <= a;
    outputs(5451) <= a;
    outputs(5452) <= b and not a;
    outputs(5453) <= not b;
    outputs(5454) <= b;
    outputs(5455) <= not (a xor b);
    outputs(5456) <= a and not b;
    outputs(5457) <= not a;
    outputs(5458) <= b;
    outputs(5459) <= b;
    outputs(5460) <= a and not b;
    outputs(5461) <= b;
    outputs(5462) <= b and not a;
    outputs(5463) <= a xor b;
    outputs(5464) <= a;
    outputs(5465) <= not b;
    outputs(5466) <= a xor b;
    outputs(5467) <= b;
    outputs(5468) <= not b;
    outputs(5469) <= a and not b;
    outputs(5470) <= a or b;
    outputs(5471) <= not (a xor b);
    outputs(5472) <= a and not b;
    outputs(5473) <= a xor b;
    outputs(5474) <= not a;
    outputs(5475) <= not (a xor b);
    outputs(5476) <= a;
    outputs(5477) <= not (a or b);
    outputs(5478) <= a and b;
    outputs(5479) <= not a;
    outputs(5480) <= a and not b;
    outputs(5481) <= not (a xor b);
    outputs(5482) <= not b;
    outputs(5483) <= a xor b;
    outputs(5484) <= not (a xor b);
    outputs(5485) <= b;
    outputs(5486) <= not (a xor b);
    outputs(5487) <= not (a xor b);
    outputs(5488) <= a xor b;
    outputs(5489) <= not (a xor b);
    outputs(5490) <= a and not b;
    outputs(5491) <= a xor b;
    outputs(5492) <= not a;
    outputs(5493) <= not a or b;
    outputs(5494) <= a xor b;
    outputs(5495) <= not a;
    outputs(5496) <= a;
    outputs(5497) <= b;
    outputs(5498) <= not b;
    outputs(5499) <= b;
    outputs(5500) <= not a;
    outputs(5501) <= a;
    outputs(5502) <= not (a or b);
    outputs(5503) <= a xor b;
    outputs(5504) <= not a;
    outputs(5505) <= a xor b;
    outputs(5506) <= a xor b;
    outputs(5507) <= a or b;
    outputs(5508) <= b;
    outputs(5509) <= a and not b;
    outputs(5510) <= not b;
    outputs(5511) <= b;
    outputs(5512) <= b;
    outputs(5513) <= not b;
    outputs(5514) <= b;
    outputs(5515) <= not a;
    outputs(5516) <= b;
    outputs(5517) <= b and not a;
    outputs(5518) <= b;
    outputs(5519) <= not b;
    outputs(5520) <= not (a or b);
    outputs(5521) <= a and not b;
    outputs(5522) <= not (a or b);
    outputs(5523) <= b;
    outputs(5524) <= b and not a;
    outputs(5525) <= not a or b;
    outputs(5526) <= not (a xor b);
    outputs(5527) <= not (a or b);
    outputs(5528) <= not a;
    outputs(5529) <= not a;
    outputs(5530) <= not (a xor b);
    outputs(5531) <= a and not b;
    outputs(5532) <= a xor b;
    outputs(5533) <= b;
    outputs(5534) <= a or b;
    outputs(5535) <= b;
    outputs(5536) <= a;
    outputs(5537) <= a;
    outputs(5538) <= not a or b;
    outputs(5539) <= not a;
    outputs(5540) <= b;
    outputs(5541) <= not (a or b);
    outputs(5542) <= a or b;
    outputs(5543) <= not a;
    outputs(5544) <= b;
    outputs(5545) <= not b;
    outputs(5546) <= not (a xor b);
    outputs(5547) <= a;
    outputs(5548) <= a;
    outputs(5549) <= not (a xor b);
    outputs(5550) <= not (a or b);
    outputs(5551) <= not a;
    outputs(5552) <= not (a xor b);
    outputs(5553) <= not a;
    outputs(5554) <= not a;
    outputs(5555) <= a and not b;
    outputs(5556) <= not b or a;
    outputs(5557) <= not b;
    outputs(5558) <= b and not a;
    outputs(5559) <= not b;
    outputs(5560) <= a xor b;
    outputs(5561) <= not (a xor b);
    outputs(5562) <= not a;
    outputs(5563) <= not a;
    outputs(5564) <= not (a or b);
    outputs(5565) <= a and b;
    outputs(5566) <= not a;
    outputs(5567) <= a and not b;
    outputs(5568) <= not (a xor b);
    outputs(5569) <= a and b;
    outputs(5570) <= not (a xor b);
    outputs(5571) <= a;
    outputs(5572) <= not b;
    outputs(5573) <= b;
    outputs(5574) <= a and b;
    outputs(5575) <= b;
    outputs(5576) <= b;
    outputs(5577) <= not (a xor b);
    outputs(5578) <= not b;
    outputs(5579) <= not (a or b);
    outputs(5580) <= not (a xor b);
    outputs(5581) <= b;
    outputs(5582) <= b;
    outputs(5583) <= a xor b;
    outputs(5584) <= a and not b;
    outputs(5585) <= not a or b;
    outputs(5586) <= b;
    outputs(5587) <= a xor b;
    outputs(5588) <= b;
    outputs(5589) <= not (a or b);
    outputs(5590) <= b;
    outputs(5591) <= b and not a;
    outputs(5592) <= a;
    outputs(5593) <= not a;
    outputs(5594) <= not a;
    outputs(5595) <= not b;
    outputs(5596) <= not b;
    outputs(5597) <= a xor b;
    outputs(5598) <= a xor b;
    outputs(5599) <= not (a xor b);
    outputs(5600) <= a and b;
    outputs(5601) <= a;
    outputs(5602) <= b;
    outputs(5603) <= a;
    outputs(5604) <= b;
    outputs(5605) <= not b;
    outputs(5606) <= a;
    outputs(5607) <= a xor b;
    outputs(5608) <= a;
    outputs(5609) <= a xor b;
    outputs(5610) <= a xor b;
    outputs(5611) <= not a;
    outputs(5612) <= not b;
    outputs(5613) <= not (a or b);
    outputs(5614) <= a and b;
    outputs(5615) <= not (a or b);
    outputs(5616) <= not (a xor b);
    outputs(5617) <= not b;
    outputs(5618) <= not (a or b);
    outputs(5619) <= b and not a;
    outputs(5620) <= a;
    outputs(5621) <= not (a xor b);
    outputs(5622) <= a;
    outputs(5623) <= b;
    outputs(5624) <= a xor b;
    outputs(5625) <= not b;
    outputs(5626) <= not a;
    outputs(5627) <= a xor b;
    outputs(5628) <= a and b;
    outputs(5629) <= a xor b;
    outputs(5630) <= a or b;
    outputs(5631) <= a xor b;
    outputs(5632) <= a and not b;
    outputs(5633) <= a and b;
    outputs(5634) <= not (a xor b);
    outputs(5635) <= not (a xor b);
    outputs(5636) <= a xor b;
    outputs(5637) <= not (a and b);
    outputs(5638) <= b;
    outputs(5639) <= not (a xor b);
    outputs(5640) <= b;
    outputs(5641) <= not a;
    outputs(5642) <= not (a xor b);
    outputs(5643) <= a;
    outputs(5644) <= a;
    outputs(5645) <= not b;
    outputs(5646) <= a;
    outputs(5647) <= a or b;
    outputs(5648) <= not a;
    outputs(5649) <= not a;
    outputs(5650) <= b;
    outputs(5651) <= not a;
    outputs(5652) <= a;
    outputs(5653) <= not (a xor b);
    outputs(5654) <= not (a xor b);
    outputs(5655) <= not (a xor b);
    outputs(5656) <= a xor b;
    outputs(5657) <= a and not b;
    outputs(5658) <= a;
    outputs(5659) <= b and not a;
    outputs(5660) <= a and b;
    outputs(5661) <= not (a xor b);
    outputs(5662) <= a and b;
    outputs(5663) <= not (a or b);
    outputs(5664) <= not (a xor b);
    outputs(5665) <= not (a and b);
    outputs(5666) <= b;
    outputs(5667) <= not (a xor b);
    outputs(5668) <= a and b;
    outputs(5669) <= not (a xor b);
    outputs(5670) <= not b or a;
    outputs(5671) <= not (a xor b);
    outputs(5672) <= b;
    outputs(5673) <= not (a xor b);
    outputs(5674) <= not (a xor b);
    outputs(5675) <= b;
    outputs(5676) <= not a;
    outputs(5677) <= a xor b;
    outputs(5678) <= not a;
    outputs(5679) <= a and b;
    outputs(5680) <= a xor b;
    outputs(5681) <= not b;
    outputs(5682) <= not (a xor b);
    outputs(5683) <= not b or a;
    outputs(5684) <= a xor b;
    outputs(5685) <= not (a or b);
    outputs(5686) <= a;
    outputs(5687) <= a and b;
    outputs(5688) <= not a;
    outputs(5689) <= not a;
    outputs(5690) <= a and b;
    outputs(5691) <= b;
    outputs(5692) <= a or b;
    outputs(5693) <= a xor b;
    outputs(5694) <= not a or b;
    outputs(5695) <= not (a xor b);
    outputs(5696) <= not (a or b);
    outputs(5697) <= a xor b;
    outputs(5698) <= not a or b;
    outputs(5699) <= not (a xor b);
    outputs(5700) <= not b;
    outputs(5701) <= a xor b;
    outputs(5702) <= a and b;
    outputs(5703) <= a;
    outputs(5704) <= a xor b;
    outputs(5705) <= not (a xor b);
    outputs(5706) <= a xor b;
    outputs(5707) <= a xor b;
    outputs(5708) <= not (a xor b);
    outputs(5709) <= b;
    outputs(5710) <= not (a or b);
    outputs(5711) <= b;
    outputs(5712) <= not b;
    outputs(5713) <= a;
    outputs(5714) <= a;
    outputs(5715) <= not a;
    outputs(5716) <= a;
    outputs(5717) <= not b;
    outputs(5718) <= a and not b;
    outputs(5719) <= not (a xor b);
    outputs(5720) <= not (a or b);
    outputs(5721) <= not (a xor b);
    outputs(5722) <= b;
    outputs(5723) <= not (a or b);
    outputs(5724) <= b;
    outputs(5725) <= a;
    outputs(5726) <= not a;
    outputs(5727) <= not (a xor b);
    outputs(5728) <= a and not b;
    outputs(5729) <= a xor b;
    outputs(5730) <= b;
    outputs(5731) <= a and not b;
    outputs(5732) <= b;
    outputs(5733) <= b;
    outputs(5734) <= not (a or b);
    outputs(5735) <= not (a or b);
    outputs(5736) <= b;
    outputs(5737) <= a and b;
    outputs(5738) <= not a;
    outputs(5739) <= not b;
    outputs(5740) <= a xor b;
    outputs(5741) <= a xor b;
    outputs(5742) <= not (a or b);
    outputs(5743) <= not b or a;
    outputs(5744) <= a xor b;
    outputs(5745) <= a xor b;
    outputs(5746) <= a xor b;
    outputs(5747) <= a and b;
    outputs(5748) <= not (a xor b);
    outputs(5749) <= not b;
    outputs(5750) <= a and b;
    outputs(5751) <= a and not b;
    outputs(5752) <= not b;
    outputs(5753) <= b;
    outputs(5754) <= not (a xor b);
    outputs(5755) <= a xor b;
    outputs(5756) <= not (a or b);
    outputs(5757) <= not (a xor b);
    outputs(5758) <= b;
    outputs(5759) <= not b;
    outputs(5760) <= not a;
    outputs(5761) <= not (a or b);
    outputs(5762) <= not (a or b);
    outputs(5763) <= a and not b;
    outputs(5764) <= b;
    outputs(5765) <= a and not b;
    outputs(5766) <= b and not a;
    outputs(5767) <= not (a xor b);
    outputs(5768) <= a xor b;
    outputs(5769) <= not (a xor b);
    outputs(5770) <= b;
    outputs(5771) <= not (a xor b);
    outputs(5772) <= not a;
    outputs(5773) <= a and b;
    outputs(5774) <= not (a and b);
    outputs(5775) <= not (a or b);
    outputs(5776) <= not b;
    outputs(5777) <= a;
    outputs(5778) <= a;
    outputs(5779) <= a and b;
    outputs(5780) <= not (a xor b);
    outputs(5781) <= not (a xor b);
    outputs(5782) <= not (a xor b);
    outputs(5783) <= a and b;
    outputs(5784) <= not b;
    outputs(5785) <= a;
    outputs(5786) <= not b;
    outputs(5787) <= not a;
    outputs(5788) <= not (a and b);
    outputs(5789) <= a;
    outputs(5790) <= not a;
    outputs(5791) <= not (a xor b);
    outputs(5792) <= not b;
    outputs(5793) <= not a or b;
    outputs(5794) <= not a or b;
    outputs(5795) <= not b;
    outputs(5796) <= a and b;
    outputs(5797) <= not (a or b);
    outputs(5798) <= a;
    outputs(5799) <= not a;
    outputs(5800) <= b;
    outputs(5801) <= a and b;
    outputs(5802) <= not a or b;
    outputs(5803) <= a;
    outputs(5804) <= not a;
    outputs(5805) <= b;
    outputs(5806) <= not a;
    outputs(5807) <= not a;
    outputs(5808) <= not (a xor b);
    outputs(5809) <= not a;
    outputs(5810) <= a;
    outputs(5811) <= not (a xor b);
    outputs(5812) <= not a;
    outputs(5813) <= a;
    outputs(5814) <= not (a or b);
    outputs(5815) <= not b;
    outputs(5816) <= b;
    outputs(5817) <= not b;
    outputs(5818) <= not a;
    outputs(5819) <= b;
    outputs(5820) <= b;
    outputs(5821) <= not b;
    outputs(5822) <= a xor b;
    outputs(5823) <= not a;
    outputs(5824) <= a and not b;
    outputs(5825) <= not b;
    outputs(5826) <= not a or b;
    outputs(5827) <= a and not b;
    outputs(5828) <= a;
    outputs(5829) <= not a;
    outputs(5830) <= not a;
    outputs(5831) <= not (a xor b);
    outputs(5832) <= b;
    outputs(5833) <= a;
    outputs(5834) <= b;
    outputs(5835) <= not b;
    outputs(5836) <= not (a xor b);
    outputs(5837) <= b;
    outputs(5838) <= a xor b;
    outputs(5839) <= a xor b;
    outputs(5840) <= a and not b;
    outputs(5841) <= a xor b;
    outputs(5842) <= b;
    outputs(5843) <= not (a xor b);
    outputs(5844) <= not b;
    outputs(5845) <= not b or a;
    outputs(5846) <= b and not a;
    outputs(5847) <= a xor b;
    outputs(5848) <= b;
    outputs(5849) <= not b;
    outputs(5850) <= b and not a;
    outputs(5851) <= a and not b;
    outputs(5852) <= not (a xor b);
    outputs(5853) <= not (a xor b);
    outputs(5854) <= not a;
    outputs(5855) <= not b;
    outputs(5856) <= a xor b;
    outputs(5857) <= not b;
    outputs(5858) <= a xor b;
    outputs(5859) <= not (a or b);
    outputs(5860) <= a;
    outputs(5861) <= b;
    outputs(5862) <= not (a or b);
    outputs(5863) <= a xor b;
    outputs(5864) <= not a;
    outputs(5865) <= not (a xor b);
    outputs(5866) <= not a;
    outputs(5867) <= not a;
    outputs(5868) <= not (a xor b);
    outputs(5869) <= a and b;
    outputs(5870) <= not (a xor b);
    outputs(5871) <= a;
    outputs(5872) <= a and not b;
    outputs(5873) <= b;
    outputs(5874) <= not b;
    outputs(5875) <= not a;
    outputs(5876) <= a;
    outputs(5877) <= b and not a;
    outputs(5878) <= a;
    outputs(5879) <= b and not a;
    outputs(5880) <= a and b;
    outputs(5881) <= not (a xor b);
    outputs(5882) <= not b;
    outputs(5883) <= a;
    outputs(5884) <= not (a or b);
    outputs(5885) <= a xor b;
    outputs(5886) <= not (a xor b);
    outputs(5887) <= b;
    outputs(5888) <= not a;
    outputs(5889) <= a xor b;
    outputs(5890) <= not a;
    outputs(5891) <= a and not b;
    outputs(5892) <= a or b;
    outputs(5893) <= not (a xor b);
    outputs(5894) <= a xor b;
    outputs(5895) <= not b;
    outputs(5896) <= b;
    outputs(5897) <= not b;
    outputs(5898) <= not (a xor b);
    outputs(5899) <= a;
    outputs(5900) <= not b;
    outputs(5901) <= not (a xor b);
    outputs(5902) <= a;
    outputs(5903) <= a;
    outputs(5904) <= not (a or b);
    outputs(5905) <= b;
    outputs(5906) <= not b or a;
    outputs(5907) <= b and not a;
    outputs(5908) <= b and not a;
    outputs(5909) <= a xor b;
    outputs(5910) <= not (a xor b);
    outputs(5911) <= not a;
    outputs(5912) <= not b;
    outputs(5913) <= b;
    outputs(5914) <= not (a or b);
    outputs(5915) <= not (a xor b);
    outputs(5916) <= not a or b;
    outputs(5917) <= not (a xor b);
    outputs(5918) <= a xor b;
    outputs(5919) <= a xor b;
    outputs(5920) <= a xor b;
    outputs(5921) <= not a;
    outputs(5922) <= a;
    outputs(5923) <= b;
    outputs(5924) <= not (a or b);
    outputs(5925) <= not a;
    outputs(5926) <= not b;
    outputs(5927) <= not a;
    outputs(5928) <= not a or b;
    outputs(5929) <= b;
    outputs(5930) <= not b;
    outputs(5931) <= not (a or b);
    outputs(5932) <= not a;
    outputs(5933) <= a and not b;
    outputs(5934) <= not (a or b);
    outputs(5935) <= not b;
    outputs(5936) <= b and not a;
    outputs(5937) <= a and not b;
    outputs(5938) <= a and b;
    outputs(5939) <= a;
    outputs(5940) <= a and not b;
    outputs(5941) <= not (a xor b);
    outputs(5942) <= not b;
    outputs(5943) <= not a;
    outputs(5944) <= not (a xor b);
    outputs(5945) <= a xor b;
    outputs(5946) <= b and not a;
    outputs(5947) <= a xor b;
    outputs(5948) <= a xor b;
    outputs(5949) <= a;
    outputs(5950) <= a;
    outputs(5951) <= b and not a;
    outputs(5952) <= a xor b;
    outputs(5953) <= not (a or b);
    outputs(5954) <= not a;
    outputs(5955) <= b;
    outputs(5956) <= not a;
    outputs(5957) <= not (a xor b);
    outputs(5958) <= not a;
    outputs(5959) <= not b;
    outputs(5960) <= a and b;
    outputs(5961) <= b and not a;
    outputs(5962) <= not a or b;
    outputs(5963) <= a;
    outputs(5964) <= not (a xor b);
    outputs(5965) <= not (a xor b);
    outputs(5966) <= a and not b;
    outputs(5967) <= a xor b;
    outputs(5968) <= not (a xor b);
    outputs(5969) <= not a;
    outputs(5970) <= not b;
    outputs(5971) <= a and not b;
    outputs(5972) <= a xor b;
    outputs(5973) <= not (a xor b);
    outputs(5974) <= b and not a;
    outputs(5975) <= not b;
    outputs(5976) <= a or b;
    outputs(5977) <= not (a xor b);
    outputs(5978) <= a;
    outputs(5979) <= b;
    outputs(5980) <= b;
    outputs(5981) <= a;
    outputs(5982) <= not b;
    outputs(5983) <= a xor b;
    outputs(5984) <= not a;
    outputs(5985) <= a xor b;
    outputs(5986) <= b and not a;
    outputs(5987) <= not (a xor b);
    outputs(5988) <= not (a xor b);
    outputs(5989) <= not b;
    outputs(5990) <= not a;
    outputs(5991) <= not a;
    outputs(5992) <= a and b;
    outputs(5993) <= a xor b;
    outputs(5994) <= not (a xor b);
    outputs(5995) <= a and not b;
    outputs(5996) <= not (a xor b);
    outputs(5997) <= a xor b;
    outputs(5998) <= not b;
    outputs(5999) <= b;
    outputs(6000) <= not (a xor b);
    outputs(6001) <= a and not b;
    outputs(6002) <= not b;
    outputs(6003) <= not (a xor b);
    outputs(6004) <= not (a xor b);
    outputs(6005) <= not b;
    outputs(6006) <= a and b;
    outputs(6007) <= b and not a;
    outputs(6008) <= not (a xor b);
    outputs(6009) <= a and not b;
    outputs(6010) <= not (a xor b);
    outputs(6011) <= not b;
    outputs(6012) <= b;
    outputs(6013) <= b;
    outputs(6014) <= a;
    outputs(6015) <= a xor b;
    outputs(6016) <= b and not a;
    outputs(6017) <= not (a xor b);
    outputs(6018) <= b;
    outputs(6019) <= b;
    outputs(6020) <= a xor b;
    outputs(6021) <= not (a xor b);
    outputs(6022) <= not (a xor b);
    outputs(6023) <= not (a xor b);
    outputs(6024) <= a;
    outputs(6025) <= not a;
    outputs(6026) <= b;
    outputs(6027) <= not (a xor b);
    outputs(6028) <= b;
    outputs(6029) <= not a;
    outputs(6030) <= b;
    outputs(6031) <= b;
    outputs(6032) <= not b;
    outputs(6033) <= not a;
    outputs(6034) <= a xor b;
    outputs(6035) <= b;
    outputs(6036) <= a and b;
    outputs(6037) <= a and b;
    outputs(6038) <= not b;
    outputs(6039) <= b;
    outputs(6040) <= a;
    outputs(6041) <= not (a or b);
    outputs(6042) <= not a or b;
    outputs(6043) <= not (a or b);
    outputs(6044) <= a xor b;
    outputs(6045) <= a xor b;
    outputs(6046) <= a;
    outputs(6047) <= not b;
    outputs(6048) <= not (a xor b);
    outputs(6049) <= b and not a;
    outputs(6050) <= not a;
    outputs(6051) <= not a;
    outputs(6052) <= a xor b;
    outputs(6053) <= a xor b;
    outputs(6054) <= not (a xor b);
    outputs(6055) <= a and not b;
    outputs(6056) <= a;
    outputs(6057) <= b and not a;
    outputs(6058) <= a and b;
    outputs(6059) <= b;
    outputs(6060) <= a xor b;
    outputs(6061) <= a;
    outputs(6062) <= b;
    outputs(6063) <= not b;
    outputs(6064) <= not a;
    outputs(6065) <= a or b;
    outputs(6066) <= a;
    outputs(6067) <= not a;
    outputs(6068) <= not (a xor b);
    outputs(6069) <= not (a or b);
    outputs(6070) <= a xor b;
    outputs(6071) <= not (a xor b);
    outputs(6072) <= a or b;
    outputs(6073) <= a xor b;
    outputs(6074) <= a;
    outputs(6075) <= a;
    outputs(6076) <= not (a or b);
    outputs(6077) <= a and b;
    outputs(6078) <= not a;
    outputs(6079) <= a and not b;
    outputs(6080) <= not a or b;
    outputs(6081) <= b;
    outputs(6082) <= not (a or b);
    outputs(6083) <= a;
    outputs(6084) <= b and not a;
    outputs(6085) <= a and not b;
    outputs(6086) <= a xor b;
    outputs(6087) <= a and b;
    outputs(6088) <= not b or a;
    outputs(6089) <= b and not a;
    outputs(6090) <= a xor b;
    outputs(6091) <= a and not b;
    outputs(6092) <= a;
    outputs(6093) <= a and b;
    outputs(6094) <= a;
    outputs(6095) <= a xor b;
    outputs(6096) <= a;
    outputs(6097) <= not (a or b);
    outputs(6098) <= not a;
    outputs(6099) <= a and b;
    outputs(6100) <= not a;
    outputs(6101) <= not b;
    outputs(6102) <= not (a or b);
    outputs(6103) <= not (a xor b);
    outputs(6104) <= a;
    outputs(6105) <= a and b;
    outputs(6106) <= not b;
    outputs(6107) <= not (a xor b);
    outputs(6108) <= not (a xor b);
    outputs(6109) <= not (a xor b);
    outputs(6110) <= b and not a;
    outputs(6111) <= b;
    outputs(6112) <= b and not a;
    outputs(6113) <= b;
    outputs(6114) <= a xor b;
    outputs(6115) <= not a;
    outputs(6116) <= not (a or b);
    outputs(6117) <= b and not a;
    outputs(6118) <= not (a and b);
    outputs(6119) <= a and b;
    outputs(6120) <= a xor b;
    outputs(6121) <= a xor b;
    outputs(6122) <= b;
    outputs(6123) <= a and not b;
    outputs(6124) <= a xor b;
    outputs(6125) <= not (a xor b);
    outputs(6126) <= a;
    outputs(6127) <= b and not a;
    outputs(6128) <= not a or b;
    outputs(6129) <= not (a and b);
    outputs(6130) <= b and not a;
    outputs(6131) <= a and b;
    outputs(6132) <= not (a xor b);
    outputs(6133) <= not b;
    outputs(6134) <= not a;
    outputs(6135) <= not b;
    outputs(6136) <= b;
    outputs(6137) <= not (a or b);
    outputs(6138) <= a;
    outputs(6139) <= not (a xor b);
    outputs(6140) <= not (a xor b);
    outputs(6141) <= b;
    outputs(6142) <= not (a xor b);
    outputs(6143) <= not (a or b);
    outputs(6144) <= not (a xor b);
    outputs(6145) <= not (a xor b);
    outputs(6146) <= not (a xor b);
    outputs(6147) <= not b;
    outputs(6148) <= b;
    outputs(6149) <= not a;
    outputs(6150) <= a;
    outputs(6151) <= a xor b;
    outputs(6152) <= not (a or b);
    outputs(6153) <= b and not a;
    outputs(6154) <= b and not a;
    outputs(6155) <= a;
    outputs(6156) <= a xor b;
    outputs(6157) <= a xor b;
    outputs(6158) <= not (a xor b);
    outputs(6159) <= a xor b;
    outputs(6160) <= a xor b;
    outputs(6161) <= not (a xor b);
    outputs(6162) <= not b;
    outputs(6163) <= not (a xor b);
    outputs(6164) <= b;
    outputs(6165) <= not a;
    outputs(6166) <= not (a xor b);
    outputs(6167) <= not a or b;
    outputs(6168) <= not b;
    outputs(6169) <= a;
    outputs(6170) <= a xor b;
    outputs(6171) <= not b or a;
    outputs(6172) <= not (a xor b);
    outputs(6173) <= not b;
    outputs(6174) <= a xor b;
    outputs(6175) <= b;
    outputs(6176) <= not (a or b);
    outputs(6177) <= not b;
    outputs(6178) <= not b or a;
    outputs(6179) <= not a;
    outputs(6180) <= not b;
    outputs(6181) <= b;
    outputs(6182) <= not (a and b);
    outputs(6183) <= not b or a;
    outputs(6184) <= not (a xor b);
    outputs(6185) <= not b;
    outputs(6186) <= not (a or b);
    outputs(6187) <= not (a xor b);
    outputs(6188) <= not a or b;
    outputs(6189) <= not (a xor b);
    outputs(6190) <= not (a or b);
    outputs(6191) <= b;
    outputs(6192) <= b;
    outputs(6193) <= not (a and b);
    outputs(6194) <= a and b;
    outputs(6195) <= a;
    outputs(6196) <= not a;
    outputs(6197) <= a or b;
    outputs(6198) <= b;
    outputs(6199) <= not a;
    outputs(6200) <= not (a or b);
    outputs(6201) <= not (a or b);
    outputs(6202) <= a xor b;
    outputs(6203) <= a;
    outputs(6204) <= not b;
    outputs(6205) <= a;
    outputs(6206) <= not b;
    outputs(6207) <= b;
    outputs(6208) <= a xor b;
    outputs(6209) <= b;
    outputs(6210) <= not (a xor b);
    outputs(6211) <= not (a or b);
    outputs(6212) <= a and not b;
    outputs(6213) <= not b;
    outputs(6214) <= not b;
    outputs(6215) <= not a;
    outputs(6216) <= not (a xor b);
    outputs(6217) <= b;
    outputs(6218) <= not (a xor b);
    outputs(6219) <= a xor b;
    outputs(6220) <= a;
    outputs(6221) <= not (a and b);
    outputs(6222) <= not a or b;
    outputs(6223) <= a;
    outputs(6224) <= b and not a;
    outputs(6225) <= a;
    outputs(6226) <= a xor b;
    outputs(6227) <= not a or b;
    outputs(6228) <= b;
    outputs(6229) <= a or b;
    outputs(6230) <= not (a or b);
    outputs(6231) <= a xor b;
    outputs(6232) <= a xor b;
    outputs(6233) <= a;
    outputs(6234) <= a and not b;
    outputs(6235) <= not a or b;
    outputs(6236) <= not a or b;
    outputs(6237) <= a;
    outputs(6238) <= not b or a;
    outputs(6239) <= a;
    outputs(6240) <= not (a xor b);
    outputs(6241) <= b;
    outputs(6242) <= not b;
    outputs(6243) <= not a;
    outputs(6244) <= a and b;
    outputs(6245) <= not b;
    outputs(6246) <= not (a xor b);
    outputs(6247) <= not (a xor b);
    outputs(6248) <= a;
    outputs(6249) <= a xor b;
    outputs(6250) <= not (a and b);
    outputs(6251) <= a;
    outputs(6252) <= not a;
    outputs(6253) <= a or b;
    outputs(6254) <= a xor b;
    outputs(6255) <= not (a or b);
    outputs(6256) <= not b;
    outputs(6257) <= not (a xor b);
    outputs(6258) <= not (a xor b);
    outputs(6259) <= a and not b;
    outputs(6260) <= not a;
    outputs(6261) <= b;
    outputs(6262) <= not (a xor b);
    outputs(6263) <= b;
    outputs(6264) <= not a;
    outputs(6265) <= b;
    outputs(6266) <= a xor b;
    outputs(6267) <= not (a and b);
    outputs(6268) <= b and not a;
    outputs(6269) <= b;
    outputs(6270) <= a xor b;
    outputs(6271) <= a xor b;
    outputs(6272) <= a xor b;
    outputs(6273) <= not a;
    outputs(6274) <= b;
    outputs(6275) <= not b;
    outputs(6276) <= not b;
    outputs(6277) <= not (a xor b);
    outputs(6278) <= b;
    outputs(6279) <= not a;
    outputs(6280) <= not (a xor b);
    outputs(6281) <= a xor b;
    outputs(6282) <= not (a xor b);
    outputs(6283) <= a xor b;
    outputs(6284) <= not a or b;
    outputs(6285) <= b;
    outputs(6286) <= not (a or b);
    outputs(6287) <= a xor b;
    outputs(6288) <= b;
    outputs(6289) <= not a;
    outputs(6290) <= not a;
    outputs(6291) <= not (a xor b);
    outputs(6292) <= not b or a;
    outputs(6293) <= not (a or b);
    outputs(6294) <= not b or a;
    outputs(6295) <= a xor b;
    outputs(6296) <= a;
    outputs(6297) <= a or b;
    outputs(6298) <= a;
    outputs(6299) <= not b;
    outputs(6300) <= a;
    outputs(6301) <= not a;
    outputs(6302) <= a xor b;
    outputs(6303) <= b;
    outputs(6304) <= not (a xor b);
    outputs(6305) <= a xor b;
    outputs(6306) <= a;
    outputs(6307) <= a or b;
    outputs(6308) <= a;
    outputs(6309) <= a;
    outputs(6310) <= a;
    outputs(6311) <= not b;
    outputs(6312) <= not (a or b);
    outputs(6313) <= a;
    outputs(6314) <= not b;
    outputs(6315) <= a xor b;
    outputs(6316) <= not a or b;
    outputs(6317) <= not (a xor b);
    outputs(6318) <= not b;
    outputs(6319) <= a and b;
    outputs(6320) <= not b;
    outputs(6321) <= b;
    outputs(6322) <= a xor b;
    outputs(6323) <= not b;
    outputs(6324) <= a;
    outputs(6325) <= not b;
    outputs(6326) <= a;
    outputs(6327) <= not (a or b);
    outputs(6328) <= not a;
    outputs(6329) <= a xor b;
    outputs(6330) <= b;
    outputs(6331) <= a or b;
    outputs(6332) <= not (a xor b);
    outputs(6333) <= not b;
    outputs(6334) <= b;
    outputs(6335) <= a and b;
    outputs(6336) <= a;
    outputs(6337) <= a;
    outputs(6338) <= a;
    outputs(6339) <= not (a and b);
    outputs(6340) <= not (a and b);
    outputs(6341) <= a or b;
    outputs(6342) <= not b;
    outputs(6343) <= a;
    outputs(6344) <= not (a xor b);
    outputs(6345) <= a and b;
    outputs(6346) <= a xor b;
    outputs(6347) <= a;
    outputs(6348) <= not (a xor b);
    outputs(6349) <= not (a xor b);
    outputs(6350) <= a and b;
    outputs(6351) <= not (a and b);
    outputs(6352) <= a xor b;
    outputs(6353) <= not (a xor b);
    outputs(6354) <= a;
    outputs(6355) <= a xor b;
    outputs(6356) <= a xor b;
    outputs(6357) <= not (a xor b);
    outputs(6358) <= not b;
    outputs(6359) <= a xor b;
    outputs(6360) <= not a;
    outputs(6361) <= not b;
    outputs(6362) <= not b or a;
    outputs(6363) <= not (a xor b);
    outputs(6364) <= b;
    outputs(6365) <= not (a xor b);
    outputs(6366) <= a and b;
    outputs(6367) <= b;
    outputs(6368) <= a;
    outputs(6369) <= not a;
    outputs(6370) <= not b;
    outputs(6371) <= b;
    outputs(6372) <= not b;
    outputs(6373) <= not a;
    outputs(6374) <= not (a xor b);
    outputs(6375) <= not b;
    outputs(6376) <= not a;
    outputs(6377) <= b;
    outputs(6378) <= not a or b;
    outputs(6379) <= not (a and b);
    outputs(6380) <= not b;
    outputs(6381) <= a and b;
    outputs(6382) <= a xor b;
    outputs(6383) <= b;
    outputs(6384) <= not b;
    outputs(6385) <= a xor b;
    outputs(6386) <= a xor b;
    outputs(6387) <= not (a and b);
    outputs(6388) <= not b;
    outputs(6389) <= a xor b;
    outputs(6390) <= b and not a;
    outputs(6391) <= not b;
    outputs(6392) <= not b;
    outputs(6393) <= a;
    outputs(6394) <= not (a xor b);
    outputs(6395) <= not (a xor b);
    outputs(6396) <= a;
    outputs(6397) <= not (a and b);
    outputs(6398) <= not (a xor b);
    outputs(6399) <= a;
    outputs(6400) <= a xor b;
    outputs(6401) <= not b;
    outputs(6402) <= not b;
    outputs(6403) <= a;
    outputs(6404) <= a xor b;
    outputs(6405) <= not a;
    outputs(6406) <= not a or b;
    outputs(6407) <= not b;
    outputs(6408) <= a and b;
    outputs(6409) <= a xor b;
    outputs(6410) <= not (a xor b);
    outputs(6411) <= b;
    outputs(6412) <= not (a xor b);
    outputs(6413) <= not b;
    outputs(6414) <= b;
    outputs(6415) <= not (a xor b);
    outputs(6416) <= b and not a;
    outputs(6417) <= not (a xor b);
    outputs(6418) <= not (a xor b);
    outputs(6419) <= not a;
    outputs(6420) <= a xor b;
    outputs(6421) <= a and not b;
    outputs(6422) <= b;
    outputs(6423) <= a or b;
    outputs(6424) <= not a;
    outputs(6425) <= not a;
    outputs(6426) <= b;
    outputs(6427) <= b;
    outputs(6428) <= a xor b;
    outputs(6429) <= a xor b;
    outputs(6430) <= b;
    outputs(6431) <= b;
    outputs(6432) <= b and not a;
    outputs(6433) <= b;
    outputs(6434) <= not (a xor b);
    outputs(6435) <= b;
    outputs(6436) <= not (a or b);
    outputs(6437) <= not a or b;
    outputs(6438) <= not a;
    outputs(6439) <= not a or b;
    outputs(6440) <= a;
    outputs(6441) <= b;
    outputs(6442) <= not a;
    outputs(6443) <= not (a and b);
    outputs(6444) <= a;
    outputs(6445) <= not b;
    outputs(6446) <= not (a xor b);
    outputs(6447) <= not (a and b);
    outputs(6448) <= a xor b;
    outputs(6449) <= not b;
    outputs(6450) <= not a;
    outputs(6451) <= a or b;
    outputs(6452) <= a xor b;
    outputs(6453) <= not (a and b);
    outputs(6454) <= b;
    outputs(6455) <= not b or a;
    outputs(6456) <= not a;
    outputs(6457) <= a xor b;
    outputs(6458) <= not b;
    outputs(6459) <= a;
    outputs(6460) <= not a;
    outputs(6461) <= a xor b;
    outputs(6462) <= not (a or b);
    outputs(6463) <= a and b;
    outputs(6464) <= a;
    outputs(6465) <= a xor b;
    outputs(6466) <= a xor b;
    outputs(6467) <= not (a and b);
    outputs(6468) <= not b or a;
    outputs(6469) <= not b;
    outputs(6470) <= not a or b;
    outputs(6471) <= a xor b;
    outputs(6472) <= not (a xor b);
    outputs(6473) <= b;
    outputs(6474) <= not b;
    outputs(6475) <= not a or b;
    outputs(6476) <= not (a xor b);
    outputs(6477) <= a;
    outputs(6478) <= a xor b;
    outputs(6479) <= not a;
    outputs(6480) <= not b;
    outputs(6481) <= not a or b;
    outputs(6482) <= not a;
    outputs(6483) <= not b;
    outputs(6484) <= not (a xor b);
    outputs(6485) <= a;
    outputs(6486) <= not b;
    outputs(6487) <= not a;
    outputs(6488) <= not a;
    outputs(6489) <= not a or b;
    outputs(6490) <= not b;
    outputs(6491) <= a and not b;
    outputs(6492) <= not (a xor b);
    outputs(6493) <= not (a xor b);
    outputs(6494) <= a or b;
    outputs(6495) <= a;
    outputs(6496) <= not (a xor b);
    outputs(6497) <= a and b;
    outputs(6498) <= not (a xor b);
    outputs(6499) <= a xor b;
    outputs(6500) <= b;
    outputs(6501) <= b;
    outputs(6502) <= not b;
    outputs(6503) <= a xor b;
    outputs(6504) <= a and b;
    outputs(6505) <= not b;
    outputs(6506) <= a xor b;
    outputs(6507) <= not b;
    outputs(6508) <= b;
    outputs(6509) <= not (a xor b);
    outputs(6510) <= not a or b;
    outputs(6511) <= a and not b;
    outputs(6512) <= not a;
    outputs(6513) <= a and not b;
    outputs(6514) <= not a;
    outputs(6515) <= not (a xor b);
    outputs(6516) <= b;
    outputs(6517) <= a;
    outputs(6518) <= a xor b;
    outputs(6519) <= not a;
    outputs(6520) <= not (a xor b);
    outputs(6521) <= not (a xor b);
    outputs(6522) <= a or b;
    outputs(6523) <= a xor b;
    outputs(6524) <= b;
    outputs(6525) <= not a;
    outputs(6526) <= b;
    outputs(6527) <= not (a xor b);
    outputs(6528) <= b;
    outputs(6529) <= b;
    outputs(6530) <= not b;
    outputs(6531) <= a;
    outputs(6532) <= b and not a;
    outputs(6533) <= a or b;
    outputs(6534) <= b;
    outputs(6535) <= not a or b;
    outputs(6536) <= a and b;
    outputs(6537) <= b and not a;
    outputs(6538) <= a and b;
    outputs(6539) <= a xor b;
    outputs(6540) <= a;
    outputs(6541) <= a;
    outputs(6542) <= a;
    outputs(6543) <= not (a xor b);
    outputs(6544) <= b;
    outputs(6545) <= a xor b;
    outputs(6546) <= not (a xor b);
    outputs(6547) <= not b or a;
    outputs(6548) <= not (a xor b);
    outputs(6549) <= not (a and b);
    outputs(6550) <= a;
    outputs(6551) <= a;
    outputs(6552) <= a;
    outputs(6553) <= not a;
    outputs(6554) <= not a or b;
    outputs(6555) <= b;
    outputs(6556) <= not a or b;
    outputs(6557) <= b;
    outputs(6558) <= a xor b;
    outputs(6559) <= a xor b;
    outputs(6560) <= not b;
    outputs(6561) <= not a;
    outputs(6562) <= b;
    outputs(6563) <= not (a and b);
    outputs(6564) <= not b;
    outputs(6565) <= not a;
    outputs(6566) <= not (a xor b);
    outputs(6567) <= not (a xor b);
    outputs(6568) <= a;
    outputs(6569) <= not (a xor b);
    outputs(6570) <= b and not a;
    outputs(6571) <= not a;
    outputs(6572) <= a or b;
    outputs(6573) <= b;
    outputs(6574) <= a;
    outputs(6575) <= not (a xor b);
    outputs(6576) <= b;
    outputs(6577) <= a;
    outputs(6578) <= not (a xor b);
    outputs(6579) <= a;
    outputs(6580) <= not a;
    outputs(6581) <= not b;
    outputs(6582) <= not (a xor b);
    outputs(6583) <= not b;
    outputs(6584) <= not (a xor b);
    outputs(6585) <= not (a xor b);
    outputs(6586) <= not (a xor b);
    outputs(6587) <= b;
    outputs(6588) <= a xor b;
    outputs(6589) <= not a;
    outputs(6590) <= not a;
    outputs(6591) <= not (a xor b);
    outputs(6592) <= a or b;
    outputs(6593) <= a;
    outputs(6594) <= b;
    outputs(6595) <= not a;
    outputs(6596) <= not (a or b);
    outputs(6597) <= a and not b;
    outputs(6598) <= not (a or b);
    outputs(6599) <= a or b;
    outputs(6600) <= b and not a;
    outputs(6601) <= not b;
    outputs(6602) <= not (a or b);
    outputs(6603) <= a xor b;
    outputs(6604) <= not (a xor b);
    outputs(6605) <= not b or a;
    outputs(6606) <= not (a xor b);
    outputs(6607) <= b;
    outputs(6608) <= not (a xor b);
    outputs(6609) <= not (a xor b);
    outputs(6610) <= a;
    outputs(6611) <= a xor b;
    outputs(6612) <= a;
    outputs(6613) <= not (a and b);
    outputs(6614) <= a xor b;
    outputs(6615) <= not (a xor b);
    outputs(6616) <= a xor b;
    outputs(6617) <= a;
    outputs(6618) <= not a;
    outputs(6619) <= a;
    outputs(6620) <= a xor b;
    outputs(6621) <= not b or a;
    outputs(6622) <= b and not a;
    outputs(6623) <= not (a xor b);
    outputs(6624) <= a;
    outputs(6625) <= a;
    outputs(6626) <= b;
    outputs(6627) <= a xor b;
    outputs(6628) <= b;
    outputs(6629) <= a;
    outputs(6630) <= not a;
    outputs(6631) <= not a;
    outputs(6632) <= not (a xor b);
    outputs(6633) <= not a or b;
    outputs(6634) <= a and not b;
    outputs(6635) <= not a;
    outputs(6636) <= a xor b;
    outputs(6637) <= a;
    outputs(6638) <= b;
    outputs(6639) <= not a or b;
    outputs(6640) <= a xor b;
    outputs(6641) <= b and not a;
    outputs(6642) <= a xor b;
    outputs(6643) <= b and not a;
    outputs(6644) <= not a;
    outputs(6645) <= not a;
    outputs(6646) <= not (a or b);
    outputs(6647) <= not (a or b);
    outputs(6648) <= not a or b;
    outputs(6649) <= not a or b;
    outputs(6650) <= not (a and b);
    outputs(6651) <= b;
    outputs(6652) <= a;
    outputs(6653) <= b;
    outputs(6654) <= not (a xor b);
    outputs(6655) <= not a;
    outputs(6656) <= not a;
    outputs(6657) <= b and not a;
    outputs(6658) <= not b;
    outputs(6659) <= not (a or b);
    outputs(6660) <= b;
    outputs(6661) <= a xor b;
    outputs(6662) <= a or b;
    outputs(6663) <= a;
    outputs(6664) <= b and not a;
    outputs(6665) <= b;
    outputs(6666) <= not (a xor b);
    outputs(6667) <= a;
    outputs(6668) <= a xor b;
    outputs(6669) <= not a;
    outputs(6670) <= a and not b;
    outputs(6671) <= not (a or b);
    outputs(6672) <= not (a xor b);
    outputs(6673) <= a xor b;
    outputs(6674) <= a xor b;
    outputs(6675) <= a;
    outputs(6676) <= not (a xor b);
    outputs(6677) <= not b;
    outputs(6678) <= not b;
    outputs(6679) <= not (a xor b);
    outputs(6680) <= not a;
    outputs(6681) <= not a or b;
    outputs(6682) <= not a;
    outputs(6683) <= not (a xor b);
    outputs(6684) <= not b;
    outputs(6685) <= not a;
    outputs(6686) <= b and not a;
    outputs(6687) <= a and b;
    outputs(6688) <= a xor b;
    outputs(6689) <= a;
    outputs(6690) <= b and not a;
    outputs(6691) <= b and not a;
    outputs(6692) <= not a;
    outputs(6693) <= a;
    outputs(6694) <= not (a or b);
    outputs(6695) <= not b;
    outputs(6696) <= not (a xor b);
    outputs(6697) <= not b;
    outputs(6698) <= not b;
    outputs(6699) <= not b;
    outputs(6700) <= a and not b;
    outputs(6701) <= not b or a;
    outputs(6702) <= a xor b;
    outputs(6703) <= not b;
    outputs(6704) <= not (a xor b);
    outputs(6705) <= b;
    outputs(6706) <= not b or a;
    outputs(6707) <= not b;
    outputs(6708) <= a and not b;
    outputs(6709) <= not b or a;
    outputs(6710) <= not b;
    outputs(6711) <= a xor b;
    outputs(6712) <= b;
    outputs(6713) <= b and not a;
    outputs(6714) <= a and b;
    outputs(6715) <= not (a xor b);
    outputs(6716) <= a;
    outputs(6717) <= not (a or b);
    outputs(6718) <= a;
    outputs(6719) <= not a;
    outputs(6720) <= not a;
    outputs(6721) <= b;
    outputs(6722) <= a;
    outputs(6723) <= not a;
    outputs(6724) <= not (a and b);
    outputs(6725) <= not (a or b);
    outputs(6726) <= a;
    outputs(6727) <= not a or b;
    outputs(6728) <= a xor b;
    outputs(6729) <= a xor b;
    outputs(6730) <= a;
    outputs(6731) <= a xor b;
    outputs(6732) <= not b or a;
    outputs(6733) <= a xor b;
    outputs(6734) <= not b or a;
    outputs(6735) <= a xor b;
    outputs(6736) <= a;
    outputs(6737) <= not (a or b);
    outputs(6738) <= a xor b;
    outputs(6739) <= a;
    outputs(6740) <= a xor b;
    outputs(6741) <= not a or b;
    outputs(6742) <= not (a xor b);
    outputs(6743) <= a xor b;
    outputs(6744) <= not a;
    outputs(6745) <= not (a xor b);
    outputs(6746) <= not (a and b);
    outputs(6747) <= not (a and b);
    outputs(6748) <= a xor b;
    outputs(6749) <= not (a and b);
    outputs(6750) <= not (a xor b);
    outputs(6751) <= not (a xor b);
    outputs(6752) <= not a or b;
    outputs(6753) <= b and not a;
    outputs(6754) <= b;
    outputs(6755) <= not a;
    outputs(6756) <= not (a or b);
    outputs(6757) <= a xor b;
    outputs(6758) <= not a or b;
    outputs(6759) <= not (a or b);
    outputs(6760) <= a xor b;
    outputs(6761) <= not a or b;
    outputs(6762) <= a or b;
    outputs(6763) <= a xor b;
    outputs(6764) <= a xor b;
    outputs(6765) <= not (a xor b);
    outputs(6766) <= a;
    outputs(6767) <= not a;
    outputs(6768) <= not b or a;
    outputs(6769) <= not (a or b);
    outputs(6770) <= a or b;
    outputs(6771) <= not a;
    outputs(6772) <= not b;
    outputs(6773) <= not a;
    outputs(6774) <= b;
    outputs(6775) <= not (a xor b);
    outputs(6776) <= a xor b;
    outputs(6777) <= not a;
    outputs(6778) <= a or b;
    outputs(6779) <= not a;
    outputs(6780) <= a;
    outputs(6781) <= a xor b;
    outputs(6782) <= a and not b;
    outputs(6783) <= b;
    outputs(6784) <= not (a xor b);
    outputs(6785) <= not a;
    outputs(6786) <= a xor b;
    outputs(6787) <= a xor b;
    outputs(6788) <= a xor b;
    outputs(6789) <= not a or b;
    outputs(6790) <= not b;
    outputs(6791) <= not (a xor b);
    outputs(6792) <= not (a or b);
    outputs(6793) <= a xor b;
    outputs(6794) <= not b;
    outputs(6795) <= a;
    outputs(6796) <= not (a xor b);
    outputs(6797) <= not (a xor b);
    outputs(6798) <= not b;
    outputs(6799) <= b and not a;
    outputs(6800) <= a xor b;
    outputs(6801) <= not b;
    outputs(6802) <= not b;
    outputs(6803) <= a xor b;
    outputs(6804) <= b;
    outputs(6805) <= not (a xor b);
    outputs(6806) <= not (a xor b);
    outputs(6807) <= not a or b;
    outputs(6808) <= b;
    outputs(6809) <= a xor b;
    outputs(6810) <= not (a or b);
    outputs(6811) <= not b or a;
    outputs(6812) <= not (a xor b);
    outputs(6813) <= a or b;
    outputs(6814) <= not a;
    outputs(6815) <= not a;
    outputs(6816) <= not b or a;
    outputs(6817) <= not a;
    outputs(6818) <= not (a xor b);
    outputs(6819) <= a;
    outputs(6820) <= not (a xor b);
    outputs(6821) <= a and not b;
    outputs(6822) <= not a or b;
    outputs(6823) <= not (a xor b);
    outputs(6824) <= not b or a;
    outputs(6825) <= not a;
    outputs(6826) <= a;
    outputs(6827) <= not (a xor b);
    outputs(6828) <= a xor b;
    outputs(6829) <= not a;
    outputs(6830) <= a xor b;
    outputs(6831) <= a;
    outputs(6832) <= not (a xor b);
    outputs(6833) <= not (a xor b);
    outputs(6834) <= a xor b;
    outputs(6835) <= not (a xor b);
    outputs(6836) <= a;
    outputs(6837) <= a xor b;
    outputs(6838) <= not (a xor b);
    outputs(6839) <= not (a or b);
    outputs(6840) <= a xor b;
    outputs(6841) <= a xor b;
    outputs(6842) <= not (a xor b);
    outputs(6843) <= a;
    outputs(6844) <= not a;
    outputs(6845) <= not b;
    outputs(6846) <= a;
    outputs(6847) <= a;
    outputs(6848) <= not (a xor b);
    outputs(6849) <= b and not a;
    outputs(6850) <= a or b;
    outputs(6851) <= not b;
    outputs(6852) <= a;
    outputs(6853) <= a or b;
    outputs(6854) <= a;
    outputs(6855) <= a xor b;
    outputs(6856) <= a xor b;
    outputs(6857) <= not b;
    outputs(6858) <= b;
    outputs(6859) <= not (a xor b);
    outputs(6860) <= not a;
    outputs(6861) <= not (a and b);
    outputs(6862) <= not b;
    outputs(6863) <= not b;
    outputs(6864) <= a xor b;
    outputs(6865) <= b and not a;
    outputs(6866) <= not (a xor b);
    outputs(6867) <= not a;
    outputs(6868) <= not (a and b);
    outputs(6869) <= b;
    outputs(6870) <= b;
    outputs(6871) <= a;
    outputs(6872) <= a or b;
    outputs(6873) <= not b;
    outputs(6874) <= a xor b;
    outputs(6875) <= not b;
    outputs(6876) <= a and not b;
    outputs(6877) <= not (a or b);
    outputs(6878) <= b and not a;
    outputs(6879) <= not b;
    outputs(6880) <= a and b;
    outputs(6881) <= a or b;
    outputs(6882) <= not (a or b);
    outputs(6883) <= a xor b;
    outputs(6884) <= not a;
    outputs(6885) <= not (a xor b);
    outputs(6886) <= a;
    outputs(6887) <= not a;
    outputs(6888) <= a xor b;
    outputs(6889) <= a xor b;
    outputs(6890) <= a or b;
    outputs(6891) <= not (a xor b);
    outputs(6892) <= not a;
    outputs(6893) <= not (a or b);
    outputs(6894) <= a xor b;
    outputs(6895) <= not (a and b);
    outputs(6896) <= b;
    outputs(6897) <= a xor b;
    outputs(6898) <= a;
    outputs(6899) <= not (a xor b);
    outputs(6900) <= not b;
    outputs(6901) <= not a;
    outputs(6902) <= a xor b;
    outputs(6903) <= not (a xor b);
    outputs(6904) <= a xor b;
    outputs(6905) <= b;
    outputs(6906) <= a xor b;
    outputs(6907) <= not (a xor b);
    outputs(6908) <= b and not a;
    outputs(6909) <= not b;
    outputs(6910) <= not (a xor b);
    outputs(6911) <= not (a xor b);
    outputs(6912) <= not b;
    outputs(6913) <= not (a xor b);
    outputs(6914) <= b;
    outputs(6915) <= not (a xor b);
    outputs(6916) <= a and not b;
    outputs(6917) <= a;
    outputs(6918) <= '1';
    outputs(6919) <= not (a or b);
    outputs(6920) <= not b;
    outputs(6921) <= not (a xor b);
    outputs(6922) <= not a;
    outputs(6923) <= not (a or b);
    outputs(6924) <= b;
    outputs(6925) <= a;
    outputs(6926) <= a;
    outputs(6927) <= not a;
    outputs(6928) <= a and b;
    outputs(6929) <= b;
    outputs(6930) <= a and not b;
    outputs(6931) <= not a or b;
    outputs(6932) <= a and not b;
    outputs(6933) <= b and not a;
    outputs(6934) <= not (a xor b);
    outputs(6935) <= a xor b;
    outputs(6936) <= not a;
    outputs(6937) <= not b;
    outputs(6938) <= not (a xor b);
    outputs(6939) <= b;
    outputs(6940) <= not (a xor b);
    outputs(6941) <= a xor b;
    outputs(6942) <= not a;
    outputs(6943) <= not (a xor b);
    outputs(6944) <= b;
    outputs(6945) <= a and not b;
    outputs(6946) <= not b or a;
    outputs(6947) <= a xor b;
    outputs(6948) <= not a or b;
    outputs(6949) <= a;
    outputs(6950) <= not (a xor b);
    outputs(6951) <= a xor b;
    outputs(6952) <= a xor b;
    outputs(6953) <= not b;
    outputs(6954) <= b;
    outputs(6955) <= not b;
    outputs(6956) <= not (a or b);
    outputs(6957) <= b;
    outputs(6958) <= a xor b;
    outputs(6959) <= not (a xor b);
    outputs(6960) <= not b;
    outputs(6961) <= not a;
    outputs(6962) <= b and not a;
    outputs(6963) <= not a;
    outputs(6964) <= b and not a;
    outputs(6965) <= not b;
    outputs(6966) <= a and not b;
    outputs(6967) <= not a;
    outputs(6968) <= a and b;
    outputs(6969) <= b;
    outputs(6970) <= a;
    outputs(6971) <= not (a xor b);
    outputs(6972) <= not b;
    outputs(6973) <= not (a xor b);
    outputs(6974) <= not (a or b);
    outputs(6975) <= not (a xor b);
    outputs(6976) <= a xor b;
    outputs(6977) <= not (a xor b);
    outputs(6978) <= a and not b;
    outputs(6979) <= not b or a;
    outputs(6980) <= b and not a;
    outputs(6981) <= not (a xor b);
    outputs(6982) <= not a;
    outputs(6983) <= a and not b;
    outputs(6984) <= not (a xor b);
    outputs(6985) <= a or b;
    outputs(6986) <= a xor b;
    outputs(6987) <= b;
    outputs(6988) <= not b;
    outputs(6989) <= not b;
    outputs(6990) <= not b;
    outputs(6991) <= b;
    outputs(6992) <= a or b;
    outputs(6993) <= not a;
    outputs(6994) <= not (a or b);
    outputs(6995) <= b;
    outputs(6996) <= not b;
    outputs(6997) <= a;
    outputs(6998) <= a;
    outputs(6999) <= not b or a;
    outputs(7000) <= a;
    outputs(7001) <= not (a xor b);
    outputs(7002) <= not a;
    outputs(7003) <= a;
    outputs(7004) <= not (a or b);
    outputs(7005) <= not (a or b);
    outputs(7006) <= b;
    outputs(7007) <= a and b;
    outputs(7008) <= a;
    outputs(7009) <= b and not a;
    outputs(7010) <= a xor b;
    outputs(7011) <= b;
    outputs(7012) <= b;
    outputs(7013) <= a;
    outputs(7014) <= not (a xor b);
    outputs(7015) <= a;
    outputs(7016) <= not (a xor b);
    outputs(7017) <= a xor b;
    outputs(7018) <= not b;
    outputs(7019) <= not (a xor b);
    outputs(7020) <= a xor b;
    outputs(7021) <= not (a xor b);
    outputs(7022) <= b;
    outputs(7023) <= b and not a;
    outputs(7024) <= b;
    outputs(7025) <= not a or b;
    outputs(7026) <= a and not b;
    outputs(7027) <= not a;
    outputs(7028) <= a;
    outputs(7029) <= b and not a;
    outputs(7030) <= not b;
    outputs(7031) <= b;
    outputs(7032) <= not a;
    outputs(7033) <= a xor b;
    outputs(7034) <= b;
    outputs(7035) <= a and b;
    outputs(7036) <= a and not b;
    outputs(7037) <= not (a xor b);
    outputs(7038) <= not a or b;
    outputs(7039) <= a;
    outputs(7040) <= not a;
    outputs(7041) <= b;
    outputs(7042) <= a and not b;
    outputs(7043) <= not b;
    outputs(7044) <= a;
    outputs(7045) <= not a or b;
    outputs(7046) <= b;
    outputs(7047) <= not b;
    outputs(7048) <= a or b;
    outputs(7049) <= a or b;
    outputs(7050) <= a xor b;
    outputs(7051) <= not (a xor b);
    outputs(7052) <= not (a or b);
    outputs(7053) <= a xor b;
    outputs(7054) <= b;
    outputs(7055) <= not (a xor b);
    outputs(7056) <= a and b;
    outputs(7057) <= a xor b;
    outputs(7058) <= not (a xor b);
    outputs(7059) <= not a;
    outputs(7060) <= b and not a;
    outputs(7061) <= a and not b;
    outputs(7062) <= not b;
    outputs(7063) <= a or b;
    outputs(7064) <= not b;
    outputs(7065) <= a xor b;
    outputs(7066) <= not a or b;
    outputs(7067) <= a or b;
    outputs(7068) <= a xor b;
    outputs(7069) <= a and not b;
    outputs(7070) <= a or b;
    outputs(7071) <= not a or b;
    outputs(7072) <= a xor b;
    outputs(7073) <= not b or a;
    outputs(7074) <= not a or b;
    outputs(7075) <= not a;
    outputs(7076) <= not (a or b);
    outputs(7077) <= not (a xor b);
    outputs(7078) <= a xor b;
    outputs(7079) <= b;
    outputs(7080) <= not (a or b);
    outputs(7081) <= not (a xor b);
    outputs(7082) <= a and b;
    outputs(7083) <= b;
    outputs(7084) <= not b;
    outputs(7085) <= a;
    outputs(7086) <= a xor b;
    outputs(7087) <= not a;
    outputs(7088) <= b;
    outputs(7089) <= not (a xor b);
    outputs(7090) <= a;
    outputs(7091) <= not (a xor b);
    outputs(7092) <= not (a xor b);
    outputs(7093) <= a;
    outputs(7094) <= a xor b;
    outputs(7095) <= a;
    outputs(7096) <= not (a and b);
    outputs(7097) <= a;
    outputs(7098) <= a and b;
    outputs(7099) <= not (a xor b);
    outputs(7100) <= not b;
    outputs(7101) <= a and b;
    outputs(7102) <= not a;
    outputs(7103) <= a xor b;
    outputs(7104) <= a xor b;
    outputs(7105) <= a;
    outputs(7106) <= b;
    outputs(7107) <= a xor b;
    outputs(7108) <= not (a xor b);
    outputs(7109) <= a;
    outputs(7110) <= b;
    outputs(7111) <= a xor b;
    outputs(7112) <= not a;
    outputs(7113) <= a and b;
    outputs(7114) <= a and b;
    outputs(7115) <= not b;
    outputs(7116) <= not a;
    outputs(7117) <= not b;
    outputs(7118) <= a or b;
    outputs(7119) <= a;
    outputs(7120) <= b;
    outputs(7121) <= b;
    outputs(7122) <= b;
    outputs(7123) <= not b;
    outputs(7124) <= b;
    outputs(7125) <= a xor b;
    outputs(7126) <= not (a or b);
    outputs(7127) <= b;
    outputs(7128) <= not a;
    outputs(7129) <= not b;
    outputs(7130) <= b;
    outputs(7131) <= b;
    outputs(7132) <= not b or a;
    outputs(7133) <= not a;
    outputs(7134) <= not b;
    outputs(7135) <= a xor b;
    outputs(7136) <= a xor b;
    outputs(7137) <= b;
    outputs(7138) <= not (a xor b);
    outputs(7139) <= not a;
    outputs(7140) <= not a;
    outputs(7141) <= not a;
    outputs(7142) <= a and b;
    outputs(7143) <= not (a and b);
    outputs(7144) <= not a or b;
    outputs(7145) <= not (a xor b);
    outputs(7146) <= not a;
    outputs(7147) <= a xor b;
    outputs(7148) <= not a;
    outputs(7149) <= a;
    outputs(7150) <= not (a xor b);
    outputs(7151) <= not a;
    outputs(7152) <= a and not b;
    outputs(7153) <= a xor b;
    outputs(7154) <= a xor b;
    outputs(7155) <= not (a xor b);
    outputs(7156) <= b;
    outputs(7157) <= not a or b;
    outputs(7158) <= a and not b;
    outputs(7159) <= not (a xor b);
    outputs(7160) <= a xor b;
    outputs(7161) <= not (a and b);
    outputs(7162) <= not (a xor b);
    outputs(7163) <= not b;
    outputs(7164) <= b;
    outputs(7165) <= b and not a;
    outputs(7166) <= b;
    outputs(7167) <= b;
    outputs(7168) <= not (a xor b);
    outputs(7169) <= not (a and b);
    outputs(7170) <= not a;
    outputs(7171) <= not a or b;
    outputs(7172) <= not (a xor b);
    outputs(7173) <= b;
    outputs(7174) <= not b;
    outputs(7175) <= not (a or b);
    outputs(7176) <= not b;
    outputs(7177) <= not (a or b);
    outputs(7178) <= not (a or b);
    outputs(7179) <= a;
    outputs(7180) <= a;
    outputs(7181) <= not (a xor b);
    outputs(7182) <= a or b;
    outputs(7183) <= b;
    outputs(7184) <= not (a xor b);
    outputs(7185) <= a;
    outputs(7186) <= a xor b;
    outputs(7187) <= not (a xor b);
    outputs(7188) <= not a;
    outputs(7189) <= not (a or b);
    outputs(7190) <= not a;
    outputs(7191) <= a xor b;
    outputs(7192) <= a xor b;
    outputs(7193) <= not (a xor b);
    outputs(7194) <= not (a xor b);
    outputs(7195) <= a xor b;
    outputs(7196) <= not (a or b);
    outputs(7197) <= not a;
    outputs(7198) <= not a;
    outputs(7199) <= a xor b;
    outputs(7200) <= not (a xor b);
    outputs(7201) <= b;
    outputs(7202) <= not b;
    outputs(7203) <= a xor b;
    outputs(7204) <= a xor b;
    outputs(7205) <= not a;
    outputs(7206) <= a;
    outputs(7207) <= not b;
    outputs(7208) <= not (a and b);
    outputs(7209) <= not a;
    outputs(7210) <= not (a xor b);
    outputs(7211) <= a xor b;
    outputs(7212) <= b;
    outputs(7213) <= not a;
    outputs(7214) <= b;
    outputs(7215) <= not b or a;
    outputs(7216) <= a or b;
    outputs(7217) <= a and b;
    outputs(7218) <= a xor b;
    outputs(7219) <= b and not a;
    outputs(7220) <= a xor b;
    outputs(7221) <= not b;
    outputs(7222) <= a xor b;
    outputs(7223) <= not a;
    outputs(7224) <= a xor b;
    outputs(7225) <= not b;
    outputs(7226) <= not (a or b);
    outputs(7227) <= a and b;
    outputs(7228) <= b and not a;
    outputs(7229) <= a xor b;
    outputs(7230) <= not (a xor b);
    outputs(7231) <= not (a xor b);
    outputs(7232) <= a;
    outputs(7233) <= not b;
    outputs(7234) <= a;
    outputs(7235) <= not (a or b);
    outputs(7236) <= a xor b;
    outputs(7237) <= not a;
    outputs(7238) <= not (a and b);
    outputs(7239) <= not a;
    outputs(7240) <= not a;
    outputs(7241) <= a;
    outputs(7242) <= b;
    outputs(7243) <= a and b;
    outputs(7244) <= a xor b;
    outputs(7245) <= not b;
    outputs(7246) <= a;
    outputs(7247) <= b and not a;
    outputs(7248) <= a xor b;
    outputs(7249) <= a and b;
    outputs(7250) <= b and not a;
    outputs(7251) <= a xor b;
    outputs(7252) <= a and b;
    outputs(7253) <= not b;
    outputs(7254) <= not (a xor b);
    outputs(7255) <= not (a xor b);
    outputs(7256) <= not b;
    outputs(7257) <= b and not a;
    outputs(7258) <= not a;
    outputs(7259) <= a and not b;
    outputs(7260) <= not (a xor b);
    outputs(7261) <= not a;
    outputs(7262) <= a xor b;
    outputs(7263) <= not a;
    outputs(7264) <= a xor b;
    outputs(7265) <= b;
    outputs(7266) <= b;
    outputs(7267) <= a xor b;
    outputs(7268) <= a xor b;
    outputs(7269) <= not a;
    outputs(7270) <= b;
    outputs(7271) <= a;
    outputs(7272) <= not (a xor b);
    outputs(7273) <= a xor b;
    outputs(7274) <= a and not b;
    outputs(7275) <= not (a or b);
    outputs(7276) <= a;
    outputs(7277) <= not (a or b);
    outputs(7278) <= not b;
    outputs(7279) <= a xor b;
    outputs(7280) <= not (a and b);
    outputs(7281) <= not a;
    outputs(7282) <= b and not a;
    outputs(7283) <= a and b;
    outputs(7284) <= a xor b;
    outputs(7285) <= not a;
    outputs(7286) <= a;
    outputs(7287) <= not (a xor b);
    outputs(7288) <= a xor b;
    outputs(7289) <= not a;
    outputs(7290) <= not a;
    outputs(7291) <= b and not a;
    outputs(7292) <= not (a xor b);
    outputs(7293) <= a xor b;
    outputs(7294) <= not a;
    outputs(7295) <= not (a xor b);
    outputs(7296) <= b;
    outputs(7297) <= not (a xor b);
    outputs(7298) <= not b;
    outputs(7299) <= not (a and b);
    outputs(7300) <= a xor b;
    outputs(7301) <= not b;
    outputs(7302) <= a;
    outputs(7303) <= a and not b;
    outputs(7304) <= not a;
    outputs(7305) <= b;
    outputs(7306) <= b;
    outputs(7307) <= a xor b;
    outputs(7308) <= not a;
    outputs(7309) <= a xor b;
    outputs(7310) <= a;
    outputs(7311) <= not (a xor b);
    outputs(7312) <= not (a xor b);
    outputs(7313) <= not a;
    outputs(7314) <= b;
    outputs(7315) <= a xor b;
    outputs(7316) <= not a;
    outputs(7317) <= not (a xor b);
    outputs(7318) <= not b;
    outputs(7319) <= not b;
    outputs(7320) <= not a;
    outputs(7321) <= b;
    outputs(7322) <= not (a or b);
    outputs(7323) <= b and not a;
    outputs(7324) <= a or b;
    outputs(7325) <= not (a xor b);
    outputs(7326) <= not (a and b);
    outputs(7327) <= not (a xor b);
    outputs(7328) <= not (a xor b);
    outputs(7329) <= a xor b;
    outputs(7330) <= a and b;
    outputs(7331) <= not b;
    outputs(7332) <= not (a xor b);
    outputs(7333) <= not a;
    outputs(7334) <= b;
    outputs(7335) <= a;
    outputs(7336) <= not (a xor b);
    outputs(7337) <= not (a xor b);
    outputs(7338) <= a and not b;
    outputs(7339) <= not (a xor b);
    outputs(7340) <= not (a xor b);
    outputs(7341) <= b;
    outputs(7342) <= not b;
    outputs(7343) <= not b;
    outputs(7344) <= a;
    outputs(7345) <= b;
    outputs(7346) <= a xor b;
    outputs(7347) <= a xor b;
    outputs(7348) <= not (a xor b);
    outputs(7349) <= a;
    outputs(7350) <= a xor b;
    outputs(7351) <= a xor b;
    outputs(7352) <= a xor b;
    outputs(7353) <= a xor b;
    outputs(7354) <= not a;
    outputs(7355) <= not (a xor b);
    outputs(7356) <= not a or b;
    outputs(7357) <= not (a xor b);
    outputs(7358) <= b;
    outputs(7359) <= not a;
    outputs(7360) <= not b;
    outputs(7361) <= not a;
    outputs(7362) <= not (a or b);
    outputs(7363) <= not a;
    outputs(7364) <= not a;
    outputs(7365) <= a xor b;
    outputs(7366) <= a and not b;
    outputs(7367) <= a xor b;
    outputs(7368) <= a xor b;
    outputs(7369) <= a or b;
    outputs(7370) <= b;
    outputs(7371) <= a;
    outputs(7372) <= b;
    outputs(7373) <= not b;
    outputs(7374) <= a and not b;
    outputs(7375) <= a;
    outputs(7376) <= not (a xor b);
    outputs(7377) <= a;
    outputs(7378) <= a and b;
    outputs(7379) <= a;
    outputs(7380) <= b;
    outputs(7381) <= a and b;
    outputs(7382) <= b and not a;
    outputs(7383) <= not b;
    outputs(7384) <= not b;
    outputs(7385) <= b;
    outputs(7386) <= not (a and b);
    outputs(7387) <= not (a xor b);
    outputs(7388) <= a and not b;
    outputs(7389) <= not (a and b);
    outputs(7390) <= b;
    outputs(7391) <= a or b;
    outputs(7392) <= b and not a;
    outputs(7393) <= not b;
    outputs(7394) <= not (a xor b);
    outputs(7395) <= a;
    outputs(7396) <= b;
    outputs(7397) <= not (a xor b);
    outputs(7398) <= a;
    outputs(7399) <= not b;
    outputs(7400) <= not a;
    outputs(7401) <= not (a xor b);
    outputs(7402) <= a xor b;
    outputs(7403) <= not a;
    outputs(7404) <= a xor b;
    outputs(7405) <= a xor b;
    outputs(7406) <= a;
    outputs(7407) <= a or b;
    outputs(7408) <= a and not b;
    outputs(7409) <= not (a xor b);
    outputs(7410) <= not b;
    outputs(7411) <= b and not a;
    outputs(7412) <= b;
    outputs(7413) <= b;
    outputs(7414) <= a xor b;
    outputs(7415) <= not (a xor b);
    outputs(7416) <= not (a xor b);
    outputs(7417) <= not b;
    outputs(7418) <= not b;
    outputs(7419) <= not a;
    outputs(7420) <= not (a xor b);
    outputs(7421) <= a xor b;
    outputs(7422) <= a and not b;
    outputs(7423) <= not a;
    outputs(7424) <= a;
    outputs(7425) <= not b;
    outputs(7426) <= not b;
    outputs(7427) <= a xor b;
    outputs(7428) <= not a;
    outputs(7429) <= a xor b;
    outputs(7430) <= not (a or b);
    outputs(7431) <= a xor b;
    outputs(7432) <= b and not a;
    outputs(7433) <= not (a and b);
    outputs(7434) <= not a;
    outputs(7435) <= not (a and b);
    outputs(7436) <= b;
    outputs(7437) <= not a or b;
    outputs(7438) <= b;
    outputs(7439) <= b;
    outputs(7440) <= b and not a;
    outputs(7441) <= a or b;
    outputs(7442) <= not b;
    outputs(7443) <= b;
    outputs(7444) <= not b;
    outputs(7445) <= not a or b;
    outputs(7446) <= not a;
    outputs(7447) <= a xor b;
    outputs(7448) <= a;
    outputs(7449) <= not (a xor b);
    outputs(7450) <= a;
    outputs(7451) <= b and not a;
    outputs(7452) <= not (a xor b);
    outputs(7453) <= not (a xor b);
    outputs(7454) <= not b;
    outputs(7455) <= a;
    outputs(7456) <= not (a xor b);
    outputs(7457) <= a;
    outputs(7458) <= a;
    outputs(7459) <= a;
    outputs(7460) <= not (a xor b);
    outputs(7461) <= a xor b;
    outputs(7462) <= not a;
    outputs(7463) <= b;
    outputs(7464) <= a and b;
    outputs(7465) <= not a;
    outputs(7466) <= b and not a;
    outputs(7467) <= not a or b;
    outputs(7468) <= not b;
    outputs(7469) <= not b;
    outputs(7470) <= not (a xor b);
    outputs(7471) <= not b;
    outputs(7472) <= a;
    outputs(7473) <= not (a and b);
    outputs(7474) <= not (a xor b);
    outputs(7475) <= not b or a;
    outputs(7476) <= not (a xor b);
    outputs(7477) <= not a;
    outputs(7478) <= not (a xor b);
    outputs(7479) <= not a or b;
    outputs(7480) <= not (a xor b);
    outputs(7481) <= a xor b;
    outputs(7482) <= not a;
    outputs(7483) <= a xor b;
    outputs(7484) <= not b or a;
    outputs(7485) <= a xor b;
    outputs(7486) <= a and b;
    outputs(7487) <= a xor b;
    outputs(7488) <= a xor b;
    outputs(7489) <= not a;
    outputs(7490) <= a or b;
    outputs(7491) <= not (a xor b);
    outputs(7492) <= a and b;
    outputs(7493) <= not a;
    outputs(7494) <= not b;
    outputs(7495) <= not (a xor b);
    outputs(7496) <= not a;
    outputs(7497) <= a and not b;
    outputs(7498) <= a xor b;
    outputs(7499) <= a and not b;
    outputs(7500) <= not b;
    outputs(7501) <= a xor b;
    outputs(7502) <= a xor b;
    outputs(7503) <= not b;
    outputs(7504) <= not b or a;
    outputs(7505) <= a and not b;
    outputs(7506) <= b;
    outputs(7507) <= not (a xor b);
    outputs(7508) <= not b;
    outputs(7509) <= not a;
    outputs(7510) <= a and not b;
    outputs(7511) <= not (a or b);
    outputs(7512) <= not a;
    outputs(7513) <= not (a xor b);
    outputs(7514) <= b;
    outputs(7515) <= a;
    outputs(7516) <= b and not a;
    outputs(7517) <= a xor b;
    outputs(7518) <= not (a or b);
    outputs(7519) <= not a;
    outputs(7520) <= not a;
    outputs(7521) <= a or b;
    outputs(7522) <= b;
    outputs(7523) <= a and b;
    outputs(7524) <= not b;
    outputs(7525) <= a and b;
    outputs(7526) <= not (a xor b);
    outputs(7527) <= not (a xor b);
    outputs(7528) <= not (a or b);
    outputs(7529) <= not (a xor b);
    outputs(7530) <= a xor b;
    outputs(7531) <= not b or a;
    outputs(7532) <= not (a xor b);
    outputs(7533) <= not b or a;
    outputs(7534) <= b;
    outputs(7535) <= a xor b;
    outputs(7536) <= a and not b;
    outputs(7537) <= a xor b;
    outputs(7538) <= a xor b;
    outputs(7539) <= a xor b;
    outputs(7540) <= b;
    outputs(7541) <= a xor b;
    outputs(7542) <= a xor b;
    outputs(7543) <= b and not a;
    outputs(7544) <= a and not b;
    outputs(7545) <= not (a or b);
    outputs(7546) <= not b;
    outputs(7547) <= a xor b;
    outputs(7548) <= a;
    outputs(7549) <= b and not a;
    outputs(7550) <= a and b;
    outputs(7551) <= a and not b;
    outputs(7552) <= not (a or b);
    outputs(7553) <= a xor b;
    outputs(7554) <= not (a and b);
    outputs(7555) <= a;
    outputs(7556) <= not (a or b);
    outputs(7557) <= not b;
    outputs(7558) <= b;
    outputs(7559) <= b and not a;
    outputs(7560) <= b and not a;
    outputs(7561) <= not (a or b);
    outputs(7562) <= not (a xor b);
    outputs(7563) <= a or b;
    outputs(7564) <= not b;
    outputs(7565) <= not (a xor b);
    outputs(7566) <= not (a xor b);
    outputs(7567) <= not b;
    outputs(7568) <= a and b;
    outputs(7569) <= not a;
    outputs(7570) <= not a;
    outputs(7571) <= a xor b;
    outputs(7572) <= a and b;
    outputs(7573) <= not (a xor b);
    outputs(7574) <= not a;
    outputs(7575) <= not (a xor b);
    outputs(7576) <= not b;
    outputs(7577) <= a;
    outputs(7578) <= '1';
    outputs(7579) <= b;
    outputs(7580) <= not (a xor b);
    outputs(7581) <= not (a xor b);
    outputs(7582) <= not (a xor b);
    outputs(7583) <= a;
    outputs(7584) <= not b;
    outputs(7585) <= a xor b;
    outputs(7586) <= not b;
    outputs(7587) <= not (a and b);
    outputs(7588) <= a xor b;
    outputs(7589) <= not b;
    outputs(7590) <= a;
    outputs(7591) <= b;
    outputs(7592) <= a and b;
    outputs(7593) <= a and b;
    outputs(7594) <= a xor b;
    outputs(7595) <= not (a xor b);
    outputs(7596) <= a and not b;
    outputs(7597) <= not a;
    outputs(7598) <= a xor b;
    outputs(7599) <= not (a xor b);
    outputs(7600) <= a or b;
    outputs(7601) <= a xor b;
    outputs(7602) <= not (a xor b);
    outputs(7603) <= a and b;
    outputs(7604) <= not a;
    outputs(7605) <= not (a xor b);
    outputs(7606) <= not (a or b);
    outputs(7607) <= b;
    outputs(7608) <= b and not a;
    outputs(7609) <= b;
    outputs(7610) <= not b;
    outputs(7611) <= b and not a;
    outputs(7612) <= a;
    outputs(7613) <= a;
    outputs(7614) <= a or b;
    outputs(7615) <= not b;
    outputs(7616) <= not a;
    outputs(7617) <= b and not a;
    outputs(7618) <= a xor b;
    outputs(7619) <= a;
    outputs(7620) <= a xor b;
    outputs(7621) <= a xor b;
    outputs(7622) <= a;
    outputs(7623) <= not a;
    outputs(7624) <= not b;
    outputs(7625) <= not (a xor b);
    outputs(7626) <= not b;
    outputs(7627) <= not a;
    outputs(7628) <= not (a xor b);
    outputs(7629) <= not (a or b);
    outputs(7630) <= b and not a;
    outputs(7631) <= b;
    outputs(7632) <= not (a xor b);
    outputs(7633) <= not (a or b);
    outputs(7634) <= not b;
    outputs(7635) <= not (a xor b);
    outputs(7636) <= not (a xor b);
    outputs(7637) <= b;
    outputs(7638) <= a xor b;
    outputs(7639) <= not (a xor b);
    outputs(7640) <= not b;
    outputs(7641) <= not b;
    outputs(7642) <= not (a and b);
    outputs(7643) <= a xor b;
    outputs(7644) <= not a;
    outputs(7645) <= not (a xor b);
    outputs(7646) <= a xor b;
    outputs(7647) <= not (a xor b);
    outputs(7648) <= b;
    outputs(7649) <= not (a xor b);
    outputs(7650) <= not (a or b);
    outputs(7651) <= not (a or b);
    outputs(7652) <= b;
    outputs(7653) <= a and not b;
    outputs(7654) <= b;
    outputs(7655) <= not (a or b);
    outputs(7656) <= not a;
    outputs(7657) <= not b or a;
    outputs(7658) <= not (a xor b);
    outputs(7659) <= a and not b;
    outputs(7660) <= not b;
    outputs(7661) <= not (a xor b);
    outputs(7662) <= b;
    outputs(7663) <= not (a or b);
    outputs(7664) <= a and b;
    outputs(7665) <= a and b;
    outputs(7666) <= a;
    outputs(7667) <= not (a xor b);
    outputs(7668) <= b;
    outputs(7669) <= a xor b;
    outputs(7670) <= a xor b;
    outputs(7671) <= b;
    outputs(7672) <= a and not b;
    outputs(7673) <= b;
    outputs(7674) <= not (a xor b);
    outputs(7675) <= a;
    outputs(7676) <= a xor b;
    outputs(7677) <= not a;
    outputs(7678) <= a and not b;
    outputs(7679) <= b and not a;
end Behavioral;
