library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(2559 downto 0);
    signal layer1_outputs: std_logic_vector(2559 downto 0);
    signal layer2_outputs: std_logic_vector(2559 downto 0);

begin
    layer0_outputs(0) <= not b or a;
    layer0_outputs(1) <= not (a or b);
    layer0_outputs(2) <= not (a xor b);
    layer0_outputs(3) <= b and not a;
    layer0_outputs(4) <= not b or a;
    layer0_outputs(5) <= b and not a;
    layer0_outputs(6) <= 1'b0;
    layer0_outputs(7) <= b;
    layer0_outputs(8) <= not a or b;
    layer0_outputs(9) <= a and b;
    layer0_outputs(10) <= not (a or b);
    layer0_outputs(11) <= not b or a;
    layer0_outputs(12) <= 1'b1;
    layer0_outputs(13) <= a;
    layer0_outputs(14) <= not a;
    layer0_outputs(15) <= a and not b;
    layer0_outputs(16) <= not b or a;
    layer0_outputs(17) <= a xor b;
    layer0_outputs(18) <= a xor b;
    layer0_outputs(19) <= not (a or b);
    layer0_outputs(20) <= not (a or b);
    layer0_outputs(21) <= a and b;
    layer0_outputs(22) <= b and not a;
    layer0_outputs(23) <= not (a and b);
    layer0_outputs(24) <= 1'b1;
    layer0_outputs(25) <= not (a and b);
    layer0_outputs(26) <= b and not a;
    layer0_outputs(27) <= not (a or b);
    layer0_outputs(28) <= a or b;
    layer0_outputs(29) <= not a;
    layer0_outputs(30) <= b;
    layer0_outputs(31) <= not (a and b);
    layer0_outputs(32) <= not b;
    layer0_outputs(33) <= not b or a;
    layer0_outputs(34) <= not b;
    layer0_outputs(35) <= not (a or b);
    layer0_outputs(36) <= not (a xor b);
    layer0_outputs(37) <= 1'b0;
    layer0_outputs(38) <= not a or b;
    layer0_outputs(39) <= not b or a;
    layer0_outputs(40) <= not (a or b);
    layer0_outputs(41) <= not a or b;
    layer0_outputs(42) <= not b;
    layer0_outputs(43) <= not b or a;
    layer0_outputs(44) <= a or b;
    layer0_outputs(45) <= not a;
    layer0_outputs(46) <= not (a xor b);
    layer0_outputs(47) <= not a;
    layer0_outputs(48) <= not a;
    layer0_outputs(49) <= b;
    layer0_outputs(50) <= b and not a;
    layer0_outputs(51) <= 1'b0;
    layer0_outputs(52) <= not (a and b);
    layer0_outputs(53) <= not a;
    layer0_outputs(54) <= a and not b;
    layer0_outputs(55) <= a xor b;
    layer0_outputs(56) <= a or b;
    layer0_outputs(57) <= a or b;
    layer0_outputs(58) <= a;
    layer0_outputs(59) <= not a or b;
    layer0_outputs(60) <= not (a or b);
    layer0_outputs(61) <= b and not a;
    layer0_outputs(62) <= not (a xor b);
    layer0_outputs(63) <= 1'b1;
    layer0_outputs(64) <= not (a or b);
    layer0_outputs(65) <= 1'b0;
    layer0_outputs(66) <= a;
    layer0_outputs(67) <= b;
    layer0_outputs(68) <= a and b;
    layer0_outputs(69) <= not b or a;
    layer0_outputs(70) <= a and not b;
    layer0_outputs(71) <= not a;
    layer0_outputs(72) <= b and not a;
    layer0_outputs(73) <= a;
    layer0_outputs(74) <= a or b;
    layer0_outputs(75) <= a and not b;
    layer0_outputs(76) <= a or b;
    layer0_outputs(77) <= b and not a;
    layer0_outputs(78) <= not a;
    layer0_outputs(79) <= not a or b;
    layer0_outputs(80) <= b;
    layer0_outputs(81) <= a and not b;
    layer0_outputs(82) <= not (a or b);
    layer0_outputs(83) <= not a or b;
    layer0_outputs(84) <= a and not b;
    layer0_outputs(85) <= a xor b;
    layer0_outputs(86) <= not (a xor b);
    layer0_outputs(87) <= not a or b;
    layer0_outputs(88) <= not a;
    layer0_outputs(89) <= b and not a;
    layer0_outputs(90) <= a;
    layer0_outputs(91) <= a xor b;
    layer0_outputs(92) <= a and b;
    layer0_outputs(93) <= 1'b1;
    layer0_outputs(94) <= 1'b0;
    layer0_outputs(95) <= not (a xor b);
    layer0_outputs(96) <= a and not b;
    layer0_outputs(97) <= a xor b;
    layer0_outputs(98) <= not a or b;
    layer0_outputs(99) <= not a;
    layer0_outputs(100) <= not (a or b);
    layer0_outputs(101) <= a;
    layer0_outputs(102) <= a or b;
    layer0_outputs(103) <= b and not a;
    layer0_outputs(104) <= not b;
    layer0_outputs(105) <= not (a xor b);
    layer0_outputs(106) <= b;
    layer0_outputs(107) <= not a or b;
    layer0_outputs(108) <= a or b;
    layer0_outputs(109) <= not b;
    layer0_outputs(110) <= a or b;
    layer0_outputs(111) <= b and not a;
    layer0_outputs(112) <= not (a xor b);
    layer0_outputs(113) <= a or b;
    layer0_outputs(114) <= not b or a;
    layer0_outputs(115) <= not a;
    layer0_outputs(116) <= not (a xor b);
    layer0_outputs(117) <= a;
    layer0_outputs(118) <= not a;
    layer0_outputs(119) <= a and b;
    layer0_outputs(120) <= a and b;
    layer0_outputs(121) <= b and not a;
    layer0_outputs(122) <= b and not a;
    layer0_outputs(123) <= 1'b0;
    layer0_outputs(124) <= a;
    layer0_outputs(125) <= not b;
    layer0_outputs(126) <= not (a and b);
    layer0_outputs(127) <= a xor b;
    layer0_outputs(128) <= not (a xor b);
    layer0_outputs(129) <= a and b;
    layer0_outputs(130) <= 1'b0;
    layer0_outputs(131) <= not (a and b);
    layer0_outputs(132) <= not (a xor b);
    layer0_outputs(133) <= b;
    layer0_outputs(134) <= a or b;
    layer0_outputs(135) <= not (a xor b);
    layer0_outputs(136) <= not (a xor b);
    layer0_outputs(137) <= a xor b;
    layer0_outputs(138) <= not a;
    layer0_outputs(139) <= not b;
    layer0_outputs(140) <= not (a or b);
    layer0_outputs(141) <= not a or b;
    layer0_outputs(142) <= a;
    layer0_outputs(143) <= a or b;
    layer0_outputs(144) <= b;
    layer0_outputs(145) <= a or b;
    layer0_outputs(146) <= a and not b;
    layer0_outputs(147) <= not a or b;
    layer0_outputs(148) <= not a;
    layer0_outputs(149) <= not a;
    layer0_outputs(150) <= a;
    layer0_outputs(151) <= not a or b;
    layer0_outputs(152) <= a;
    layer0_outputs(153) <= b;
    layer0_outputs(154) <= 1'b1;
    layer0_outputs(155) <= not a or b;
    layer0_outputs(156) <= 1'b1;
    layer0_outputs(157) <= not (a or b);
    layer0_outputs(158) <= not a or b;
    layer0_outputs(159) <= not (a and b);
    layer0_outputs(160) <= a and not b;
    layer0_outputs(161) <= a xor b;
    layer0_outputs(162) <= b and not a;
    layer0_outputs(163) <= b;
    layer0_outputs(164) <= not (a or b);
    layer0_outputs(165) <= not (a xor b);
    layer0_outputs(166) <= not (a or b);
    layer0_outputs(167) <= not b;
    layer0_outputs(168) <= not b or a;
    layer0_outputs(169) <= a xor b;
    layer0_outputs(170) <= a or b;
    layer0_outputs(171) <= not (a and b);
    layer0_outputs(172) <= not b or a;
    layer0_outputs(173) <= not b;
    layer0_outputs(174) <= 1'b1;
    layer0_outputs(175) <= b and not a;
    layer0_outputs(176) <= a;
    layer0_outputs(177) <= a;
    layer0_outputs(178) <= a or b;
    layer0_outputs(179) <= b and not a;
    layer0_outputs(180) <= b and not a;
    layer0_outputs(181) <= not b;
    layer0_outputs(182) <= not (a or b);
    layer0_outputs(183) <= not (a or b);
    layer0_outputs(184) <= not b or a;
    layer0_outputs(185) <= a or b;
    layer0_outputs(186) <= not (a and b);
    layer0_outputs(187) <= a or b;
    layer0_outputs(188) <= b;
    layer0_outputs(189) <= b;
    layer0_outputs(190) <= 1'b1;
    layer0_outputs(191) <= a or b;
    layer0_outputs(192) <= not b;
    layer0_outputs(193) <= a or b;
    layer0_outputs(194) <= not a;
    layer0_outputs(195) <= not (a or b);
    layer0_outputs(196) <= a and b;
    layer0_outputs(197) <= not (a or b);
    layer0_outputs(198) <= a or b;
    layer0_outputs(199) <= a xor b;
    layer0_outputs(200) <= not a;
    layer0_outputs(201) <= b and not a;
    layer0_outputs(202) <= a xor b;
    layer0_outputs(203) <= a or b;
    layer0_outputs(204) <= a or b;
    layer0_outputs(205) <= not b;
    layer0_outputs(206) <= b;
    layer0_outputs(207) <= a;
    layer0_outputs(208) <= a or b;
    layer0_outputs(209) <= not b;
    layer0_outputs(210) <= not a or b;
    layer0_outputs(211) <= not a;
    layer0_outputs(212) <= a;
    layer0_outputs(213) <= not a;
    layer0_outputs(214) <= not (a xor b);
    layer0_outputs(215) <= not b;
    layer0_outputs(216) <= not b;
    layer0_outputs(217) <= b;
    layer0_outputs(218) <= a and not b;
    layer0_outputs(219) <= not (a or b);
    layer0_outputs(220) <= not (a and b);
    layer0_outputs(221) <= not a or b;
    layer0_outputs(222) <= a xor b;
    layer0_outputs(223) <= a and not b;
    layer0_outputs(224) <= b and not a;
    layer0_outputs(225) <= not a;
    layer0_outputs(226) <= a xor b;
    layer0_outputs(227) <= b;
    layer0_outputs(228) <= not (a and b);
    layer0_outputs(229) <= not b or a;
    layer0_outputs(230) <= not (a xor b);
    layer0_outputs(231) <= not b or a;
    layer0_outputs(232) <= not b or a;
    layer0_outputs(233) <= not b;
    layer0_outputs(234) <= b and not a;
    layer0_outputs(235) <= b and not a;
    layer0_outputs(236) <= 1'b0;
    layer0_outputs(237) <= not a or b;
    layer0_outputs(238) <= not a;
    layer0_outputs(239) <= a xor b;
    layer0_outputs(240) <= not b or a;
    layer0_outputs(241) <= b and not a;
    layer0_outputs(242) <= a or b;
    layer0_outputs(243) <= b;
    layer0_outputs(244) <= not (a or b);
    layer0_outputs(245) <= not b or a;
    layer0_outputs(246) <= not b or a;
    layer0_outputs(247) <= b;
    layer0_outputs(248) <= a and not b;
    layer0_outputs(249) <= a or b;
    layer0_outputs(250) <= not b;
    layer0_outputs(251) <= not a;
    layer0_outputs(252) <= not (a xor b);
    layer0_outputs(253) <= 1'b1;
    layer0_outputs(254) <= a or b;
    layer0_outputs(255) <= not (a and b);
    layer0_outputs(256) <= b and not a;
    layer0_outputs(257) <= not (a or b);
    layer0_outputs(258) <= a or b;
    layer0_outputs(259) <= not (a xor b);
    layer0_outputs(260) <= a xor b;
    layer0_outputs(261) <= not a or b;
    layer0_outputs(262) <= 1'b1;
    layer0_outputs(263) <= not a;
    layer0_outputs(264) <= not (a or b);
    layer0_outputs(265) <= 1'b0;
    layer0_outputs(266) <= b;
    layer0_outputs(267) <= a and not b;
    layer0_outputs(268) <= a and not b;
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= not (a or b);
    layer0_outputs(271) <= 1'b1;
    layer0_outputs(272) <= a or b;
    layer0_outputs(273) <= not a or b;
    layer0_outputs(274) <= a xor b;
    layer0_outputs(275) <= not a;
    layer0_outputs(276) <= 1'b1;
    layer0_outputs(277) <= 1'b1;
    layer0_outputs(278) <= not a or b;
    layer0_outputs(279) <= not a;
    layer0_outputs(280) <= not a;
    layer0_outputs(281) <= not b;
    layer0_outputs(282) <= b and not a;
    layer0_outputs(283) <= not b or a;
    layer0_outputs(284) <= 1'b0;
    layer0_outputs(285) <= b;
    layer0_outputs(286) <= a or b;
    layer0_outputs(287) <= a or b;
    layer0_outputs(288) <= b and not a;
    layer0_outputs(289) <= not (a or b);
    layer0_outputs(290) <= not (a and b);
    layer0_outputs(291) <= not (a or b);
    layer0_outputs(292) <= a or b;
    layer0_outputs(293) <= not a or b;
    layer0_outputs(294) <= not (a or b);
    layer0_outputs(295) <= not (a xor b);
    layer0_outputs(296) <= b;
    layer0_outputs(297) <= not (a xor b);
    layer0_outputs(298) <= not a;
    layer0_outputs(299) <= not (a or b);
    layer0_outputs(300) <= b;
    layer0_outputs(301) <= a or b;
    layer0_outputs(302) <= not b or a;
    layer0_outputs(303) <= a or b;
    layer0_outputs(304) <= a and not b;
    layer0_outputs(305) <= not a or b;
    layer0_outputs(306) <= not b;
    layer0_outputs(307) <= a or b;
    layer0_outputs(308) <= a;
    layer0_outputs(309) <= not a;
    layer0_outputs(310) <= a or b;
    layer0_outputs(311) <= b;
    layer0_outputs(312) <= a and not b;
    layer0_outputs(313) <= b and not a;
    layer0_outputs(314) <= a or b;
    layer0_outputs(315) <= not b;
    layer0_outputs(316) <= not (a or b);
    layer0_outputs(317) <= not (a xor b);
    layer0_outputs(318) <= b;
    layer0_outputs(319) <= a or b;
    layer0_outputs(320) <= not a;
    layer0_outputs(321) <= a or b;
    layer0_outputs(322) <= a and not b;
    layer0_outputs(323) <= not (a xor b);
    layer0_outputs(324) <= b and not a;
    layer0_outputs(325) <= not a or b;
    layer0_outputs(326) <= a and not b;
    layer0_outputs(327) <= not b or a;
    layer0_outputs(328) <= a and b;
    layer0_outputs(329) <= not b;
    layer0_outputs(330) <= not b or a;
    layer0_outputs(331) <= not b;
    layer0_outputs(332) <= b and not a;
    layer0_outputs(333) <= not a;
    layer0_outputs(334) <= not (a or b);
    layer0_outputs(335) <= b and not a;
    layer0_outputs(336) <= 1'b1;
    layer0_outputs(337) <= not b or a;
    layer0_outputs(338) <= a;
    layer0_outputs(339) <= a and not b;
    layer0_outputs(340) <= a and b;
    layer0_outputs(341) <= a xor b;
    layer0_outputs(342) <= a or b;
    layer0_outputs(343) <= a;
    layer0_outputs(344) <= a xor b;
    layer0_outputs(345) <= 1'b0;
    layer0_outputs(346) <= not (a or b);
    layer0_outputs(347) <= a xor b;
    layer0_outputs(348) <= a or b;
    layer0_outputs(349) <= a and not b;
    layer0_outputs(350) <= not (a or b);
    layer0_outputs(351) <= a or b;
    layer0_outputs(352) <= a or b;
    layer0_outputs(353) <= not b;
    layer0_outputs(354) <= b and not a;
    layer0_outputs(355) <= not b;
    layer0_outputs(356) <= 1'b1;
    layer0_outputs(357) <= not b or a;
    layer0_outputs(358) <= not a or b;
    layer0_outputs(359) <= not b or a;
    layer0_outputs(360) <= not (a or b);
    layer0_outputs(361) <= not (a or b);
    layer0_outputs(362) <= not b or a;
    layer0_outputs(363) <= not b;
    layer0_outputs(364) <= not (a xor b);
    layer0_outputs(365) <= not a or b;
    layer0_outputs(366) <= a;
    layer0_outputs(367) <= a or b;
    layer0_outputs(368) <= a xor b;
    layer0_outputs(369) <= not b;
    layer0_outputs(370) <= not a or b;
    layer0_outputs(371) <= not (a or b);
    layer0_outputs(372) <= a;
    layer0_outputs(373) <= not (a or b);
    layer0_outputs(374) <= a xor b;
    layer0_outputs(375) <= a and not b;
    layer0_outputs(376) <= not a;
    layer0_outputs(377) <= not b or a;
    layer0_outputs(378) <= a or b;
    layer0_outputs(379) <= a or b;
    layer0_outputs(380) <= not a;
    layer0_outputs(381) <= not (a or b);
    layer0_outputs(382) <= not a;
    layer0_outputs(383) <= not (a and b);
    layer0_outputs(384) <= a or b;
    layer0_outputs(385) <= 1'b1;
    layer0_outputs(386) <= a and not b;
    layer0_outputs(387) <= not a or b;
    layer0_outputs(388) <= a;
    layer0_outputs(389) <= a and not b;
    layer0_outputs(390) <= not (a and b);
    layer0_outputs(391) <= a xor b;
    layer0_outputs(392) <= a and not b;
    layer0_outputs(393) <= 1'b0;
    layer0_outputs(394) <= not (a and b);
    layer0_outputs(395) <= not a or b;
    layer0_outputs(396) <= a xor b;
    layer0_outputs(397) <= a;
    layer0_outputs(398) <= not (a xor b);
    layer0_outputs(399) <= a or b;
    layer0_outputs(400) <= b and not a;
    layer0_outputs(401) <= a and not b;
    layer0_outputs(402) <= 1'b1;
    layer0_outputs(403) <= not (a xor b);
    layer0_outputs(404) <= a xor b;
    layer0_outputs(405) <= not (a or b);
    layer0_outputs(406) <= a or b;
    layer0_outputs(407) <= not (a or b);
    layer0_outputs(408) <= not (a xor b);
    layer0_outputs(409) <= a;
    layer0_outputs(410) <= not b or a;
    layer0_outputs(411) <= a and not b;
    layer0_outputs(412) <= a or b;
    layer0_outputs(413) <= b;
    layer0_outputs(414) <= a and not b;
    layer0_outputs(415) <= a and not b;
    layer0_outputs(416) <= a or b;
    layer0_outputs(417) <= a or b;
    layer0_outputs(418) <= not b or a;
    layer0_outputs(419) <= not (a and b);
    layer0_outputs(420) <= a and b;
    layer0_outputs(421) <= b;
    layer0_outputs(422) <= not a;
    layer0_outputs(423) <= b;
    layer0_outputs(424) <= not b or a;
    layer0_outputs(425) <= a xor b;
    layer0_outputs(426) <= a or b;
    layer0_outputs(427) <= a;
    layer0_outputs(428) <= 1'b0;
    layer0_outputs(429) <= b;
    layer0_outputs(430) <= a and b;
    layer0_outputs(431) <= not (a and b);
    layer0_outputs(432) <= not b;
    layer0_outputs(433) <= not b;
    layer0_outputs(434) <= a and not b;
    layer0_outputs(435) <= a or b;
    layer0_outputs(436) <= not (a or b);
    layer0_outputs(437) <= not b or a;
    layer0_outputs(438) <= not b;
    layer0_outputs(439) <= a or b;
    layer0_outputs(440) <= a;
    layer0_outputs(441) <= not b or a;
    layer0_outputs(442) <= not b or a;
    layer0_outputs(443) <= a xor b;
    layer0_outputs(444) <= not a;
    layer0_outputs(445) <= b;
    layer0_outputs(446) <= a xor b;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= not (a or b);
    layer0_outputs(449) <= not (a or b);
    layer0_outputs(450) <= a;
    layer0_outputs(451) <= 1'b0;
    layer0_outputs(452) <= a xor b;
    layer0_outputs(453) <= not b or a;
    layer0_outputs(454) <= not (a and b);
    layer0_outputs(455) <= not (a xor b);
    layer0_outputs(456) <= not b;
    layer0_outputs(457) <= a;
    layer0_outputs(458) <= a xor b;
    layer0_outputs(459) <= 1'b0;
    layer0_outputs(460) <= a xor b;
    layer0_outputs(461) <= a or b;
    layer0_outputs(462) <= a xor b;
    layer0_outputs(463) <= a;
    layer0_outputs(464) <= not (a xor b);
    layer0_outputs(465) <= b and not a;
    layer0_outputs(466) <= not (a or b);
    layer0_outputs(467) <= a xor b;
    layer0_outputs(468) <= not b;
    layer0_outputs(469) <= not a;
    layer0_outputs(470) <= not (a or b);
    layer0_outputs(471) <= a xor b;
    layer0_outputs(472) <= a xor b;
    layer0_outputs(473) <= not (a or b);
    layer0_outputs(474) <= not b or a;
    layer0_outputs(475) <= a;
    layer0_outputs(476) <= b and not a;
    layer0_outputs(477) <= a and b;
    layer0_outputs(478) <= b;
    layer0_outputs(479) <= not (a or b);
    layer0_outputs(480) <= not a or b;
    layer0_outputs(481) <= not a or b;
    layer0_outputs(482) <= not (a xor b);
    layer0_outputs(483) <= not (a or b);
    layer0_outputs(484) <= a and b;
    layer0_outputs(485) <= a;
    layer0_outputs(486) <= a and not b;
    layer0_outputs(487) <= not (a or b);
    layer0_outputs(488) <= not a;
    layer0_outputs(489) <= not b;
    layer0_outputs(490) <= a or b;
    layer0_outputs(491) <= b and not a;
    layer0_outputs(492) <= a or b;
    layer0_outputs(493) <= not a;
    layer0_outputs(494) <= a;
    layer0_outputs(495) <= b and not a;
    layer0_outputs(496) <= not (a or b);
    layer0_outputs(497) <= a;
    layer0_outputs(498) <= not a;
    layer0_outputs(499) <= b;
    layer0_outputs(500) <= not b;
    layer0_outputs(501) <= a or b;
    layer0_outputs(502) <= a and not b;
    layer0_outputs(503) <= b and not a;
    layer0_outputs(504) <= b and not a;
    layer0_outputs(505) <= not (a and b);
    layer0_outputs(506) <= a or b;
    layer0_outputs(507) <= not a;
    layer0_outputs(508) <= not b or a;
    layer0_outputs(509) <= not a or b;
    layer0_outputs(510) <= not b;
    layer0_outputs(511) <= not a or b;
    layer0_outputs(512) <= not a or b;
    layer0_outputs(513) <= a or b;
    layer0_outputs(514) <= a and b;
    layer0_outputs(515) <= a or b;
    layer0_outputs(516) <= a and not b;
    layer0_outputs(517) <= b and not a;
    layer0_outputs(518) <= a and not b;
    layer0_outputs(519) <= a and b;
    layer0_outputs(520) <= b;
    layer0_outputs(521) <= b;
    layer0_outputs(522) <= not b or a;
    layer0_outputs(523) <= b and not a;
    layer0_outputs(524) <= not b or a;
    layer0_outputs(525) <= not b;
    layer0_outputs(526) <= not a;
    layer0_outputs(527) <= a and not b;
    layer0_outputs(528) <= a;
    layer0_outputs(529) <= not b;
    layer0_outputs(530) <= a and not b;
    layer0_outputs(531) <= b;
    layer0_outputs(532) <= not (a xor b);
    layer0_outputs(533) <= not (a xor b);
    layer0_outputs(534) <= a and not b;
    layer0_outputs(535) <= b and not a;
    layer0_outputs(536) <= not (a xor b);
    layer0_outputs(537) <= a and not b;
    layer0_outputs(538) <= a;
    layer0_outputs(539) <= 1'b0;
    layer0_outputs(540) <= 1'b1;
    layer0_outputs(541) <= a and b;
    layer0_outputs(542) <= b;
    layer0_outputs(543) <= not b;
    layer0_outputs(544) <= 1'b0;
    layer0_outputs(545) <= a;
    layer0_outputs(546) <= not b or a;
    layer0_outputs(547) <= not a;
    layer0_outputs(548) <= not b;
    layer0_outputs(549) <= not (a or b);
    layer0_outputs(550) <= not (a xor b);
    layer0_outputs(551) <= b and not a;
    layer0_outputs(552) <= not b or a;
    layer0_outputs(553) <= b;
    layer0_outputs(554) <= a or b;
    layer0_outputs(555) <= not (a or b);
    layer0_outputs(556) <= a and not b;
    layer0_outputs(557) <= b;
    layer0_outputs(558) <= not (a or b);
    layer0_outputs(559) <= a and not b;
    layer0_outputs(560) <= not (a or b);
    layer0_outputs(561) <= a;
    layer0_outputs(562) <= not b;
    layer0_outputs(563) <= a;
    layer0_outputs(564) <= a or b;
    layer0_outputs(565) <= a;
    layer0_outputs(566) <= 1'b1;
    layer0_outputs(567) <= not a or b;
    layer0_outputs(568) <= b and not a;
    layer0_outputs(569) <= a and not b;
    layer0_outputs(570) <= not (a and b);
    layer0_outputs(571) <= a or b;
    layer0_outputs(572) <= not b or a;
    layer0_outputs(573) <= a;
    layer0_outputs(574) <= a or b;
    layer0_outputs(575) <= a xor b;
    layer0_outputs(576) <= not (a or b);
    layer0_outputs(577) <= a and b;
    layer0_outputs(578) <= a xor b;
    layer0_outputs(579) <= not (a xor b);
    layer0_outputs(580) <= b and not a;
    layer0_outputs(581) <= a;
    layer0_outputs(582) <= not (a and b);
    layer0_outputs(583) <= a or b;
    layer0_outputs(584) <= a or b;
    layer0_outputs(585) <= not (a or b);
    layer0_outputs(586) <= 1'b0;
    layer0_outputs(587) <= a;
    layer0_outputs(588) <= not b or a;
    layer0_outputs(589) <= b and not a;
    layer0_outputs(590) <= 1'b1;
    layer0_outputs(591) <= a and not b;
    layer0_outputs(592) <= 1'b0;
    layer0_outputs(593) <= not a or b;
    layer0_outputs(594) <= a and b;
    layer0_outputs(595) <= b and not a;
    layer0_outputs(596) <= not a;
    layer0_outputs(597) <= a;
    layer0_outputs(598) <= not a;
    layer0_outputs(599) <= a or b;
    layer0_outputs(600) <= not (a or b);
    layer0_outputs(601) <= not (a or b);
    layer0_outputs(602) <= a or b;
    layer0_outputs(603) <= not (a xor b);
    layer0_outputs(604) <= a;
    layer0_outputs(605) <= a;
    layer0_outputs(606) <= 1'b0;
    layer0_outputs(607) <= a and b;
    layer0_outputs(608) <= b and not a;
    layer0_outputs(609) <= a xor b;
    layer0_outputs(610) <= a or b;
    layer0_outputs(611) <= b and not a;
    layer0_outputs(612) <= a or b;
    layer0_outputs(613) <= not a or b;
    layer0_outputs(614) <= 1'b0;
    layer0_outputs(615) <= not a or b;
    layer0_outputs(616) <= not (a or b);
    layer0_outputs(617) <= not b;
    layer0_outputs(618) <= not a;
    layer0_outputs(619) <= b;
    layer0_outputs(620) <= 1'b0;
    layer0_outputs(621) <= not (a or b);
    layer0_outputs(622) <= b and not a;
    layer0_outputs(623) <= not a or b;
    layer0_outputs(624) <= a and b;
    layer0_outputs(625) <= not b or a;
    layer0_outputs(626) <= b and not a;
    layer0_outputs(627) <= not (a xor b);
    layer0_outputs(628) <= a xor b;
    layer0_outputs(629) <= b and not a;
    layer0_outputs(630) <= not (a or b);
    layer0_outputs(631) <= 1'b1;
    layer0_outputs(632) <= a or b;
    layer0_outputs(633) <= a xor b;
    layer0_outputs(634) <= a and not b;
    layer0_outputs(635) <= 1'b1;
    layer0_outputs(636) <= not (a or b);
    layer0_outputs(637) <= not (a or b);
    layer0_outputs(638) <= a xor b;
    layer0_outputs(639) <= not b;
    layer0_outputs(640) <= not (a xor b);
    layer0_outputs(641) <= not (a xor b);
    layer0_outputs(642) <= a or b;
    layer0_outputs(643) <= a or b;
    layer0_outputs(644) <= not b or a;
    layer0_outputs(645) <= not b or a;
    layer0_outputs(646) <= a or b;
    layer0_outputs(647) <= a or b;
    layer0_outputs(648) <= b and not a;
    layer0_outputs(649) <= a or b;
    layer0_outputs(650) <= a or b;
    layer0_outputs(651) <= a;
    layer0_outputs(652) <= b;
    layer0_outputs(653) <= not (a or b);
    layer0_outputs(654) <= b;
    layer0_outputs(655) <= not (a or b);
    layer0_outputs(656) <= b;
    layer0_outputs(657) <= a or b;
    layer0_outputs(658) <= b;
    layer0_outputs(659) <= a and b;
    layer0_outputs(660) <= a and not b;
    layer0_outputs(661) <= not b or a;
    layer0_outputs(662) <= not (a or b);
    layer0_outputs(663) <= b;
    layer0_outputs(664) <= not b;
    layer0_outputs(665) <= not b;
    layer0_outputs(666) <= a and not b;
    layer0_outputs(667) <= not a or b;
    layer0_outputs(668) <= not (a or b);
    layer0_outputs(669) <= not b;
    layer0_outputs(670) <= a xor b;
    layer0_outputs(671) <= not a;
    layer0_outputs(672) <= a and not b;
    layer0_outputs(673) <= 1'b0;
    layer0_outputs(674) <= b;
    layer0_outputs(675) <= b;
    layer0_outputs(676) <= b;
    layer0_outputs(677) <= 1'b0;
    layer0_outputs(678) <= not a;
    layer0_outputs(679) <= 1'b0;
    layer0_outputs(680) <= not (a xor b);
    layer0_outputs(681) <= not b;
    layer0_outputs(682) <= b;
    layer0_outputs(683) <= a or b;
    layer0_outputs(684) <= b and not a;
    layer0_outputs(685) <= not b;
    layer0_outputs(686) <= not a;
    layer0_outputs(687) <= a or b;
    layer0_outputs(688) <= not (a xor b);
    layer0_outputs(689) <= a or b;
    layer0_outputs(690) <= not (a or b);
    layer0_outputs(691) <= a;
    layer0_outputs(692) <= not a or b;
    layer0_outputs(693) <= a;
    layer0_outputs(694) <= a or b;
    layer0_outputs(695) <= not (a xor b);
    layer0_outputs(696) <= not (a xor b);
    layer0_outputs(697) <= a or b;
    layer0_outputs(698) <= not a or b;
    layer0_outputs(699) <= b;
    layer0_outputs(700) <= not (a xor b);
    layer0_outputs(701) <= b;
    layer0_outputs(702) <= a and b;
    layer0_outputs(703) <= not (a or b);
    layer0_outputs(704) <= not b;
    layer0_outputs(705) <= not (a or b);
    layer0_outputs(706) <= a and not b;
    layer0_outputs(707) <= not (a xor b);
    layer0_outputs(708) <= not a or b;
    layer0_outputs(709) <= 1'b1;
    layer0_outputs(710) <= b;
    layer0_outputs(711) <= not (a xor b);
    layer0_outputs(712) <= not a;
    layer0_outputs(713) <= not a or b;
    layer0_outputs(714) <= 1'b1;
    layer0_outputs(715) <= not (a or b);
    layer0_outputs(716) <= not a or b;
    layer0_outputs(717) <= b;
    layer0_outputs(718) <= not (a or b);
    layer0_outputs(719) <= a or b;
    layer0_outputs(720) <= b;
    layer0_outputs(721) <= b and not a;
    layer0_outputs(722) <= not (a xor b);
    layer0_outputs(723) <= not b;
    layer0_outputs(724) <= 1'b1;
    layer0_outputs(725) <= not b;
    layer0_outputs(726) <= not b or a;
    layer0_outputs(727) <= not (a or b);
    layer0_outputs(728) <= not a;
    layer0_outputs(729) <= a or b;
    layer0_outputs(730) <= not (a or b);
    layer0_outputs(731) <= b;
    layer0_outputs(732) <= not (a or b);
    layer0_outputs(733) <= not (a or b);
    layer0_outputs(734) <= 1'b1;
    layer0_outputs(735) <= a xor b;
    layer0_outputs(736) <= not a;
    layer0_outputs(737) <= not a;
    layer0_outputs(738) <= b;
    layer0_outputs(739) <= not b or a;
    layer0_outputs(740) <= 1'b0;
    layer0_outputs(741) <= 1'b1;
    layer0_outputs(742) <= not b or a;
    layer0_outputs(743) <= b and not a;
    layer0_outputs(744) <= a;
    layer0_outputs(745) <= not a;
    layer0_outputs(746) <= not a or b;
    layer0_outputs(747) <= b and not a;
    layer0_outputs(748) <= not (a or b);
    layer0_outputs(749) <= not a or b;
    layer0_outputs(750) <= not (a xor b);
    layer0_outputs(751) <= not b or a;
    layer0_outputs(752) <= a;
    layer0_outputs(753) <= not b;
    layer0_outputs(754) <= a and b;
    layer0_outputs(755) <= a;
    layer0_outputs(756) <= b;
    layer0_outputs(757) <= b;
    layer0_outputs(758) <= a xor b;
    layer0_outputs(759) <= b and not a;
    layer0_outputs(760) <= a or b;
    layer0_outputs(761) <= not (a xor b);
    layer0_outputs(762) <= a or b;
    layer0_outputs(763) <= not a;
    layer0_outputs(764) <= a and not b;
    layer0_outputs(765) <= not b;
    layer0_outputs(766) <= not b;
    layer0_outputs(767) <= a or b;
    layer0_outputs(768) <= not a;
    layer0_outputs(769) <= a or b;
    layer0_outputs(770) <= not b;
    layer0_outputs(771) <= not (a or b);
    layer0_outputs(772) <= not (a and b);
    layer0_outputs(773) <= not b;
    layer0_outputs(774) <= 1'b1;
    layer0_outputs(775) <= a;
    layer0_outputs(776) <= not (a and b);
    layer0_outputs(777) <= not (a or b);
    layer0_outputs(778) <= b;
    layer0_outputs(779) <= a and not b;
    layer0_outputs(780) <= b;
    layer0_outputs(781) <= not (a xor b);
    layer0_outputs(782) <= a or b;
    layer0_outputs(783) <= not b;
    layer0_outputs(784) <= not (a or b);
    layer0_outputs(785) <= not a or b;
    layer0_outputs(786) <= b and not a;
    layer0_outputs(787) <= a and b;
    layer0_outputs(788) <= not (a or b);
    layer0_outputs(789) <= 1'b0;
    layer0_outputs(790) <= a;
    layer0_outputs(791) <= b;
    layer0_outputs(792) <= not (a xor b);
    layer0_outputs(793) <= a;
    layer0_outputs(794) <= not (a and b);
    layer0_outputs(795) <= not (a or b);
    layer0_outputs(796) <= 1'b0;
    layer0_outputs(797) <= a and not b;
    layer0_outputs(798) <= b and not a;
    layer0_outputs(799) <= not (a or b);
    layer0_outputs(800) <= not (a or b);
    layer0_outputs(801) <= not (a or b);
    layer0_outputs(802) <= b and not a;
    layer0_outputs(803) <= a or b;
    layer0_outputs(804) <= a and not b;
    layer0_outputs(805) <= a and b;
    layer0_outputs(806) <= a and not b;
    layer0_outputs(807) <= not (a or b);
    layer0_outputs(808) <= not (a or b);
    layer0_outputs(809) <= b and not a;
    layer0_outputs(810) <= not a;
    layer0_outputs(811) <= not (a or b);
    layer0_outputs(812) <= b;
    layer0_outputs(813) <= not b;
    layer0_outputs(814) <= not b;
    layer0_outputs(815) <= not (a or b);
    layer0_outputs(816) <= a;
    layer0_outputs(817) <= a and b;
    layer0_outputs(818) <= 1'b0;
    layer0_outputs(819) <= not b or a;
    layer0_outputs(820) <= not (a or b);
    layer0_outputs(821) <= 1'b1;
    layer0_outputs(822) <= 1'b0;
    layer0_outputs(823) <= a xor b;
    layer0_outputs(824) <= not (a or b);
    layer0_outputs(825) <= b;
    layer0_outputs(826) <= b and not a;
    layer0_outputs(827) <= a and not b;
    layer0_outputs(828) <= not b or a;
    layer0_outputs(829) <= not (a or b);
    layer0_outputs(830) <= not a or b;
    layer0_outputs(831) <= a xor b;
    layer0_outputs(832) <= a and not b;
    layer0_outputs(833) <= b;
    layer0_outputs(834) <= b;
    layer0_outputs(835) <= a;
    layer0_outputs(836) <= a or b;
    layer0_outputs(837) <= a;
    layer0_outputs(838) <= b;
    layer0_outputs(839) <= not a or b;
    layer0_outputs(840) <= a or b;
    layer0_outputs(841) <= not (a and b);
    layer0_outputs(842) <= not a;
    layer0_outputs(843) <= not b or a;
    layer0_outputs(844) <= not (a or b);
    layer0_outputs(845) <= not b;
    layer0_outputs(846) <= not b or a;
    layer0_outputs(847) <= a and not b;
    layer0_outputs(848) <= 1'b1;
    layer0_outputs(849) <= not (a or b);
    layer0_outputs(850) <= b;
    layer0_outputs(851) <= not (a or b);
    layer0_outputs(852) <= a or b;
    layer0_outputs(853) <= not a or b;
    layer0_outputs(854) <= a;
    layer0_outputs(855) <= a or b;
    layer0_outputs(856) <= not b or a;
    layer0_outputs(857) <= not (a or b);
    layer0_outputs(858) <= a and not b;
    layer0_outputs(859) <= not (a or b);
    layer0_outputs(860) <= a or b;
    layer0_outputs(861) <= not (a or b);
    layer0_outputs(862) <= a and b;
    layer0_outputs(863) <= a and not b;
    layer0_outputs(864) <= b;
    layer0_outputs(865) <= not (a or b);
    layer0_outputs(866) <= not (a and b);
    layer0_outputs(867) <= not b;
    layer0_outputs(868) <= a and not b;
    layer0_outputs(869) <= not b or a;
    layer0_outputs(870) <= a;
    layer0_outputs(871) <= not (a xor b);
    layer0_outputs(872) <= not a or b;
    layer0_outputs(873) <= a and not b;
    layer0_outputs(874) <= not a or b;
    layer0_outputs(875) <= not (a and b);
    layer0_outputs(876) <= a or b;
    layer0_outputs(877) <= 1'b1;
    layer0_outputs(878) <= b;
    layer0_outputs(879) <= not a;
    layer0_outputs(880) <= a or b;
    layer0_outputs(881) <= not (a or b);
    layer0_outputs(882) <= a and not b;
    layer0_outputs(883) <= a and not b;
    layer0_outputs(884) <= a;
    layer0_outputs(885) <= a or b;
    layer0_outputs(886) <= 1'b0;
    layer0_outputs(887) <= a;
    layer0_outputs(888) <= not b;
    layer0_outputs(889) <= 1'b1;
    layer0_outputs(890) <= not a;
    layer0_outputs(891) <= a and b;
    layer0_outputs(892) <= b and not a;
    layer0_outputs(893) <= not (a or b);
    layer0_outputs(894) <= not (a xor b);
    layer0_outputs(895) <= not (a and b);
    layer0_outputs(896) <= a;
    layer0_outputs(897) <= a;
    layer0_outputs(898) <= not b;
    layer0_outputs(899) <= not (a or b);
    layer0_outputs(900) <= not (a and b);
    layer0_outputs(901) <= not b;
    layer0_outputs(902) <= not (a or b);
    layer0_outputs(903) <= not b;
    layer0_outputs(904) <= b;
    layer0_outputs(905) <= not (a and b);
    layer0_outputs(906) <= a xor b;
    layer0_outputs(907) <= not (a xor b);
    layer0_outputs(908) <= not a;
    layer0_outputs(909) <= a or b;
    layer0_outputs(910) <= a or b;
    layer0_outputs(911) <= not a or b;
    layer0_outputs(912) <= not (a or b);
    layer0_outputs(913) <= b;
    layer0_outputs(914) <= not b;
    layer0_outputs(915) <= not (a or b);
    layer0_outputs(916) <= not (a or b);
    layer0_outputs(917) <= a and b;
    layer0_outputs(918) <= a;
    layer0_outputs(919) <= a;
    layer0_outputs(920) <= not b or a;
    layer0_outputs(921) <= not b or a;
    layer0_outputs(922) <= not b;
    layer0_outputs(923) <= b and not a;
    layer0_outputs(924) <= b;
    layer0_outputs(925) <= not b or a;
    layer0_outputs(926) <= b;
    layer0_outputs(927) <= not (a and b);
    layer0_outputs(928) <= a;
    layer0_outputs(929) <= not (a or b);
    layer0_outputs(930) <= not a;
    layer0_outputs(931) <= not (a xor b);
    layer0_outputs(932) <= a;
    layer0_outputs(933) <= a and not b;
    layer0_outputs(934) <= not b or a;
    layer0_outputs(935) <= a or b;
    layer0_outputs(936) <= a;
    layer0_outputs(937) <= b;
    layer0_outputs(938) <= not (a or b);
    layer0_outputs(939) <= a xor b;
    layer0_outputs(940) <= not a;
    layer0_outputs(941) <= a and b;
    layer0_outputs(942) <= 1'b1;
    layer0_outputs(943) <= not a;
    layer0_outputs(944) <= not b or a;
    layer0_outputs(945) <= b;
    layer0_outputs(946) <= b and not a;
    layer0_outputs(947) <= not (a or b);
    layer0_outputs(948) <= b and not a;
    layer0_outputs(949) <= not (a or b);
    layer0_outputs(950) <= not (a and b);
    layer0_outputs(951) <= not b or a;
    layer0_outputs(952) <= a or b;
    layer0_outputs(953) <= a and b;
    layer0_outputs(954) <= a;
    layer0_outputs(955) <= not (a or b);
    layer0_outputs(956) <= not (a or b);
    layer0_outputs(957) <= not a or b;
    layer0_outputs(958) <= not (a or b);
    layer0_outputs(959) <= a or b;
    layer0_outputs(960) <= not (a and b);
    layer0_outputs(961) <= b and not a;
    layer0_outputs(962) <= not b;
    layer0_outputs(963) <= b;
    layer0_outputs(964) <= a;
    layer0_outputs(965) <= not (a and b);
    layer0_outputs(966) <= a and b;
    layer0_outputs(967) <= not (a or b);
    layer0_outputs(968) <= not (a or b);
    layer0_outputs(969) <= not (a and b);
    layer0_outputs(970) <= a or b;
    layer0_outputs(971) <= 1'b0;
    layer0_outputs(972) <= not b;
    layer0_outputs(973) <= a xor b;
    layer0_outputs(974) <= not b;
    layer0_outputs(975) <= a or b;
    layer0_outputs(976) <= a xor b;
    layer0_outputs(977) <= not (a or b);
    layer0_outputs(978) <= not (a and b);
    layer0_outputs(979) <= not (a xor b);
    layer0_outputs(980) <= not a;
    layer0_outputs(981) <= b;
    layer0_outputs(982) <= not a;
    layer0_outputs(983) <= 1'b0;
    layer0_outputs(984) <= a and not b;
    layer0_outputs(985) <= a or b;
    layer0_outputs(986) <= not b;
    layer0_outputs(987) <= not (a xor b);
    layer0_outputs(988) <= a or b;
    layer0_outputs(989) <= b;
    layer0_outputs(990) <= not b or a;
    layer0_outputs(991) <= b and not a;
    layer0_outputs(992) <= a;
    layer0_outputs(993) <= not a or b;
    layer0_outputs(994) <= not (a xor b);
    layer0_outputs(995) <= not (a xor b);
    layer0_outputs(996) <= b;
    layer0_outputs(997) <= not b;
    layer0_outputs(998) <= not b or a;
    layer0_outputs(999) <= a and b;
    layer0_outputs(1000) <= not a;
    layer0_outputs(1001) <= a;
    layer0_outputs(1002) <= a;
    layer0_outputs(1003) <= not b or a;
    layer0_outputs(1004) <= b and not a;
    layer0_outputs(1005) <= not (a xor b);
    layer0_outputs(1006) <= not (a or b);
    layer0_outputs(1007) <= not (a xor b);
    layer0_outputs(1008) <= not a;
    layer0_outputs(1009) <= not (a xor b);
    layer0_outputs(1010) <= not (a or b);
    layer0_outputs(1011) <= b;
    layer0_outputs(1012) <= not (a xor b);
    layer0_outputs(1013) <= b and not a;
    layer0_outputs(1014) <= a;
    layer0_outputs(1015) <= not b;
    layer0_outputs(1016) <= not (a xor b);
    layer0_outputs(1017) <= not b or a;
    layer0_outputs(1018) <= not a or b;
    layer0_outputs(1019) <= b;
    layer0_outputs(1020) <= b;
    layer0_outputs(1021) <= not (a xor b);
    layer0_outputs(1022) <= not (a or b);
    layer0_outputs(1023) <= not (a or b);
    layer0_outputs(1024) <= a and not b;
    layer0_outputs(1025) <= not a;
    layer0_outputs(1026) <= a or b;
    layer0_outputs(1027) <= b;
    layer0_outputs(1028) <= not a;
    layer0_outputs(1029) <= 1'b1;
    layer0_outputs(1030) <= not (a and b);
    layer0_outputs(1031) <= not a;
    layer0_outputs(1032) <= not a;
    layer0_outputs(1033) <= b and not a;
    layer0_outputs(1034) <= not a;
    layer0_outputs(1035) <= not b;
    layer0_outputs(1036) <= not b;
    layer0_outputs(1037) <= b and not a;
    layer0_outputs(1038) <= b and not a;
    layer0_outputs(1039) <= a or b;
    layer0_outputs(1040) <= not a;
    layer0_outputs(1041) <= not (a and b);
    layer0_outputs(1042) <= not (a xor b);
    layer0_outputs(1043) <= b and not a;
    layer0_outputs(1044) <= a;
    layer0_outputs(1045) <= not (a or b);
    layer0_outputs(1046) <= b;
    layer0_outputs(1047) <= 1'b1;
    layer0_outputs(1048) <= not b;
    layer0_outputs(1049) <= not a or b;
    layer0_outputs(1050) <= a or b;
    layer0_outputs(1051) <= not a;
    layer0_outputs(1052) <= not (a and b);
    layer0_outputs(1053) <= not a or b;
    layer0_outputs(1054) <= b;
    layer0_outputs(1055) <= a or b;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= b;
    layer0_outputs(1058) <= a or b;
    layer0_outputs(1059) <= a xor b;
    layer0_outputs(1060) <= not a;
    layer0_outputs(1061) <= not a;
    layer0_outputs(1062) <= a and b;
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= a;
    layer0_outputs(1065) <= not b or a;
    layer0_outputs(1066) <= not (a or b);
    layer0_outputs(1067) <= a;
    layer0_outputs(1068) <= a xor b;
    layer0_outputs(1069) <= not (a or b);
    layer0_outputs(1070) <= b and not a;
    layer0_outputs(1071) <= not b;
    layer0_outputs(1072) <= b;
    layer0_outputs(1073) <= not b;
    layer0_outputs(1074) <= b;
    layer0_outputs(1075) <= a or b;
    layer0_outputs(1076) <= 1'b0;
    layer0_outputs(1077) <= not b or a;
    layer0_outputs(1078) <= b;
    layer0_outputs(1079) <= a;
    layer0_outputs(1080) <= 1'b1;
    layer0_outputs(1081) <= not (a and b);
    layer0_outputs(1082) <= not b;
    layer0_outputs(1083) <= a xor b;
    layer0_outputs(1084) <= a or b;
    layer0_outputs(1085) <= not a or b;
    layer0_outputs(1086) <= not (a xor b);
    layer0_outputs(1087) <= not a;
    layer0_outputs(1088) <= not a;
    layer0_outputs(1089) <= not a or b;
    layer0_outputs(1090) <= not b;
    layer0_outputs(1091) <= not (a or b);
    layer0_outputs(1092) <= b;
    layer0_outputs(1093) <= a;
    layer0_outputs(1094) <= not (a xor b);
    layer0_outputs(1095) <= a and not b;
    layer0_outputs(1096) <= a;
    layer0_outputs(1097) <= not b or a;
    layer0_outputs(1098) <= not b or a;
    layer0_outputs(1099) <= a and b;
    layer0_outputs(1100) <= a;
    layer0_outputs(1101) <= not a or b;
    layer0_outputs(1102) <= not a or b;
    layer0_outputs(1103) <= a and not b;
    layer0_outputs(1104) <= a;
    layer0_outputs(1105) <= b and not a;
    layer0_outputs(1106) <= a xor b;
    layer0_outputs(1107) <= a and not b;
    layer0_outputs(1108) <= b;
    layer0_outputs(1109) <= not a;
    layer0_outputs(1110) <= a or b;
    layer0_outputs(1111) <= not b;
    layer0_outputs(1112) <= a;
    layer0_outputs(1113) <= a and not b;
    layer0_outputs(1114) <= not a or b;
    layer0_outputs(1115) <= a;
    layer0_outputs(1116) <= a;
    layer0_outputs(1117) <= not (a or b);
    layer0_outputs(1118) <= b;
    layer0_outputs(1119) <= not a or b;
    layer0_outputs(1120) <= b and not a;
    layer0_outputs(1121) <= b;
    layer0_outputs(1122) <= b;
    layer0_outputs(1123) <= not b;
    layer0_outputs(1124) <= a xor b;
    layer0_outputs(1125) <= b;
    layer0_outputs(1126) <= not (a or b);
    layer0_outputs(1127) <= a;
    layer0_outputs(1128) <= a or b;
    layer0_outputs(1129) <= not (a or b);
    layer0_outputs(1130) <= 1'b1;
    layer0_outputs(1131) <= not (a xor b);
    layer0_outputs(1132) <= a;
    layer0_outputs(1133) <= b;
    layer0_outputs(1134) <= b and not a;
    layer0_outputs(1135) <= b;
    layer0_outputs(1136) <= not (a or b);
    layer0_outputs(1137) <= a xor b;
    layer0_outputs(1138) <= a;
    layer0_outputs(1139) <= a and not b;
    layer0_outputs(1140) <= b;
    layer0_outputs(1141) <= b;
    layer0_outputs(1142) <= not b;
    layer0_outputs(1143) <= b and not a;
    layer0_outputs(1144) <= b and not a;
    layer0_outputs(1145) <= not a or b;
    layer0_outputs(1146) <= not (a or b);
    layer0_outputs(1147) <= not b;
    layer0_outputs(1148) <= a xor b;
    layer0_outputs(1149) <= a;
    layer0_outputs(1150) <= not b or a;
    layer0_outputs(1151) <= not (a or b);
    layer0_outputs(1152) <= a xor b;
    layer0_outputs(1153) <= not (a or b);
    layer0_outputs(1154) <= not (a and b);
    layer0_outputs(1155) <= b and not a;
    layer0_outputs(1156) <= b;
    layer0_outputs(1157) <= b and not a;
    layer0_outputs(1158) <= a and b;
    layer0_outputs(1159) <= not b or a;
    layer0_outputs(1160) <= a;
    layer0_outputs(1161) <= a xor b;
    layer0_outputs(1162) <= a and not b;
    layer0_outputs(1163) <= not a or b;
    layer0_outputs(1164) <= not b;
    layer0_outputs(1165) <= a and not b;
    layer0_outputs(1166) <= a and not b;
    layer0_outputs(1167) <= not (a xor b);
    layer0_outputs(1168) <= a xor b;
    layer0_outputs(1169) <= a and b;
    layer0_outputs(1170) <= b and not a;
    layer0_outputs(1171) <= a and not b;
    layer0_outputs(1172) <= not b;
    layer0_outputs(1173) <= a or b;
    layer0_outputs(1174) <= a;
    layer0_outputs(1175) <= not a or b;
    layer0_outputs(1176) <= not a or b;
    layer0_outputs(1177) <= not a or b;
    layer0_outputs(1178) <= not a or b;
    layer0_outputs(1179) <= 1'b0;
    layer0_outputs(1180) <= not a or b;
    layer0_outputs(1181) <= a and b;
    layer0_outputs(1182) <= a or b;
    layer0_outputs(1183) <= a xor b;
    layer0_outputs(1184) <= a xor b;
    layer0_outputs(1185) <= a;
    layer0_outputs(1186) <= not b or a;
    layer0_outputs(1187) <= 1'b0;
    layer0_outputs(1188) <= b;
    layer0_outputs(1189) <= a xor b;
    layer0_outputs(1190) <= a or b;
    layer0_outputs(1191) <= not b;
    layer0_outputs(1192) <= a or b;
    layer0_outputs(1193) <= 1'b1;
    layer0_outputs(1194) <= a and not b;
    layer0_outputs(1195) <= not (a and b);
    layer0_outputs(1196) <= b and not a;
    layer0_outputs(1197) <= not (a or b);
    layer0_outputs(1198) <= not (a or b);
    layer0_outputs(1199) <= not (a xor b);
    layer0_outputs(1200) <= not b;
    layer0_outputs(1201) <= a xor b;
    layer0_outputs(1202) <= b;
    layer0_outputs(1203) <= a;
    layer0_outputs(1204) <= not a;
    layer0_outputs(1205) <= 1'b0;
    layer0_outputs(1206) <= a or b;
    layer0_outputs(1207) <= not a;
    layer0_outputs(1208) <= not (a or b);
    layer0_outputs(1209) <= 1'b0;
    layer0_outputs(1210) <= not b or a;
    layer0_outputs(1211) <= not a or b;
    layer0_outputs(1212) <= a or b;
    layer0_outputs(1213) <= 1'b0;
    layer0_outputs(1214) <= not a;
    layer0_outputs(1215) <= not a or b;
    layer0_outputs(1216) <= b;
    layer0_outputs(1217) <= a;
    layer0_outputs(1218) <= a or b;
    layer0_outputs(1219) <= a or b;
    layer0_outputs(1220) <= a or b;
    layer0_outputs(1221) <= a;
    layer0_outputs(1222) <= not (a or b);
    layer0_outputs(1223) <= not a;
    layer0_outputs(1224) <= a;
    layer0_outputs(1225) <= a or b;
    layer0_outputs(1226) <= a or b;
    layer0_outputs(1227) <= a;
    layer0_outputs(1228) <= a and not b;
    layer0_outputs(1229) <= a;
    layer0_outputs(1230) <= not (a and b);
    layer0_outputs(1231) <= a;
    layer0_outputs(1232) <= a and not b;
    layer0_outputs(1233) <= not a or b;
    layer0_outputs(1234) <= a xor b;
    layer0_outputs(1235) <= a or b;
    layer0_outputs(1236) <= not b;
    layer0_outputs(1237) <= b;
    layer0_outputs(1238) <= 1'b0;
    layer0_outputs(1239) <= a or b;
    layer0_outputs(1240) <= a or b;
    layer0_outputs(1241) <= a xor b;
    layer0_outputs(1242) <= not (a or b);
    layer0_outputs(1243) <= a xor b;
    layer0_outputs(1244) <= not a or b;
    layer0_outputs(1245) <= not b;
    layer0_outputs(1246) <= not (a or b);
    layer0_outputs(1247) <= not (a or b);
    layer0_outputs(1248) <= not (a or b);
    layer0_outputs(1249) <= 1'b1;
    layer0_outputs(1250) <= b and not a;
    layer0_outputs(1251) <= 1'b0;
    layer0_outputs(1252) <= not a;
    layer0_outputs(1253) <= 1'b0;
    layer0_outputs(1254) <= a xor b;
    layer0_outputs(1255) <= 1'b1;
    layer0_outputs(1256) <= 1'b1;
    layer0_outputs(1257) <= not b or a;
    layer0_outputs(1258) <= a;
    layer0_outputs(1259) <= not (a or b);
    layer0_outputs(1260) <= a xor b;
    layer0_outputs(1261) <= not b;
    layer0_outputs(1262) <= a xor b;
    layer0_outputs(1263) <= not b or a;
    layer0_outputs(1264) <= a;
    layer0_outputs(1265) <= a;
    layer0_outputs(1266) <= b;
    layer0_outputs(1267) <= not b or a;
    layer0_outputs(1268) <= a xor b;
    layer0_outputs(1269) <= b and not a;
    layer0_outputs(1270) <= not (a xor b);
    layer0_outputs(1271) <= not (a or b);
    layer0_outputs(1272) <= not (a or b);
    layer0_outputs(1273) <= not (a xor b);
    layer0_outputs(1274) <= b;
    layer0_outputs(1275) <= not (a and b);
    layer0_outputs(1276) <= not b or a;
    layer0_outputs(1277) <= a or b;
    layer0_outputs(1278) <= 1'b0;
    layer0_outputs(1279) <= not a or b;
    layer0_outputs(1280) <= a xor b;
    layer0_outputs(1281) <= a or b;
    layer0_outputs(1282) <= not (a or b);
    layer0_outputs(1283) <= not a or b;
    layer0_outputs(1284) <= a or b;
    layer0_outputs(1285) <= b and not a;
    layer0_outputs(1286) <= not (a or b);
    layer0_outputs(1287) <= a;
    layer0_outputs(1288) <= not (a or b);
    layer0_outputs(1289) <= not a;
    layer0_outputs(1290) <= not a;
    layer0_outputs(1291) <= a xor b;
    layer0_outputs(1292) <= 1'b0;
    layer0_outputs(1293) <= not (a or b);
    layer0_outputs(1294) <= not (a xor b);
    layer0_outputs(1295) <= not b;
    layer0_outputs(1296) <= a and not b;
    layer0_outputs(1297) <= not a;
    layer0_outputs(1298) <= 1'b0;
    layer0_outputs(1299) <= 1'b1;
    layer0_outputs(1300) <= not b;
    layer0_outputs(1301) <= a or b;
    layer0_outputs(1302) <= not (a xor b);
    layer0_outputs(1303) <= not a;
    layer0_outputs(1304) <= b;
    layer0_outputs(1305) <= not b;
    layer0_outputs(1306) <= b;
    layer0_outputs(1307) <= 1'b0;
    layer0_outputs(1308) <= not a;
    layer0_outputs(1309) <= a and b;
    layer0_outputs(1310) <= not (a or b);
    layer0_outputs(1311) <= not a or b;
    layer0_outputs(1312) <= a and not b;
    layer0_outputs(1313) <= not b;
    layer0_outputs(1314) <= not a or b;
    layer0_outputs(1315) <= 1'b1;
    layer0_outputs(1316) <= not (a and b);
    layer0_outputs(1317) <= not a or b;
    layer0_outputs(1318) <= a and not b;
    layer0_outputs(1319) <= a or b;
    layer0_outputs(1320) <= a or b;
    layer0_outputs(1321) <= 1'b0;
    layer0_outputs(1322) <= a xor b;
    layer0_outputs(1323) <= b;
    layer0_outputs(1324) <= 1'b1;
    layer0_outputs(1325) <= a or b;
    layer0_outputs(1326) <= not a or b;
    layer0_outputs(1327) <= a xor b;
    layer0_outputs(1328) <= b and not a;
    layer0_outputs(1329) <= a or b;
    layer0_outputs(1330) <= not a or b;
    layer0_outputs(1331) <= b and not a;
    layer0_outputs(1332) <= not a or b;
    layer0_outputs(1333) <= 1'b0;
    layer0_outputs(1334) <= a;
    layer0_outputs(1335) <= a and not b;
    layer0_outputs(1336) <= a;
    layer0_outputs(1337) <= a or b;
    layer0_outputs(1338) <= a xor b;
    layer0_outputs(1339) <= a or b;
    layer0_outputs(1340) <= 1'b1;
    layer0_outputs(1341) <= a xor b;
    layer0_outputs(1342) <= a xor b;
    layer0_outputs(1343) <= not b or a;
    layer0_outputs(1344) <= not (a xor b);
    layer0_outputs(1345) <= 1'b0;
    layer0_outputs(1346) <= not (a or b);
    layer0_outputs(1347) <= 1'b0;
    layer0_outputs(1348) <= not a or b;
    layer0_outputs(1349) <= not b;
    layer0_outputs(1350) <= a;
    layer0_outputs(1351) <= not b;
    layer0_outputs(1352) <= b and not a;
    layer0_outputs(1353) <= not (a xor b);
    layer0_outputs(1354) <= not b or a;
    layer0_outputs(1355) <= not a;
    layer0_outputs(1356) <= b and not a;
    layer0_outputs(1357) <= not a;
    layer0_outputs(1358) <= b;
    layer0_outputs(1359) <= b;
    layer0_outputs(1360) <= a;
    layer0_outputs(1361) <= not (a or b);
    layer0_outputs(1362) <= 1'b1;
    layer0_outputs(1363) <= a;
    layer0_outputs(1364) <= b and not a;
    layer0_outputs(1365) <= a or b;
    layer0_outputs(1366) <= a;
    layer0_outputs(1367) <= not b or a;
    layer0_outputs(1368) <= 1'b1;
    layer0_outputs(1369) <= a or b;
    layer0_outputs(1370) <= not (a or b);
    layer0_outputs(1371) <= not (a and b);
    layer0_outputs(1372) <= a or b;
    layer0_outputs(1373) <= 1'b0;
    layer0_outputs(1374) <= not b or a;
    layer0_outputs(1375) <= a and not b;
    layer0_outputs(1376) <= not a;
    layer0_outputs(1377) <= not (a or b);
    layer0_outputs(1378) <= not b;
    layer0_outputs(1379) <= a or b;
    layer0_outputs(1380) <= a or b;
    layer0_outputs(1381) <= a or b;
    layer0_outputs(1382) <= a xor b;
    layer0_outputs(1383) <= a and not b;
    layer0_outputs(1384) <= not (a or b);
    layer0_outputs(1385) <= 1'b1;
    layer0_outputs(1386) <= not (a xor b);
    layer0_outputs(1387) <= a xor b;
    layer0_outputs(1388) <= not (a or b);
    layer0_outputs(1389) <= a xor b;
    layer0_outputs(1390) <= not a;
    layer0_outputs(1391) <= not (a or b);
    layer0_outputs(1392) <= not (a or b);
    layer0_outputs(1393) <= a or b;
    layer0_outputs(1394) <= not (a or b);
    layer0_outputs(1395) <= not (a and b);
    layer0_outputs(1396) <= not (a xor b);
    layer0_outputs(1397) <= 1'b1;
    layer0_outputs(1398) <= b;
    layer0_outputs(1399) <= b;
    layer0_outputs(1400) <= not b or a;
    layer0_outputs(1401) <= not (a or b);
    layer0_outputs(1402) <= 1'b0;
    layer0_outputs(1403) <= b;
    layer0_outputs(1404) <= a xor b;
    layer0_outputs(1405) <= a;
    layer0_outputs(1406) <= a or b;
    layer0_outputs(1407) <= not b;
    layer0_outputs(1408) <= 1'b1;
    layer0_outputs(1409) <= not a or b;
    layer0_outputs(1410) <= a and not b;
    layer0_outputs(1411) <= a xor b;
    layer0_outputs(1412) <= not a;
    layer0_outputs(1413) <= b and not a;
    layer0_outputs(1414) <= a and not b;
    layer0_outputs(1415) <= not a or b;
    layer0_outputs(1416) <= a or b;
    layer0_outputs(1417) <= b and not a;
    layer0_outputs(1418) <= a and not b;
    layer0_outputs(1419) <= not b or a;
    layer0_outputs(1420) <= a and not b;
    layer0_outputs(1421) <= not (a and b);
    layer0_outputs(1422) <= not (a or b);
    layer0_outputs(1423) <= not a or b;
    layer0_outputs(1424) <= a;
    layer0_outputs(1425) <= a;
    layer0_outputs(1426) <= 1'b0;
    layer0_outputs(1427) <= not (a and b);
    layer0_outputs(1428) <= 1'b0;
    layer0_outputs(1429) <= not a or b;
    layer0_outputs(1430) <= not a;
    layer0_outputs(1431) <= b;
    layer0_outputs(1432) <= not (a and b);
    layer0_outputs(1433) <= not b or a;
    layer0_outputs(1434) <= a or b;
    layer0_outputs(1435) <= a and not b;
    layer0_outputs(1436) <= not (a or b);
    layer0_outputs(1437) <= not b or a;
    layer0_outputs(1438) <= b and not a;
    layer0_outputs(1439) <= b and not a;
    layer0_outputs(1440) <= b;
    layer0_outputs(1441) <= a and b;
    layer0_outputs(1442) <= not b;
    layer0_outputs(1443) <= not (a or b);
    layer0_outputs(1444) <= a;
    layer0_outputs(1445) <= a;
    layer0_outputs(1446) <= 1'b1;
    layer0_outputs(1447) <= a and not b;
    layer0_outputs(1448) <= b;
    layer0_outputs(1449) <= 1'b0;
    layer0_outputs(1450) <= a and not b;
    layer0_outputs(1451) <= b and not a;
    layer0_outputs(1452) <= not b;
    layer0_outputs(1453) <= b and not a;
    layer0_outputs(1454) <= not (a and b);
    layer0_outputs(1455) <= a and not b;
    layer0_outputs(1456) <= not b or a;
    layer0_outputs(1457) <= not (a or b);
    layer0_outputs(1458) <= not b or a;
    layer0_outputs(1459) <= not (a or b);
    layer0_outputs(1460) <= a or b;
    layer0_outputs(1461) <= a and not b;
    layer0_outputs(1462) <= not (a or b);
    layer0_outputs(1463) <= b;
    layer0_outputs(1464) <= b;
    layer0_outputs(1465) <= not b;
    layer0_outputs(1466) <= not a;
    layer0_outputs(1467) <= not (a xor b);
    layer0_outputs(1468) <= not b;
    layer0_outputs(1469) <= 1'b1;
    layer0_outputs(1470) <= not (a xor b);
    layer0_outputs(1471) <= b and not a;
    layer0_outputs(1472) <= b;
    layer0_outputs(1473) <= a;
    layer0_outputs(1474) <= 1'b1;
    layer0_outputs(1475) <= not (a or b);
    layer0_outputs(1476) <= b and not a;
    layer0_outputs(1477) <= b;
    layer0_outputs(1478) <= a or b;
    layer0_outputs(1479) <= not (a xor b);
    layer0_outputs(1480) <= not (a and b);
    layer0_outputs(1481) <= not b;
    layer0_outputs(1482) <= a;
    layer0_outputs(1483) <= not (a or b);
    layer0_outputs(1484) <= a and not b;
    layer0_outputs(1485) <= b and not a;
    layer0_outputs(1486) <= a xor b;
    layer0_outputs(1487) <= not a;
    layer0_outputs(1488) <= 1'b1;
    layer0_outputs(1489) <= b and not a;
    layer0_outputs(1490) <= a and not b;
    layer0_outputs(1491) <= b;
    layer0_outputs(1492) <= not b;
    layer0_outputs(1493) <= a;
    layer0_outputs(1494) <= not b;
    layer0_outputs(1495) <= not a;
    layer0_outputs(1496) <= a;
    layer0_outputs(1497) <= not a or b;
    layer0_outputs(1498) <= not b or a;
    layer0_outputs(1499) <= a and not b;
    layer0_outputs(1500) <= not (a xor b);
    layer0_outputs(1501) <= not (a and b);
    layer0_outputs(1502) <= a xor b;
    layer0_outputs(1503) <= a;
    layer0_outputs(1504) <= not a;
    layer0_outputs(1505) <= a or b;
    layer0_outputs(1506) <= not b;
    layer0_outputs(1507) <= b;
    layer0_outputs(1508) <= not a or b;
    layer0_outputs(1509) <= not (a or b);
    layer0_outputs(1510) <= not (a or b);
    layer0_outputs(1511) <= b;
    layer0_outputs(1512) <= not a or b;
    layer0_outputs(1513) <= b and not a;
    layer0_outputs(1514) <= a or b;
    layer0_outputs(1515) <= not (a or b);
    layer0_outputs(1516) <= a or b;
    layer0_outputs(1517) <= 1'b1;
    layer0_outputs(1518) <= a xor b;
    layer0_outputs(1519) <= a or b;
    layer0_outputs(1520) <= a or b;
    layer0_outputs(1521) <= not b or a;
    layer0_outputs(1522) <= a xor b;
    layer0_outputs(1523) <= not b;
    layer0_outputs(1524) <= a or b;
    layer0_outputs(1525) <= not (a or b);
    layer0_outputs(1526) <= a;
    layer0_outputs(1527) <= a or b;
    layer0_outputs(1528) <= not (a or b);
    layer0_outputs(1529) <= not a or b;
    layer0_outputs(1530) <= not (a xor b);
    layer0_outputs(1531) <= b;
    layer0_outputs(1532) <= not (a xor b);
    layer0_outputs(1533) <= a or b;
    layer0_outputs(1534) <= not b or a;
    layer0_outputs(1535) <= a or b;
    layer0_outputs(1536) <= b and not a;
    layer0_outputs(1537) <= a xor b;
    layer0_outputs(1538) <= a or b;
    layer0_outputs(1539) <= not a;
    layer0_outputs(1540) <= a or b;
    layer0_outputs(1541) <= not b;
    layer0_outputs(1542) <= a and not b;
    layer0_outputs(1543) <= a;
    layer0_outputs(1544) <= b;
    layer0_outputs(1545) <= not a;
    layer0_outputs(1546) <= b;
    layer0_outputs(1547) <= b and not a;
    layer0_outputs(1548) <= not b or a;
    layer0_outputs(1549) <= not (a or b);
    layer0_outputs(1550) <= not a;
    layer0_outputs(1551) <= not b;
    layer0_outputs(1552) <= a xor b;
    layer0_outputs(1553) <= a and b;
    layer0_outputs(1554) <= not b;
    layer0_outputs(1555) <= not b or a;
    layer0_outputs(1556) <= a or b;
    layer0_outputs(1557) <= not a;
    layer0_outputs(1558) <= not b or a;
    layer0_outputs(1559) <= not (a or b);
    layer0_outputs(1560) <= not (a or b);
    layer0_outputs(1561) <= not b;
    layer0_outputs(1562) <= b;
    layer0_outputs(1563) <= a and not b;
    layer0_outputs(1564) <= not (a or b);
    layer0_outputs(1565) <= not (a or b);
    layer0_outputs(1566) <= a or b;
    layer0_outputs(1567) <= a;
    layer0_outputs(1568) <= not (a xor b);
    layer0_outputs(1569) <= not (a xor b);
    layer0_outputs(1570) <= a or b;
    layer0_outputs(1571) <= b and not a;
    layer0_outputs(1572) <= b;
    layer0_outputs(1573) <= b;
    layer0_outputs(1574) <= not b;
    layer0_outputs(1575) <= not (a xor b);
    layer0_outputs(1576) <= not a or b;
    layer0_outputs(1577) <= a and not b;
    layer0_outputs(1578) <= not (a or b);
    layer0_outputs(1579) <= not b;
    layer0_outputs(1580) <= b;
    layer0_outputs(1581) <= not a;
    layer0_outputs(1582) <= not b or a;
    layer0_outputs(1583) <= not (a or b);
    layer0_outputs(1584) <= a and b;
    layer0_outputs(1585) <= not (a or b);
    layer0_outputs(1586) <= a and not b;
    layer0_outputs(1587) <= a or b;
    layer0_outputs(1588) <= not b or a;
    layer0_outputs(1589) <= a xor b;
    layer0_outputs(1590) <= not a or b;
    layer0_outputs(1591) <= not a;
    layer0_outputs(1592) <= 1'b0;
    layer0_outputs(1593) <= not (a xor b);
    layer0_outputs(1594) <= a;
    layer0_outputs(1595) <= b;
    layer0_outputs(1596) <= not a;
    layer0_outputs(1597) <= not b;
    layer0_outputs(1598) <= not (a and b);
    layer0_outputs(1599) <= a;
    layer0_outputs(1600) <= not b or a;
    layer0_outputs(1601) <= not (a xor b);
    layer0_outputs(1602) <= a and not b;
    layer0_outputs(1603) <= a xor b;
    layer0_outputs(1604) <= a;
    layer0_outputs(1605) <= a or b;
    layer0_outputs(1606) <= a or b;
    layer0_outputs(1607) <= 1'b0;
    layer0_outputs(1608) <= a and not b;
    layer0_outputs(1609) <= not b or a;
    layer0_outputs(1610) <= b;
    layer0_outputs(1611) <= not b;
    layer0_outputs(1612) <= a or b;
    layer0_outputs(1613) <= not (a or b);
    layer0_outputs(1614) <= 1'b0;
    layer0_outputs(1615) <= a and not b;
    layer0_outputs(1616) <= not a or b;
    layer0_outputs(1617) <= b and not a;
    layer0_outputs(1618) <= 1'b1;
    layer0_outputs(1619) <= b and not a;
    layer0_outputs(1620) <= not a;
    layer0_outputs(1621) <= not a;
    layer0_outputs(1622) <= not (a or b);
    layer0_outputs(1623) <= not b;
    layer0_outputs(1624) <= a xor b;
    layer0_outputs(1625) <= not (a or b);
    layer0_outputs(1626) <= b;
    layer0_outputs(1627) <= 1'b1;
    layer0_outputs(1628) <= b;
    layer0_outputs(1629) <= not b or a;
    layer0_outputs(1630) <= b and not a;
    layer0_outputs(1631) <= not a or b;
    layer0_outputs(1632) <= a and b;
    layer0_outputs(1633) <= not (a and b);
    layer0_outputs(1634) <= not b or a;
    layer0_outputs(1635) <= a xor b;
    layer0_outputs(1636) <= a and not b;
    layer0_outputs(1637) <= b and not a;
    layer0_outputs(1638) <= b and not a;
    layer0_outputs(1639) <= a;
    layer0_outputs(1640) <= not a or b;
    layer0_outputs(1641) <= not (a or b);
    layer0_outputs(1642) <= not a or b;
    layer0_outputs(1643) <= not a;
    layer0_outputs(1644) <= b and not a;
    layer0_outputs(1645) <= b;
    layer0_outputs(1646) <= not b;
    layer0_outputs(1647) <= a or b;
    layer0_outputs(1648) <= not a;
    layer0_outputs(1649) <= b and not a;
    layer0_outputs(1650) <= not a;
    layer0_outputs(1651) <= a and b;
    layer0_outputs(1652) <= not a;
    layer0_outputs(1653) <= not b or a;
    layer0_outputs(1654) <= a and not b;
    layer0_outputs(1655) <= a and not b;
    layer0_outputs(1656) <= a;
    layer0_outputs(1657) <= b and not a;
    layer0_outputs(1658) <= not b or a;
    layer0_outputs(1659) <= a or b;
    layer0_outputs(1660) <= not a;
    layer0_outputs(1661) <= not a;
    layer0_outputs(1662) <= not a or b;
    layer0_outputs(1663) <= not a or b;
    layer0_outputs(1664) <= not b;
    layer0_outputs(1665) <= not b;
    layer0_outputs(1666) <= a xor b;
    layer0_outputs(1667) <= not (a xor b);
    layer0_outputs(1668) <= a or b;
    layer0_outputs(1669) <= not b or a;
    layer0_outputs(1670) <= b;
    layer0_outputs(1671) <= a;
    layer0_outputs(1672) <= a and not b;
    layer0_outputs(1673) <= not a;
    layer0_outputs(1674) <= a;
    layer0_outputs(1675) <= a;
    layer0_outputs(1676) <= b and not a;
    layer0_outputs(1677) <= not a or b;
    layer0_outputs(1678) <= 1'b1;
    layer0_outputs(1679) <= not a;
    layer0_outputs(1680) <= not b;
    layer0_outputs(1681) <= not b;
    layer0_outputs(1682) <= 1'b0;
    layer0_outputs(1683) <= a or b;
    layer0_outputs(1684) <= a and not b;
    layer0_outputs(1685) <= not b;
    layer0_outputs(1686) <= b;
    layer0_outputs(1687) <= a or b;
    layer0_outputs(1688) <= b;
    layer0_outputs(1689) <= b;
    layer0_outputs(1690) <= b and not a;
    layer0_outputs(1691) <= not b;
    layer0_outputs(1692) <= a or b;
    layer0_outputs(1693) <= not (a or b);
    layer0_outputs(1694) <= b;
    layer0_outputs(1695) <= a and not b;
    layer0_outputs(1696) <= a or b;
    layer0_outputs(1697) <= not b;
    layer0_outputs(1698) <= a and not b;
    layer0_outputs(1699) <= not (a xor b);
    layer0_outputs(1700) <= not a;
    layer0_outputs(1701) <= not (a or b);
    layer0_outputs(1702) <= 1'b1;
    layer0_outputs(1703) <= not (a and b);
    layer0_outputs(1704) <= a and not b;
    layer0_outputs(1705) <= b;
    layer0_outputs(1706) <= not (a or b);
    layer0_outputs(1707) <= b;
    layer0_outputs(1708) <= a xor b;
    layer0_outputs(1709) <= not (a or b);
    layer0_outputs(1710) <= not a;
    layer0_outputs(1711) <= b;
    layer0_outputs(1712) <= b;
    layer0_outputs(1713) <= not (a or b);
    layer0_outputs(1714) <= not a or b;
    layer0_outputs(1715) <= not b or a;
    layer0_outputs(1716) <= not a or b;
    layer0_outputs(1717) <= not (a xor b);
    layer0_outputs(1718) <= not (a or b);
    layer0_outputs(1719) <= 1'b1;
    layer0_outputs(1720) <= not a;
    layer0_outputs(1721) <= not b;
    layer0_outputs(1722) <= a;
    layer0_outputs(1723) <= not b;
    layer0_outputs(1724) <= not b;
    layer0_outputs(1725) <= not a;
    layer0_outputs(1726) <= not (a xor b);
    layer0_outputs(1727) <= not (a and b);
    layer0_outputs(1728) <= not (a or b);
    layer0_outputs(1729) <= not b or a;
    layer0_outputs(1730) <= b and not a;
    layer0_outputs(1731) <= not (a or b);
    layer0_outputs(1732) <= b;
    layer0_outputs(1733) <= not a or b;
    layer0_outputs(1734) <= a or b;
    layer0_outputs(1735) <= b and not a;
    layer0_outputs(1736) <= not (a xor b);
    layer0_outputs(1737) <= a or b;
    layer0_outputs(1738) <= not (a or b);
    layer0_outputs(1739) <= a or b;
    layer0_outputs(1740) <= not b;
    layer0_outputs(1741) <= not (a or b);
    layer0_outputs(1742) <= a;
    layer0_outputs(1743) <= not a or b;
    layer0_outputs(1744) <= a and not b;
    layer0_outputs(1745) <= a and b;
    layer0_outputs(1746) <= b and not a;
    layer0_outputs(1747) <= not (a xor b);
    layer0_outputs(1748) <= 1'b1;
    layer0_outputs(1749) <= not (a or b);
    layer0_outputs(1750) <= a or b;
    layer0_outputs(1751) <= not (a xor b);
    layer0_outputs(1752) <= b;
    layer0_outputs(1753) <= not a or b;
    layer0_outputs(1754) <= not b;
    layer0_outputs(1755) <= b and not a;
    layer0_outputs(1756) <= not (a and b);
    layer0_outputs(1757) <= a xor b;
    layer0_outputs(1758) <= b;
    layer0_outputs(1759) <= not a;
    layer0_outputs(1760) <= a or b;
    layer0_outputs(1761) <= b;
    layer0_outputs(1762) <= not a;
    layer0_outputs(1763) <= not (a or b);
    layer0_outputs(1764) <= a xor b;
    layer0_outputs(1765) <= not (a or b);
    layer0_outputs(1766) <= not a or b;
    layer0_outputs(1767) <= b and not a;
    layer0_outputs(1768) <= b and not a;
    layer0_outputs(1769) <= not a or b;
    layer0_outputs(1770) <= a;
    layer0_outputs(1771) <= b;
    layer0_outputs(1772) <= b and not a;
    layer0_outputs(1773) <= a and not b;
    layer0_outputs(1774) <= a;
    layer0_outputs(1775) <= not b or a;
    layer0_outputs(1776) <= b and not a;
    layer0_outputs(1777) <= a and b;
    layer0_outputs(1778) <= a or b;
    layer0_outputs(1779) <= not b;
    layer0_outputs(1780) <= a or b;
    layer0_outputs(1781) <= not a or b;
    layer0_outputs(1782) <= 1'b1;
    layer0_outputs(1783) <= not a or b;
    layer0_outputs(1784) <= not (a xor b);
    layer0_outputs(1785) <= not a or b;
    layer0_outputs(1786) <= 1'b0;
    layer0_outputs(1787) <= not (a or b);
    layer0_outputs(1788) <= not b;
    layer0_outputs(1789) <= not (a or b);
    layer0_outputs(1790) <= not a;
    layer0_outputs(1791) <= b and not a;
    layer0_outputs(1792) <= a;
    layer0_outputs(1793) <= not b or a;
    layer0_outputs(1794) <= not (a or b);
    layer0_outputs(1795) <= a and not b;
    layer0_outputs(1796) <= not b or a;
    layer0_outputs(1797) <= not (a xor b);
    layer0_outputs(1798) <= not (a or b);
    layer0_outputs(1799) <= not (a or b);
    layer0_outputs(1800) <= a;
    layer0_outputs(1801) <= 1'b0;
    layer0_outputs(1802) <= not (a or b);
    layer0_outputs(1803) <= 1'b1;
    layer0_outputs(1804) <= a or b;
    layer0_outputs(1805) <= a xor b;
    layer0_outputs(1806) <= a or b;
    layer0_outputs(1807) <= a or b;
    layer0_outputs(1808) <= b and not a;
    layer0_outputs(1809) <= a or b;
    layer0_outputs(1810) <= not (a or b);
    layer0_outputs(1811) <= not b or a;
    layer0_outputs(1812) <= not a;
    layer0_outputs(1813) <= a or b;
    layer0_outputs(1814) <= a xor b;
    layer0_outputs(1815) <= a or b;
    layer0_outputs(1816) <= a or b;
    layer0_outputs(1817) <= not b;
    layer0_outputs(1818) <= not (a or b);
    layer0_outputs(1819) <= not (a or b);
    layer0_outputs(1820) <= a or b;
    layer0_outputs(1821) <= a or b;
    layer0_outputs(1822) <= not b or a;
    layer0_outputs(1823) <= 1'b1;
    layer0_outputs(1824) <= not a;
    layer0_outputs(1825) <= a xor b;
    layer0_outputs(1826) <= a;
    layer0_outputs(1827) <= b;
    layer0_outputs(1828) <= not (a xor b);
    layer0_outputs(1829) <= b and not a;
    layer0_outputs(1830) <= not b or a;
    layer0_outputs(1831) <= 1'b0;
    layer0_outputs(1832) <= not (a xor b);
    layer0_outputs(1833) <= b;
    layer0_outputs(1834) <= b and not a;
    layer0_outputs(1835) <= a or b;
    layer0_outputs(1836) <= not b or a;
    layer0_outputs(1837) <= 1'b1;
    layer0_outputs(1838) <= not b;
    layer0_outputs(1839) <= not (a and b);
    layer0_outputs(1840) <= not b;
    layer0_outputs(1841) <= a;
    layer0_outputs(1842) <= not (a or b);
    layer0_outputs(1843) <= a xor b;
    layer0_outputs(1844) <= a xor b;
    layer0_outputs(1845) <= 1'b1;
    layer0_outputs(1846) <= a or b;
    layer0_outputs(1847) <= a or b;
    layer0_outputs(1848) <= a and not b;
    layer0_outputs(1849) <= not b or a;
    layer0_outputs(1850) <= 1'b0;
    layer0_outputs(1851) <= not (a or b);
    layer0_outputs(1852) <= b and not a;
    layer0_outputs(1853) <= not b;
    layer0_outputs(1854) <= not (a or b);
    layer0_outputs(1855) <= b and not a;
    layer0_outputs(1856) <= not b;
    layer0_outputs(1857) <= not (a or b);
    layer0_outputs(1858) <= a or b;
    layer0_outputs(1859) <= not a;
    layer0_outputs(1860) <= not (a xor b);
    layer0_outputs(1861) <= not a;
    layer0_outputs(1862) <= b;
    layer0_outputs(1863) <= not b;
    layer0_outputs(1864) <= a or b;
    layer0_outputs(1865) <= a xor b;
    layer0_outputs(1866) <= b;
    layer0_outputs(1867) <= not a or b;
    layer0_outputs(1868) <= 1'b1;
    layer0_outputs(1869) <= not a;
    layer0_outputs(1870) <= not a;
    layer0_outputs(1871) <= not a;
    layer0_outputs(1872) <= not b;
    layer0_outputs(1873) <= b;
    layer0_outputs(1874) <= not (a or b);
    layer0_outputs(1875) <= a;
    layer0_outputs(1876) <= a or b;
    layer0_outputs(1877) <= not a or b;
    layer0_outputs(1878) <= not a or b;
    layer0_outputs(1879) <= a;
    layer0_outputs(1880) <= not b;
    layer0_outputs(1881) <= a xor b;
    layer0_outputs(1882) <= not (a or b);
    layer0_outputs(1883) <= not b;
    layer0_outputs(1884) <= not b;
    layer0_outputs(1885) <= a or b;
    layer0_outputs(1886) <= not (a xor b);
    layer0_outputs(1887) <= not a or b;
    layer0_outputs(1888) <= b;
    layer0_outputs(1889) <= not b;
    layer0_outputs(1890) <= not b;
    layer0_outputs(1891) <= a;
    layer0_outputs(1892) <= not a;
    layer0_outputs(1893) <= a;
    layer0_outputs(1894) <= not (a or b);
    layer0_outputs(1895) <= a;
    layer0_outputs(1896) <= not b or a;
    layer0_outputs(1897) <= a and not b;
    layer0_outputs(1898) <= a and b;
    layer0_outputs(1899) <= a;
    layer0_outputs(1900) <= not a or b;
    layer0_outputs(1901) <= 1'b0;
    layer0_outputs(1902) <= not (a xor b);
    layer0_outputs(1903) <= a;
    layer0_outputs(1904) <= 1'b1;
    layer0_outputs(1905) <= not a;
    layer0_outputs(1906) <= not b;
    layer0_outputs(1907) <= a;
    layer0_outputs(1908) <= not a or b;
    layer0_outputs(1909) <= not a;
    layer0_outputs(1910) <= not a or b;
    layer0_outputs(1911) <= a and b;
    layer0_outputs(1912) <= a xor b;
    layer0_outputs(1913) <= not (a xor b);
    layer0_outputs(1914) <= not a;
    layer0_outputs(1915) <= not (a or b);
    layer0_outputs(1916) <= a or b;
    layer0_outputs(1917) <= not (a or b);
    layer0_outputs(1918) <= a and not b;
    layer0_outputs(1919) <= not (a xor b);
    layer0_outputs(1920) <= a or b;
    layer0_outputs(1921) <= not (a xor b);
    layer0_outputs(1922) <= a or b;
    layer0_outputs(1923) <= not a or b;
    layer0_outputs(1924) <= a;
    layer0_outputs(1925) <= not (a or b);
    layer0_outputs(1926) <= not a;
    layer0_outputs(1927) <= a and not b;
    layer0_outputs(1928) <= a or b;
    layer0_outputs(1929) <= a and not b;
    layer0_outputs(1930) <= b;
    layer0_outputs(1931) <= a;
    layer0_outputs(1932) <= not (a and b);
    layer0_outputs(1933) <= not b or a;
    layer0_outputs(1934) <= not b;
    layer0_outputs(1935) <= a or b;
    layer0_outputs(1936) <= not (a xor b);
    layer0_outputs(1937) <= not (a xor b);
    layer0_outputs(1938) <= b and not a;
    layer0_outputs(1939) <= not (a xor b);
    layer0_outputs(1940) <= b;
    layer0_outputs(1941) <= not (a xor b);
    layer0_outputs(1942) <= a and b;
    layer0_outputs(1943) <= a and not b;
    layer0_outputs(1944) <= b and not a;
    layer0_outputs(1945) <= not b;
    layer0_outputs(1946) <= not (a or b);
    layer0_outputs(1947) <= not (a or b);
    layer0_outputs(1948) <= not b;
    layer0_outputs(1949) <= a or b;
    layer0_outputs(1950) <= 1'b1;
    layer0_outputs(1951) <= a;
    layer0_outputs(1952) <= not a or b;
    layer0_outputs(1953) <= b;
    layer0_outputs(1954) <= a;
    layer0_outputs(1955) <= b;
    layer0_outputs(1956) <= not a;
    layer0_outputs(1957) <= not b;
    layer0_outputs(1958) <= a or b;
    layer0_outputs(1959) <= not (a or b);
    layer0_outputs(1960) <= not (a xor b);
    layer0_outputs(1961) <= not (a and b);
    layer0_outputs(1962) <= not b or a;
    layer0_outputs(1963) <= 1'b1;
    layer0_outputs(1964) <= not b;
    layer0_outputs(1965) <= not b;
    layer0_outputs(1966) <= b;
    layer0_outputs(1967) <= a;
    layer0_outputs(1968) <= a or b;
    layer0_outputs(1969) <= not b;
    layer0_outputs(1970) <= not (a or b);
    layer0_outputs(1971) <= a and not b;
    layer0_outputs(1972) <= b;
    layer0_outputs(1973) <= a or b;
    layer0_outputs(1974) <= not a;
    layer0_outputs(1975) <= a and b;
    layer0_outputs(1976) <= not (a or b);
    layer0_outputs(1977) <= not b;
    layer0_outputs(1978) <= a;
    layer0_outputs(1979) <= a xor b;
    layer0_outputs(1980) <= 1'b0;
    layer0_outputs(1981) <= a or b;
    layer0_outputs(1982) <= not b or a;
    layer0_outputs(1983) <= a and not b;
    layer0_outputs(1984) <= a and not b;
    layer0_outputs(1985) <= not (a and b);
    layer0_outputs(1986) <= 1'b0;
    layer0_outputs(1987) <= b and not a;
    layer0_outputs(1988) <= a and not b;
    layer0_outputs(1989) <= a or b;
    layer0_outputs(1990) <= a or b;
    layer0_outputs(1991) <= not b;
    layer0_outputs(1992) <= not b;
    layer0_outputs(1993) <= not (a xor b);
    layer0_outputs(1994) <= not a or b;
    layer0_outputs(1995) <= a or b;
    layer0_outputs(1996) <= a and not b;
    layer0_outputs(1997) <= not b or a;
    layer0_outputs(1998) <= not b or a;
    layer0_outputs(1999) <= not a;
    layer0_outputs(2000) <= 1'b0;
    layer0_outputs(2001) <= a;
    layer0_outputs(2002) <= a xor b;
    layer0_outputs(2003) <= a or b;
    layer0_outputs(2004) <= not b or a;
    layer0_outputs(2005) <= b and not a;
    layer0_outputs(2006) <= 1'b1;
    layer0_outputs(2007) <= not (a or b);
    layer0_outputs(2008) <= b;
    layer0_outputs(2009) <= 1'b0;
    layer0_outputs(2010) <= not b or a;
    layer0_outputs(2011) <= not a or b;
    layer0_outputs(2012) <= a or b;
    layer0_outputs(2013) <= a;
    layer0_outputs(2014) <= a and not b;
    layer0_outputs(2015) <= a and not b;
    layer0_outputs(2016) <= not b;
    layer0_outputs(2017) <= not a;
    layer0_outputs(2018) <= b;
    layer0_outputs(2019) <= b;
    layer0_outputs(2020) <= not b;
    layer0_outputs(2021) <= a;
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= a or b;
    layer0_outputs(2024) <= a xor b;
    layer0_outputs(2025) <= not b;
    layer0_outputs(2026) <= not (a or b);
    layer0_outputs(2027) <= a xor b;
    layer0_outputs(2028) <= a or b;
    layer0_outputs(2029) <= not (a and b);
    layer0_outputs(2030) <= not (a or b);
    layer0_outputs(2031) <= not a;
    layer0_outputs(2032) <= not (a and b);
    layer0_outputs(2033) <= 1'b0;
    layer0_outputs(2034) <= not b;
    layer0_outputs(2035) <= a;
    layer0_outputs(2036) <= a and not b;
    layer0_outputs(2037) <= not (a or b);
    layer0_outputs(2038) <= a;
    layer0_outputs(2039) <= a or b;
    layer0_outputs(2040) <= a xor b;
    layer0_outputs(2041) <= a and b;
    layer0_outputs(2042) <= not a;
    layer0_outputs(2043) <= a and not b;
    layer0_outputs(2044) <= not a or b;
    layer0_outputs(2045) <= a and not b;
    layer0_outputs(2046) <= a;
    layer0_outputs(2047) <= not a or b;
    layer0_outputs(2048) <= not b or a;
    layer0_outputs(2049) <= not a or b;
    layer0_outputs(2050) <= b;
    layer0_outputs(2051) <= a and b;
    layer0_outputs(2052) <= a or b;
    layer0_outputs(2053) <= b and not a;
    layer0_outputs(2054) <= a and not b;
    layer0_outputs(2055) <= a;
    layer0_outputs(2056) <= b and not a;
    layer0_outputs(2057) <= a;
    layer0_outputs(2058) <= not (a xor b);
    layer0_outputs(2059) <= a and b;
    layer0_outputs(2060) <= b and not a;
    layer0_outputs(2061) <= 1'b1;
    layer0_outputs(2062) <= a or b;
    layer0_outputs(2063) <= b;
    layer0_outputs(2064) <= not b;
    layer0_outputs(2065) <= not a or b;
    layer0_outputs(2066) <= a or b;
    layer0_outputs(2067) <= not b or a;
    layer0_outputs(2068) <= a;
    layer0_outputs(2069) <= a and not b;
    layer0_outputs(2070) <= b and not a;
    layer0_outputs(2071) <= not b or a;
    layer0_outputs(2072) <= 1'b1;
    layer0_outputs(2073) <= b and not a;
    layer0_outputs(2074) <= a and b;
    layer0_outputs(2075) <= 1'b1;
    layer0_outputs(2076) <= b and not a;
    layer0_outputs(2077) <= not b;
    layer0_outputs(2078) <= a or b;
    layer0_outputs(2079) <= a or b;
    layer0_outputs(2080) <= not (a or b);
    layer0_outputs(2081) <= b and not a;
    layer0_outputs(2082) <= b and not a;
    layer0_outputs(2083) <= a xor b;
    layer0_outputs(2084) <= not a or b;
    layer0_outputs(2085) <= b and not a;
    layer0_outputs(2086) <= a;
    layer0_outputs(2087) <= b;
    layer0_outputs(2088) <= b and not a;
    layer0_outputs(2089) <= a or b;
    layer0_outputs(2090) <= not b;
    layer0_outputs(2091) <= a and not b;
    layer0_outputs(2092) <= a or b;
    layer0_outputs(2093) <= not (a xor b);
    layer0_outputs(2094) <= a;
    layer0_outputs(2095) <= not a or b;
    layer0_outputs(2096) <= not (a or b);
    layer0_outputs(2097) <= not (a xor b);
    layer0_outputs(2098) <= a or b;
    layer0_outputs(2099) <= not (a or b);
    layer0_outputs(2100) <= not (a xor b);
    layer0_outputs(2101) <= b;
    layer0_outputs(2102) <= b;
    layer0_outputs(2103) <= not (a or b);
    layer0_outputs(2104) <= b and not a;
    layer0_outputs(2105) <= 1'b0;
    layer0_outputs(2106) <= b and not a;
    layer0_outputs(2107) <= not (a or b);
    layer0_outputs(2108) <= a or b;
    layer0_outputs(2109) <= a;
    layer0_outputs(2110) <= a or b;
    layer0_outputs(2111) <= not (a and b);
    layer0_outputs(2112) <= 1'b0;
    layer0_outputs(2113) <= not (a or b);
    layer0_outputs(2114) <= not a;
    layer0_outputs(2115) <= a;
    layer0_outputs(2116) <= not (a or b);
    layer0_outputs(2117) <= not a;
    layer0_outputs(2118) <= b;
    layer0_outputs(2119) <= not a or b;
    layer0_outputs(2120) <= a or b;
    layer0_outputs(2121) <= a xor b;
    layer0_outputs(2122) <= b and not a;
    layer0_outputs(2123) <= not b;
    layer0_outputs(2124) <= a xor b;
    layer0_outputs(2125) <= b and not a;
    layer0_outputs(2126) <= not a;
    layer0_outputs(2127) <= not a;
    layer0_outputs(2128) <= a and not b;
    layer0_outputs(2129) <= a and not b;
    layer0_outputs(2130) <= not (a or b);
    layer0_outputs(2131) <= not a or b;
    layer0_outputs(2132) <= not a;
    layer0_outputs(2133) <= 1'b1;
    layer0_outputs(2134) <= b;
    layer0_outputs(2135) <= a and not b;
    layer0_outputs(2136) <= a or b;
    layer0_outputs(2137) <= a xor b;
    layer0_outputs(2138) <= not b;
    layer0_outputs(2139) <= not (a or b);
    layer0_outputs(2140) <= not (a xor b);
    layer0_outputs(2141) <= a or b;
    layer0_outputs(2142) <= not (a xor b);
    layer0_outputs(2143) <= not a;
    layer0_outputs(2144) <= not a or b;
    layer0_outputs(2145) <= b;
    layer0_outputs(2146) <= a;
    layer0_outputs(2147) <= a xor b;
    layer0_outputs(2148) <= a xor b;
    layer0_outputs(2149) <= a and not b;
    layer0_outputs(2150) <= not a;
    layer0_outputs(2151) <= not a;
    layer0_outputs(2152) <= a or b;
    layer0_outputs(2153) <= a and not b;
    layer0_outputs(2154) <= 1'b0;
    layer0_outputs(2155) <= b and not a;
    layer0_outputs(2156) <= b;
    layer0_outputs(2157) <= not b or a;
    layer0_outputs(2158) <= not a;
    layer0_outputs(2159) <= a xor b;
    layer0_outputs(2160) <= not a or b;
    layer0_outputs(2161) <= not (a or b);
    layer0_outputs(2162) <= not (a xor b);
    layer0_outputs(2163) <= not (a xor b);
    layer0_outputs(2164) <= a;
    layer0_outputs(2165) <= b;
    layer0_outputs(2166) <= a or b;
    layer0_outputs(2167) <= not (a or b);
    layer0_outputs(2168) <= a or b;
    layer0_outputs(2169) <= not (a or b);
    layer0_outputs(2170) <= a;
    layer0_outputs(2171) <= a;
    layer0_outputs(2172) <= a and not b;
    layer0_outputs(2173) <= b;
    layer0_outputs(2174) <= a or b;
    layer0_outputs(2175) <= a;
    layer0_outputs(2176) <= b;
    layer0_outputs(2177) <= a or b;
    layer0_outputs(2178) <= a xor b;
    layer0_outputs(2179) <= a and b;
    layer0_outputs(2180) <= a or b;
    layer0_outputs(2181) <= not (a or b);
    layer0_outputs(2182) <= not a;
    layer0_outputs(2183) <= a or b;
    layer0_outputs(2184) <= not (a or b);
    layer0_outputs(2185) <= 1'b1;
    layer0_outputs(2186) <= a;
    layer0_outputs(2187) <= not (a xor b);
    layer0_outputs(2188) <= not a;
    layer0_outputs(2189) <= b;
    layer0_outputs(2190) <= a xor b;
    layer0_outputs(2191) <= a xor b;
    layer0_outputs(2192) <= not a;
    layer0_outputs(2193) <= a or b;
    layer0_outputs(2194) <= not b;
    layer0_outputs(2195) <= not (a or b);
    layer0_outputs(2196) <= not (a or b);
    layer0_outputs(2197) <= not (a or b);
    layer0_outputs(2198) <= not (a or b);
    layer0_outputs(2199) <= a and not b;
    layer0_outputs(2200) <= not b or a;
    layer0_outputs(2201) <= not (a or b);
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= not (a or b);
    layer0_outputs(2204) <= not a;
    layer0_outputs(2205) <= not (a xor b);
    layer0_outputs(2206) <= b and not a;
    layer0_outputs(2207) <= not (a or b);
    layer0_outputs(2208) <= not (a and b);
    layer0_outputs(2209) <= not b;
    layer0_outputs(2210) <= not (a xor b);
    layer0_outputs(2211) <= not (a and b);
    layer0_outputs(2212) <= a xor b;
    layer0_outputs(2213) <= b;
    layer0_outputs(2214) <= not b;
    layer0_outputs(2215) <= a or b;
    layer0_outputs(2216) <= not b or a;
    layer0_outputs(2217) <= a or b;
    layer0_outputs(2218) <= a xor b;
    layer0_outputs(2219) <= a;
    layer0_outputs(2220) <= not b or a;
    layer0_outputs(2221) <= a;
    layer0_outputs(2222) <= not (a and b);
    layer0_outputs(2223) <= not (a or b);
    layer0_outputs(2224) <= a;
    layer0_outputs(2225) <= not a;
    layer0_outputs(2226) <= not a or b;
    layer0_outputs(2227) <= not a;
    layer0_outputs(2228) <= a xor b;
    layer0_outputs(2229) <= a;
    layer0_outputs(2230) <= not b or a;
    layer0_outputs(2231) <= not (a and b);
    layer0_outputs(2232) <= not a;
    layer0_outputs(2233) <= a;
    layer0_outputs(2234) <= 1'b1;
    layer0_outputs(2235) <= a;
    layer0_outputs(2236) <= a and not b;
    layer0_outputs(2237) <= not (a xor b);
    layer0_outputs(2238) <= b and not a;
    layer0_outputs(2239) <= not a or b;
    layer0_outputs(2240) <= a;
    layer0_outputs(2241) <= not (a or b);
    layer0_outputs(2242) <= a and not b;
    layer0_outputs(2243) <= not b or a;
    layer0_outputs(2244) <= a;
    layer0_outputs(2245) <= not a;
    layer0_outputs(2246) <= not b;
    layer0_outputs(2247) <= a or b;
    layer0_outputs(2248) <= a xor b;
    layer0_outputs(2249) <= not b;
    layer0_outputs(2250) <= not (a xor b);
    layer0_outputs(2251) <= b;
    layer0_outputs(2252) <= not a or b;
    layer0_outputs(2253) <= a or b;
    layer0_outputs(2254) <= not b or a;
    layer0_outputs(2255) <= not (a xor b);
    layer0_outputs(2256) <= a xor b;
    layer0_outputs(2257) <= not (a xor b);
    layer0_outputs(2258) <= not b or a;
    layer0_outputs(2259) <= not (a or b);
    layer0_outputs(2260) <= a and not b;
    layer0_outputs(2261) <= b;
    layer0_outputs(2262) <= not (a or b);
    layer0_outputs(2263) <= a or b;
    layer0_outputs(2264) <= a or b;
    layer0_outputs(2265) <= not a or b;
    layer0_outputs(2266) <= a or b;
    layer0_outputs(2267) <= a;
    layer0_outputs(2268) <= not (a and b);
    layer0_outputs(2269) <= not b or a;
    layer0_outputs(2270) <= not (a or b);
    layer0_outputs(2271) <= a xor b;
    layer0_outputs(2272) <= not (a or b);
    layer0_outputs(2273) <= not b or a;
    layer0_outputs(2274) <= a or b;
    layer0_outputs(2275) <= a;
    layer0_outputs(2276) <= a and b;
    layer0_outputs(2277) <= not (a or b);
    layer0_outputs(2278) <= not b or a;
    layer0_outputs(2279) <= a;
    layer0_outputs(2280) <= 1'b1;
    layer0_outputs(2281) <= not (a or b);
    layer0_outputs(2282) <= a;
    layer0_outputs(2283) <= a;
    layer0_outputs(2284) <= b;
    layer0_outputs(2285) <= b and not a;
    layer0_outputs(2286) <= a or b;
    layer0_outputs(2287) <= 1'b1;
    layer0_outputs(2288) <= not b;
    layer0_outputs(2289) <= a or b;
    layer0_outputs(2290) <= b;
    layer0_outputs(2291) <= b and not a;
    layer0_outputs(2292) <= a and not b;
    layer0_outputs(2293) <= not (a or b);
    layer0_outputs(2294) <= a or b;
    layer0_outputs(2295) <= not (a or b);
    layer0_outputs(2296) <= b;
    layer0_outputs(2297) <= a and not b;
    layer0_outputs(2298) <= not (a xor b);
    layer0_outputs(2299) <= not (a xor b);
    layer0_outputs(2300) <= not a or b;
    layer0_outputs(2301) <= b;
    layer0_outputs(2302) <= 1'b0;
    layer0_outputs(2303) <= a xor b;
    layer0_outputs(2304) <= a or b;
    layer0_outputs(2305) <= a and b;
    layer0_outputs(2306) <= b;
    layer0_outputs(2307) <= b and not a;
    layer0_outputs(2308) <= not (a or b);
    layer0_outputs(2309) <= a and not b;
    layer0_outputs(2310) <= a xor b;
    layer0_outputs(2311) <= not b;
    layer0_outputs(2312) <= b;
    layer0_outputs(2313) <= a or b;
    layer0_outputs(2314) <= b and not a;
    layer0_outputs(2315) <= a or b;
    layer0_outputs(2316) <= 1'b0;
    layer0_outputs(2317) <= a or b;
    layer0_outputs(2318) <= b and not a;
    layer0_outputs(2319) <= not b or a;
    layer0_outputs(2320) <= not a;
    layer0_outputs(2321) <= a and not b;
    layer0_outputs(2322) <= 1'b0;
    layer0_outputs(2323) <= not (a and b);
    layer0_outputs(2324) <= a and not b;
    layer0_outputs(2325) <= b;
    layer0_outputs(2326) <= not (a and b);
    layer0_outputs(2327) <= not (a or b);
    layer0_outputs(2328) <= not a or b;
    layer0_outputs(2329) <= b;
    layer0_outputs(2330) <= not b;
    layer0_outputs(2331) <= b and not a;
    layer0_outputs(2332) <= b;
    layer0_outputs(2333) <= b;
    layer0_outputs(2334) <= not (a or b);
    layer0_outputs(2335) <= not (a or b);
    layer0_outputs(2336) <= b;
    layer0_outputs(2337) <= a or b;
    layer0_outputs(2338) <= not (a or b);
    layer0_outputs(2339) <= not (a or b);
    layer0_outputs(2340) <= a xor b;
    layer0_outputs(2341) <= not b;
    layer0_outputs(2342) <= not (a or b);
    layer0_outputs(2343) <= not (a and b);
    layer0_outputs(2344) <= 1'b1;
    layer0_outputs(2345) <= 1'b0;
    layer0_outputs(2346) <= b and not a;
    layer0_outputs(2347) <= not a or b;
    layer0_outputs(2348) <= not b;
    layer0_outputs(2349) <= not (a or b);
    layer0_outputs(2350) <= a or b;
    layer0_outputs(2351) <= a;
    layer0_outputs(2352) <= not b;
    layer0_outputs(2353) <= a or b;
    layer0_outputs(2354) <= b;
    layer0_outputs(2355) <= a or b;
    layer0_outputs(2356) <= a;
    layer0_outputs(2357) <= 1'b1;
    layer0_outputs(2358) <= not b;
    layer0_outputs(2359) <= not (a or b);
    layer0_outputs(2360) <= a xor b;
    layer0_outputs(2361) <= a and not b;
    layer0_outputs(2362) <= not a;
    layer0_outputs(2363) <= a or b;
    layer0_outputs(2364) <= a and b;
    layer0_outputs(2365) <= b;
    layer0_outputs(2366) <= b and not a;
    layer0_outputs(2367) <= a or b;
    layer0_outputs(2368) <= a and not b;
    layer0_outputs(2369) <= not a;
    layer0_outputs(2370) <= not b or a;
    layer0_outputs(2371) <= not a or b;
    layer0_outputs(2372) <= not (a or b);
    layer0_outputs(2373) <= a and not b;
    layer0_outputs(2374) <= a or b;
    layer0_outputs(2375) <= not a or b;
    layer0_outputs(2376) <= a and b;
    layer0_outputs(2377) <= not b;
    layer0_outputs(2378) <= not (a and b);
    layer0_outputs(2379) <= a or b;
    layer0_outputs(2380) <= not (a or b);
    layer0_outputs(2381) <= a;
    layer0_outputs(2382) <= a and not b;
    layer0_outputs(2383) <= 1'b1;
    layer0_outputs(2384) <= not a;
    layer0_outputs(2385) <= not b;
    layer0_outputs(2386) <= 1'b0;
    layer0_outputs(2387) <= b;
    layer0_outputs(2388) <= a xor b;
    layer0_outputs(2389) <= not (a or b);
    layer0_outputs(2390) <= b;
    layer0_outputs(2391) <= not (a or b);
    layer0_outputs(2392) <= not b or a;
    layer0_outputs(2393) <= not a;
    layer0_outputs(2394) <= a and not b;
    layer0_outputs(2395) <= a and b;
    layer0_outputs(2396) <= a or b;
    layer0_outputs(2397) <= not (a xor b);
    layer0_outputs(2398) <= b;
    layer0_outputs(2399) <= a and not b;
    layer0_outputs(2400) <= not a;
    layer0_outputs(2401) <= not (a xor b);
    layer0_outputs(2402) <= not b;
    layer0_outputs(2403) <= a and not b;
    layer0_outputs(2404) <= a or b;
    layer0_outputs(2405) <= a;
    layer0_outputs(2406) <= not b or a;
    layer0_outputs(2407) <= not b;
    layer0_outputs(2408) <= not a or b;
    layer0_outputs(2409) <= not a;
    layer0_outputs(2410) <= not a or b;
    layer0_outputs(2411) <= not (a or b);
    layer0_outputs(2412) <= not b or a;
    layer0_outputs(2413) <= not (a or b);
    layer0_outputs(2414) <= a;
    layer0_outputs(2415) <= 1'b1;
    layer0_outputs(2416) <= b;
    layer0_outputs(2417) <= not (a xor b);
    layer0_outputs(2418) <= b and not a;
    layer0_outputs(2419) <= a or b;
    layer0_outputs(2420) <= not (a xor b);
    layer0_outputs(2421) <= b;
    layer0_outputs(2422) <= not a;
    layer0_outputs(2423) <= b;
    layer0_outputs(2424) <= not a or b;
    layer0_outputs(2425) <= not (a xor b);
    layer0_outputs(2426) <= b;
    layer0_outputs(2427) <= not (a or b);
    layer0_outputs(2428) <= not b;
    layer0_outputs(2429) <= not a or b;
    layer0_outputs(2430) <= not b;
    layer0_outputs(2431) <= not (a or b);
    layer0_outputs(2432) <= not b;
    layer0_outputs(2433) <= not a or b;
    layer0_outputs(2434) <= not b or a;
    layer0_outputs(2435) <= a xor b;
    layer0_outputs(2436) <= b;
    layer0_outputs(2437) <= a;
    layer0_outputs(2438) <= a;
    layer0_outputs(2439) <= b and not a;
    layer0_outputs(2440) <= b;
    layer0_outputs(2441) <= b;
    layer0_outputs(2442) <= not (a or b);
    layer0_outputs(2443) <= a;
    layer0_outputs(2444) <= b;
    layer0_outputs(2445) <= a and not b;
    layer0_outputs(2446) <= not b or a;
    layer0_outputs(2447) <= a and not b;
    layer0_outputs(2448) <= a or b;
    layer0_outputs(2449) <= not (a and b);
    layer0_outputs(2450) <= not (a or b);
    layer0_outputs(2451) <= a;
    layer0_outputs(2452) <= a and not b;
    layer0_outputs(2453) <= b;
    layer0_outputs(2454) <= not (a xor b);
    layer0_outputs(2455) <= not b;
    layer0_outputs(2456) <= 1'b1;
    layer0_outputs(2457) <= not (a or b);
    layer0_outputs(2458) <= a and not b;
    layer0_outputs(2459) <= a or b;
    layer0_outputs(2460) <= b and not a;
    layer0_outputs(2461) <= not a;
    layer0_outputs(2462) <= 1'b1;
    layer0_outputs(2463) <= a;
    layer0_outputs(2464) <= not a or b;
    layer0_outputs(2465) <= a and not b;
    layer0_outputs(2466) <= not b or a;
    layer0_outputs(2467) <= not (a or b);
    layer0_outputs(2468) <= not b;
    layer0_outputs(2469) <= a;
    layer0_outputs(2470) <= a or b;
    layer0_outputs(2471) <= not a;
    layer0_outputs(2472) <= b and not a;
    layer0_outputs(2473) <= b and not a;
    layer0_outputs(2474) <= a or b;
    layer0_outputs(2475) <= not (a xor b);
    layer0_outputs(2476) <= not b;
    layer0_outputs(2477) <= a;
    layer0_outputs(2478) <= not (a xor b);
    layer0_outputs(2479) <= b;
    layer0_outputs(2480) <= a;
    layer0_outputs(2481) <= not (a or b);
    layer0_outputs(2482) <= a or b;
    layer0_outputs(2483) <= not (a xor b);
    layer0_outputs(2484) <= not b or a;
    layer0_outputs(2485) <= not a;
    layer0_outputs(2486) <= not b or a;
    layer0_outputs(2487) <= not (a or b);
    layer0_outputs(2488) <= a or b;
    layer0_outputs(2489) <= a;
    layer0_outputs(2490) <= not b;
    layer0_outputs(2491) <= 1'b0;
    layer0_outputs(2492) <= not (a xor b);
    layer0_outputs(2493) <= not (a or b);
    layer0_outputs(2494) <= b;
    layer0_outputs(2495) <= not (a xor b);
    layer0_outputs(2496) <= a or b;
    layer0_outputs(2497) <= a and not b;
    layer0_outputs(2498) <= not b;
    layer0_outputs(2499) <= a or b;
    layer0_outputs(2500) <= a and not b;
    layer0_outputs(2501) <= b;
    layer0_outputs(2502) <= not (a or b);
    layer0_outputs(2503) <= not (a xor b);
    layer0_outputs(2504) <= a;
    layer0_outputs(2505) <= not (a or b);
    layer0_outputs(2506) <= a;
    layer0_outputs(2507) <= a or b;
    layer0_outputs(2508) <= not a;
    layer0_outputs(2509) <= a;
    layer0_outputs(2510) <= not (a xor b);
    layer0_outputs(2511) <= not b or a;
    layer0_outputs(2512) <= not (a or b);
    layer0_outputs(2513) <= not a;
    layer0_outputs(2514) <= a or b;
    layer0_outputs(2515) <= not (a or b);
    layer0_outputs(2516) <= not (a xor b);
    layer0_outputs(2517) <= not (a or b);
    layer0_outputs(2518) <= not b;
    layer0_outputs(2519) <= not (a or b);
    layer0_outputs(2520) <= b and not a;
    layer0_outputs(2521) <= a or b;
    layer0_outputs(2522) <= not a;
    layer0_outputs(2523) <= a and not b;
    layer0_outputs(2524) <= b;
    layer0_outputs(2525) <= a and not b;
    layer0_outputs(2526) <= not a or b;
    layer0_outputs(2527) <= a or b;
    layer0_outputs(2528) <= not b or a;
    layer0_outputs(2529) <= a;
    layer0_outputs(2530) <= not a;
    layer0_outputs(2531) <= b;
    layer0_outputs(2532) <= a xor b;
    layer0_outputs(2533) <= 1'b1;
    layer0_outputs(2534) <= not (a or b);
    layer0_outputs(2535) <= not b or a;
    layer0_outputs(2536) <= 1'b0;
    layer0_outputs(2537) <= not b;
    layer0_outputs(2538) <= not b;
    layer0_outputs(2539) <= not a or b;
    layer0_outputs(2540) <= not (a xor b);
    layer0_outputs(2541) <= a;
    layer0_outputs(2542) <= b;
    layer0_outputs(2543) <= a xor b;
    layer0_outputs(2544) <= not a;
    layer0_outputs(2545) <= not (a or b);
    layer0_outputs(2546) <= not a;
    layer0_outputs(2547) <= a or b;
    layer0_outputs(2548) <= not (a xor b);
    layer0_outputs(2549) <= not (a xor b);
    layer0_outputs(2550) <= not (a or b);
    layer0_outputs(2551) <= not (a xor b);
    layer0_outputs(2552) <= not a or b;
    layer0_outputs(2553) <= a or b;
    layer0_outputs(2554) <= b;
    layer0_outputs(2555) <= not b;
    layer0_outputs(2556) <= b and not a;
    layer0_outputs(2557) <= not b or a;
    layer0_outputs(2558) <= not (a or b);
    layer0_outputs(2559) <= 1'b1;
    layer1_outputs(0) <= a;
    layer1_outputs(1) <= not (a and b);
    layer1_outputs(2) <= a and b;
    layer1_outputs(3) <= b and not a;
    layer1_outputs(4) <= a or b;
    layer1_outputs(5) <= not a;
    layer1_outputs(6) <= not b;
    layer1_outputs(7) <= a and not b;
    layer1_outputs(8) <= not (a xor b);
    layer1_outputs(9) <= a and b;
    layer1_outputs(10) <= not (a and b);
    layer1_outputs(11) <= not (a or b);
    layer1_outputs(12) <= a;
    layer1_outputs(13) <= not b;
    layer1_outputs(14) <= a;
    layer1_outputs(15) <= not (a and b);
    layer1_outputs(16) <= not (a or b);
    layer1_outputs(17) <= not (a and b);
    layer1_outputs(18) <= a and b;
    layer1_outputs(19) <= not b;
    layer1_outputs(20) <= a or b;
    layer1_outputs(21) <= not (a and b);
    layer1_outputs(22) <= b and not a;
    layer1_outputs(23) <= not a;
    layer1_outputs(24) <= a and not b;
    layer1_outputs(25) <= not a or b;
    layer1_outputs(26) <= not b;
    layer1_outputs(27) <= a;
    layer1_outputs(28) <= b and not a;
    layer1_outputs(29) <= not (a or b);
    layer1_outputs(30) <= not a;
    layer1_outputs(31) <= a;
    layer1_outputs(32) <= a and b;
    layer1_outputs(33) <= b;
    layer1_outputs(34) <= not b;
    layer1_outputs(35) <= not (a and b);
    layer1_outputs(36) <= a and b;
    layer1_outputs(37) <= not (a and b);
    layer1_outputs(38) <= a and not b;
    layer1_outputs(39) <= a xor b;
    layer1_outputs(40) <= not (a and b);
    layer1_outputs(41) <= b and not a;
    layer1_outputs(42) <= a and b;
    layer1_outputs(43) <= b;
    layer1_outputs(44) <= b;
    layer1_outputs(45) <= not (a xor b);
    layer1_outputs(46) <= a or b;
    layer1_outputs(47) <= not a or b;
    layer1_outputs(48) <= a xor b;
    layer1_outputs(49) <= a;
    layer1_outputs(50) <= a and b;
    layer1_outputs(51) <= b;
    layer1_outputs(52) <= a and not b;
    layer1_outputs(53) <= b and not a;
    layer1_outputs(54) <= not b or a;
    layer1_outputs(55) <= a;
    layer1_outputs(56) <= a;
    layer1_outputs(57) <= a;
    layer1_outputs(58) <= a and not b;
    layer1_outputs(59) <= not a;
    layer1_outputs(60) <= 1'b1;
    layer1_outputs(61) <= b;
    layer1_outputs(62) <= not (a xor b);
    layer1_outputs(63) <= a;
    layer1_outputs(64) <= a xor b;
    layer1_outputs(65) <= a and b;
    layer1_outputs(66) <= a;
    layer1_outputs(67) <= a and not b;
    layer1_outputs(68) <= a xor b;
    layer1_outputs(69) <= a and not b;
    layer1_outputs(70) <= not (a xor b);
    layer1_outputs(71) <= b and not a;
    layer1_outputs(72) <= a;
    layer1_outputs(73) <= a xor b;
    layer1_outputs(74) <= not a;
    layer1_outputs(75) <= a or b;
    layer1_outputs(76) <= a or b;
    layer1_outputs(77) <= b and not a;
    layer1_outputs(78) <= not a or b;
    layer1_outputs(79) <= not a;
    layer1_outputs(80) <= a xor b;
    layer1_outputs(81) <= not a;
    layer1_outputs(82) <= a and b;
    layer1_outputs(83) <= b;
    layer1_outputs(84) <= a or b;
    layer1_outputs(85) <= a xor b;
    layer1_outputs(86) <= not a;
    layer1_outputs(87) <= b;
    layer1_outputs(88) <= not (a xor b);
    layer1_outputs(89) <= a or b;
    layer1_outputs(90) <= b and not a;
    layer1_outputs(91) <= b and not a;
    layer1_outputs(92) <= 1'b0;
    layer1_outputs(93) <= a or b;
    layer1_outputs(94) <= not (a or b);
    layer1_outputs(95) <= not a or b;
    layer1_outputs(96) <= not b;
    layer1_outputs(97) <= not b;
    layer1_outputs(98) <= not b or a;
    layer1_outputs(99) <= not (a and b);
    layer1_outputs(100) <= not b;
    layer1_outputs(101) <= a and b;
    layer1_outputs(102) <= not b or a;
    layer1_outputs(103) <= not b;
    layer1_outputs(104) <= a and b;
    layer1_outputs(105) <= a and not b;
    layer1_outputs(106) <= a;
    layer1_outputs(107) <= a;
    layer1_outputs(108) <= a or b;
    layer1_outputs(109) <= a or b;
    layer1_outputs(110) <= b and not a;
    layer1_outputs(111) <= not a;
    layer1_outputs(112) <= a or b;
    layer1_outputs(113) <= a and not b;
    layer1_outputs(114) <= not b or a;
    layer1_outputs(115) <= a and not b;
    layer1_outputs(116) <= not (a or b);
    layer1_outputs(117) <= not (a or b);
    layer1_outputs(118) <= b and not a;
    layer1_outputs(119) <= not a or b;
    layer1_outputs(120) <= not a or b;
    layer1_outputs(121) <= a or b;
    layer1_outputs(122) <= not (a or b);
    layer1_outputs(123) <= a xor b;
    layer1_outputs(124) <= a and not b;
    layer1_outputs(125) <= a or b;
    layer1_outputs(126) <= not b;
    layer1_outputs(127) <= not b;
    layer1_outputs(128) <= not b;
    layer1_outputs(129) <= a xor b;
    layer1_outputs(130) <= not (a or b);
    layer1_outputs(131) <= a and not b;
    layer1_outputs(132) <= b;
    layer1_outputs(133) <= not b or a;
    layer1_outputs(134) <= not (a or b);
    layer1_outputs(135) <= a xor b;
    layer1_outputs(136) <= b and not a;
    layer1_outputs(137) <= not a;
    layer1_outputs(138) <= b;
    layer1_outputs(139) <= a and b;
    layer1_outputs(140) <= b;
    layer1_outputs(141) <= not b;
    layer1_outputs(142) <= b;
    layer1_outputs(143) <= a and b;
    layer1_outputs(144) <= a and b;
    layer1_outputs(145) <= a and b;
    layer1_outputs(146) <= a xor b;
    layer1_outputs(147) <= not (a xor b);
    layer1_outputs(148) <= a or b;
    layer1_outputs(149) <= not a;
    layer1_outputs(150) <= a and b;
    layer1_outputs(151) <= not b or a;
    layer1_outputs(152) <= a or b;
    layer1_outputs(153) <= not (a xor b);
    layer1_outputs(154) <= a or b;
    layer1_outputs(155) <= not a or b;
    layer1_outputs(156) <= not a;
    layer1_outputs(157) <= not b;
    layer1_outputs(158) <= a;
    layer1_outputs(159) <= not (a and b);
    layer1_outputs(160) <= b and not a;
    layer1_outputs(161) <= not (a or b);
    layer1_outputs(162) <= not a or b;
    layer1_outputs(163) <= a and not b;
    layer1_outputs(164) <= not b or a;
    layer1_outputs(165) <= not (a or b);
    layer1_outputs(166) <= not (a or b);
    layer1_outputs(167) <= not a;
    layer1_outputs(168) <= 1'b0;
    layer1_outputs(169) <= not b;
    layer1_outputs(170) <= b;
    layer1_outputs(171) <= not (a xor b);
    layer1_outputs(172) <= a and not b;
    layer1_outputs(173) <= a;
    layer1_outputs(174) <= a;
    layer1_outputs(175) <= not (a and b);
    layer1_outputs(176) <= a and not b;
    layer1_outputs(177) <= a or b;
    layer1_outputs(178) <= a xor b;
    layer1_outputs(179) <= not b or a;
    layer1_outputs(180) <= not (a or b);
    layer1_outputs(181) <= a or b;
    layer1_outputs(182) <= not (a xor b);
    layer1_outputs(183) <= not b;
    layer1_outputs(184) <= 1'b1;
    layer1_outputs(185) <= b and not a;
    layer1_outputs(186) <= not (a or b);
    layer1_outputs(187) <= a and b;
    layer1_outputs(188) <= a and b;
    layer1_outputs(189) <= not b;
    layer1_outputs(190) <= a and b;
    layer1_outputs(191) <= a;
    layer1_outputs(192) <= not b;
    layer1_outputs(193) <= 1'b1;
    layer1_outputs(194) <= 1'b0;
    layer1_outputs(195) <= a xor b;
    layer1_outputs(196) <= not a or b;
    layer1_outputs(197) <= a;
    layer1_outputs(198) <= not (a xor b);
    layer1_outputs(199) <= not (a xor b);
    layer1_outputs(200) <= 1'b1;
    layer1_outputs(201) <= a;
    layer1_outputs(202) <= not a;
    layer1_outputs(203) <= a;
    layer1_outputs(204) <= not (a and b);
    layer1_outputs(205) <= not (a or b);
    layer1_outputs(206) <= not a;
    layer1_outputs(207) <= a and b;
    layer1_outputs(208) <= a xor b;
    layer1_outputs(209) <= b;
    layer1_outputs(210) <= b and not a;
    layer1_outputs(211) <= not (a xor b);
    layer1_outputs(212) <= a;
    layer1_outputs(213) <= not a or b;
    layer1_outputs(214) <= a;
    layer1_outputs(215) <= b and not a;
    layer1_outputs(216) <= not b;
    layer1_outputs(217) <= not b or a;
    layer1_outputs(218) <= not a;
    layer1_outputs(219) <= a and not b;
    layer1_outputs(220) <= not b or a;
    layer1_outputs(221) <= b and not a;
    layer1_outputs(222) <= 1'b0;
    layer1_outputs(223) <= a or b;
    layer1_outputs(224) <= not b or a;
    layer1_outputs(225) <= not a;
    layer1_outputs(226) <= not (a or b);
    layer1_outputs(227) <= not (a and b);
    layer1_outputs(228) <= a;
    layer1_outputs(229) <= not a;
    layer1_outputs(230) <= a or b;
    layer1_outputs(231) <= not b or a;
    layer1_outputs(232) <= not a;
    layer1_outputs(233) <= not a;
    layer1_outputs(234) <= not (a or b);
    layer1_outputs(235) <= not a;
    layer1_outputs(236) <= not b or a;
    layer1_outputs(237) <= 1'b1;
    layer1_outputs(238) <= b and not a;
    layer1_outputs(239) <= a;
    layer1_outputs(240) <= a;
    layer1_outputs(241) <= not b;
    layer1_outputs(242) <= a and not b;
    layer1_outputs(243) <= not b or a;
    layer1_outputs(244) <= a and not b;
    layer1_outputs(245) <= a or b;
    layer1_outputs(246) <= not (a or b);
    layer1_outputs(247) <= not b;
    layer1_outputs(248) <= b;
    layer1_outputs(249) <= not (a xor b);
    layer1_outputs(250) <= not a;
    layer1_outputs(251) <= 1'b1;
    layer1_outputs(252) <= not (a and b);
    layer1_outputs(253) <= 1'b0;
    layer1_outputs(254) <= not (a and b);
    layer1_outputs(255) <= not (a or b);
    layer1_outputs(256) <= a xor b;
    layer1_outputs(257) <= b;
    layer1_outputs(258) <= not (a and b);
    layer1_outputs(259) <= not a;
    layer1_outputs(260) <= not (a and b);
    layer1_outputs(261) <= a;
    layer1_outputs(262) <= not b or a;
    layer1_outputs(263) <= not a;
    layer1_outputs(264) <= not (a or b);
    layer1_outputs(265) <= a xor b;
    layer1_outputs(266) <= a or b;
    layer1_outputs(267) <= b;
    layer1_outputs(268) <= not a or b;
    layer1_outputs(269) <= not a;
    layer1_outputs(270) <= b and not a;
    layer1_outputs(271) <= a;
    layer1_outputs(272) <= not a;
    layer1_outputs(273) <= a or b;
    layer1_outputs(274) <= b;
    layer1_outputs(275) <= 1'b1;
    layer1_outputs(276) <= not (a and b);
    layer1_outputs(277) <= a;
    layer1_outputs(278) <= not (a or b);
    layer1_outputs(279) <= a and b;
    layer1_outputs(280) <= 1'b1;
    layer1_outputs(281) <= not b or a;
    layer1_outputs(282) <= a and b;
    layer1_outputs(283) <= not (a and b);
    layer1_outputs(284) <= a or b;
    layer1_outputs(285) <= 1'b0;
    layer1_outputs(286) <= a or b;
    layer1_outputs(287) <= not a;
    layer1_outputs(288) <= a;
    layer1_outputs(289) <= not a;
    layer1_outputs(290) <= b and not a;
    layer1_outputs(291) <= a and b;
    layer1_outputs(292) <= not (a xor b);
    layer1_outputs(293) <= b;
    layer1_outputs(294) <= a or b;
    layer1_outputs(295) <= b;
    layer1_outputs(296) <= not (a or b);
    layer1_outputs(297) <= not (a xor b);
    layer1_outputs(298) <= not b;
    layer1_outputs(299) <= not (a or b);
    layer1_outputs(300) <= not (a or b);
    layer1_outputs(301) <= not a or b;
    layer1_outputs(302) <= not a or b;
    layer1_outputs(303) <= not a or b;
    layer1_outputs(304) <= not b or a;
    layer1_outputs(305) <= not b;
    layer1_outputs(306) <= a and not b;
    layer1_outputs(307) <= b;
    layer1_outputs(308) <= not (a or b);
    layer1_outputs(309) <= not b or a;
    layer1_outputs(310) <= a;
    layer1_outputs(311) <= b;
    layer1_outputs(312) <= not b;
    layer1_outputs(313) <= not (a or b);
    layer1_outputs(314) <= a;
    layer1_outputs(315) <= not (a and b);
    layer1_outputs(316) <= a xor b;
    layer1_outputs(317) <= not (a and b);
    layer1_outputs(318) <= not b or a;
    layer1_outputs(319) <= a xor b;
    layer1_outputs(320) <= not a;
    layer1_outputs(321) <= not b or a;
    layer1_outputs(322) <= 1'b1;
    layer1_outputs(323) <= b;
    layer1_outputs(324) <= not a or b;
    layer1_outputs(325) <= not (a and b);
    layer1_outputs(326) <= a and not b;
    layer1_outputs(327) <= 1'b0;
    layer1_outputs(328) <= b;
    layer1_outputs(329) <= not b;
    layer1_outputs(330) <= a xor b;
    layer1_outputs(331) <= b and not a;
    layer1_outputs(332) <= a and not b;
    layer1_outputs(333) <= a and b;
    layer1_outputs(334) <= not (a or b);
    layer1_outputs(335) <= not (a or b);
    layer1_outputs(336) <= not a;
    layer1_outputs(337) <= not a or b;
    layer1_outputs(338) <= not b or a;
    layer1_outputs(339) <= not (a or b);
    layer1_outputs(340) <= not b;
    layer1_outputs(341) <= 1'b1;
    layer1_outputs(342) <= a or b;
    layer1_outputs(343) <= not (a or b);
    layer1_outputs(344) <= b and not a;
    layer1_outputs(345) <= b and not a;
    layer1_outputs(346) <= not (a and b);
    layer1_outputs(347) <= not a;
    layer1_outputs(348) <= not (a or b);
    layer1_outputs(349) <= a;
    layer1_outputs(350) <= not a;
    layer1_outputs(351) <= a;
    layer1_outputs(352) <= not a;
    layer1_outputs(353) <= b;
    layer1_outputs(354) <= not (a xor b);
    layer1_outputs(355) <= a or b;
    layer1_outputs(356) <= a and not b;
    layer1_outputs(357) <= not b or a;
    layer1_outputs(358) <= not a;
    layer1_outputs(359) <= not (a or b);
    layer1_outputs(360) <= not (a and b);
    layer1_outputs(361) <= not b;
    layer1_outputs(362) <= not b or a;
    layer1_outputs(363) <= b;
    layer1_outputs(364) <= not (a xor b);
    layer1_outputs(365) <= a and b;
    layer1_outputs(366) <= not (a and b);
    layer1_outputs(367) <= not (a or b);
    layer1_outputs(368) <= b;
    layer1_outputs(369) <= a and not b;
    layer1_outputs(370) <= not b or a;
    layer1_outputs(371) <= not a or b;
    layer1_outputs(372) <= not a;
    layer1_outputs(373) <= not b;
    layer1_outputs(374) <= a;
    layer1_outputs(375) <= not (a xor b);
    layer1_outputs(376) <= a or b;
    layer1_outputs(377) <= not b or a;
    layer1_outputs(378) <= not b;
    layer1_outputs(379) <= a or b;
    layer1_outputs(380) <= a or b;
    layer1_outputs(381) <= not b;
    layer1_outputs(382) <= b;
    layer1_outputs(383) <= not (a and b);
    layer1_outputs(384) <= not a;
    layer1_outputs(385) <= a and b;
    layer1_outputs(386) <= not (a or b);
    layer1_outputs(387) <= not (a or b);
    layer1_outputs(388) <= not b;
    layer1_outputs(389) <= not a;
    layer1_outputs(390) <= a and not b;
    layer1_outputs(391) <= not a;
    layer1_outputs(392) <= not a or b;
    layer1_outputs(393) <= a xor b;
    layer1_outputs(394) <= not (a or b);
    layer1_outputs(395) <= 1'b0;
    layer1_outputs(396) <= b;
    layer1_outputs(397) <= a and b;
    layer1_outputs(398) <= a or b;
    layer1_outputs(399) <= not (a and b);
    layer1_outputs(400) <= not b;
    layer1_outputs(401) <= b and not a;
    layer1_outputs(402) <= not b;
    layer1_outputs(403) <= not a or b;
    layer1_outputs(404) <= b and not a;
    layer1_outputs(405) <= not b;
    layer1_outputs(406) <= b;
    layer1_outputs(407) <= not b or a;
    layer1_outputs(408) <= not b;
    layer1_outputs(409) <= b and not a;
    layer1_outputs(410) <= not (a or b);
    layer1_outputs(411) <= b and not a;
    layer1_outputs(412) <= a and not b;
    layer1_outputs(413) <= not b;
    layer1_outputs(414) <= a xor b;
    layer1_outputs(415) <= not (a and b);
    layer1_outputs(416) <= not a or b;
    layer1_outputs(417) <= a or b;
    layer1_outputs(418) <= not b or a;
    layer1_outputs(419) <= not b or a;
    layer1_outputs(420) <= b;
    layer1_outputs(421) <= b;
    layer1_outputs(422) <= b;
    layer1_outputs(423) <= a and not b;
    layer1_outputs(424) <= not a or b;
    layer1_outputs(425) <= not (a xor b);
    layer1_outputs(426) <= a or b;
    layer1_outputs(427) <= a and b;
    layer1_outputs(428) <= a;
    layer1_outputs(429) <= b;
    layer1_outputs(430) <= not b or a;
    layer1_outputs(431) <= not a;
    layer1_outputs(432) <= not a or b;
    layer1_outputs(433) <= not a or b;
    layer1_outputs(434) <= a or b;
    layer1_outputs(435) <= not a;
    layer1_outputs(436) <= a and not b;
    layer1_outputs(437) <= b and not a;
    layer1_outputs(438) <= not (a or b);
    layer1_outputs(439) <= not a or b;
    layer1_outputs(440) <= a or b;
    layer1_outputs(441) <= a;
    layer1_outputs(442) <= a;
    layer1_outputs(443) <= not a or b;
    layer1_outputs(444) <= not a;
    layer1_outputs(445) <= b and not a;
    layer1_outputs(446) <= not a;
    layer1_outputs(447) <= a and not b;
    layer1_outputs(448) <= b;
    layer1_outputs(449) <= a and not b;
    layer1_outputs(450) <= b;
    layer1_outputs(451) <= a or b;
    layer1_outputs(452) <= a or b;
    layer1_outputs(453) <= a;
    layer1_outputs(454) <= b;
    layer1_outputs(455) <= not (a xor b);
    layer1_outputs(456) <= 1'b1;
    layer1_outputs(457) <= not b or a;
    layer1_outputs(458) <= b and not a;
    layer1_outputs(459) <= b;
    layer1_outputs(460) <= not (a xor b);
    layer1_outputs(461) <= a or b;
    layer1_outputs(462) <= not a or b;
    layer1_outputs(463) <= not (a or b);
    layer1_outputs(464) <= a and not b;
    layer1_outputs(465) <= not a;
    layer1_outputs(466) <= not a or b;
    layer1_outputs(467) <= a and b;
    layer1_outputs(468) <= not (a xor b);
    layer1_outputs(469) <= not a or b;
    layer1_outputs(470) <= 1'b0;
    layer1_outputs(471) <= not (a xor b);
    layer1_outputs(472) <= not b;
    layer1_outputs(473) <= a and b;
    layer1_outputs(474) <= not (a xor b);
    layer1_outputs(475) <= not a or b;
    layer1_outputs(476) <= not (a xor b);
    layer1_outputs(477) <= not b;
    layer1_outputs(478) <= not (a xor b);
    layer1_outputs(479) <= not (a and b);
    layer1_outputs(480) <= a;
    layer1_outputs(481) <= a and not b;
    layer1_outputs(482) <= not a or b;
    layer1_outputs(483) <= not (a xor b);
    layer1_outputs(484) <= a or b;
    layer1_outputs(485) <= a;
    layer1_outputs(486) <= not (a or b);
    layer1_outputs(487) <= a;
    layer1_outputs(488) <= a and b;
    layer1_outputs(489) <= a;
    layer1_outputs(490) <= b;
    layer1_outputs(491) <= not b or a;
    layer1_outputs(492) <= a;
    layer1_outputs(493) <= not (a or b);
    layer1_outputs(494) <= b;
    layer1_outputs(495) <= not b;
    layer1_outputs(496) <= b;
    layer1_outputs(497) <= a and b;
    layer1_outputs(498) <= b;
    layer1_outputs(499) <= not (a or b);
    layer1_outputs(500) <= not a or b;
    layer1_outputs(501) <= a and not b;
    layer1_outputs(502) <= a and not b;
    layer1_outputs(503) <= not a;
    layer1_outputs(504) <= a or b;
    layer1_outputs(505) <= a and not b;
    layer1_outputs(506) <= a xor b;
    layer1_outputs(507) <= a and b;
    layer1_outputs(508) <= b;
    layer1_outputs(509) <= not (a and b);
    layer1_outputs(510) <= a and not b;
    layer1_outputs(511) <= b;
    layer1_outputs(512) <= b and not a;
    layer1_outputs(513) <= a;
    layer1_outputs(514) <= b and not a;
    layer1_outputs(515) <= 1'b1;
    layer1_outputs(516) <= a xor b;
    layer1_outputs(517) <= b;
    layer1_outputs(518) <= b and not a;
    layer1_outputs(519) <= not b or a;
    layer1_outputs(520) <= a xor b;
    layer1_outputs(521) <= not (a and b);
    layer1_outputs(522) <= not (a and b);
    layer1_outputs(523) <= not (a and b);
    layer1_outputs(524) <= a or b;
    layer1_outputs(525) <= a;
    layer1_outputs(526) <= not b or a;
    layer1_outputs(527) <= b and not a;
    layer1_outputs(528) <= not a;
    layer1_outputs(529) <= a;
    layer1_outputs(530) <= not a;
    layer1_outputs(531) <= b;
    layer1_outputs(532) <= not a;
    layer1_outputs(533) <= a xor b;
    layer1_outputs(534) <= not (a or b);
    layer1_outputs(535) <= not (a and b);
    layer1_outputs(536) <= not a;
    layer1_outputs(537) <= b and not a;
    layer1_outputs(538) <= not a;
    layer1_outputs(539) <= not a or b;
    layer1_outputs(540) <= b and not a;
    layer1_outputs(541) <= not b;
    layer1_outputs(542) <= not b or a;
    layer1_outputs(543) <= not a;
    layer1_outputs(544) <= b and not a;
    layer1_outputs(545) <= a and not b;
    layer1_outputs(546) <= not (a xor b);
    layer1_outputs(547) <= not a or b;
    layer1_outputs(548) <= a;
    layer1_outputs(549) <= b and not a;
    layer1_outputs(550) <= not b;
    layer1_outputs(551) <= b;
    layer1_outputs(552) <= not (a and b);
    layer1_outputs(553) <= a xor b;
    layer1_outputs(554) <= a or b;
    layer1_outputs(555) <= not b;
    layer1_outputs(556) <= not a or b;
    layer1_outputs(557) <= b and not a;
    layer1_outputs(558) <= a;
    layer1_outputs(559) <= b;
    layer1_outputs(560) <= a and b;
    layer1_outputs(561) <= b and not a;
    layer1_outputs(562) <= a and not b;
    layer1_outputs(563) <= not (a and b);
    layer1_outputs(564) <= not b;
    layer1_outputs(565) <= b;
    layer1_outputs(566) <= b and not a;
    layer1_outputs(567) <= not a;
    layer1_outputs(568) <= not a or b;
    layer1_outputs(569) <= a xor b;
    layer1_outputs(570) <= 1'b0;
    layer1_outputs(571) <= a and b;
    layer1_outputs(572) <= a or b;
    layer1_outputs(573) <= b and not a;
    layer1_outputs(574) <= not (a and b);
    layer1_outputs(575) <= not (a and b);
    layer1_outputs(576) <= a and b;
    layer1_outputs(577) <= a;
    layer1_outputs(578) <= a and not b;
    layer1_outputs(579) <= b;
    layer1_outputs(580) <= not b or a;
    layer1_outputs(581) <= a or b;
    layer1_outputs(582) <= not a;
    layer1_outputs(583) <= not b or a;
    layer1_outputs(584) <= not b or a;
    layer1_outputs(585) <= b;
    layer1_outputs(586) <= a and b;
    layer1_outputs(587) <= not a or b;
    layer1_outputs(588) <= not (a xor b);
    layer1_outputs(589) <= a or b;
    layer1_outputs(590) <= a;
    layer1_outputs(591) <= b;
    layer1_outputs(592) <= not b or a;
    layer1_outputs(593) <= not (a or b);
    layer1_outputs(594) <= not b;
    layer1_outputs(595) <= a or b;
    layer1_outputs(596) <= a and b;
    layer1_outputs(597) <= not (a or b);
    layer1_outputs(598) <= not (a or b);
    layer1_outputs(599) <= a or b;
    layer1_outputs(600) <= not a;
    layer1_outputs(601) <= 1'b1;
    layer1_outputs(602) <= not (a or b);
    layer1_outputs(603) <= not a;
    layer1_outputs(604) <= a or b;
    layer1_outputs(605) <= a and not b;
    layer1_outputs(606) <= not (a or b);
    layer1_outputs(607) <= a;
    layer1_outputs(608) <= b;
    layer1_outputs(609) <= not a or b;
    layer1_outputs(610) <= a;
    layer1_outputs(611) <= a;
    layer1_outputs(612) <= not a;
    layer1_outputs(613) <= not a or b;
    layer1_outputs(614) <= a xor b;
    layer1_outputs(615) <= not (a and b);
    layer1_outputs(616) <= 1'b0;
    layer1_outputs(617) <= a xor b;
    layer1_outputs(618) <= a and not b;
    layer1_outputs(619) <= not b;
    layer1_outputs(620) <= a and not b;
    layer1_outputs(621) <= not b or a;
    layer1_outputs(622) <= b and not a;
    layer1_outputs(623) <= a or b;
    layer1_outputs(624) <= not b or a;
    layer1_outputs(625) <= b;
    layer1_outputs(626) <= 1'b0;
    layer1_outputs(627) <= a;
    layer1_outputs(628) <= a or b;
    layer1_outputs(629) <= a and b;
    layer1_outputs(630) <= not (a or b);
    layer1_outputs(631) <= a and b;
    layer1_outputs(632) <= not (a xor b);
    layer1_outputs(633) <= a and b;
    layer1_outputs(634) <= b;
    layer1_outputs(635) <= 1'b1;
    layer1_outputs(636) <= not (a xor b);
    layer1_outputs(637) <= a;
    layer1_outputs(638) <= not b;
    layer1_outputs(639) <= not (a xor b);
    layer1_outputs(640) <= b;
    layer1_outputs(641) <= a or b;
    layer1_outputs(642) <= a xor b;
    layer1_outputs(643) <= 1'b1;
    layer1_outputs(644) <= a;
    layer1_outputs(645) <= a;
    layer1_outputs(646) <= not (a or b);
    layer1_outputs(647) <= not (a and b);
    layer1_outputs(648) <= not b or a;
    layer1_outputs(649) <= not (a or b);
    layer1_outputs(650) <= a;
    layer1_outputs(651) <= a;
    layer1_outputs(652) <= not a;
    layer1_outputs(653) <= 1'b1;
    layer1_outputs(654) <= a or b;
    layer1_outputs(655) <= a and b;
    layer1_outputs(656) <= a and not b;
    layer1_outputs(657) <= a xor b;
    layer1_outputs(658) <= a xor b;
    layer1_outputs(659) <= not b or a;
    layer1_outputs(660) <= b;
    layer1_outputs(661) <= a xor b;
    layer1_outputs(662) <= b;
    layer1_outputs(663) <= a or b;
    layer1_outputs(664) <= a and not b;
    layer1_outputs(665) <= not a or b;
    layer1_outputs(666) <= b;
    layer1_outputs(667) <= not a;
    layer1_outputs(668) <= not b;
    layer1_outputs(669) <= not (a or b);
    layer1_outputs(670) <= not b or a;
    layer1_outputs(671) <= not b;
    layer1_outputs(672) <= not (a and b);
    layer1_outputs(673) <= a and b;
    layer1_outputs(674) <= b and not a;
    layer1_outputs(675) <= a or b;
    layer1_outputs(676) <= not (a and b);
    layer1_outputs(677) <= a xor b;
    layer1_outputs(678) <= b and not a;
    layer1_outputs(679) <= not b;
    layer1_outputs(680) <= not b;
    layer1_outputs(681) <= b and not a;
    layer1_outputs(682) <= b;
    layer1_outputs(683) <= a or b;
    layer1_outputs(684) <= 1'b0;
    layer1_outputs(685) <= a or b;
    layer1_outputs(686) <= a;
    layer1_outputs(687) <= not a;
    layer1_outputs(688) <= a and b;
    layer1_outputs(689) <= a xor b;
    layer1_outputs(690) <= a;
    layer1_outputs(691) <= a and b;
    layer1_outputs(692) <= not (a and b);
    layer1_outputs(693) <= not (a or b);
    layer1_outputs(694) <= a or b;
    layer1_outputs(695) <= b;
    layer1_outputs(696) <= b;
    layer1_outputs(697) <= not a or b;
    layer1_outputs(698) <= not (a and b);
    layer1_outputs(699) <= b;
    layer1_outputs(700) <= a xor b;
    layer1_outputs(701) <= b;
    layer1_outputs(702) <= not (a xor b);
    layer1_outputs(703) <= not a;
    layer1_outputs(704) <= not a;
    layer1_outputs(705) <= not (a and b);
    layer1_outputs(706) <= not a;
    layer1_outputs(707) <= not b;
    layer1_outputs(708) <= b;
    layer1_outputs(709) <= a or b;
    layer1_outputs(710) <= b;
    layer1_outputs(711) <= a and not b;
    layer1_outputs(712) <= not b;
    layer1_outputs(713) <= not (a xor b);
    layer1_outputs(714) <= not b or a;
    layer1_outputs(715) <= a xor b;
    layer1_outputs(716) <= b;
    layer1_outputs(717) <= not (a and b);
    layer1_outputs(718) <= not a;
    layer1_outputs(719) <= not (a or b);
    layer1_outputs(720) <= not (a or b);
    layer1_outputs(721) <= not a;
    layer1_outputs(722) <= not (a xor b);
    layer1_outputs(723) <= a and b;
    layer1_outputs(724) <= a;
    layer1_outputs(725) <= not a;
    layer1_outputs(726) <= not b or a;
    layer1_outputs(727) <= b;
    layer1_outputs(728) <= b and not a;
    layer1_outputs(729) <= a and not b;
    layer1_outputs(730) <= 1'b0;
    layer1_outputs(731) <= not a or b;
    layer1_outputs(732) <= a and b;
    layer1_outputs(733) <= 1'b1;
    layer1_outputs(734) <= not b or a;
    layer1_outputs(735) <= not b;
    layer1_outputs(736) <= b;
    layer1_outputs(737) <= a and b;
    layer1_outputs(738) <= not (a or b);
    layer1_outputs(739) <= not (a xor b);
    layer1_outputs(740) <= a or b;
    layer1_outputs(741) <= not b;
    layer1_outputs(742) <= a or b;
    layer1_outputs(743) <= not (a or b);
    layer1_outputs(744) <= b;
    layer1_outputs(745) <= a;
    layer1_outputs(746) <= not b;
    layer1_outputs(747) <= not (a xor b);
    layer1_outputs(748) <= a or b;
    layer1_outputs(749) <= a and b;
    layer1_outputs(750) <= not a or b;
    layer1_outputs(751) <= a or b;
    layer1_outputs(752) <= a;
    layer1_outputs(753) <= not b or a;
    layer1_outputs(754) <= a xor b;
    layer1_outputs(755) <= not a;
    layer1_outputs(756) <= a;
    layer1_outputs(757) <= a;
    layer1_outputs(758) <= a;
    layer1_outputs(759) <= a xor b;
    layer1_outputs(760) <= a;
    layer1_outputs(761) <= b;
    layer1_outputs(762) <= 1'b1;
    layer1_outputs(763) <= not a or b;
    layer1_outputs(764) <= not b;
    layer1_outputs(765) <= a and b;
    layer1_outputs(766) <= not (a or b);
    layer1_outputs(767) <= a and not b;
    layer1_outputs(768) <= b and not a;
    layer1_outputs(769) <= not b;
    layer1_outputs(770) <= not a;
    layer1_outputs(771) <= 1'b1;
    layer1_outputs(772) <= not b or a;
    layer1_outputs(773) <= not a or b;
    layer1_outputs(774) <= a or b;
    layer1_outputs(775) <= not b or a;
    layer1_outputs(776) <= not a or b;
    layer1_outputs(777) <= a or b;
    layer1_outputs(778) <= a or b;
    layer1_outputs(779) <= not b or a;
    layer1_outputs(780) <= b and not a;
    layer1_outputs(781) <= a and b;
    layer1_outputs(782) <= not (a and b);
    layer1_outputs(783) <= a or b;
    layer1_outputs(784) <= b and not a;
    layer1_outputs(785) <= not b or a;
    layer1_outputs(786) <= not b;
    layer1_outputs(787) <= a;
    layer1_outputs(788) <= a and b;
    layer1_outputs(789) <= b;
    layer1_outputs(790) <= b;
    layer1_outputs(791) <= b and not a;
    layer1_outputs(792) <= not a or b;
    layer1_outputs(793) <= b and not a;
    layer1_outputs(794) <= not (a and b);
    layer1_outputs(795) <= a and not b;
    layer1_outputs(796) <= a xor b;
    layer1_outputs(797) <= b;
    layer1_outputs(798) <= not (a and b);
    layer1_outputs(799) <= not b or a;
    layer1_outputs(800) <= a or b;
    layer1_outputs(801) <= not b;
    layer1_outputs(802) <= not b;
    layer1_outputs(803) <= a and b;
    layer1_outputs(804) <= b and not a;
    layer1_outputs(805) <= a;
    layer1_outputs(806) <= not b;
    layer1_outputs(807) <= not b;
    layer1_outputs(808) <= not b;
    layer1_outputs(809) <= not (a or b);
    layer1_outputs(810) <= b;
    layer1_outputs(811) <= a xor b;
    layer1_outputs(812) <= b;
    layer1_outputs(813) <= not b or a;
    layer1_outputs(814) <= a and b;
    layer1_outputs(815) <= a or b;
    layer1_outputs(816) <= b and not a;
    layer1_outputs(817) <= not (a xor b);
    layer1_outputs(818) <= not (a and b);
    layer1_outputs(819) <= a and b;
    layer1_outputs(820) <= not a;
    layer1_outputs(821) <= a;
    layer1_outputs(822) <= not a;
    layer1_outputs(823) <= a and not b;
    layer1_outputs(824) <= b and not a;
    layer1_outputs(825) <= not (a and b);
    layer1_outputs(826) <= not b;
    layer1_outputs(827) <= not (a and b);
    layer1_outputs(828) <= b;
    layer1_outputs(829) <= not b;
    layer1_outputs(830) <= not a or b;
    layer1_outputs(831) <= not (a xor b);
    layer1_outputs(832) <= not (a and b);
    layer1_outputs(833) <= a;
    layer1_outputs(834) <= not a;
    layer1_outputs(835) <= b;
    layer1_outputs(836) <= not a or b;
    layer1_outputs(837) <= a;
    layer1_outputs(838) <= not b;
    layer1_outputs(839) <= a;
    layer1_outputs(840) <= not b;
    layer1_outputs(841) <= not b;
    layer1_outputs(842) <= a and b;
    layer1_outputs(843) <= not b or a;
    layer1_outputs(844) <= a;
    layer1_outputs(845) <= a and b;
    layer1_outputs(846) <= not b;
    layer1_outputs(847) <= not b;
    layer1_outputs(848) <= not a or b;
    layer1_outputs(849) <= not b;
    layer1_outputs(850) <= a or b;
    layer1_outputs(851) <= a or b;
    layer1_outputs(852) <= a;
    layer1_outputs(853) <= not b or a;
    layer1_outputs(854) <= a;
    layer1_outputs(855) <= b;
    layer1_outputs(856) <= a and b;
    layer1_outputs(857) <= not a or b;
    layer1_outputs(858) <= not a;
    layer1_outputs(859) <= not b or a;
    layer1_outputs(860) <= a and not b;
    layer1_outputs(861) <= not (a and b);
    layer1_outputs(862) <= not (a or b);
    layer1_outputs(863) <= not a or b;
    layer1_outputs(864) <= b;
    layer1_outputs(865) <= a;
    layer1_outputs(866) <= not a or b;
    layer1_outputs(867) <= not (a or b);
    layer1_outputs(868) <= not a;
    layer1_outputs(869) <= b and not a;
    layer1_outputs(870) <= not (a or b);
    layer1_outputs(871) <= not (a xor b);
    layer1_outputs(872) <= not b;
    layer1_outputs(873) <= b and not a;
    layer1_outputs(874) <= not a;
    layer1_outputs(875) <= b;
    layer1_outputs(876) <= not b;
    layer1_outputs(877) <= b;
    layer1_outputs(878) <= not b or a;
    layer1_outputs(879) <= b;
    layer1_outputs(880) <= a;
    layer1_outputs(881) <= a or b;
    layer1_outputs(882) <= a and b;
    layer1_outputs(883) <= not (a and b);
    layer1_outputs(884) <= b;
    layer1_outputs(885) <= b;
    layer1_outputs(886) <= not (a or b);
    layer1_outputs(887) <= 1'b0;
    layer1_outputs(888) <= a or b;
    layer1_outputs(889) <= a;
    layer1_outputs(890) <= not (a or b);
    layer1_outputs(891) <= not (a or b);
    layer1_outputs(892) <= a;
    layer1_outputs(893) <= not b;
    layer1_outputs(894) <= a or b;
    layer1_outputs(895) <= not (a xor b);
    layer1_outputs(896) <= not b;
    layer1_outputs(897) <= a and b;
    layer1_outputs(898) <= a;
    layer1_outputs(899) <= not b or a;
    layer1_outputs(900) <= not (a or b);
    layer1_outputs(901) <= not b;
    layer1_outputs(902) <= b;
    layer1_outputs(903) <= a and b;
    layer1_outputs(904) <= not a or b;
    layer1_outputs(905) <= not a or b;
    layer1_outputs(906) <= not b;
    layer1_outputs(907) <= not a or b;
    layer1_outputs(908) <= a;
    layer1_outputs(909) <= a or b;
    layer1_outputs(910) <= not b or a;
    layer1_outputs(911) <= not b or a;
    layer1_outputs(912) <= a and not b;
    layer1_outputs(913) <= not b;
    layer1_outputs(914) <= a and b;
    layer1_outputs(915) <= not (a and b);
    layer1_outputs(916) <= b;
    layer1_outputs(917) <= a and b;
    layer1_outputs(918) <= a or b;
    layer1_outputs(919) <= not b or a;
    layer1_outputs(920) <= a or b;
    layer1_outputs(921) <= not (a and b);
    layer1_outputs(922) <= b and not a;
    layer1_outputs(923) <= a or b;
    layer1_outputs(924) <= not b or a;
    layer1_outputs(925) <= b and not a;
    layer1_outputs(926) <= a;
    layer1_outputs(927) <= a;
    layer1_outputs(928) <= b;
    layer1_outputs(929) <= a and b;
    layer1_outputs(930) <= 1'b0;
    layer1_outputs(931) <= not b or a;
    layer1_outputs(932) <= not (a xor b);
    layer1_outputs(933) <= not b;
    layer1_outputs(934) <= b;
    layer1_outputs(935) <= b;
    layer1_outputs(936) <= not (a and b);
    layer1_outputs(937) <= not b or a;
    layer1_outputs(938) <= a;
    layer1_outputs(939) <= a;
    layer1_outputs(940) <= not (a xor b);
    layer1_outputs(941) <= not a;
    layer1_outputs(942) <= not (a or b);
    layer1_outputs(943) <= not (a and b);
    layer1_outputs(944) <= 1'b1;
    layer1_outputs(945) <= b and not a;
    layer1_outputs(946) <= 1'b1;
    layer1_outputs(947) <= b;
    layer1_outputs(948) <= not a or b;
    layer1_outputs(949) <= a or b;
    layer1_outputs(950) <= a or b;
    layer1_outputs(951) <= not (a xor b);
    layer1_outputs(952) <= not a;
    layer1_outputs(953) <= not a;
    layer1_outputs(954) <= a or b;
    layer1_outputs(955) <= not a or b;
    layer1_outputs(956) <= not b or a;
    layer1_outputs(957) <= not b;
    layer1_outputs(958) <= not a;
    layer1_outputs(959) <= not b;
    layer1_outputs(960) <= not (a and b);
    layer1_outputs(961) <= a and b;
    layer1_outputs(962) <= a;
    layer1_outputs(963) <= 1'b1;
    layer1_outputs(964) <= not b;
    layer1_outputs(965) <= not a;
    layer1_outputs(966) <= not b;
    layer1_outputs(967) <= b;
    layer1_outputs(968) <= not b;
    layer1_outputs(969) <= a;
    layer1_outputs(970) <= not a;
    layer1_outputs(971) <= not (a xor b);
    layer1_outputs(972) <= not b;
    layer1_outputs(973) <= a and b;
    layer1_outputs(974) <= not (a xor b);
    layer1_outputs(975) <= a;
    layer1_outputs(976) <= a or b;
    layer1_outputs(977) <= b and not a;
    layer1_outputs(978) <= a and not b;
    layer1_outputs(979) <= a xor b;
    layer1_outputs(980) <= a and not b;
    layer1_outputs(981) <= b and not a;
    layer1_outputs(982) <= not b;
    layer1_outputs(983) <= b;
    layer1_outputs(984) <= a and not b;
    layer1_outputs(985) <= not (a and b);
    layer1_outputs(986) <= not b;
    layer1_outputs(987) <= a;
    layer1_outputs(988) <= not b;
    layer1_outputs(989) <= not (a xor b);
    layer1_outputs(990) <= not (a or b);
    layer1_outputs(991) <= not b or a;
    layer1_outputs(992) <= not (a xor b);
    layer1_outputs(993) <= not a or b;
    layer1_outputs(994) <= not (a and b);
    layer1_outputs(995) <= not (a xor b);
    layer1_outputs(996) <= a and b;
    layer1_outputs(997) <= a xor b;
    layer1_outputs(998) <= not (a or b);
    layer1_outputs(999) <= not a or b;
    layer1_outputs(1000) <= a or b;
    layer1_outputs(1001) <= not a;
    layer1_outputs(1002) <= b;
    layer1_outputs(1003) <= not b;
    layer1_outputs(1004) <= b and not a;
    layer1_outputs(1005) <= not a or b;
    layer1_outputs(1006) <= not a;
    layer1_outputs(1007) <= a;
    layer1_outputs(1008) <= b;
    layer1_outputs(1009) <= not (a xor b);
    layer1_outputs(1010) <= b and not a;
    layer1_outputs(1011) <= a;
    layer1_outputs(1012) <= b;
    layer1_outputs(1013) <= not (a xor b);
    layer1_outputs(1014) <= not (a xor b);
    layer1_outputs(1015) <= a and b;
    layer1_outputs(1016) <= a or b;
    layer1_outputs(1017) <= not a or b;
    layer1_outputs(1018) <= a;
    layer1_outputs(1019) <= not a or b;
    layer1_outputs(1020) <= not (a or b);
    layer1_outputs(1021) <= b;
    layer1_outputs(1022) <= not a;
    layer1_outputs(1023) <= a;
    layer1_outputs(1024) <= b and not a;
    layer1_outputs(1025) <= not b;
    layer1_outputs(1026) <= a and b;
    layer1_outputs(1027) <= not (a and b);
    layer1_outputs(1028) <= not (a xor b);
    layer1_outputs(1029) <= not b or a;
    layer1_outputs(1030) <= not (a and b);
    layer1_outputs(1031) <= a;
    layer1_outputs(1032) <= b;
    layer1_outputs(1033) <= a and not b;
    layer1_outputs(1034) <= not (a or b);
    layer1_outputs(1035) <= 1'b1;
    layer1_outputs(1036) <= a;
    layer1_outputs(1037) <= b and not a;
    layer1_outputs(1038) <= b and not a;
    layer1_outputs(1039) <= not a;
    layer1_outputs(1040) <= b;
    layer1_outputs(1041) <= b;
    layer1_outputs(1042) <= b;
    layer1_outputs(1043) <= not b or a;
    layer1_outputs(1044) <= 1'b0;
    layer1_outputs(1045) <= not a or b;
    layer1_outputs(1046) <= b;
    layer1_outputs(1047) <= 1'b1;
    layer1_outputs(1048) <= a xor b;
    layer1_outputs(1049) <= a or b;
    layer1_outputs(1050) <= not b or a;
    layer1_outputs(1051) <= not (a or b);
    layer1_outputs(1052) <= a xor b;
    layer1_outputs(1053) <= a;
    layer1_outputs(1054) <= not a;
    layer1_outputs(1055) <= b;
    layer1_outputs(1056) <= not (a and b);
    layer1_outputs(1057) <= not a;
    layer1_outputs(1058) <= not b or a;
    layer1_outputs(1059) <= b;
    layer1_outputs(1060) <= a and b;
    layer1_outputs(1061) <= b and not a;
    layer1_outputs(1062) <= not a;
    layer1_outputs(1063) <= b and not a;
    layer1_outputs(1064) <= a and not b;
    layer1_outputs(1065) <= not b or a;
    layer1_outputs(1066) <= 1'b0;
    layer1_outputs(1067) <= a xor b;
    layer1_outputs(1068) <= a xor b;
    layer1_outputs(1069) <= not (a or b);
    layer1_outputs(1070) <= not a or b;
    layer1_outputs(1071) <= not (a xor b);
    layer1_outputs(1072) <= not (a and b);
    layer1_outputs(1073) <= a;
    layer1_outputs(1074) <= a or b;
    layer1_outputs(1075) <= a or b;
    layer1_outputs(1076) <= not (a and b);
    layer1_outputs(1077) <= 1'b0;
    layer1_outputs(1078) <= not a or b;
    layer1_outputs(1079) <= not b or a;
    layer1_outputs(1080) <= not a or b;
    layer1_outputs(1081) <= not (a and b);
    layer1_outputs(1082) <= not (a or b);
    layer1_outputs(1083) <= not a or b;
    layer1_outputs(1084) <= a xor b;
    layer1_outputs(1085) <= b;
    layer1_outputs(1086) <= a or b;
    layer1_outputs(1087) <= a and b;
    layer1_outputs(1088) <= a xor b;
    layer1_outputs(1089) <= a;
    layer1_outputs(1090) <= a;
    layer1_outputs(1091) <= b;
    layer1_outputs(1092) <= not b;
    layer1_outputs(1093) <= a and not b;
    layer1_outputs(1094) <= not a;
    layer1_outputs(1095) <= not (a xor b);
    layer1_outputs(1096) <= a and not b;
    layer1_outputs(1097) <= not a or b;
    layer1_outputs(1098) <= not b;
    layer1_outputs(1099) <= a and b;
    layer1_outputs(1100) <= a;
    layer1_outputs(1101) <= a and not b;
    layer1_outputs(1102) <= not (a and b);
    layer1_outputs(1103) <= 1'b0;
    layer1_outputs(1104) <= a;
    layer1_outputs(1105) <= not (a and b);
    layer1_outputs(1106) <= not (a and b);
    layer1_outputs(1107) <= not b;
    layer1_outputs(1108) <= a;
    layer1_outputs(1109) <= not a or b;
    layer1_outputs(1110) <= a and not b;
    layer1_outputs(1111) <= not a or b;
    layer1_outputs(1112) <= not a or b;
    layer1_outputs(1113) <= not b;
    layer1_outputs(1114) <= a and not b;
    layer1_outputs(1115) <= not a or b;
    layer1_outputs(1116) <= a and not b;
    layer1_outputs(1117) <= not a or b;
    layer1_outputs(1118) <= not (a xor b);
    layer1_outputs(1119) <= b and not a;
    layer1_outputs(1120) <= a;
    layer1_outputs(1121) <= 1'b1;
    layer1_outputs(1122) <= not a or b;
    layer1_outputs(1123) <= not (a or b);
    layer1_outputs(1124) <= a and b;
    layer1_outputs(1125) <= not (a and b);
    layer1_outputs(1126) <= a xor b;
    layer1_outputs(1127) <= not (a xor b);
    layer1_outputs(1128) <= a;
    layer1_outputs(1129) <= not (a xor b);
    layer1_outputs(1130) <= a and b;
    layer1_outputs(1131) <= b;
    layer1_outputs(1132) <= not b;
    layer1_outputs(1133) <= not b;
    layer1_outputs(1134) <= b;
    layer1_outputs(1135) <= a and not b;
    layer1_outputs(1136) <= not a;
    layer1_outputs(1137) <= a and b;
    layer1_outputs(1138) <= a and b;
    layer1_outputs(1139) <= 1'b1;
    layer1_outputs(1140) <= a;
    layer1_outputs(1141) <= not a or b;
    layer1_outputs(1142) <= b;
    layer1_outputs(1143) <= b;
    layer1_outputs(1144) <= b and not a;
    layer1_outputs(1145) <= not (a or b);
    layer1_outputs(1146) <= a;
    layer1_outputs(1147) <= a or b;
    layer1_outputs(1148) <= not (a or b);
    layer1_outputs(1149) <= b and not a;
    layer1_outputs(1150) <= b;
    layer1_outputs(1151) <= not b;
    layer1_outputs(1152) <= b and not a;
    layer1_outputs(1153) <= not b or a;
    layer1_outputs(1154) <= not a or b;
    layer1_outputs(1155) <= not b or a;
    layer1_outputs(1156) <= a or b;
    layer1_outputs(1157) <= not b or a;
    layer1_outputs(1158) <= a;
    layer1_outputs(1159) <= not a;
    layer1_outputs(1160) <= a and not b;
    layer1_outputs(1161) <= a or b;
    layer1_outputs(1162) <= not (a and b);
    layer1_outputs(1163) <= b;
    layer1_outputs(1164) <= not (a or b);
    layer1_outputs(1165) <= a and not b;
    layer1_outputs(1166) <= not a;
    layer1_outputs(1167) <= a and b;
    layer1_outputs(1168) <= not b;
    layer1_outputs(1169) <= not (a or b);
    layer1_outputs(1170) <= a or b;
    layer1_outputs(1171) <= not a or b;
    layer1_outputs(1172) <= a;
    layer1_outputs(1173) <= not (a and b);
    layer1_outputs(1174) <= a;
    layer1_outputs(1175) <= b;
    layer1_outputs(1176) <= a and not b;
    layer1_outputs(1177) <= b;
    layer1_outputs(1178) <= not b;
    layer1_outputs(1179) <= not (a or b);
    layer1_outputs(1180) <= not a or b;
    layer1_outputs(1181) <= not (a xor b);
    layer1_outputs(1182) <= a or b;
    layer1_outputs(1183) <= a and not b;
    layer1_outputs(1184) <= a;
    layer1_outputs(1185) <= not (a xor b);
    layer1_outputs(1186) <= not (a or b);
    layer1_outputs(1187) <= not b or a;
    layer1_outputs(1188) <= not b or a;
    layer1_outputs(1189) <= not a;
    layer1_outputs(1190) <= b;
    layer1_outputs(1191) <= b and not a;
    layer1_outputs(1192) <= not (a or b);
    layer1_outputs(1193) <= not b;
    layer1_outputs(1194) <= not (a xor b);
    layer1_outputs(1195) <= not a;
    layer1_outputs(1196) <= not b;
    layer1_outputs(1197) <= a and not b;
    layer1_outputs(1198) <= b and not a;
    layer1_outputs(1199) <= not a or b;
    layer1_outputs(1200) <= not a;
    layer1_outputs(1201) <= b;
    layer1_outputs(1202) <= a and b;
    layer1_outputs(1203) <= not (a and b);
    layer1_outputs(1204) <= b and not a;
    layer1_outputs(1205) <= a;
    layer1_outputs(1206) <= b and not a;
    layer1_outputs(1207) <= a;
    layer1_outputs(1208) <= 1'b0;
    layer1_outputs(1209) <= a xor b;
    layer1_outputs(1210) <= not a;
    layer1_outputs(1211) <= a and not b;
    layer1_outputs(1212) <= a and not b;
    layer1_outputs(1213) <= not a;
    layer1_outputs(1214) <= a and not b;
    layer1_outputs(1215) <= a or b;
    layer1_outputs(1216) <= not a;
    layer1_outputs(1217) <= 1'b1;
    layer1_outputs(1218) <= b;
    layer1_outputs(1219) <= not a or b;
    layer1_outputs(1220) <= a or b;
    layer1_outputs(1221) <= b;
    layer1_outputs(1222) <= not (a and b);
    layer1_outputs(1223) <= a or b;
    layer1_outputs(1224) <= 1'b1;
    layer1_outputs(1225) <= a and b;
    layer1_outputs(1226) <= not (a and b);
    layer1_outputs(1227) <= a and b;
    layer1_outputs(1228) <= not (a and b);
    layer1_outputs(1229) <= 1'b1;
    layer1_outputs(1230) <= b;
    layer1_outputs(1231) <= 1'b1;
    layer1_outputs(1232) <= not (a and b);
    layer1_outputs(1233) <= not a;
    layer1_outputs(1234) <= a xor b;
    layer1_outputs(1235) <= not (a or b);
    layer1_outputs(1236) <= a or b;
    layer1_outputs(1237) <= b;
    layer1_outputs(1238) <= 1'b0;
    layer1_outputs(1239) <= not b;
    layer1_outputs(1240) <= a and not b;
    layer1_outputs(1241) <= a xor b;
    layer1_outputs(1242) <= not a;
    layer1_outputs(1243) <= a and not b;
    layer1_outputs(1244) <= a and b;
    layer1_outputs(1245) <= not (a xor b);
    layer1_outputs(1246) <= a;
    layer1_outputs(1247) <= not (a or b);
    layer1_outputs(1248) <= a;
    layer1_outputs(1249) <= not a;
    layer1_outputs(1250) <= b;
    layer1_outputs(1251) <= not b or a;
    layer1_outputs(1252) <= b and not a;
    layer1_outputs(1253) <= a and not b;
    layer1_outputs(1254) <= 1'b1;
    layer1_outputs(1255) <= not a;
    layer1_outputs(1256) <= b;
    layer1_outputs(1257) <= a;
    layer1_outputs(1258) <= not (a xor b);
    layer1_outputs(1259) <= b;
    layer1_outputs(1260) <= not a or b;
    layer1_outputs(1261) <= b;
    layer1_outputs(1262) <= b;
    layer1_outputs(1263) <= a or b;
    layer1_outputs(1264) <= b;
    layer1_outputs(1265) <= not (a xor b);
    layer1_outputs(1266) <= a and b;
    layer1_outputs(1267) <= not b;
    layer1_outputs(1268) <= b and not a;
    layer1_outputs(1269) <= not b or a;
    layer1_outputs(1270) <= a;
    layer1_outputs(1271) <= b;
    layer1_outputs(1272) <= a or b;
    layer1_outputs(1273) <= not a or b;
    layer1_outputs(1274) <= a;
    layer1_outputs(1275) <= a or b;
    layer1_outputs(1276) <= a;
    layer1_outputs(1277) <= not (a or b);
    layer1_outputs(1278) <= a and b;
    layer1_outputs(1279) <= 1'b1;
    layer1_outputs(1280) <= a or b;
    layer1_outputs(1281) <= not b;
    layer1_outputs(1282) <= a and not b;
    layer1_outputs(1283) <= not a or b;
    layer1_outputs(1284) <= not a or b;
    layer1_outputs(1285) <= not b;
    layer1_outputs(1286) <= a and not b;
    layer1_outputs(1287) <= a xor b;
    layer1_outputs(1288) <= not (a and b);
    layer1_outputs(1289) <= not b or a;
    layer1_outputs(1290) <= not (a and b);
    layer1_outputs(1291) <= a;
    layer1_outputs(1292) <= b;
    layer1_outputs(1293) <= not b or a;
    layer1_outputs(1294) <= a and b;
    layer1_outputs(1295) <= b and not a;
    layer1_outputs(1296) <= a and not b;
    layer1_outputs(1297) <= 1'b0;
    layer1_outputs(1298) <= not b;
    layer1_outputs(1299) <= not b;
    layer1_outputs(1300) <= not a;
    layer1_outputs(1301) <= 1'b0;
    layer1_outputs(1302) <= a and b;
    layer1_outputs(1303) <= a;
    layer1_outputs(1304) <= 1'b1;
    layer1_outputs(1305) <= not b;
    layer1_outputs(1306) <= not (a xor b);
    layer1_outputs(1307) <= not a or b;
    layer1_outputs(1308) <= 1'b1;
    layer1_outputs(1309) <= b;
    layer1_outputs(1310) <= not (a or b);
    layer1_outputs(1311) <= not (a or b);
    layer1_outputs(1312) <= b and not a;
    layer1_outputs(1313) <= not (a or b);
    layer1_outputs(1314) <= a;
    layer1_outputs(1315) <= a;
    layer1_outputs(1316) <= a and not b;
    layer1_outputs(1317) <= a;
    layer1_outputs(1318) <= not (a or b);
    layer1_outputs(1319) <= not b;
    layer1_outputs(1320) <= not (a xor b);
    layer1_outputs(1321) <= a or b;
    layer1_outputs(1322) <= not b;
    layer1_outputs(1323) <= b and not a;
    layer1_outputs(1324) <= not (a or b);
    layer1_outputs(1325) <= a xor b;
    layer1_outputs(1326) <= not (a xor b);
    layer1_outputs(1327) <= not (a and b);
    layer1_outputs(1328) <= not (a xor b);
    layer1_outputs(1329) <= a or b;
    layer1_outputs(1330) <= not a or b;
    layer1_outputs(1331) <= b and not a;
    layer1_outputs(1332) <= b and not a;
    layer1_outputs(1333) <= a and not b;
    layer1_outputs(1334) <= a and b;
    layer1_outputs(1335) <= not a;
    layer1_outputs(1336) <= not b or a;
    layer1_outputs(1337) <= b;
    layer1_outputs(1338) <= not b or a;
    layer1_outputs(1339) <= not b;
    layer1_outputs(1340) <= not (a or b);
    layer1_outputs(1341) <= not a or b;
    layer1_outputs(1342) <= a and not b;
    layer1_outputs(1343) <= a xor b;
    layer1_outputs(1344) <= not (a and b);
    layer1_outputs(1345) <= b;
    layer1_outputs(1346) <= b;
    layer1_outputs(1347) <= a;
    layer1_outputs(1348) <= not a;
    layer1_outputs(1349) <= a and not b;
    layer1_outputs(1350) <= not a or b;
    layer1_outputs(1351) <= b;
    layer1_outputs(1352) <= b and not a;
    layer1_outputs(1353) <= not a;
    layer1_outputs(1354) <= not (a and b);
    layer1_outputs(1355) <= not (a and b);
    layer1_outputs(1356) <= b;
    layer1_outputs(1357) <= a and b;
    layer1_outputs(1358) <= not (a and b);
    layer1_outputs(1359) <= not (a and b);
    layer1_outputs(1360) <= not a or b;
    layer1_outputs(1361) <= not (a and b);
    layer1_outputs(1362) <= a xor b;
    layer1_outputs(1363) <= not (a and b);
    layer1_outputs(1364) <= not (a and b);
    layer1_outputs(1365) <= a and b;
    layer1_outputs(1366) <= a and b;
    layer1_outputs(1367) <= not a;
    layer1_outputs(1368) <= not b;
    layer1_outputs(1369) <= a xor b;
    layer1_outputs(1370) <= not a or b;
    layer1_outputs(1371) <= not (a or b);
    layer1_outputs(1372) <= a;
    layer1_outputs(1373) <= not b or a;
    layer1_outputs(1374) <= not b;
    layer1_outputs(1375) <= b;
    layer1_outputs(1376) <= not (a or b);
    layer1_outputs(1377) <= not a;
    layer1_outputs(1378) <= not a;
    layer1_outputs(1379) <= not (a and b);
    layer1_outputs(1380) <= not b or a;
    layer1_outputs(1381) <= a;
    layer1_outputs(1382) <= a or b;
    layer1_outputs(1383) <= not b or a;
    layer1_outputs(1384) <= b;
    layer1_outputs(1385) <= 1'b1;
    layer1_outputs(1386) <= a or b;
    layer1_outputs(1387) <= 1'b0;
    layer1_outputs(1388) <= a xor b;
    layer1_outputs(1389) <= b;
    layer1_outputs(1390) <= a and b;
    layer1_outputs(1391) <= a or b;
    layer1_outputs(1392) <= a and b;
    layer1_outputs(1393) <= not (a xor b);
    layer1_outputs(1394) <= not (a or b);
    layer1_outputs(1395) <= not (a and b);
    layer1_outputs(1396) <= not (a and b);
    layer1_outputs(1397) <= not a;
    layer1_outputs(1398) <= a;
    layer1_outputs(1399) <= b;
    layer1_outputs(1400) <= not (a and b);
    layer1_outputs(1401) <= a;
    layer1_outputs(1402) <= a or b;
    layer1_outputs(1403) <= b;
    layer1_outputs(1404) <= a and not b;
    layer1_outputs(1405) <= a and not b;
    layer1_outputs(1406) <= not a or b;
    layer1_outputs(1407) <= b;
    layer1_outputs(1408) <= not (a and b);
    layer1_outputs(1409) <= not (a or b);
    layer1_outputs(1410) <= not (a and b);
    layer1_outputs(1411) <= a and not b;
    layer1_outputs(1412) <= a and b;
    layer1_outputs(1413) <= a;
    layer1_outputs(1414) <= a or b;
    layer1_outputs(1415) <= a and b;
    layer1_outputs(1416) <= a xor b;
    layer1_outputs(1417) <= a or b;
    layer1_outputs(1418) <= not b;
    layer1_outputs(1419) <= a xor b;
    layer1_outputs(1420) <= not b;
    layer1_outputs(1421) <= 1'b0;
    layer1_outputs(1422) <= not b or a;
    layer1_outputs(1423) <= b and not a;
    layer1_outputs(1424) <= not a;
    layer1_outputs(1425) <= a and not b;
    layer1_outputs(1426) <= a;
    layer1_outputs(1427) <= b and not a;
    layer1_outputs(1428) <= a and not b;
    layer1_outputs(1429) <= b and not a;
    layer1_outputs(1430) <= a and not b;
    layer1_outputs(1431) <= b;
    layer1_outputs(1432) <= b;
    layer1_outputs(1433) <= a and b;
    layer1_outputs(1434) <= not (a and b);
    layer1_outputs(1435) <= a xor b;
    layer1_outputs(1436) <= not a or b;
    layer1_outputs(1437) <= b;
    layer1_outputs(1438) <= not b or a;
    layer1_outputs(1439) <= b and not a;
    layer1_outputs(1440) <= 1'b0;
    layer1_outputs(1441) <= not a or b;
    layer1_outputs(1442) <= not a;
    layer1_outputs(1443) <= not a;
    layer1_outputs(1444) <= not (a or b);
    layer1_outputs(1445) <= not b or a;
    layer1_outputs(1446) <= not a;
    layer1_outputs(1447) <= not (a xor b);
    layer1_outputs(1448) <= b;
    layer1_outputs(1449) <= a;
    layer1_outputs(1450) <= a;
    layer1_outputs(1451) <= a or b;
    layer1_outputs(1452) <= not a;
    layer1_outputs(1453) <= a and not b;
    layer1_outputs(1454) <= not (a xor b);
    layer1_outputs(1455) <= not a;
    layer1_outputs(1456) <= not a or b;
    layer1_outputs(1457) <= not (a or b);
    layer1_outputs(1458) <= a xor b;
    layer1_outputs(1459) <= not a;
    layer1_outputs(1460) <= not b;
    layer1_outputs(1461) <= b and not a;
    layer1_outputs(1462) <= a or b;
    layer1_outputs(1463) <= a;
    layer1_outputs(1464) <= a and not b;
    layer1_outputs(1465) <= not a or b;
    layer1_outputs(1466) <= a;
    layer1_outputs(1467) <= a xor b;
    layer1_outputs(1468) <= a or b;
    layer1_outputs(1469) <= not b or a;
    layer1_outputs(1470) <= a;
    layer1_outputs(1471) <= a xor b;
    layer1_outputs(1472) <= a or b;
    layer1_outputs(1473) <= a xor b;
    layer1_outputs(1474) <= a xor b;
    layer1_outputs(1475) <= not b;
    layer1_outputs(1476) <= b and not a;
    layer1_outputs(1477) <= not b;
    layer1_outputs(1478) <= a;
    layer1_outputs(1479) <= not (a and b);
    layer1_outputs(1480) <= not (a or b);
    layer1_outputs(1481) <= not (a and b);
    layer1_outputs(1482) <= b;
    layer1_outputs(1483) <= not (a xor b);
    layer1_outputs(1484) <= 1'b1;
    layer1_outputs(1485) <= a and b;
    layer1_outputs(1486) <= not a;
    layer1_outputs(1487) <= a;
    layer1_outputs(1488) <= b;
    layer1_outputs(1489) <= not (a xor b);
    layer1_outputs(1490) <= not a or b;
    layer1_outputs(1491) <= a;
    layer1_outputs(1492) <= a xor b;
    layer1_outputs(1493) <= a;
    layer1_outputs(1494) <= b;
    layer1_outputs(1495) <= b and not a;
    layer1_outputs(1496) <= a and b;
    layer1_outputs(1497) <= not b;
    layer1_outputs(1498) <= not (a or b);
    layer1_outputs(1499) <= a or b;
    layer1_outputs(1500) <= a or b;
    layer1_outputs(1501) <= b;
    layer1_outputs(1502) <= not b or a;
    layer1_outputs(1503) <= a xor b;
    layer1_outputs(1504) <= a xor b;
    layer1_outputs(1505) <= not a or b;
    layer1_outputs(1506) <= a;
    layer1_outputs(1507) <= not a;
    layer1_outputs(1508) <= not (a xor b);
    layer1_outputs(1509) <= not a;
    layer1_outputs(1510) <= not a or b;
    layer1_outputs(1511) <= not a;
    layer1_outputs(1512) <= not (a xor b);
    layer1_outputs(1513) <= not a or b;
    layer1_outputs(1514) <= b;
    layer1_outputs(1515) <= not b;
    layer1_outputs(1516) <= a and b;
    layer1_outputs(1517) <= a and not b;
    layer1_outputs(1518) <= not b or a;
    layer1_outputs(1519) <= a xor b;
    layer1_outputs(1520) <= a;
    layer1_outputs(1521) <= not (a and b);
    layer1_outputs(1522) <= not (a xor b);
    layer1_outputs(1523) <= b;
    layer1_outputs(1524) <= b;
    layer1_outputs(1525) <= not b;
    layer1_outputs(1526) <= not b or a;
    layer1_outputs(1527) <= not b;
    layer1_outputs(1528) <= not (a xor b);
    layer1_outputs(1529) <= not a;
    layer1_outputs(1530) <= not b or a;
    layer1_outputs(1531) <= b;
    layer1_outputs(1532) <= a and not b;
    layer1_outputs(1533) <= b;
    layer1_outputs(1534) <= a and b;
    layer1_outputs(1535) <= a;
    layer1_outputs(1536) <= 1'b1;
    layer1_outputs(1537) <= a and b;
    layer1_outputs(1538) <= not (a and b);
    layer1_outputs(1539) <= a;
    layer1_outputs(1540) <= b;
    layer1_outputs(1541) <= a and b;
    layer1_outputs(1542) <= not a;
    layer1_outputs(1543) <= a;
    layer1_outputs(1544) <= a;
    layer1_outputs(1545) <= not b or a;
    layer1_outputs(1546) <= not a;
    layer1_outputs(1547) <= a and not b;
    layer1_outputs(1548) <= b and not a;
    layer1_outputs(1549) <= not b or a;
    layer1_outputs(1550) <= not a;
    layer1_outputs(1551) <= not (a and b);
    layer1_outputs(1552) <= not (a or b);
    layer1_outputs(1553) <= not a or b;
    layer1_outputs(1554) <= b and not a;
    layer1_outputs(1555) <= not (a or b);
    layer1_outputs(1556) <= not (a xor b);
    layer1_outputs(1557) <= b and not a;
    layer1_outputs(1558) <= a and not b;
    layer1_outputs(1559) <= not a or b;
    layer1_outputs(1560) <= a and not b;
    layer1_outputs(1561) <= a and b;
    layer1_outputs(1562) <= not b or a;
    layer1_outputs(1563) <= a;
    layer1_outputs(1564) <= not b;
    layer1_outputs(1565) <= a and b;
    layer1_outputs(1566) <= a;
    layer1_outputs(1567) <= not (a or b);
    layer1_outputs(1568) <= not a;
    layer1_outputs(1569) <= b and not a;
    layer1_outputs(1570) <= not a;
    layer1_outputs(1571) <= not (a and b);
    layer1_outputs(1572) <= not (a or b);
    layer1_outputs(1573) <= not a;
    layer1_outputs(1574) <= not a;
    layer1_outputs(1575) <= not (a or b);
    layer1_outputs(1576) <= a;
    layer1_outputs(1577) <= a xor b;
    layer1_outputs(1578) <= not (a and b);
    layer1_outputs(1579) <= not a or b;
    layer1_outputs(1580) <= not (a or b);
    layer1_outputs(1581) <= a or b;
    layer1_outputs(1582) <= b;
    layer1_outputs(1583) <= not (a and b);
    layer1_outputs(1584) <= a or b;
    layer1_outputs(1585) <= b;
    layer1_outputs(1586) <= not b;
    layer1_outputs(1587) <= not (a or b);
    layer1_outputs(1588) <= not a;
    layer1_outputs(1589) <= a or b;
    layer1_outputs(1590) <= not (a and b);
    layer1_outputs(1591) <= not a;
    layer1_outputs(1592) <= a;
    layer1_outputs(1593) <= b and not a;
    layer1_outputs(1594) <= b;
    layer1_outputs(1595) <= not (a and b);
    layer1_outputs(1596) <= not b;
    layer1_outputs(1597) <= not a;
    layer1_outputs(1598) <= not b;
    layer1_outputs(1599) <= not b;
    layer1_outputs(1600) <= b and not a;
    layer1_outputs(1601) <= 1'b1;
    layer1_outputs(1602) <= a;
    layer1_outputs(1603) <= not a;
    layer1_outputs(1604) <= b;
    layer1_outputs(1605) <= not (a xor b);
    layer1_outputs(1606) <= a and b;
    layer1_outputs(1607) <= b and not a;
    layer1_outputs(1608) <= a;
    layer1_outputs(1609) <= a and not b;
    layer1_outputs(1610) <= not (a xor b);
    layer1_outputs(1611) <= 1'b0;
    layer1_outputs(1612) <= not b;
    layer1_outputs(1613) <= a or b;
    layer1_outputs(1614) <= not a or b;
    layer1_outputs(1615) <= a or b;
    layer1_outputs(1616) <= b;
    layer1_outputs(1617) <= not (a and b);
    layer1_outputs(1618) <= not (a and b);
    layer1_outputs(1619) <= a xor b;
    layer1_outputs(1620) <= not b;
    layer1_outputs(1621) <= not (a xor b);
    layer1_outputs(1622) <= not (a xor b);
    layer1_outputs(1623) <= b;
    layer1_outputs(1624) <= not b or a;
    layer1_outputs(1625) <= not b;
    layer1_outputs(1626) <= not a or b;
    layer1_outputs(1627) <= not a;
    layer1_outputs(1628) <= a and b;
    layer1_outputs(1629) <= a or b;
    layer1_outputs(1630) <= a and b;
    layer1_outputs(1631) <= 1'b0;
    layer1_outputs(1632) <= a or b;
    layer1_outputs(1633) <= a and not b;
    layer1_outputs(1634) <= not b or a;
    layer1_outputs(1635) <= b;
    layer1_outputs(1636) <= b and not a;
    layer1_outputs(1637) <= a and b;
    layer1_outputs(1638) <= 1'b1;
    layer1_outputs(1639) <= not a or b;
    layer1_outputs(1640) <= a and b;
    layer1_outputs(1641) <= not b or a;
    layer1_outputs(1642) <= a and not b;
    layer1_outputs(1643) <= not a;
    layer1_outputs(1644) <= not b;
    layer1_outputs(1645) <= b and not a;
    layer1_outputs(1646) <= a;
    layer1_outputs(1647) <= not a or b;
    layer1_outputs(1648) <= b;
    layer1_outputs(1649) <= b;
    layer1_outputs(1650) <= not b;
    layer1_outputs(1651) <= a and not b;
    layer1_outputs(1652) <= not a or b;
    layer1_outputs(1653) <= a or b;
    layer1_outputs(1654) <= not (a and b);
    layer1_outputs(1655) <= a and b;
    layer1_outputs(1656) <= not a;
    layer1_outputs(1657) <= a;
    layer1_outputs(1658) <= a and not b;
    layer1_outputs(1659) <= not a;
    layer1_outputs(1660) <= a;
    layer1_outputs(1661) <= not (a and b);
    layer1_outputs(1662) <= not (a and b);
    layer1_outputs(1663) <= 1'b1;
    layer1_outputs(1664) <= a and not b;
    layer1_outputs(1665) <= not a;
    layer1_outputs(1666) <= b;
    layer1_outputs(1667) <= not a or b;
    layer1_outputs(1668) <= not b or a;
    layer1_outputs(1669) <= a;
    layer1_outputs(1670) <= a;
    layer1_outputs(1671) <= a or b;
    layer1_outputs(1672) <= a xor b;
    layer1_outputs(1673) <= b and not a;
    layer1_outputs(1674) <= a and b;
    layer1_outputs(1675) <= not b or a;
    layer1_outputs(1676) <= not (a and b);
    layer1_outputs(1677) <= a and not b;
    layer1_outputs(1678) <= a and not b;
    layer1_outputs(1679) <= a;
    layer1_outputs(1680) <= a or b;
    layer1_outputs(1681) <= not (a and b);
    layer1_outputs(1682) <= 1'b0;
    layer1_outputs(1683) <= a;
    layer1_outputs(1684) <= not a or b;
    layer1_outputs(1685) <= not b or a;
    layer1_outputs(1686) <= a or b;
    layer1_outputs(1687) <= not b;
    layer1_outputs(1688) <= not (a xor b);
    layer1_outputs(1689) <= not b;
    layer1_outputs(1690) <= a or b;
    layer1_outputs(1691) <= a or b;
    layer1_outputs(1692) <= not (a or b);
    layer1_outputs(1693) <= not a or b;
    layer1_outputs(1694) <= not b or a;
    layer1_outputs(1695) <= a and not b;
    layer1_outputs(1696) <= not b;
    layer1_outputs(1697) <= not b;
    layer1_outputs(1698) <= not b;
    layer1_outputs(1699) <= 1'b0;
    layer1_outputs(1700) <= a and b;
    layer1_outputs(1701) <= a;
    layer1_outputs(1702) <= not b or a;
    layer1_outputs(1703) <= a;
    layer1_outputs(1704) <= a or b;
    layer1_outputs(1705) <= b and not a;
    layer1_outputs(1706) <= b and not a;
    layer1_outputs(1707) <= a or b;
    layer1_outputs(1708) <= 1'b0;
    layer1_outputs(1709) <= not (a and b);
    layer1_outputs(1710) <= a and not b;
    layer1_outputs(1711) <= not b;
    layer1_outputs(1712) <= not (a or b);
    layer1_outputs(1713) <= b and not a;
    layer1_outputs(1714) <= not b;
    layer1_outputs(1715) <= not (a or b);
    layer1_outputs(1716) <= not b;
    layer1_outputs(1717) <= a xor b;
    layer1_outputs(1718) <= not (a and b);
    layer1_outputs(1719) <= a and b;
    layer1_outputs(1720) <= a;
    layer1_outputs(1721) <= b;
    layer1_outputs(1722) <= not a;
    layer1_outputs(1723) <= not b or a;
    layer1_outputs(1724) <= 1'b1;
    layer1_outputs(1725) <= b;
    layer1_outputs(1726) <= a and not b;
    layer1_outputs(1727) <= a and not b;
    layer1_outputs(1728) <= not a;
    layer1_outputs(1729) <= not a;
    layer1_outputs(1730) <= not b or a;
    layer1_outputs(1731) <= b;
    layer1_outputs(1732) <= not a or b;
    layer1_outputs(1733) <= not b or a;
    layer1_outputs(1734) <= not b or a;
    layer1_outputs(1735) <= not b;
    layer1_outputs(1736) <= b and not a;
    layer1_outputs(1737) <= b;
    layer1_outputs(1738) <= not (a and b);
    layer1_outputs(1739) <= not a or b;
    layer1_outputs(1740) <= not a;
    layer1_outputs(1741) <= not (a and b);
    layer1_outputs(1742) <= not (a xor b);
    layer1_outputs(1743) <= not b or a;
    layer1_outputs(1744) <= not a or b;
    layer1_outputs(1745) <= a and b;
    layer1_outputs(1746) <= not (a and b);
    layer1_outputs(1747) <= not b or a;
    layer1_outputs(1748) <= a;
    layer1_outputs(1749) <= a xor b;
    layer1_outputs(1750) <= 1'b0;
    layer1_outputs(1751) <= not a;
    layer1_outputs(1752) <= a and not b;
    layer1_outputs(1753) <= not b;
    layer1_outputs(1754) <= a and not b;
    layer1_outputs(1755) <= not a or b;
    layer1_outputs(1756) <= b and not a;
    layer1_outputs(1757) <= not (a xor b);
    layer1_outputs(1758) <= not (a xor b);
    layer1_outputs(1759) <= a xor b;
    layer1_outputs(1760) <= not (a or b);
    layer1_outputs(1761) <= b;
    layer1_outputs(1762) <= a;
    layer1_outputs(1763) <= a and not b;
    layer1_outputs(1764) <= not b;
    layer1_outputs(1765) <= a;
    layer1_outputs(1766) <= a;
    layer1_outputs(1767) <= not (a xor b);
    layer1_outputs(1768) <= not b;
    layer1_outputs(1769) <= not (a or b);
    layer1_outputs(1770) <= b and not a;
    layer1_outputs(1771) <= a or b;
    layer1_outputs(1772) <= not a;
    layer1_outputs(1773) <= a or b;
    layer1_outputs(1774) <= a;
    layer1_outputs(1775) <= not b or a;
    layer1_outputs(1776) <= b;
    layer1_outputs(1777) <= not a;
    layer1_outputs(1778) <= b;
    layer1_outputs(1779) <= not a;
    layer1_outputs(1780) <= not (a xor b);
    layer1_outputs(1781) <= not (a or b);
    layer1_outputs(1782) <= a;
    layer1_outputs(1783) <= b;
    layer1_outputs(1784) <= not b;
    layer1_outputs(1785) <= b;
    layer1_outputs(1786) <= not b or a;
    layer1_outputs(1787) <= b;
    layer1_outputs(1788) <= a;
    layer1_outputs(1789) <= b and not a;
    layer1_outputs(1790) <= a and not b;
    layer1_outputs(1791) <= not a;
    layer1_outputs(1792) <= not (a and b);
    layer1_outputs(1793) <= b;
    layer1_outputs(1794) <= b;
    layer1_outputs(1795) <= not b;
    layer1_outputs(1796) <= a xor b;
    layer1_outputs(1797) <= not b or a;
    layer1_outputs(1798) <= 1'b1;
    layer1_outputs(1799) <= b;
    layer1_outputs(1800) <= not b;
    layer1_outputs(1801) <= b;
    layer1_outputs(1802) <= 1'b1;
    layer1_outputs(1803) <= not b;
    layer1_outputs(1804) <= b and not a;
    layer1_outputs(1805) <= not a;
    layer1_outputs(1806) <= a or b;
    layer1_outputs(1807) <= not (a xor b);
    layer1_outputs(1808) <= not (a and b);
    layer1_outputs(1809) <= not b;
    layer1_outputs(1810) <= a and not b;
    layer1_outputs(1811) <= not (a or b);
    layer1_outputs(1812) <= 1'b0;
    layer1_outputs(1813) <= a and b;
    layer1_outputs(1814) <= not b;
    layer1_outputs(1815) <= a xor b;
    layer1_outputs(1816) <= not a or b;
    layer1_outputs(1817) <= not (a and b);
    layer1_outputs(1818) <= not b;
    layer1_outputs(1819) <= b and not a;
    layer1_outputs(1820) <= not a or b;
    layer1_outputs(1821) <= a and not b;
    layer1_outputs(1822) <= a;
    layer1_outputs(1823) <= a or b;
    layer1_outputs(1824) <= b;
    layer1_outputs(1825) <= b;
    layer1_outputs(1826) <= a and b;
    layer1_outputs(1827) <= not b;
    layer1_outputs(1828) <= a and not b;
    layer1_outputs(1829) <= not (a or b);
    layer1_outputs(1830) <= not b or a;
    layer1_outputs(1831) <= a;
    layer1_outputs(1832) <= not (a or b);
    layer1_outputs(1833) <= not (a and b);
    layer1_outputs(1834) <= 1'b1;
    layer1_outputs(1835) <= not b;
    layer1_outputs(1836) <= not (a and b);
    layer1_outputs(1837) <= a;
    layer1_outputs(1838) <= not b;
    layer1_outputs(1839) <= not a;
    layer1_outputs(1840) <= b and not a;
    layer1_outputs(1841) <= b;
    layer1_outputs(1842) <= a;
    layer1_outputs(1843) <= b;
    layer1_outputs(1844) <= a xor b;
    layer1_outputs(1845) <= a or b;
    layer1_outputs(1846) <= not b;
    layer1_outputs(1847) <= b;
    layer1_outputs(1848) <= not b or a;
    layer1_outputs(1849) <= b and not a;
    layer1_outputs(1850) <= b;
    layer1_outputs(1851) <= b and not a;
    layer1_outputs(1852) <= a;
    layer1_outputs(1853) <= a;
    layer1_outputs(1854) <= 1'b1;
    layer1_outputs(1855) <= not b;
    layer1_outputs(1856) <= a and b;
    layer1_outputs(1857) <= not (a xor b);
    layer1_outputs(1858) <= not b;
    layer1_outputs(1859) <= a;
    layer1_outputs(1860) <= not (a or b);
    layer1_outputs(1861) <= b;
    layer1_outputs(1862) <= a or b;
    layer1_outputs(1863) <= a and not b;
    layer1_outputs(1864) <= a and b;
    layer1_outputs(1865) <= not (a or b);
    layer1_outputs(1866) <= not b or a;
    layer1_outputs(1867) <= a;
    layer1_outputs(1868) <= not a;
    layer1_outputs(1869) <= not a;
    layer1_outputs(1870) <= not a or b;
    layer1_outputs(1871) <= not (a and b);
    layer1_outputs(1872) <= a xor b;
    layer1_outputs(1873) <= a and not b;
    layer1_outputs(1874) <= not (a and b);
    layer1_outputs(1875) <= a and b;
    layer1_outputs(1876) <= not a;
    layer1_outputs(1877) <= not a;
    layer1_outputs(1878) <= not (a or b);
    layer1_outputs(1879) <= a and not b;
    layer1_outputs(1880) <= not a or b;
    layer1_outputs(1881) <= not b;
    layer1_outputs(1882) <= b and not a;
    layer1_outputs(1883) <= not a;
    layer1_outputs(1884) <= not b or a;
    layer1_outputs(1885) <= a and not b;
    layer1_outputs(1886) <= not (a and b);
    layer1_outputs(1887) <= b and not a;
    layer1_outputs(1888) <= a;
    layer1_outputs(1889) <= a and not b;
    layer1_outputs(1890) <= not (a and b);
    layer1_outputs(1891) <= not b;
    layer1_outputs(1892) <= a;
    layer1_outputs(1893) <= not (a or b);
    layer1_outputs(1894) <= b;
    layer1_outputs(1895) <= a;
    layer1_outputs(1896) <= not a;
    layer1_outputs(1897) <= a and not b;
    layer1_outputs(1898) <= b and not a;
    layer1_outputs(1899) <= a and b;
    layer1_outputs(1900) <= a or b;
    layer1_outputs(1901) <= not b;
    layer1_outputs(1902) <= not b or a;
    layer1_outputs(1903) <= a;
    layer1_outputs(1904) <= not b or a;
    layer1_outputs(1905) <= b;
    layer1_outputs(1906) <= a and not b;
    layer1_outputs(1907) <= not b;
    layer1_outputs(1908) <= not (a and b);
    layer1_outputs(1909) <= a;
    layer1_outputs(1910) <= a or b;
    layer1_outputs(1911) <= not a;
    layer1_outputs(1912) <= a and b;
    layer1_outputs(1913) <= not (a xor b);
    layer1_outputs(1914) <= a and b;
    layer1_outputs(1915) <= not (a and b);
    layer1_outputs(1916) <= a and not b;
    layer1_outputs(1917) <= not (a and b);
    layer1_outputs(1918) <= a and b;
    layer1_outputs(1919) <= b and not a;
    layer1_outputs(1920) <= b;
    layer1_outputs(1921) <= not b;
    layer1_outputs(1922) <= b;
    layer1_outputs(1923) <= not a or b;
    layer1_outputs(1924) <= a xor b;
    layer1_outputs(1925) <= not (a and b);
    layer1_outputs(1926) <= a xor b;
    layer1_outputs(1927) <= a and not b;
    layer1_outputs(1928) <= not b;
    layer1_outputs(1929) <= a or b;
    layer1_outputs(1930) <= not (a xor b);
    layer1_outputs(1931) <= b and not a;
    layer1_outputs(1932) <= a or b;
    layer1_outputs(1933) <= b;
    layer1_outputs(1934) <= not (a xor b);
    layer1_outputs(1935) <= not (a or b);
    layer1_outputs(1936) <= a or b;
    layer1_outputs(1937) <= not (a and b);
    layer1_outputs(1938) <= not b;
    layer1_outputs(1939) <= not b or a;
    layer1_outputs(1940) <= a xor b;
    layer1_outputs(1941) <= not (a and b);
    layer1_outputs(1942) <= a;
    layer1_outputs(1943) <= a and not b;
    layer1_outputs(1944) <= b;
    layer1_outputs(1945) <= a;
    layer1_outputs(1946) <= a and not b;
    layer1_outputs(1947) <= not b;
    layer1_outputs(1948) <= not (a or b);
    layer1_outputs(1949) <= a xor b;
    layer1_outputs(1950) <= not (a xor b);
    layer1_outputs(1951) <= not b;
    layer1_outputs(1952) <= not b;
    layer1_outputs(1953) <= not (a or b);
    layer1_outputs(1954) <= not b or a;
    layer1_outputs(1955) <= a xor b;
    layer1_outputs(1956) <= a and not b;
    layer1_outputs(1957) <= not b;
    layer1_outputs(1958) <= not a;
    layer1_outputs(1959) <= a xor b;
    layer1_outputs(1960) <= not a or b;
    layer1_outputs(1961) <= a and b;
    layer1_outputs(1962) <= a xor b;
    layer1_outputs(1963) <= not (a xor b);
    layer1_outputs(1964) <= not b or a;
    layer1_outputs(1965) <= a and not b;
    layer1_outputs(1966) <= not (a or b);
    layer1_outputs(1967) <= b;
    layer1_outputs(1968) <= not b or a;
    layer1_outputs(1969) <= a xor b;
    layer1_outputs(1970) <= not (a xor b);
    layer1_outputs(1971) <= a xor b;
    layer1_outputs(1972) <= not b or a;
    layer1_outputs(1973) <= not a;
    layer1_outputs(1974) <= not a;
    layer1_outputs(1975) <= not (a and b);
    layer1_outputs(1976) <= a;
    layer1_outputs(1977) <= not a;
    layer1_outputs(1978) <= not a;
    layer1_outputs(1979) <= a;
    layer1_outputs(1980) <= b;
    layer1_outputs(1981) <= b;
    layer1_outputs(1982) <= a and b;
    layer1_outputs(1983) <= b;
    layer1_outputs(1984) <= a and not b;
    layer1_outputs(1985) <= a or b;
    layer1_outputs(1986) <= a and b;
    layer1_outputs(1987) <= a and not b;
    layer1_outputs(1988) <= not b;
    layer1_outputs(1989) <= not a or b;
    layer1_outputs(1990) <= not b;
    layer1_outputs(1991) <= not a or b;
    layer1_outputs(1992) <= b and not a;
    layer1_outputs(1993) <= not (a or b);
    layer1_outputs(1994) <= b and not a;
    layer1_outputs(1995) <= not (a or b);
    layer1_outputs(1996) <= not (a or b);
    layer1_outputs(1997) <= not b or a;
    layer1_outputs(1998) <= not (a or b);
    layer1_outputs(1999) <= 1'b0;
    layer1_outputs(2000) <= not a or b;
    layer1_outputs(2001) <= not b or a;
    layer1_outputs(2002) <= a or b;
    layer1_outputs(2003) <= not a;
    layer1_outputs(2004) <= not b;
    layer1_outputs(2005) <= not b;
    layer1_outputs(2006) <= a and b;
    layer1_outputs(2007) <= b;
    layer1_outputs(2008) <= a or b;
    layer1_outputs(2009) <= 1'b1;
    layer1_outputs(2010) <= not b or a;
    layer1_outputs(2011) <= b;
    layer1_outputs(2012) <= not (a or b);
    layer1_outputs(2013) <= a;
    layer1_outputs(2014) <= not a;
    layer1_outputs(2015) <= a and not b;
    layer1_outputs(2016) <= not b or a;
    layer1_outputs(2017) <= not b;
    layer1_outputs(2018) <= not a or b;
    layer1_outputs(2019) <= not b;
    layer1_outputs(2020) <= b;
    layer1_outputs(2021) <= not b;
    layer1_outputs(2022) <= not a or b;
    layer1_outputs(2023) <= a or b;
    layer1_outputs(2024) <= not a or b;
    layer1_outputs(2025) <= not a;
    layer1_outputs(2026) <= not (a or b);
    layer1_outputs(2027) <= a;
    layer1_outputs(2028) <= not a;
    layer1_outputs(2029) <= not b or a;
    layer1_outputs(2030) <= not (a or b);
    layer1_outputs(2031) <= 1'b0;
    layer1_outputs(2032) <= not a or b;
    layer1_outputs(2033) <= not b;
    layer1_outputs(2034) <= not a or b;
    layer1_outputs(2035) <= not b;
    layer1_outputs(2036) <= b and not a;
    layer1_outputs(2037) <= not (a xor b);
    layer1_outputs(2038) <= not a;
    layer1_outputs(2039) <= b;
    layer1_outputs(2040) <= a and not b;
    layer1_outputs(2041) <= not b or a;
    layer1_outputs(2042) <= 1'b0;
    layer1_outputs(2043) <= not b;
    layer1_outputs(2044) <= a;
    layer1_outputs(2045) <= not b;
    layer1_outputs(2046) <= not a or b;
    layer1_outputs(2047) <= not a;
    layer1_outputs(2048) <= not b or a;
    layer1_outputs(2049) <= b;
    layer1_outputs(2050) <= not (a or b);
    layer1_outputs(2051) <= b;
    layer1_outputs(2052) <= 1'b0;
    layer1_outputs(2053) <= a or b;
    layer1_outputs(2054) <= not b or a;
    layer1_outputs(2055) <= a;
    layer1_outputs(2056) <= a and b;
    layer1_outputs(2057) <= not (a and b);
    layer1_outputs(2058) <= not a or b;
    layer1_outputs(2059) <= not (a and b);
    layer1_outputs(2060) <= not b;
    layer1_outputs(2061) <= a and b;
    layer1_outputs(2062) <= b;
    layer1_outputs(2063) <= not (a or b);
    layer1_outputs(2064) <= not a;
    layer1_outputs(2065) <= not (a xor b);
    layer1_outputs(2066) <= not b or a;
    layer1_outputs(2067) <= b and not a;
    layer1_outputs(2068) <= a xor b;
    layer1_outputs(2069) <= a and not b;
    layer1_outputs(2070) <= not (a xor b);
    layer1_outputs(2071) <= a or b;
    layer1_outputs(2072) <= a;
    layer1_outputs(2073) <= not b;
    layer1_outputs(2074) <= not (a and b);
    layer1_outputs(2075) <= a;
    layer1_outputs(2076) <= not a or b;
    layer1_outputs(2077) <= a;
    layer1_outputs(2078) <= not a;
    layer1_outputs(2079) <= not a;
    layer1_outputs(2080) <= not a or b;
    layer1_outputs(2081) <= b;
    layer1_outputs(2082) <= a and b;
    layer1_outputs(2083) <= not a;
    layer1_outputs(2084) <= not (a xor b);
    layer1_outputs(2085) <= a and b;
    layer1_outputs(2086) <= a;
    layer1_outputs(2087) <= not (a xor b);
    layer1_outputs(2088) <= b;
    layer1_outputs(2089) <= a;
    layer1_outputs(2090) <= a;
    layer1_outputs(2091) <= b and not a;
    layer1_outputs(2092) <= a or b;
    layer1_outputs(2093) <= a and b;
    layer1_outputs(2094) <= not a or b;
    layer1_outputs(2095) <= a and b;
    layer1_outputs(2096) <= not (a and b);
    layer1_outputs(2097) <= 1'b0;
    layer1_outputs(2098) <= not (a xor b);
    layer1_outputs(2099) <= not a;
    layer1_outputs(2100) <= not a or b;
    layer1_outputs(2101) <= a and not b;
    layer1_outputs(2102) <= not b or a;
    layer1_outputs(2103) <= not b;
    layer1_outputs(2104) <= b;
    layer1_outputs(2105) <= b;
    layer1_outputs(2106) <= a and not b;
    layer1_outputs(2107) <= a and b;
    layer1_outputs(2108) <= not b or a;
    layer1_outputs(2109) <= not b;
    layer1_outputs(2110) <= b;
    layer1_outputs(2111) <= not a;
    layer1_outputs(2112) <= b and not a;
    layer1_outputs(2113) <= a xor b;
    layer1_outputs(2114) <= not (a or b);
    layer1_outputs(2115) <= a and not b;
    layer1_outputs(2116) <= a and b;
    layer1_outputs(2117) <= not (a xor b);
    layer1_outputs(2118) <= not a;
    layer1_outputs(2119) <= a and b;
    layer1_outputs(2120) <= not a;
    layer1_outputs(2121) <= not b;
    layer1_outputs(2122) <= a or b;
    layer1_outputs(2123) <= not a;
    layer1_outputs(2124) <= a;
    layer1_outputs(2125) <= a or b;
    layer1_outputs(2126) <= not (a or b);
    layer1_outputs(2127) <= b;
    layer1_outputs(2128) <= a and not b;
    layer1_outputs(2129) <= not b or a;
    layer1_outputs(2130) <= not a or b;
    layer1_outputs(2131) <= not (a or b);
    layer1_outputs(2132) <= not (a or b);
    layer1_outputs(2133) <= a xor b;
    layer1_outputs(2134) <= not a or b;
    layer1_outputs(2135) <= a and b;
    layer1_outputs(2136) <= not a;
    layer1_outputs(2137) <= not (a or b);
    layer1_outputs(2138) <= a and b;
    layer1_outputs(2139) <= not (a xor b);
    layer1_outputs(2140) <= not (a and b);
    layer1_outputs(2141) <= a;
    layer1_outputs(2142) <= a and not b;
    layer1_outputs(2143) <= a and not b;
    layer1_outputs(2144) <= b;
    layer1_outputs(2145) <= a and not b;
    layer1_outputs(2146) <= not b;
    layer1_outputs(2147) <= a and b;
    layer1_outputs(2148) <= not b or a;
    layer1_outputs(2149) <= not a or b;
    layer1_outputs(2150) <= a;
    layer1_outputs(2151) <= a or b;
    layer1_outputs(2152) <= a or b;
    layer1_outputs(2153) <= a;
    layer1_outputs(2154) <= b;
    layer1_outputs(2155) <= a and b;
    layer1_outputs(2156) <= 1'b1;
    layer1_outputs(2157) <= not b;
    layer1_outputs(2158) <= not a;
    layer1_outputs(2159) <= a and not b;
    layer1_outputs(2160) <= b;
    layer1_outputs(2161) <= not b;
    layer1_outputs(2162) <= not (a or b);
    layer1_outputs(2163) <= a or b;
    layer1_outputs(2164) <= a and not b;
    layer1_outputs(2165) <= a and not b;
    layer1_outputs(2166) <= not a;
    layer1_outputs(2167) <= not b or a;
    layer1_outputs(2168) <= not b;
    layer1_outputs(2169) <= 1'b1;
    layer1_outputs(2170) <= not b or a;
    layer1_outputs(2171) <= a;
    layer1_outputs(2172) <= a and b;
    layer1_outputs(2173) <= b;
    layer1_outputs(2174) <= not a;
    layer1_outputs(2175) <= b;
    layer1_outputs(2176) <= not a;
    layer1_outputs(2177) <= not (a and b);
    layer1_outputs(2178) <= a;
    layer1_outputs(2179) <= b and not a;
    layer1_outputs(2180) <= not (a xor b);
    layer1_outputs(2181) <= b;
    layer1_outputs(2182) <= not a;
    layer1_outputs(2183) <= not b;
    layer1_outputs(2184) <= not a;
    layer1_outputs(2185) <= not (a or b);
    layer1_outputs(2186) <= not (a or b);
    layer1_outputs(2187) <= b;
    layer1_outputs(2188) <= not a;
    layer1_outputs(2189) <= a and not b;
    layer1_outputs(2190) <= not (a xor b);
    layer1_outputs(2191) <= a;
    layer1_outputs(2192) <= not (a or b);
    layer1_outputs(2193) <= a;
    layer1_outputs(2194) <= a and not b;
    layer1_outputs(2195) <= a and not b;
    layer1_outputs(2196) <= not b;
    layer1_outputs(2197) <= a and not b;
    layer1_outputs(2198) <= a xor b;
    layer1_outputs(2199) <= a and b;
    layer1_outputs(2200) <= a xor b;
    layer1_outputs(2201) <= b;
    layer1_outputs(2202) <= not a or b;
    layer1_outputs(2203) <= not (a and b);
    layer1_outputs(2204) <= not (a and b);
    layer1_outputs(2205) <= a or b;
    layer1_outputs(2206) <= not (a or b);
    layer1_outputs(2207) <= not a;
    layer1_outputs(2208) <= not a;
    layer1_outputs(2209) <= not (a and b);
    layer1_outputs(2210) <= b and not a;
    layer1_outputs(2211) <= not (a and b);
    layer1_outputs(2212) <= not b or a;
    layer1_outputs(2213) <= b and not a;
    layer1_outputs(2214) <= b;
    layer1_outputs(2215) <= a and b;
    layer1_outputs(2216) <= 1'b1;
    layer1_outputs(2217) <= b;
    layer1_outputs(2218) <= not (a or b);
    layer1_outputs(2219) <= not a;
    layer1_outputs(2220) <= not (a and b);
    layer1_outputs(2221) <= b;
    layer1_outputs(2222) <= 1'b0;
    layer1_outputs(2223) <= a or b;
    layer1_outputs(2224) <= a and b;
    layer1_outputs(2225) <= not (a and b);
    layer1_outputs(2226) <= not a;
    layer1_outputs(2227) <= not a;
    layer1_outputs(2228) <= a or b;
    layer1_outputs(2229) <= not a or b;
    layer1_outputs(2230) <= a or b;
    layer1_outputs(2231) <= a xor b;
    layer1_outputs(2232) <= not a;
    layer1_outputs(2233) <= not (a xor b);
    layer1_outputs(2234) <= a and not b;
    layer1_outputs(2235) <= not (a xor b);
    layer1_outputs(2236) <= a and not b;
    layer1_outputs(2237) <= a or b;
    layer1_outputs(2238) <= not a or b;
    layer1_outputs(2239) <= a xor b;
    layer1_outputs(2240) <= not (a xor b);
    layer1_outputs(2241) <= a or b;
    layer1_outputs(2242) <= b;
    layer1_outputs(2243) <= b;
    layer1_outputs(2244) <= not b;
    layer1_outputs(2245) <= not a;
    layer1_outputs(2246) <= a;
    layer1_outputs(2247) <= not b;
    layer1_outputs(2248) <= not a;
    layer1_outputs(2249) <= a and b;
    layer1_outputs(2250) <= not (a xor b);
    layer1_outputs(2251) <= a;
    layer1_outputs(2252) <= b and not a;
    layer1_outputs(2253) <= not a;
    layer1_outputs(2254) <= 1'b1;
    layer1_outputs(2255) <= a;
    layer1_outputs(2256) <= not b;
    layer1_outputs(2257) <= b and not a;
    layer1_outputs(2258) <= b;
    layer1_outputs(2259) <= b;
    layer1_outputs(2260) <= b and not a;
    layer1_outputs(2261) <= a;
    layer1_outputs(2262) <= not (a and b);
    layer1_outputs(2263) <= b;
    layer1_outputs(2264) <= a or b;
    layer1_outputs(2265) <= not (a and b);
    layer1_outputs(2266) <= b and not a;
    layer1_outputs(2267) <= a or b;
    layer1_outputs(2268) <= b;
    layer1_outputs(2269) <= b;
    layer1_outputs(2270) <= a;
    layer1_outputs(2271) <= not b or a;
    layer1_outputs(2272) <= a;
    layer1_outputs(2273) <= not b or a;
    layer1_outputs(2274) <= not (a and b);
    layer1_outputs(2275) <= not (a and b);
    layer1_outputs(2276) <= not b;
    layer1_outputs(2277) <= b and not a;
    layer1_outputs(2278) <= a;
    layer1_outputs(2279) <= a and b;
    layer1_outputs(2280) <= not b;
    layer1_outputs(2281) <= b and not a;
    layer1_outputs(2282) <= not b;
    layer1_outputs(2283) <= b and not a;
    layer1_outputs(2284) <= a;
    layer1_outputs(2285) <= a;
    layer1_outputs(2286) <= a;
    layer1_outputs(2287) <= not a;
    layer1_outputs(2288) <= a;
    layer1_outputs(2289) <= a;
    layer1_outputs(2290) <= b;
    layer1_outputs(2291) <= a or b;
    layer1_outputs(2292) <= a or b;
    layer1_outputs(2293) <= not b;
    layer1_outputs(2294) <= a and not b;
    layer1_outputs(2295) <= not a;
    layer1_outputs(2296) <= not (a xor b);
    layer1_outputs(2297) <= b;
    layer1_outputs(2298) <= a;
    layer1_outputs(2299) <= not a;
    layer1_outputs(2300) <= not a;
    layer1_outputs(2301) <= not b or a;
    layer1_outputs(2302) <= a and b;
    layer1_outputs(2303) <= a xor b;
    layer1_outputs(2304) <= not b or a;
    layer1_outputs(2305) <= b and not a;
    layer1_outputs(2306) <= not a;
    layer1_outputs(2307) <= not a or b;
    layer1_outputs(2308) <= b and not a;
    layer1_outputs(2309) <= not b or a;
    layer1_outputs(2310) <= b;
    layer1_outputs(2311) <= not b;
    layer1_outputs(2312) <= not b;
    layer1_outputs(2313) <= not (a xor b);
    layer1_outputs(2314) <= not a;
    layer1_outputs(2315) <= b;
    layer1_outputs(2316) <= b;
    layer1_outputs(2317) <= a;
    layer1_outputs(2318) <= not (a and b);
    layer1_outputs(2319) <= not a or b;
    layer1_outputs(2320) <= a or b;
    layer1_outputs(2321) <= not a;
    layer1_outputs(2322) <= 1'b1;
    layer1_outputs(2323) <= 1'b1;
    layer1_outputs(2324) <= not b;
    layer1_outputs(2325) <= not a or b;
    layer1_outputs(2326) <= not a;
    layer1_outputs(2327) <= a;
    layer1_outputs(2328) <= a;
    layer1_outputs(2329) <= a;
    layer1_outputs(2330) <= b;
    layer1_outputs(2331) <= b;
    layer1_outputs(2332) <= b;
    layer1_outputs(2333) <= a and not b;
    layer1_outputs(2334) <= not b;
    layer1_outputs(2335) <= a xor b;
    layer1_outputs(2336) <= not b or a;
    layer1_outputs(2337) <= b and not a;
    layer1_outputs(2338) <= b;
    layer1_outputs(2339) <= not (a or b);
    layer1_outputs(2340) <= b and not a;
    layer1_outputs(2341) <= b and not a;
    layer1_outputs(2342) <= not (a xor b);
    layer1_outputs(2343) <= not (a and b);
    layer1_outputs(2344) <= not (a xor b);
    layer1_outputs(2345) <= not a;
    layer1_outputs(2346) <= a;
    layer1_outputs(2347) <= not (a xor b);
    layer1_outputs(2348) <= b;
    layer1_outputs(2349) <= not a or b;
    layer1_outputs(2350) <= not (a or b);
    layer1_outputs(2351) <= a;
    layer1_outputs(2352) <= a or b;
    layer1_outputs(2353) <= a and not b;
    layer1_outputs(2354) <= b and not a;
    layer1_outputs(2355) <= b;
    layer1_outputs(2356) <= not b or a;
    layer1_outputs(2357) <= a and not b;
    layer1_outputs(2358) <= not a;
    layer1_outputs(2359) <= a or b;
    layer1_outputs(2360) <= a;
    layer1_outputs(2361) <= not (a xor b);
    layer1_outputs(2362) <= not (a xor b);
    layer1_outputs(2363) <= b;
    layer1_outputs(2364) <= a and not b;
    layer1_outputs(2365) <= not a;
    layer1_outputs(2366) <= b;
    layer1_outputs(2367) <= not (a or b);
    layer1_outputs(2368) <= not b or a;
    layer1_outputs(2369) <= a;
    layer1_outputs(2370) <= 1'b1;
    layer1_outputs(2371) <= not (a or b);
    layer1_outputs(2372) <= a;
    layer1_outputs(2373) <= not b or a;
    layer1_outputs(2374) <= a and not b;
    layer1_outputs(2375) <= a xor b;
    layer1_outputs(2376) <= a and b;
    layer1_outputs(2377) <= b;
    layer1_outputs(2378) <= b;
    layer1_outputs(2379) <= a and b;
    layer1_outputs(2380) <= a or b;
    layer1_outputs(2381) <= b;
    layer1_outputs(2382) <= not a or b;
    layer1_outputs(2383) <= a xor b;
    layer1_outputs(2384) <= a and b;
    layer1_outputs(2385) <= a;
    layer1_outputs(2386) <= not (a and b);
    layer1_outputs(2387) <= b;
    layer1_outputs(2388) <= not b or a;
    layer1_outputs(2389) <= b and not a;
    layer1_outputs(2390) <= a or b;
    layer1_outputs(2391) <= not (a xor b);
    layer1_outputs(2392) <= not b or a;
    layer1_outputs(2393) <= b and not a;
    layer1_outputs(2394) <= not a;
    layer1_outputs(2395) <= not (a and b);
    layer1_outputs(2396) <= a and not b;
    layer1_outputs(2397) <= a or b;
    layer1_outputs(2398) <= not (a or b);
    layer1_outputs(2399) <= b;
    layer1_outputs(2400) <= a and not b;
    layer1_outputs(2401) <= not b or a;
    layer1_outputs(2402) <= a;
    layer1_outputs(2403) <= 1'b1;
    layer1_outputs(2404) <= a xor b;
    layer1_outputs(2405) <= not (a or b);
    layer1_outputs(2406) <= not a;
    layer1_outputs(2407) <= a and not b;
    layer1_outputs(2408) <= not (a or b);
    layer1_outputs(2409) <= not (a and b);
    layer1_outputs(2410) <= a or b;
    layer1_outputs(2411) <= b;
    layer1_outputs(2412) <= a or b;
    layer1_outputs(2413) <= not b;
    layer1_outputs(2414) <= not (a and b);
    layer1_outputs(2415) <= not a;
    layer1_outputs(2416) <= a xor b;
    layer1_outputs(2417) <= not (a and b);
    layer1_outputs(2418) <= a or b;
    layer1_outputs(2419) <= not a or b;
    layer1_outputs(2420) <= not b;
    layer1_outputs(2421) <= not b or a;
    layer1_outputs(2422) <= not a or b;
    layer1_outputs(2423) <= b and not a;
    layer1_outputs(2424) <= a;
    layer1_outputs(2425) <= not (a or b);
    layer1_outputs(2426) <= a or b;
    layer1_outputs(2427) <= not a or b;
    layer1_outputs(2428) <= not a;
    layer1_outputs(2429) <= a or b;
    layer1_outputs(2430) <= not b;
    layer1_outputs(2431) <= a and not b;
    layer1_outputs(2432) <= not b;
    layer1_outputs(2433) <= not b or a;
    layer1_outputs(2434) <= a;
    layer1_outputs(2435) <= not (a xor b);
    layer1_outputs(2436) <= not b;
    layer1_outputs(2437) <= not b or a;
    layer1_outputs(2438) <= not b or a;
    layer1_outputs(2439) <= not b or a;
    layer1_outputs(2440) <= not b or a;
    layer1_outputs(2441) <= b and not a;
    layer1_outputs(2442) <= b;
    layer1_outputs(2443) <= not (a xor b);
    layer1_outputs(2444) <= not b;
    layer1_outputs(2445) <= not a or b;
    layer1_outputs(2446) <= a and not b;
    layer1_outputs(2447) <= a;
    layer1_outputs(2448) <= 1'b0;
    layer1_outputs(2449) <= not (a and b);
    layer1_outputs(2450) <= b;
    layer1_outputs(2451) <= a and b;
    layer1_outputs(2452) <= not a or b;
    layer1_outputs(2453) <= not b or a;
    layer1_outputs(2454) <= a and not b;
    layer1_outputs(2455) <= not a or b;
    layer1_outputs(2456) <= a;
    layer1_outputs(2457) <= not (a and b);
    layer1_outputs(2458) <= a and b;
    layer1_outputs(2459) <= a and not b;
    layer1_outputs(2460) <= 1'b1;
    layer1_outputs(2461) <= not (a or b);
    layer1_outputs(2462) <= not b;
    layer1_outputs(2463) <= a xor b;
    layer1_outputs(2464) <= b;
    layer1_outputs(2465) <= not a or b;
    layer1_outputs(2466) <= b;
    layer1_outputs(2467) <= a;
    layer1_outputs(2468) <= a and not b;
    layer1_outputs(2469) <= a;
    layer1_outputs(2470) <= not (a and b);
    layer1_outputs(2471) <= not (a or b);
    layer1_outputs(2472) <= b and not a;
    layer1_outputs(2473) <= a xor b;
    layer1_outputs(2474) <= not a;
    layer1_outputs(2475) <= a;
    layer1_outputs(2476) <= 1'b0;
    layer1_outputs(2477) <= a;
    layer1_outputs(2478) <= not a;
    layer1_outputs(2479) <= not a;
    layer1_outputs(2480) <= not (a or b);
    layer1_outputs(2481) <= not (a and b);
    layer1_outputs(2482) <= not (a or b);
    layer1_outputs(2483) <= a;
    layer1_outputs(2484) <= not b or a;
    layer1_outputs(2485) <= a or b;
    layer1_outputs(2486) <= a and b;
    layer1_outputs(2487) <= a and b;
    layer1_outputs(2488) <= not b or a;
    layer1_outputs(2489) <= not (a xor b);
    layer1_outputs(2490) <= not b;
    layer1_outputs(2491) <= not a or b;
    layer1_outputs(2492) <= a and b;
    layer1_outputs(2493) <= not a;
    layer1_outputs(2494) <= not b;
    layer1_outputs(2495) <= not a;
    layer1_outputs(2496) <= not (a and b);
    layer1_outputs(2497) <= 1'b0;
    layer1_outputs(2498) <= a and not b;
    layer1_outputs(2499) <= not a or b;
    layer1_outputs(2500) <= a and b;
    layer1_outputs(2501) <= a xor b;
    layer1_outputs(2502) <= a and not b;
    layer1_outputs(2503) <= a;
    layer1_outputs(2504) <= a and b;
    layer1_outputs(2505) <= not b or a;
    layer1_outputs(2506) <= b;
    layer1_outputs(2507) <= a and b;
    layer1_outputs(2508) <= a or b;
    layer1_outputs(2509) <= 1'b1;
    layer1_outputs(2510) <= not (a xor b);
    layer1_outputs(2511) <= not a;
    layer1_outputs(2512) <= a and not b;
    layer1_outputs(2513) <= a;
    layer1_outputs(2514) <= a or b;
    layer1_outputs(2515) <= a and b;
    layer1_outputs(2516) <= not a;
    layer1_outputs(2517) <= not b or a;
    layer1_outputs(2518) <= not a;
    layer1_outputs(2519) <= not a or b;
    layer1_outputs(2520) <= a and not b;
    layer1_outputs(2521) <= b;
    layer1_outputs(2522) <= a and b;
    layer1_outputs(2523) <= a;
    layer1_outputs(2524) <= a xor b;
    layer1_outputs(2525) <= not a;
    layer1_outputs(2526) <= a or b;
    layer1_outputs(2527) <= b and not a;
    layer1_outputs(2528) <= not a;
    layer1_outputs(2529) <= a;
    layer1_outputs(2530) <= a xor b;
    layer1_outputs(2531) <= not (a xor b);
    layer1_outputs(2532) <= a;
    layer1_outputs(2533) <= not a or b;
    layer1_outputs(2534) <= not (a or b);
    layer1_outputs(2535) <= a;
    layer1_outputs(2536) <= not a or b;
    layer1_outputs(2537) <= b;
    layer1_outputs(2538) <= not b;
    layer1_outputs(2539) <= not b;
    layer1_outputs(2540) <= not a or b;
    layer1_outputs(2541) <= not (a xor b);
    layer1_outputs(2542) <= a and not b;
    layer1_outputs(2543) <= a;
    layer1_outputs(2544) <= not b;
    layer1_outputs(2545) <= not a or b;
    layer1_outputs(2546) <= not (a or b);
    layer1_outputs(2547) <= a xor b;
    layer1_outputs(2548) <= a and b;
    layer1_outputs(2549) <= not a;
    layer1_outputs(2550) <= a and b;
    layer1_outputs(2551) <= not a or b;
    layer1_outputs(2552) <= a and b;
    layer1_outputs(2553) <= not (a and b);
    layer1_outputs(2554) <= not a;
    layer1_outputs(2555) <= not (a or b);
    layer1_outputs(2556) <= a;
    layer1_outputs(2557) <= 1'b1;
    layer1_outputs(2558) <= a xor b;
    layer1_outputs(2559) <= not (a and b);
    layer2_outputs(0) <= b and not a;
    layer2_outputs(1) <= not a or b;
    layer2_outputs(2) <= not b;
    layer2_outputs(3) <= a xor b;
    layer2_outputs(4) <= not a or b;
    layer2_outputs(5) <= not a;
    layer2_outputs(6) <= b;
    layer2_outputs(7) <= a and not b;
    layer2_outputs(8) <= a and b;
    layer2_outputs(9) <= not (a and b);
    layer2_outputs(10) <= a;
    layer2_outputs(11) <= b;
    layer2_outputs(12) <= not a;
    layer2_outputs(13) <= not (a xor b);
    layer2_outputs(14) <= b and not a;
    layer2_outputs(15) <= a and b;
    layer2_outputs(16) <= not b;
    layer2_outputs(17) <= not b or a;
    layer2_outputs(18) <= b;
    layer2_outputs(19) <= b and not a;
    layer2_outputs(20) <= a and b;
    layer2_outputs(21) <= a;
    layer2_outputs(22) <= not (a and b);
    layer2_outputs(23) <= not (a and b);
    layer2_outputs(24) <= 1'b0;
    layer2_outputs(25) <= not b;
    layer2_outputs(26) <= a and b;
    layer2_outputs(27) <= a xor b;
    layer2_outputs(28) <= not b or a;
    layer2_outputs(29) <= not a;
    layer2_outputs(30) <= a and not b;
    layer2_outputs(31) <= 1'b1;
    layer2_outputs(32) <= b;
    layer2_outputs(33) <= a;
    layer2_outputs(34) <= a or b;
    layer2_outputs(35) <= b;
    layer2_outputs(36) <= a and b;
    layer2_outputs(37) <= a;
    layer2_outputs(38) <= not b;
    layer2_outputs(39) <= b and not a;
    layer2_outputs(40) <= not (a or b);
    layer2_outputs(41) <= not a;
    layer2_outputs(42) <= not b;
    layer2_outputs(43) <= a and b;
    layer2_outputs(44) <= not b;
    layer2_outputs(45) <= not b;
    layer2_outputs(46) <= not b;
    layer2_outputs(47) <= a and not b;
    layer2_outputs(48) <= not b;
    layer2_outputs(49) <= a and not b;
    layer2_outputs(50) <= b and not a;
    layer2_outputs(51) <= a or b;
    layer2_outputs(52) <= not b;
    layer2_outputs(53) <= a xor b;
    layer2_outputs(54) <= a;
    layer2_outputs(55) <= a xor b;
    layer2_outputs(56) <= not b;
    layer2_outputs(57) <= not b;
    layer2_outputs(58) <= not (a and b);
    layer2_outputs(59) <= a and not b;
    layer2_outputs(60) <= not a;
    layer2_outputs(61) <= not b or a;
    layer2_outputs(62) <= a xor b;
    layer2_outputs(63) <= not b;
    layer2_outputs(64) <= not (a xor b);
    layer2_outputs(65) <= not a;
    layer2_outputs(66) <= not (a and b);
    layer2_outputs(67) <= b;
    layer2_outputs(68) <= b;
    layer2_outputs(69) <= not b;
    layer2_outputs(70) <= not b or a;
    layer2_outputs(71) <= not (a and b);
    layer2_outputs(72) <= b and not a;
    layer2_outputs(73) <= a xor b;
    layer2_outputs(74) <= not a or b;
    layer2_outputs(75) <= 1'b1;
    layer2_outputs(76) <= a and not b;
    layer2_outputs(77) <= a xor b;
    layer2_outputs(78) <= b;
    layer2_outputs(79) <= not (a or b);
    layer2_outputs(80) <= b;
    layer2_outputs(81) <= not a;
    layer2_outputs(82) <= b;
    layer2_outputs(83) <= not a or b;
    layer2_outputs(84) <= b and not a;
    layer2_outputs(85) <= a or b;
    layer2_outputs(86) <= b and not a;
    layer2_outputs(87) <= not b;
    layer2_outputs(88) <= a xor b;
    layer2_outputs(89) <= not a;
    layer2_outputs(90) <= not b;
    layer2_outputs(91) <= a and not b;
    layer2_outputs(92) <= a and not b;
    layer2_outputs(93) <= b;
    layer2_outputs(94) <= b;
    layer2_outputs(95) <= not (a xor b);
    layer2_outputs(96) <= a xor b;
    layer2_outputs(97) <= not a;
    layer2_outputs(98) <= not (a xor b);
    layer2_outputs(99) <= not a;
    layer2_outputs(100) <= b;
    layer2_outputs(101) <= not b or a;
    layer2_outputs(102) <= not b or a;
    layer2_outputs(103) <= not a;
    layer2_outputs(104) <= not a;
    layer2_outputs(105) <= a or b;
    layer2_outputs(106) <= not (a and b);
    layer2_outputs(107) <= not a or b;
    layer2_outputs(108) <= not b or a;
    layer2_outputs(109) <= a;
    layer2_outputs(110) <= b;
    layer2_outputs(111) <= b and not a;
    layer2_outputs(112) <= not (a or b);
    layer2_outputs(113) <= not (a or b);
    layer2_outputs(114) <= not (a or b);
    layer2_outputs(115) <= not (a and b);
    layer2_outputs(116) <= not (a and b);
    layer2_outputs(117) <= a and not b;
    layer2_outputs(118) <= not (a and b);
    layer2_outputs(119) <= b and not a;
    layer2_outputs(120) <= a and b;
    layer2_outputs(121) <= not b;
    layer2_outputs(122) <= a;
    layer2_outputs(123) <= not a;
    layer2_outputs(124) <= b and not a;
    layer2_outputs(125) <= a;
    layer2_outputs(126) <= not (a and b);
    layer2_outputs(127) <= not b;
    layer2_outputs(128) <= not (a and b);
    layer2_outputs(129) <= not a or b;
    layer2_outputs(130) <= not b or a;
    layer2_outputs(131) <= a;
    layer2_outputs(132) <= a and not b;
    layer2_outputs(133) <= not (a or b);
    layer2_outputs(134) <= not (a and b);
    layer2_outputs(135) <= not a;
    layer2_outputs(136) <= not a;
    layer2_outputs(137) <= not (a and b);
    layer2_outputs(138) <= b;
    layer2_outputs(139) <= a xor b;
    layer2_outputs(140) <= a or b;
    layer2_outputs(141) <= a and not b;
    layer2_outputs(142) <= a or b;
    layer2_outputs(143) <= b;
    layer2_outputs(144) <= b and not a;
    layer2_outputs(145) <= a;
    layer2_outputs(146) <= b and not a;
    layer2_outputs(147) <= not a;
    layer2_outputs(148) <= not a or b;
    layer2_outputs(149) <= a xor b;
    layer2_outputs(150) <= not (a or b);
    layer2_outputs(151) <= not (a or b);
    layer2_outputs(152) <= not a;
    layer2_outputs(153) <= b;
    layer2_outputs(154) <= a and not b;
    layer2_outputs(155) <= not (a or b);
    layer2_outputs(156) <= a or b;
    layer2_outputs(157) <= not (a and b);
    layer2_outputs(158) <= not a or b;
    layer2_outputs(159) <= not b or a;
    layer2_outputs(160) <= a and not b;
    layer2_outputs(161) <= a;
    layer2_outputs(162) <= not b;
    layer2_outputs(163) <= not (a or b);
    layer2_outputs(164) <= not (a or b);
    layer2_outputs(165) <= not a or b;
    layer2_outputs(166) <= a and not b;
    layer2_outputs(167) <= not a or b;
    layer2_outputs(168) <= b;
    layer2_outputs(169) <= not a;
    layer2_outputs(170) <= not b or a;
    layer2_outputs(171) <= a or b;
    layer2_outputs(172) <= a xor b;
    layer2_outputs(173) <= 1'b0;
    layer2_outputs(174) <= not a or b;
    layer2_outputs(175) <= a and b;
    layer2_outputs(176) <= a or b;
    layer2_outputs(177) <= not b or a;
    layer2_outputs(178) <= a and b;
    layer2_outputs(179) <= a;
    layer2_outputs(180) <= not b;
    layer2_outputs(181) <= not (a or b);
    layer2_outputs(182) <= not (a xor b);
    layer2_outputs(183) <= a and b;
    layer2_outputs(184) <= a or b;
    layer2_outputs(185) <= a or b;
    layer2_outputs(186) <= a and not b;
    layer2_outputs(187) <= a and not b;
    layer2_outputs(188) <= not a or b;
    layer2_outputs(189) <= not b;
    layer2_outputs(190) <= a;
    layer2_outputs(191) <= a;
    layer2_outputs(192) <= not (a xor b);
    layer2_outputs(193) <= a or b;
    layer2_outputs(194) <= a;
    layer2_outputs(195) <= b and not a;
    layer2_outputs(196) <= not b or a;
    layer2_outputs(197) <= 1'b0;
    layer2_outputs(198) <= not (a or b);
    layer2_outputs(199) <= not b;
    layer2_outputs(200) <= a and b;
    layer2_outputs(201) <= not a;
    layer2_outputs(202) <= b;
    layer2_outputs(203) <= not b;
    layer2_outputs(204) <= b;
    layer2_outputs(205) <= not a or b;
    layer2_outputs(206) <= not b or a;
    layer2_outputs(207) <= a or b;
    layer2_outputs(208) <= a and not b;
    layer2_outputs(209) <= not (a or b);
    layer2_outputs(210) <= b;
    layer2_outputs(211) <= not b;
    layer2_outputs(212) <= a or b;
    layer2_outputs(213) <= a;
    layer2_outputs(214) <= a or b;
    layer2_outputs(215) <= not b or a;
    layer2_outputs(216) <= a and not b;
    layer2_outputs(217) <= not b or a;
    layer2_outputs(218) <= a and not b;
    layer2_outputs(219) <= not (a or b);
    layer2_outputs(220) <= a and b;
    layer2_outputs(221) <= a;
    layer2_outputs(222) <= not b;
    layer2_outputs(223) <= not b;
    layer2_outputs(224) <= not (a xor b);
    layer2_outputs(225) <= b;
    layer2_outputs(226) <= b;
    layer2_outputs(227) <= b;
    layer2_outputs(228) <= a and not b;
    layer2_outputs(229) <= b;
    layer2_outputs(230) <= not b;
    layer2_outputs(231) <= not b;
    layer2_outputs(232) <= a or b;
    layer2_outputs(233) <= b;
    layer2_outputs(234) <= a and not b;
    layer2_outputs(235) <= a or b;
    layer2_outputs(236) <= b and not a;
    layer2_outputs(237) <= b;
    layer2_outputs(238) <= a and not b;
    layer2_outputs(239) <= not (a and b);
    layer2_outputs(240) <= not (a or b);
    layer2_outputs(241) <= a;
    layer2_outputs(242) <= b and not a;
    layer2_outputs(243) <= a or b;
    layer2_outputs(244) <= not a or b;
    layer2_outputs(245) <= b and not a;
    layer2_outputs(246) <= not a;
    layer2_outputs(247) <= a xor b;
    layer2_outputs(248) <= b and not a;
    layer2_outputs(249) <= not (a and b);
    layer2_outputs(250) <= not b;
    layer2_outputs(251) <= not b or a;
    layer2_outputs(252) <= not a;
    layer2_outputs(253) <= not a;
    layer2_outputs(254) <= not a;
    layer2_outputs(255) <= not a or b;
    layer2_outputs(256) <= b;
    layer2_outputs(257) <= not b or a;
    layer2_outputs(258) <= a;
    layer2_outputs(259) <= a xor b;
    layer2_outputs(260) <= not a or b;
    layer2_outputs(261) <= not (a xor b);
    layer2_outputs(262) <= not a;
    layer2_outputs(263) <= not (a and b);
    layer2_outputs(264) <= a and b;
    layer2_outputs(265) <= a;
    layer2_outputs(266) <= b;
    layer2_outputs(267) <= not b;
    layer2_outputs(268) <= not b;
    layer2_outputs(269) <= a;
    layer2_outputs(270) <= not b or a;
    layer2_outputs(271) <= not (a xor b);
    layer2_outputs(272) <= a xor b;
    layer2_outputs(273) <= b and not a;
    layer2_outputs(274) <= a or b;
    layer2_outputs(275) <= not (a xor b);
    layer2_outputs(276) <= a xor b;
    layer2_outputs(277) <= not a;
    layer2_outputs(278) <= not a;
    layer2_outputs(279) <= b;
    layer2_outputs(280) <= not a or b;
    layer2_outputs(281) <= not b;
    layer2_outputs(282) <= not b or a;
    layer2_outputs(283) <= a xor b;
    layer2_outputs(284) <= not a;
    layer2_outputs(285) <= not b;
    layer2_outputs(286) <= not (a xor b);
    layer2_outputs(287) <= not a;
    layer2_outputs(288) <= b;
    layer2_outputs(289) <= not b;
    layer2_outputs(290) <= b;
    layer2_outputs(291) <= not (a xor b);
    layer2_outputs(292) <= a;
    layer2_outputs(293) <= not b;
    layer2_outputs(294) <= a;
    layer2_outputs(295) <= not (a and b);
    layer2_outputs(296) <= b;
    layer2_outputs(297) <= not (a or b);
    layer2_outputs(298) <= not (a xor b);
    layer2_outputs(299) <= not b or a;
    layer2_outputs(300) <= a and b;
    layer2_outputs(301) <= not b;
    layer2_outputs(302) <= a and b;
    layer2_outputs(303) <= not (a or b);
    layer2_outputs(304) <= b and not a;
    layer2_outputs(305) <= not (a or b);
    layer2_outputs(306) <= not b;
    layer2_outputs(307) <= a and not b;
    layer2_outputs(308) <= a and b;
    layer2_outputs(309) <= a xor b;
    layer2_outputs(310) <= not b;
    layer2_outputs(311) <= a and not b;
    layer2_outputs(312) <= b and not a;
    layer2_outputs(313) <= b;
    layer2_outputs(314) <= a;
    layer2_outputs(315) <= not a;
    layer2_outputs(316) <= a;
    layer2_outputs(317) <= a;
    layer2_outputs(318) <= a and not b;
    layer2_outputs(319) <= b and not a;
    layer2_outputs(320) <= a and b;
    layer2_outputs(321) <= not b;
    layer2_outputs(322) <= a;
    layer2_outputs(323) <= a or b;
    layer2_outputs(324) <= a;
    layer2_outputs(325) <= a xor b;
    layer2_outputs(326) <= a and not b;
    layer2_outputs(327) <= b;
    layer2_outputs(328) <= a or b;
    layer2_outputs(329) <= a;
    layer2_outputs(330) <= b and not a;
    layer2_outputs(331) <= a and not b;
    layer2_outputs(332) <= a;
    layer2_outputs(333) <= a or b;
    layer2_outputs(334) <= not (a xor b);
    layer2_outputs(335) <= not b;
    layer2_outputs(336) <= not (a xor b);
    layer2_outputs(337) <= not b;
    layer2_outputs(338) <= not a;
    layer2_outputs(339) <= not (a or b);
    layer2_outputs(340) <= a and b;
    layer2_outputs(341) <= a and b;
    layer2_outputs(342) <= not a;
    layer2_outputs(343) <= a and b;
    layer2_outputs(344) <= a and b;
    layer2_outputs(345) <= not b or a;
    layer2_outputs(346) <= not (a or b);
    layer2_outputs(347) <= a;
    layer2_outputs(348) <= a xor b;
    layer2_outputs(349) <= not a;
    layer2_outputs(350) <= a and not b;
    layer2_outputs(351) <= a and not b;
    layer2_outputs(352) <= a or b;
    layer2_outputs(353) <= a and b;
    layer2_outputs(354) <= not (a or b);
    layer2_outputs(355) <= a xor b;
    layer2_outputs(356) <= a or b;
    layer2_outputs(357) <= not b;
    layer2_outputs(358) <= not b;
    layer2_outputs(359) <= not a;
    layer2_outputs(360) <= not (a or b);
    layer2_outputs(361) <= a;
    layer2_outputs(362) <= not (a and b);
    layer2_outputs(363) <= not a;
    layer2_outputs(364) <= a;
    layer2_outputs(365) <= not (a and b);
    layer2_outputs(366) <= a;
    layer2_outputs(367) <= a and not b;
    layer2_outputs(368) <= not a;
    layer2_outputs(369) <= not a;
    layer2_outputs(370) <= b;
    layer2_outputs(371) <= not a;
    layer2_outputs(372) <= not b or a;
    layer2_outputs(373) <= b;
    layer2_outputs(374) <= a or b;
    layer2_outputs(375) <= a and not b;
    layer2_outputs(376) <= not a;
    layer2_outputs(377) <= b;
    layer2_outputs(378) <= b and not a;
    layer2_outputs(379) <= not (a or b);
    layer2_outputs(380) <= 1'b1;
    layer2_outputs(381) <= a or b;
    layer2_outputs(382) <= not b;
    layer2_outputs(383) <= b and not a;
    layer2_outputs(384) <= not b or a;
    layer2_outputs(385) <= not a;
    layer2_outputs(386) <= a;
    layer2_outputs(387) <= not b or a;
    layer2_outputs(388) <= not b;
    layer2_outputs(389) <= a and b;
    layer2_outputs(390) <= not (a or b);
    layer2_outputs(391) <= 1'b1;
    layer2_outputs(392) <= a and not b;
    layer2_outputs(393) <= not (a and b);
    layer2_outputs(394) <= not b;
    layer2_outputs(395) <= not b;
    layer2_outputs(396) <= not b;
    layer2_outputs(397) <= b and not a;
    layer2_outputs(398) <= a and not b;
    layer2_outputs(399) <= 1'b1;
    layer2_outputs(400) <= b;
    layer2_outputs(401) <= not (a or b);
    layer2_outputs(402) <= a;
    layer2_outputs(403) <= b and not a;
    layer2_outputs(404) <= not b;
    layer2_outputs(405) <= not (a or b);
    layer2_outputs(406) <= not a;
    layer2_outputs(407) <= b and not a;
    layer2_outputs(408) <= a or b;
    layer2_outputs(409) <= a or b;
    layer2_outputs(410) <= not b;
    layer2_outputs(411) <= not (a or b);
    layer2_outputs(412) <= a or b;
    layer2_outputs(413) <= not b;
    layer2_outputs(414) <= not b;
    layer2_outputs(415) <= a;
    layer2_outputs(416) <= not a;
    layer2_outputs(417) <= a and not b;
    layer2_outputs(418) <= a and b;
    layer2_outputs(419) <= not (a or b);
    layer2_outputs(420) <= a and b;
    layer2_outputs(421) <= b and not a;
    layer2_outputs(422) <= not a;
    layer2_outputs(423) <= not a;
    layer2_outputs(424) <= b;
    layer2_outputs(425) <= b;
    layer2_outputs(426) <= not (a xor b);
    layer2_outputs(427) <= b;
    layer2_outputs(428) <= a;
    layer2_outputs(429) <= not b or a;
    layer2_outputs(430) <= not a;
    layer2_outputs(431) <= not (a and b);
    layer2_outputs(432) <= b;
    layer2_outputs(433) <= not a;
    layer2_outputs(434) <= not (a xor b);
    layer2_outputs(435) <= a and not b;
    layer2_outputs(436) <= not (a and b);
    layer2_outputs(437) <= not (a or b);
    layer2_outputs(438) <= not (a and b);
    layer2_outputs(439) <= not (a or b);
    layer2_outputs(440) <= b;
    layer2_outputs(441) <= b and not a;
    layer2_outputs(442) <= a and b;
    layer2_outputs(443) <= not (a xor b);
    layer2_outputs(444) <= not (a xor b);
    layer2_outputs(445) <= not (a and b);
    layer2_outputs(446) <= not (a xor b);
    layer2_outputs(447) <= not a;
    layer2_outputs(448) <= not (a or b);
    layer2_outputs(449) <= a;
    layer2_outputs(450) <= a and not b;
    layer2_outputs(451) <= not b;
    layer2_outputs(452) <= b;
    layer2_outputs(453) <= not (a and b);
    layer2_outputs(454) <= b;
    layer2_outputs(455) <= a;
    layer2_outputs(456) <= not a or b;
    layer2_outputs(457) <= a;
    layer2_outputs(458) <= b;
    layer2_outputs(459) <= b and not a;
    layer2_outputs(460) <= b and not a;
    layer2_outputs(461) <= a and b;
    layer2_outputs(462) <= not a or b;
    layer2_outputs(463) <= not b;
    layer2_outputs(464) <= a;
    layer2_outputs(465) <= a;
    layer2_outputs(466) <= b and not a;
    layer2_outputs(467) <= a and b;
    layer2_outputs(468) <= a and not b;
    layer2_outputs(469) <= not b or a;
    layer2_outputs(470) <= a;
    layer2_outputs(471) <= not (a or b);
    layer2_outputs(472) <= a or b;
    layer2_outputs(473) <= not b;
    layer2_outputs(474) <= a and b;
    layer2_outputs(475) <= b;
    layer2_outputs(476) <= not a;
    layer2_outputs(477) <= b;
    layer2_outputs(478) <= b;
    layer2_outputs(479) <= not b;
    layer2_outputs(480) <= a or b;
    layer2_outputs(481) <= b;
    layer2_outputs(482) <= a or b;
    layer2_outputs(483) <= not (a xor b);
    layer2_outputs(484) <= not (a and b);
    layer2_outputs(485) <= b;
    layer2_outputs(486) <= b;
    layer2_outputs(487) <= a;
    layer2_outputs(488) <= not (a and b);
    layer2_outputs(489) <= a and not b;
    layer2_outputs(490) <= b;
    layer2_outputs(491) <= not (a or b);
    layer2_outputs(492) <= not a or b;
    layer2_outputs(493) <= a and not b;
    layer2_outputs(494) <= not (a and b);
    layer2_outputs(495) <= a;
    layer2_outputs(496) <= not a;
    layer2_outputs(497) <= a or b;
    layer2_outputs(498) <= a;
    layer2_outputs(499) <= b;
    layer2_outputs(500) <= a and b;
    layer2_outputs(501) <= b and not a;
    layer2_outputs(502) <= b and not a;
    layer2_outputs(503) <= a or b;
    layer2_outputs(504) <= b and not a;
    layer2_outputs(505) <= a xor b;
    layer2_outputs(506) <= not b;
    layer2_outputs(507) <= not a or b;
    layer2_outputs(508) <= a and not b;
    layer2_outputs(509) <= not b or a;
    layer2_outputs(510) <= not b;
    layer2_outputs(511) <= not a or b;
    layer2_outputs(512) <= b;
    layer2_outputs(513) <= not (a xor b);
    layer2_outputs(514) <= not a or b;
    layer2_outputs(515) <= a;
    layer2_outputs(516) <= a and not b;
    layer2_outputs(517) <= not b;
    layer2_outputs(518) <= not b or a;
    layer2_outputs(519) <= a;
    layer2_outputs(520) <= not (a and b);
    layer2_outputs(521) <= b;
    layer2_outputs(522) <= a or b;
    layer2_outputs(523) <= not b;
    layer2_outputs(524) <= not (a xor b);
    layer2_outputs(525) <= not b;
    layer2_outputs(526) <= not (a or b);
    layer2_outputs(527) <= not a;
    layer2_outputs(528) <= not (a or b);
    layer2_outputs(529) <= a xor b;
    layer2_outputs(530) <= a;
    layer2_outputs(531) <= not (a and b);
    layer2_outputs(532) <= not a;
    layer2_outputs(533) <= not b;
    layer2_outputs(534) <= not a or b;
    layer2_outputs(535) <= not a or b;
    layer2_outputs(536) <= not b or a;
    layer2_outputs(537) <= not a;
    layer2_outputs(538) <= a and not b;
    layer2_outputs(539) <= a and not b;
    layer2_outputs(540) <= not b;
    layer2_outputs(541) <= not (a or b);
    layer2_outputs(542) <= b and not a;
    layer2_outputs(543) <= b and not a;
    layer2_outputs(544) <= b;
    layer2_outputs(545) <= a and not b;
    layer2_outputs(546) <= not a or b;
    layer2_outputs(547) <= not (a or b);
    layer2_outputs(548) <= a and not b;
    layer2_outputs(549) <= not b;
    layer2_outputs(550) <= not (a and b);
    layer2_outputs(551) <= not b;
    layer2_outputs(552) <= not a or b;
    layer2_outputs(553) <= a xor b;
    layer2_outputs(554) <= not (a or b);
    layer2_outputs(555) <= a;
    layer2_outputs(556) <= not (a or b);
    layer2_outputs(557) <= a or b;
    layer2_outputs(558) <= a or b;
    layer2_outputs(559) <= b;
    layer2_outputs(560) <= a xor b;
    layer2_outputs(561) <= not b;
    layer2_outputs(562) <= a or b;
    layer2_outputs(563) <= not a or b;
    layer2_outputs(564) <= a xor b;
    layer2_outputs(565) <= not b or a;
    layer2_outputs(566) <= b and not a;
    layer2_outputs(567) <= not a;
    layer2_outputs(568) <= not b;
    layer2_outputs(569) <= a or b;
    layer2_outputs(570) <= not b or a;
    layer2_outputs(571) <= not b;
    layer2_outputs(572) <= b and not a;
    layer2_outputs(573) <= a;
    layer2_outputs(574) <= not a or b;
    layer2_outputs(575) <= not (a or b);
    layer2_outputs(576) <= a and b;
    layer2_outputs(577) <= not b;
    layer2_outputs(578) <= not (a or b);
    layer2_outputs(579) <= a and b;
    layer2_outputs(580) <= not (a xor b);
    layer2_outputs(581) <= not a;
    layer2_outputs(582) <= a or b;
    layer2_outputs(583) <= not a;
    layer2_outputs(584) <= not (a or b);
    layer2_outputs(585) <= b;
    layer2_outputs(586) <= not (a xor b);
    layer2_outputs(587) <= b;
    layer2_outputs(588) <= not (a or b);
    layer2_outputs(589) <= not a;
    layer2_outputs(590) <= not b or a;
    layer2_outputs(591) <= not (a and b);
    layer2_outputs(592) <= a xor b;
    layer2_outputs(593) <= not a;
    layer2_outputs(594) <= a;
    layer2_outputs(595) <= not (a or b);
    layer2_outputs(596) <= not (a xor b);
    layer2_outputs(597) <= a and b;
    layer2_outputs(598) <= not (a or b);
    layer2_outputs(599) <= not b;
    layer2_outputs(600) <= a;
    layer2_outputs(601) <= not a or b;
    layer2_outputs(602) <= a;
    layer2_outputs(603) <= b;
    layer2_outputs(604) <= not (a and b);
    layer2_outputs(605) <= a and b;
    layer2_outputs(606) <= a xor b;
    layer2_outputs(607) <= b;
    layer2_outputs(608) <= b and not a;
    layer2_outputs(609) <= b and not a;
    layer2_outputs(610) <= not a or b;
    layer2_outputs(611) <= not (a and b);
    layer2_outputs(612) <= not a;
    layer2_outputs(613) <= b;
    layer2_outputs(614) <= not (a and b);
    layer2_outputs(615) <= not b;
    layer2_outputs(616) <= not b or a;
    layer2_outputs(617) <= b;
    layer2_outputs(618) <= a;
    layer2_outputs(619) <= not b or a;
    layer2_outputs(620) <= not (a xor b);
    layer2_outputs(621) <= not a;
    layer2_outputs(622) <= a;
    layer2_outputs(623) <= a and not b;
    layer2_outputs(624) <= a;
    layer2_outputs(625) <= not (a and b);
    layer2_outputs(626) <= not b;
    layer2_outputs(627) <= not (a xor b);
    layer2_outputs(628) <= not b;
    layer2_outputs(629) <= 1'b1;
    layer2_outputs(630) <= not a or b;
    layer2_outputs(631) <= not b or a;
    layer2_outputs(632) <= a and b;
    layer2_outputs(633) <= b;
    layer2_outputs(634) <= a and b;
    layer2_outputs(635) <= not a;
    layer2_outputs(636) <= a and not b;
    layer2_outputs(637) <= not (a and b);
    layer2_outputs(638) <= a;
    layer2_outputs(639) <= not (a or b);
    layer2_outputs(640) <= a and not b;
    layer2_outputs(641) <= not b;
    layer2_outputs(642) <= not b;
    layer2_outputs(643) <= not b;
    layer2_outputs(644) <= a;
    layer2_outputs(645) <= a or b;
    layer2_outputs(646) <= not (a and b);
    layer2_outputs(647) <= b and not a;
    layer2_outputs(648) <= a and not b;
    layer2_outputs(649) <= 1'b0;
    layer2_outputs(650) <= a and not b;
    layer2_outputs(651) <= not (a or b);
    layer2_outputs(652) <= b;
    layer2_outputs(653) <= b;
    layer2_outputs(654) <= b;
    layer2_outputs(655) <= b and not a;
    layer2_outputs(656) <= b and not a;
    layer2_outputs(657) <= not a;
    layer2_outputs(658) <= b;
    layer2_outputs(659) <= not a;
    layer2_outputs(660) <= a;
    layer2_outputs(661) <= not b;
    layer2_outputs(662) <= 1'b1;
    layer2_outputs(663) <= not a;
    layer2_outputs(664) <= not b;
    layer2_outputs(665) <= not (a xor b);
    layer2_outputs(666) <= not a;
    layer2_outputs(667) <= a or b;
    layer2_outputs(668) <= not b;
    layer2_outputs(669) <= not (a xor b);
    layer2_outputs(670) <= a and b;
    layer2_outputs(671) <= not (a xor b);
    layer2_outputs(672) <= not a;
    layer2_outputs(673) <= not b or a;
    layer2_outputs(674) <= a and b;
    layer2_outputs(675) <= a;
    layer2_outputs(676) <= b;
    layer2_outputs(677) <= not b;
    layer2_outputs(678) <= a;
    layer2_outputs(679) <= b and not a;
    layer2_outputs(680) <= a;
    layer2_outputs(681) <= a;
    layer2_outputs(682) <= not a;
    layer2_outputs(683) <= not b;
    layer2_outputs(684) <= not a or b;
    layer2_outputs(685) <= a;
    layer2_outputs(686) <= not (a xor b);
    layer2_outputs(687) <= not a;
    layer2_outputs(688) <= b and not a;
    layer2_outputs(689) <= not (a or b);
    layer2_outputs(690) <= not a;
    layer2_outputs(691) <= not b;
    layer2_outputs(692) <= not b;
    layer2_outputs(693) <= b;
    layer2_outputs(694) <= not b or a;
    layer2_outputs(695) <= a and not b;
    layer2_outputs(696) <= b;
    layer2_outputs(697) <= a and not b;
    layer2_outputs(698) <= a xor b;
    layer2_outputs(699) <= a or b;
    layer2_outputs(700) <= not (a and b);
    layer2_outputs(701) <= not b;
    layer2_outputs(702) <= not (a and b);
    layer2_outputs(703) <= not b or a;
    layer2_outputs(704) <= 1'b1;
    layer2_outputs(705) <= not (a or b);
    layer2_outputs(706) <= b;
    layer2_outputs(707) <= not (a xor b);
    layer2_outputs(708) <= not a;
    layer2_outputs(709) <= b;
    layer2_outputs(710) <= not a or b;
    layer2_outputs(711) <= not a or b;
    layer2_outputs(712) <= a and not b;
    layer2_outputs(713) <= not (a xor b);
    layer2_outputs(714) <= not (a and b);
    layer2_outputs(715) <= b;
    layer2_outputs(716) <= a;
    layer2_outputs(717) <= b;
    layer2_outputs(718) <= not a;
    layer2_outputs(719) <= not a;
    layer2_outputs(720) <= not b;
    layer2_outputs(721) <= not b or a;
    layer2_outputs(722) <= not b;
    layer2_outputs(723) <= not a;
    layer2_outputs(724) <= not (a or b);
    layer2_outputs(725) <= a;
    layer2_outputs(726) <= b;
    layer2_outputs(727) <= a;
    layer2_outputs(728) <= a xor b;
    layer2_outputs(729) <= not a or b;
    layer2_outputs(730) <= not (a and b);
    layer2_outputs(731) <= a and b;
    layer2_outputs(732) <= a or b;
    layer2_outputs(733) <= not b;
    layer2_outputs(734) <= a and b;
    layer2_outputs(735) <= a and b;
    layer2_outputs(736) <= a xor b;
    layer2_outputs(737) <= not (a or b);
    layer2_outputs(738) <= not a or b;
    layer2_outputs(739) <= a or b;
    layer2_outputs(740) <= not (a xor b);
    layer2_outputs(741) <= not a or b;
    layer2_outputs(742) <= 1'b1;
    layer2_outputs(743) <= not (a and b);
    layer2_outputs(744) <= a or b;
    layer2_outputs(745) <= a or b;
    layer2_outputs(746) <= b;
    layer2_outputs(747) <= not b;
    layer2_outputs(748) <= not (a xor b);
    layer2_outputs(749) <= b;
    layer2_outputs(750) <= a and b;
    layer2_outputs(751) <= not a or b;
    layer2_outputs(752) <= not (a and b);
    layer2_outputs(753) <= not b or a;
    layer2_outputs(754) <= not (a xor b);
    layer2_outputs(755) <= not (a and b);
    layer2_outputs(756) <= not b;
    layer2_outputs(757) <= a and b;
    layer2_outputs(758) <= not a;
    layer2_outputs(759) <= not (a or b);
    layer2_outputs(760) <= b;
    layer2_outputs(761) <= b and not a;
    layer2_outputs(762) <= a xor b;
    layer2_outputs(763) <= not b;
    layer2_outputs(764) <= a;
    layer2_outputs(765) <= not a or b;
    layer2_outputs(766) <= b and not a;
    layer2_outputs(767) <= not b;
    layer2_outputs(768) <= not (a and b);
    layer2_outputs(769) <= a or b;
    layer2_outputs(770) <= b and not a;
    layer2_outputs(771) <= not (a or b);
    layer2_outputs(772) <= a;
    layer2_outputs(773) <= a;
    layer2_outputs(774) <= b and not a;
    layer2_outputs(775) <= a and not b;
    layer2_outputs(776) <= not a;
    layer2_outputs(777) <= not (a xor b);
    layer2_outputs(778) <= not a or b;
    layer2_outputs(779) <= a;
    layer2_outputs(780) <= a xor b;
    layer2_outputs(781) <= b and not a;
    layer2_outputs(782) <= a;
    layer2_outputs(783) <= not (a or b);
    layer2_outputs(784) <= a and not b;
    layer2_outputs(785) <= b and not a;
    layer2_outputs(786) <= b;
    layer2_outputs(787) <= not (a xor b);
    layer2_outputs(788) <= not (a or b);
    layer2_outputs(789) <= not a;
    layer2_outputs(790) <= not b or a;
    layer2_outputs(791) <= not (a and b);
    layer2_outputs(792) <= not (a or b);
    layer2_outputs(793) <= b;
    layer2_outputs(794) <= not (a and b);
    layer2_outputs(795) <= b;
    layer2_outputs(796) <= not (a xor b);
    layer2_outputs(797) <= a and not b;
    layer2_outputs(798) <= b;
    layer2_outputs(799) <= a and not b;
    layer2_outputs(800) <= not (a and b);
    layer2_outputs(801) <= not b or a;
    layer2_outputs(802) <= a;
    layer2_outputs(803) <= a;
    layer2_outputs(804) <= b;
    layer2_outputs(805) <= b and not a;
    layer2_outputs(806) <= a and not b;
    layer2_outputs(807) <= a or b;
    layer2_outputs(808) <= b and not a;
    layer2_outputs(809) <= a;
    layer2_outputs(810) <= not (a or b);
    layer2_outputs(811) <= not a or b;
    layer2_outputs(812) <= a or b;
    layer2_outputs(813) <= not b;
    layer2_outputs(814) <= not b;
    layer2_outputs(815) <= not a or b;
    layer2_outputs(816) <= a;
    layer2_outputs(817) <= a;
    layer2_outputs(818) <= a and not b;
    layer2_outputs(819) <= not b;
    layer2_outputs(820) <= a and not b;
    layer2_outputs(821) <= b;
    layer2_outputs(822) <= not a;
    layer2_outputs(823) <= not a or b;
    layer2_outputs(824) <= not b or a;
    layer2_outputs(825) <= b;
    layer2_outputs(826) <= b;
    layer2_outputs(827) <= b and not a;
    layer2_outputs(828) <= a;
    layer2_outputs(829) <= not b;
    layer2_outputs(830) <= a and not b;
    layer2_outputs(831) <= a and not b;
    layer2_outputs(832) <= a;
    layer2_outputs(833) <= not b;
    layer2_outputs(834) <= not b or a;
    layer2_outputs(835) <= not b;
    layer2_outputs(836) <= a or b;
    layer2_outputs(837) <= not b or a;
    layer2_outputs(838) <= not b or a;
    layer2_outputs(839) <= a and not b;
    layer2_outputs(840) <= a and b;
    layer2_outputs(841) <= not a;
    layer2_outputs(842) <= not b;
    layer2_outputs(843) <= not b or a;
    layer2_outputs(844) <= not b or a;
    layer2_outputs(845) <= not a or b;
    layer2_outputs(846) <= a and b;
    layer2_outputs(847) <= 1'b0;
    layer2_outputs(848) <= a and b;
    layer2_outputs(849) <= not a;
    layer2_outputs(850) <= not b;
    layer2_outputs(851) <= not b;
    layer2_outputs(852) <= not a;
    layer2_outputs(853) <= a;
    layer2_outputs(854) <= not b;
    layer2_outputs(855) <= a;
    layer2_outputs(856) <= a or b;
    layer2_outputs(857) <= not (a xor b);
    layer2_outputs(858) <= a xor b;
    layer2_outputs(859) <= b;
    layer2_outputs(860) <= a and not b;
    layer2_outputs(861) <= not a or b;
    layer2_outputs(862) <= a;
    layer2_outputs(863) <= a;
    layer2_outputs(864) <= b;
    layer2_outputs(865) <= not a;
    layer2_outputs(866) <= not b;
    layer2_outputs(867) <= a;
    layer2_outputs(868) <= a or b;
    layer2_outputs(869) <= not (a or b);
    layer2_outputs(870) <= b;
    layer2_outputs(871) <= not a;
    layer2_outputs(872) <= not a or b;
    layer2_outputs(873) <= not b or a;
    layer2_outputs(874) <= b and not a;
    layer2_outputs(875) <= a or b;
    layer2_outputs(876) <= a;
    layer2_outputs(877) <= not b;
    layer2_outputs(878) <= not (a and b);
    layer2_outputs(879) <= not b;
    layer2_outputs(880) <= not b;
    layer2_outputs(881) <= not b;
    layer2_outputs(882) <= a xor b;
    layer2_outputs(883) <= not (a and b);
    layer2_outputs(884) <= not b or a;
    layer2_outputs(885) <= not b or a;
    layer2_outputs(886) <= not a;
    layer2_outputs(887) <= a or b;
    layer2_outputs(888) <= a and b;
    layer2_outputs(889) <= not (a and b);
    layer2_outputs(890) <= not a;
    layer2_outputs(891) <= not a;
    layer2_outputs(892) <= not b;
    layer2_outputs(893) <= a and b;
    layer2_outputs(894) <= not (a or b);
    layer2_outputs(895) <= not b or a;
    layer2_outputs(896) <= a;
    layer2_outputs(897) <= not b or a;
    layer2_outputs(898) <= not (a and b);
    layer2_outputs(899) <= a and b;
    layer2_outputs(900) <= not b;
    layer2_outputs(901) <= b and not a;
    layer2_outputs(902) <= not b or a;
    layer2_outputs(903) <= a xor b;
    layer2_outputs(904) <= a and not b;
    layer2_outputs(905) <= b and not a;
    layer2_outputs(906) <= not (a or b);
    layer2_outputs(907) <= not b or a;
    layer2_outputs(908) <= b;
    layer2_outputs(909) <= b and not a;
    layer2_outputs(910) <= a or b;
    layer2_outputs(911) <= not b or a;
    layer2_outputs(912) <= b;
    layer2_outputs(913) <= b;
    layer2_outputs(914) <= not a;
    layer2_outputs(915) <= not a;
    layer2_outputs(916) <= not (a xor b);
    layer2_outputs(917) <= 1'b1;
    layer2_outputs(918) <= not a;
    layer2_outputs(919) <= not b or a;
    layer2_outputs(920) <= not (a or b);
    layer2_outputs(921) <= a and b;
    layer2_outputs(922) <= not b;
    layer2_outputs(923) <= not a;
    layer2_outputs(924) <= not b;
    layer2_outputs(925) <= a and b;
    layer2_outputs(926) <= 1'b1;
    layer2_outputs(927) <= b;
    layer2_outputs(928) <= a and not b;
    layer2_outputs(929) <= b;
    layer2_outputs(930) <= a;
    layer2_outputs(931) <= b and not a;
    layer2_outputs(932) <= not b or a;
    layer2_outputs(933) <= not (a and b);
    layer2_outputs(934) <= a and not b;
    layer2_outputs(935) <= not (a or b);
    layer2_outputs(936) <= not (a and b);
    layer2_outputs(937) <= not (a or b);
    layer2_outputs(938) <= b;
    layer2_outputs(939) <= a xor b;
    layer2_outputs(940) <= not a or b;
    layer2_outputs(941) <= a or b;
    layer2_outputs(942) <= not b;
    layer2_outputs(943) <= not a;
    layer2_outputs(944) <= a or b;
    layer2_outputs(945) <= not a;
    layer2_outputs(946) <= a or b;
    layer2_outputs(947) <= not a;
    layer2_outputs(948) <= b and not a;
    layer2_outputs(949) <= not b;
    layer2_outputs(950) <= not (a or b);
    layer2_outputs(951) <= a and b;
    layer2_outputs(952) <= not a;
    layer2_outputs(953) <= b;
    layer2_outputs(954) <= not a;
    layer2_outputs(955) <= not b;
    layer2_outputs(956) <= a and b;
    layer2_outputs(957) <= not b;
    layer2_outputs(958) <= not a;
    layer2_outputs(959) <= a and b;
    layer2_outputs(960) <= not b;
    layer2_outputs(961) <= not b;
    layer2_outputs(962) <= not a or b;
    layer2_outputs(963) <= not a;
    layer2_outputs(964) <= a and b;
    layer2_outputs(965) <= a and b;
    layer2_outputs(966) <= a;
    layer2_outputs(967) <= a or b;
    layer2_outputs(968) <= b and not a;
    layer2_outputs(969) <= not (a or b);
    layer2_outputs(970) <= not b;
    layer2_outputs(971) <= not b;
    layer2_outputs(972) <= not b;
    layer2_outputs(973) <= not b or a;
    layer2_outputs(974) <= not (a or b);
    layer2_outputs(975) <= not b;
    layer2_outputs(976) <= 1'b1;
    layer2_outputs(977) <= a or b;
    layer2_outputs(978) <= not b;
    layer2_outputs(979) <= a;
    layer2_outputs(980) <= a and not b;
    layer2_outputs(981) <= a and b;
    layer2_outputs(982) <= not (a or b);
    layer2_outputs(983) <= a and b;
    layer2_outputs(984) <= a and b;
    layer2_outputs(985) <= not (a xor b);
    layer2_outputs(986) <= a or b;
    layer2_outputs(987) <= not a or b;
    layer2_outputs(988) <= not a or b;
    layer2_outputs(989) <= a or b;
    layer2_outputs(990) <= b and not a;
    layer2_outputs(991) <= a;
    layer2_outputs(992) <= not (a or b);
    layer2_outputs(993) <= b and not a;
    layer2_outputs(994) <= a and not b;
    layer2_outputs(995) <= not a or b;
    layer2_outputs(996) <= 1'b1;
    layer2_outputs(997) <= not a;
    layer2_outputs(998) <= not (a xor b);
    layer2_outputs(999) <= not a or b;
    layer2_outputs(1000) <= not (a or b);
    layer2_outputs(1001) <= a and b;
    layer2_outputs(1002) <= a and not b;
    layer2_outputs(1003) <= 1'b1;
    layer2_outputs(1004) <= a xor b;
    layer2_outputs(1005) <= not a;
    layer2_outputs(1006) <= a;
    layer2_outputs(1007) <= not a;
    layer2_outputs(1008) <= not b or a;
    layer2_outputs(1009) <= 1'b1;
    layer2_outputs(1010) <= a;
    layer2_outputs(1011) <= b;
    layer2_outputs(1012) <= a xor b;
    layer2_outputs(1013) <= not a;
    layer2_outputs(1014) <= not (a or b);
    layer2_outputs(1015) <= not (a and b);
    layer2_outputs(1016) <= 1'b1;
    layer2_outputs(1017) <= not a or b;
    layer2_outputs(1018) <= a and b;
    layer2_outputs(1019) <= not a;
    layer2_outputs(1020) <= a or b;
    layer2_outputs(1021) <= not a or b;
    layer2_outputs(1022) <= not a;
    layer2_outputs(1023) <= b and not a;
    layer2_outputs(1024) <= a and not b;
    layer2_outputs(1025) <= b;
    layer2_outputs(1026) <= b;
    layer2_outputs(1027) <= a;
    layer2_outputs(1028) <= a;
    layer2_outputs(1029) <= not (a or b);
    layer2_outputs(1030) <= not b or a;
    layer2_outputs(1031) <= b;
    layer2_outputs(1032) <= a;
    layer2_outputs(1033) <= a and b;
    layer2_outputs(1034) <= not b or a;
    layer2_outputs(1035) <= not b;
    layer2_outputs(1036) <= b and not a;
    layer2_outputs(1037) <= not b;
    layer2_outputs(1038) <= not b;
    layer2_outputs(1039) <= not b;
    layer2_outputs(1040) <= a and not b;
    layer2_outputs(1041) <= a and b;
    layer2_outputs(1042) <= not a or b;
    layer2_outputs(1043) <= b;
    layer2_outputs(1044) <= not b;
    layer2_outputs(1045) <= not (a and b);
    layer2_outputs(1046) <= not b;
    layer2_outputs(1047) <= b and not a;
    layer2_outputs(1048) <= a xor b;
    layer2_outputs(1049) <= a;
    layer2_outputs(1050) <= not (a or b);
    layer2_outputs(1051) <= a or b;
    layer2_outputs(1052) <= not a;
    layer2_outputs(1053) <= not b or a;
    layer2_outputs(1054) <= b and not a;
    layer2_outputs(1055) <= not a;
    layer2_outputs(1056) <= a;
    layer2_outputs(1057) <= b;
    layer2_outputs(1058) <= not a or b;
    layer2_outputs(1059) <= b;
    layer2_outputs(1060) <= not b or a;
    layer2_outputs(1061) <= not (a or b);
    layer2_outputs(1062) <= not (a or b);
    layer2_outputs(1063) <= a and b;
    layer2_outputs(1064) <= a xor b;
    layer2_outputs(1065) <= b;
    layer2_outputs(1066) <= not a;
    layer2_outputs(1067) <= b and not a;
    layer2_outputs(1068) <= 1'b0;
    layer2_outputs(1069) <= not b;
    layer2_outputs(1070) <= a;
    layer2_outputs(1071) <= not a or b;
    layer2_outputs(1072) <= not (a or b);
    layer2_outputs(1073) <= a xor b;
    layer2_outputs(1074) <= not a;
    layer2_outputs(1075) <= a and not b;
    layer2_outputs(1076) <= not a;
    layer2_outputs(1077) <= not b;
    layer2_outputs(1078) <= not a or b;
    layer2_outputs(1079) <= not (a xor b);
    layer2_outputs(1080) <= not (a and b);
    layer2_outputs(1081) <= b;
    layer2_outputs(1082) <= not (a and b);
    layer2_outputs(1083) <= not a;
    layer2_outputs(1084) <= a or b;
    layer2_outputs(1085) <= not b or a;
    layer2_outputs(1086) <= a and b;
    layer2_outputs(1087) <= a and not b;
    layer2_outputs(1088) <= not a;
    layer2_outputs(1089) <= a and not b;
    layer2_outputs(1090) <= a;
    layer2_outputs(1091) <= a;
    layer2_outputs(1092) <= a or b;
    layer2_outputs(1093) <= not (a or b);
    layer2_outputs(1094) <= not b or a;
    layer2_outputs(1095) <= a and b;
    layer2_outputs(1096) <= a or b;
    layer2_outputs(1097) <= a or b;
    layer2_outputs(1098) <= not b or a;
    layer2_outputs(1099) <= not b;
    layer2_outputs(1100) <= not b;
    layer2_outputs(1101) <= b;
    layer2_outputs(1102) <= b;
    layer2_outputs(1103) <= a or b;
    layer2_outputs(1104) <= not (a and b);
    layer2_outputs(1105) <= not b or a;
    layer2_outputs(1106) <= a;
    layer2_outputs(1107) <= not (a and b);
    layer2_outputs(1108) <= not (a and b);
    layer2_outputs(1109) <= not b;
    layer2_outputs(1110) <= a;
    layer2_outputs(1111) <= a and b;
    layer2_outputs(1112) <= b;
    layer2_outputs(1113) <= not b;
    layer2_outputs(1114) <= b;
    layer2_outputs(1115) <= a and not b;
    layer2_outputs(1116) <= not (a and b);
    layer2_outputs(1117) <= not a;
    layer2_outputs(1118) <= a and b;
    layer2_outputs(1119) <= 1'b0;
    layer2_outputs(1120) <= b and not a;
    layer2_outputs(1121) <= not b or a;
    layer2_outputs(1122) <= a;
    layer2_outputs(1123) <= not (a or b);
    layer2_outputs(1124) <= not b;
    layer2_outputs(1125) <= a;
    layer2_outputs(1126) <= not b;
    layer2_outputs(1127) <= a xor b;
    layer2_outputs(1128) <= b;
    layer2_outputs(1129) <= a or b;
    layer2_outputs(1130) <= a and not b;
    layer2_outputs(1131) <= b;
    layer2_outputs(1132) <= not b or a;
    layer2_outputs(1133) <= a xor b;
    layer2_outputs(1134) <= not (a and b);
    layer2_outputs(1135) <= not b;
    layer2_outputs(1136) <= not a or b;
    layer2_outputs(1137) <= not a or b;
    layer2_outputs(1138) <= not b;
    layer2_outputs(1139) <= not b;
    layer2_outputs(1140) <= b and not a;
    layer2_outputs(1141) <= not a;
    layer2_outputs(1142) <= not a;
    layer2_outputs(1143) <= not a;
    layer2_outputs(1144) <= not a or b;
    layer2_outputs(1145) <= a xor b;
    layer2_outputs(1146) <= b;
    layer2_outputs(1147) <= b;
    layer2_outputs(1148) <= b;
    layer2_outputs(1149) <= not (a xor b);
    layer2_outputs(1150) <= a and not b;
    layer2_outputs(1151) <= a;
    layer2_outputs(1152) <= not b;
    layer2_outputs(1153) <= b;
    layer2_outputs(1154) <= b;
    layer2_outputs(1155) <= a and not b;
    layer2_outputs(1156) <= a;
    layer2_outputs(1157) <= b;
    layer2_outputs(1158) <= not (a or b);
    layer2_outputs(1159) <= a and b;
    layer2_outputs(1160) <= not a;
    layer2_outputs(1161) <= a and not b;
    layer2_outputs(1162) <= a or b;
    layer2_outputs(1163) <= a and not b;
    layer2_outputs(1164) <= not b or a;
    layer2_outputs(1165) <= a or b;
    layer2_outputs(1166) <= a;
    layer2_outputs(1167) <= not b or a;
    layer2_outputs(1168) <= a or b;
    layer2_outputs(1169) <= 1'b0;
    layer2_outputs(1170) <= a or b;
    layer2_outputs(1171) <= not a;
    layer2_outputs(1172) <= not a;
    layer2_outputs(1173) <= not a or b;
    layer2_outputs(1174) <= not (a and b);
    layer2_outputs(1175) <= not b;
    layer2_outputs(1176) <= not a or b;
    layer2_outputs(1177) <= b and not a;
    layer2_outputs(1178) <= b and not a;
    layer2_outputs(1179) <= a and b;
    layer2_outputs(1180) <= b;
    layer2_outputs(1181) <= not b or a;
    layer2_outputs(1182) <= a and not b;
    layer2_outputs(1183) <= not a;
    layer2_outputs(1184) <= a and b;
    layer2_outputs(1185) <= a;
    layer2_outputs(1186) <= not b;
    layer2_outputs(1187) <= b;
    layer2_outputs(1188) <= not b or a;
    layer2_outputs(1189) <= not b;
    layer2_outputs(1190) <= a xor b;
    layer2_outputs(1191) <= not b;
    layer2_outputs(1192) <= a and b;
    layer2_outputs(1193) <= b;
    layer2_outputs(1194) <= not b;
    layer2_outputs(1195) <= not (a or b);
    layer2_outputs(1196) <= not (a and b);
    layer2_outputs(1197) <= not (a or b);
    layer2_outputs(1198) <= not (a or b);
    layer2_outputs(1199) <= a and b;
    layer2_outputs(1200) <= 1'b1;
    layer2_outputs(1201) <= not (a and b);
    layer2_outputs(1202) <= not (a and b);
    layer2_outputs(1203) <= a;
    layer2_outputs(1204) <= b;
    layer2_outputs(1205) <= not b;
    layer2_outputs(1206) <= not b;
    layer2_outputs(1207) <= not (a and b);
    layer2_outputs(1208) <= not b;
    layer2_outputs(1209) <= not a or b;
    layer2_outputs(1210) <= a;
    layer2_outputs(1211) <= a;
    layer2_outputs(1212) <= a and b;
    layer2_outputs(1213) <= a;
    layer2_outputs(1214) <= a;
    layer2_outputs(1215) <= a or b;
    layer2_outputs(1216) <= not a;
    layer2_outputs(1217) <= not b;
    layer2_outputs(1218) <= not b or a;
    layer2_outputs(1219) <= b and not a;
    layer2_outputs(1220) <= not a;
    layer2_outputs(1221) <= not (a xor b);
    layer2_outputs(1222) <= b and not a;
    layer2_outputs(1223) <= not a or b;
    layer2_outputs(1224) <= not a or b;
    layer2_outputs(1225) <= b;
    layer2_outputs(1226) <= a and not b;
    layer2_outputs(1227) <= a and b;
    layer2_outputs(1228) <= not b;
    layer2_outputs(1229) <= not b or a;
    layer2_outputs(1230) <= not (a and b);
    layer2_outputs(1231) <= a and not b;
    layer2_outputs(1232) <= not b;
    layer2_outputs(1233) <= not a;
    layer2_outputs(1234) <= a;
    layer2_outputs(1235) <= not b;
    layer2_outputs(1236) <= a;
    layer2_outputs(1237) <= b;
    layer2_outputs(1238) <= a;
    layer2_outputs(1239) <= not (a or b);
    layer2_outputs(1240) <= b and not a;
    layer2_outputs(1241) <= not b or a;
    layer2_outputs(1242) <= not b or a;
    layer2_outputs(1243) <= a;
    layer2_outputs(1244) <= not b;
    layer2_outputs(1245) <= a and not b;
    layer2_outputs(1246) <= not b or a;
    layer2_outputs(1247) <= a;
    layer2_outputs(1248) <= not a or b;
    layer2_outputs(1249) <= a xor b;
    layer2_outputs(1250) <= a or b;
    layer2_outputs(1251) <= not a or b;
    layer2_outputs(1252) <= not b or a;
    layer2_outputs(1253) <= not b or a;
    layer2_outputs(1254) <= not b;
    layer2_outputs(1255) <= not a or b;
    layer2_outputs(1256) <= b and not a;
    layer2_outputs(1257) <= not a or b;
    layer2_outputs(1258) <= a;
    layer2_outputs(1259) <= a or b;
    layer2_outputs(1260) <= a;
    layer2_outputs(1261) <= a or b;
    layer2_outputs(1262) <= a xor b;
    layer2_outputs(1263) <= not b;
    layer2_outputs(1264) <= a;
    layer2_outputs(1265) <= b and not a;
    layer2_outputs(1266) <= b;
    layer2_outputs(1267) <= a;
    layer2_outputs(1268) <= not b;
    layer2_outputs(1269) <= b;
    layer2_outputs(1270) <= not b or a;
    layer2_outputs(1271) <= a;
    layer2_outputs(1272) <= not (a xor b);
    layer2_outputs(1273) <= b;
    layer2_outputs(1274) <= not a;
    layer2_outputs(1275) <= b;
    layer2_outputs(1276) <= a and b;
    layer2_outputs(1277) <= not b or a;
    layer2_outputs(1278) <= not (a and b);
    layer2_outputs(1279) <= a and not b;
    layer2_outputs(1280) <= not (a xor b);
    layer2_outputs(1281) <= not (a and b);
    layer2_outputs(1282) <= not b;
    layer2_outputs(1283) <= a or b;
    layer2_outputs(1284) <= a or b;
    layer2_outputs(1285) <= a xor b;
    layer2_outputs(1286) <= not b;
    layer2_outputs(1287) <= a or b;
    layer2_outputs(1288) <= not b;
    layer2_outputs(1289) <= not (a or b);
    layer2_outputs(1290) <= a or b;
    layer2_outputs(1291) <= a and b;
    layer2_outputs(1292) <= not b or a;
    layer2_outputs(1293) <= a and not b;
    layer2_outputs(1294) <= not (a or b);
    layer2_outputs(1295) <= 1'b1;
    layer2_outputs(1296) <= a;
    layer2_outputs(1297) <= not a or b;
    layer2_outputs(1298) <= not (a xor b);
    layer2_outputs(1299) <= not a or b;
    layer2_outputs(1300) <= a and not b;
    layer2_outputs(1301) <= not (a and b);
    layer2_outputs(1302) <= not (a and b);
    layer2_outputs(1303) <= not b or a;
    layer2_outputs(1304) <= not (a and b);
    layer2_outputs(1305) <= b and not a;
    layer2_outputs(1306) <= not (a or b);
    layer2_outputs(1307) <= not (a xor b);
    layer2_outputs(1308) <= not a or b;
    layer2_outputs(1309) <= b;
    layer2_outputs(1310) <= a and not b;
    layer2_outputs(1311) <= not (a or b);
    layer2_outputs(1312) <= not (a or b);
    layer2_outputs(1313) <= b;
    layer2_outputs(1314) <= not a or b;
    layer2_outputs(1315) <= not (a or b);
    layer2_outputs(1316) <= a or b;
    layer2_outputs(1317) <= a;
    layer2_outputs(1318) <= not (a or b);
    layer2_outputs(1319) <= not a;
    layer2_outputs(1320) <= not (a and b);
    layer2_outputs(1321) <= b and not a;
    layer2_outputs(1322) <= not (a or b);
    layer2_outputs(1323) <= not a;
    layer2_outputs(1324) <= not (a and b);
    layer2_outputs(1325) <= not (a xor b);
    layer2_outputs(1326) <= a xor b;
    layer2_outputs(1327) <= not b;
    layer2_outputs(1328) <= not b;
    layer2_outputs(1329) <= a and b;
    layer2_outputs(1330) <= not a;
    layer2_outputs(1331) <= not a or b;
    layer2_outputs(1332) <= a and not b;
    layer2_outputs(1333) <= not b;
    layer2_outputs(1334) <= a and not b;
    layer2_outputs(1335) <= b;
    layer2_outputs(1336) <= a;
    layer2_outputs(1337) <= not a or b;
    layer2_outputs(1338) <= not b;
    layer2_outputs(1339) <= not b or a;
    layer2_outputs(1340) <= not b or a;
    layer2_outputs(1341) <= b and not a;
    layer2_outputs(1342) <= b and not a;
    layer2_outputs(1343) <= b and not a;
    layer2_outputs(1344) <= not b;
    layer2_outputs(1345) <= not (a or b);
    layer2_outputs(1346) <= not (a xor b);
    layer2_outputs(1347) <= a and not b;
    layer2_outputs(1348) <= b and not a;
    layer2_outputs(1349) <= not b;
    layer2_outputs(1350) <= a or b;
    layer2_outputs(1351) <= not b or a;
    layer2_outputs(1352) <= not b or a;
    layer2_outputs(1353) <= not (a or b);
    layer2_outputs(1354) <= a xor b;
    layer2_outputs(1355) <= not (a or b);
    layer2_outputs(1356) <= a;
    layer2_outputs(1357) <= not b or a;
    layer2_outputs(1358) <= b;
    layer2_outputs(1359) <= not (a or b);
    layer2_outputs(1360) <= not (a or b);
    layer2_outputs(1361) <= not b or a;
    layer2_outputs(1362) <= b;
    layer2_outputs(1363) <= b;
    layer2_outputs(1364) <= not a;
    layer2_outputs(1365) <= a;
    layer2_outputs(1366) <= b;
    layer2_outputs(1367) <= not a;
    layer2_outputs(1368) <= a and not b;
    layer2_outputs(1369) <= not (a xor b);
    layer2_outputs(1370) <= not (a xor b);
    layer2_outputs(1371) <= not (a or b);
    layer2_outputs(1372) <= a xor b;
    layer2_outputs(1373) <= a xor b;
    layer2_outputs(1374) <= a or b;
    layer2_outputs(1375) <= not b;
    layer2_outputs(1376) <= not b;
    layer2_outputs(1377) <= b;
    layer2_outputs(1378) <= not (a xor b);
    layer2_outputs(1379) <= a;
    layer2_outputs(1380) <= a;
    layer2_outputs(1381) <= not (a and b);
    layer2_outputs(1382) <= a and b;
    layer2_outputs(1383) <= not (a xor b);
    layer2_outputs(1384) <= b;
    layer2_outputs(1385) <= not a or b;
    layer2_outputs(1386) <= b and not a;
    layer2_outputs(1387) <= a and b;
    layer2_outputs(1388) <= b;
    layer2_outputs(1389) <= not a or b;
    layer2_outputs(1390) <= b;
    layer2_outputs(1391) <= not a;
    layer2_outputs(1392) <= not (a or b);
    layer2_outputs(1393) <= not b;
    layer2_outputs(1394) <= a;
    layer2_outputs(1395) <= not (a or b);
    layer2_outputs(1396) <= a xor b;
    layer2_outputs(1397) <= a xor b;
    layer2_outputs(1398) <= not b;
    layer2_outputs(1399) <= a xor b;
    layer2_outputs(1400) <= b and not a;
    layer2_outputs(1401) <= not a;
    layer2_outputs(1402) <= not b;
    layer2_outputs(1403) <= not (a or b);
    layer2_outputs(1404) <= a and b;
    layer2_outputs(1405) <= not (a or b);
    layer2_outputs(1406) <= not b;
    layer2_outputs(1407) <= a xor b;
    layer2_outputs(1408) <= not b;
    layer2_outputs(1409) <= a xor b;
    layer2_outputs(1410) <= not a or b;
    layer2_outputs(1411) <= a;
    layer2_outputs(1412) <= not a;
    layer2_outputs(1413) <= a;
    layer2_outputs(1414) <= not (a and b);
    layer2_outputs(1415) <= not (a or b);
    layer2_outputs(1416) <= a xor b;
    layer2_outputs(1417) <= not a;
    layer2_outputs(1418) <= not b;
    layer2_outputs(1419) <= not b;
    layer2_outputs(1420) <= not b;
    layer2_outputs(1421) <= b;
    layer2_outputs(1422) <= not b;
    layer2_outputs(1423) <= a or b;
    layer2_outputs(1424) <= a;
    layer2_outputs(1425) <= a;
    layer2_outputs(1426) <= a;
    layer2_outputs(1427) <= not a;
    layer2_outputs(1428) <= a;
    layer2_outputs(1429) <= not (a and b);
    layer2_outputs(1430) <= a;
    layer2_outputs(1431) <= not (a xor b);
    layer2_outputs(1432) <= a and not b;
    layer2_outputs(1433) <= not a;
    layer2_outputs(1434) <= b;
    layer2_outputs(1435) <= a and not b;
    layer2_outputs(1436) <= b and not a;
    layer2_outputs(1437) <= not a;
    layer2_outputs(1438) <= not a or b;
    layer2_outputs(1439) <= b;
    layer2_outputs(1440) <= not (a and b);
    layer2_outputs(1441) <= a xor b;
    layer2_outputs(1442) <= a;
    layer2_outputs(1443) <= a and not b;
    layer2_outputs(1444) <= a xor b;
    layer2_outputs(1445) <= not a or b;
    layer2_outputs(1446) <= not b;
    layer2_outputs(1447) <= not a;
    layer2_outputs(1448) <= b;
    layer2_outputs(1449) <= a;
    layer2_outputs(1450) <= a and b;
    layer2_outputs(1451) <= a or b;
    layer2_outputs(1452) <= a;
    layer2_outputs(1453) <= a;
    layer2_outputs(1454) <= a and not b;
    layer2_outputs(1455) <= not b;
    layer2_outputs(1456) <= not (a xor b);
    layer2_outputs(1457) <= not a;
    layer2_outputs(1458) <= not a;
    layer2_outputs(1459) <= not a;
    layer2_outputs(1460) <= not a;
    layer2_outputs(1461) <= a;
    layer2_outputs(1462) <= not a;
    layer2_outputs(1463) <= not (a or b);
    layer2_outputs(1464) <= not b;
    layer2_outputs(1465) <= b;
    layer2_outputs(1466) <= a and not b;
    layer2_outputs(1467) <= a xor b;
    layer2_outputs(1468) <= a or b;
    layer2_outputs(1469) <= a and b;
    layer2_outputs(1470) <= not a;
    layer2_outputs(1471) <= not b;
    layer2_outputs(1472) <= b and not a;
    layer2_outputs(1473) <= 1'b1;
    layer2_outputs(1474) <= not (a or b);
    layer2_outputs(1475) <= a;
    layer2_outputs(1476) <= not b;
    layer2_outputs(1477) <= not (a and b);
    layer2_outputs(1478) <= not a;
    layer2_outputs(1479) <= a or b;
    layer2_outputs(1480) <= b and not a;
    layer2_outputs(1481) <= not (a or b);
    layer2_outputs(1482) <= not a or b;
    layer2_outputs(1483) <= not a;
    layer2_outputs(1484) <= not a;
    layer2_outputs(1485) <= not (a or b);
    layer2_outputs(1486) <= a;
    layer2_outputs(1487) <= not (a and b);
    layer2_outputs(1488) <= b;
    layer2_outputs(1489) <= a and not b;
    layer2_outputs(1490) <= not (a or b);
    layer2_outputs(1491) <= not b;
    layer2_outputs(1492) <= b;
    layer2_outputs(1493) <= not (a or b);
    layer2_outputs(1494) <= a or b;
    layer2_outputs(1495) <= not b;
    layer2_outputs(1496) <= a;
    layer2_outputs(1497) <= not a;
    layer2_outputs(1498) <= not (a and b);
    layer2_outputs(1499) <= not (a or b);
    layer2_outputs(1500) <= not (a or b);
    layer2_outputs(1501) <= not b or a;
    layer2_outputs(1502) <= a and b;
    layer2_outputs(1503) <= a;
    layer2_outputs(1504) <= not b;
    layer2_outputs(1505) <= a and not b;
    layer2_outputs(1506) <= not (a and b);
    layer2_outputs(1507) <= a xor b;
    layer2_outputs(1508) <= b;
    layer2_outputs(1509) <= not (a or b);
    layer2_outputs(1510) <= a and b;
    layer2_outputs(1511) <= not b or a;
    layer2_outputs(1512) <= not (a xor b);
    layer2_outputs(1513) <= a and not b;
    layer2_outputs(1514) <= not b or a;
    layer2_outputs(1515) <= b;
    layer2_outputs(1516) <= a;
    layer2_outputs(1517) <= a and not b;
    layer2_outputs(1518) <= not a;
    layer2_outputs(1519) <= a and not b;
    layer2_outputs(1520) <= a;
    layer2_outputs(1521) <= b and not a;
    layer2_outputs(1522) <= not (a or b);
    layer2_outputs(1523) <= a or b;
    layer2_outputs(1524) <= not a;
    layer2_outputs(1525) <= not b or a;
    layer2_outputs(1526) <= b;
    layer2_outputs(1527) <= b and not a;
    layer2_outputs(1528) <= a;
    layer2_outputs(1529) <= not b or a;
    layer2_outputs(1530) <= not (a or b);
    layer2_outputs(1531) <= a and not b;
    layer2_outputs(1532) <= b;
    layer2_outputs(1533) <= b;
    layer2_outputs(1534) <= a and not b;
    layer2_outputs(1535) <= a;
    layer2_outputs(1536) <= a and b;
    layer2_outputs(1537) <= not a;
    layer2_outputs(1538) <= not (a xor b);
    layer2_outputs(1539) <= b and not a;
    layer2_outputs(1540) <= b;
    layer2_outputs(1541) <= not (a or b);
    layer2_outputs(1542) <= 1'b1;
    layer2_outputs(1543) <= a;
    layer2_outputs(1544) <= a xor b;
    layer2_outputs(1545) <= a and not b;
    layer2_outputs(1546) <= not a or b;
    layer2_outputs(1547) <= a and b;
    layer2_outputs(1548) <= not a;
    layer2_outputs(1549) <= not b;
    layer2_outputs(1550) <= not b or a;
    layer2_outputs(1551) <= not (a or b);
    layer2_outputs(1552) <= not (a or b);
    layer2_outputs(1553) <= a;
    layer2_outputs(1554) <= b and not a;
    layer2_outputs(1555) <= a and b;
    layer2_outputs(1556) <= not (a or b);
    layer2_outputs(1557) <= a;
    layer2_outputs(1558) <= not (a and b);
    layer2_outputs(1559) <= not a or b;
    layer2_outputs(1560) <= b;
    layer2_outputs(1561) <= not b or a;
    layer2_outputs(1562) <= b and not a;
    layer2_outputs(1563) <= a;
    layer2_outputs(1564) <= not b or a;
    layer2_outputs(1565) <= not (a xor b);
    layer2_outputs(1566) <= a and not b;
    layer2_outputs(1567) <= not a;
    layer2_outputs(1568) <= a;
    layer2_outputs(1569) <= a or b;
    layer2_outputs(1570) <= not (a xor b);
    layer2_outputs(1571) <= not a;
    layer2_outputs(1572) <= a xor b;
    layer2_outputs(1573) <= a or b;
    layer2_outputs(1574) <= a or b;
    layer2_outputs(1575) <= b;
    layer2_outputs(1576) <= b;
    layer2_outputs(1577) <= b and not a;
    layer2_outputs(1578) <= b and not a;
    layer2_outputs(1579) <= a and not b;
    layer2_outputs(1580) <= a and not b;
    layer2_outputs(1581) <= b;
    layer2_outputs(1582) <= not b;
    layer2_outputs(1583) <= b and not a;
    layer2_outputs(1584) <= a or b;
    layer2_outputs(1585) <= not b or a;
    layer2_outputs(1586) <= a;
    layer2_outputs(1587) <= not b;
    layer2_outputs(1588) <= not b or a;
    layer2_outputs(1589) <= not b;
    layer2_outputs(1590) <= not b;
    layer2_outputs(1591) <= b and not a;
    layer2_outputs(1592) <= a or b;
    layer2_outputs(1593) <= not b or a;
    layer2_outputs(1594) <= not a;
    layer2_outputs(1595) <= a and b;
    layer2_outputs(1596) <= not a;
    layer2_outputs(1597) <= a;
    layer2_outputs(1598) <= not b;
    layer2_outputs(1599) <= a or b;
    layer2_outputs(1600) <= not b;
    layer2_outputs(1601) <= not a;
    layer2_outputs(1602) <= 1'b1;
    layer2_outputs(1603) <= not b or a;
    layer2_outputs(1604) <= not a;
    layer2_outputs(1605) <= a and b;
    layer2_outputs(1606) <= not (a xor b);
    layer2_outputs(1607) <= a xor b;
    layer2_outputs(1608) <= b and not a;
    layer2_outputs(1609) <= b;
    layer2_outputs(1610) <= not a or b;
    layer2_outputs(1611) <= a xor b;
    layer2_outputs(1612) <= not (a xor b);
    layer2_outputs(1613) <= a;
    layer2_outputs(1614) <= a or b;
    layer2_outputs(1615) <= a or b;
    layer2_outputs(1616) <= not a or b;
    layer2_outputs(1617) <= a;
    layer2_outputs(1618) <= a xor b;
    layer2_outputs(1619) <= a;
    layer2_outputs(1620) <= not a;
    layer2_outputs(1621) <= not a or b;
    layer2_outputs(1622) <= a and b;
    layer2_outputs(1623) <= 1'b0;
    layer2_outputs(1624) <= b and not a;
    layer2_outputs(1625) <= not b;
    layer2_outputs(1626) <= b and not a;
    layer2_outputs(1627) <= not (a xor b);
    layer2_outputs(1628) <= b and not a;
    layer2_outputs(1629) <= b;
    layer2_outputs(1630) <= a and b;
    layer2_outputs(1631) <= not a or b;
    layer2_outputs(1632) <= not b;
    layer2_outputs(1633) <= a or b;
    layer2_outputs(1634) <= not a;
    layer2_outputs(1635) <= not a;
    layer2_outputs(1636) <= b;
    layer2_outputs(1637) <= not (a xor b);
    layer2_outputs(1638) <= a and b;
    layer2_outputs(1639) <= not a or b;
    layer2_outputs(1640) <= a;
    layer2_outputs(1641) <= b and not a;
    layer2_outputs(1642) <= b;
    layer2_outputs(1643) <= a xor b;
    layer2_outputs(1644) <= not (a or b);
    layer2_outputs(1645) <= not b;
    layer2_outputs(1646) <= not b;
    layer2_outputs(1647) <= a;
    layer2_outputs(1648) <= not (a or b);
    layer2_outputs(1649) <= a and not b;
    layer2_outputs(1650) <= not b;
    layer2_outputs(1651) <= a;
    layer2_outputs(1652) <= b;
    layer2_outputs(1653) <= not b or a;
    layer2_outputs(1654) <= not a;
    layer2_outputs(1655) <= a;
    layer2_outputs(1656) <= not a;
    layer2_outputs(1657) <= not a or b;
    layer2_outputs(1658) <= not b;
    layer2_outputs(1659) <= not a or b;
    layer2_outputs(1660) <= a or b;
    layer2_outputs(1661) <= not b;
    layer2_outputs(1662) <= a or b;
    layer2_outputs(1663) <= a or b;
    layer2_outputs(1664) <= not (a and b);
    layer2_outputs(1665) <= a and b;
    layer2_outputs(1666) <= b;
    layer2_outputs(1667) <= a and b;
    layer2_outputs(1668) <= not a;
    layer2_outputs(1669) <= not a;
    layer2_outputs(1670) <= not (a or b);
    layer2_outputs(1671) <= not (a or b);
    layer2_outputs(1672) <= not b or a;
    layer2_outputs(1673) <= a or b;
    layer2_outputs(1674) <= b;
    layer2_outputs(1675) <= not b or a;
    layer2_outputs(1676) <= b;
    layer2_outputs(1677) <= a;
    layer2_outputs(1678) <= not (a and b);
    layer2_outputs(1679) <= not a or b;
    layer2_outputs(1680) <= not b or a;
    layer2_outputs(1681) <= a;
    layer2_outputs(1682) <= b;
    layer2_outputs(1683) <= a and not b;
    layer2_outputs(1684) <= not (a and b);
    layer2_outputs(1685) <= a;
    layer2_outputs(1686) <= a or b;
    layer2_outputs(1687) <= a and b;
    layer2_outputs(1688) <= not a;
    layer2_outputs(1689) <= not (a or b);
    layer2_outputs(1690) <= a xor b;
    layer2_outputs(1691) <= not b;
    layer2_outputs(1692) <= a;
    layer2_outputs(1693) <= not a or b;
    layer2_outputs(1694) <= not b;
    layer2_outputs(1695) <= b;
    layer2_outputs(1696) <= not b;
    layer2_outputs(1697) <= not (a xor b);
    layer2_outputs(1698) <= a and not b;
    layer2_outputs(1699) <= not a;
    layer2_outputs(1700) <= not a;
    layer2_outputs(1701) <= a and b;
    layer2_outputs(1702) <= a and not b;
    layer2_outputs(1703) <= a or b;
    layer2_outputs(1704) <= not (a and b);
    layer2_outputs(1705) <= not (a xor b);
    layer2_outputs(1706) <= not b or a;
    layer2_outputs(1707) <= a and not b;
    layer2_outputs(1708) <= not a;
    layer2_outputs(1709) <= b;
    layer2_outputs(1710) <= a xor b;
    layer2_outputs(1711) <= not (a or b);
    layer2_outputs(1712) <= a;
    layer2_outputs(1713) <= a or b;
    layer2_outputs(1714) <= a;
    layer2_outputs(1715) <= not a;
    layer2_outputs(1716) <= not b;
    layer2_outputs(1717) <= not a;
    layer2_outputs(1718) <= a;
    layer2_outputs(1719) <= not b or a;
    layer2_outputs(1720) <= not (a and b);
    layer2_outputs(1721) <= not a or b;
    layer2_outputs(1722) <= not b;
    layer2_outputs(1723) <= 1'b0;
    layer2_outputs(1724) <= a and b;
    layer2_outputs(1725) <= not (a xor b);
    layer2_outputs(1726) <= not b;
    layer2_outputs(1727) <= b and not a;
    layer2_outputs(1728) <= not (a and b);
    layer2_outputs(1729) <= not a;
    layer2_outputs(1730) <= 1'b1;
    layer2_outputs(1731) <= not a or b;
    layer2_outputs(1732) <= a;
    layer2_outputs(1733) <= not (a or b);
    layer2_outputs(1734) <= a;
    layer2_outputs(1735) <= a;
    layer2_outputs(1736) <= not (a and b);
    layer2_outputs(1737) <= not a or b;
    layer2_outputs(1738) <= a or b;
    layer2_outputs(1739) <= not b or a;
    layer2_outputs(1740) <= not b;
    layer2_outputs(1741) <= not a;
    layer2_outputs(1742) <= not a;
    layer2_outputs(1743) <= not a;
    layer2_outputs(1744) <= a;
    layer2_outputs(1745) <= b;
    layer2_outputs(1746) <= not (a and b);
    layer2_outputs(1747) <= not a;
    layer2_outputs(1748) <= a xor b;
    layer2_outputs(1749) <= not a;
    layer2_outputs(1750) <= a;
    layer2_outputs(1751) <= not (a or b);
    layer2_outputs(1752) <= not a;
    layer2_outputs(1753) <= a or b;
    layer2_outputs(1754) <= a or b;
    layer2_outputs(1755) <= a or b;
    layer2_outputs(1756) <= not (a xor b);
    layer2_outputs(1757) <= not b;
    layer2_outputs(1758) <= 1'b0;
    layer2_outputs(1759) <= a;
    layer2_outputs(1760) <= a and b;
    layer2_outputs(1761) <= a and b;
    layer2_outputs(1762) <= b;
    layer2_outputs(1763) <= not b;
    layer2_outputs(1764) <= not a or b;
    layer2_outputs(1765) <= not b or a;
    layer2_outputs(1766) <= not b;
    layer2_outputs(1767) <= b;
    layer2_outputs(1768) <= not (a or b);
    layer2_outputs(1769) <= a and not b;
    layer2_outputs(1770) <= a;
    layer2_outputs(1771) <= b;
    layer2_outputs(1772) <= a xor b;
    layer2_outputs(1773) <= not a or b;
    layer2_outputs(1774) <= not b or a;
    layer2_outputs(1775) <= b and not a;
    layer2_outputs(1776) <= not a;
    layer2_outputs(1777) <= not b;
    layer2_outputs(1778) <= b;
    layer2_outputs(1779) <= not a or b;
    layer2_outputs(1780) <= a or b;
    layer2_outputs(1781) <= a or b;
    layer2_outputs(1782) <= not b or a;
    layer2_outputs(1783) <= b;
    layer2_outputs(1784) <= a xor b;
    layer2_outputs(1785) <= a or b;
    layer2_outputs(1786) <= a or b;
    layer2_outputs(1787) <= b and not a;
    layer2_outputs(1788) <= not a;
    layer2_outputs(1789) <= not (a and b);
    layer2_outputs(1790) <= b;
    layer2_outputs(1791) <= not b or a;
    layer2_outputs(1792) <= not (a or b);
    layer2_outputs(1793) <= a or b;
    layer2_outputs(1794) <= not b;
    layer2_outputs(1795) <= a and not b;
    layer2_outputs(1796) <= b and not a;
    layer2_outputs(1797) <= a;
    layer2_outputs(1798) <= a and b;
    layer2_outputs(1799) <= b and not a;
    layer2_outputs(1800) <= a and not b;
    layer2_outputs(1801) <= a;
    layer2_outputs(1802) <= a;
    layer2_outputs(1803) <= a;
    layer2_outputs(1804) <= a and b;
    layer2_outputs(1805) <= a or b;
    layer2_outputs(1806) <= not b;
    layer2_outputs(1807) <= not b or a;
    layer2_outputs(1808) <= a;
    layer2_outputs(1809) <= a or b;
    layer2_outputs(1810) <= not a;
    layer2_outputs(1811) <= not b;
    layer2_outputs(1812) <= not a or b;
    layer2_outputs(1813) <= a;
    layer2_outputs(1814) <= not (a and b);
    layer2_outputs(1815) <= not b;
    layer2_outputs(1816) <= b and not a;
    layer2_outputs(1817) <= a;
    layer2_outputs(1818) <= b;
    layer2_outputs(1819) <= not (a and b);
    layer2_outputs(1820) <= b;
    layer2_outputs(1821) <= a;
    layer2_outputs(1822) <= b and not a;
    layer2_outputs(1823) <= not (a or b);
    layer2_outputs(1824) <= a;
    layer2_outputs(1825) <= b;
    layer2_outputs(1826) <= not a;
    layer2_outputs(1827) <= b;
    layer2_outputs(1828) <= not (a or b);
    layer2_outputs(1829) <= b;
    layer2_outputs(1830) <= a and not b;
    layer2_outputs(1831) <= b;
    layer2_outputs(1832) <= b;
    layer2_outputs(1833) <= a or b;
    layer2_outputs(1834) <= b;
    layer2_outputs(1835) <= a or b;
    layer2_outputs(1836) <= not a or b;
    layer2_outputs(1837) <= a and not b;
    layer2_outputs(1838) <= a and b;
    layer2_outputs(1839) <= a or b;
    layer2_outputs(1840) <= not b or a;
    layer2_outputs(1841) <= not (a and b);
    layer2_outputs(1842) <= not b;
    layer2_outputs(1843) <= a;
    layer2_outputs(1844) <= b;
    layer2_outputs(1845) <= not (a or b);
    layer2_outputs(1846) <= a;
    layer2_outputs(1847) <= b;
    layer2_outputs(1848) <= b;
    layer2_outputs(1849) <= not b;
    layer2_outputs(1850) <= b;
    layer2_outputs(1851) <= not (a or b);
    layer2_outputs(1852) <= not a or b;
    layer2_outputs(1853) <= not b or a;
    layer2_outputs(1854) <= b;
    layer2_outputs(1855) <= a xor b;
    layer2_outputs(1856) <= b;
    layer2_outputs(1857) <= not (a or b);
    layer2_outputs(1858) <= a;
    layer2_outputs(1859) <= a xor b;
    layer2_outputs(1860) <= a;
    layer2_outputs(1861) <= b and not a;
    layer2_outputs(1862) <= a and b;
    layer2_outputs(1863) <= not a;
    layer2_outputs(1864) <= not a or b;
    layer2_outputs(1865) <= a xor b;
    layer2_outputs(1866) <= not (a or b);
    layer2_outputs(1867) <= not (a xor b);
    layer2_outputs(1868) <= a;
    layer2_outputs(1869) <= b;
    layer2_outputs(1870) <= a;
    layer2_outputs(1871) <= b;
    layer2_outputs(1872) <= a;
    layer2_outputs(1873) <= not b;
    layer2_outputs(1874) <= a;
    layer2_outputs(1875) <= not a;
    layer2_outputs(1876) <= not (a or b);
    layer2_outputs(1877) <= not a or b;
    layer2_outputs(1878) <= not a;
    layer2_outputs(1879) <= a or b;
    layer2_outputs(1880) <= b and not a;
    layer2_outputs(1881) <= not b;
    layer2_outputs(1882) <= a or b;
    layer2_outputs(1883) <= not (a and b);
    layer2_outputs(1884) <= not a or b;
    layer2_outputs(1885) <= not (a or b);
    layer2_outputs(1886) <= not b or a;
    layer2_outputs(1887) <= not (a xor b);
    layer2_outputs(1888) <= b;
    layer2_outputs(1889) <= not b;
    layer2_outputs(1890) <= not (a xor b);
    layer2_outputs(1891) <= not a or b;
    layer2_outputs(1892) <= not a;
    layer2_outputs(1893) <= not a or b;
    layer2_outputs(1894) <= not a or b;
    layer2_outputs(1895) <= b;
    layer2_outputs(1896) <= not a;
    layer2_outputs(1897) <= not (a xor b);
    layer2_outputs(1898) <= b;
    layer2_outputs(1899) <= b;
    layer2_outputs(1900) <= not (a or b);
    layer2_outputs(1901) <= not (a and b);
    layer2_outputs(1902) <= b;
    layer2_outputs(1903) <= not (a or b);
    layer2_outputs(1904) <= b;
    layer2_outputs(1905) <= b;
    layer2_outputs(1906) <= not a;
    layer2_outputs(1907) <= a;
    layer2_outputs(1908) <= not (a or b);
    layer2_outputs(1909) <= not a;
    layer2_outputs(1910) <= not b;
    layer2_outputs(1911) <= a and not b;
    layer2_outputs(1912) <= a and not b;
    layer2_outputs(1913) <= not (a or b);
    layer2_outputs(1914) <= not a;
    layer2_outputs(1915) <= b and not a;
    layer2_outputs(1916) <= b and not a;
    layer2_outputs(1917) <= not a;
    layer2_outputs(1918) <= a xor b;
    layer2_outputs(1919) <= a;
    layer2_outputs(1920) <= a and b;
    layer2_outputs(1921) <= not a or b;
    layer2_outputs(1922) <= b and not a;
    layer2_outputs(1923) <= a and not b;
    layer2_outputs(1924) <= a and not b;
    layer2_outputs(1925) <= not (a xor b);
    layer2_outputs(1926) <= a and not b;
    layer2_outputs(1927) <= not b;
    layer2_outputs(1928) <= not b;
    layer2_outputs(1929) <= not b or a;
    layer2_outputs(1930) <= a and not b;
    layer2_outputs(1931) <= a and b;
    layer2_outputs(1932) <= b;
    layer2_outputs(1933) <= a xor b;
    layer2_outputs(1934) <= a and b;
    layer2_outputs(1935) <= b and not a;
    layer2_outputs(1936) <= a xor b;
    layer2_outputs(1937) <= not b;
    layer2_outputs(1938) <= a and not b;
    layer2_outputs(1939) <= not (a and b);
    layer2_outputs(1940) <= not a;
    layer2_outputs(1941) <= not b;
    layer2_outputs(1942) <= not (a or b);
    layer2_outputs(1943) <= a or b;
    layer2_outputs(1944) <= not (a and b);
    layer2_outputs(1945) <= a;
    layer2_outputs(1946) <= a;
    layer2_outputs(1947) <= not b;
    layer2_outputs(1948) <= not b;
    layer2_outputs(1949) <= a and not b;
    layer2_outputs(1950) <= b and not a;
    layer2_outputs(1951) <= a xor b;
    layer2_outputs(1952) <= not b;
    layer2_outputs(1953) <= not b or a;
    layer2_outputs(1954) <= a;
    layer2_outputs(1955) <= a and b;
    layer2_outputs(1956) <= not a or b;
    layer2_outputs(1957) <= not a or b;
    layer2_outputs(1958) <= not (a and b);
    layer2_outputs(1959) <= b;
    layer2_outputs(1960) <= a or b;
    layer2_outputs(1961) <= not b;
    layer2_outputs(1962) <= not b;
    layer2_outputs(1963) <= a and b;
    layer2_outputs(1964) <= not (a and b);
    layer2_outputs(1965) <= not (a and b);
    layer2_outputs(1966) <= a and b;
    layer2_outputs(1967) <= not (a and b);
    layer2_outputs(1968) <= a;
    layer2_outputs(1969) <= a and not b;
    layer2_outputs(1970) <= not (a and b);
    layer2_outputs(1971) <= a;
    layer2_outputs(1972) <= not b;
    layer2_outputs(1973) <= 1'b1;
    layer2_outputs(1974) <= a and b;
    layer2_outputs(1975) <= b and not a;
    layer2_outputs(1976) <= not (a and b);
    layer2_outputs(1977) <= not a;
    layer2_outputs(1978) <= not b or a;
    layer2_outputs(1979) <= not b;
    layer2_outputs(1980) <= not (a and b);
    layer2_outputs(1981) <= a and not b;
    layer2_outputs(1982) <= not a;
    layer2_outputs(1983) <= a and not b;
    layer2_outputs(1984) <= a or b;
    layer2_outputs(1985) <= not b;
    layer2_outputs(1986) <= not (a or b);
    layer2_outputs(1987) <= not (a or b);
    layer2_outputs(1988) <= b;
    layer2_outputs(1989) <= a;
    layer2_outputs(1990) <= a and b;
    layer2_outputs(1991) <= not b;
    layer2_outputs(1992) <= not (a and b);
    layer2_outputs(1993) <= b;
    layer2_outputs(1994) <= b;
    layer2_outputs(1995) <= not (a and b);
    layer2_outputs(1996) <= not (a xor b);
    layer2_outputs(1997) <= a xor b;
    layer2_outputs(1998) <= a or b;
    layer2_outputs(1999) <= not a or b;
    layer2_outputs(2000) <= not (a xor b);
    layer2_outputs(2001) <= b;
    layer2_outputs(2002) <= 1'b0;
    layer2_outputs(2003) <= not a;
    layer2_outputs(2004) <= a xor b;
    layer2_outputs(2005) <= not a;
    layer2_outputs(2006) <= a;
    layer2_outputs(2007) <= a xor b;
    layer2_outputs(2008) <= b;
    layer2_outputs(2009) <= a and not b;
    layer2_outputs(2010) <= not (a or b);
    layer2_outputs(2011) <= b;
    layer2_outputs(2012) <= not b or a;
    layer2_outputs(2013) <= b;
    layer2_outputs(2014) <= not b or a;
    layer2_outputs(2015) <= not a or b;
    layer2_outputs(2016) <= b;
    layer2_outputs(2017) <= a xor b;
    layer2_outputs(2018) <= a xor b;
    layer2_outputs(2019) <= not b or a;
    layer2_outputs(2020) <= a or b;
    layer2_outputs(2021) <= not a or b;
    layer2_outputs(2022) <= b and not a;
    layer2_outputs(2023) <= not (a and b);
    layer2_outputs(2024) <= not (a xor b);
    layer2_outputs(2025) <= a;
    layer2_outputs(2026) <= not (a and b);
    layer2_outputs(2027) <= not a;
    layer2_outputs(2028) <= b and not a;
    layer2_outputs(2029) <= not b or a;
    layer2_outputs(2030) <= b;
    layer2_outputs(2031) <= a and b;
    layer2_outputs(2032) <= b;
    layer2_outputs(2033) <= not a;
    layer2_outputs(2034) <= not (a or b);
    layer2_outputs(2035) <= not (a xor b);
    layer2_outputs(2036) <= b and not a;
    layer2_outputs(2037) <= not b;
    layer2_outputs(2038) <= not b or a;
    layer2_outputs(2039) <= not b or a;
    layer2_outputs(2040) <= not (a and b);
    layer2_outputs(2041) <= b;
    layer2_outputs(2042) <= b;
    layer2_outputs(2043) <= a or b;
    layer2_outputs(2044) <= not a;
    layer2_outputs(2045) <= a and b;
    layer2_outputs(2046) <= not (a and b);
    layer2_outputs(2047) <= not (a or b);
    layer2_outputs(2048) <= b and not a;
    layer2_outputs(2049) <= not a;
    layer2_outputs(2050) <= b;
    layer2_outputs(2051) <= not (a xor b);
    layer2_outputs(2052) <= b and not a;
    layer2_outputs(2053) <= not (a and b);
    layer2_outputs(2054) <= a;
    layer2_outputs(2055) <= a and b;
    layer2_outputs(2056) <= b;
    layer2_outputs(2057) <= a and b;
    layer2_outputs(2058) <= not b;
    layer2_outputs(2059) <= not b;
    layer2_outputs(2060) <= a and b;
    layer2_outputs(2061) <= b and not a;
    layer2_outputs(2062) <= not a or b;
    layer2_outputs(2063) <= not a;
    layer2_outputs(2064) <= not b or a;
    layer2_outputs(2065) <= not a or b;
    layer2_outputs(2066) <= b;
    layer2_outputs(2067) <= not b or a;
    layer2_outputs(2068) <= a and not b;
    layer2_outputs(2069) <= not a;
    layer2_outputs(2070) <= not (a or b);
    layer2_outputs(2071) <= b;
    layer2_outputs(2072) <= b;
    layer2_outputs(2073) <= 1'b0;
    layer2_outputs(2074) <= a;
    layer2_outputs(2075) <= not b;
    layer2_outputs(2076) <= a xor b;
    layer2_outputs(2077) <= a and b;
    layer2_outputs(2078) <= 1'b0;
    layer2_outputs(2079) <= not (a or b);
    layer2_outputs(2080) <= not (a or b);
    layer2_outputs(2081) <= not a;
    layer2_outputs(2082) <= not a;
    layer2_outputs(2083) <= not b;
    layer2_outputs(2084) <= not a;
    layer2_outputs(2085) <= not b;
    layer2_outputs(2086) <= not a or b;
    layer2_outputs(2087) <= not b;
    layer2_outputs(2088) <= a and b;
    layer2_outputs(2089) <= b;
    layer2_outputs(2090) <= not (a or b);
    layer2_outputs(2091) <= a and b;
    layer2_outputs(2092) <= not a;
    layer2_outputs(2093) <= b;
    layer2_outputs(2094) <= not a;
    layer2_outputs(2095) <= not b;
    layer2_outputs(2096) <= not a or b;
    layer2_outputs(2097) <= b;
    layer2_outputs(2098) <= not a;
    layer2_outputs(2099) <= not b or a;
    layer2_outputs(2100) <= not b;
    layer2_outputs(2101) <= not a;
    layer2_outputs(2102) <= not (a or b);
    layer2_outputs(2103) <= a and b;
    layer2_outputs(2104) <= not a or b;
    layer2_outputs(2105) <= not b;
    layer2_outputs(2106) <= a and b;
    layer2_outputs(2107) <= not a or b;
    layer2_outputs(2108) <= not a;
    layer2_outputs(2109) <= not b;
    layer2_outputs(2110) <= not b or a;
    layer2_outputs(2111) <= b;
    layer2_outputs(2112) <= a;
    layer2_outputs(2113) <= b;
    layer2_outputs(2114) <= not (a xor b);
    layer2_outputs(2115) <= not b;
    layer2_outputs(2116) <= b;
    layer2_outputs(2117) <= a and b;
    layer2_outputs(2118) <= not b;
    layer2_outputs(2119) <= b;
    layer2_outputs(2120) <= not a;
    layer2_outputs(2121) <= not b;
    layer2_outputs(2122) <= not (a xor b);
    layer2_outputs(2123) <= not (a or b);
    layer2_outputs(2124) <= not (a or b);
    layer2_outputs(2125) <= not a;
    layer2_outputs(2126) <= a and not b;
    layer2_outputs(2127) <= not (a xor b);
    layer2_outputs(2128) <= not a;
    layer2_outputs(2129) <= a and b;
    layer2_outputs(2130) <= not a;
    layer2_outputs(2131) <= not b or a;
    layer2_outputs(2132) <= b and not a;
    layer2_outputs(2133) <= b;
    layer2_outputs(2134) <= a or b;
    layer2_outputs(2135) <= not (a and b);
    layer2_outputs(2136) <= a xor b;
    layer2_outputs(2137) <= a and not b;
    layer2_outputs(2138) <= a;
    layer2_outputs(2139) <= not (a and b);
    layer2_outputs(2140) <= a and not b;
    layer2_outputs(2141) <= not (a and b);
    layer2_outputs(2142) <= a or b;
    layer2_outputs(2143) <= a and not b;
    layer2_outputs(2144) <= not (a and b);
    layer2_outputs(2145) <= a and not b;
    layer2_outputs(2146) <= b;
    layer2_outputs(2147) <= a and b;
    layer2_outputs(2148) <= not a;
    layer2_outputs(2149) <= b;
    layer2_outputs(2150) <= b;
    layer2_outputs(2151) <= not b;
    layer2_outputs(2152) <= b;
    layer2_outputs(2153) <= not b;
    layer2_outputs(2154) <= not a;
    layer2_outputs(2155) <= a;
    layer2_outputs(2156) <= not (a or b);
    layer2_outputs(2157) <= not a;
    layer2_outputs(2158) <= a and not b;
    layer2_outputs(2159) <= not (a or b);
    layer2_outputs(2160) <= not a or b;
    layer2_outputs(2161) <= not a or b;
    layer2_outputs(2162) <= a and not b;
    layer2_outputs(2163) <= a;
    layer2_outputs(2164) <= not (a or b);
    layer2_outputs(2165) <= a or b;
    layer2_outputs(2166) <= not (a and b);
    layer2_outputs(2167) <= a and not b;
    layer2_outputs(2168) <= a;
    layer2_outputs(2169) <= not b;
    layer2_outputs(2170) <= not (a or b);
    layer2_outputs(2171) <= not b;
    layer2_outputs(2172) <= b and not a;
    layer2_outputs(2173) <= a and not b;
    layer2_outputs(2174) <= a and b;
    layer2_outputs(2175) <= not a;
    layer2_outputs(2176) <= b;
    layer2_outputs(2177) <= not b;
    layer2_outputs(2178) <= not a;
    layer2_outputs(2179) <= a xor b;
    layer2_outputs(2180) <= not b or a;
    layer2_outputs(2181) <= not (a and b);
    layer2_outputs(2182) <= a xor b;
    layer2_outputs(2183) <= not (a or b);
    layer2_outputs(2184) <= b;
    layer2_outputs(2185) <= not a or b;
    layer2_outputs(2186) <= not (a or b);
    layer2_outputs(2187) <= a;
    layer2_outputs(2188) <= not a;
    layer2_outputs(2189) <= not b or a;
    layer2_outputs(2190) <= a;
    layer2_outputs(2191) <= a and b;
    layer2_outputs(2192) <= b;
    layer2_outputs(2193) <= not (a xor b);
    layer2_outputs(2194) <= not b or a;
    layer2_outputs(2195) <= not a;
    layer2_outputs(2196) <= a and b;
    layer2_outputs(2197) <= not (a or b);
    layer2_outputs(2198) <= not (a xor b);
    layer2_outputs(2199) <= not (a or b);
    layer2_outputs(2200) <= not a or b;
    layer2_outputs(2201) <= a;
    layer2_outputs(2202) <= not a;
    layer2_outputs(2203) <= b;
    layer2_outputs(2204) <= a;
    layer2_outputs(2205) <= a xor b;
    layer2_outputs(2206) <= not (a and b);
    layer2_outputs(2207) <= b and not a;
    layer2_outputs(2208) <= not (a or b);
    layer2_outputs(2209) <= b;
    layer2_outputs(2210) <= a xor b;
    layer2_outputs(2211) <= not a or b;
    layer2_outputs(2212) <= not a or b;
    layer2_outputs(2213) <= a xor b;
    layer2_outputs(2214) <= not (a and b);
    layer2_outputs(2215) <= b and not a;
    layer2_outputs(2216) <= not a;
    layer2_outputs(2217) <= not (a xor b);
    layer2_outputs(2218) <= not b;
    layer2_outputs(2219) <= b;
    layer2_outputs(2220) <= not b;
    layer2_outputs(2221) <= not a;
    layer2_outputs(2222) <= a and b;
    layer2_outputs(2223) <= a;
    layer2_outputs(2224) <= b;
    layer2_outputs(2225) <= a and b;
    layer2_outputs(2226) <= a;
    layer2_outputs(2227) <= not a;
    layer2_outputs(2228) <= not (a or b);
    layer2_outputs(2229) <= not (a or b);
    layer2_outputs(2230) <= not b;
    layer2_outputs(2231) <= not (a and b);
    layer2_outputs(2232) <= not b or a;
    layer2_outputs(2233) <= b;
    layer2_outputs(2234) <= 1'b1;
    layer2_outputs(2235) <= not a;
    layer2_outputs(2236) <= b and not a;
    layer2_outputs(2237) <= a;
    layer2_outputs(2238) <= a and not b;
    layer2_outputs(2239) <= b;
    layer2_outputs(2240) <= not a;
    layer2_outputs(2241) <= not a;
    layer2_outputs(2242) <= not a;
    layer2_outputs(2243) <= not (a xor b);
    layer2_outputs(2244) <= b and not a;
    layer2_outputs(2245) <= a;
    layer2_outputs(2246) <= not a;
    layer2_outputs(2247) <= a xor b;
    layer2_outputs(2248) <= a;
    layer2_outputs(2249) <= b and not a;
    layer2_outputs(2250) <= a and not b;
    layer2_outputs(2251) <= not (a and b);
    layer2_outputs(2252) <= b;
    layer2_outputs(2253) <= b and not a;
    layer2_outputs(2254) <= not (a and b);
    layer2_outputs(2255) <= not a;
    layer2_outputs(2256) <= not a or b;
    layer2_outputs(2257) <= a and b;
    layer2_outputs(2258) <= not (a and b);
    layer2_outputs(2259) <= b and not a;
    layer2_outputs(2260) <= not a;
    layer2_outputs(2261) <= not (a and b);
    layer2_outputs(2262) <= not (a and b);
    layer2_outputs(2263) <= a and b;
    layer2_outputs(2264) <= not (a or b);
    layer2_outputs(2265) <= not (a or b);
    layer2_outputs(2266) <= a and b;
    layer2_outputs(2267) <= not a;
    layer2_outputs(2268) <= a;
    layer2_outputs(2269) <= not (a or b);
    layer2_outputs(2270) <= a or b;
    layer2_outputs(2271) <= a;
    layer2_outputs(2272) <= b;
    layer2_outputs(2273) <= not a;
    layer2_outputs(2274) <= not a or b;
    layer2_outputs(2275) <= not a or b;
    layer2_outputs(2276) <= not b;
    layer2_outputs(2277) <= b and not a;
    layer2_outputs(2278) <= not a;
    layer2_outputs(2279) <= a and b;
    layer2_outputs(2280) <= not b;
    layer2_outputs(2281) <= not b;
    layer2_outputs(2282) <= not (a or b);
    layer2_outputs(2283) <= a;
    layer2_outputs(2284) <= b and not a;
    layer2_outputs(2285) <= not b;
    layer2_outputs(2286) <= not a or b;
    layer2_outputs(2287) <= not b;
    layer2_outputs(2288) <= not b;
    layer2_outputs(2289) <= b;
    layer2_outputs(2290) <= a or b;
    layer2_outputs(2291) <= b and not a;
    layer2_outputs(2292) <= a and b;
    layer2_outputs(2293) <= a and b;
    layer2_outputs(2294) <= not b;
    layer2_outputs(2295) <= not b or a;
    layer2_outputs(2296) <= not b;
    layer2_outputs(2297) <= a and not b;
    layer2_outputs(2298) <= not (a xor b);
    layer2_outputs(2299) <= a;
    layer2_outputs(2300) <= a xor b;
    layer2_outputs(2301) <= b and not a;
    layer2_outputs(2302) <= a xor b;
    layer2_outputs(2303) <= not b or a;
    layer2_outputs(2304) <= not (a and b);
    layer2_outputs(2305) <= not b;
    layer2_outputs(2306) <= a;
    layer2_outputs(2307) <= not (a and b);
    layer2_outputs(2308) <= a;
    layer2_outputs(2309) <= not b;
    layer2_outputs(2310) <= not a;
    layer2_outputs(2311) <= b;
    layer2_outputs(2312) <= not b;
    layer2_outputs(2313) <= a;
    layer2_outputs(2314) <= not (a and b);
    layer2_outputs(2315) <= not (a or b);
    layer2_outputs(2316) <= not (a and b);
    layer2_outputs(2317) <= b and not a;
    layer2_outputs(2318) <= a or b;
    layer2_outputs(2319) <= a;
    layer2_outputs(2320) <= not a;
    layer2_outputs(2321) <= a;
    layer2_outputs(2322) <= a;
    layer2_outputs(2323) <= not (a xor b);
    layer2_outputs(2324) <= not a;
    layer2_outputs(2325) <= b and not a;
    layer2_outputs(2326) <= 1'b0;
    layer2_outputs(2327) <= b;
    layer2_outputs(2328) <= a;
    layer2_outputs(2329) <= a and not b;
    layer2_outputs(2330) <= b;
    layer2_outputs(2331) <= a;
    layer2_outputs(2332) <= not b;
    layer2_outputs(2333) <= a;
    layer2_outputs(2334) <= not (a or b);
    layer2_outputs(2335) <= not a;
    layer2_outputs(2336) <= a and not b;
    layer2_outputs(2337) <= 1'b0;
    layer2_outputs(2338) <= a;
    layer2_outputs(2339) <= a and not b;
    layer2_outputs(2340) <= not (a or b);
    layer2_outputs(2341) <= b and not a;
    layer2_outputs(2342) <= a xor b;
    layer2_outputs(2343) <= a;
    layer2_outputs(2344) <= not a or b;
    layer2_outputs(2345) <= a and b;
    layer2_outputs(2346) <= not b or a;
    layer2_outputs(2347) <= not (a or b);
    layer2_outputs(2348) <= a and not b;
    layer2_outputs(2349) <= not a;
    layer2_outputs(2350) <= not (a xor b);
    layer2_outputs(2351) <= not a or b;
    layer2_outputs(2352) <= not b or a;
    layer2_outputs(2353) <= b;
    layer2_outputs(2354) <= 1'b1;
    layer2_outputs(2355) <= b and not a;
    layer2_outputs(2356) <= not a;
    layer2_outputs(2357) <= 1'b1;
    layer2_outputs(2358) <= not a;
    layer2_outputs(2359) <= not (a and b);
    layer2_outputs(2360) <= not a or b;
    layer2_outputs(2361) <= not (a and b);
    layer2_outputs(2362) <= not b;
    layer2_outputs(2363) <= not b;
    layer2_outputs(2364) <= not a;
    layer2_outputs(2365) <= not b;
    layer2_outputs(2366) <= not a;
    layer2_outputs(2367) <= not b;
    layer2_outputs(2368) <= not (a and b);
    layer2_outputs(2369) <= not b or a;
    layer2_outputs(2370) <= b;
    layer2_outputs(2371) <= 1'b0;
    layer2_outputs(2372) <= not (a and b);
    layer2_outputs(2373) <= not b;
    layer2_outputs(2374) <= a and b;
    layer2_outputs(2375) <= not a;
    layer2_outputs(2376) <= b and not a;
    layer2_outputs(2377) <= not b or a;
    layer2_outputs(2378) <= not (a or b);
    layer2_outputs(2379) <= not (a xor b);
    layer2_outputs(2380) <= not (a or b);
    layer2_outputs(2381) <= not b or a;
    layer2_outputs(2382) <= not (a or b);
    layer2_outputs(2383) <= a and b;
    layer2_outputs(2384) <= not b;
    layer2_outputs(2385) <= not (a or b);
    layer2_outputs(2386) <= not (a or b);
    layer2_outputs(2387) <= not a;
    layer2_outputs(2388) <= b and not a;
    layer2_outputs(2389) <= not a or b;
    layer2_outputs(2390) <= b and not a;
    layer2_outputs(2391) <= b;
    layer2_outputs(2392) <= a;
    layer2_outputs(2393) <= b;
    layer2_outputs(2394) <= a or b;
    layer2_outputs(2395) <= not (a xor b);
    layer2_outputs(2396) <= not (a and b);
    layer2_outputs(2397) <= not b;
    layer2_outputs(2398) <= not b or a;
    layer2_outputs(2399) <= not (a or b);
    layer2_outputs(2400) <= b and not a;
    layer2_outputs(2401) <= not b;
    layer2_outputs(2402) <= a or b;
    layer2_outputs(2403) <= not (a xor b);
    layer2_outputs(2404) <= not a;
    layer2_outputs(2405) <= not b or a;
    layer2_outputs(2406) <= a or b;
    layer2_outputs(2407) <= a or b;
    layer2_outputs(2408) <= not (a or b);
    layer2_outputs(2409) <= not (a or b);
    layer2_outputs(2410) <= not (a or b);
    layer2_outputs(2411) <= not b or a;
    layer2_outputs(2412) <= not (a and b);
    layer2_outputs(2413) <= not a or b;
    layer2_outputs(2414) <= not b;
    layer2_outputs(2415) <= not (a or b);
    layer2_outputs(2416) <= not (a and b);
    layer2_outputs(2417) <= not b;
    layer2_outputs(2418) <= a;
    layer2_outputs(2419) <= not (a or b);
    layer2_outputs(2420) <= not a;
    layer2_outputs(2421) <= a or b;
    layer2_outputs(2422) <= not (a or b);
    layer2_outputs(2423) <= a and not b;
    layer2_outputs(2424) <= b;
    layer2_outputs(2425) <= not b;
    layer2_outputs(2426) <= not b;
    layer2_outputs(2427) <= b and not a;
    layer2_outputs(2428) <= a and not b;
    layer2_outputs(2429) <= b and not a;
    layer2_outputs(2430) <= b;
    layer2_outputs(2431) <= a;
    layer2_outputs(2432) <= not (a and b);
    layer2_outputs(2433) <= not a;
    layer2_outputs(2434) <= not b;
    layer2_outputs(2435) <= not (a and b);
    layer2_outputs(2436) <= not a or b;
    layer2_outputs(2437) <= a and not b;
    layer2_outputs(2438) <= a and not b;
    layer2_outputs(2439) <= a;
    layer2_outputs(2440) <= a and b;
    layer2_outputs(2441) <= a and not b;
    layer2_outputs(2442) <= b and not a;
    layer2_outputs(2443) <= a and not b;
    layer2_outputs(2444) <= a;
    layer2_outputs(2445) <= not a;
    layer2_outputs(2446) <= not a;
    layer2_outputs(2447) <= a and not b;
    layer2_outputs(2448) <= a or b;
    layer2_outputs(2449) <= not b;
    layer2_outputs(2450) <= b;
    layer2_outputs(2451) <= a xor b;
    layer2_outputs(2452) <= not a;
    layer2_outputs(2453) <= not a;
    layer2_outputs(2454) <= a;
    layer2_outputs(2455) <= not (a or b);
    layer2_outputs(2456) <= b;
    layer2_outputs(2457) <= not b or a;
    layer2_outputs(2458) <= not (a and b);
    layer2_outputs(2459) <= a and b;
    layer2_outputs(2460) <= a and not b;
    layer2_outputs(2461) <= b and not a;
    layer2_outputs(2462) <= a and not b;
    layer2_outputs(2463) <= not b or a;
    layer2_outputs(2464) <= not (a and b);
    layer2_outputs(2465) <= not b;
    layer2_outputs(2466) <= a or b;
    layer2_outputs(2467) <= not a or b;
    layer2_outputs(2468) <= b and not a;
    layer2_outputs(2469) <= not a or b;
    layer2_outputs(2470) <= a xor b;
    layer2_outputs(2471) <= not (a or b);
    layer2_outputs(2472) <= a;
    layer2_outputs(2473) <= not a;
    layer2_outputs(2474) <= a;
    layer2_outputs(2475) <= not a or b;
    layer2_outputs(2476) <= not a;
    layer2_outputs(2477) <= a and not b;
    layer2_outputs(2478) <= b;
    layer2_outputs(2479) <= not a;
    layer2_outputs(2480) <= b;
    layer2_outputs(2481) <= b;
    layer2_outputs(2482) <= a;
    layer2_outputs(2483) <= not a;
    layer2_outputs(2484) <= not a;
    layer2_outputs(2485) <= not a;
    layer2_outputs(2486) <= b and not a;
    layer2_outputs(2487) <= not (a or b);
    layer2_outputs(2488) <= not a or b;
    layer2_outputs(2489) <= not (a and b);
    layer2_outputs(2490) <= not a or b;
    layer2_outputs(2491) <= a;
    layer2_outputs(2492) <= not (a or b);
    layer2_outputs(2493) <= a;
    layer2_outputs(2494) <= b;
    layer2_outputs(2495) <= not a or b;
    layer2_outputs(2496) <= b;
    layer2_outputs(2497) <= a and b;
    layer2_outputs(2498) <= not b;
    layer2_outputs(2499) <= b and not a;
    layer2_outputs(2500) <= a and not b;
    layer2_outputs(2501) <= not b or a;
    layer2_outputs(2502) <= 1'b0;
    layer2_outputs(2503) <= not (a and b);
    layer2_outputs(2504) <= not (a xor b);
    layer2_outputs(2505) <= b and not a;
    layer2_outputs(2506) <= not (a or b);
    layer2_outputs(2507) <= not (a and b);
    layer2_outputs(2508) <= not a or b;
    layer2_outputs(2509) <= not b;
    layer2_outputs(2510) <= b and not a;
    layer2_outputs(2511) <= not b or a;
    layer2_outputs(2512) <= b;
    layer2_outputs(2513) <= a;
    layer2_outputs(2514) <= a and b;
    layer2_outputs(2515) <= a and b;
    layer2_outputs(2516) <= not (a or b);
    layer2_outputs(2517) <= not b or a;
    layer2_outputs(2518) <= a xor b;
    layer2_outputs(2519) <= a xor b;
    layer2_outputs(2520) <= b and not a;
    layer2_outputs(2521) <= not a;
    layer2_outputs(2522) <= a;
    layer2_outputs(2523) <= not a;
    layer2_outputs(2524) <= a xor b;
    layer2_outputs(2525) <= b and not a;
    layer2_outputs(2526) <= not (a xor b);
    layer2_outputs(2527) <= not a or b;
    layer2_outputs(2528) <= not b;
    layer2_outputs(2529) <= a and not b;
    layer2_outputs(2530) <= not a;
    layer2_outputs(2531) <= not (a or b);
    layer2_outputs(2532) <= not b;
    layer2_outputs(2533) <= a and not b;
    layer2_outputs(2534) <= a or b;
    layer2_outputs(2535) <= a or b;
    layer2_outputs(2536) <= not (a or b);
    layer2_outputs(2537) <= not b;
    layer2_outputs(2538) <= not b;
    layer2_outputs(2539) <= b;
    layer2_outputs(2540) <= a;
    layer2_outputs(2541) <= not (a xor b);
    layer2_outputs(2542) <= a;
    layer2_outputs(2543) <= not b;
    layer2_outputs(2544) <= b and not a;
    layer2_outputs(2545) <= not b;
    layer2_outputs(2546) <= b and not a;
    layer2_outputs(2547) <= not a;
    layer2_outputs(2548) <= not b or a;
    layer2_outputs(2549) <= not (a and b);
    layer2_outputs(2550) <= not b;
    layer2_outputs(2551) <= not b;
    layer2_outputs(2552) <= not (a and b);
    layer2_outputs(2553) <= b;
    layer2_outputs(2554) <= a or b;
    layer2_outputs(2555) <= not a;
    layer2_outputs(2556) <= not a;
    layer2_outputs(2557) <= a xor b;
    layer2_outputs(2558) <= a and not b;
    layer2_outputs(2559) <= a and not b;
    outputs(0) <= a and b;
    outputs(1) <= not b or a;
    outputs(2) <= not (a and b);
    outputs(3) <= not a;
    outputs(4) <= not b;
    outputs(5) <= a;
    outputs(6) <= a and b;
    outputs(7) <= not b or a;
    outputs(8) <= not b;
    outputs(9) <= b and not a;
    outputs(10) <= not a;
    outputs(11) <= not b or a;
    outputs(12) <= b and not a;
    outputs(13) <= a and not b;
    outputs(14) <= not b;
    outputs(15) <= a;
    outputs(16) <= not b or a;
    outputs(17) <= not (a or b);
    outputs(18) <= not (a or b);
    outputs(19) <= a;
    outputs(20) <= a;
    outputs(21) <= a and b;
    outputs(22) <= not b;
    outputs(23) <= b;
    outputs(24) <= not a;
    outputs(25) <= not a;
    outputs(26) <= a and not b;
    outputs(27) <= b;
    outputs(28) <= a and not b;
    outputs(29) <= a;
    outputs(30) <= not b;
    outputs(31) <= not b;
    outputs(32) <= a;
    outputs(33) <= not b;
    outputs(34) <= not a or b;
    outputs(35) <= a and not b;
    outputs(36) <= a;
    outputs(37) <= not a;
    outputs(38) <= a;
    outputs(39) <= b;
    outputs(40) <= not b;
    outputs(41) <= not b;
    outputs(42) <= a;
    outputs(43) <= not a;
    outputs(44) <= a and not b;
    outputs(45) <= not b or a;
    outputs(46) <= not b;
    outputs(47) <= a;
    outputs(48) <= a and b;
    outputs(49) <= b;
    outputs(50) <= not (a and b);
    outputs(51) <= not a;
    outputs(52) <= b;
    outputs(53) <= not b;
    outputs(54) <= b;
    outputs(55) <= not (a xor b);
    outputs(56) <= not a;
    outputs(57) <= not b;
    outputs(58) <= a xor b;
    outputs(59) <= b;
    outputs(60) <= not b or a;
    outputs(61) <= not (a or b);
    outputs(62) <= not a or b;
    outputs(63) <= not a;
    outputs(64) <= a and not b;
    outputs(65) <= a and not b;
    outputs(66) <= not a or b;
    outputs(67) <= not a;
    outputs(68) <= not a;
    outputs(69) <= a and b;
    outputs(70) <= a;
    outputs(71) <= not b;
    outputs(72) <= a;
    outputs(73) <= not b or a;
    outputs(74) <= not (a and b);
    outputs(75) <= b;
    outputs(76) <= a;
    outputs(77) <= b;
    outputs(78) <= not (a or b);
    outputs(79) <= a;
    outputs(80) <= a;
    outputs(81) <= a and b;
    outputs(82) <= not b;
    outputs(83) <= b;
    outputs(84) <= a and not b;
    outputs(85) <= a xor b;
    outputs(86) <= not b;
    outputs(87) <= not a;
    outputs(88) <= not b;
    outputs(89) <= b and not a;
    outputs(90) <= a;
    outputs(91) <= not (a and b);
    outputs(92) <= not a;
    outputs(93) <= b;
    outputs(94) <= a and b;
    outputs(95) <= not (a or b);
    outputs(96) <= b;
    outputs(97) <= not (a and b);
    outputs(98) <= not a or b;
    outputs(99) <= not a or b;
    outputs(100) <= a xor b;
    outputs(101) <= not a;
    outputs(102) <= a and not b;
    outputs(103) <= not (a or b);
    outputs(104) <= not (a and b);
    outputs(105) <= b;
    outputs(106) <= b and not a;
    outputs(107) <= a and not b;
    outputs(108) <= not b or a;
    outputs(109) <= a and not b;
    outputs(110) <= a or b;
    outputs(111) <= a xor b;
    outputs(112) <= not (a or b);
    outputs(113) <= a and not b;
    outputs(114) <= a;
    outputs(115) <= a and not b;
    outputs(116) <= not (a or b);
    outputs(117) <= not a;
    outputs(118) <= not (a and b);
    outputs(119) <= b;
    outputs(120) <= a or b;
    outputs(121) <= not b or a;
    outputs(122) <= a and not b;
    outputs(123) <= a;
    outputs(124) <= not a;
    outputs(125) <= not (a or b);
    outputs(126) <= b;
    outputs(127) <= not a;
    outputs(128) <= not b;
    outputs(129) <= b;
    outputs(130) <= not (a or b);
    outputs(131) <= a or b;
    outputs(132) <= a;
    outputs(133) <= b and not a;
    outputs(134) <= not b;
    outputs(135) <= a;
    outputs(136) <= b and not a;
    outputs(137) <= not b;
    outputs(138) <= b and not a;
    outputs(139) <= b;
    outputs(140) <= a;
    outputs(141) <= b;
    outputs(142) <= not b;
    outputs(143) <= not a;
    outputs(144) <= b and not a;
    outputs(145) <= not (a and b);
    outputs(146) <= b;
    outputs(147) <= not a;
    outputs(148) <= not a or b;
    outputs(149) <= not b;
    outputs(150) <= a or b;
    outputs(151) <= not (a and b);
    outputs(152) <= a and not b;
    outputs(153) <= not b;
    outputs(154) <= not (a xor b);
    outputs(155) <= not (a xor b);
    outputs(156) <= a;
    outputs(157) <= not b or a;
    outputs(158) <= not b or a;
    outputs(159) <= not a;
    outputs(160) <= a xor b;
    outputs(161) <= a;
    outputs(162) <= not b;
    outputs(163) <= not a;
    outputs(164) <= b;
    outputs(165) <= b;
    outputs(166) <= a;
    outputs(167) <= not (a xor b);
    outputs(168) <= b and not a;
    outputs(169) <= not b;
    outputs(170) <= a;
    outputs(171) <= a;
    outputs(172) <= not b;
    outputs(173) <= not b;
    outputs(174) <= a xor b;
    outputs(175) <= a;
    outputs(176) <= b and not a;
    outputs(177) <= a;
    outputs(178) <= a and not b;
    outputs(179) <= a xor b;
    outputs(180) <= a and not b;
    outputs(181) <= a or b;
    outputs(182) <= a;
    outputs(183) <= b;
    outputs(184) <= a;
    outputs(185) <= not a;
    outputs(186) <= not (a xor b);
    outputs(187) <= a;
    outputs(188) <= not (a or b);
    outputs(189) <= b;
    outputs(190) <= not a;
    outputs(191) <= not a or b;
    outputs(192) <= b and not a;
    outputs(193) <= b and not a;
    outputs(194) <= b;
    outputs(195) <= a and not b;
    outputs(196) <= not a;
    outputs(197) <= a and not b;
    outputs(198) <= not a;
    outputs(199) <= not a;
    outputs(200) <= not b;
    outputs(201) <= not a;
    outputs(202) <= not (a or b);
    outputs(203) <= a;
    outputs(204) <= a;
    outputs(205) <= a or b;
    outputs(206) <= not (a and b);
    outputs(207) <= a;
    outputs(208) <= b;
    outputs(209) <= not (a and b);
    outputs(210) <= not a or b;
    outputs(211) <= not (a or b);
    outputs(212) <= not b;
    outputs(213) <= not (a or b);
    outputs(214) <= not b or a;
    outputs(215) <= b and not a;
    outputs(216) <= not (a xor b);
    outputs(217) <= a and not b;
    outputs(218) <= b;
    outputs(219) <= b;
    outputs(220) <= not a or b;
    outputs(221) <= not (a and b);
    outputs(222) <= a xor b;
    outputs(223) <= not a;
    outputs(224) <= a;
    outputs(225) <= a;
    outputs(226) <= not a;
    outputs(227) <= not b;
    outputs(228) <= not b or a;
    outputs(229) <= a;
    outputs(230) <= b;
    outputs(231) <= b;
    outputs(232) <= a;
    outputs(233) <= a;
    outputs(234) <= b;
    outputs(235) <= not b;
    outputs(236) <= a;
    outputs(237) <= not b;
    outputs(238) <= not (a or b);
    outputs(239) <= a or b;
    outputs(240) <= a xor b;
    outputs(241) <= b and not a;
    outputs(242) <= a;
    outputs(243) <= not (a or b);
    outputs(244) <= not b;
    outputs(245) <= b;
    outputs(246) <= not a;
    outputs(247) <= a xor b;
    outputs(248) <= a;
    outputs(249) <= not a or b;
    outputs(250) <= a or b;
    outputs(251) <= b and not a;
    outputs(252) <= a;
    outputs(253) <= not (a xor b);
    outputs(254) <= a xor b;
    outputs(255) <= a;
    outputs(256) <= a and not b;
    outputs(257) <= not a;
    outputs(258) <= a and b;
    outputs(259) <= not (a xor b);
    outputs(260) <= a;
    outputs(261) <= b and not a;
    outputs(262) <= not (a or b);
    outputs(263) <= a and not b;
    outputs(264) <= a xor b;
    outputs(265) <= b and not a;
    outputs(266) <= not b;
    outputs(267) <= not a;
    outputs(268) <= a;
    outputs(269) <= a and not b;
    outputs(270) <= a and not b;
    outputs(271) <= b;
    outputs(272) <= b;
    outputs(273) <= a and b;
    outputs(274) <= a and not b;
    outputs(275) <= b;
    outputs(276) <= a and not b;
    outputs(277) <= a and b;
    outputs(278) <= a;
    outputs(279) <= b and not a;
    outputs(280) <= not (a or b);
    outputs(281) <= a and not b;
    outputs(282) <= not a;
    outputs(283) <= a;
    outputs(284) <= b and not a;
    outputs(285) <= a xor b;
    outputs(286) <= not (a or b);
    outputs(287) <= not (a or b);
    outputs(288) <= not (a or b);
    outputs(289) <= a and b;
    outputs(290) <= a and not b;
    outputs(291) <= a and b;
    outputs(292) <= not b or a;
    outputs(293) <= a and b;
    outputs(294) <= not b;
    outputs(295) <= not b;
    outputs(296) <= not b;
    outputs(297) <= b and not a;
    outputs(298) <= a and b;
    outputs(299) <= not (a or b);
    outputs(300) <= b;
    outputs(301) <= a and not b;
    outputs(302) <= a and b;
    outputs(303) <= a and b;
    outputs(304) <= a xor b;
    outputs(305) <= not (a or b);
    outputs(306) <= b and not a;
    outputs(307) <= not b;
    outputs(308) <= b;
    outputs(309) <= b;
    outputs(310) <= not (a or b);
    outputs(311) <= b and not a;
    outputs(312) <= b and not a;
    outputs(313) <= not a;
    outputs(314) <= not (a or b);
    outputs(315) <= a and not b;
    outputs(316) <= a;
    outputs(317) <= a and not b;
    outputs(318) <= a and b;
    outputs(319) <= a and not b;
    outputs(320) <= not (a or b);
    outputs(321) <= b;
    outputs(322) <= a and not b;
    outputs(323) <= a and b;
    outputs(324) <= a and b;
    outputs(325) <= b and not a;
    outputs(326) <= a xor b;
    outputs(327) <= not a or b;
    outputs(328) <= b and not a;
    outputs(329) <= a and b;
    outputs(330) <= a and b;
    outputs(331) <= not b;
    outputs(332) <= b and not a;
    outputs(333) <= a and not b;
    outputs(334) <= not b;
    outputs(335) <= not (a or b);
    outputs(336) <= not a;
    outputs(337) <= a and not b;
    outputs(338) <= not (a or b);
    outputs(339) <= a and not b;
    outputs(340) <= not b;
    outputs(341) <= a and not b;
    outputs(342) <= a and b;
    outputs(343) <= not (a or b);
    outputs(344) <= a and not b;
    outputs(345) <= not (a or b);
    outputs(346) <= b and not a;
    outputs(347) <= a and b;
    outputs(348) <= not b;
    outputs(349) <= not a;
    outputs(350) <= not a;
    outputs(351) <= a and not b;
    outputs(352) <= not a;
    outputs(353) <= a and b;
    outputs(354) <= not (a or b);
    outputs(355) <= b and not a;
    outputs(356) <= a and not b;
    outputs(357) <= a and b;
    outputs(358) <= not (a xor b);
    outputs(359) <= a and not b;
    outputs(360) <= b and not a;
    outputs(361) <= not (a or b);
    outputs(362) <= b and not a;
    outputs(363) <= b and not a;
    outputs(364) <= b and not a;
    outputs(365) <= b;
    outputs(366) <= a;
    outputs(367) <= not a;
    outputs(368) <= a and b;
    outputs(369) <= a and b;
    outputs(370) <= a and not b;
    outputs(371) <= not (a or b);
    outputs(372) <= a xor b;
    outputs(373) <= not a;
    outputs(374) <= a and not b;
    outputs(375) <= a;
    outputs(376) <= a and not b;
    outputs(377) <= not b or a;
    outputs(378) <= a and not b;
    outputs(379) <= a and not b;
    outputs(380) <= a and b;
    outputs(381) <= b;
    outputs(382) <= b and not a;
    outputs(383) <= b;
    outputs(384) <= a;
    outputs(385) <= a and not b;
    outputs(386) <= a;
    outputs(387) <= a and b;
    outputs(388) <= a and not b;
    outputs(389) <= not (a or b);
    outputs(390) <= not (a or b);
    outputs(391) <= a and not b;
    outputs(392) <= a and not b;
    outputs(393) <= b and not a;
    outputs(394) <= a xor b;
    outputs(395) <= a and not b;
    outputs(396) <= a and not b;
    outputs(397) <= b and not a;
    outputs(398) <= b and not a;
    outputs(399) <= a and not b;
    outputs(400) <= a;
    outputs(401) <= b and not a;
    outputs(402) <= not (a or b);
    outputs(403) <= a and b;
    outputs(404) <= not (a or b);
    outputs(405) <= a and b;
    outputs(406) <= b and not a;
    outputs(407) <= a and not b;
    outputs(408) <= a and not b;
    outputs(409) <= a and not b;
    outputs(410) <= a and b;
    outputs(411) <= not (a or b);
    outputs(412) <= a and b;
    outputs(413) <= b and not a;
    outputs(414) <= b and not a;
    outputs(415) <= not b;
    outputs(416) <= a and not b;
    outputs(417) <= not (a or b);
    outputs(418) <= b and not a;
    outputs(419) <= a xor b;
    outputs(420) <= b and not a;
    outputs(421) <= b and not a;
    outputs(422) <= b and not a;
    outputs(423) <= b and not a;
    outputs(424) <= not (a or b);
    outputs(425) <= a;
    outputs(426) <= a and b;
    outputs(427) <= a and b;
    outputs(428) <= a and b;
    outputs(429) <= b;
    outputs(430) <= a and not b;
    outputs(431) <= b and not a;
    outputs(432) <= a and b;
    outputs(433) <= a and b;
    outputs(434) <= not a;
    outputs(435) <= not (a or b);
    outputs(436) <= b and not a;
    outputs(437) <= b and not a;
    outputs(438) <= a and not b;
    outputs(439) <= a;
    outputs(440) <= a;
    outputs(441) <= b and not a;
    outputs(442) <= not b;
    outputs(443) <= b and not a;
    outputs(444) <= a;
    outputs(445) <= not (a or b);
    outputs(446) <= a;
    outputs(447) <= b and not a;
    outputs(448) <= b and not a;
    outputs(449) <= not (a or b);
    outputs(450) <= a and b;
    outputs(451) <= not (a or b);
    outputs(452) <= b;
    outputs(453) <= a and not b;
    outputs(454) <= not (a or b);
    outputs(455) <= b;
    outputs(456) <= a and not b;
    outputs(457) <= b;
    outputs(458) <= a and not b;
    outputs(459) <= b and not a;
    outputs(460) <= not a;
    outputs(461) <= not (a xor b);
    outputs(462) <= a;
    outputs(463) <= b and not a;
    outputs(464) <= not a;
    outputs(465) <= a and not b;
    outputs(466) <= a and not b;
    outputs(467) <= not (a or b);
    outputs(468) <= a;
    outputs(469) <= a and not b;
    outputs(470) <= b and not a;
    outputs(471) <= a and b;
    outputs(472) <= a and b;
    outputs(473) <= a xor b;
    outputs(474) <= b;
    outputs(475) <= a;
    outputs(476) <= b and not a;
    outputs(477) <= not b;
    outputs(478) <= not a;
    outputs(479) <= a and b;
    outputs(480) <= a and b;
    outputs(481) <= a and b;
    outputs(482) <= a and not b;
    outputs(483) <= a and not b;
    outputs(484) <= b;
    outputs(485) <= not b;
    outputs(486) <= b;
    outputs(487) <= a and not b;
    outputs(488) <= a and not b;
    outputs(489) <= a;
    outputs(490) <= a and not b;
    outputs(491) <= a;
    outputs(492) <= b and not a;
    outputs(493) <= a and not b;
    outputs(494) <= b and not a;
    outputs(495) <= a and b;
    outputs(496) <= a and b;
    outputs(497) <= a and b;
    outputs(498) <= a and b;
    outputs(499) <= b;
    outputs(500) <= not (a xor b);
    outputs(501) <= a and b;
    outputs(502) <= b and not a;
    outputs(503) <= not (a or b);
    outputs(504) <= not b;
    outputs(505) <= not b;
    outputs(506) <= not (a or b);
    outputs(507) <= a;
    outputs(508) <= not (a xor b);
    outputs(509) <= not a;
    outputs(510) <= not (a or b);
    outputs(511) <= not a;
    outputs(512) <= not a;
    outputs(513) <= not a;
    outputs(514) <= b;
    outputs(515) <= a and b;
    outputs(516) <= not a;
    outputs(517) <= not a;
    outputs(518) <= not (a xor b);
    outputs(519) <= not b or a;
    outputs(520) <= b and not a;
    outputs(521) <= not b;
    outputs(522) <= a or b;
    outputs(523) <= b;
    outputs(524) <= a;
    outputs(525) <= not b;
    outputs(526) <= b and not a;
    outputs(527) <= a;
    outputs(528) <= a;
    outputs(529) <= a or b;
    outputs(530) <= b;
    outputs(531) <= b;
    outputs(532) <= a or b;
    outputs(533) <= a;
    outputs(534) <= a and b;
    outputs(535) <= a and not b;
    outputs(536) <= not (a xor b);
    outputs(537) <= not a;
    outputs(538) <= b;
    outputs(539) <= not a;
    outputs(540) <= not b;
    outputs(541) <= a;
    outputs(542) <= a and not b;
    outputs(543) <= not (a or b);
    outputs(544) <= not (a and b);
    outputs(545) <= a;
    outputs(546) <= a or b;
    outputs(547) <= b;
    outputs(548) <= not (a or b);
    outputs(549) <= a or b;
    outputs(550) <= not (a and b);
    outputs(551) <= b and not a;
    outputs(552) <= not a;
    outputs(553) <= b and not a;
    outputs(554) <= a;
    outputs(555) <= not b;
    outputs(556) <= a and b;
    outputs(557) <= b and not a;
    outputs(558) <= b;
    outputs(559) <= a and b;
    outputs(560) <= not (a or b);
    outputs(561) <= not (a xor b);
    outputs(562) <= b;
    outputs(563) <= a or b;
    outputs(564) <= not (a or b);
    outputs(565) <= not a;
    outputs(566) <= a and b;
    outputs(567) <= a and b;
    outputs(568) <= not b;
    outputs(569) <= not (a or b);
    outputs(570) <= b;
    outputs(571) <= not (a xor b);
    outputs(572) <= not (a or b);
    outputs(573) <= not a;
    outputs(574) <= a or b;
    outputs(575) <= not a;
    outputs(576) <= a;
    outputs(577) <= a;
    outputs(578) <= a and b;
    outputs(579) <= a;
    outputs(580) <= not b;
    outputs(581) <= a and not b;
    outputs(582) <= b and not a;
    outputs(583) <= not (a xor b);
    outputs(584) <= not a;
    outputs(585) <= a xor b;
    outputs(586) <= not a or b;
    outputs(587) <= a or b;
    outputs(588) <= a;
    outputs(589) <= not (a and b);
    outputs(590) <= b;
    outputs(591) <= not a;
    outputs(592) <= a;
    outputs(593) <= not a;
    outputs(594) <= not a;
    outputs(595) <= b and not a;
    outputs(596) <= not b or a;
    outputs(597) <= a;
    outputs(598) <= not b;
    outputs(599) <= not b;
    outputs(600) <= not a;
    outputs(601) <= a and b;
    outputs(602) <= not b or a;
    outputs(603) <= not a;
    outputs(604) <= not b or a;
    outputs(605) <= not (a or b);
    outputs(606) <= not a or b;
    outputs(607) <= not (a xor b);
    outputs(608) <= a xor b;
    outputs(609) <= b and not a;
    outputs(610) <= not a;
    outputs(611) <= not (a or b);
    outputs(612) <= b;
    outputs(613) <= not (a or b);
    outputs(614) <= not b;
    outputs(615) <= not a;
    outputs(616) <= not (a or b);
    outputs(617) <= a or b;
    outputs(618) <= not (a and b);
    outputs(619) <= b;
    outputs(620) <= b and not a;
    outputs(621) <= a or b;
    outputs(622) <= not b or a;
    outputs(623) <= not a or b;
    outputs(624) <= not a;
    outputs(625) <= not (a or b);
    outputs(626) <= a;
    outputs(627) <= a;
    outputs(628) <= b;
    outputs(629) <= a;
    outputs(630) <= a and not b;
    outputs(631) <= a;
    outputs(632) <= not b;
    outputs(633) <= b;
    outputs(634) <= b;
    outputs(635) <= a;
    outputs(636) <= not (a xor b);
    outputs(637) <= not (a or b);
    outputs(638) <= not a;
    outputs(639) <= a and not b;
    outputs(640) <= a and not b;
    outputs(641) <= b and not a;
    outputs(642) <= a and b;
    outputs(643) <= b;
    outputs(644) <= not (a or b);
    outputs(645) <= not b;
    outputs(646) <= not b;
    outputs(647) <= a and not b;
    outputs(648) <= b;
    outputs(649) <= a and b;
    outputs(650) <= not b;
    outputs(651) <= a and not b;
    outputs(652) <= b;
    outputs(653) <= a and not b;
    outputs(654) <= b;
    outputs(655) <= not b;
    outputs(656) <= not b;
    outputs(657) <= not b;
    outputs(658) <= b;
    outputs(659) <= not (a or b);
    outputs(660) <= not b;
    outputs(661) <= not b;
    outputs(662) <= not b or a;
    outputs(663) <= not (a or b);
    outputs(664) <= b and not a;
    outputs(665) <= not b;
    outputs(666) <= b;
    outputs(667) <= a and not b;
    outputs(668) <= not (a xor b);
    outputs(669) <= a and not b;
    outputs(670) <= not b;
    outputs(671) <= a;
    outputs(672) <= not (a xor b);
    outputs(673) <= not (a xor b);
    outputs(674) <= b;
    outputs(675) <= not a;
    outputs(676) <= not b;
    outputs(677) <= not b;
    outputs(678) <= not b;
    outputs(679) <= b and not a;
    outputs(680) <= not b;
    outputs(681) <= b;
    outputs(682) <= not b or a;
    outputs(683) <= not a;
    outputs(684) <= b;
    outputs(685) <= a;
    outputs(686) <= not (a xor b);
    outputs(687) <= not b;
    outputs(688) <= b and not a;
    outputs(689) <= not a;
    outputs(690) <= not a;
    outputs(691) <= not a;
    outputs(692) <= b;
    outputs(693) <= a and not b;
    outputs(694) <= a and not b;
    outputs(695) <= b and not a;
    outputs(696) <= b;
    outputs(697) <= b;
    outputs(698) <= not a or b;
    outputs(699) <= a xor b;
    outputs(700) <= not b;
    outputs(701) <= not a;
    outputs(702) <= not b;
    outputs(703) <= not (a or b);
    outputs(704) <= a;
    outputs(705) <= b and not a;
    outputs(706) <= a and b;
    outputs(707) <= a;
    outputs(708) <= not a;
    outputs(709) <= not b;
    outputs(710) <= b;
    outputs(711) <= a;
    outputs(712) <= not (a or b);
    outputs(713) <= not (a xor b);
    outputs(714) <= a;
    outputs(715) <= a or b;
    outputs(716) <= a or b;
    outputs(717) <= not b or a;
    outputs(718) <= not b;
    outputs(719) <= a;
    outputs(720) <= not (a or b);
    outputs(721) <= a or b;
    outputs(722) <= not b;
    outputs(723) <= b and not a;
    outputs(724) <= b and not a;
    outputs(725) <= a and b;
    outputs(726) <= b;
    outputs(727) <= a or b;
    outputs(728) <= b and not a;
    outputs(729) <= not b;
    outputs(730) <= b;
    outputs(731) <= a;
    outputs(732) <= not a or b;
    outputs(733) <= a;
    outputs(734) <= not b or a;
    outputs(735) <= not b or a;
    outputs(736) <= not b or a;
    outputs(737) <= a xor b;
    outputs(738) <= a;
    outputs(739) <= b;
    outputs(740) <= b and not a;
    outputs(741) <= b;
    outputs(742) <= not (a or b);
    outputs(743) <= b;
    outputs(744) <= b;
    outputs(745) <= not (a xor b);
    outputs(746) <= not b or a;
    outputs(747) <= b;
    outputs(748) <= a and not b;
    outputs(749) <= b;
    outputs(750) <= not b;
    outputs(751) <= not b;
    outputs(752) <= not (a and b);
    outputs(753) <= b;
    outputs(754) <= not (a and b);
    outputs(755) <= a;
    outputs(756) <= a and b;
    outputs(757) <= not (a or b);
    outputs(758) <= a and b;
    outputs(759) <= a;
    outputs(760) <= not b or a;
    outputs(761) <= a;
    outputs(762) <= a and not b;
    outputs(763) <= not b or a;
    outputs(764) <= a;
    outputs(765) <= not a;
    outputs(766) <= not b;
    outputs(767) <= a and not b;
    outputs(768) <= a or b;
    outputs(769) <= a;
    outputs(770) <= a and not b;
    outputs(771) <= b;
    outputs(772) <= a and b;
    outputs(773) <= not b or a;
    outputs(774) <= a and b;
    outputs(775) <= not (a or b);
    outputs(776) <= not a;
    outputs(777) <= not a or b;
    outputs(778) <= b and not a;
    outputs(779) <= not (a and b);
    outputs(780) <= not (a or b);
    outputs(781) <= not (a or b);
    outputs(782) <= not b;
    outputs(783) <= not (a or b);
    outputs(784) <= a;
    outputs(785) <= a and b;
    outputs(786) <= b;
    outputs(787) <= not b;
    outputs(788) <= not a;
    outputs(789) <= not (a or b);
    outputs(790) <= a and b;
    outputs(791) <= a and not b;
    outputs(792) <= not a;
    outputs(793) <= not (a or b);
    outputs(794) <= b and not a;
    outputs(795) <= a and b;
    outputs(796) <= a;
    outputs(797) <= a xor b;
    outputs(798) <= not a or b;
    outputs(799) <= not (a or b);
    outputs(800) <= not b;
    outputs(801) <= a;
    outputs(802) <= a and not b;
    outputs(803) <= not b or a;
    outputs(804) <= not (a xor b);
    outputs(805) <= a and not b;
    outputs(806) <= b;
    outputs(807) <= not a;
    outputs(808) <= a xor b;
    outputs(809) <= not b or a;
    outputs(810) <= b and not a;
    outputs(811) <= not b;
    outputs(812) <= not (a and b);
    outputs(813) <= b and not a;
    outputs(814) <= not b;
    outputs(815) <= not b;
    outputs(816) <= not (a and b);
    outputs(817) <= b and not a;
    outputs(818) <= a;
    outputs(819) <= not (a or b);
    outputs(820) <= not a;
    outputs(821) <= not a;
    outputs(822) <= a;
    outputs(823) <= not b;
    outputs(824) <= not (a or b);
    outputs(825) <= a and b;
    outputs(826) <= not a;
    outputs(827) <= not (a and b);
    outputs(828) <= not (a and b);
    outputs(829) <= a and not b;
    outputs(830) <= b and not a;
    outputs(831) <= b and not a;
    outputs(832) <= b and not a;
    outputs(833) <= not b;
    outputs(834) <= not a or b;
    outputs(835) <= a;
    outputs(836) <= not b;
    outputs(837) <= a xor b;
    outputs(838) <= not (a xor b);
    outputs(839) <= b and not a;
    outputs(840) <= a and b;
    outputs(841) <= not a;
    outputs(842) <= not a;
    outputs(843) <= not a or b;
    outputs(844) <= a and b;
    outputs(845) <= b;
    outputs(846) <= a or b;
    outputs(847) <= b;
    outputs(848) <= not (a and b);
    outputs(849) <= b;
    outputs(850) <= a or b;
    outputs(851) <= b;
    outputs(852) <= not b;
    outputs(853) <= a xor b;
    outputs(854) <= not a;
    outputs(855) <= a and not b;
    outputs(856) <= not (a or b);
    outputs(857) <= not b;
    outputs(858) <= not b;
    outputs(859) <= a and not b;
    outputs(860) <= b;
    outputs(861) <= not a;
    outputs(862) <= a;
    outputs(863) <= a and not b;
    outputs(864) <= not (a xor b);
    outputs(865) <= a and b;
    outputs(866) <= a and not b;
    outputs(867) <= not (a xor b);
    outputs(868) <= not a;
    outputs(869) <= b;
    outputs(870) <= b;
    outputs(871) <= not (a or b);
    outputs(872) <= a;
    outputs(873) <= a and not b;
    outputs(874) <= a;
    outputs(875) <= b and not a;
    outputs(876) <= not a;
    outputs(877) <= a;
    outputs(878) <= not (a or b);
    outputs(879) <= not b or a;
    outputs(880) <= a xor b;
    outputs(881) <= not a;
    outputs(882) <= not (a and b);
    outputs(883) <= not a;
    outputs(884) <= b;
    outputs(885) <= not a;
    outputs(886) <= not a;
    outputs(887) <= a and b;
    outputs(888) <= not a;
    outputs(889) <= not b;
    outputs(890) <= a;
    outputs(891) <= not b;
    outputs(892) <= not a or b;
    outputs(893) <= a and b;
    outputs(894) <= not a or b;
    outputs(895) <= b;
    outputs(896) <= b;
    outputs(897) <= a and not b;
    outputs(898) <= not a;
    outputs(899) <= not a or b;
    outputs(900) <= not (a xor b);
    outputs(901) <= not b;
    outputs(902) <= a or b;
    outputs(903) <= a;
    outputs(904) <= b;
    outputs(905) <= a and b;
    outputs(906) <= a or b;
    outputs(907) <= not a;
    outputs(908) <= b and not a;
    outputs(909) <= a and b;
    outputs(910) <= not b or a;
    outputs(911) <= not a;
    outputs(912) <= not (a xor b);
    outputs(913) <= a or b;
    outputs(914) <= not (a or b);
    outputs(915) <= a or b;
    outputs(916) <= a and not b;
    outputs(917) <= a and not b;
    outputs(918) <= b;
    outputs(919) <= not (a or b);
    outputs(920) <= not b or a;
    outputs(921) <= not a or b;
    outputs(922) <= a;
    outputs(923) <= a;
    outputs(924) <= not a;
    outputs(925) <= a and not b;
    outputs(926) <= a;
    outputs(927) <= b;
    outputs(928) <= a and not b;
    outputs(929) <= a xor b;
    outputs(930) <= b and not a;
    outputs(931) <= b and not a;
    outputs(932) <= not (a xor b);
    outputs(933) <= b;
    outputs(934) <= not a;
    outputs(935) <= a and b;
    outputs(936) <= b;
    outputs(937) <= not b;
    outputs(938) <= not b;
    outputs(939) <= a;
    outputs(940) <= a;
    outputs(941) <= b and not a;
    outputs(942) <= not (a or b);
    outputs(943) <= b;
    outputs(944) <= a;
    outputs(945) <= b;
    outputs(946) <= not (a xor b);
    outputs(947) <= a and not b;
    outputs(948) <= a xor b;
    outputs(949) <= a and b;
    outputs(950) <= b;
    outputs(951) <= not b;
    outputs(952) <= not (a xor b);
    outputs(953) <= not (a xor b);
    outputs(954) <= not (a xor b);
    outputs(955) <= b;
    outputs(956) <= b and not a;
    outputs(957) <= not (a or b);
    outputs(958) <= b and not a;
    outputs(959) <= b;
    outputs(960) <= a or b;
    outputs(961) <= not (a or b);
    outputs(962) <= b;
    outputs(963) <= b;
    outputs(964) <= b and not a;
    outputs(965) <= not a or b;
    outputs(966) <= a;
    outputs(967) <= a or b;
    outputs(968) <= a or b;
    outputs(969) <= b;
    outputs(970) <= not (a xor b);
    outputs(971) <= a;
    outputs(972) <= b and not a;
    outputs(973) <= b and not a;
    outputs(974) <= a xor b;
    outputs(975) <= b;
    outputs(976) <= a and b;
    outputs(977) <= not a;
    outputs(978) <= not a or b;
    outputs(979) <= a or b;
    outputs(980) <= not (a or b);
    outputs(981) <= not b;
    outputs(982) <= not b;
    outputs(983) <= not a or b;
    outputs(984) <= not a;
    outputs(985) <= not a;
    outputs(986) <= b and not a;
    outputs(987) <= b;
    outputs(988) <= a and b;
    outputs(989) <= not a;
    outputs(990) <= not b;
    outputs(991) <= a and b;
    outputs(992) <= a;
    outputs(993) <= not (a and b);
    outputs(994) <= b;
    outputs(995) <= not (a or b);
    outputs(996) <= not b;
    outputs(997) <= not b;
    outputs(998) <= a;
    outputs(999) <= not b;
    outputs(1000) <= a or b;
    outputs(1001) <= not (a or b);
    outputs(1002) <= a;
    outputs(1003) <= not (a or b);
    outputs(1004) <= a and b;
    outputs(1005) <= a xor b;
    outputs(1006) <= b;
    outputs(1007) <= a xor b;
    outputs(1008) <= b and not a;
    outputs(1009) <= a and b;
    outputs(1010) <= b;
    outputs(1011) <= a and not b;
    outputs(1012) <= not (a or b);
    outputs(1013) <= a;
    outputs(1014) <= not (a or b);
    outputs(1015) <= not b;
    outputs(1016) <= b;
    outputs(1017) <= not a;
    outputs(1018) <= not b;
    outputs(1019) <= not (a or b);
    outputs(1020) <= not a;
    outputs(1021) <= b;
    outputs(1022) <= not a;
    outputs(1023) <= not b;
    outputs(1024) <= not (a or b);
    outputs(1025) <= not a;
    outputs(1026) <= b;
    outputs(1027) <= b;
    outputs(1028) <= a xor b;
    outputs(1029) <= b and not a;
    outputs(1030) <= not b;
    outputs(1031) <= a and not b;
    outputs(1032) <= not a;
    outputs(1033) <= b;
    outputs(1034) <= a;
    outputs(1035) <= not a;
    outputs(1036) <= a;
    outputs(1037) <= not b or a;
    outputs(1038) <= not (a or b);
    outputs(1039) <= b;
    outputs(1040) <= not a;
    outputs(1041) <= a;
    outputs(1042) <= b;
    outputs(1043) <= not (a or b);
    outputs(1044) <= not (a or b);
    outputs(1045) <= b;
    outputs(1046) <= b and not a;
    outputs(1047) <= not a;
    outputs(1048) <= a;
    outputs(1049) <= b;
    outputs(1050) <= not a;
    outputs(1051) <= a and not b;
    outputs(1052) <= not (a xor b);
    outputs(1053) <= not b;
    outputs(1054) <= not a;
    outputs(1055) <= b and not a;
    outputs(1056) <= not a;
    outputs(1057) <= not b;
    outputs(1058) <= not (a or b);
    outputs(1059) <= b and not a;
    outputs(1060) <= a;
    outputs(1061) <= a and b;
    outputs(1062) <= a;
    outputs(1063) <= a and not b;
    outputs(1064) <= b;
    outputs(1065) <= b;
    outputs(1066) <= not a;
    outputs(1067) <= a and b;
    outputs(1068) <= a and b;
    outputs(1069) <= not b;
    outputs(1070) <= not (a and b);
    outputs(1071) <= a and b;
    outputs(1072) <= a and not b;
    outputs(1073) <= a and b;
    outputs(1074) <= a xor b;
    outputs(1075) <= a;
    outputs(1076) <= a and not b;
    outputs(1077) <= a;
    outputs(1078) <= b and not a;
    outputs(1079) <= not b;
    outputs(1080) <= a and not b;
    outputs(1081) <= a;
    outputs(1082) <= not (a or b);
    outputs(1083) <= b and not a;
    outputs(1084) <= a;
    outputs(1085) <= a and b;
    outputs(1086) <= a and not b;
    outputs(1087) <= not a;
    outputs(1088) <= not a;
    outputs(1089) <= a;
    outputs(1090) <= a or b;
    outputs(1091) <= not a;
    outputs(1092) <= a and not b;
    outputs(1093) <= a and not b;
    outputs(1094) <= a and b;
    outputs(1095) <= not (a xor b);
    outputs(1096) <= not a;
    outputs(1097) <= not b;
    outputs(1098) <= b;
    outputs(1099) <= a and b;
    outputs(1100) <= not (a or b);
    outputs(1101) <= a;
    outputs(1102) <= b and not a;
    outputs(1103) <= a and not b;
    outputs(1104) <= not (a or b);
    outputs(1105) <= not b or a;
    outputs(1106) <= a;
    outputs(1107) <= a xor b;
    outputs(1108) <= a xor b;
    outputs(1109) <= a and b;
    outputs(1110) <= not a;
    outputs(1111) <= a xor b;
    outputs(1112) <= not (a and b);
    outputs(1113) <= not b;
    outputs(1114) <= b and not a;
    outputs(1115) <= not b;
    outputs(1116) <= not a;
    outputs(1117) <= b;
    outputs(1118) <= a;
    outputs(1119) <= a;
    outputs(1120) <= not (a xor b);
    outputs(1121) <= not (a or b);
    outputs(1122) <= b;
    outputs(1123) <= not (a xor b);
    outputs(1124) <= b and not a;
    outputs(1125) <= a xor b;
    outputs(1126) <= b;
    outputs(1127) <= a;
    outputs(1128) <= a;
    outputs(1129) <= a and not b;
    outputs(1130) <= not (a or b);
    outputs(1131) <= a and b;
    outputs(1132) <= not (a or b);
    outputs(1133) <= a xor b;
    outputs(1134) <= a and b;
    outputs(1135) <= a xor b;
    outputs(1136) <= b and not a;
    outputs(1137) <= b;
    outputs(1138) <= not a;
    outputs(1139) <= a xor b;
    outputs(1140) <= a;
    outputs(1141) <= not b;
    outputs(1142) <= not (a or b);
    outputs(1143) <= b and not a;
    outputs(1144) <= not (a xor b);
    outputs(1145) <= a;
    outputs(1146) <= a and not b;
    outputs(1147) <= a and not b;
    outputs(1148) <= not b;
    outputs(1149) <= a;
    outputs(1150) <= a and not b;
    outputs(1151) <= not (a or b);
    outputs(1152) <= not b;
    outputs(1153) <= a and not b;
    outputs(1154) <= not b;
    outputs(1155) <= b and not a;
    outputs(1156) <= b;
    outputs(1157) <= a and b;
    outputs(1158) <= not (a and b);
    outputs(1159) <= a and b;
    outputs(1160) <= a;
    outputs(1161) <= not b;
    outputs(1162) <= a;
    outputs(1163) <= not b or a;
    outputs(1164) <= not a or b;
    outputs(1165) <= not b;
    outputs(1166) <= not (a or b);
    outputs(1167) <= a and not b;
    outputs(1168) <= b;
    outputs(1169) <= not (a xor b);
    outputs(1170) <= b and not a;
    outputs(1171) <= not a;
    outputs(1172) <= not a;
    outputs(1173) <= a xor b;
    outputs(1174) <= b and not a;
    outputs(1175) <= b and not a;
    outputs(1176) <= not b;
    outputs(1177) <= b;
    outputs(1178) <= b;
    outputs(1179) <= not (a xor b);
    outputs(1180) <= a xor b;
    outputs(1181) <= a;
    outputs(1182) <= a and not b;
    outputs(1183) <= not (a xor b);
    outputs(1184) <= a;
    outputs(1185) <= not b;
    outputs(1186) <= not a;
    outputs(1187) <= not (a or b);
    outputs(1188) <= not (a or b);
    outputs(1189) <= b and not a;
    outputs(1190) <= not (a or b);
    outputs(1191) <= a;
    outputs(1192) <= not b;
    outputs(1193) <= b and not a;
    outputs(1194) <= b;
    outputs(1195) <= not b;
    outputs(1196) <= not b;
    outputs(1197) <= not (a or b);
    outputs(1198) <= a and b;
    outputs(1199) <= not (a xor b);
    outputs(1200) <= not (a or b);
    outputs(1201) <= a and not b;
    outputs(1202) <= not (a and b);
    outputs(1203) <= b and not a;
    outputs(1204) <= a;
    outputs(1205) <= b and not a;
    outputs(1206) <= not a;
    outputs(1207) <= a;
    outputs(1208) <= a and b;
    outputs(1209) <= b;
    outputs(1210) <= a and not b;
    outputs(1211) <= a and b;
    outputs(1212) <= not (a xor b);
    outputs(1213) <= not a;
    outputs(1214) <= not b;
    outputs(1215) <= not b;
    outputs(1216) <= a and not b;
    outputs(1217) <= b;
    outputs(1218) <= a and not b;
    outputs(1219) <= a;
    outputs(1220) <= a and not b;
    outputs(1221) <= a xor b;
    outputs(1222) <= a and not b;
    outputs(1223) <= a xor b;
    outputs(1224) <= b;
    outputs(1225) <= not b;
    outputs(1226) <= a and not b;
    outputs(1227) <= not a;
    outputs(1228) <= not (a or b);
    outputs(1229) <= a xor b;
    outputs(1230) <= not (a xor b);
    outputs(1231) <= not a;
    outputs(1232) <= not (a or b);
    outputs(1233) <= b;
    outputs(1234) <= b and not a;
    outputs(1235) <= a;
    outputs(1236) <= a;
    outputs(1237) <= not b;
    outputs(1238) <= not a;
    outputs(1239) <= a;
    outputs(1240) <= a xor b;
    outputs(1241) <= not (a or b);
    outputs(1242) <= a;
    outputs(1243) <= b and not a;
    outputs(1244) <= a;
    outputs(1245) <= b and not a;
    outputs(1246) <= a and not b;
    outputs(1247) <= b;
    outputs(1248) <= a xor b;
    outputs(1249) <= a;
    outputs(1250) <= a and not b;
    outputs(1251) <= b;
    outputs(1252) <= b and not a;
    outputs(1253) <= a and b;
    outputs(1254) <= b;
    outputs(1255) <= not (a xor b);
    outputs(1256) <= a and b;
    outputs(1257) <= a and b;
    outputs(1258) <= not b;
    outputs(1259) <= a and not b;
    outputs(1260) <= b and not a;
    outputs(1261) <= a or b;
    outputs(1262) <= a;
    outputs(1263) <= not a;
    outputs(1264) <= b and not a;
    outputs(1265) <= b;
    outputs(1266) <= b;
    outputs(1267) <= b and not a;
    outputs(1268) <= not a;
    outputs(1269) <= a and b;
    outputs(1270) <= a xor b;
    outputs(1271) <= b and not a;
    outputs(1272) <= b;
    outputs(1273) <= not (a or b);
    outputs(1274) <= a and not b;
    outputs(1275) <= not a or b;
    outputs(1276) <= a and b;
    outputs(1277) <= b;
    outputs(1278) <= not b;
    outputs(1279) <= not (a or b);
    outputs(1280) <= a;
    outputs(1281) <= not b;
    outputs(1282) <= not a;
    outputs(1283) <= b;
    outputs(1284) <= b;
    outputs(1285) <= a xor b;
    outputs(1286) <= not a;
    outputs(1287) <= a xor b;
    outputs(1288) <= b;
    outputs(1289) <= not b;
    outputs(1290) <= not b;
    outputs(1291) <= not (a xor b);
    outputs(1292) <= not a;
    outputs(1293) <= not a;
    outputs(1294) <= a and b;
    outputs(1295) <= not a;
    outputs(1296) <= b;
    outputs(1297) <= not (a or b);
    outputs(1298) <= a xor b;
    outputs(1299) <= not (a or b);
    outputs(1300) <= not (a xor b);
    outputs(1301) <= b;
    outputs(1302) <= b and not a;
    outputs(1303) <= b;
    outputs(1304) <= not (a and b);
    outputs(1305) <= not b or a;
    outputs(1306) <= a and not b;
    outputs(1307) <= not b;
    outputs(1308) <= not (a or b);
    outputs(1309) <= b;
    outputs(1310) <= b;
    outputs(1311) <= a and b;
    outputs(1312) <= not b;
    outputs(1313) <= a and not b;
    outputs(1314) <= not a or b;
    outputs(1315) <= not a or b;
    outputs(1316) <= not b;
    outputs(1317) <= not (a or b);
    outputs(1318) <= not (a and b);
    outputs(1319) <= not b;
    outputs(1320) <= not b;
    outputs(1321) <= a;
    outputs(1322) <= a xor b;
    outputs(1323) <= not (a or b);
    outputs(1324) <= a or b;
    outputs(1325) <= not a;
    outputs(1326) <= b;
    outputs(1327) <= b and not a;
    outputs(1328) <= not a;
    outputs(1329) <= not a;
    outputs(1330) <= not b;
    outputs(1331) <= not (a or b);
    outputs(1332) <= not b;
    outputs(1333) <= a;
    outputs(1334) <= b and not a;
    outputs(1335) <= not a;
    outputs(1336) <= b;
    outputs(1337) <= not (a xor b);
    outputs(1338) <= not (a or b);
    outputs(1339) <= not (a xor b);
    outputs(1340) <= not (a xor b);
    outputs(1341) <= not b;
    outputs(1342) <= not a;
    outputs(1343) <= b;
    outputs(1344) <= not a;
    outputs(1345) <= a;
    outputs(1346) <= a and b;
    outputs(1347) <= not a;
    outputs(1348) <= b;
    outputs(1349) <= a;
    outputs(1350) <= not a;
    outputs(1351) <= not b or a;
    outputs(1352) <= not a;
    outputs(1353) <= a;
    outputs(1354) <= not b;
    outputs(1355) <= not (a and b);
    outputs(1356) <= not b;
    outputs(1357) <= not (a xor b);
    outputs(1358) <= a and b;
    outputs(1359) <= a;
    outputs(1360) <= b;
    outputs(1361) <= a or b;
    outputs(1362) <= not a;
    outputs(1363) <= not (a and b);
    outputs(1364) <= not b;
    outputs(1365) <= b and not a;
    outputs(1366) <= a and b;
    outputs(1367) <= not (a xor b);
    outputs(1368) <= not b;
    outputs(1369) <= not (a xor b);
    outputs(1370) <= a or b;
    outputs(1371) <= not a;
    outputs(1372) <= not a or b;
    outputs(1373) <= not b;
    outputs(1374) <= a;
    outputs(1375) <= a;
    outputs(1376) <= a and b;
    outputs(1377) <= not (a or b);
    outputs(1378) <= not b or a;
    outputs(1379) <= not b;
    outputs(1380) <= not a;
    outputs(1381) <= not (a xor b);
    outputs(1382) <= not b;
    outputs(1383) <= a and b;
    outputs(1384) <= not b;
    outputs(1385) <= b;
    outputs(1386) <= a and b;
    outputs(1387) <= not a or b;
    outputs(1388) <= a and b;
    outputs(1389) <= not a;
    outputs(1390) <= not b;
    outputs(1391) <= a;
    outputs(1392) <= b;
    outputs(1393) <= a xor b;
    outputs(1394) <= a and not b;
    outputs(1395) <= not b;
    outputs(1396) <= b;
    outputs(1397) <= a and b;
    outputs(1398) <= not b;
    outputs(1399) <= b;
    outputs(1400) <= a;
    outputs(1401) <= not a;
    outputs(1402) <= not a;
    outputs(1403) <= a and not b;
    outputs(1404) <= not a;
    outputs(1405) <= b;
    outputs(1406) <= a xor b;
    outputs(1407) <= not b or a;
    outputs(1408) <= b and not a;
    outputs(1409) <= b and not a;
    outputs(1410) <= not (a or b);
    outputs(1411) <= a xor b;
    outputs(1412) <= a and not b;
    outputs(1413) <= a or b;
    outputs(1414) <= b and not a;
    outputs(1415) <= a and b;
    outputs(1416) <= a;
    outputs(1417) <= not (a and b);
    outputs(1418) <= a and b;
    outputs(1419) <= not (a xor b);
    outputs(1420) <= not (a xor b);
    outputs(1421) <= b and not a;
    outputs(1422) <= a and b;
    outputs(1423) <= a and not b;
    outputs(1424) <= b and not a;
    outputs(1425) <= a xor b;
    outputs(1426) <= b and not a;
    outputs(1427) <= a and b;
    outputs(1428) <= not b;
    outputs(1429) <= a and b;
    outputs(1430) <= a and b;
    outputs(1431) <= not b;
    outputs(1432) <= not (a xor b);
    outputs(1433) <= not a;
    outputs(1434) <= not b;
    outputs(1435) <= not (a or b);
    outputs(1436) <= a and b;
    outputs(1437) <= not a;
    outputs(1438) <= not a;
    outputs(1439) <= a and b;
    outputs(1440) <= b;
    outputs(1441) <= not b;
    outputs(1442) <= not a;
    outputs(1443) <= a and not b;
    outputs(1444) <= a xor b;
    outputs(1445) <= not (a or b);
    outputs(1446) <= not a;
    outputs(1447) <= not (a xor b);
    outputs(1448) <= not (a or b);
    outputs(1449) <= not a;
    outputs(1450) <= a;
    outputs(1451) <= not b;
    outputs(1452) <= not a;
    outputs(1453) <= a xor b;
    outputs(1454) <= a;
    outputs(1455) <= a;
    outputs(1456) <= a;
    outputs(1457) <= a xor b;
    outputs(1458) <= not (a xor b);
    outputs(1459) <= not a or b;
    outputs(1460) <= not b or a;
    outputs(1461) <= a and not b;
    outputs(1462) <= b;
    outputs(1463) <= b and not a;
    outputs(1464) <= not a;
    outputs(1465) <= a;
    outputs(1466) <= b and not a;
    outputs(1467) <= b;
    outputs(1468) <= a xor b;
    outputs(1469) <= not (a xor b);
    outputs(1470) <= a xor b;
    outputs(1471) <= not a;
    outputs(1472) <= a and not b;
    outputs(1473) <= not b;
    outputs(1474) <= a and not b;
    outputs(1475) <= a xor b;
    outputs(1476) <= a xor b;
    outputs(1477) <= a and b;
    outputs(1478) <= not (a xor b);
    outputs(1479) <= not (a xor b);
    outputs(1480) <= not (a xor b);
    outputs(1481) <= not (a or b);
    outputs(1482) <= not (a xor b);
    outputs(1483) <= not a;
    outputs(1484) <= a;
    outputs(1485) <= b;
    outputs(1486) <= a or b;
    outputs(1487) <= not b or a;
    outputs(1488) <= b;
    outputs(1489) <= not b or a;
    outputs(1490) <= b;
    outputs(1491) <= b;
    outputs(1492) <= b and not a;
    outputs(1493) <= not a;
    outputs(1494) <= a xor b;
    outputs(1495) <= b;
    outputs(1496) <= a and b;
    outputs(1497) <= b and not a;
    outputs(1498) <= not (a xor b);
    outputs(1499) <= b and not a;
    outputs(1500) <= not a;
    outputs(1501) <= not (a or b);
    outputs(1502) <= a xor b;
    outputs(1503) <= a and b;
    outputs(1504) <= not a;
    outputs(1505) <= a xor b;
    outputs(1506) <= not (a or b);
    outputs(1507) <= b;
    outputs(1508) <= b and not a;
    outputs(1509) <= not b;
    outputs(1510) <= a and not b;
    outputs(1511) <= a;
    outputs(1512) <= a and not b;
    outputs(1513) <= not (a xor b);
    outputs(1514) <= a;
    outputs(1515) <= not b;
    outputs(1516) <= b;
    outputs(1517) <= b;
    outputs(1518) <= b;
    outputs(1519) <= b and not a;
    outputs(1520) <= a and not b;
    outputs(1521) <= a xor b;
    outputs(1522) <= not (a xor b);
    outputs(1523) <= not (a or b);
    outputs(1524) <= not a;
    outputs(1525) <= a and b;
    outputs(1526) <= not a;
    outputs(1527) <= b;
    outputs(1528) <= not (a and b);
    outputs(1529) <= a;
    outputs(1530) <= not (a xor b);
    outputs(1531) <= b;
    outputs(1532) <= a;
    outputs(1533) <= not b;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= a;
    outputs(1536) <= not b;
    outputs(1537) <= not b;
    outputs(1538) <= b and not a;
    outputs(1539) <= not a;
    outputs(1540) <= a;
    outputs(1541) <= a;
    outputs(1542) <= b and not a;
    outputs(1543) <= a and not b;
    outputs(1544) <= not a;
    outputs(1545) <= b;
    outputs(1546) <= not a;
    outputs(1547) <= not b;
    outputs(1548) <= a and not b;
    outputs(1549) <= a;
    outputs(1550) <= not (a or b);
    outputs(1551) <= a and b;
    outputs(1552) <= not (a or b);
    outputs(1553) <= not a or b;
    outputs(1554) <= b;
    outputs(1555) <= a xor b;
    outputs(1556) <= b;
    outputs(1557) <= a and b;
    outputs(1558) <= not a;
    outputs(1559) <= b and not a;
    outputs(1560) <= a and b;
    outputs(1561) <= b;
    outputs(1562) <= a xor b;
    outputs(1563) <= a and b;
    outputs(1564) <= a or b;
    outputs(1565) <= a;
    outputs(1566) <= a or b;
    outputs(1567) <= a or b;
    outputs(1568) <= not (a xor b);
    outputs(1569) <= a;
    outputs(1570) <= not b or a;
    outputs(1571) <= not a;
    outputs(1572) <= b and not a;
    outputs(1573) <= b and not a;
    outputs(1574) <= a xor b;
    outputs(1575) <= a and not b;
    outputs(1576) <= not b or a;
    outputs(1577) <= b;
    outputs(1578) <= b;
    outputs(1579) <= not (a or b);
    outputs(1580) <= b and not a;
    outputs(1581) <= not (a or b);
    outputs(1582) <= not b;
    outputs(1583) <= a;
    outputs(1584) <= a and b;
    outputs(1585) <= not b;
    outputs(1586) <= a;
    outputs(1587) <= a;
    outputs(1588) <= a;
    outputs(1589) <= not (a and b);
    outputs(1590) <= not (a or b);
    outputs(1591) <= a xor b;
    outputs(1592) <= not b;
    outputs(1593) <= b and not a;
    outputs(1594) <= a and not b;
    outputs(1595) <= b;
    outputs(1596) <= not (a and b);
    outputs(1597) <= not a;
    outputs(1598) <= not b;
    outputs(1599) <= a xor b;
    outputs(1600) <= not b;
    outputs(1601) <= a and not b;
    outputs(1602) <= not b;
    outputs(1603) <= not a;
    outputs(1604) <= a;
    outputs(1605) <= b;
    outputs(1606) <= b;
    outputs(1607) <= b;
    outputs(1608) <= a or b;
    outputs(1609) <= not (a and b);
    outputs(1610) <= not b;
    outputs(1611) <= b and not a;
    outputs(1612) <= a;
    outputs(1613) <= b;
    outputs(1614) <= b and not a;
    outputs(1615) <= not a;
    outputs(1616) <= b;
    outputs(1617) <= not a;
    outputs(1618) <= b;
    outputs(1619) <= b and not a;
    outputs(1620) <= not a;
    outputs(1621) <= not (a or b);
    outputs(1622) <= a xor b;
    outputs(1623) <= not (a or b);
    outputs(1624) <= not a;
    outputs(1625) <= b;
    outputs(1626) <= b;
    outputs(1627) <= not a;
    outputs(1628) <= a;
    outputs(1629) <= b;
    outputs(1630) <= a or b;
    outputs(1631) <= not b;
    outputs(1632) <= a and not b;
    outputs(1633) <= b;
    outputs(1634) <= a;
    outputs(1635) <= b and not a;
    outputs(1636) <= a;
    outputs(1637) <= not a;
    outputs(1638) <= a and not b;
    outputs(1639) <= a and not b;
    outputs(1640) <= a;
    outputs(1641) <= b and not a;
    outputs(1642) <= not (a xor b);
    outputs(1643) <= not a or b;
    outputs(1644) <= b;
    outputs(1645) <= not a or b;
    outputs(1646) <= b and not a;
    outputs(1647) <= not (a or b);
    outputs(1648) <= not a;
    outputs(1649) <= a or b;
    outputs(1650) <= not (a or b);
    outputs(1651) <= b;
    outputs(1652) <= not (a xor b);
    outputs(1653) <= b;
    outputs(1654) <= not a;
    outputs(1655) <= not (a or b);
    outputs(1656) <= not b or a;
    outputs(1657) <= b;
    outputs(1658) <= b and not a;
    outputs(1659) <= b and not a;
    outputs(1660) <= b and not a;
    outputs(1661) <= a;
    outputs(1662) <= b and not a;
    outputs(1663) <= b and not a;
    outputs(1664) <= not (a and b);
    outputs(1665) <= not (a or b);
    outputs(1666) <= a or b;
    outputs(1667) <= b;
    outputs(1668) <= not (a or b);
    outputs(1669) <= not (a and b);
    outputs(1670) <= not (a or b);
    outputs(1671) <= b;
    outputs(1672) <= not a;
    outputs(1673) <= b and not a;
    outputs(1674) <= b and not a;
    outputs(1675) <= a and b;
    outputs(1676) <= not a;
    outputs(1677) <= a xor b;
    outputs(1678) <= a;
    outputs(1679) <= a;
    outputs(1680) <= a and b;
    outputs(1681) <= not (a or b);
    outputs(1682) <= b;
    outputs(1683) <= not a;
    outputs(1684) <= a and b;
    outputs(1685) <= not (a or b);
    outputs(1686) <= a;
    outputs(1687) <= b and not a;
    outputs(1688) <= a;
    outputs(1689) <= b;
    outputs(1690) <= not (a or b);
    outputs(1691) <= b;
    outputs(1692) <= b and not a;
    outputs(1693) <= not (a or b);
    outputs(1694) <= a;
    outputs(1695) <= b and not a;
    outputs(1696) <= not (a or b);
    outputs(1697) <= a and not b;
    outputs(1698) <= a xor b;
    outputs(1699) <= b and not a;
    outputs(1700) <= not (a or b);
    outputs(1701) <= not b;
    outputs(1702) <= a and not b;
    outputs(1703) <= a xor b;
    outputs(1704) <= b;
    outputs(1705) <= not b or a;
    outputs(1706) <= not a;
    outputs(1707) <= not b;
    outputs(1708) <= not b;
    outputs(1709) <= not (a and b);
    outputs(1710) <= not (a or b);
    outputs(1711) <= a and b;
    outputs(1712) <= b;
    outputs(1713) <= not b;
    outputs(1714) <= not (a xor b);
    outputs(1715) <= not (a or b);
    outputs(1716) <= not (a or b);
    outputs(1717) <= not a;
    outputs(1718) <= b;
    outputs(1719) <= b;
    outputs(1720) <= a;
    outputs(1721) <= not a;
    outputs(1722) <= not a or b;
    outputs(1723) <= b and not a;
    outputs(1724) <= not (a xor b);
    outputs(1725) <= a and b;
    outputs(1726) <= not b;
    outputs(1727) <= not a;
    outputs(1728) <= a and b;
    outputs(1729) <= not a;
    outputs(1730) <= not b;
    outputs(1731) <= b and not a;
    outputs(1732) <= a and b;
    outputs(1733) <= not b;
    outputs(1734) <= b;
    outputs(1735) <= not a or b;
    outputs(1736) <= b;
    outputs(1737) <= not (a xor b);
    outputs(1738) <= a xor b;
    outputs(1739) <= not a;
    outputs(1740) <= a and b;
    outputs(1741) <= a;
    outputs(1742) <= not a or b;
    outputs(1743) <= b and not a;
    outputs(1744) <= a;
    outputs(1745) <= a and not b;
    outputs(1746) <= b;
    outputs(1747) <= a and not b;
    outputs(1748) <= a;
    outputs(1749) <= not b;
    outputs(1750) <= b;
    outputs(1751) <= b and not a;
    outputs(1752) <= a and not b;
    outputs(1753) <= not b;
    outputs(1754) <= a and not b;
    outputs(1755) <= not b;
    outputs(1756) <= a;
    outputs(1757) <= not b;
    outputs(1758) <= a;
    outputs(1759) <= not a;
    outputs(1760) <= a;
    outputs(1761) <= a and b;
    outputs(1762) <= not (a xor b);
    outputs(1763) <= b;
    outputs(1764) <= b and not a;
    outputs(1765) <= not b;
    outputs(1766) <= not b;
    outputs(1767) <= a;
    outputs(1768) <= not b;
    outputs(1769) <= not b;
    outputs(1770) <= a and b;
    outputs(1771) <= not (a xor b);
    outputs(1772) <= not a;
    outputs(1773) <= b and not a;
    outputs(1774) <= not a;
    outputs(1775) <= a and not b;
    outputs(1776) <= b and not a;
    outputs(1777) <= b;
    outputs(1778) <= a xor b;
    outputs(1779) <= not a;
    outputs(1780) <= a;
    outputs(1781) <= a and not b;
    outputs(1782) <= a and b;
    outputs(1783) <= a;
    outputs(1784) <= not a;
    outputs(1785) <= b and not a;
    outputs(1786) <= a;
    outputs(1787) <= a and not b;
    outputs(1788) <= not a;
    outputs(1789) <= a and b;
    outputs(1790) <= a xor b;
    outputs(1791) <= not b;
    outputs(1792) <= a xor b;
    outputs(1793) <= not (a or b);
    outputs(1794) <= not (a or b);
    outputs(1795) <= a xor b;
    outputs(1796) <= not b;
    outputs(1797) <= b and not a;
    outputs(1798) <= b;
    outputs(1799) <= not (a or b);
    outputs(1800) <= a or b;
    outputs(1801) <= b;
    outputs(1802) <= b;
    outputs(1803) <= not b;
    outputs(1804) <= b;
    outputs(1805) <= a and b;
    outputs(1806) <= a and b;
    outputs(1807) <= a;
    outputs(1808) <= not b;
    outputs(1809) <= not a;
    outputs(1810) <= not b or a;
    outputs(1811) <= not b;
    outputs(1812) <= a and not b;
    outputs(1813) <= not (a or b);
    outputs(1814) <= a and b;
    outputs(1815) <= a;
    outputs(1816) <= a;
    outputs(1817) <= a;
    outputs(1818) <= not b;
    outputs(1819) <= not b;
    outputs(1820) <= not a;
    outputs(1821) <= b;
    outputs(1822) <= b;
    outputs(1823) <= b and not a;
    outputs(1824) <= b;
    outputs(1825) <= a;
    outputs(1826) <= a and b;
    outputs(1827) <= not a;
    outputs(1828) <= not a;
    outputs(1829) <= a and not b;
    outputs(1830) <= not a;
    outputs(1831) <= a;
    outputs(1832) <= b and not a;
    outputs(1833) <= not (a or b);
    outputs(1834) <= not (a or b);
    outputs(1835) <= a xor b;
    outputs(1836) <= not a;
    outputs(1837) <= not (a or b);
    outputs(1838) <= a;
    outputs(1839) <= b and not a;
    outputs(1840) <= not b;
    outputs(1841) <= not (a xor b);
    outputs(1842) <= a;
    outputs(1843) <= b and not a;
    outputs(1844) <= a;
    outputs(1845) <= not (a or b);
    outputs(1846) <= not b or a;
    outputs(1847) <= not b or a;
    outputs(1848) <= not (a or b);
    outputs(1849) <= b and not a;
    outputs(1850) <= not (a xor b);
    outputs(1851) <= b;
    outputs(1852) <= a and not b;
    outputs(1853) <= b;
    outputs(1854) <= b;
    outputs(1855) <= b;
    outputs(1856) <= a or b;
    outputs(1857) <= a and not b;
    outputs(1858) <= not (a or b);
    outputs(1859) <= b;
    outputs(1860) <= a and not b;
    outputs(1861) <= not a;
    outputs(1862) <= not b;
    outputs(1863) <= b;
    outputs(1864) <= b and not a;
    outputs(1865) <= not (a or b);
    outputs(1866) <= not (a and b);
    outputs(1867) <= b and not a;
    outputs(1868) <= a;
    outputs(1869) <= not a or b;
    outputs(1870) <= not a;
    outputs(1871) <= b and not a;
    outputs(1872) <= a and not b;
    outputs(1873) <= b and not a;
    outputs(1874) <= not (a or b);
    outputs(1875) <= b;
    outputs(1876) <= not b;
    outputs(1877) <= a xor b;
    outputs(1878) <= not b;
    outputs(1879) <= not (a or b);
    outputs(1880) <= a;
    outputs(1881) <= b and not a;
    outputs(1882) <= a and b;
    outputs(1883) <= not (a or b);
    outputs(1884) <= a and not b;
    outputs(1885) <= not (a xor b);
    outputs(1886) <= b and not a;
    outputs(1887) <= b;
    outputs(1888) <= not b;
    outputs(1889) <= not a;
    outputs(1890) <= a and not b;
    outputs(1891) <= not b;
    outputs(1892) <= a and b;
    outputs(1893) <= a and b;
    outputs(1894) <= not b;
    outputs(1895) <= b;
    outputs(1896) <= not a or b;
    outputs(1897) <= not (a or b);
    outputs(1898) <= not (a xor b);
    outputs(1899) <= a and b;
    outputs(1900) <= a and b;
    outputs(1901) <= b and not a;
    outputs(1902) <= b and not a;
    outputs(1903) <= not a;
    outputs(1904) <= not (a xor b);
    outputs(1905) <= not b;
    outputs(1906) <= a and not b;
    outputs(1907) <= not (a or b);
    outputs(1908) <= a;
    outputs(1909) <= not b;
    outputs(1910) <= not b;
    outputs(1911) <= not b;
    outputs(1912) <= not (a xor b);
    outputs(1913) <= not a;
    outputs(1914) <= not b or a;
    outputs(1915) <= a;
    outputs(1916) <= a and not b;
    outputs(1917) <= not (a or b);
    outputs(1918) <= not a;
    outputs(1919) <= not (a or b);
    outputs(1920) <= b;
    outputs(1921) <= b and not a;
    outputs(1922) <= not a;
    outputs(1923) <= a and b;
    outputs(1924) <= a;
    outputs(1925) <= b and not a;
    outputs(1926) <= a and not b;
    outputs(1927) <= a;
    outputs(1928) <= b and not a;
    outputs(1929) <= a;
    outputs(1930) <= not b;
    outputs(1931) <= not (a xor b);
    outputs(1932) <= not a;
    outputs(1933) <= a or b;
    outputs(1934) <= not b;
    outputs(1935) <= not a;
    outputs(1936) <= not (a or b);
    outputs(1937) <= b;
    outputs(1938) <= not (a or b);
    outputs(1939) <= a and b;
    outputs(1940) <= not a;
    outputs(1941) <= not b;
    outputs(1942) <= b;
    outputs(1943) <= a;
    outputs(1944) <= not a;
    outputs(1945) <= a xor b;
    outputs(1946) <= not (a or b);
    outputs(1947) <= a and not b;
    outputs(1948) <= not (a or b);
    outputs(1949) <= a xor b;
    outputs(1950) <= not b;
    outputs(1951) <= a;
    outputs(1952) <= a and not b;
    outputs(1953) <= not (a or b);
    outputs(1954) <= a;
    outputs(1955) <= a;
    outputs(1956) <= not a or b;
    outputs(1957) <= b;
    outputs(1958) <= a;
    outputs(1959) <= a and b;
    outputs(1960) <= b;
    outputs(1961) <= a and b;
    outputs(1962) <= b;
    outputs(1963) <= a and b;
    outputs(1964) <= not (a or b);
    outputs(1965) <= not (a and b);
    outputs(1966) <= not (a xor b);
    outputs(1967) <= not a;
    outputs(1968) <= b;
    outputs(1969) <= a and not b;
    outputs(1970) <= not a;
    outputs(1971) <= b and not a;
    outputs(1972) <= b and not a;
    outputs(1973) <= b and not a;
    outputs(1974) <= a and b;
    outputs(1975) <= b;
    outputs(1976) <= a and not b;
    outputs(1977) <= b;
    outputs(1978) <= not (a xor b);
    outputs(1979) <= a;
    outputs(1980) <= a and not b;
    outputs(1981) <= a and b;
    outputs(1982) <= a and not b;
    outputs(1983) <= b;
    outputs(1984) <= not b or a;
    outputs(1985) <= a;
    outputs(1986) <= not a or b;
    outputs(1987) <= a or b;
    outputs(1988) <= a xor b;
    outputs(1989) <= not a;
    outputs(1990) <= a xor b;
    outputs(1991) <= a xor b;
    outputs(1992) <= a and not b;
    outputs(1993) <= a and b;
    outputs(1994) <= not b or a;
    outputs(1995) <= not b;
    outputs(1996) <= a;
    outputs(1997) <= b and not a;
    outputs(1998) <= not b;
    outputs(1999) <= a;
    outputs(2000) <= not a;
    outputs(2001) <= a and not b;
    outputs(2002) <= b and not a;
    outputs(2003) <= not (a xor b);
    outputs(2004) <= b and not a;
    outputs(2005) <= a or b;
    outputs(2006) <= b;
    outputs(2007) <= not b;
    outputs(2008) <= not (a xor b);
    outputs(2009) <= not (a or b);
    outputs(2010) <= not b;
    outputs(2011) <= a and not b;
    outputs(2012) <= not a;
    outputs(2013) <= b;
    outputs(2014) <= a and b;
    outputs(2015) <= b;
    outputs(2016) <= not a or b;
    outputs(2017) <= a xor b;
    outputs(2018) <= b;
    outputs(2019) <= not a;
    outputs(2020) <= b and not a;
    outputs(2021) <= not a;
    outputs(2022) <= not b;
    outputs(2023) <= b;
    outputs(2024) <= a and b;
    outputs(2025) <= not (a xor b);
    outputs(2026) <= not a;
    outputs(2027) <= not (a xor b);
    outputs(2028) <= a and not b;
    outputs(2029) <= not (a xor b);
    outputs(2030) <= not a;
    outputs(2031) <= not b;
    outputs(2032) <= not a;
    outputs(2033) <= not (a or b);
    outputs(2034) <= a and b;
    outputs(2035) <= b and not a;
    outputs(2036) <= a and b;
    outputs(2037) <= not a;
    outputs(2038) <= b;
    outputs(2039) <= b;
    outputs(2040) <= not a;
    outputs(2041) <= a and b;
    outputs(2042) <= not (a xor b);
    outputs(2043) <= b and not a;
    outputs(2044) <= not a or b;
    outputs(2045) <= not b;
    outputs(2046) <= not (a or b);
    outputs(2047) <= not (a or b);
    outputs(2048) <= a and not b;
    outputs(2049) <= not a;
    outputs(2050) <= not b;
    outputs(2051) <= not b;
    outputs(2052) <= a;
    outputs(2053) <= not (a xor b);
    outputs(2054) <= not b;
    outputs(2055) <= not (a or b);
    outputs(2056) <= a and b;
    outputs(2057) <= not b;
    outputs(2058) <= a and b;
    outputs(2059) <= not (a or b);
    outputs(2060) <= a xor b;
    outputs(2061) <= a and b;
    outputs(2062) <= not a or b;
    outputs(2063) <= not (a or b);
    outputs(2064) <= not (a and b);
    outputs(2065) <= a and not b;
    outputs(2066) <= not (a xor b);
    outputs(2067) <= not (a or b);
    outputs(2068) <= b;
    outputs(2069) <= not b;
    outputs(2070) <= not a;
    outputs(2071) <= a and not b;
    outputs(2072) <= b;
    outputs(2073) <= a;
    outputs(2074) <= not (a or b);
    outputs(2075) <= not b or a;
    outputs(2076) <= not (a or b);
    outputs(2077) <= not (a or b);
    outputs(2078) <= a xor b;
    outputs(2079) <= not (a or b);
    outputs(2080) <= a and not b;
    outputs(2081) <= not b;
    outputs(2082) <= not b or a;
    outputs(2083) <= a xor b;
    outputs(2084) <= not b;
    outputs(2085) <= a and not b;
    outputs(2086) <= not b;
    outputs(2087) <= b;
    outputs(2088) <= not a or b;
    outputs(2089) <= not b;
    outputs(2090) <= a or b;
    outputs(2091) <= not b;
    outputs(2092) <= a xor b;
    outputs(2093) <= not (a or b);
    outputs(2094) <= not (a or b);
    outputs(2095) <= not a or b;
    outputs(2096) <= a xor b;
    outputs(2097) <= not a;
    outputs(2098) <= not b;
    outputs(2099) <= not b;
    outputs(2100) <= a;
    outputs(2101) <= not b;
    outputs(2102) <= b;
    outputs(2103) <= not a;
    outputs(2104) <= not (a and b);
    outputs(2105) <= a or b;
    outputs(2106) <= not (a xor b);
    outputs(2107) <= a;
    outputs(2108) <= not b;
    outputs(2109) <= b and not a;
    outputs(2110) <= not (a xor b);
    outputs(2111) <= a;
    outputs(2112) <= b and not a;
    outputs(2113) <= not b;
    outputs(2114) <= a;
    outputs(2115) <= b;
    outputs(2116) <= a and b;
    outputs(2117) <= not a;
    outputs(2118) <= a or b;
    outputs(2119) <= b and not a;
    outputs(2120) <= not (a or b);
    outputs(2121) <= b and not a;
    outputs(2122) <= not a;
    outputs(2123) <= a;
    outputs(2124) <= not (a or b);
    outputs(2125) <= a and b;
    outputs(2126) <= not b;
    outputs(2127) <= not (a xor b);
    outputs(2128) <= b;
    outputs(2129) <= b;
    outputs(2130) <= not (a or b);
    outputs(2131) <= a;
    outputs(2132) <= a;
    outputs(2133) <= a and b;
    outputs(2134) <= not (a or b);
    outputs(2135) <= b;
    outputs(2136) <= b;
    outputs(2137) <= a;
    outputs(2138) <= not (a or b);
    outputs(2139) <= a xor b;
    outputs(2140) <= a and b;
    outputs(2141) <= a and b;
    outputs(2142) <= a;
    outputs(2143) <= a;
    outputs(2144) <= a and b;
    outputs(2145) <= a and not b;
    outputs(2146) <= b;
    outputs(2147) <= not b;
    outputs(2148) <= not (a and b);
    outputs(2149) <= not b;
    outputs(2150) <= not b or a;
    outputs(2151) <= not (a xor b);
    outputs(2152) <= not (a and b);
    outputs(2153) <= b and not a;
    outputs(2154) <= not b or a;
    outputs(2155) <= not (a xor b);
    outputs(2156) <= b;
    outputs(2157) <= a;
    outputs(2158) <= not (a or b);
    outputs(2159) <= not (a xor b);
    outputs(2160) <= b;
    outputs(2161) <= not b;
    outputs(2162) <= a xor b;
    outputs(2163) <= not a;
    outputs(2164) <= b and not a;
    outputs(2165) <= a;
    outputs(2166) <= not (a or b);
    outputs(2167) <= not a;
    outputs(2168) <= b and not a;
    outputs(2169) <= a and b;
    outputs(2170) <= b;
    outputs(2171) <= b and not a;
    outputs(2172) <= b;
    outputs(2173) <= not (a and b);
    outputs(2174) <= b;
    outputs(2175) <= not b;
    outputs(2176) <= not (a or b);
    outputs(2177) <= a and not b;
    outputs(2178) <= a;
    outputs(2179) <= not a;
    outputs(2180) <= not (a or b);
    outputs(2181) <= not (a xor b);
    outputs(2182) <= b;
    outputs(2183) <= a;
    outputs(2184) <= a;
    outputs(2185) <= b and not a;
    outputs(2186) <= a and b;
    outputs(2187) <= not a or b;
    outputs(2188) <= a and b;
    outputs(2189) <= not (a and b);
    outputs(2190) <= a;
    outputs(2191) <= a;
    outputs(2192) <= not b;
    outputs(2193) <= a;
    outputs(2194) <= not b;
    outputs(2195) <= not a;
    outputs(2196) <= a xor b;
    outputs(2197) <= a;
    outputs(2198) <= not b or a;
    outputs(2199) <= not (a xor b);
    outputs(2200) <= not (a or b);
    outputs(2201) <= b and not a;
    outputs(2202) <= not a or b;
    outputs(2203) <= not (a and b);
    outputs(2204) <= not (a xor b);
    outputs(2205) <= not (a or b);
    outputs(2206) <= not a;
    outputs(2207) <= not (a xor b);
    outputs(2208) <= a or b;
    outputs(2209) <= a and not b;
    outputs(2210) <= not b;
    outputs(2211) <= not (a or b);
    outputs(2212) <= not (a xor b);
    outputs(2213) <= not b or a;
    outputs(2214) <= not (a or b);
    outputs(2215) <= b;
    outputs(2216) <= a or b;
    outputs(2217) <= not a or b;
    outputs(2218) <= b;
    outputs(2219) <= a or b;
    outputs(2220) <= a and not b;
    outputs(2221) <= b;
    outputs(2222) <= a or b;
    outputs(2223) <= not b;
    outputs(2224) <= a and not b;
    outputs(2225) <= a;
    outputs(2226) <= not (a or b);
    outputs(2227) <= a;
    outputs(2228) <= not b;
    outputs(2229) <= b and not a;
    outputs(2230) <= not a or b;
    outputs(2231) <= not (a or b);
    outputs(2232) <= a;
    outputs(2233) <= not b or a;
    outputs(2234) <= b and not a;
    outputs(2235) <= not b;
    outputs(2236) <= not (a xor b);
    outputs(2237) <= b;
    outputs(2238) <= not a;
    outputs(2239) <= not (a xor b);
    outputs(2240) <= not (a or b);
    outputs(2241) <= not (a and b);
    outputs(2242) <= a xor b;
    outputs(2243) <= a and not b;
    outputs(2244) <= b;
    outputs(2245) <= a or b;
    outputs(2246) <= not b;
    outputs(2247) <= a;
    outputs(2248) <= not (a xor b);
    outputs(2249) <= not a;
    outputs(2250) <= a;
    outputs(2251) <= a or b;
    outputs(2252) <= not a;
    outputs(2253) <= not b;
    outputs(2254) <= a;
    outputs(2255) <= b;
    outputs(2256) <= not b;
    outputs(2257) <= not (a or b);
    outputs(2258) <= not (a or b);
    outputs(2259) <= a;
    outputs(2260) <= b and not a;
    outputs(2261) <= not b;
    outputs(2262) <= a xor b;
    outputs(2263) <= not a;
    outputs(2264) <= b and not a;
    outputs(2265) <= not b;
    outputs(2266) <= not (a xor b);
    outputs(2267) <= not (a xor b);
    outputs(2268) <= a;
    outputs(2269) <= b and not a;
    outputs(2270) <= a and not b;
    outputs(2271) <= a and b;
    outputs(2272) <= not (a or b);
    outputs(2273) <= a;
    outputs(2274) <= a xor b;
    outputs(2275) <= not (a xor b);
    outputs(2276) <= not (a or b);
    outputs(2277) <= a and b;
    outputs(2278) <= not b;
    outputs(2279) <= not b;
    outputs(2280) <= a xor b;
    outputs(2281) <= b;
    outputs(2282) <= not a or b;
    outputs(2283) <= b;
    outputs(2284) <= a xor b;
    outputs(2285) <= a xor b;
    outputs(2286) <= a;
    outputs(2287) <= a;
    outputs(2288) <= not (a and b);
    outputs(2289) <= a;
    outputs(2290) <= a xor b;
    outputs(2291) <= a xor b;
    outputs(2292) <= a and b;
    outputs(2293) <= not a;
    outputs(2294) <= b;
    outputs(2295) <= not a;
    outputs(2296) <= a and b;
    outputs(2297) <= a and b;
    outputs(2298) <= a and not b;
    outputs(2299) <= not a;
    outputs(2300) <= not b;
    outputs(2301) <= not a;
    outputs(2302) <= not (a or b);
    outputs(2303) <= not a;
    outputs(2304) <= not b;
    outputs(2305) <= not (a or b);
    outputs(2306) <= not a;
    outputs(2307) <= a;
    outputs(2308) <= b and not a;
    outputs(2309) <= a and not b;
    outputs(2310) <= b and not a;
    outputs(2311) <= a or b;
    outputs(2312) <= b;
    outputs(2313) <= b;
    outputs(2314) <= a and not b;
    outputs(2315) <= not a;
    outputs(2316) <= b;
    outputs(2317) <= a and b;
    outputs(2318) <= not a;
    outputs(2319) <= not (a or b);
    outputs(2320) <= a xor b;
    outputs(2321) <= not (a and b);
    outputs(2322) <= a and not b;
    outputs(2323) <= a;
    outputs(2324) <= a and not b;
    outputs(2325) <= not a;
    outputs(2326) <= a and not b;
    outputs(2327) <= a xor b;
    outputs(2328) <= not (a or b);
    outputs(2329) <= not (a or b);
    outputs(2330) <= a and b;
    outputs(2331) <= not (a or b);
    outputs(2332) <= not a;
    outputs(2333) <= a and not b;
    outputs(2334) <= a and not b;
    outputs(2335) <= not a or b;
    outputs(2336) <= not b;
    outputs(2337) <= not (a or b);
    outputs(2338) <= not a;
    outputs(2339) <= a and b;
    outputs(2340) <= not a;
    outputs(2341) <= a and not b;
    outputs(2342) <= b and not a;
    outputs(2343) <= a and not b;
    outputs(2344) <= b and not a;
    outputs(2345) <= not b;
    outputs(2346) <= a;
    outputs(2347) <= not (a or b);
    outputs(2348) <= a and not b;
    outputs(2349) <= a and b;
    outputs(2350) <= not (a or b);
    outputs(2351) <= not b;
    outputs(2352) <= b and not a;
    outputs(2353) <= b;
    outputs(2354) <= not b;
    outputs(2355) <= not a;
    outputs(2356) <= not b or a;
    outputs(2357) <= b and not a;
    outputs(2358) <= a and b;
    outputs(2359) <= not (a xor b);
    outputs(2360) <= not (a or b);
    outputs(2361) <= a;
    outputs(2362) <= not (a xor b);
    outputs(2363) <= not b;
    outputs(2364) <= not a;
    outputs(2365) <= not (a xor b);
    outputs(2366) <= not a or b;
    outputs(2367) <= a;
    outputs(2368) <= a and b;
    outputs(2369) <= not (a or b);
    outputs(2370) <= not (a or b);
    outputs(2371) <= not a;
    outputs(2372) <= a and b;
    outputs(2373) <= not (a or b);
    outputs(2374) <= not (a xor b);
    outputs(2375) <= b and not a;
    outputs(2376) <= b and not a;
    outputs(2377) <= not (a or b);
    outputs(2378) <= not (a or b);
    outputs(2379) <= a and b;
    outputs(2380) <= not (a and b);
    outputs(2381) <= a and b;
    outputs(2382) <= not a or b;
    outputs(2383) <= not b;
    outputs(2384) <= not b;
    outputs(2385) <= a and not b;
    outputs(2386) <= not (a and b);
    outputs(2387) <= not a;
    outputs(2388) <= not a;
    outputs(2389) <= b and not a;
    outputs(2390) <= b and not a;
    outputs(2391) <= not a;
    outputs(2392) <= a;
    outputs(2393) <= b and not a;
    outputs(2394) <= a xor b;
    outputs(2395) <= b and not a;
    outputs(2396) <= a and not b;
    outputs(2397) <= not b or a;
    outputs(2398) <= a xor b;
    outputs(2399) <= not b;
    outputs(2400) <= a xor b;
    outputs(2401) <= a and b;
    outputs(2402) <= a and not b;
    outputs(2403) <= not a;
    outputs(2404) <= not b;
    outputs(2405) <= a and not b;
    outputs(2406) <= not (a or b);
    outputs(2407) <= a and not b;
    outputs(2408) <= b and not a;
    outputs(2409) <= a and b;
    outputs(2410) <= not (a or b);
    outputs(2411) <= a xor b;
    outputs(2412) <= a xor b;
    outputs(2413) <= not a or b;
    outputs(2414) <= not (a xor b);
    outputs(2415) <= a and b;
    outputs(2416) <= a and b;
    outputs(2417) <= a;
    outputs(2418) <= a;
    outputs(2419) <= not a;
    outputs(2420) <= not (a or b);
    outputs(2421) <= b and not a;
    outputs(2422) <= a and b;
    outputs(2423) <= a and not b;
    outputs(2424) <= b and not a;
    outputs(2425) <= not (a or b);
    outputs(2426) <= a and not b;
    outputs(2427) <= not (a or b);
    outputs(2428) <= b;
    outputs(2429) <= not a;
    outputs(2430) <= b;
    outputs(2431) <= not a;
    outputs(2432) <= b and not a;
    outputs(2433) <= a and not b;
    outputs(2434) <= not (a or b);
    outputs(2435) <= a and not b;
    outputs(2436) <= b and not a;
    outputs(2437) <= a;
    outputs(2438) <= b;
    outputs(2439) <= not (a or b);
    outputs(2440) <= b;
    outputs(2441) <= a or b;
    outputs(2442) <= not (a or b);
    outputs(2443) <= a;
    outputs(2444) <= a;
    outputs(2445) <= a and not b;
    outputs(2446) <= a;
    outputs(2447) <= b and not a;
    outputs(2448) <= a and not b;
    outputs(2449) <= a and b;
    outputs(2450) <= not b;
    outputs(2451) <= a;
    outputs(2452) <= a and not b;
    outputs(2453) <= b;
    outputs(2454) <= not a;
    outputs(2455) <= b and not a;
    outputs(2456) <= a and not b;
    outputs(2457) <= b;
    outputs(2458) <= b and not a;
    outputs(2459) <= a and b;
    outputs(2460) <= b and not a;
    outputs(2461) <= a;
    outputs(2462) <= not b;
    outputs(2463) <= not b;
    outputs(2464) <= not (a or b);
    outputs(2465) <= a xor b;
    outputs(2466) <= a and not b;
    outputs(2467) <= not a;
    outputs(2468) <= not b;
    outputs(2469) <= a;
    outputs(2470) <= not a;
    outputs(2471) <= not a;
    outputs(2472) <= not b;
    outputs(2473) <= not (a xor b);
    outputs(2474) <= b;
    outputs(2475) <= not a;
    outputs(2476) <= not b;
    outputs(2477) <= b;
    outputs(2478) <= not (a or b);
    outputs(2479) <= not b;
    outputs(2480) <= not a;
    outputs(2481) <= a;
    outputs(2482) <= a and b;
    outputs(2483) <= a;
    outputs(2484) <= 1'b0;
    outputs(2485) <= not a;
    outputs(2486) <= a and b;
    outputs(2487) <= b;
    outputs(2488) <= a;
    outputs(2489) <= not a;
    outputs(2490) <= a and b;
    outputs(2491) <= not (a xor b);
    outputs(2492) <= b and not a;
    outputs(2493) <= not (a or b);
    outputs(2494) <= not a;
    outputs(2495) <= a xor b;
    outputs(2496) <= not (a or b);
    outputs(2497) <= a and not b;
    outputs(2498) <= a and b;
    outputs(2499) <= not (a or b);
    outputs(2500) <= not b or a;
    outputs(2501) <= b;
    outputs(2502) <= not b;
    outputs(2503) <= a and not b;
    outputs(2504) <= b and not a;
    outputs(2505) <= not b;
    outputs(2506) <= not (a or b);
    outputs(2507) <= a xor b;
    outputs(2508) <= a and b;
    outputs(2509) <= not a;
    outputs(2510) <= not (a xor b);
    outputs(2511) <= a and b;
    outputs(2512) <= a;
    outputs(2513) <= not a;
    outputs(2514) <= b and not a;
    outputs(2515) <= not (a xor b);
    outputs(2516) <= a xor b;
    outputs(2517) <= a and b;
    outputs(2518) <= a;
    outputs(2519) <= not b;
    outputs(2520) <= not b;
    outputs(2521) <= a;
    outputs(2522) <= not a;
    outputs(2523) <= a and not b;
    outputs(2524) <= not b;
    outputs(2525) <= not (a or b);
    outputs(2526) <= b and not a;
    outputs(2527) <= not a;
    outputs(2528) <= not a;
    outputs(2529) <= a or b;
    outputs(2530) <= not (a xor b);
    outputs(2531) <= b and not a;
    outputs(2532) <= a and not b;
    outputs(2533) <= a and not b;
    outputs(2534) <= not (a or b);
    outputs(2535) <= a and b;
    outputs(2536) <= not (a or b);
    outputs(2537) <= a;
    outputs(2538) <= not (a xor b);
    outputs(2539) <= b and not a;
    outputs(2540) <= not b;
    outputs(2541) <= b;
    outputs(2542) <= not b;
    outputs(2543) <= b and not a;
    outputs(2544) <= a and not b;
    outputs(2545) <= a and not b;
    outputs(2546) <= b and not a;
    outputs(2547) <= a and b;
    outputs(2548) <= not a;
    outputs(2549) <= a and not b;
    outputs(2550) <= b and not a;
    outputs(2551) <= b and not a;
    outputs(2552) <= a and b;
    outputs(2553) <= not (a or b);
    outputs(2554) <= not (a or b);
    outputs(2555) <= a and b;
    outputs(2556) <= a xor b;
    outputs(2557) <= not (a or b);
    outputs(2558) <= not a;
    outputs(2559) <= not b;
end Behavioral;
