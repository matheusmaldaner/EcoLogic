module logic_network(
    input wire [255:0] inputs,
    output wire [10239:0] outputs
);

    wire [10239:0] layer0_outputs;

    assign layer0_outputs[0] = ~((inputs[100]) | (inputs[42]));
    assign layer0_outputs[1] = ~(inputs[235]);
    assign layer0_outputs[2] = ~(inputs[246]) | (inputs[241]);
    assign layer0_outputs[3] = ~(inputs[184]) | (inputs[146]);
    assign layer0_outputs[4] = ~((inputs[162]) | (inputs[216]));
    assign layer0_outputs[5] = ~(inputs[94]) | (inputs[161]);
    assign layer0_outputs[6] = (inputs[133]) | (inputs[1]);
    assign layer0_outputs[7] = ~((inputs[53]) ^ (inputs[160]));
    assign layer0_outputs[8] = ~((inputs[189]) & (inputs[254]));
    assign layer0_outputs[9] = (inputs[65]) | (inputs[227]);
    assign layer0_outputs[10] = ~(inputs[168]) | (inputs[33]);
    assign layer0_outputs[11] = (inputs[75]) ^ (inputs[18]);
    assign layer0_outputs[12] = ~(inputs[58]) | (inputs[243]);
    assign layer0_outputs[13] = ~((inputs[104]) | (inputs[253]));
    assign layer0_outputs[14] = (inputs[213]) & ~(inputs[103]);
    assign layer0_outputs[15] = ~((inputs[160]) | (inputs[214]));
    assign layer0_outputs[16] = ~(inputs[46]);
    assign layer0_outputs[17] = inputs[0];
    assign layer0_outputs[18] = ~((inputs[109]) | (inputs[50]));
    assign layer0_outputs[19] = (inputs[175]) & ~(inputs[141]);
    assign layer0_outputs[20] = (inputs[229]) & ~(inputs[130]);
    assign layer0_outputs[21] = ~(inputs[212]) | (inputs[46]);
    assign layer0_outputs[22] = ~((inputs[100]) & (inputs[135]));
    assign layer0_outputs[23] = (inputs[115]) & (inputs[112]);
    assign layer0_outputs[24] = (inputs[227]) & ~(inputs[113]);
    assign layer0_outputs[25] = ~(inputs[236]) | (inputs[15]);
    assign layer0_outputs[26] = (inputs[123]) & (inputs[48]);
    assign layer0_outputs[27] = (inputs[187]) | (inputs[62]);
    assign layer0_outputs[28] = (inputs[10]) & ~(inputs[192]);
    assign layer0_outputs[29] = (inputs[220]) ^ (inputs[64]);
    assign layer0_outputs[30] = inputs[215];
    assign layer0_outputs[31] = ~((inputs[63]) | (inputs[83]));
    assign layer0_outputs[32] = (inputs[200]) | (inputs[155]);
    assign layer0_outputs[33] = inputs[94];
    assign layer0_outputs[34] = (inputs[57]) | (inputs[34]);
    assign layer0_outputs[35] = ~((inputs[60]) | (inputs[15]));
    assign layer0_outputs[36] = ~(inputs[74]) | (inputs[96]);
    assign layer0_outputs[37] = ~((inputs[116]) | (inputs[188]));
    assign layer0_outputs[38] = 1'b0;
    assign layer0_outputs[39] = inputs[119];
    assign layer0_outputs[40] = (inputs[180]) & ~(inputs[66]);
    assign layer0_outputs[41] = (inputs[41]) | (inputs[247]);
    assign layer0_outputs[42] = ~(inputs[164]);
    assign layer0_outputs[43] = (inputs[171]) | (inputs[140]);
    assign layer0_outputs[44] = ~(inputs[179]);
    assign layer0_outputs[45] = ~((inputs[139]) | (inputs[188]));
    assign layer0_outputs[46] = ~(inputs[228]);
    assign layer0_outputs[47] = ~(inputs[14]);
    assign layer0_outputs[48] = ~(inputs[16]) | (inputs[242]);
    assign layer0_outputs[49] = ~(inputs[28]) | (inputs[206]);
    assign layer0_outputs[50] = ~(inputs[14]) | (inputs[171]);
    assign layer0_outputs[51] = ~(inputs[152]) | (inputs[203]);
    assign layer0_outputs[52] = (inputs[170]) & ~(inputs[213]);
    assign layer0_outputs[53] = (inputs[196]) | (inputs[203]);
    assign layer0_outputs[54] = ~((inputs[98]) | (inputs[137]));
    assign layer0_outputs[55] = ~(inputs[17]);
    assign layer0_outputs[56] = ~(inputs[228]);
    assign layer0_outputs[57] = ~(inputs[23]) | (inputs[125]);
    assign layer0_outputs[58] = ~(inputs[159]);
    assign layer0_outputs[59] = ~((inputs[237]) ^ (inputs[181]));
    assign layer0_outputs[60] = ~((inputs[8]) | (inputs[107]));
    assign layer0_outputs[61] = ~((inputs[182]) ^ (inputs[152]));
    assign layer0_outputs[62] = (inputs[105]) & ~(inputs[176]);
    assign layer0_outputs[63] = (inputs[221]) | (inputs[160]);
    assign layer0_outputs[64] = ~(inputs[32]) | (inputs[244]);
    assign layer0_outputs[65] = (inputs[244]) & ~(inputs[158]);
    assign layer0_outputs[66] = inputs[197];
    assign layer0_outputs[67] = ~(inputs[3]);
    assign layer0_outputs[68] = ~((inputs[165]) | (inputs[145]));
    assign layer0_outputs[69] = (inputs[21]) | (inputs[84]);
    assign layer0_outputs[70] = ~(inputs[72]);
    assign layer0_outputs[71] = ~((inputs[54]) | (inputs[140]));
    assign layer0_outputs[72] = ~((inputs[233]) & (inputs[174]));
    assign layer0_outputs[73] = inputs[98];
    assign layer0_outputs[74] = ~((inputs[155]) ^ (inputs[178]));
    assign layer0_outputs[75] = inputs[119];
    assign layer0_outputs[76] = inputs[193];
    assign layer0_outputs[77] = inputs[92];
    assign layer0_outputs[78] = ~(inputs[248]) | (inputs[235]);
    assign layer0_outputs[79] = (inputs[228]) | (inputs[128]);
    assign layer0_outputs[80] = ~(inputs[11]);
    assign layer0_outputs[81] = ~(inputs[95]);
    assign layer0_outputs[82] = inputs[153];
    assign layer0_outputs[83] = ~((inputs[108]) ^ (inputs[103]));
    assign layer0_outputs[84] = ~((inputs[155]) ^ (inputs[124]));
    assign layer0_outputs[85] = ~((inputs[19]) | (inputs[33]));
    assign layer0_outputs[86] = ~(inputs[109]);
    assign layer0_outputs[87] = (inputs[251]) & ~(inputs[72]);
    assign layer0_outputs[88] = (inputs[61]) | (inputs[89]);
    assign layer0_outputs[89] = (inputs[62]) | (inputs[54]);
    assign layer0_outputs[90] = (inputs[139]) | (inputs[252]);
    assign layer0_outputs[91] = 1'b1;
    assign layer0_outputs[92] = ~(inputs[49]);
    assign layer0_outputs[93] = ~((inputs[210]) | (inputs[0]));
    assign layer0_outputs[94] = (inputs[165]) ^ (inputs[177]);
    assign layer0_outputs[95] = ~((inputs[209]) | (inputs[21]));
    assign layer0_outputs[96] = (inputs[89]) ^ (inputs[153]);
    assign layer0_outputs[97] = (inputs[27]) & ~(inputs[191]);
    assign layer0_outputs[98] = ~(inputs[108]);
    assign layer0_outputs[99] = ~((inputs[99]) | (inputs[15]));
    assign layer0_outputs[100] = (inputs[116]) & (inputs[93]);
    assign layer0_outputs[101] = ~((inputs[39]) | (inputs[9]));
    assign layer0_outputs[102] = (inputs[26]) ^ (inputs[207]);
    assign layer0_outputs[103] = inputs[247];
    assign layer0_outputs[104] = ~((inputs[52]) ^ (inputs[114]));
    assign layer0_outputs[105] = ~((inputs[111]) | (inputs[50]));
    assign layer0_outputs[106] = ~((inputs[238]) | (inputs[72]));
    assign layer0_outputs[107] = ~(inputs[97]);
    assign layer0_outputs[108] = (inputs[12]) ^ (inputs[141]);
    assign layer0_outputs[109] = ~(inputs[170]) | (inputs[151]);
    assign layer0_outputs[110] = inputs[217];
    assign layer0_outputs[111] = inputs[230];
    assign layer0_outputs[112] = inputs[166];
    assign layer0_outputs[113] = ~(inputs[245]) | (inputs[153]);
    assign layer0_outputs[114] = (inputs[28]) | (inputs[73]);
    assign layer0_outputs[115] = (inputs[137]) & ~(inputs[158]);
    assign layer0_outputs[116] = inputs[44];
    assign layer0_outputs[117] = ~(inputs[99]) | (inputs[27]);
    assign layer0_outputs[118] = inputs[114];
    assign layer0_outputs[119] = ~((inputs[165]) | (inputs[253]));
    assign layer0_outputs[120] = (inputs[21]) ^ (inputs[85]);
    assign layer0_outputs[121] = (inputs[51]) & ~(inputs[191]);
    assign layer0_outputs[122] = ~(inputs[42]) | (inputs[157]);
    assign layer0_outputs[123] = (inputs[120]) & ~(inputs[95]);
    assign layer0_outputs[124] = ~((inputs[125]) ^ (inputs[122]));
    assign layer0_outputs[125] = inputs[224];
    assign layer0_outputs[126] = ~(inputs[98]) | (inputs[190]);
    assign layer0_outputs[127] = ~((inputs[207]) ^ (inputs[60]));
    assign layer0_outputs[128] = (inputs[235]) ^ (inputs[124]);
    assign layer0_outputs[129] = (inputs[3]) | (inputs[136]);
    assign layer0_outputs[130] = 1'b0;
    assign layer0_outputs[131] = ~(inputs[125]);
    assign layer0_outputs[132] = ~((inputs[42]) | (inputs[4]));
    assign layer0_outputs[133] = ~((inputs[66]) | (inputs[204]));
    assign layer0_outputs[134] = ~((inputs[51]) & (inputs[102]));
    assign layer0_outputs[135] = ~(inputs[152]) | (inputs[159]);
    assign layer0_outputs[136] = ~(inputs[179]);
    assign layer0_outputs[137] = (inputs[62]) & ~(inputs[117]);
    assign layer0_outputs[138] = inputs[132];
    assign layer0_outputs[139] = ~((inputs[204]) ^ (inputs[124]));
    assign layer0_outputs[140] = ~((inputs[48]) | (inputs[167]));
    assign layer0_outputs[141] = ~((inputs[42]) ^ (inputs[102]));
    assign layer0_outputs[142] = ~((inputs[244]) ^ (inputs[250]));
    assign layer0_outputs[143] = ~(inputs[166]);
    assign layer0_outputs[144] = (inputs[38]) & ~(inputs[235]);
    assign layer0_outputs[145] = ~((inputs[129]) ^ (inputs[39]));
    assign layer0_outputs[146] = inputs[73];
    assign layer0_outputs[147] = (inputs[213]) ^ (inputs[38]);
    assign layer0_outputs[148] = inputs[185];
    assign layer0_outputs[149] = inputs[140];
    assign layer0_outputs[150] = ~(inputs[175]);
    assign layer0_outputs[151] = ~((inputs[25]) | (inputs[49]));
    assign layer0_outputs[152] = ~(inputs[43]) | (inputs[46]);
    assign layer0_outputs[153] = ~(inputs[138]);
    assign layer0_outputs[154] = ~(inputs[206]) | (inputs[174]);
    assign layer0_outputs[155] = (inputs[248]) | (inputs[144]);
    assign layer0_outputs[156] = ~((inputs[85]) ^ (inputs[145]));
    assign layer0_outputs[157] = ~(inputs[170]) | (inputs[44]);
    assign layer0_outputs[158] = 1'b0;
    assign layer0_outputs[159] = (inputs[180]) & (inputs[70]);
    assign layer0_outputs[160] = ~(inputs[245]) | (inputs[150]);
    assign layer0_outputs[161] = inputs[21];
    assign layer0_outputs[162] = (inputs[153]) & ~(inputs[193]);
    assign layer0_outputs[163] = inputs[67];
    assign layer0_outputs[164] = ~((inputs[147]) | (inputs[152]));
    assign layer0_outputs[165] = ~((inputs[242]) ^ (inputs[179]));
    assign layer0_outputs[166] = ~((inputs[212]) | (inputs[60]));
    assign layer0_outputs[167] = inputs[213];
    assign layer0_outputs[168] = (inputs[60]) | (inputs[192]);
    assign layer0_outputs[169] = ~(inputs[106]);
    assign layer0_outputs[170] = ~((inputs[16]) | (inputs[40]));
    assign layer0_outputs[171] = (inputs[125]) & (inputs[123]);
    assign layer0_outputs[172] = (inputs[237]) | (inputs[160]);
    assign layer0_outputs[173] = inputs[128];
    assign layer0_outputs[174] = (inputs[225]) & ~(inputs[79]);
    assign layer0_outputs[175] = (inputs[130]) | (inputs[237]);
    assign layer0_outputs[176] = inputs[41];
    assign layer0_outputs[177] = ~((inputs[185]) | (inputs[144]));
    assign layer0_outputs[178] = 1'b0;
    assign layer0_outputs[179] = (inputs[104]) & (inputs[33]);
    assign layer0_outputs[180] = ~(inputs[254]) | (inputs[156]);
    assign layer0_outputs[181] = (inputs[155]) ^ (inputs[148]);
    assign layer0_outputs[182] = inputs[132];
    assign layer0_outputs[183] = (inputs[214]) | (inputs[129]);
    assign layer0_outputs[184] = ~((inputs[64]) | (inputs[180]));
    assign layer0_outputs[185] = ~(inputs[178]);
    assign layer0_outputs[186] = ~((inputs[145]) | (inputs[80]));
    assign layer0_outputs[187] = inputs[120];
    assign layer0_outputs[188] = (inputs[213]) & ~(inputs[53]);
    assign layer0_outputs[189] = inputs[122];
    assign layer0_outputs[190] = (inputs[90]) | (inputs[21]);
    assign layer0_outputs[191] = (inputs[222]) & ~(inputs[206]);
    assign layer0_outputs[192] = (inputs[102]) | (inputs[43]);
    assign layer0_outputs[193] = inputs[117];
    assign layer0_outputs[194] = ~((inputs[158]) | (inputs[47]));
    assign layer0_outputs[195] = ~((inputs[45]) | (inputs[110]));
    assign layer0_outputs[196] = (inputs[37]) | (inputs[22]);
    assign layer0_outputs[197] = ~((inputs[66]) | (inputs[14]));
    assign layer0_outputs[198] = ~((inputs[50]) ^ (inputs[221]));
    assign layer0_outputs[199] = ~(inputs[84]);
    assign layer0_outputs[200] = ~(inputs[8]) | (inputs[39]);
    assign layer0_outputs[201] = inputs[214];
    assign layer0_outputs[202] = ~((inputs[199]) ^ (inputs[200]));
    assign layer0_outputs[203] = inputs[152];
    assign layer0_outputs[204] = inputs[214];
    assign layer0_outputs[205] = ~(inputs[56]) | (inputs[81]);
    assign layer0_outputs[206] = ~((inputs[152]) ^ (inputs[201]));
    assign layer0_outputs[207] = (inputs[179]) ^ (inputs[35]);
    assign layer0_outputs[208] = ~((inputs[134]) | (inputs[122]));
    assign layer0_outputs[209] = ~((inputs[121]) | (inputs[192]));
    assign layer0_outputs[210] = (inputs[231]) ^ (inputs[152]);
    assign layer0_outputs[211] = 1'b0;
    assign layer0_outputs[212] = (inputs[146]) | (inputs[196]);
    assign layer0_outputs[213] = ~(inputs[242]);
    assign layer0_outputs[214] = (inputs[231]) & ~(inputs[64]);
    assign layer0_outputs[215] = (inputs[125]) & ~(inputs[198]);
    assign layer0_outputs[216] = ~(inputs[237]);
    assign layer0_outputs[217] = 1'b1;
    assign layer0_outputs[218] = (inputs[154]) & (inputs[160]);
    assign layer0_outputs[219] = ~((inputs[49]) | (inputs[254]));
    assign layer0_outputs[220] = 1'b0;
    assign layer0_outputs[221] = ~(inputs[92]);
    assign layer0_outputs[222] = ~((inputs[44]) ^ (inputs[231]));
    assign layer0_outputs[223] = ~((inputs[129]) ^ (inputs[185]));
    assign layer0_outputs[224] = (inputs[42]) | (inputs[208]);
    assign layer0_outputs[225] = (inputs[13]) | (inputs[237]);
    assign layer0_outputs[226] = (inputs[182]) ^ (inputs[138]);
    assign layer0_outputs[227] = ~(inputs[218]) | (inputs[31]);
    assign layer0_outputs[228] = (inputs[220]) & ~(inputs[97]);
    assign layer0_outputs[229] = (inputs[143]) | (inputs[223]);
    assign layer0_outputs[230] = inputs[213];
    assign layer0_outputs[231] = (inputs[62]) & ~(inputs[139]);
    assign layer0_outputs[232] = (inputs[167]) & ~(inputs[211]);
    assign layer0_outputs[233] = (inputs[121]) & (inputs[153]);
    assign layer0_outputs[234] = ~((inputs[59]) | (inputs[4]));
    assign layer0_outputs[235] = ~(inputs[244]) | (inputs[168]);
    assign layer0_outputs[236] = (inputs[163]) | (inputs[206]);
    assign layer0_outputs[237] = ~(inputs[56]) | (inputs[50]);
    assign layer0_outputs[238] = ~((inputs[117]) ^ (inputs[174]));
    assign layer0_outputs[239] = 1'b1;
    assign layer0_outputs[240] = ~(inputs[3]);
    assign layer0_outputs[241] = inputs[72];
    assign layer0_outputs[242] = inputs[174];
    assign layer0_outputs[243] = (inputs[94]) ^ (inputs[187]);
    assign layer0_outputs[244] = ~((inputs[213]) | (inputs[229]));
    assign layer0_outputs[245] = ~((inputs[161]) ^ (inputs[130]));
    assign layer0_outputs[246] = (inputs[193]) | (inputs[210]);
    assign layer0_outputs[247] = ~((inputs[144]) | (inputs[220]));
    assign layer0_outputs[248] = ~((inputs[36]) | (inputs[167]));
    assign layer0_outputs[249] = inputs[21];
    assign layer0_outputs[250] = (inputs[70]) ^ (inputs[90]);
    assign layer0_outputs[251] = ~(inputs[40]) | (inputs[217]);
    assign layer0_outputs[252] = ~(inputs[224]) | (inputs[19]);
    assign layer0_outputs[253] = ~((inputs[124]) | (inputs[96]));
    assign layer0_outputs[254] = ~((inputs[216]) ^ (inputs[148]));
    assign layer0_outputs[255] = (inputs[226]) | (inputs[233]);
    assign layer0_outputs[256] = (inputs[215]) & ~(inputs[46]);
    assign layer0_outputs[257] = ~((inputs[65]) ^ (inputs[204]));
    assign layer0_outputs[258] = inputs[84];
    assign layer0_outputs[259] = (inputs[230]) & ~(inputs[121]);
    assign layer0_outputs[260] = (inputs[159]) ^ (inputs[218]);
    assign layer0_outputs[261] = inputs[200];
    assign layer0_outputs[262] = inputs[122];
    assign layer0_outputs[263] = (inputs[69]) ^ (inputs[81]);
    assign layer0_outputs[264] = ~(inputs[114]) | (inputs[233]);
    assign layer0_outputs[265] = inputs[18];
    assign layer0_outputs[266] = ~((inputs[31]) | (inputs[234]));
    assign layer0_outputs[267] = (inputs[141]) ^ (inputs[29]);
    assign layer0_outputs[268] = inputs[252];
    assign layer0_outputs[269] = inputs[90];
    assign layer0_outputs[270] = ~(inputs[60]);
    assign layer0_outputs[271] = ~(inputs[226]);
    assign layer0_outputs[272] = ~((inputs[111]) ^ (inputs[88]));
    assign layer0_outputs[273] = inputs[194];
    assign layer0_outputs[274] = ~(inputs[90]);
    assign layer0_outputs[275] = ~(inputs[233]);
    assign layer0_outputs[276] = ~(inputs[17]) | (inputs[175]);
    assign layer0_outputs[277] = ~((inputs[3]) | (inputs[3]));
    assign layer0_outputs[278] = inputs[50];
    assign layer0_outputs[279] = 1'b0;
    assign layer0_outputs[280] = ~(inputs[22]) | (inputs[161]);
    assign layer0_outputs[281] = inputs[27];
    assign layer0_outputs[282] = inputs[8];
    assign layer0_outputs[283] = ~((inputs[55]) ^ (inputs[8]));
    assign layer0_outputs[284] = ~(inputs[118]);
    assign layer0_outputs[285] = (inputs[238]) & (inputs[140]);
    assign layer0_outputs[286] = (inputs[4]) | (inputs[188]);
    assign layer0_outputs[287] = ~(inputs[193]) | (inputs[71]);
    assign layer0_outputs[288] = 1'b0;
    assign layer0_outputs[289] = ~(inputs[250]) | (inputs[185]);
    assign layer0_outputs[290] = ~(inputs[126]) | (inputs[93]);
    assign layer0_outputs[291] = ~(inputs[187]) | (inputs[134]);
    assign layer0_outputs[292] = inputs[40];
    assign layer0_outputs[293] = ~(inputs[38]);
    assign layer0_outputs[294] = (inputs[102]) ^ (inputs[52]);
    assign layer0_outputs[295] = ~(inputs[14]);
    assign layer0_outputs[296] = ~((inputs[158]) ^ (inputs[218]));
    assign layer0_outputs[297] = (inputs[144]) ^ (inputs[198]);
    assign layer0_outputs[298] = ~(inputs[36]);
    assign layer0_outputs[299] = ~((inputs[99]) ^ (inputs[82]));
    assign layer0_outputs[300] = ~((inputs[24]) | (inputs[211]));
    assign layer0_outputs[301] = (inputs[226]) | (inputs[207]);
    assign layer0_outputs[302] = ~((inputs[221]) | (inputs[212]));
    assign layer0_outputs[303] = inputs[31];
    assign layer0_outputs[304] = ~((inputs[172]) | (inputs[215]));
    assign layer0_outputs[305] = ~(inputs[202]);
    assign layer0_outputs[306] = ~(inputs[167]) | (inputs[79]);
    assign layer0_outputs[307] = ~((inputs[244]) | (inputs[172]));
    assign layer0_outputs[308] = inputs[241];
    assign layer0_outputs[309] = inputs[121];
    assign layer0_outputs[310] = (inputs[5]) | (inputs[78]);
    assign layer0_outputs[311] = (inputs[231]) & ~(inputs[31]);
    assign layer0_outputs[312] = (inputs[88]) & ~(inputs[224]);
    assign layer0_outputs[313] = inputs[15];
    assign layer0_outputs[314] = (inputs[191]) ^ (inputs[183]);
    assign layer0_outputs[315] = (inputs[102]) & ~(inputs[125]);
    assign layer0_outputs[316] = ~(inputs[153]);
    assign layer0_outputs[317] = (inputs[111]) | (inputs[94]);
    assign layer0_outputs[318] = (inputs[29]) | (inputs[16]);
    assign layer0_outputs[319] = ~(inputs[116]);
    assign layer0_outputs[320] = (inputs[124]) | (inputs[4]);
    assign layer0_outputs[321] = ~(inputs[178]);
    assign layer0_outputs[322] = ~(inputs[177]);
    assign layer0_outputs[323] = inputs[33];
    assign layer0_outputs[324] = inputs[105];
    assign layer0_outputs[325] = ~((inputs[39]) | (inputs[48]));
    assign layer0_outputs[326] = inputs[213];
    assign layer0_outputs[327] = ~(inputs[86]) | (inputs[188]);
    assign layer0_outputs[328] = ~(inputs[21]);
    assign layer0_outputs[329] = (inputs[117]) ^ (inputs[221]);
    assign layer0_outputs[330] = (inputs[5]) ^ (inputs[70]);
    assign layer0_outputs[331] = ~((inputs[1]) | (inputs[120]));
    assign layer0_outputs[332] = ~((inputs[143]) | (inputs[243]));
    assign layer0_outputs[333] = (inputs[71]) & ~(inputs[18]);
    assign layer0_outputs[334] = ~((inputs[98]) ^ (inputs[81]));
    assign layer0_outputs[335] = (inputs[74]) | (inputs[129]);
    assign layer0_outputs[336] = (inputs[168]) | (inputs[253]);
    assign layer0_outputs[337] = (inputs[18]) | (inputs[34]);
    assign layer0_outputs[338] = (inputs[132]) & ~(inputs[227]);
    assign layer0_outputs[339] = (inputs[144]) ^ (inputs[181]);
    assign layer0_outputs[340] = 1'b0;
    assign layer0_outputs[341] = inputs[128];
    assign layer0_outputs[342] = ~(inputs[202]);
    assign layer0_outputs[343] = inputs[100];
    assign layer0_outputs[344] = ~((inputs[119]) & (inputs[9]));
    assign layer0_outputs[345] = (inputs[217]) & ~(inputs[235]);
    assign layer0_outputs[346] = ~(inputs[85]);
    assign layer0_outputs[347] = (inputs[239]) | (inputs[238]);
    assign layer0_outputs[348] = inputs[49];
    assign layer0_outputs[349] = (inputs[84]) | (inputs[45]);
    assign layer0_outputs[350] = inputs[105];
    assign layer0_outputs[351] = ~(inputs[254]) | (inputs[252]);
    assign layer0_outputs[352] = (inputs[105]) & ~(inputs[34]);
    assign layer0_outputs[353] = (inputs[8]) & ~(inputs[244]);
    assign layer0_outputs[354] = ~((inputs[59]) ^ (inputs[33]));
    assign layer0_outputs[355] = ~((inputs[137]) | (inputs[153]));
    assign layer0_outputs[356] = ~(inputs[129]) | (inputs[102]);
    assign layer0_outputs[357] = ~((inputs[122]) ^ (inputs[157]));
    assign layer0_outputs[358] = (inputs[225]) | (inputs[197]);
    assign layer0_outputs[359] = inputs[132];
    assign layer0_outputs[360] = ~((inputs[24]) & (inputs[72]));
    assign layer0_outputs[361] = ~(inputs[57]);
    assign layer0_outputs[362] = ~((inputs[211]) | (inputs[188]));
    assign layer0_outputs[363] = ~(inputs[58]);
    assign layer0_outputs[364] = ~((inputs[68]) ^ (inputs[80]));
    assign layer0_outputs[365] = ~(inputs[84]);
    assign layer0_outputs[366] = ~((inputs[234]) ^ (inputs[206]));
    assign layer0_outputs[367] = ~(inputs[73]);
    assign layer0_outputs[368] = inputs[192];
    assign layer0_outputs[369] = ~(inputs[82]);
    assign layer0_outputs[370] = ~(inputs[227]);
    assign layer0_outputs[371] = (inputs[206]) | (inputs[109]);
    assign layer0_outputs[372] = inputs[50];
    assign layer0_outputs[373] = ~((inputs[193]) ^ (inputs[58]));
    assign layer0_outputs[374] = (inputs[156]) & ~(inputs[252]);
    assign layer0_outputs[375] = ~((inputs[197]) | (inputs[82]));
    assign layer0_outputs[376] = (inputs[182]) | (inputs[34]);
    assign layer0_outputs[377] = ~(inputs[174]);
    assign layer0_outputs[378] = ~((inputs[24]) ^ (inputs[191]));
    assign layer0_outputs[379] = ~(inputs[83]) | (inputs[65]);
    assign layer0_outputs[380] = (inputs[61]) & ~(inputs[113]);
    assign layer0_outputs[381] = ~((inputs[21]) ^ (inputs[142]));
    assign layer0_outputs[382] = (inputs[136]) & ~(inputs[202]);
    assign layer0_outputs[383] = inputs[110];
    assign layer0_outputs[384] = ~(inputs[77]);
    assign layer0_outputs[385] = inputs[150];
    assign layer0_outputs[386] = ~(inputs[26]) | (inputs[216]);
    assign layer0_outputs[387] = ~((inputs[108]) ^ (inputs[111]));
    assign layer0_outputs[388] = ~((inputs[18]) | (inputs[152]));
    assign layer0_outputs[389] = ~((inputs[255]) | (inputs[192]));
    assign layer0_outputs[390] = ~(inputs[210]);
    assign layer0_outputs[391] = (inputs[31]) & (inputs[211]);
    assign layer0_outputs[392] = ~(inputs[155]) | (inputs[131]);
    assign layer0_outputs[393] = ~((inputs[133]) & (inputs[68]));
    assign layer0_outputs[394] = (inputs[39]) & ~(inputs[161]);
    assign layer0_outputs[395] = ~(inputs[111]) | (inputs[253]);
    assign layer0_outputs[396] = ~((inputs[126]) | (inputs[179]));
    assign layer0_outputs[397] = ~((inputs[20]) ^ (inputs[159]));
    assign layer0_outputs[398] = inputs[189];
    assign layer0_outputs[399] = inputs[165];
    assign layer0_outputs[400] = ~((inputs[99]) | (inputs[3]));
    assign layer0_outputs[401] = ~(inputs[53]);
    assign layer0_outputs[402] = (inputs[38]) & (inputs[69]);
    assign layer0_outputs[403] = ~((inputs[87]) ^ (inputs[60]));
    assign layer0_outputs[404] = (inputs[136]) | (inputs[43]);
    assign layer0_outputs[405] = (inputs[234]) & ~(inputs[126]);
    assign layer0_outputs[406] = ~(inputs[104]);
    assign layer0_outputs[407] = ~(inputs[132]);
    assign layer0_outputs[408] = ~((inputs[168]) | (inputs[236]));
    assign layer0_outputs[409] = ~((inputs[8]) & (inputs[133]));
    assign layer0_outputs[410] = ~((inputs[183]) | (inputs[63]));
    assign layer0_outputs[411] = ~(inputs[116]);
    assign layer0_outputs[412] = 1'b0;
    assign layer0_outputs[413] = 1'b1;
    assign layer0_outputs[414] = (inputs[160]) | (inputs[179]);
    assign layer0_outputs[415] = ~((inputs[251]) | (inputs[185]));
    assign layer0_outputs[416] = (inputs[40]) | (inputs[109]);
    assign layer0_outputs[417] = ~((inputs[113]) ^ (inputs[16]));
    assign layer0_outputs[418] = ~((inputs[174]) & (inputs[159]));
    assign layer0_outputs[419] = ~(inputs[150]);
    assign layer0_outputs[420] = (inputs[209]) & ~(inputs[205]);
    assign layer0_outputs[421] = ~((inputs[104]) | (inputs[208]));
    assign layer0_outputs[422] = ~(inputs[53]) | (inputs[190]);
    assign layer0_outputs[423] = ~((inputs[135]) ^ (inputs[194]));
    assign layer0_outputs[424] = (inputs[70]) ^ (inputs[33]);
    assign layer0_outputs[425] = ~((inputs[198]) | (inputs[185]));
    assign layer0_outputs[426] = ~(inputs[120]);
    assign layer0_outputs[427] = (inputs[183]) & (inputs[108]);
    assign layer0_outputs[428] = (inputs[180]) & ~(inputs[74]);
    assign layer0_outputs[429] = ~((inputs[187]) ^ (inputs[241]));
    assign layer0_outputs[430] = (inputs[178]) & ~(inputs[43]);
    assign layer0_outputs[431] = (inputs[165]) ^ (inputs[146]);
    assign layer0_outputs[432] = ~(inputs[83]) | (inputs[72]);
    assign layer0_outputs[433] = (inputs[44]) & ~(inputs[15]);
    assign layer0_outputs[434] = (inputs[140]) & (inputs[139]);
    assign layer0_outputs[435] = ~((inputs[131]) ^ (inputs[100]));
    assign layer0_outputs[436] = ~((inputs[216]) & (inputs[187]));
    assign layer0_outputs[437] = (inputs[214]) & ~(inputs[96]);
    assign layer0_outputs[438] = ~(inputs[252]);
    assign layer0_outputs[439] = ~(inputs[245]) | (inputs[15]);
    assign layer0_outputs[440] = (inputs[72]) & (inputs[44]);
    assign layer0_outputs[441] = ~((inputs[60]) | (inputs[130]));
    assign layer0_outputs[442] = (inputs[173]) | (inputs[80]);
    assign layer0_outputs[443] = inputs[154];
    assign layer0_outputs[444] = ~((inputs[143]) | (inputs[225]));
    assign layer0_outputs[445] = ~((inputs[213]) | (inputs[37]));
    assign layer0_outputs[446] = ~((inputs[184]) & (inputs[201]));
    assign layer0_outputs[447] = ~(inputs[188]);
    assign layer0_outputs[448] = ~((inputs[2]) & (inputs[175]));
    assign layer0_outputs[449] = (inputs[10]) | (inputs[0]);
    assign layer0_outputs[450] = ~(inputs[93]);
    assign layer0_outputs[451] = 1'b1;
    assign layer0_outputs[452] = (inputs[61]) & (inputs[20]);
    assign layer0_outputs[453] = ~((inputs[132]) | (inputs[186]));
    assign layer0_outputs[454] = inputs[171];
    assign layer0_outputs[455] = ~((inputs[177]) | (inputs[194]));
    assign layer0_outputs[456] = ~(inputs[145]) | (inputs[57]);
    assign layer0_outputs[457] = ~(inputs[228]);
    assign layer0_outputs[458] = inputs[30];
    assign layer0_outputs[459] = ~(inputs[120]);
    assign layer0_outputs[460] = inputs[180];
    assign layer0_outputs[461] = ~((inputs[133]) | (inputs[101]));
    assign layer0_outputs[462] = ~((inputs[207]) | (inputs[220]));
    assign layer0_outputs[463] = ~((inputs[142]) | (inputs[79]));
    assign layer0_outputs[464] = (inputs[106]) ^ (inputs[232]);
    assign layer0_outputs[465] = inputs[100];
    assign layer0_outputs[466] = inputs[25];
    assign layer0_outputs[467] = (inputs[70]) ^ (inputs[65]);
    assign layer0_outputs[468] = ~((inputs[223]) | (inputs[5]));
    assign layer0_outputs[469] = inputs[215];
    assign layer0_outputs[470] = inputs[22];
    assign layer0_outputs[471] = ~(inputs[221]);
    assign layer0_outputs[472] = ~((inputs[191]) | (inputs[176]));
    assign layer0_outputs[473] = inputs[34];
    assign layer0_outputs[474] = ~(inputs[213]);
    assign layer0_outputs[475] = ~(inputs[132]) | (inputs[48]);
    assign layer0_outputs[476] = ~((inputs[82]) | (inputs[111]));
    assign layer0_outputs[477] = ~(inputs[217]);
    assign layer0_outputs[478] = inputs[233];
    assign layer0_outputs[479] = ~((inputs[9]) ^ (inputs[4]));
    assign layer0_outputs[480] = ~((inputs[161]) ^ (inputs[245]));
    assign layer0_outputs[481] = (inputs[244]) & (inputs[55]);
    assign layer0_outputs[482] = (inputs[245]) & ~(inputs[48]);
    assign layer0_outputs[483] = ~((inputs[225]) | (inputs[64]));
    assign layer0_outputs[484] = (inputs[227]) & ~(inputs[20]);
    assign layer0_outputs[485] = inputs[89];
    assign layer0_outputs[486] = (inputs[22]) | (inputs[123]);
    assign layer0_outputs[487] = ~(inputs[153]);
    assign layer0_outputs[488] = ~(inputs[152]);
    assign layer0_outputs[489] = 1'b1;
    assign layer0_outputs[490] = ~((inputs[147]) | (inputs[232]));
    assign layer0_outputs[491] = inputs[68];
    assign layer0_outputs[492] = ~((inputs[230]) | (inputs[228]));
    assign layer0_outputs[493] = ~((inputs[144]) ^ (inputs[81]));
    assign layer0_outputs[494] = (inputs[103]) & ~(inputs[199]);
    assign layer0_outputs[495] = (inputs[245]) & (inputs[11]);
    assign layer0_outputs[496] = ~(inputs[123]);
    assign layer0_outputs[497] = (inputs[107]) & ~(inputs[235]);
    assign layer0_outputs[498] = ~(inputs[210]) | (inputs[48]);
    assign layer0_outputs[499] = inputs[24];
    assign layer0_outputs[500] = ~((inputs[47]) ^ (inputs[238]));
    assign layer0_outputs[501] = ~((inputs[87]) ^ (inputs[115]));
    assign layer0_outputs[502] = ~((inputs[135]) ^ (inputs[36]));
    assign layer0_outputs[503] = inputs[165];
    assign layer0_outputs[504] = inputs[215];
    assign layer0_outputs[505] = ~(inputs[6]) | (inputs[214]);
    assign layer0_outputs[506] = ~(inputs[89]);
    assign layer0_outputs[507] = 1'b1;
    assign layer0_outputs[508] = (inputs[176]) ^ (inputs[144]);
    assign layer0_outputs[509] = inputs[152];
    assign layer0_outputs[510] = (inputs[170]) & ~(inputs[249]);
    assign layer0_outputs[511] = (inputs[112]) ^ (inputs[219]);
    assign layer0_outputs[512] = ~(inputs[19]);
    assign layer0_outputs[513] = inputs[90];
    assign layer0_outputs[514] = (inputs[252]) & (inputs[159]);
    assign layer0_outputs[515] = ~(inputs[242]);
    assign layer0_outputs[516] = (inputs[17]) & ~(inputs[175]);
    assign layer0_outputs[517] = (inputs[249]) | (inputs[94]);
    assign layer0_outputs[518] = ~(inputs[70]) | (inputs[173]);
    assign layer0_outputs[519] = ~(inputs[163]);
    assign layer0_outputs[520] = ~(inputs[231]);
    assign layer0_outputs[521] = (inputs[145]) | (inputs[91]);
    assign layer0_outputs[522] = (inputs[76]) & ~(inputs[30]);
    assign layer0_outputs[523] = ~((inputs[233]) ^ (inputs[168]));
    assign layer0_outputs[524] = (inputs[170]) ^ (inputs[122]);
    assign layer0_outputs[525] = ~(inputs[3]) | (inputs[161]);
    assign layer0_outputs[526] = (inputs[136]) & ~(inputs[64]);
    assign layer0_outputs[527] = ~((inputs[79]) ^ (inputs[91]));
    assign layer0_outputs[528] = (inputs[189]) | (inputs[130]);
    assign layer0_outputs[529] = (inputs[148]) & ~(inputs[202]);
    assign layer0_outputs[530] = ~((inputs[147]) ^ (inputs[67]));
    assign layer0_outputs[531] = ~(inputs[73]);
    assign layer0_outputs[532] = ~(inputs[125]);
    assign layer0_outputs[533] = ~(inputs[0]);
    assign layer0_outputs[534] = inputs[215];
    assign layer0_outputs[535] = inputs[130];
    assign layer0_outputs[536] = (inputs[154]) | (inputs[45]);
    assign layer0_outputs[537] = ~((inputs[178]) | (inputs[207]));
    assign layer0_outputs[538] = (inputs[40]) | (inputs[116]);
    assign layer0_outputs[539] = ~(inputs[31]);
    assign layer0_outputs[540] = ~((inputs[141]) | (inputs[26]));
    assign layer0_outputs[541] = ~((inputs[210]) | (inputs[95]));
    assign layer0_outputs[542] = (inputs[78]) & ~(inputs[2]);
    assign layer0_outputs[543] = ~((inputs[167]) | (inputs[151]));
    assign layer0_outputs[544] = inputs[200];
    assign layer0_outputs[545] = ~((inputs[237]) | (inputs[29]));
    assign layer0_outputs[546] = (inputs[150]) & ~(inputs[99]);
    assign layer0_outputs[547] = inputs[141];
    assign layer0_outputs[548] = ~(inputs[200]);
    assign layer0_outputs[549] = ~(inputs[20]);
    assign layer0_outputs[550] = ~(inputs[187]);
    assign layer0_outputs[551] = (inputs[129]) ^ (inputs[83]);
    assign layer0_outputs[552] = ~((inputs[155]) | (inputs[84]));
    assign layer0_outputs[553] = (inputs[186]) & ~(inputs[3]);
    assign layer0_outputs[554] = (inputs[216]) & ~(inputs[105]);
    assign layer0_outputs[555] = (inputs[167]) & ~(inputs[5]);
    assign layer0_outputs[556] = (inputs[1]) & ~(inputs[4]);
    assign layer0_outputs[557] = 1'b0;
    assign layer0_outputs[558] = (inputs[25]) & ~(inputs[225]);
    assign layer0_outputs[559] = (inputs[8]) ^ (inputs[47]);
    assign layer0_outputs[560] = ~((inputs[216]) | (inputs[171]));
    assign layer0_outputs[561] = inputs[131];
    assign layer0_outputs[562] = (inputs[176]) | (inputs[60]);
    assign layer0_outputs[563] = inputs[42];
    assign layer0_outputs[564] = ~(inputs[182]);
    assign layer0_outputs[565] = (inputs[80]) | (inputs[172]);
    assign layer0_outputs[566] = ~(inputs[122]);
    assign layer0_outputs[567] = inputs[47];
    assign layer0_outputs[568] = ~(inputs[198]) | (inputs[192]);
    assign layer0_outputs[569] = ~(inputs[153]) | (inputs[118]);
    assign layer0_outputs[570] = ~((inputs[50]) & (inputs[89]));
    assign layer0_outputs[571] = inputs[38];
    assign layer0_outputs[572] = (inputs[239]) ^ (inputs[132]);
    assign layer0_outputs[573] = ~(inputs[21]) | (inputs[29]);
    assign layer0_outputs[574] = ~((inputs[100]) ^ (inputs[147]));
    assign layer0_outputs[575] = ~(inputs[37]);
    assign layer0_outputs[576] = (inputs[177]) | (inputs[165]);
    assign layer0_outputs[577] = inputs[85];
    assign layer0_outputs[578] = (inputs[84]) & ~(inputs[109]);
    assign layer0_outputs[579] = inputs[205];
    assign layer0_outputs[580] = ~(inputs[100]);
    assign layer0_outputs[581] = ~(inputs[104]) | (inputs[176]);
    assign layer0_outputs[582] = ~((inputs[65]) | (inputs[87]));
    assign layer0_outputs[583] = ~(inputs[21]);
    assign layer0_outputs[584] = inputs[113];
    assign layer0_outputs[585] = (inputs[247]) ^ (inputs[58]);
    assign layer0_outputs[586] = ~((inputs[0]) | (inputs[215]));
    assign layer0_outputs[587] = (inputs[15]) & ~(inputs[137]);
    assign layer0_outputs[588] = ~((inputs[171]) & (inputs[195]));
    assign layer0_outputs[589] = (inputs[44]) | (inputs[6]);
    assign layer0_outputs[590] = inputs[16];
    assign layer0_outputs[591] = ~(inputs[74]) | (inputs[236]);
    assign layer0_outputs[592] = (inputs[59]) & ~(inputs[71]);
    assign layer0_outputs[593] = ~(inputs[247]);
    assign layer0_outputs[594] = inputs[53];
    assign layer0_outputs[595] = inputs[6];
    assign layer0_outputs[596] = inputs[168];
    assign layer0_outputs[597] = ~(inputs[78]);
    assign layer0_outputs[598] = ~((inputs[249]) | (inputs[18]));
    assign layer0_outputs[599] = inputs[145];
    assign layer0_outputs[600] = (inputs[140]) & ~(inputs[50]);
    assign layer0_outputs[601] = (inputs[230]) & ~(inputs[75]);
    assign layer0_outputs[602] = ~(inputs[118]);
    assign layer0_outputs[603] = inputs[163];
    assign layer0_outputs[604] = ~(inputs[218]);
    assign layer0_outputs[605] = inputs[31];
    assign layer0_outputs[606] = inputs[161];
    assign layer0_outputs[607] = inputs[139];
    assign layer0_outputs[608] = (inputs[128]) & ~(inputs[143]);
    assign layer0_outputs[609] = (inputs[243]) ^ (inputs[216]);
    assign layer0_outputs[610] = ~(inputs[25]);
    assign layer0_outputs[611] = ~((inputs[72]) ^ (inputs[108]));
    assign layer0_outputs[612] = ~(inputs[131]);
    assign layer0_outputs[613] = inputs[114];
    assign layer0_outputs[614] = ~((inputs[129]) ^ (inputs[116]));
    assign layer0_outputs[615] = ~(inputs[87]);
    assign layer0_outputs[616] = (inputs[76]) | (inputs[192]);
    assign layer0_outputs[617] = inputs[108];
    assign layer0_outputs[618] = (inputs[191]) ^ (inputs[165]);
    assign layer0_outputs[619] = (inputs[169]) | (inputs[18]);
    assign layer0_outputs[620] = ~(inputs[195]);
    assign layer0_outputs[621] = ~(inputs[88]);
    assign layer0_outputs[622] = inputs[165];
    assign layer0_outputs[623] = (inputs[96]) | (inputs[95]);
    assign layer0_outputs[624] = ~(inputs[105]);
    assign layer0_outputs[625] = inputs[184];
    assign layer0_outputs[626] = (inputs[113]) | (inputs[111]);
    assign layer0_outputs[627] = ~((inputs[37]) | (inputs[52]));
    assign layer0_outputs[628] = (inputs[186]) & ~(inputs[97]);
    assign layer0_outputs[629] = inputs[128];
    assign layer0_outputs[630] = ~((inputs[51]) | (inputs[108]));
    assign layer0_outputs[631] = inputs[56];
    assign layer0_outputs[632] = ~((inputs[126]) ^ (inputs[199]));
    assign layer0_outputs[633] = (inputs[152]) & ~(inputs[211]);
    assign layer0_outputs[634] = ~(inputs[61]);
    assign layer0_outputs[635] = (inputs[166]) & ~(inputs[81]);
    assign layer0_outputs[636] = ~(inputs[86]);
    assign layer0_outputs[637] = (inputs[87]) ^ (inputs[43]);
    assign layer0_outputs[638] = (inputs[140]) ^ (inputs[204]);
    assign layer0_outputs[639] = ~((inputs[203]) ^ (inputs[104]));
    assign layer0_outputs[640] = ~(inputs[103]) | (inputs[125]);
    assign layer0_outputs[641] = (inputs[205]) & (inputs[185]);
    assign layer0_outputs[642] = (inputs[210]) ^ (inputs[92]);
    assign layer0_outputs[643] = (inputs[73]) | (inputs[140]);
    assign layer0_outputs[644] = ~(inputs[146]);
    assign layer0_outputs[645] = ~((inputs[64]) | (inputs[232]));
    assign layer0_outputs[646] = ~(inputs[218]);
    assign layer0_outputs[647] = inputs[98];
    assign layer0_outputs[648] = ~((inputs[28]) | (inputs[238]));
    assign layer0_outputs[649] = ~((inputs[57]) | (inputs[241]));
    assign layer0_outputs[650] = 1'b0;
    assign layer0_outputs[651] = inputs[6];
    assign layer0_outputs[652] = ~((inputs[222]) ^ (inputs[60]));
    assign layer0_outputs[653] = ~(inputs[91]);
    assign layer0_outputs[654] = ~((inputs[0]) | (inputs[40]));
    assign layer0_outputs[655] = (inputs[170]) ^ (inputs[191]);
    assign layer0_outputs[656] = ~(inputs[214]) | (inputs[131]);
    assign layer0_outputs[657] = ~((inputs[33]) | (inputs[187]));
    assign layer0_outputs[658] = ~((inputs[172]) | (inputs[222]));
    assign layer0_outputs[659] = ~((inputs[244]) ^ (inputs[36]));
    assign layer0_outputs[660] = ~(inputs[207]) | (inputs[81]);
    assign layer0_outputs[661] = (inputs[38]) | (inputs[255]);
    assign layer0_outputs[662] = (inputs[61]) | (inputs[58]);
    assign layer0_outputs[663] = ~(inputs[180]);
    assign layer0_outputs[664] = ~(inputs[146]);
    assign layer0_outputs[665] = inputs[162];
    assign layer0_outputs[666] = ~((inputs[177]) ^ (inputs[220]));
    assign layer0_outputs[667] = inputs[124];
    assign layer0_outputs[668] = inputs[164];
    assign layer0_outputs[669] = 1'b1;
    assign layer0_outputs[670] = (inputs[17]) ^ (inputs[135]);
    assign layer0_outputs[671] = (inputs[19]) ^ (inputs[253]);
    assign layer0_outputs[672] = (inputs[199]) | (inputs[184]);
    assign layer0_outputs[673] = ~((inputs[28]) | (inputs[95]));
    assign layer0_outputs[674] = (inputs[210]) | (inputs[247]);
    assign layer0_outputs[675] = (inputs[126]) & ~(inputs[246]);
    assign layer0_outputs[676] = inputs[51];
    assign layer0_outputs[677] = ~(inputs[151]);
    assign layer0_outputs[678] = (inputs[254]) ^ (inputs[99]);
    assign layer0_outputs[679] = ~(inputs[73]);
    assign layer0_outputs[680] = (inputs[75]) & ~(inputs[163]);
    assign layer0_outputs[681] = (inputs[106]) & ~(inputs[229]);
    assign layer0_outputs[682] = ~(inputs[18]);
    assign layer0_outputs[683] = ~((inputs[141]) | (inputs[157]));
    assign layer0_outputs[684] = ~((inputs[150]) ^ (inputs[80]));
    assign layer0_outputs[685] = inputs[228];
    assign layer0_outputs[686] = inputs[22];
    assign layer0_outputs[687] = (inputs[9]) | (inputs[116]);
    assign layer0_outputs[688] = (inputs[111]) | (inputs[97]);
    assign layer0_outputs[689] = (inputs[233]) & ~(inputs[64]);
    assign layer0_outputs[690] = inputs[128];
    assign layer0_outputs[691] = (inputs[183]) & ~(inputs[42]);
    assign layer0_outputs[692] = (inputs[112]) ^ (inputs[170]);
    assign layer0_outputs[693] = (inputs[52]) ^ (inputs[54]);
    assign layer0_outputs[694] = inputs[189];
    assign layer0_outputs[695] = ~(inputs[219]);
    assign layer0_outputs[696] = 1'b0;
    assign layer0_outputs[697] = ~((inputs[97]) ^ (inputs[159]));
    assign layer0_outputs[698] = (inputs[112]) & ~(inputs[32]);
    assign layer0_outputs[699] = (inputs[134]) & (inputs[94]);
    assign layer0_outputs[700] = (inputs[104]) ^ (inputs[3]);
    assign layer0_outputs[701] = (inputs[144]) ^ (inputs[168]);
    assign layer0_outputs[702] = (inputs[158]) | (inputs[73]);
    assign layer0_outputs[703] = (inputs[64]) & ~(inputs[59]);
    assign layer0_outputs[704] = inputs[133];
    assign layer0_outputs[705] = inputs[106];
    assign layer0_outputs[706] = (inputs[93]) ^ (inputs[153]);
    assign layer0_outputs[707] = (inputs[38]) | (inputs[54]);
    assign layer0_outputs[708] = (inputs[0]) | (inputs[63]);
    assign layer0_outputs[709] = ~((inputs[41]) ^ (inputs[160]));
    assign layer0_outputs[710] = ~((inputs[217]) ^ (inputs[41]));
    assign layer0_outputs[711] = (inputs[134]) & ~(inputs[72]);
    assign layer0_outputs[712] = (inputs[120]) & ~(inputs[219]);
    assign layer0_outputs[713] = ~((inputs[242]) | (inputs[103]));
    assign layer0_outputs[714] = (inputs[139]) & (inputs[75]);
    assign layer0_outputs[715] = ~(inputs[84]) | (inputs[157]);
    assign layer0_outputs[716] = inputs[44];
    assign layer0_outputs[717] = (inputs[127]) | (inputs[66]);
    assign layer0_outputs[718] = ~((inputs[110]) | (inputs[145]));
    assign layer0_outputs[719] = ~((inputs[156]) | (inputs[1]));
    assign layer0_outputs[720] = (inputs[226]) & ~(inputs[131]);
    assign layer0_outputs[721] = (inputs[145]) | (inputs[48]);
    assign layer0_outputs[722] = (inputs[237]) ^ (inputs[52]);
    assign layer0_outputs[723] = (inputs[65]) & (inputs[179]);
    assign layer0_outputs[724] = (inputs[25]) ^ (inputs[110]);
    assign layer0_outputs[725] = (inputs[45]) ^ (inputs[81]);
    assign layer0_outputs[726] = ~((inputs[191]) | (inputs[36]));
    assign layer0_outputs[727] = (inputs[3]) | (inputs[212]);
    assign layer0_outputs[728] = ~(inputs[64]);
    assign layer0_outputs[729] = (inputs[230]) | (inputs[4]);
    assign layer0_outputs[730] = ~((inputs[4]) ^ (inputs[102]));
    assign layer0_outputs[731] = ~((inputs[229]) | (inputs[175]));
    assign layer0_outputs[732] = ~((inputs[253]) & (inputs[236]));
    assign layer0_outputs[733] = (inputs[49]) | (inputs[124]);
    assign layer0_outputs[734] = (inputs[63]) | (inputs[8]);
    assign layer0_outputs[735] = inputs[164];
    assign layer0_outputs[736] = ~((inputs[66]) | (inputs[67]));
    assign layer0_outputs[737] = (inputs[207]) & ~(inputs[241]);
    assign layer0_outputs[738] = ~((inputs[197]) ^ (inputs[14]));
    assign layer0_outputs[739] = ~(inputs[252]) | (inputs[197]);
    assign layer0_outputs[740] = ~((inputs[165]) & (inputs[151]));
    assign layer0_outputs[741] = ~((inputs[85]) | (inputs[35]));
    assign layer0_outputs[742] = ~(inputs[226]) | (inputs[141]);
    assign layer0_outputs[743] = ~((inputs[183]) ^ (inputs[149]));
    assign layer0_outputs[744] = (inputs[222]) & ~(inputs[155]);
    assign layer0_outputs[745] = (inputs[57]) | (inputs[120]);
    assign layer0_outputs[746] = ~((inputs[240]) & (inputs[147]));
    assign layer0_outputs[747] = ~((inputs[106]) & (inputs[10]));
    assign layer0_outputs[748] = ~(inputs[85]);
    assign layer0_outputs[749] = ~(inputs[104]);
    assign layer0_outputs[750] = (inputs[183]) & ~(inputs[144]);
    assign layer0_outputs[751] = inputs[166];
    assign layer0_outputs[752] = ~((inputs[200]) & (inputs[228]));
    assign layer0_outputs[753] = (inputs[178]) | (inputs[146]);
    assign layer0_outputs[754] = (inputs[192]) & ~(inputs[241]);
    assign layer0_outputs[755] = ~((inputs[188]) | (inputs[34]));
    assign layer0_outputs[756] = (inputs[221]) & (inputs[202]);
    assign layer0_outputs[757] = (inputs[146]) ^ (inputs[215]);
    assign layer0_outputs[758] = ~((inputs[8]) ^ (inputs[217]));
    assign layer0_outputs[759] = 1'b1;
    assign layer0_outputs[760] = inputs[226];
    assign layer0_outputs[761] = (inputs[71]) ^ (inputs[83]);
    assign layer0_outputs[762] = (inputs[159]) | (inputs[126]);
    assign layer0_outputs[763] = (inputs[127]) | (inputs[148]);
    assign layer0_outputs[764] = ~((inputs[57]) | (inputs[49]));
    assign layer0_outputs[765] = inputs[198];
    assign layer0_outputs[766] = ~(inputs[67]) | (inputs[221]);
    assign layer0_outputs[767] = ~((inputs[92]) | (inputs[49]));
    assign layer0_outputs[768] = inputs[78];
    assign layer0_outputs[769] = ~((inputs[39]) & (inputs[115]));
    assign layer0_outputs[770] = (inputs[243]) ^ (inputs[13]);
    assign layer0_outputs[771] = ~(inputs[120]);
    assign layer0_outputs[772] = (inputs[146]) | (inputs[162]);
    assign layer0_outputs[773] = (inputs[246]) & ~(inputs[161]);
    assign layer0_outputs[774] = (inputs[68]) & ~(inputs[247]);
    assign layer0_outputs[775] = (inputs[213]) & ~(inputs[164]);
    assign layer0_outputs[776] = ~((inputs[199]) | (inputs[104]));
    assign layer0_outputs[777] = (inputs[222]) | (inputs[36]);
    assign layer0_outputs[778] = ~(inputs[81]);
    assign layer0_outputs[779] = inputs[173];
    assign layer0_outputs[780] = ~(inputs[98]);
    assign layer0_outputs[781] = (inputs[104]) ^ (inputs[42]);
    assign layer0_outputs[782] = ~(inputs[150]);
    assign layer0_outputs[783] = ~((inputs[170]) ^ (inputs[233]));
    assign layer0_outputs[784] = ~(inputs[39]) | (inputs[124]);
    assign layer0_outputs[785] = ~(inputs[177]);
    assign layer0_outputs[786] = inputs[225];
    assign layer0_outputs[787] = (inputs[66]) | (inputs[43]);
    assign layer0_outputs[788] = (inputs[125]) | (inputs[3]);
    assign layer0_outputs[789] = ~((inputs[162]) | (inputs[251]));
    assign layer0_outputs[790] = inputs[26];
    assign layer0_outputs[791] = (inputs[193]) | (inputs[68]);
    assign layer0_outputs[792] = 1'b0;
    assign layer0_outputs[793] = ~((inputs[134]) ^ (inputs[167]));
    assign layer0_outputs[794] = (inputs[117]) ^ (inputs[129]);
    assign layer0_outputs[795] = ~(inputs[99]);
    assign layer0_outputs[796] = ~((inputs[53]) | (inputs[47]));
    assign layer0_outputs[797] = (inputs[98]) & ~(inputs[250]);
    assign layer0_outputs[798] = ~(inputs[83]);
    assign layer0_outputs[799] = inputs[203];
    assign layer0_outputs[800] = ~(inputs[173]) | (inputs[128]);
    assign layer0_outputs[801] = ~(inputs[202]);
    assign layer0_outputs[802] = (inputs[135]) | (inputs[245]);
    assign layer0_outputs[803] = ~(inputs[200]) | (inputs[228]);
    assign layer0_outputs[804] = ~(inputs[21]);
    assign layer0_outputs[805] = ~(inputs[11]);
    assign layer0_outputs[806] = (inputs[242]) ^ (inputs[74]);
    assign layer0_outputs[807] = inputs[184];
    assign layer0_outputs[808] = (inputs[140]) ^ (inputs[170]);
    assign layer0_outputs[809] = (inputs[88]) ^ (inputs[93]);
    assign layer0_outputs[810] = inputs[195];
    assign layer0_outputs[811] = inputs[179];
    assign layer0_outputs[812] = (inputs[191]) & (inputs[151]);
    assign layer0_outputs[813] = ~(inputs[108]);
    assign layer0_outputs[814] = ~((inputs[148]) & (inputs[159]));
    assign layer0_outputs[815] = inputs[157];
    assign layer0_outputs[816] = (inputs[140]) ^ (inputs[27]);
    assign layer0_outputs[817] = (inputs[154]) & ~(inputs[167]);
    assign layer0_outputs[818] = inputs[200];
    assign layer0_outputs[819] = (inputs[136]) & ~(inputs[4]);
    assign layer0_outputs[820] = inputs[128];
    assign layer0_outputs[821] = ~(inputs[212]) | (inputs[83]);
    assign layer0_outputs[822] = ~(inputs[71]);
    assign layer0_outputs[823] = ~(inputs[56]);
    assign layer0_outputs[824] = inputs[61];
    assign layer0_outputs[825] = (inputs[5]) | (inputs[241]);
    assign layer0_outputs[826] = (inputs[50]) | (inputs[76]);
    assign layer0_outputs[827] = ~((inputs[75]) | (inputs[10]));
    assign layer0_outputs[828] = ~(inputs[136]);
    assign layer0_outputs[829] = (inputs[49]) & ~(inputs[46]);
    assign layer0_outputs[830] = inputs[88];
    assign layer0_outputs[831] = ~((inputs[241]) ^ (inputs[1]));
    assign layer0_outputs[832] = (inputs[108]) & ~(inputs[83]);
    assign layer0_outputs[833] = (inputs[61]) | (inputs[98]);
    assign layer0_outputs[834] = ~((inputs[220]) | (inputs[174]));
    assign layer0_outputs[835] = ~(inputs[33]) | (inputs[127]);
    assign layer0_outputs[836] = ~((inputs[206]) ^ (inputs[110]));
    assign layer0_outputs[837] = (inputs[233]) | (inputs[202]);
    assign layer0_outputs[838] = (inputs[14]) | (inputs[100]);
    assign layer0_outputs[839] = ~((inputs[6]) | (inputs[33]));
    assign layer0_outputs[840] = inputs[169];
    assign layer0_outputs[841] = 1'b1;
    assign layer0_outputs[842] = inputs[148];
    assign layer0_outputs[843] = ~(inputs[8]);
    assign layer0_outputs[844] = ~((inputs[110]) | (inputs[75]));
    assign layer0_outputs[845] = (inputs[74]) & ~(inputs[35]);
    assign layer0_outputs[846] = inputs[133];
    assign layer0_outputs[847] = (inputs[126]) | (inputs[12]);
    assign layer0_outputs[848] = (inputs[79]) ^ (inputs[21]);
    assign layer0_outputs[849] = inputs[134];
    assign layer0_outputs[850] = (inputs[73]) & ~(inputs[193]);
    assign layer0_outputs[851] = ~(inputs[233]) | (inputs[253]);
    assign layer0_outputs[852] = ~(inputs[20]);
    assign layer0_outputs[853] = ~(inputs[113]) | (inputs[55]);
    assign layer0_outputs[854] = ~((inputs[46]) ^ (inputs[133]));
    assign layer0_outputs[855] = ~((inputs[238]) | (inputs[40]));
    assign layer0_outputs[856] = ~(inputs[142]) | (inputs[121]);
    assign layer0_outputs[857] = ~(inputs[244]) | (inputs[103]);
    assign layer0_outputs[858] = ~(inputs[99]) | (inputs[15]);
    assign layer0_outputs[859] = ~(inputs[108]) | (inputs[207]);
    assign layer0_outputs[860] = ~((inputs[251]) | (inputs[159]));
    assign layer0_outputs[861] = inputs[68];
    assign layer0_outputs[862] = inputs[195];
    assign layer0_outputs[863] = (inputs[208]) | (inputs[217]);
    assign layer0_outputs[864] = ~(inputs[190]);
    assign layer0_outputs[865] = (inputs[252]) | (inputs[230]);
    assign layer0_outputs[866] = ~(inputs[203]) | (inputs[118]);
    assign layer0_outputs[867] = ~((inputs[41]) & (inputs[44]));
    assign layer0_outputs[868] = inputs[201];
    assign layer0_outputs[869] = (inputs[9]) & ~(inputs[65]);
    assign layer0_outputs[870] = ~((inputs[251]) | (inputs[133]));
    assign layer0_outputs[871] = (inputs[153]) | (inputs[17]);
    assign layer0_outputs[872] = ~(inputs[117]) | (inputs[62]);
    assign layer0_outputs[873] = inputs[89];
    assign layer0_outputs[874] = ~((inputs[38]) | (inputs[193]));
    assign layer0_outputs[875] = ~(inputs[123]);
    assign layer0_outputs[876] = ~(inputs[244]);
    assign layer0_outputs[877] = (inputs[81]) | (inputs[103]);
    assign layer0_outputs[878] = ~((inputs[67]) ^ (inputs[84]));
    assign layer0_outputs[879] = ~(inputs[143]);
    assign layer0_outputs[880] = ~((inputs[245]) ^ (inputs[214]));
    assign layer0_outputs[881] = inputs[236];
    assign layer0_outputs[882] = (inputs[218]) ^ (inputs[209]);
    assign layer0_outputs[883] = ~(inputs[122]);
    assign layer0_outputs[884] = ~(inputs[98]);
    assign layer0_outputs[885] = inputs[196];
    assign layer0_outputs[886] = 1'b1;
    assign layer0_outputs[887] = (inputs[104]) & ~(inputs[152]);
    assign layer0_outputs[888] = inputs[162];
    assign layer0_outputs[889] = (inputs[87]) & ~(inputs[16]);
    assign layer0_outputs[890] = ~((inputs[15]) ^ (inputs[150]));
    assign layer0_outputs[891] = ~(inputs[43]);
    assign layer0_outputs[892] = ~((inputs[44]) & (inputs[12]));
    assign layer0_outputs[893] = ~(inputs[242]);
    assign layer0_outputs[894] = (inputs[28]) & (inputs[9]);
    assign layer0_outputs[895] = inputs[159];
    assign layer0_outputs[896] = ~(inputs[118]) | (inputs[160]);
    assign layer0_outputs[897] = ~((inputs[134]) ^ (inputs[163]));
    assign layer0_outputs[898] = ~((inputs[203]) & (inputs[224]));
    assign layer0_outputs[899] = ~((inputs[143]) ^ (inputs[233]));
    assign layer0_outputs[900] = inputs[67];
    assign layer0_outputs[901] = ~(inputs[116]);
    assign layer0_outputs[902] = inputs[56];
    assign layer0_outputs[903] = (inputs[180]) | (inputs[209]);
    assign layer0_outputs[904] = ~(inputs[203]);
    assign layer0_outputs[905] = (inputs[23]) ^ (inputs[211]);
    assign layer0_outputs[906] = inputs[112];
    assign layer0_outputs[907] = (inputs[149]) & ~(inputs[20]);
    assign layer0_outputs[908] = (inputs[45]) | (inputs[244]);
    assign layer0_outputs[909] = (inputs[163]) & (inputs[227]);
    assign layer0_outputs[910] = inputs[14];
    assign layer0_outputs[911] = (inputs[223]) | (inputs[212]);
    assign layer0_outputs[912] = ~((inputs[116]) ^ (inputs[122]));
    assign layer0_outputs[913] = ~((inputs[183]) | (inputs[62]));
    assign layer0_outputs[914] = ~(inputs[132]);
    assign layer0_outputs[915] = ~(inputs[20]) | (inputs[69]);
    assign layer0_outputs[916] = inputs[228];
    assign layer0_outputs[917] = (inputs[60]) & ~(inputs[214]);
    assign layer0_outputs[918] = (inputs[150]) & ~(inputs[113]);
    assign layer0_outputs[919] = ~(inputs[133]);
    assign layer0_outputs[920] = ~((inputs[201]) | (inputs[190]));
    assign layer0_outputs[921] = ~(inputs[51]) | (inputs[110]);
    assign layer0_outputs[922] = ~(inputs[218]);
    assign layer0_outputs[923] = (inputs[5]) | (inputs[206]);
    assign layer0_outputs[924] = 1'b0;
    assign layer0_outputs[925] = (inputs[89]) & ~(inputs[31]);
    assign layer0_outputs[926] = ~(inputs[131]);
    assign layer0_outputs[927] = ~(inputs[184]);
    assign layer0_outputs[928] = ~((inputs[5]) ^ (inputs[169]));
    assign layer0_outputs[929] = inputs[197];
    assign layer0_outputs[930] = ~((inputs[109]) ^ (inputs[156]));
    assign layer0_outputs[931] = (inputs[163]) ^ (inputs[125]);
    assign layer0_outputs[932] = (inputs[27]) ^ (inputs[145]);
    assign layer0_outputs[933] = ~(inputs[166]) | (inputs[225]);
    assign layer0_outputs[934] = (inputs[7]) | (inputs[22]);
    assign layer0_outputs[935] = (inputs[120]) & (inputs[113]);
    assign layer0_outputs[936] = ~((inputs[115]) | (inputs[162]));
    assign layer0_outputs[937] = ~((inputs[76]) & (inputs[107]));
    assign layer0_outputs[938] = 1'b0;
    assign layer0_outputs[939] = ~(inputs[147]);
    assign layer0_outputs[940] = inputs[145];
    assign layer0_outputs[941] = ~((inputs[86]) | (inputs[100]));
    assign layer0_outputs[942] = 1'b1;
    assign layer0_outputs[943] = ~((inputs[142]) | (inputs[207]));
    assign layer0_outputs[944] = ~((inputs[221]) | (inputs[17]));
    assign layer0_outputs[945] = ~((inputs[64]) | (inputs[66]));
    assign layer0_outputs[946] = (inputs[92]) & ~(inputs[67]);
    assign layer0_outputs[947] = (inputs[92]) ^ (inputs[1]);
    assign layer0_outputs[948] = ~(inputs[19]);
    assign layer0_outputs[949] = (inputs[16]) | (inputs[85]);
    assign layer0_outputs[950] = inputs[133];
    assign layer0_outputs[951] = ~(inputs[81]) | (inputs[156]);
    assign layer0_outputs[952] = (inputs[151]) ^ (inputs[194]);
    assign layer0_outputs[953] = (inputs[150]) ^ (inputs[103]);
    assign layer0_outputs[954] = ~((inputs[224]) | (inputs[77]));
    assign layer0_outputs[955] = ~(inputs[232]);
    assign layer0_outputs[956] = ~(inputs[223]) | (inputs[226]);
    assign layer0_outputs[957] = inputs[111];
    assign layer0_outputs[958] = inputs[52];
    assign layer0_outputs[959] = ~((inputs[143]) | (inputs[67]));
    assign layer0_outputs[960] = (inputs[93]) & ~(inputs[240]);
    assign layer0_outputs[961] = (inputs[235]) & ~(inputs[132]);
    assign layer0_outputs[962] = (inputs[131]) & ~(inputs[203]);
    assign layer0_outputs[963] = ~((inputs[42]) | (inputs[124]));
    assign layer0_outputs[964] = ~((inputs[150]) | (inputs[176]));
    assign layer0_outputs[965] = (inputs[210]) | (inputs[240]);
    assign layer0_outputs[966] = inputs[230];
    assign layer0_outputs[967] = (inputs[25]) | (inputs[65]);
    assign layer0_outputs[968] = (inputs[119]) & ~(inputs[170]);
    assign layer0_outputs[969] = (inputs[228]) | (inputs[191]);
    assign layer0_outputs[970] = (inputs[249]) & ~(inputs[239]);
    assign layer0_outputs[971] = (inputs[135]) | (inputs[65]);
    assign layer0_outputs[972] = inputs[49];
    assign layer0_outputs[973] = ~(inputs[21]);
    assign layer0_outputs[974] = (inputs[43]) ^ (inputs[181]);
    assign layer0_outputs[975] = (inputs[77]) | (inputs[93]);
    assign layer0_outputs[976] = 1'b1;
    assign layer0_outputs[977] = (inputs[97]) & ~(inputs[224]);
    assign layer0_outputs[978] = inputs[162];
    assign layer0_outputs[979] = inputs[253];
    assign layer0_outputs[980] = (inputs[71]) ^ (inputs[83]);
    assign layer0_outputs[981] = inputs[39];
    assign layer0_outputs[982] = ~(inputs[169]);
    assign layer0_outputs[983] = inputs[144];
    assign layer0_outputs[984] = inputs[38];
    assign layer0_outputs[985] = ~(inputs[109]) | (inputs[9]);
    assign layer0_outputs[986] = inputs[130];
    assign layer0_outputs[987] = ~(inputs[214]);
    assign layer0_outputs[988] = 1'b0;
    assign layer0_outputs[989] = ~(inputs[251]);
    assign layer0_outputs[990] = inputs[163];
    assign layer0_outputs[991] = ~(inputs[248]);
    assign layer0_outputs[992] = (inputs[117]) ^ (inputs[234]);
    assign layer0_outputs[993] = (inputs[18]) ^ (inputs[9]);
    assign layer0_outputs[994] = 1'b0;
    assign layer0_outputs[995] = ~((inputs[0]) & (inputs[184]));
    assign layer0_outputs[996] = inputs[23];
    assign layer0_outputs[997] = ~(inputs[247]) | (inputs[7]);
    assign layer0_outputs[998] = ~(inputs[212]);
    assign layer0_outputs[999] = ~((inputs[196]) | (inputs[176]));
    assign layer0_outputs[1000] = ~(inputs[138]) | (inputs[236]);
    assign layer0_outputs[1001] = ~(inputs[107]);
    assign layer0_outputs[1002] = (inputs[217]) & ~(inputs[65]);
    assign layer0_outputs[1003] = inputs[68];
    assign layer0_outputs[1004] = (inputs[217]) & ~(inputs[237]);
    assign layer0_outputs[1005] = inputs[211];
    assign layer0_outputs[1006] = inputs[209];
    assign layer0_outputs[1007] = ~((inputs[250]) | (inputs[109]));
    assign layer0_outputs[1008] = ~((inputs[105]) | (inputs[106]));
    assign layer0_outputs[1009] = ~((inputs[33]) & (inputs[227]));
    assign layer0_outputs[1010] = (inputs[107]) ^ (inputs[197]);
    assign layer0_outputs[1011] = ~(inputs[83]);
    assign layer0_outputs[1012] = ~(inputs[38]);
    assign layer0_outputs[1013] = inputs[216];
    assign layer0_outputs[1014] = (inputs[52]) | (inputs[28]);
    assign layer0_outputs[1015] = (inputs[193]) & ~(inputs[50]);
    assign layer0_outputs[1016] = (inputs[156]) & (inputs[59]);
    assign layer0_outputs[1017] = ~(inputs[51]);
    assign layer0_outputs[1018] = (inputs[109]) & ~(inputs[207]);
    assign layer0_outputs[1019] = (inputs[99]) ^ (inputs[73]);
    assign layer0_outputs[1020] = ~(inputs[111]);
    assign layer0_outputs[1021] = ~((inputs[77]) | (inputs[35]));
    assign layer0_outputs[1022] = inputs[89];
    assign layer0_outputs[1023] = inputs[82];
    assign layer0_outputs[1024] = ~((inputs[238]) | (inputs[50]));
    assign layer0_outputs[1025] = 1'b0;
    assign layer0_outputs[1026] = inputs[101];
    assign layer0_outputs[1027] = ~((inputs[204]) | (inputs[240]));
    assign layer0_outputs[1028] = 1'b1;
    assign layer0_outputs[1029] = (inputs[152]) & ~(inputs[28]);
    assign layer0_outputs[1030] = (inputs[80]) ^ (inputs[167]);
    assign layer0_outputs[1031] = inputs[232];
    assign layer0_outputs[1032] = ~((inputs[195]) | (inputs[245]));
    assign layer0_outputs[1033] = ~(inputs[113]);
    assign layer0_outputs[1034] = ~(inputs[126]);
    assign layer0_outputs[1035] = ~((inputs[11]) | (inputs[31]));
    assign layer0_outputs[1036] = inputs[90];
    assign layer0_outputs[1037] = inputs[147];
    assign layer0_outputs[1038] = (inputs[240]) | (inputs[24]);
    assign layer0_outputs[1039] = (inputs[10]) & ~(inputs[88]);
    assign layer0_outputs[1040] = (inputs[60]) | (inputs[195]);
    assign layer0_outputs[1041] = (inputs[39]) | (inputs[35]);
    assign layer0_outputs[1042] = ~(inputs[167]);
    assign layer0_outputs[1043] = 1'b1;
    assign layer0_outputs[1044] = ~((inputs[174]) | (inputs[176]));
    assign layer0_outputs[1045] = ~(inputs[75]);
    assign layer0_outputs[1046] = ~(inputs[252]);
    assign layer0_outputs[1047] = (inputs[129]) | (inputs[59]);
    assign layer0_outputs[1048] = ~(inputs[227]);
    assign layer0_outputs[1049] = (inputs[61]) & (inputs[11]);
    assign layer0_outputs[1050] = inputs[163];
    assign layer0_outputs[1051] = ~((inputs[65]) | (inputs[47]));
    assign layer0_outputs[1052] = inputs[66];
    assign layer0_outputs[1053] = (inputs[89]) ^ (inputs[232]);
    assign layer0_outputs[1054] = (inputs[13]) & ~(inputs[191]);
    assign layer0_outputs[1055] = ~((inputs[225]) ^ (inputs[26]));
    assign layer0_outputs[1056] = ~(inputs[191]);
    assign layer0_outputs[1057] = ~((inputs[89]) ^ (inputs[134]));
    assign layer0_outputs[1058] = 1'b1;
    assign layer0_outputs[1059] = ~((inputs[127]) | (inputs[182]));
    assign layer0_outputs[1060] = ~((inputs[47]) | (inputs[23]));
    assign layer0_outputs[1061] = ~(inputs[95]);
    assign layer0_outputs[1062] = ~(inputs[214]);
    assign layer0_outputs[1063] = (inputs[162]) | (inputs[190]);
    assign layer0_outputs[1064] = inputs[2];
    assign layer0_outputs[1065] = (inputs[183]) ^ (inputs[109]);
    assign layer0_outputs[1066] = (inputs[252]) | (inputs[54]);
    assign layer0_outputs[1067] = inputs[251];
    assign layer0_outputs[1068] = ~(inputs[121]) | (inputs[129]);
    assign layer0_outputs[1069] = inputs[190];
    assign layer0_outputs[1070] = ~((inputs[118]) | (inputs[248]));
    assign layer0_outputs[1071] = (inputs[184]) & (inputs[241]);
    assign layer0_outputs[1072] = inputs[234];
    assign layer0_outputs[1073] = ~(inputs[37]) | (inputs[234]);
    assign layer0_outputs[1074] = (inputs[111]) | (inputs[1]);
    assign layer0_outputs[1075] = (inputs[254]) | (inputs[146]);
    assign layer0_outputs[1076] = (inputs[179]) | (inputs[49]);
    assign layer0_outputs[1077] = ~(inputs[231]);
    assign layer0_outputs[1078] = (inputs[86]) | (inputs[109]);
    assign layer0_outputs[1079] = (inputs[219]) | (inputs[2]);
    assign layer0_outputs[1080] = ~(inputs[44]);
    assign layer0_outputs[1081] = ~(inputs[120]);
    assign layer0_outputs[1082] = (inputs[179]) & ~(inputs[78]);
    assign layer0_outputs[1083] = ~((inputs[35]) | (inputs[247]));
    assign layer0_outputs[1084] = inputs[16];
    assign layer0_outputs[1085] = ~(inputs[206]) | (inputs[48]);
    assign layer0_outputs[1086] = ~(inputs[106]) | (inputs[235]);
    assign layer0_outputs[1087] = ~(inputs[107]);
    assign layer0_outputs[1088] = ~(inputs[50]) | (inputs[61]);
    assign layer0_outputs[1089] = (inputs[173]) & ~(inputs[247]);
    assign layer0_outputs[1090] = ~(inputs[74]);
    assign layer0_outputs[1091] = (inputs[27]) | (inputs[57]);
    assign layer0_outputs[1092] = ~((inputs[51]) & (inputs[7]));
    assign layer0_outputs[1093] = ~((inputs[173]) ^ (inputs[83]));
    assign layer0_outputs[1094] = ~(inputs[174]);
    assign layer0_outputs[1095] = (inputs[53]) | (inputs[9]);
    assign layer0_outputs[1096] = ~((inputs[152]) ^ (inputs[165]));
    assign layer0_outputs[1097] = ~(inputs[167]);
    assign layer0_outputs[1098] = ~(inputs[229]);
    assign layer0_outputs[1099] = ~(inputs[203]) | (inputs[32]);
    assign layer0_outputs[1100] = inputs[79];
    assign layer0_outputs[1101] = inputs[114];
    assign layer0_outputs[1102] = (inputs[85]) ^ (inputs[113]);
    assign layer0_outputs[1103] = (inputs[123]) ^ (inputs[57]);
    assign layer0_outputs[1104] = (inputs[56]) & ~(inputs[205]);
    assign layer0_outputs[1105] = (inputs[82]) & ~(inputs[152]);
    assign layer0_outputs[1106] = (inputs[190]) ^ (inputs[125]);
    assign layer0_outputs[1107] = (inputs[146]) ^ (inputs[194]);
    assign layer0_outputs[1108] = ~((inputs[79]) | (inputs[164]));
    assign layer0_outputs[1109] = (inputs[84]) & ~(inputs[160]);
    assign layer0_outputs[1110] = (inputs[184]) & ~(inputs[205]);
    assign layer0_outputs[1111] = 1'b1;
    assign layer0_outputs[1112] = 1'b1;
    assign layer0_outputs[1113] = inputs[129];
    assign layer0_outputs[1114] = ~((inputs[255]) | (inputs[185]));
    assign layer0_outputs[1115] = inputs[92];
    assign layer0_outputs[1116] = ~(inputs[139]) | (inputs[248]);
    assign layer0_outputs[1117] = ~(inputs[120]);
    assign layer0_outputs[1118] = (inputs[77]) & ~(inputs[99]);
    assign layer0_outputs[1119] = inputs[107];
    assign layer0_outputs[1120] = inputs[212];
    assign layer0_outputs[1121] = ~((inputs[139]) ^ (inputs[254]));
    assign layer0_outputs[1122] = ~(inputs[139]);
    assign layer0_outputs[1123] = ~((inputs[116]) ^ (inputs[144]));
    assign layer0_outputs[1124] = ~(inputs[119]) | (inputs[141]);
    assign layer0_outputs[1125] = ~(inputs[232]) | (inputs[1]);
    assign layer0_outputs[1126] = ~((inputs[201]) ^ (inputs[249]));
    assign layer0_outputs[1127] = inputs[224];
    assign layer0_outputs[1128] = ~(inputs[135]) | (inputs[143]);
    assign layer0_outputs[1129] = (inputs[82]) ^ (inputs[36]);
    assign layer0_outputs[1130] = (inputs[168]) ^ (inputs[119]);
    assign layer0_outputs[1131] = inputs[191];
    assign layer0_outputs[1132] = (inputs[63]) | (inputs[119]);
    assign layer0_outputs[1133] = ~((inputs[162]) | (inputs[126]));
    assign layer0_outputs[1134] = (inputs[166]) ^ (inputs[0]);
    assign layer0_outputs[1135] = (inputs[245]) ^ (inputs[38]);
    assign layer0_outputs[1136] = (inputs[157]) ^ (inputs[21]);
    assign layer0_outputs[1137] = ~(inputs[217]);
    assign layer0_outputs[1138] = (inputs[42]) & ~(inputs[120]);
    assign layer0_outputs[1139] = inputs[63];
    assign layer0_outputs[1140] = (inputs[251]) & ~(inputs[160]);
    assign layer0_outputs[1141] = ~((inputs[4]) | (inputs[195]));
    assign layer0_outputs[1142] = inputs[19];
    assign layer0_outputs[1143] = inputs[238];
    assign layer0_outputs[1144] = (inputs[249]) | (inputs[172]);
    assign layer0_outputs[1145] = ~(inputs[194]);
    assign layer0_outputs[1146] = ~((inputs[232]) ^ (inputs[22]));
    assign layer0_outputs[1147] = ~((inputs[230]) | (inputs[206]));
    assign layer0_outputs[1148] = ~(inputs[220]) | (inputs[240]);
    assign layer0_outputs[1149] = ~(inputs[75]) | (inputs[102]);
    assign layer0_outputs[1150] = inputs[126];
    assign layer0_outputs[1151] = ~((inputs[210]) | (inputs[25]));
    assign layer0_outputs[1152] = (inputs[116]) ^ (inputs[169]);
    assign layer0_outputs[1153] = inputs[209];
    assign layer0_outputs[1154] = ~((inputs[144]) | (inputs[32]));
    assign layer0_outputs[1155] = inputs[79];
    assign layer0_outputs[1156] = ~(inputs[158]) | (inputs[87]);
    assign layer0_outputs[1157] = ~((inputs[192]) | (inputs[77]));
    assign layer0_outputs[1158] = ~(inputs[30]) | (inputs[242]);
    assign layer0_outputs[1159] = (inputs[136]) & ~(inputs[143]);
    assign layer0_outputs[1160] = ~((inputs[14]) ^ (inputs[13]));
    assign layer0_outputs[1161] = (inputs[186]) & ~(inputs[69]);
    assign layer0_outputs[1162] = inputs[194];
    assign layer0_outputs[1163] = (inputs[28]) ^ (inputs[37]);
    assign layer0_outputs[1164] = ~((inputs[238]) | (inputs[5]));
    assign layer0_outputs[1165] = ~((inputs[154]) | (inputs[88]));
    assign layer0_outputs[1166] = ~(inputs[149]);
    assign layer0_outputs[1167] = (inputs[167]) & ~(inputs[31]);
    assign layer0_outputs[1168] = ~((inputs[161]) ^ (inputs[249]));
    assign layer0_outputs[1169] = ~(inputs[4]);
    assign layer0_outputs[1170] = ~((inputs[209]) | (inputs[114]));
    assign layer0_outputs[1171] = (inputs[146]) & ~(inputs[149]);
    assign layer0_outputs[1172] = (inputs[247]) ^ (inputs[220]);
    assign layer0_outputs[1173] = ~((inputs[230]) ^ (inputs[162]));
    assign layer0_outputs[1174] = ~((inputs[228]) & (inputs[210]));
    assign layer0_outputs[1175] = ~(inputs[83]) | (inputs[248]);
    assign layer0_outputs[1176] = ~(inputs[160]);
    assign layer0_outputs[1177] = ~((inputs[112]) ^ (inputs[86]));
    assign layer0_outputs[1178] = (inputs[53]) | (inputs[6]);
    assign layer0_outputs[1179] = (inputs[164]) & ~(inputs[45]);
    assign layer0_outputs[1180] = 1'b1;
    assign layer0_outputs[1181] = ~((inputs[67]) | (inputs[215]));
    assign layer0_outputs[1182] = ~((inputs[19]) | (inputs[75]));
    assign layer0_outputs[1183] = ~(inputs[227]);
    assign layer0_outputs[1184] = ~(inputs[217]) | (inputs[1]);
    assign layer0_outputs[1185] = ~((inputs[197]) ^ (inputs[162]));
    assign layer0_outputs[1186] = ~(inputs[97]);
    assign layer0_outputs[1187] = (inputs[242]) & ~(inputs[129]);
    assign layer0_outputs[1188] = ~(inputs[101]);
    assign layer0_outputs[1189] = (inputs[127]) & ~(inputs[169]);
    assign layer0_outputs[1190] = ~(inputs[212]);
    assign layer0_outputs[1191] = (inputs[24]) & ~(inputs[192]);
    assign layer0_outputs[1192] = ~(inputs[56]) | (inputs[201]);
    assign layer0_outputs[1193] = ~((inputs[12]) ^ (inputs[36]));
    assign layer0_outputs[1194] = inputs[222];
    assign layer0_outputs[1195] = inputs[41];
    assign layer0_outputs[1196] = inputs[63];
    assign layer0_outputs[1197] = (inputs[246]) & ~(inputs[0]);
    assign layer0_outputs[1198] = inputs[115];
    assign layer0_outputs[1199] = ~((inputs[198]) ^ (inputs[244]));
    assign layer0_outputs[1200] = ~((inputs[225]) | (inputs[5]));
    assign layer0_outputs[1201] = ~(inputs[108]) | (inputs[240]);
    assign layer0_outputs[1202] = (inputs[17]) ^ (inputs[11]);
    assign layer0_outputs[1203] = inputs[74];
    assign layer0_outputs[1204] = ~((inputs[194]) | (inputs[241]));
    assign layer0_outputs[1205] = (inputs[177]) ^ (inputs[118]);
    assign layer0_outputs[1206] = ~((inputs[220]) ^ (inputs[21]));
    assign layer0_outputs[1207] = ~((inputs[205]) | (inputs[224]));
    assign layer0_outputs[1208] = ~(inputs[86]) | (inputs[127]);
    assign layer0_outputs[1209] = (inputs[247]) & (inputs[222]);
    assign layer0_outputs[1210] = ~((inputs[79]) | (inputs[242]));
    assign layer0_outputs[1211] = (inputs[178]) | (inputs[146]);
    assign layer0_outputs[1212] = (inputs[23]) & ~(inputs[227]);
    assign layer0_outputs[1213] = ~((inputs[77]) | (inputs[226]));
    assign layer0_outputs[1214] = inputs[35];
    assign layer0_outputs[1215] = (inputs[26]) & ~(inputs[89]);
    assign layer0_outputs[1216] = ~((inputs[55]) ^ (inputs[244]));
    assign layer0_outputs[1217] = ~(inputs[57]) | (inputs[151]);
    assign layer0_outputs[1218] = ~((inputs[117]) ^ (inputs[26]));
    assign layer0_outputs[1219] = 1'b1;
    assign layer0_outputs[1220] = inputs[194];
    assign layer0_outputs[1221] = 1'b0;
    assign layer0_outputs[1222] = (inputs[231]) & ~(inputs[13]);
    assign layer0_outputs[1223] = ~(inputs[113]);
    assign layer0_outputs[1224] = (inputs[22]) ^ (inputs[156]);
    assign layer0_outputs[1225] = inputs[88];
    assign layer0_outputs[1226] = ~(inputs[220]);
    assign layer0_outputs[1227] = ~(inputs[117]);
    assign layer0_outputs[1228] = inputs[246];
    assign layer0_outputs[1229] = (inputs[251]) ^ (inputs[196]);
    assign layer0_outputs[1230] = (inputs[110]) ^ (inputs[37]);
    assign layer0_outputs[1231] = ~(inputs[90]) | (inputs[164]);
    assign layer0_outputs[1232] = ~(inputs[8]);
    assign layer0_outputs[1233] = (inputs[59]) | (inputs[238]);
    assign layer0_outputs[1234] = (inputs[10]) & ~(inputs[220]);
    assign layer0_outputs[1235] = (inputs[193]) ^ (inputs[96]);
    assign layer0_outputs[1236] = (inputs[118]) & ~(inputs[33]);
    assign layer0_outputs[1237] = (inputs[39]) & ~(inputs[192]);
    assign layer0_outputs[1238] = ~(inputs[121]) | (inputs[55]);
    assign layer0_outputs[1239] = (inputs[132]) ^ (inputs[71]);
    assign layer0_outputs[1240] = inputs[147];
    assign layer0_outputs[1241] = (inputs[221]) ^ (inputs[202]);
    assign layer0_outputs[1242] = ~((inputs[60]) ^ (inputs[189]));
    assign layer0_outputs[1243] = ~((inputs[203]) & (inputs[162]));
    assign layer0_outputs[1244] = ~((inputs[95]) | (inputs[191]));
    assign layer0_outputs[1245] = ~((inputs[53]) | (inputs[216]));
    assign layer0_outputs[1246] = ~(inputs[204]);
    assign layer0_outputs[1247] = inputs[213];
    assign layer0_outputs[1248] = ~(inputs[165]);
    assign layer0_outputs[1249] = ~((inputs[186]) ^ (inputs[106]));
    assign layer0_outputs[1250] = inputs[107];
    assign layer0_outputs[1251] = inputs[67];
    assign layer0_outputs[1252] = ~(inputs[183]) | (inputs[158]);
    assign layer0_outputs[1253] = (inputs[254]) | (inputs[177]);
    assign layer0_outputs[1254] = (inputs[175]) ^ (inputs[119]);
    assign layer0_outputs[1255] = ~(inputs[101]);
    assign layer0_outputs[1256] = ~(inputs[180]) | (inputs[63]);
    assign layer0_outputs[1257] = ~(inputs[113]);
    assign layer0_outputs[1258] = (inputs[49]) | (inputs[6]);
    assign layer0_outputs[1259] = (inputs[170]) | (inputs[146]);
    assign layer0_outputs[1260] = ~(inputs[138]);
    assign layer0_outputs[1261] = ~(inputs[180]);
    assign layer0_outputs[1262] = (inputs[152]) ^ (inputs[255]);
    assign layer0_outputs[1263] = ~((inputs[235]) | (inputs[227]));
    assign layer0_outputs[1264] = inputs[147];
    assign layer0_outputs[1265] = inputs[72];
    assign layer0_outputs[1266] = ~(inputs[198]);
    assign layer0_outputs[1267] = inputs[115];
    assign layer0_outputs[1268] = ~(inputs[39]);
    assign layer0_outputs[1269] = ~(inputs[46]);
    assign layer0_outputs[1270] = ~(inputs[155]);
    assign layer0_outputs[1271] = ~((inputs[53]) & (inputs[43]));
    assign layer0_outputs[1272] = ~((inputs[24]) | (inputs[157]));
    assign layer0_outputs[1273] = inputs[10];
    assign layer0_outputs[1274] = ~(inputs[229]) | (inputs[151]);
    assign layer0_outputs[1275] = ~((inputs[92]) ^ (inputs[159]));
    assign layer0_outputs[1276] = ~(inputs[24]);
    assign layer0_outputs[1277] = (inputs[213]) ^ (inputs[128]);
    assign layer0_outputs[1278] = ~(inputs[151]);
    assign layer0_outputs[1279] = (inputs[76]) & ~(inputs[62]);
    assign layer0_outputs[1280] = ~((inputs[66]) & (inputs[4]));
    assign layer0_outputs[1281] = ~(inputs[25]);
    assign layer0_outputs[1282] = (inputs[0]) | (inputs[243]);
    assign layer0_outputs[1283] = ~(inputs[115]);
    assign layer0_outputs[1284] = (inputs[144]) | (inputs[186]);
    assign layer0_outputs[1285] = inputs[2];
    assign layer0_outputs[1286] = ~(inputs[81]) | (inputs[177]);
    assign layer0_outputs[1287] = (inputs[159]) | (inputs[172]);
    assign layer0_outputs[1288] = inputs[40];
    assign layer0_outputs[1289] = (inputs[86]) ^ (inputs[105]);
    assign layer0_outputs[1290] = inputs[52];
    assign layer0_outputs[1291] = (inputs[165]) | (inputs[180]);
    assign layer0_outputs[1292] = (inputs[51]) | (inputs[254]);
    assign layer0_outputs[1293] = ~((inputs[47]) ^ (inputs[15]));
    assign layer0_outputs[1294] = ~((inputs[6]) ^ (inputs[157]));
    assign layer0_outputs[1295] = ~(inputs[122]);
    assign layer0_outputs[1296] = (inputs[62]) ^ (inputs[189]);
    assign layer0_outputs[1297] = ~((inputs[241]) ^ (inputs[80]));
    assign layer0_outputs[1298] = (inputs[210]) & ~(inputs[8]);
    assign layer0_outputs[1299] = ~((inputs[57]) | (inputs[224]));
    assign layer0_outputs[1300] = ~((inputs[242]) | (inputs[199]));
    assign layer0_outputs[1301] = ~(inputs[150]) | (inputs[138]);
    assign layer0_outputs[1302] = ~(inputs[214]);
    assign layer0_outputs[1303] = (inputs[33]) & ~(inputs[82]);
    assign layer0_outputs[1304] = (inputs[62]) | (inputs[185]);
    assign layer0_outputs[1305] = inputs[206];
    assign layer0_outputs[1306] = (inputs[43]) ^ (inputs[87]);
    assign layer0_outputs[1307] = (inputs[73]) & ~(inputs[181]);
    assign layer0_outputs[1308] = ~(inputs[136]);
    assign layer0_outputs[1309] = ~((inputs[230]) & (inputs[232]));
    assign layer0_outputs[1310] = ~(inputs[144]) | (inputs[63]);
    assign layer0_outputs[1311] = ~(inputs[225]);
    assign layer0_outputs[1312] = ~(inputs[235]);
    assign layer0_outputs[1313] = inputs[66];
    assign layer0_outputs[1314] = (inputs[176]) & ~(inputs[142]);
    assign layer0_outputs[1315] = ~((inputs[30]) | (inputs[190]));
    assign layer0_outputs[1316] = ~(inputs[195]) | (inputs[81]);
    assign layer0_outputs[1317] = (inputs[44]) | (inputs[92]);
    assign layer0_outputs[1318] = ~((inputs[70]) | (inputs[130]));
    assign layer0_outputs[1319] = ~((inputs[234]) & (inputs[231]));
    assign layer0_outputs[1320] = ~(inputs[11]);
    assign layer0_outputs[1321] = ~((inputs[212]) ^ (inputs[82]));
    assign layer0_outputs[1322] = inputs[111];
    assign layer0_outputs[1323] = ~(inputs[52]) | (inputs[159]);
    assign layer0_outputs[1324] = ~((inputs[66]) ^ (inputs[36]));
    assign layer0_outputs[1325] = ~(inputs[47]) | (inputs[170]);
    assign layer0_outputs[1326] = ~((inputs[249]) & (inputs[248]));
    assign layer0_outputs[1327] = inputs[248];
    assign layer0_outputs[1328] = ~(inputs[98]);
    assign layer0_outputs[1329] = (inputs[101]) & ~(inputs[96]);
    assign layer0_outputs[1330] = ~((inputs[72]) ^ (inputs[60]));
    assign layer0_outputs[1331] = ~((inputs[32]) ^ (inputs[70]));
    assign layer0_outputs[1332] = ~((inputs[3]) | (inputs[41]));
    assign layer0_outputs[1333] = ~(inputs[241]) | (inputs[183]);
    assign layer0_outputs[1334] = ~(inputs[152]);
    assign layer0_outputs[1335] = inputs[107];
    assign layer0_outputs[1336] = (inputs[13]) | (inputs[111]);
    assign layer0_outputs[1337] = (inputs[122]) & ~(inputs[28]);
    assign layer0_outputs[1338] = inputs[238];
    assign layer0_outputs[1339] = inputs[209];
    assign layer0_outputs[1340] = ~((inputs[163]) ^ (inputs[80]));
    assign layer0_outputs[1341] = (inputs[94]) | (inputs[210]);
    assign layer0_outputs[1342] = inputs[47];
    assign layer0_outputs[1343] = (inputs[201]) | (inputs[129]);
    assign layer0_outputs[1344] = ~((inputs[219]) | (inputs[198]));
    assign layer0_outputs[1345] = inputs[214];
    assign layer0_outputs[1346] = (inputs[227]) & ~(inputs[122]);
    assign layer0_outputs[1347] = (inputs[8]) & ~(inputs[5]);
    assign layer0_outputs[1348] = ~(inputs[24]) | (inputs[158]);
    assign layer0_outputs[1349] = ~((inputs[123]) | (inputs[186]));
    assign layer0_outputs[1350] = (inputs[107]) ^ (inputs[49]);
    assign layer0_outputs[1351] = ~(inputs[242]) | (inputs[150]);
    assign layer0_outputs[1352] = inputs[199];
    assign layer0_outputs[1353] = (inputs[21]) ^ (inputs[95]);
    assign layer0_outputs[1354] = (inputs[220]) & ~(inputs[49]);
    assign layer0_outputs[1355] = ~(inputs[98]) | (inputs[225]);
    assign layer0_outputs[1356] = ~((inputs[69]) | (inputs[78]));
    assign layer0_outputs[1357] = ~((inputs[236]) | (inputs[47]));
    assign layer0_outputs[1358] = (inputs[229]) & ~(inputs[108]);
    assign layer0_outputs[1359] = (inputs[49]) | (inputs[104]);
    assign layer0_outputs[1360] = ~(inputs[88]);
    assign layer0_outputs[1361] = ~(inputs[115]) | (inputs[57]);
    assign layer0_outputs[1362] = ~(inputs[136]);
    assign layer0_outputs[1363] = ~(inputs[150]);
    assign layer0_outputs[1364] = (inputs[149]) | (inputs[181]);
    assign layer0_outputs[1365] = ~(inputs[77]);
    assign layer0_outputs[1366] = (inputs[140]) ^ (inputs[189]);
    assign layer0_outputs[1367] = (inputs[190]) & ~(inputs[58]);
    assign layer0_outputs[1368] = ~(inputs[66]) | (inputs[128]);
    assign layer0_outputs[1369] = ~(inputs[194]) | (inputs[244]);
    assign layer0_outputs[1370] = ~((inputs[198]) | (inputs[168]));
    assign layer0_outputs[1371] = ~((inputs[112]) | (inputs[139]));
    assign layer0_outputs[1372] = (inputs[49]) | (inputs[83]);
    assign layer0_outputs[1373] = ~(inputs[101]);
    assign layer0_outputs[1374] = (inputs[71]) & ~(inputs[175]);
    assign layer0_outputs[1375] = (inputs[225]) | (inputs[116]);
    assign layer0_outputs[1376] = 1'b1;
    assign layer0_outputs[1377] = ~(inputs[229]) | (inputs[94]);
    assign layer0_outputs[1378] = (inputs[72]) & (inputs[138]);
    assign layer0_outputs[1379] = inputs[25];
    assign layer0_outputs[1380] = inputs[115];
    assign layer0_outputs[1381] = ~(inputs[154]);
    assign layer0_outputs[1382] = inputs[44];
    assign layer0_outputs[1383] = (inputs[166]) | (inputs[252]);
    assign layer0_outputs[1384] = ~(inputs[255]) | (inputs[48]);
    assign layer0_outputs[1385] = (inputs[93]) | (inputs[148]);
    assign layer0_outputs[1386] = (inputs[171]) & ~(inputs[77]);
    assign layer0_outputs[1387] = (inputs[94]) ^ (inputs[240]);
    assign layer0_outputs[1388] = ~(inputs[242]);
    assign layer0_outputs[1389] = ~(inputs[52]);
    assign layer0_outputs[1390] = ~((inputs[63]) ^ (inputs[156]));
    assign layer0_outputs[1391] = (inputs[98]) & ~(inputs[170]);
    assign layer0_outputs[1392] = ~(inputs[161]);
    assign layer0_outputs[1393] = inputs[82];
    assign layer0_outputs[1394] = ~((inputs[85]) | (inputs[148]));
    assign layer0_outputs[1395] = ~(inputs[254]);
    assign layer0_outputs[1396] = inputs[16];
    assign layer0_outputs[1397] = ~((inputs[131]) | (inputs[83]));
    assign layer0_outputs[1398] = inputs[122];
    assign layer0_outputs[1399] = (inputs[41]) & ~(inputs[226]);
    assign layer0_outputs[1400] = ~(inputs[121]) | (inputs[252]);
    assign layer0_outputs[1401] = inputs[230];
    assign layer0_outputs[1402] = (inputs[135]) | (inputs[199]);
    assign layer0_outputs[1403] = inputs[197];
    assign layer0_outputs[1404] = ~((inputs[19]) ^ (inputs[85]));
    assign layer0_outputs[1405] = ~((inputs[217]) | (inputs[244]));
    assign layer0_outputs[1406] = ~(inputs[122]) | (inputs[206]);
    assign layer0_outputs[1407] = inputs[76];
    assign layer0_outputs[1408] = 1'b0;
    assign layer0_outputs[1409] = inputs[44];
    assign layer0_outputs[1410] = ~((inputs[30]) & (inputs[210]));
    assign layer0_outputs[1411] = ~((inputs[172]) ^ (inputs[17]));
    assign layer0_outputs[1412] = (inputs[98]) & ~(inputs[140]);
    assign layer0_outputs[1413] = inputs[208];
    assign layer0_outputs[1414] = (inputs[81]) | (inputs[9]);
    assign layer0_outputs[1415] = (inputs[242]) & (inputs[90]);
    assign layer0_outputs[1416] = ~(inputs[243]);
    assign layer0_outputs[1417] = (inputs[226]) ^ (inputs[158]);
    assign layer0_outputs[1418] = (inputs[237]) & ~(inputs[157]);
    assign layer0_outputs[1419] = (inputs[40]) | (inputs[32]);
    assign layer0_outputs[1420] = (inputs[19]) & ~(inputs[66]);
    assign layer0_outputs[1421] = (inputs[50]) & (inputs[234]);
    assign layer0_outputs[1422] = (inputs[9]) | (inputs[165]);
    assign layer0_outputs[1423] = (inputs[247]) | (inputs[144]);
    assign layer0_outputs[1424] = (inputs[142]) ^ (inputs[74]);
    assign layer0_outputs[1425] = (inputs[88]) ^ (inputs[152]);
    assign layer0_outputs[1426] = ~(inputs[101]);
    assign layer0_outputs[1427] = ~(inputs[165]);
    assign layer0_outputs[1428] = ~((inputs[153]) | (inputs[198]));
    assign layer0_outputs[1429] = (inputs[101]) ^ (inputs[206]);
    assign layer0_outputs[1430] = (inputs[193]) ^ (inputs[161]);
    assign layer0_outputs[1431] = ~((inputs[27]) | (inputs[26]));
    assign layer0_outputs[1432] = ~((inputs[252]) | (inputs[7]));
    assign layer0_outputs[1433] = (inputs[225]) | (inputs[227]);
    assign layer0_outputs[1434] = (inputs[163]) & ~(inputs[1]);
    assign layer0_outputs[1435] = ~(inputs[105]);
    assign layer0_outputs[1436] = ~(inputs[246]);
    assign layer0_outputs[1437] = inputs[209];
    assign layer0_outputs[1438] = inputs[240];
    assign layer0_outputs[1439] = ~(inputs[178]) | (inputs[47]);
    assign layer0_outputs[1440] = ~(inputs[187]) | (inputs[67]);
    assign layer0_outputs[1441] = ~(inputs[130]);
    assign layer0_outputs[1442] = (inputs[105]) & ~(inputs[95]);
    assign layer0_outputs[1443] = ~((inputs[111]) ^ (inputs[200]));
    assign layer0_outputs[1444] = (inputs[29]) | (inputs[120]);
    assign layer0_outputs[1445] = inputs[43];
    assign layer0_outputs[1446] = inputs[30];
    assign layer0_outputs[1447] = (inputs[154]) & ~(inputs[65]);
    assign layer0_outputs[1448] = 1'b1;
    assign layer0_outputs[1449] = ~((inputs[232]) ^ (inputs[22]));
    assign layer0_outputs[1450] = (inputs[124]) | (inputs[189]);
    assign layer0_outputs[1451] = ~((inputs[56]) ^ (inputs[59]));
    assign layer0_outputs[1452] = 1'b0;
    assign layer0_outputs[1453] = (inputs[85]) ^ (inputs[253]);
    assign layer0_outputs[1454] = ~(inputs[245]) | (inputs[17]);
    assign layer0_outputs[1455] = ~(inputs[214]);
    assign layer0_outputs[1456] = ~(inputs[166]);
    assign layer0_outputs[1457] = ~((inputs[91]) ^ (inputs[105]));
    assign layer0_outputs[1458] = (inputs[111]) & (inputs[218]);
    assign layer0_outputs[1459] = ~(inputs[117]);
    assign layer0_outputs[1460] = inputs[7];
    assign layer0_outputs[1461] = ~(inputs[76]) | (inputs[212]);
    assign layer0_outputs[1462] = (inputs[12]) | (inputs[50]);
    assign layer0_outputs[1463] = ~((inputs[144]) | (inputs[165]));
    assign layer0_outputs[1464] = 1'b1;
    assign layer0_outputs[1465] = inputs[118];
    assign layer0_outputs[1466] = ~(inputs[14]) | (inputs[221]);
    assign layer0_outputs[1467] = ~((inputs[21]) | (inputs[84]));
    assign layer0_outputs[1468] = 1'b1;
    assign layer0_outputs[1469] = ~(inputs[174]);
    assign layer0_outputs[1470] = ~((inputs[211]) ^ (inputs[128]));
    assign layer0_outputs[1471] = inputs[121];
    assign layer0_outputs[1472] = ~((inputs[206]) | (inputs[86]));
    assign layer0_outputs[1473] = (inputs[168]) ^ (inputs[161]);
    assign layer0_outputs[1474] = (inputs[50]) & (inputs[159]);
    assign layer0_outputs[1475] = ~(inputs[71]);
    assign layer0_outputs[1476] = ~(inputs[232]) | (inputs[125]);
    assign layer0_outputs[1477] = (inputs[222]) & ~(inputs[55]);
    assign layer0_outputs[1478] = (inputs[188]) & ~(inputs[36]);
    assign layer0_outputs[1479] = (inputs[229]) & ~(inputs[131]);
    assign layer0_outputs[1480] = ~(inputs[77]);
    assign layer0_outputs[1481] = ~(inputs[173]) | (inputs[113]);
    assign layer0_outputs[1482] = (inputs[57]) & ~(inputs[20]);
    assign layer0_outputs[1483] = ~((inputs[185]) | (inputs[142]));
    assign layer0_outputs[1484] = (inputs[201]) ^ (inputs[31]);
    assign layer0_outputs[1485] = ~((inputs[195]) & (inputs[156]));
    assign layer0_outputs[1486] = inputs[85];
    assign layer0_outputs[1487] = (inputs[170]) ^ (inputs[226]);
    assign layer0_outputs[1488] = ~(inputs[75]);
    assign layer0_outputs[1489] = inputs[224];
    assign layer0_outputs[1490] = ~(inputs[252]);
    assign layer0_outputs[1491] = (inputs[27]) & ~(inputs[163]);
    assign layer0_outputs[1492] = (inputs[115]) & ~(inputs[226]);
    assign layer0_outputs[1493] = ~(inputs[79]);
    assign layer0_outputs[1494] = ~((inputs[254]) ^ (inputs[182]));
    assign layer0_outputs[1495] = ~((inputs[151]) & (inputs[41]));
    assign layer0_outputs[1496] = ~(inputs[100]);
    assign layer0_outputs[1497] = (inputs[148]) | (inputs[117]);
    assign layer0_outputs[1498] = ~(inputs[90]);
    assign layer0_outputs[1499] = ~((inputs[19]) ^ (inputs[232]));
    assign layer0_outputs[1500] = (inputs[138]) & ~(inputs[2]);
    assign layer0_outputs[1501] = (inputs[13]) & ~(inputs[244]);
    assign layer0_outputs[1502] = ~(inputs[115]);
    assign layer0_outputs[1503] = ~((inputs[252]) ^ (inputs[182]));
    assign layer0_outputs[1504] = ~((inputs[192]) | (inputs[12]));
    assign layer0_outputs[1505] = (inputs[182]) & ~(inputs[108]);
    assign layer0_outputs[1506] = ~((inputs[79]) | (inputs[187]));
    assign layer0_outputs[1507] = inputs[226];
    assign layer0_outputs[1508] = inputs[201];
    assign layer0_outputs[1509] = (inputs[85]) & ~(inputs[5]);
    assign layer0_outputs[1510] = inputs[233];
    assign layer0_outputs[1511] = (inputs[48]) ^ (inputs[186]);
    assign layer0_outputs[1512] = 1'b1;
    assign layer0_outputs[1513] = (inputs[49]) | (inputs[35]);
    assign layer0_outputs[1514] = ~(inputs[114]) | (inputs[65]);
    assign layer0_outputs[1515] = inputs[103];
    assign layer0_outputs[1516] = ~((inputs[126]) | (inputs[18]));
    assign layer0_outputs[1517] = (inputs[121]) | (inputs[133]);
    assign layer0_outputs[1518] = ~((inputs[255]) ^ (inputs[93]));
    assign layer0_outputs[1519] = ~(inputs[69]) | (inputs[243]);
    assign layer0_outputs[1520] = (inputs[192]) ^ (inputs[246]);
    assign layer0_outputs[1521] = ~(inputs[80]) | (inputs[73]);
    assign layer0_outputs[1522] = 1'b1;
    assign layer0_outputs[1523] = (inputs[205]) ^ (inputs[4]);
    assign layer0_outputs[1524] = ~(inputs[237]) | (inputs[103]);
    assign layer0_outputs[1525] = (inputs[5]) & ~(inputs[250]);
    assign layer0_outputs[1526] = ~((inputs[147]) | (inputs[52]));
    assign layer0_outputs[1527] = (inputs[61]) & ~(inputs[114]);
    assign layer0_outputs[1528] = ~((inputs[42]) & (inputs[21]));
    assign layer0_outputs[1529] = ~((inputs[148]) ^ (inputs[108]));
    assign layer0_outputs[1530] = ~((inputs[35]) | (inputs[223]));
    assign layer0_outputs[1531] = (inputs[123]) | (inputs[178]);
    assign layer0_outputs[1532] = (inputs[184]) & (inputs[251]);
    assign layer0_outputs[1533] = (inputs[81]) | (inputs[91]);
    assign layer0_outputs[1534] = ~(inputs[67]);
    assign layer0_outputs[1535] = ~(inputs[196]) | (inputs[91]);
    assign layer0_outputs[1536] = ~(inputs[79]);
    assign layer0_outputs[1537] = inputs[152];
    assign layer0_outputs[1538] = (inputs[29]) & ~(inputs[255]);
    assign layer0_outputs[1539] = (inputs[86]) & ~(inputs[94]);
    assign layer0_outputs[1540] = (inputs[211]) ^ (inputs[119]);
    assign layer0_outputs[1541] = ~((inputs[28]) & (inputs[205]));
    assign layer0_outputs[1542] = (inputs[26]) & ~(inputs[249]);
    assign layer0_outputs[1543] = ~((inputs[46]) | (inputs[9]));
    assign layer0_outputs[1544] = (inputs[218]) & ~(inputs[190]);
    assign layer0_outputs[1545] = inputs[29];
    assign layer0_outputs[1546] = ~(inputs[89]);
    assign layer0_outputs[1547] = ~(inputs[218]);
    assign layer0_outputs[1548] = ~(inputs[214]);
    assign layer0_outputs[1549] = (inputs[175]) | (inputs[56]);
    assign layer0_outputs[1550] = (inputs[176]) | (inputs[177]);
    assign layer0_outputs[1551] = (inputs[116]) ^ (inputs[196]);
    assign layer0_outputs[1552] = ~(inputs[238]);
    assign layer0_outputs[1553] = ~(inputs[51]) | (inputs[2]);
    assign layer0_outputs[1554] = (inputs[113]) & ~(inputs[78]);
    assign layer0_outputs[1555] = (inputs[214]) ^ (inputs[242]);
    assign layer0_outputs[1556] = ~((inputs[161]) ^ (inputs[22]));
    assign layer0_outputs[1557] = ~(inputs[76]);
    assign layer0_outputs[1558] = (inputs[44]) & ~(inputs[25]);
    assign layer0_outputs[1559] = (inputs[77]) | (inputs[228]);
    assign layer0_outputs[1560] = (inputs[17]) ^ (inputs[97]);
    assign layer0_outputs[1561] = (inputs[19]) & ~(inputs[176]);
    assign layer0_outputs[1562] = inputs[11];
    assign layer0_outputs[1563] = ~(inputs[179]);
    assign layer0_outputs[1564] = (inputs[58]) ^ (inputs[233]);
    assign layer0_outputs[1565] = inputs[176];
    assign layer0_outputs[1566] = ~(inputs[201]);
    assign layer0_outputs[1567] = (inputs[64]) & ~(inputs[20]);
    assign layer0_outputs[1568] = ~((inputs[248]) | (inputs[81]));
    assign layer0_outputs[1569] = inputs[226];
    assign layer0_outputs[1570] = ~((inputs[76]) | (inputs[81]));
    assign layer0_outputs[1571] = (inputs[255]) ^ (inputs[225]);
    assign layer0_outputs[1572] = ~(inputs[84]);
    assign layer0_outputs[1573] = (inputs[196]) & ~(inputs[46]);
    assign layer0_outputs[1574] = ~(inputs[56]) | (inputs[70]);
    assign layer0_outputs[1575] = (inputs[41]) & ~(inputs[87]);
    assign layer0_outputs[1576] = ~(inputs[212]) | (inputs[198]);
    assign layer0_outputs[1577] = ~(inputs[7]);
    assign layer0_outputs[1578] = (inputs[137]) & ~(inputs[218]);
    assign layer0_outputs[1579] = (inputs[182]) & ~(inputs[107]);
    assign layer0_outputs[1580] = ~((inputs[51]) | (inputs[93]));
    assign layer0_outputs[1581] = (inputs[206]) & ~(inputs[239]);
    assign layer0_outputs[1582] = ~(inputs[55]);
    assign layer0_outputs[1583] = ~(inputs[41]) | (inputs[128]);
    assign layer0_outputs[1584] = ~(inputs[11]);
    assign layer0_outputs[1585] = (inputs[61]) | (inputs[119]);
    assign layer0_outputs[1586] = (inputs[145]) | (inputs[3]);
    assign layer0_outputs[1587] = (inputs[74]) & ~(inputs[204]);
    assign layer0_outputs[1588] = inputs[211];
    assign layer0_outputs[1589] = ~(inputs[150]);
    assign layer0_outputs[1590] = (inputs[174]) & ~(inputs[127]);
    assign layer0_outputs[1591] = 1'b1;
    assign layer0_outputs[1592] = (inputs[148]) ^ (inputs[247]);
    assign layer0_outputs[1593] = inputs[159];
    assign layer0_outputs[1594] = ~((inputs[153]) | (inputs[13]));
    assign layer0_outputs[1595] = ~(inputs[188]) | (inputs[232]);
    assign layer0_outputs[1596] = ~((inputs[151]) | (inputs[3]));
    assign layer0_outputs[1597] = inputs[130];
    assign layer0_outputs[1598] = inputs[146];
    assign layer0_outputs[1599] = (inputs[37]) ^ (inputs[73]);
    assign layer0_outputs[1600] = (inputs[135]) | (inputs[146]);
    assign layer0_outputs[1601] = (inputs[210]) & ~(inputs[16]);
    assign layer0_outputs[1602] = ~((inputs[229]) | (inputs[84]));
    assign layer0_outputs[1603] = (inputs[127]) | (inputs[190]);
    assign layer0_outputs[1604] = ~(inputs[217]) | (inputs[113]);
    assign layer0_outputs[1605] = (inputs[185]) ^ (inputs[246]);
    assign layer0_outputs[1606] = (inputs[154]) ^ (inputs[19]);
    assign layer0_outputs[1607] = ~((inputs[229]) | (inputs[213]));
    assign layer0_outputs[1608] = (inputs[124]) | (inputs[19]);
    assign layer0_outputs[1609] = ~((inputs[52]) | (inputs[2]));
    assign layer0_outputs[1610] = ~(inputs[205]);
    assign layer0_outputs[1611] = ~(inputs[21]) | (inputs[102]);
    assign layer0_outputs[1612] = ~((inputs[51]) | (inputs[66]));
    assign layer0_outputs[1613] = inputs[169];
    assign layer0_outputs[1614] = (inputs[198]) & (inputs[60]);
    assign layer0_outputs[1615] = ~(inputs[10]);
    assign layer0_outputs[1616] = inputs[244];
    assign layer0_outputs[1617] = ~(inputs[212]) | (inputs[95]);
    assign layer0_outputs[1618] = ~(inputs[89]) | (inputs[34]);
    assign layer0_outputs[1619] = (inputs[115]) & ~(inputs[93]);
    assign layer0_outputs[1620] = (inputs[58]) | (inputs[20]);
    assign layer0_outputs[1621] = ~((inputs[154]) & (inputs[176]));
    assign layer0_outputs[1622] = ~(inputs[44]);
    assign layer0_outputs[1623] = ~((inputs[249]) | (inputs[211]));
    assign layer0_outputs[1624] = (inputs[47]) | (inputs[138]);
    assign layer0_outputs[1625] = inputs[97];
    assign layer0_outputs[1626] = (inputs[90]) | (inputs[17]);
    assign layer0_outputs[1627] = inputs[99];
    assign layer0_outputs[1628] = ~(inputs[140]);
    assign layer0_outputs[1629] = inputs[182];
    assign layer0_outputs[1630] = ~(inputs[0]);
    assign layer0_outputs[1631] = inputs[173];
    assign layer0_outputs[1632] = inputs[221];
    assign layer0_outputs[1633] = (inputs[64]) | (inputs[233]);
    assign layer0_outputs[1634] = (inputs[150]) & (inputs[86]);
    assign layer0_outputs[1635] = ~(inputs[188]);
    assign layer0_outputs[1636] = inputs[193];
    assign layer0_outputs[1637] = (inputs[80]) ^ (inputs[248]);
    assign layer0_outputs[1638] = (inputs[194]) & ~(inputs[13]);
    assign layer0_outputs[1639] = (inputs[2]) ^ (inputs[192]);
    assign layer0_outputs[1640] = ~((inputs[32]) | (inputs[190]));
    assign layer0_outputs[1641] = ~(inputs[161]);
    assign layer0_outputs[1642] = inputs[230];
    assign layer0_outputs[1643] = ~(inputs[122]) | (inputs[33]);
    assign layer0_outputs[1644] = ~((inputs[245]) | (inputs[218]));
    assign layer0_outputs[1645] = (inputs[121]) & ~(inputs[84]);
    assign layer0_outputs[1646] = (inputs[11]) & ~(inputs[81]);
    assign layer0_outputs[1647] = inputs[97];
    assign layer0_outputs[1648] = ~((inputs[15]) | (inputs[73]));
    assign layer0_outputs[1649] = inputs[91];
    assign layer0_outputs[1650] = (inputs[151]) | (inputs[135]);
    assign layer0_outputs[1651] = ~((inputs[49]) | (inputs[36]));
    assign layer0_outputs[1652] = inputs[74];
    assign layer0_outputs[1653] = ~((inputs[17]) | (inputs[148]));
    assign layer0_outputs[1654] = inputs[136];
    assign layer0_outputs[1655] = inputs[151];
    assign layer0_outputs[1656] = (inputs[143]) & ~(inputs[50]);
    assign layer0_outputs[1657] = ~((inputs[234]) | (inputs[206]));
    assign layer0_outputs[1658] = ~(inputs[153]);
    assign layer0_outputs[1659] = ~((inputs[252]) ^ (inputs[53]));
    assign layer0_outputs[1660] = inputs[117];
    assign layer0_outputs[1661] = ~((inputs[47]) | (inputs[40]));
    assign layer0_outputs[1662] = ~((inputs[222]) | (inputs[220]));
    assign layer0_outputs[1663] = (inputs[28]) & ~(inputs[202]);
    assign layer0_outputs[1664] = inputs[156];
    assign layer0_outputs[1665] = ~(inputs[228]);
    assign layer0_outputs[1666] = (inputs[37]) & ~(inputs[214]);
    assign layer0_outputs[1667] = 1'b0;
    assign layer0_outputs[1668] = (inputs[181]) | (inputs[48]);
    assign layer0_outputs[1669] = (inputs[188]) | (inputs[145]);
    assign layer0_outputs[1670] = (inputs[22]) & ~(inputs[159]);
    assign layer0_outputs[1671] = ~(inputs[7]) | (inputs[29]);
    assign layer0_outputs[1672] = ~(inputs[174]);
    assign layer0_outputs[1673] = inputs[107];
    assign layer0_outputs[1674] = (inputs[182]) & ~(inputs[192]);
    assign layer0_outputs[1675] = ~((inputs[161]) ^ (inputs[163]));
    assign layer0_outputs[1676] = ~(inputs[148]);
    assign layer0_outputs[1677] = ~(inputs[200]) | (inputs[125]);
    assign layer0_outputs[1678] = (inputs[238]) ^ (inputs[204]);
    assign layer0_outputs[1679] = (inputs[27]) ^ (inputs[109]);
    assign layer0_outputs[1680] = (inputs[48]) | (inputs[162]);
    assign layer0_outputs[1681] = (inputs[152]) | (inputs[107]);
    assign layer0_outputs[1682] = (inputs[138]) ^ (inputs[188]);
    assign layer0_outputs[1683] = 1'b0;
    assign layer0_outputs[1684] = (inputs[73]) & ~(inputs[14]);
    assign layer0_outputs[1685] = inputs[221];
    assign layer0_outputs[1686] = (inputs[127]) | (inputs[94]);
    assign layer0_outputs[1687] = ~(inputs[182]);
    assign layer0_outputs[1688] = ~(inputs[205]);
    assign layer0_outputs[1689] = (inputs[161]) ^ (inputs[69]);
    assign layer0_outputs[1690] = ~(inputs[62]);
    assign layer0_outputs[1691] = ~(inputs[73]) | (inputs[34]);
    assign layer0_outputs[1692] = inputs[136];
    assign layer0_outputs[1693] = ~((inputs[189]) ^ (inputs[113]));
    assign layer0_outputs[1694] = ~(inputs[217]);
    assign layer0_outputs[1695] = inputs[105];
    assign layer0_outputs[1696] = (inputs[183]) & ~(inputs[91]);
    assign layer0_outputs[1697] = (inputs[22]) & ~(inputs[79]);
    assign layer0_outputs[1698] = inputs[140];
    assign layer0_outputs[1699] = ~(inputs[98]);
    assign layer0_outputs[1700] = ~((inputs[188]) ^ (inputs[16]));
    assign layer0_outputs[1701] = (inputs[110]) & ~(inputs[226]);
    assign layer0_outputs[1702] = 1'b0;
    assign layer0_outputs[1703] = ~((inputs[3]) ^ (inputs[49]));
    assign layer0_outputs[1704] = ~((inputs[238]) | (inputs[94]));
    assign layer0_outputs[1705] = ~((inputs[33]) | (inputs[186]));
    assign layer0_outputs[1706] = inputs[14];
    assign layer0_outputs[1707] = (inputs[19]) & ~(inputs[82]);
    assign layer0_outputs[1708] = (inputs[20]) & (inputs[223]);
    assign layer0_outputs[1709] = ~(inputs[227]) | (inputs[26]);
    assign layer0_outputs[1710] = ~(inputs[4]);
    assign layer0_outputs[1711] = (inputs[59]) | (inputs[70]);
    assign layer0_outputs[1712] = inputs[215];
    assign layer0_outputs[1713] = inputs[107];
    assign layer0_outputs[1714] = ~((inputs[150]) | (inputs[238]));
    assign layer0_outputs[1715] = (inputs[68]) & ~(inputs[112]);
    assign layer0_outputs[1716] = ~(inputs[14]);
    assign layer0_outputs[1717] = inputs[14];
    assign layer0_outputs[1718] = ~(inputs[50]);
    assign layer0_outputs[1719] = (inputs[89]) & ~(inputs[226]);
    assign layer0_outputs[1720] = 1'b1;
    assign layer0_outputs[1721] = ~((inputs[220]) | (inputs[178]));
    assign layer0_outputs[1722] = (inputs[221]) | (inputs[33]);
    assign layer0_outputs[1723] = (inputs[179]) & ~(inputs[144]);
    assign layer0_outputs[1724] = (inputs[158]) & ~(inputs[185]);
    assign layer0_outputs[1725] = (inputs[94]) ^ (inputs[75]);
    assign layer0_outputs[1726] = (inputs[156]) & ~(inputs[41]);
    assign layer0_outputs[1727] = (inputs[78]) ^ (inputs[108]);
    assign layer0_outputs[1728] = ~(inputs[189]) | (inputs[211]);
    assign layer0_outputs[1729] = inputs[250];
    assign layer0_outputs[1730] = (inputs[161]) | (inputs[221]);
    assign layer0_outputs[1731] = ~(inputs[121]) | (inputs[209]);
    assign layer0_outputs[1732] = ~((inputs[69]) & (inputs[203]));
    assign layer0_outputs[1733] = (inputs[127]) | (inputs[122]);
    assign layer0_outputs[1734] = inputs[92];
    assign layer0_outputs[1735] = ~(inputs[12]) | (inputs[161]);
    assign layer0_outputs[1736] = (inputs[196]) ^ (inputs[32]);
    assign layer0_outputs[1737] = (inputs[49]) ^ (inputs[53]);
    assign layer0_outputs[1738] = inputs[176];
    assign layer0_outputs[1739] = ~((inputs[137]) ^ (inputs[190]));
    assign layer0_outputs[1740] = inputs[129];
    assign layer0_outputs[1741] = (inputs[74]) | (inputs[1]);
    assign layer0_outputs[1742] = (inputs[200]) & ~(inputs[94]);
    assign layer0_outputs[1743] = ~(inputs[212]) | (inputs[75]);
    assign layer0_outputs[1744] = inputs[25];
    assign layer0_outputs[1745] = inputs[92];
    assign layer0_outputs[1746] = (inputs[44]) & ~(inputs[186]);
    assign layer0_outputs[1747] = ~(inputs[171]);
    assign layer0_outputs[1748] = ~(inputs[228]);
    assign layer0_outputs[1749] = ~(inputs[67]);
    assign layer0_outputs[1750] = inputs[190];
    assign layer0_outputs[1751] = (inputs[12]) & ~(inputs[35]);
    assign layer0_outputs[1752] = (inputs[38]) | (inputs[155]);
    assign layer0_outputs[1753] = ~(inputs[105]);
    assign layer0_outputs[1754] = ~(inputs[183]);
    assign layer0_outputs[1755] = inputs[57];
    assign layer0_outputs[1756] = (inputs[2]) ^ (inputs[237]);
    assign layer0_outputs[1757] = ~(inputs[150]) | (inputs[170]);
    assign layer0_outputs[1758] = 1'b1;
    assign layer0_outputs[1759] = ~(inputs[129]) | (inputs[72]);
    assign layer0_outputs[1760] = inputs[21];
    assign layer0_outputs[1761] = ~((inputs[119]) | (inputs[34]));
    assign layer0_outputs[1762] = (inputs[25]) | (inputs[10]);
    assign layer0_outputs[1763] = (inputs[253]) | (inputs[89]);
    assign layer0_outputs[1764] = (inputs[10]) & ~(inputs[215]);
    assign layer0_outputs[1765] = (inputs[128]) | (inputs[191]);
    assign layer0_outputs[1766] = ~((inputs[52]) | (inputs[218]));
    assign layer0_outputs[1767] = inputs[167];
    assign layer0_outputs[1768] = ~(inputs[221]) | (inputs[158]);
    assign layer0_outputs[1769] = ~((inputs[42]) ^ (inputs[50]));
    assign layer0_outputs[1770] = ~(inputs[224]) | (inputs[26]);
    assign layer0_outputs[1771] = inputs[129];
    assign layer0_outputs[1772] = ~(inputs[151]);
    assign layer0_outputs[1773] = ~(inputs[105]) | (inputs[190]);
    assign layer0_outputs[1774] = (inputs[44]) | (inputs[204]);
    assign layer0_outputs[1775] = inputs[145];
    assign layer0_outputs[1776] = inputs[210];
    assign layer0_outputs[1777] = 1'b1;
    assign layer0_outputs[1778] = ~(inputs[62]);
    assign layer0_outputs[1779] = ~(inputs[198]) | (inputs[39]);
    assign layer0_outputs[1780] = ~(inputs[58]) | (inputs[239]);
    assign layer0_outputs[1781] = ~((inputs[102]) ^ (inputs[23]));
    assign layer0_outputs[1782] = ~((inputs[141]) ^ (inputs[81]));
    assign layer0_outputs[1783] = inputs[212];
    assign layer0_outputs[1784] = ~((inputs[173]) ^ (inputs[25]));
    assign layer0_outputs[1785] = ~((inputs[209]) ^ (inputs[239]));
    assign layer0_outputs[1786] = ~(inputs[11]) | (inputs[218]);
    assign layer0_outputs[1787] = (inputs[82]) | (inputs[195]);
    assign layer0_outputs[1788] = ~(inputs[178]) | (inputs[17]);
    assign layer0_outputs[1789] = (inputs[102]) & (inputs[66]);
    assign layer0_outputs[1790] = (inputs[180]) & ~(inputs[114]);
    assign layer0_outputs[1791] = ~(inputs[38]);
    assign layer0_outputs[1792] = 1'b0;
    assign layer0_outputs[1793] = (inputs[117]) ^ (inputs[189]);
    assign layer0_outputs[1794] = inputs[147];
    assign layer0_outputs[1795] = ~(inputs[130]);
    assign layer0_outputs[1796] = inputs[147];
    assign layer0_outputs[1797] = ~((inputs[77]) | (inputs[84]));
    assign layer0_outputs[1798] = (inputs[191]) | (inputs[189]);
    assign layer0_outputs[1799] = ~(inputs[179]);
    assign layer0_outputs[1800] = ~(inputs[51]);
    assign layer0_outputs[1801] = ~((inputs[82]) & (inputs[71]));
    assign layer0_outputs[1802] = 1'b1;
    assign layer0_outputs[1803] = (inputs[224]) | (inputs[174]);
    assign layer0_outputs[1804] = inputs[29];
    assign layer0_outputs[1805] = ~((inputs[101]) | (inputs[99]));
    assign layer0_outputs[1806] = ~(inputs[210]) | (inputs[74]);
    assign layer0_outputs[1807] = ~((inputs[61]) | (inputs[104]));
    assign layer0_outputs[1808] = inputs[213];
    assign layer0_outputs[1809] = (inputs[20]) ^ (inputs[112]);
    assign layer0_outputs[1810] = inputs[28];
    assign layer0_outputs[1811] = ~((inputs[51]) ^ (inputs[196]));
    assign layer0_outputs[1812] = (inputs[137]) ^ (inputs[171]);
    assign layer0_outputs[1813] = ~((inputs[167]) | (inputs[2]));
    assign layer0_outputs[1814] = (inputs[111]) ^ (inputs[84]);
    assign layer0_outputs[1815] = (inputs[6]) & (inputs[127]);
    assign layer0_outputs[1816] = (inputs[244]) & ~(inputs[4]);
    assign layer0_outputs[1817] = inputs[101];
    assign layer0_outputs[1818] = ~((inputs[142]) | (inputs[218]));
    assign layer0_outputs[1819] = ~(inputs[230]);
    assign layer0_outputs[1820] = ~((inputs[94]) | (inputs[170]));
    assign layer0_outputs[1821] = ~((inputs[70]) ^ (inputs[205]));
    assign layer0_outputs[1822] = ~((inputs[42]) | (inputs[227]));
    assign layer0_outputs[1823] = inputs[202];
    assign layer0_outputs[1824] = ~((inputs[0]) | (inputs[69]));
    assign layer0_outputs[1825] = (inputs[163]) ^ (inputs[110]);
    assign layer0_outputs[1826] = ~(inputs[231]) | (inputs[48]);
    assign layer0_outputs[1827] = ~(inputs[138]) | (inputs[205]);
    assign layer0_outputs[1828] = inputs[119];
    assign layer0_outputs[1829] = inputs[221];
    assign layer0_outputs[1830] = ~((inputs[46]) | (inputs[93]));
    assign layer0_outputs[1831] = ~((inputs[92]) | (inputs[78]));
    assign layer0_outputs[1832] = ~(inputs[166]);
    assign layer0_outputs[1833] = inputs[129];
    assign layer0_outputs[1834] = inputs[83];
    assign layer0_outputs[1835] = (inputs[191]) | (inputs[216]);
    assign layer0_outputs[1836] = (inputs[26]) & ~(inputs[184]);
    assign layer0_outputs[1837] = (inputs[96]) | (inputs[237]);
    assign layer0_outputs[1838] = (inputs[196]) | (inputs[187]);
    assign layer0_outputs[1839] = ~((inputs[246]) ^ (inputs[79]));
    assign layer0_outputs[1840] = ~((inputs[217]) & (inputs[44]));
    assign layer0_outputs[1841] = ~(inputs[22]);
    assign layer0_outputs[1842] = ~((inputs[212]) | (inputs[41]));
    assign layer0_outputs[1843] = ~(inputs[90]);
    assign layer0_outputs[1844] = (inputs[65]) | (inputs[47]);
    assign layer0_outputs[1845] = ~(inputs[127]);
    assign layer0_outputs[1846] = ~(inputs[145]) | (inputs[13]);
    assign layer0_outputs[1847] = ~((inputs[235]) | (inputs[217]));
    assign layer0_outputs[1848] = ~((inputs[96]) ^ (inputs[118]));
    assign layer0_outputs[1849] = inputs[118];
    assign layer0_outputs[1850] = ~((inputs[138]) | (inputs[241]));
    assign layer0_outputs[1851] = inputs[165];
    assign layer0_outputs[1852] = ~(inputs[22]);
    assign layer0_outputs[1853] = inputs[170];
    assign layer0_outputs[1854] = ~((inputs[20]) ^ (inputs[65]));
    assign layer0_outputs[1855] = (inputs[205]) ^ (inputs[151]);
    assign layer0_outputs[1856] = ~((inputs[18]) | (inputs[18]));
    assign layer0_outputs[1857] = ~((inputs[202]) | (inputs[243]));
    assign layer0_outputs[1858] = ~(inputs[137]);
    assign layer0_outputs[1859] = (inputs[163]) & (inputs[117]);
    assign layer0_outputs[1860] = ~((inputs[69]) ^ (inputs[68]));
    assign layer0_outputs[1861] = inputs[197];
    assign layer0_outputs[1862] = ~(inputs[98]);
    assign layer0_outputs[1863] = (inputs[182]) | (inputs[0]);
    assign layer0_outputs[1864] = inputs[79];
    assign layer0_outputs[1865] = (inputs[169]) & (inputs[81]);
    assign layer0_outputs[1866] = inputs[234];
    assign layer0_outputs[1867] = ~((inputs[42]) & (inputs[39]));
    assign layer0_outputs[1868] = ~(inputs[58]) | (inputs[71]);
    assign layer0_outputs[1869] = inputs[133];
    assign layer0_outputs[1870] = ~(inputs[179]) | (inputs[112]);
    assign layer0_outputs[1871] = ~(inputs[225]);
    assign layer0_outputs[1872] = ~(inputs[9]);
    assign layer0_outputs[1873] = ~(inputs[147]);
    assign layer0_outputs[1874] = ~((inputs[58]) | (inputs[127]));
    assign layer0_outputs[1875] = inputs[216];
    assign layer0_outputs[1876] = inputs[161];
    assign layer0_outputs[1877] = inputs[133];
    assign layer0_outputs[1878] = inputs[39];
    assign layer0_outputs[1879] = ~((inputs[97]) ^ (inputs[149]));
    assign layer0_outputs[1880] = ~((inputs[251]) & (inputs[111]));
    assign layer0_outputs[1881] = (inputs[44]) ^ (inputs[76]);
    assign layer0_outputs[1882] = (inputs[59]) & ~(inputs[38]);
    assign layer0_outputs[1883] = (inputs[117]) & (inputs[68]);
    assign layer0_outputs[1884] = (inputs[118]) ^ (inputs[215]);
    assign layer0_outputs[1885] = ~((inputs[92]) ^ (inputs[74]));
    assign layer0_outputs[1886] = inputs[7];
    assign layer0_outputs[1887] = (inputs[20]) & ~(inputs[11]);
    assign layer0_outputs[1888] = (inputs[136]) & ~(inputs[91]);
    assign layer0_outputs[1889] = (inputs[175]) & ~(inputs[138]);
    assign layer0_outputs[1890] = ~((inputs[32]) ^ (inputs[245]));
    assign layer0_outputs[1891] = (inputs[156]) & ~(inputs[95]);
    assign layer0_outputs[1892] = ~((inputs[246]) ^ (inputs[92]));
    assign layer0_outputs[1893] = ~(inputs[149]) | (inputs[78]);
    assign layer0_outputs[1894] = ~(inputs[52]);
    assign layer0_outputs[1895] = ~(inputs[74]);
    assign layer0_outputs[1896] = ~((inputs[108]) ^ (inputs[144]));
    assign layer0_outputs[1897] = (inputs[180]) & ~(inputs[142]);
    assign layer0_outputs[1898] = ~((inputs[228]) & (inputs[173]));
    assign layer0_outputs[1899] = inputs[146];
    assign layer0_outputs[1900] = ~((inputs[88]) ^ (inputs[167]));
    assign layer0_outputs[1901] = ~((inputs[11]) | (inputs[79]));
    assign layer0_outputs[1902] = (inputs[154]) & ~(inputs[236]);
    assign layer0_outputs[1903] = (inputs[56]) & ~(inputs[186]);
    assign layer0_outputs[1904] = ~(inputs[54]);
    assign layer0_outputs[1905] = (inputs[55]) & ~(inputs[171]);
    assign layer0_outputs[1906] = ~(inputs[152]) | (inputs[66]);
    assign layer0_outputs[1907] = inputs[230];
    assign layer0_outputs[1908] = ~(inputs[230]);
    assign layer0_outputs[1909] = ~(inputs[13]);
    assign layer0_outputs[1910] = ~(inputs[101]);
    assign layer0_outputs[1911] = inputs[186];
    assign layer0_outputs[1912] = ~((inputs[96]) | (inputs[100]));
    assign layer0_outputs[1913] = inputs[233];
    assign layer0_outputs[1914] = ~(inputs[39]);
    assign layer0_outputs[1915] = ~(inputs[77]) | (inputs[158]);
    assign layer0_outputs[1916] = ~(inputs[149]) | (inputs[35]);
    assign layer0_outputs[1917] = ~((inputs[156]) ^ (inputs[206]));
    assign layer0_outputs[1918] = (inputs[153]) & ~(inputs[98]);
    assign layer0_outputs[1919] = inputs[135];
    assign layer0_outputs[1920] = inputs[170];
    assign layer0_outputs[1921] = (inputs[222]) ^ (inputs[228]);
    assign layer0_outputs[1922] = inputs[193];
    assign layer0_outputs[1923] = inputs[25];
    assign layer0_outputs[1924] = (inputs[113]) ^ (inputs[99]);
    assign layer0_outputs[1925] = ~((inputs[238]) | (inputs[29]));
    assign layer0_outputs[1926] = (inputs[125]) | (inputs[250]);
    assign layer0_outputs[1927] = inputs[75];
    assign layer0_outputs[1928] = inputs[108];
    assign layer0_outputs[1929] = (inputs[255]) ^ (inputs[10]);
    assign layer0_outputs[1930] = ~((inputs[220]) | (inputs[170]));
    assign layer0_outputs[1931] = ~((inputs[184]) ^ (inputs[233]));
    assign layer0_outputs[1932] = (inputs[150]) ^ (inputs[47]);
    assign layer0_outputs[1933] = ~((inputs[126]) | (inputs[82]));
    assign layer0_outputs[1934] = inputs[102];
    assign layer0_outputs[1935] = ~(inputs[78]);
    assign layer0_outputs[1936] = ~((inputs[193]) | (inputs[210]));
    assign layer0_outputs[1937] = (inputs[89]) ^ (inputs[152]);
    assign layer0_outputs[1938] = ~((inputs[108]) | (inputs[84]));
    assign layer0_outputs[1939] = (inputs[244]) & ~(inputs[96]);
    assign layer0_outputs[1940] = ~((inputs[58]) ^ (inputs[179]));
    assign layer0_outputs[1941] = inputs[253];
    assign layer0_outputs[1942] = ~((inputs[244]) & (inputs[31]));
    assign layer0_outputs[1943] = (inputs[27]) & ~(inputs[17]);
    assign layer0_outputs[1944] = (inputs[182]) & ~(inputs[190]);
    assign layer0_outputs[1945] = 1'b0;
    assign layer0_outputs[1946] = inputs[132];
    assign layer0_outputs[1947] = ~(inputs[156]);
    assign layer0_outputs[1948] = ~((inputs[97]) & (inputs[154]));
    assign layer0_outputs[1949] = ~((inputs[53]) ^ (inputs[92]));
    assign layer0_outputs[1950] = (inputs[194]) ^ (inputs[241]);
    assign layer0_outputs[1951] = inputs[237];
    assign layer0_outputs[1952] = (inputs[120]) ^ (inputs[25]);
    assign layer0_outputs[1953] = ~((inputs[233]) ^ (inputs[185]));
    assign layer0_outputs[1954] = ~(inputs[112]);
    assign layer0_outputs[1955] = (inputs[200]) & (inputs[165]);
    assign layer0_outputs[1956] = (inputs[103]) & ~(inputs[77]);
    assign layer0_outputs[1957] = ~(inputs[253]) | (inputs[43]);
    assign layer0_outputs[1958] = (inputs[36]) ^ (inputs[126]);
    assign layer0_outputs[1959] = ~(inputs[233]);
    assign layer0_outputs[1960] = inputs[44];
    assign layer0_outputs[1961] = inputs[113];
    assign layer0_outputs[1962] = ~(inputs[90]);
    assign layer0_outputs[1963] = ~(inputs[234]) | (inputs[172]);
    assign layer0_outputs[1964] = (inputs[151]) & ~(inputs[3]);
    assign layer0_outputs[1965] = ~(inputs[247]);
    assign layer0_outputs[1966] = ~((inputs[222]) ^ (inputs[6]));
    assign layer0_outputs[1967] = (inputs[90]) | (inputs[60]);
    assign layer0_outputs[1968] = ~((inputs[6]) | (inputs[166]));
    assign layer0_outputs[1969] = (inputs[8]) ^ (inputs[112]);
    assign layer0_outputs[1970] = ~((inputs[62]) | (inputs[160]));
    assign layer0_outputs[1971] = ~(inputs[168]);
    assign layer0_outputs[1972] = inputs[229];
    assign layer0_outputs[1973] = ~((inputs[223]) ^ (inputs[13]));
    assign layer0_outputs[1974] = ~(inputs[232]);
    assign layer0_outputs[1975] = (inputs[73]) & ~(inputs[225]);
    assign layer0_outputs[1976] = (inputs[146]) ^ (inputs[242]);
    assign layer0_outputs[1977] = (inputs[218]) | (inputs[4]);
    assign layer0_outputs[1978] = inputs[181];
    assign layer0_outputs[1979] = ~(inputs[176]);
    assign layer0_outputs[1980] = (inputs[211]) & ~(inputs[105]);
    assign layer0_outputs[1981] = 1'b0;
    assign layer0_outputs[1982] = inputs[9];
    assign layer0_outputs[1983] = ~((inputs[90]) | (inputs[254]));
    assign layer0_outputs[1984] = ~((inputs[10]) | (inputs[224]));
    assign layer0_outputs[1985] = (inputs[159]) & ~(inputs[131]);
    assign layer0_outputs[1986] = (inputs[154]) | (inputs[140]);
    assign layer0_outputs[1987] = ~(inputs[203]);
    assign layer0_outputs[1988] = (inputs[247]) | (inputs[97]);
    assign layer0_outputs[1989] = ~(inputs[126]);
    assign layer0_outputs[1990] = (inputs[212]) | (inputs[205]);
    assign layer0_outputs[1991] = (inputs[159]) | (inputs[212]);
    assign layer0_outputs[1992] = ~(inputs[24]);
    assign layer0_outputs[1993] = inputs[22];
    assign layer0_outputs[1994] = ~((inputs[88]) ^ (inputs[139]));
    assign layer0_outputs[1995] = ~((inputs[250]) ^ (inputs[156]));
    assign layer0_outputs[1996] = ~((inputs[246]) | (inputs[173]));
    assign layer0_outputs[1997] = inputs[29];
    assign layer0_outputs[1998] = (inputs[177]) & ~(inputs[141]);
    assign layer0_outputs[1999] = (inputs[251]) ^ (inputs[173]);
    assign layer0_outputs[2000] = ~((inputs[96]) ^ (inputs[108]));
    assign layer0_outputs[2001] = ~(inputs[90]) | (inputs[222]);
    assign layer0_outputs[2002] = inputs[143];
    assign layer0_outputs[2003] = (inputs[126]) & ~(inputs[190]);
    assign layer0_outputs[2004] = (inputs[25]) & ~(inputs[162]);
    assign layer0_outputs[2005] = (inputs[192]) ^ (inputs[206]);
    assign layer0_outputs[2006] = ~(inputs[70]) | (inputs[18]);
    assign layer0_outputs[2007] = inputs[50];
    assign layer0_outputs[2008] = ~((inputs[137]) ^ (inputs[58]));
    assign layer0_outputs[2009] = (inputs[160]) ^ (inputs[115]);
    assign layer0_outputs[2010] = ~((inputs[7]) ^ (inputs[59]));
    assign layer0_outputs[2011] = ~((inputs[146]) | (inputs[148]));
    assign layer0_outputs[2012] = (inputs[49]) ^ (inputs[101]);
    assign layer0_outputs[2013] = inputs[208];
    assign layer0_outputs[2014] = (inputs[127]) & ~(inputs[95]);
    assign layer0_outputs[2015] = ~(inputs[156]);
    assign layer0_outputs[2016] = (inputs[225]) & ~(inputs[15]);
    assign layer0_outputs[2017] = (inputs[213]) & ~(inputs[174]);
    assign layer0_outputs[2018] = ~(inputs[8]) | (inputs[126]);
    assign layer0_outputs[2019] = ~(inputs[242]);
    assign layer0_outputs[2020] = ~(inputs[218]) | (inputs[75]);
    assign layer0_outputs[2021] = (inputs[240]) & (inputs[134]);
    assign layer0_outputs[2022] = (inputs[156]) | (inputs[9]);
    assign layer0_outputs[2023] = ~((inputs[140]) & (inputs[78]));
    assign layer0_outputs[2024] = (inputs[16]) | (inputs[2]);
    assign layer0_outputs[2025] = (inputs[74]) | (inputs[108]);
    assign layer0_outputs[2026] = (inputs[173]) & ~(inputs[95]);
    assign layer0_outputs[2027] = ~(inputs[136]) | (inputs[205]);
    assign layer0_outputs[2028] = ~((inputs[172]) ^ (inputs[184]));
    assign layer0_outputs[2029] = inputs[235];
    assign layer0_outputs[2030] = ~(inputs[244]);
    assign layer0_outputs[2031] = (inputs[243]) | (inputs[225]);
    assign layer0_outputs[2032] = (inputs[39]) | (inputs[116]);
    assign layer0_outputs[2033] = (inputs[101]) ^ (inputs[69]);
    assign layer0_outputs[2034] = ~(inputs[147]);
    assign layer0_outputs[2035] = (inputs[189]) & ~(inputs[95]);
    assign layer0_outputs[2036] = inputs[221];
    assign layer0_outputs[2037] = (inputs[234]) & ~(inputs[91]);
    assign layer0_outputs[2038] = (inputs[194]) & ~(inputs[223]);
    assign layer0_outputs[2039] = inputs[67];
    assign layer0_outputs[2040] = (inputs[183]) & ~(inputs[180]);
    assign layer0_outputs[2041] = ~((inputs[161]) | (inputs[75]));
    assign layer0_outputs[2042] = (inputs[85]) & ~(inputs[223]);
    assign layer0_outputs[2043] = inputs[62];
    assign layer0_outputs[2044] = (inputs[87]) ^ (inputs[125]);
    assign layer0_outputs[2045] = ~((inputs[236]) ^ (inputs[195]));
    assign layer0_outputs[2046] = ~(inputs[158]);
    assign layer0_outputs[2047] = (inputs[43]) | (inputs[97]);
    assign layer0_outputs[2048] = ~(inputs[122]);
    assign layer0_outputs[2049] = ~(inputs[145]);
    assign layer0_outputs[2050] = ~((inputs[130]) | (inputs[244]));
    assign layer0_outputs[2051] = ~(inputs[87]);
    assign layer0_outputs[2052] = ~((inputs[201]) ^ (inputs[221]));
    assign layer0_outputs[2053] = (inputs[143]) & ~(inputs[96]);
    assign layer0_outputs[2054] = (inputs[106]) & ~(inputs[20]);
    assign layer0_outputs[2055] = (inputs[7]) & ~(inputs[175]);
    assign layer0_outputs[2056] = inputs[59];
    assign layer0_outputs[2057] = (inputs[137]) | (inputs[104]);
    assign layer0_outputs[2058] = inputs[30];
    assign layer0_outputs[2059] = ~(inputs[36]) | (inputs[143]);
    assign layer0_outputs[2060] = (inputs[106]) & ~(inputs[204]);
    assign layer0_outputs[2061] = (inputs[91]) ^ (inputs[245]);
    assign layer0_outputs[2062] = ~(inputs[135]);
    assign layer0_outputs[2063] = inputs[150];
    assign layer0_outputs[2064] = ~(inputs[23]);
    assign layer0_outputs[2065] = (inputs[141]) | (inputs[57]);
    assign layer0_outputs[2066] = inputs[3];
    assign layer0_outputs[2067] = ~((inputs[168]) ^ (inputs[232]));
    assign layer0_outputs[2068] = ~(inputs[9]);
    assign layer0_outputs[2069] = inputs[122];
    assign layer0_outputs[2070] = ~((inputs[58]) | (inputs[176]));
    assign layer0_outputs[2071] = inputs[38];
    assign layer0_outputs[2072] = inputs[23];
    assign layer0_outputs[2073] = ~(inputs[147]);
    assign layer0_outputs[2074] = ~(inputs[68]);
    assign layer0_outputs[2075] = ~(inputs[180]) | (inputs[79]);
    assign layer0_outputs[2076] = inputs[247];
    assign layer0_outputs[2077] = inputs[109];
    assign layer0_outputs[2078] = ~(inputs[233]) | (inputs[86]);
    assign layer0_outputs[2079] = (inputs[158]) & ~(inputs[48]);
    assign layer0_outputs[2080] = (inputs[222]) | (inputs[31]);
    assign layer0_outputs[2081] = (inputs[132]) ^ (inputs[122]);
    assign layer0_outputs[2082] = ~(inputs[235]);
    assign layer0_outputs[2083] = (inputs[134]) & ~(inputs[17]);
    assign layer0_outputs[2084] = (inputs[66]) | (inputs[93]);
    assign layer0_outputs[2085] = inputs[225];
    assign layer0_outputs[2086] = ~(inputs[176]) | (inputs[95]);
    assign layer0_outputs[2087] = ~(inputs[137]);
    assign layer0_outputs[2088] = ~((inputs[17]) ^ (inputs[30]));
    assign layer0_outputs[2089] = inputs[20];
    assign layer0_outputs[2090] = ~(inputs[230]);
    assign layer0_outputs[2091] = (inputs[124]) | (inputs[68]);
    assign layer0_outputs[2092] = ~((inputs[206]) & (inputs[241]));
    assign layer0_outputs[2093] = ~((inputs[68]) ^ (inputs[195]));
    assign layer0_outputs[2094] = ~((inputs[14]) | (inputs[115]));
    assign layer0_outputs[2095] = ~(inputs[6]);
    assign layer0_outputs[2096] = (inputs[98]) ^ (inputs[218]);
    assign layer0_outputs[2097] = (inputs[101]) & ~(inputs[207]);
    assign layer0_outputs[2098] = (inputs[49]) | (inputs[93]);
    assign layer0_outputs[2099] = ~((inputs[124]) ^ (inputs[117]));
    assign layer0_outputs[2100] = ~(inputs[181]) | (inputs[240]);
    assign layer0_outputs[2101] = (inputs[147]) ^ (inputs[85]);
    assign layer0_outputs[2102] = inputs[118];
    assign layer0_outputs[2103] = ~(inputs[107]);
    assign layer0_outputs[2104] = (inputs[255]) | (inputs[204]);
    assign layer0_outputs[2105] = ~((inputs[155]) | (inputs[162]));
    assign layer0_outputs[2106] = (inputs[211]) | (inputs[71]);
    assign layer0_outputs[2107] = 1'b0;
    assign layer0_outputs[2108] = (inputs[15]) & (inputs[153]);
    assign layer0_outputs[2109] = ~((inputs[210]) | (inputs[41]));
    assign layer0_outputs[2110] = inputs[150];
    assign layer0_outputs[2111] = (inputs[189]) & ~(inputs[83]);
    assign layer0_outputs[2112] = (inputs[84]) & ~(inputs[42]);
    assign layer0_outputs[2113] = ~(inputs[7]);
    assign layer0_outputs[2114] = (inputs[63]) | (inputs[201]);
    assign layer0_outputs[2115] = ~(inputs[166]);
    assign layer0_outputs[2116] = ~((inputs[121]) ^ (inputs[162]));
    assign layer0_outputs[2117] = (inputs[197]) & ~(inputs[124]);
    assign layer0_outputs[2118] = inputs[147];
    assign layer0_outputs[2119] = ~(inputs[127]) | (inputs[152]);
    assign layer0_outputs[2120] = ~((inputs[159]) ^ (inputs[1]));
    assign layer0_outputs[2121] = inputs[101];
    assign layer0_outputs[2122] = (inputs[120]) & ~(inputs[76]);
    assign layer0_outputs[2123] = inputs[3];
    assign layer0_outputs[2124] = (inputs[165]) & ~(inputs[223]);
    assign layer0_outputs[2125] = ~(inputs[194]);
    assign layer0_outputs[2126] = ~(inputs[120]);
    assign layer0_outputs[2127] = ~(inputs[213]);
    assign layer0_outputs[2128] = ~(inputs[98]);
    assign layer0_outputs[2129] = ~(inputs[116]);
    assign layer0_outputs[2130] = ~(inputs[182]);
    assign layer0_outputs[2131] = ~((inputs[198]) | (inputs[3]));
    assign layer0_outputs[2132] = inputs[247];
    assign layer0_outputs[2133] = inputs[192];
    assign layer0_outputs[2134] = ~(inputs[114]) | (inputs[172]);
    assign layer0_outputs[2135] = (inputs[71]) & ~(inputs[150]);
    assign layer0_outputs[2136] = ~(inputs[229]);
    assign layer0_outputs[2137] = (inputs[233]) | (inputs[187]);
    assign layer0_outputs[2138] = ~((inputs[66]) | (inputs[184]));
    assign layer0_outputs[2139] = inputs[13];
    assign layer0_outputs[2140] = ~(inputs[231]);
    assign layer0_outputs[2141] = (inputs[67]) ^ (inputs[24]);
    assign layer0_outputs[2142] = (inputs[172]) & ~(inputs[64]);
    assign layer0_outputs[2143] = ~(inputs[92]) | (inputs[159]);
    assign layer0_outputs[2144] = inputs[210];
    assign layer0_outputs[2145] = ~(inputs[135]);
    assign layer0_outputs[2146] = ~((inputs[90]) ^ (inputs[206]));
    assign layer0_outputs[2147] = ~(inputs[105]);
    assign layer0_outputs[2148] = (inputs[151]) | (inputs[98]);
    assign layer0_outputs[2149] = ~((inputs[89]) | (inputs[148]));
    assign layer0_outputs[2150] = inputs[228];
    assign layer0_outputs[2151] = (inputs[250]) | (inputs[44]);
    assign layer0_outputs[2152] = (inputs[23]) & ~(inputs[196]);
    assign layer0_outputs[2153] = (inputs[86]) ^ (inputs[154]);
    assign layer0_outputs[2154] = ~(inputs[150]) | (inputs[14]);
    assign layer0_outputs[2155] = ~((inputs[76]) | (inputs[140]));
    assign layer0_outputs[2156] = ~((inputs[28]) | (inputs[96]));
    assign layer0_outputs[2157] = ~(inputs[167]);
    assign layer0_outputs[2158] = ~(inputs[119]);
    assign layer0_outputs[2159] = (inputs[96]) | (inputs[246]);
    assign layer0_outputs[2160] = inputs[139];
    assign layer0_outputs[2161] = inputs[233];
    assign layer0_outputs[2162] = ~(inputs[214]) | (inputs[162]);
    assign layer0_outputs[2163] = (inputs[153]) | (inputs[151]);
    assign layer0_outputs[2164] = (inputs[167]) & ~(inputs[255]);
    assign layer0_outputs[2165] = ~(inputs[59]);
    assign layer0_outputs[2166] = (inputs[123]) | (inputs[140]);
    assign layer0_outputs[2167] = ~(inputs[207]);
    assign layer0_outputs[2168] = (inputs[233]) & ~(inputs[62]);
    assign layer0_outputs[2169] = (inputs[216]) & ~(inputs[104]);
    assign layer0_outputs[2170] = ~((inputs[165]) | (inputs[166]));
    assign layer0_outputs[2171] = inputs[239];
    assign layer0_outputs[2172] = inputs[39];
    assign layer0_outputs[2173] = ~((inputs[53]) | (inputs[8]));
    assign layer0_outputs[2174] = (inputs[202]) | (inputs[11]);
    assign layer0_outputs[2175] = (inputs[26]) & ~(inputs[213]);
    assign layer0_outputs[2176] = ~(inputs[119]);
    assign layer0_outputs[2177] = 1'b0;
    assign layer0_outputs[2178] = inputs[190];
    assign layer0_outputs[2179] = (inputs[104]) & ~(inputs[155]);
    assign layer0_outputs[2180] = ~(inputs[101]) | (inputs[160]);
    assign layer0_outputs[2181] = ~(inputs[22]);
    assign layer0_outputs[2182] = ~(inputs[248]) | (inputs[77]);
    assign layer0_outputs[2183] = ~(inputs[44]);
    assign layer0_outputs[2184] = ~(inputs[221]);
    assign layer0_outputs[2185] = ~(inputs[216]) | (inputs[69]);
    assign layer0_outputs[2186] = inputs[232];
    assign layer0_outputs[2187] = ~(inputs[4]) | (inputs[218]);
    assign layer0_outputs[2188] = inputs[134];
    assign layer0_outputs[2189] = (inputs[166]) & ~(inputs[191]);
    assign layer0_outputs[2190] = (inputs[132]) ^ (inputs[102]);
    assign layer0_outputs[2191] = ~((inputs[215]) ^ (inputs[199]));
    assign layer0_outputs[2192] = ~((inputs[29]) ^ (inputs[132]));
    assign layer0_outputs[2193] = ~(inputs[71]) | (inputs[46]);
    assign layer0_outputs[2194] = ~(inputs[236]) | (inputs[81]);
    assign layer0_outputs[2195] = ~((inputs[39]) & (inputs[112]));
    assign layer0_outputs[2196] = (inputs[234]) & ~(inputs[123]);
    assign layer0_outputs[2197] = ~((inputs[117]) | (inputs[83]));
    assign layer0_outputs[2198] = (inputs[37]) & ~(inputs[124]);
    assign layer0_outputs[2199] = ~((inputs[175]) | (inputs[198]));
    assign layer0_outputs[2200] = (inputs[147]) | (inputs[163]);
    assign layer0_outputs[2201] = 1'b1;
    assign layer0_outputs[2202] = inputs[62];
    assign layer0_outputs[2203] = ~(inputs[254]);
    assign layer0_outputs[2204] = (inputs[30]) | (inputs[26]);
    assign layer0_outputs[2205] = ~(inputs[231]) | (inputs[63]);
    assign layer0_outputs[2206] = inputs[86];
    assign layer0_outputs[2207] = (inputs[119]) & ~(inputs[52]);
    assign layer0_outputs[2208] = inputs[230];
    assign layer0_outputs[2209] = ~(inputs[229]);
    assign layer0_outputs[2210] = inputs[144];
    assign layer0_outputs[2211] = ~((inputs[91]) ^ (inputs[108]));
    assign layer0_outputs[2212] = (inputs[90]) & ~(inputs[116]);
    assign layer0_outputs[2213] = ~(inputs[38]);
    assign layer0_outputs[2214] = ~((inputs[158]) | (inputs[129]));
    assign layer0_outputs[2215] = (inputs[40]) | (inputs[32]);
    assign layer0_outputs[2216] = (inputs[177]) & ~(inputs[48]);
    assign layer0_outputs[2217] = inputs[59];
    assign layer0_outputs[2218] = (inputs[180]) | (inputs[236]);
    assign layer0_outputs[2219] = (inputs[85]) & (inputs[225]);
    assign layer0_outputs[2220] = (inputs[198]) & ~(inputs[123]);
    assign layer0_outputs[2221] = 1'b1;
    assign layer0_outputs[2222] = inputs[25];
    assign layer0_outputs[2223] = ~((inputs[107]) | (inputs[33]));
    assign layer0_outputs[2224] = 1'b1;
    assign layer0_outputs[2225] = (inputs[148]) & ~(inputs[108]);
    assign layer0_outputs[2226] = inputs[188];
    assign layer0_outputs[2227] = (inputs[209]) & ~(inputs[15]);
    assign layer0_outputs[2228] = (inputs[169]) | (inputs[127]);
    assign layer0_outputs[2229] = (inputs[184]) | (inputs[82]);
    assign layer0_outputs[2230] = (inputs[136]) | (inputs[91]);
    assign layer0_outputs[2231] = ~(inputs[166]);
    assign layer0_outputs[2232] = (inputs[190]) | (inputs[198]);
    assign layer0_outputs[2233] = (inputs[68]) & ~(inputs[175]);
    assign layer0_outputs[2234] = ~(inputs[233]);
    assign layer0_outputs[2235] = (inputs[254]) | (inputs[151]);
    assign layer0_outputs[2236] = ~(inputs[248]) | (inputs[64]);
    assign layer0_outputs[2237] = ~(inputs[152]) | (inputs[27]);
    assign layer0_outputs[2238] = ~((inputs[139]) ^ (inputs[24]));
    assign layer0_outputs[2239] = ~(inputs[101]);
    assign layer0_outputs[2240] = ~(inputs[124]);
    assign layer0_outputs[2241] = (inputs[162]) & ~(inputs[56]);
    assign layer0_outputs[2242] = inputs[200];
    assign layer0_outputs[2243] = inputs[6];
    assign layer0_outputs[2244] = (inputs[219]) & ~(inputs[82]);
    assign layer0_outputs[2245] = (inputs[133]) & (inputs[246]);
    assign layer0_outputs[2246] = ~(inputs[85]);
    assign layer0_outputs[2247] = ~(inputs[162]);
    assign layer0_outputs[2248] = (inputs[77]) | (inputs[191]);
    assign layer0_outputs[2249] = inputs[103];
    assign layer0_outputs[2250] = ~((inputs[147]) ^ (inputs[177]));
    assign layer0_outputs[2251] = ~((inputs[189]) | (inputs[221]));
    assign layer0_outputs[2252] = ~((inputs[51]) | (inputs[114]));
    assign layer0_outputs[2253] = ~((inputs[100]) | (inputs[127]));
    assign layer0_outputs[2254] = ~(inputs[146]) | (inputs[186]);
    assign layer0_outputs[2255] = inputs[223];
    assign layer0_outputs[2256] = inputs[43];
    assign layer0_outputs[2257] = ~(inputs[233]) | (inputs[10]);
    assign layer0_outputs[2258] = (inputs[50]) & ~(inputs[81]);
    assign layer0_outputs[2259] = (inputs[48]) ^ (inputs[203]);
    assign layer0_outputs[2260] = (inputs[36]) | (inputs[132]);
    assign layer0_outputs[2261] = ~((inputs[79]) ^ (inputs[178]));
    assign layer0_outputs[2262] = 1'b0;
    assign layer0_outputs[2263] = (inputs[77]) & ~(inputs[2]);
    assign layer0_outputs[2264] = ~(inputs[188]) | (inputs[93]);
    assign layer0_outputs[2265] = (inputs[117]) ^ (inputs[69]);
    assign layer0_outputs[2266] = 1'b1;
    assign layer0_outputs[2267] = (inputs[157]) | (inputs[87]);
    assign layer0_outputs[2268] = (inputs[51]) & ~(inputs[132]);
    assign layer0_outputs[2269] = ~((inputs[157]) | (inputs[242]));
    assign layer0_outputs[2270] = ~(inputs[163]);
    assign layer0_outputs[2271] = inputs[198];
    assign layer0_outputs[2272] = ~((inputs[109]) ^ (inputs[181]));
    assign layer0_outputs[2273] = (inputs[238]) & ~(inputs[224]);
    assign layer0_outputs[2274] = ~((inputs[124]) | (inputs[148]));
    assign layer0_outputs[2275] = (inputs[87]) & ~(inputs[177]);
    assign layer0_outputs[2276] = ~(inputs[174]);
    assign layer0_outputs[2277] = inputs[238];
    assign layer0_outputs[2278] = ~((inputs[61]) ^ (inputs[23]));
    assign layer0_outputs[2279] = (inputs[111]) ^ (inputs[230]);
    assign layer0_outputs[2280] = ~(inputs[188]) | (inputs[12]);
    assign layer0_outputs[2281] = ~(inputs[101]) | (inputs[3]);
    assign layer0_outputs[2282] = ~((inputs[78]) | (inputs[191]));
    assign layer0_outputs[2283] = 1'b1;
    assign layer0_outputs[2284] = (inputs[5]) ^ (inputs[159]);
    assign layer0_outputs[2285] = (inputs[104]) & ~(inputs[164]);
    assign layer0_outputs[2286] = ~(inputs[102]);
    assign layer0_outputs[2287] = ~(inputs[218]) | (inputs[12]);
    assign layer0_outputs[2288] = inputs[77];
    assign layer0_outputs[2289] = (inputs[140]) ^ (inputs[164]);
    assign layer0_outputs[2290] = (inputs[88]) & ~(inputs[157]);
    assign layer0_outputs[2291] = (inputs[0]) & (inputs[34]);
    assign layer0_outputs[2292] = (inputs[157]) & ~(inputs[153]);
    assign layer0_outputs[2293] = ~(inputs[226]);
    assign layer0_outputs[2294] = (inputs[83]) ^ (inputs[169]);
    assign layer0_outputs[2295] = ~(inputs[72]) | (inputs[151]);
    assign layer0_outputs[2296] = 1'b1;
    assign layer0_outputs[2297] = ~(inputs[169]) | (inputs[12]);
    assign layer0_outputs[2298] = (inputs[139]) & ~(inputs[34]);
    assign layer0_outputs[2299] = 1'b0;
    assign layer0_outputs[2300] = ~(inputs[134]) | (inputs[108]);
    assign layer0_outputs[2301] = inputs[214];
    assign layer0_outputs[2302] = inputs[185];
    assign layer0_outputs[2303] = (inputs[122]) ^ (inputs[158]);
    assign layer0_outputs[2304] = ~((inputs[88]) | (inputs[252]));
    assign layer0_outputs[2305] = ~(inputs[231]);
    assign layer0_outputs[2306] = inputs[103];
    assign layer0_outputs[2307] = (inputs[246]) ^ (inputs[112]);
    assign layer0_outputs[2308] = ~((inputs[2]) | (inputs[32]));
    assign layer0_outputs[2309] = ~(inputs[0]);
    assign layer0_outputs[2310] = (inputs[155]) & ~(inputs[5]);
    assign layer0_outputs[2311] = (inputs[109]) & ~(inputs[115]);
    assign layer0_outputs[2312] = inputs[18];
    assign layer0_outputs[2313] = ~(inputs[48]);
    assign layer0_outputs[2314] = (inputs[181]) & ~(inputs[162]);
    assign layer0_outputs[2315] = ~(inputs[152]);
    assign layer0_outputs[2316] = (inputs[172]) | (inputs[251]);
    assign layer0_outputs[2317] = ~((inputs[147]) ^ (inputs[190]));
    assign layer0_outputs[2318] = inputs[232];
    assign layer0_outputs[2319] = ~((inputs[235]) | (inputs[37]));
    assign layer0_outputs[2320] = ~((inputs[144]) ^ (inputs[211]));
    assign layer0_outputs[2321] = ~((inputs[241]) | (inputs[249]));
    assign layer0_outputs[2322] = (inputs[100]) & ~(inputs[224]);
    assign layer0_outputs[2323] = inputs[217];
    assign layer0_outputs[2324] = 1'b1;
    assign layer0_outputs[2325] = ~((inputs[168]) | (inputs[1]));
    assign layer0_outputs[2326] = (inputs[1]) & (inputs[15]);
    assign layer0_outputs[2327] = ~((inputs[29]) | (inputs[15]));
    assign layer0_outputs[2328] = ~((inputs[99]) | (inputs[165]));
    assign layer0_outputs[2329] = inputs[180];
    assign layer0_outputs[2330] = ~(inputs[103]) | (inputs[179]);
    assign layer0_outputs[2331] = ~(inputs[108]);
    assign layer0_outputs[2332] = inputs[132];
    assign layer0_outputs[2333] = ~((inputs[192]) | (inputs[6]));
    assign layer0_outputs[2334] = ~(inputs[119]);
    assign layer0_outputs[2335] = (inputs[172]) ^ (inputs[221]);
    assign layer0_outputs[2336] = (inputs[113]) | (inputs[99]);
    assign layer0_outputs[2337] = ~(inputs[211]);
    assign layer0_outputs[2338] = ~(inputs[212]);
    assign layer0_outputs[2339] = (inputs[104]) & ~(inputs[206]);
    assign layer0_outputs[2340] = ~((inputs[235]) & (inputs[218]));
    assign layer0_outputs[2341] = ~((inputs[209]) | (inputs[5]));
    assign layer0_outputs[2342] = (inputs[154]) & ~(inputs[250]);
    assign layer0_outputs[2343] = (inputs[138]) ^ (inputs[13]);
    assign layer0_outputs[2344] = (inputs[196]) | (inputs[252]);
    assign layer0_outputs[2345] = ~(inputs[231]);
    assign layer0_outputs[2346] = (inputs[206]) & (inputs[183]);
    assign layer0_outputs[2347] = ~((inputs[157]) & (inputs[77]));
    assign layer0_outputs[2348] = (inputs[34]) ^ (inputs[168]);
    assign layer0_outputs[2349] = ~(inputs[197]);
    assign layer0_outputs[2350] = ~(inputs[184]);
    assign layer0_outputs[2351] = (inputs[138]) ^ (inputs[136]);
    assign layer0_outputs[2352] = ~((inputs[223]) | (inputs[41]));
    assign layer0_outputs[2353] = inputs[40];
    assign layer0_outputs[2354] = (inputs[135]) | (inputs[134]);
    assign layer0_outputs[2355] = (inputs[142]) & (inputs[236]);
    assign layer0_outputs[2356] = ~((inputs[70]) ^ (inputs[109]));
    assign layer0_outputs[2357] = (inputs[149]) & ~(inputs[80]);
    assign layer0_outputs[2358] = inputs[195];
    assign layer0_outputs[2359] = ~((inputs[161]) | (inputs[212]));
    assign layer0_outputs[2360] = (inputs[61]) ^ (inputs[23]);
    assign layer0_outputs[2361] = ~((inputs[249]) ^ (inputs[102]));
    assign layer0_outputs[2362] = ~(inputs[108]);
    assign layer0_outputs[2363] = ~(inputs[181]) | (inputs[171]);
    assign layer0_outputs[2364] = ~((inputs[156]) ^ (inputs[8]));
    assign layer0_outputs[2365] = inputs[57];
    assign layer0_outputs[2366] = ~((inputs[79]) | (inputs[23]));
    assign layer0_outputs[2367] = ~((inputs[59]) & (inputs[106]));
    assign layer0_outputs[2368] = ~(inputs[34]) | (inputs[77]);
    assign layer0_outputs[2369] = ~((inputs[189]) ^ (inputs[27]));
    assign layer0_outputs[2370] = inputs[34];
    assign layer0_outputs[2371] = ~((inputs[229]) | (inputs[33]));
    assign layer0_outputs[2372] = (inputs[100]) & ~(inputs[110]);
    assign layer0_outputs[2373] = (inputs[220]) | (inputs[212]);
    assign layer0_outputs[2374] = ~(inputs[210]);
    assign layer0_outputs[2375] = (inputs[29]) & ~(inputs[189]);
    assign layer0_outputs[2376] = inputs[149];
    assign layer0_outputs[2377] = inputs[27];
    assign layer0_outputs[2378] = ~(inputs[41]);
    assign layer0_outputs[2379] = (inputs[68]) & ~(inputs[17]);
    assign layer0_outputs[2380] = ~(inputs[93]) | (inputs[181]);
    assign layer0_outputs[2381] = ~(inputs[75]) | (inputs[255]);
    assign layer0_outputs[2382] = (inputs[102]) ^ (inputs[148]);
    assign layer0_outputs[2383] = ~(inputs[148]);
    assign layer0_outputs[2384] = ~(inputs[241]);
    assign layer0_outputs[2385] = (inputs[246]) | (inputs[249]);
    assign layer0_outputs[2386] = ~((inputs[63]) ^ (inputs[16]));
    assign layer0_outputs[2387] = ~(inputs[152]) | (inputs[216]);
    assign layer0_outputs[2388] = (inputs[218]) | (inputs[207]);
    assign layer0_outputs[2389] = ~((inputs[54]) & (inputs[37]));
    assign layer0_outputs[2390] = inputs[118];
    assign layer0_outputs[2391] = inputs[91];
    assign layer0_outputs[2392] = ~(inputs[253]);
    assign layer0_outputs[2393] = ~((inputs[32]) ^ (inputs[14]));
    assign layer0_outputs[2394] = inputs[128];
    assign layer0_outputs[2395] = ~(inputs[251]);
    assign layer0_outputs[2396] = ~(inputs[24]);
    assign layer0_outputs[2397] = ~(inputs[244]) | (inputs[4]);
    assign layer0_outputs[2398] = ~(inputs[99]);
    assign layer0_outputs[2399] = (inputs[160]) & ~(inputs[254]);
    assign layer0_outputs[2400] = inputs[219];
    assign layer0_outputs[2401] = ~((inputs[32]) & (inputs[240]));
    assign layer0_outputs[2402] = inputs[131];
    assign layer0_outputs[2403] = ~((inputs[216]) | (inputs[201]));
    assign layer0_outputs[2404] = (inputs[107]) & ~(inputs[255]);
    assign layer0_outputs[2405] = inputs[77];
    assign layer0_outputs[2406] = ~(inputs[106]);
    assign layer0_outputs[2407] = (inputs[46]) & (inputs[107]);
    assign layer0_outputs[2408] = ~(inputs[148]) | (inputs[34]);
    assign layer0_outputs[2409] = ~((inputs[82]) ^ (inputs[182]));
    assign layer0_outputs[2410] = ~(inputs[30]) | (inputs[206]);
    assign layer0_outputs[2411] = (inputs[44]) & (inputs[191]);
    assign layer0_outputs[2412] = inputs[210];
    assign layer0_outputs[2413] = ~(inputs[106]);
    assign layer0_outputs[2414] = ~(inputs[88]) | (inputs[143]);
    assign layer0_outputs[2415] = (inputs[232]) & (inputs[164]);
    assign layer0_outputs[2416] = ~((inputs[25]) | (inputs[189]));
    assign layer0_outputs[2417] = inputs[191];
    assign layer0_outputs[2418] = inputs[40];
    assign layer0_outputs[2419] = inputs[41];
    assign layer0_outputs[2420] = ~((inputs[232]) ^ (inputs[155]));
    assign layer0_outputs[2421] = ~(inputs[105]);
    assign layer0_outputs[2422] = ~(inputs[216]);
    assign layer0_outputs[2423] = (inputs[39]) & ~(inputs[157]);
    assign layer0_outputs[2424] = (inputs[85]) & (inputs[88]);
    assign layer0_outputs[2425] = (inputs[93]) | (inputs[126]);
    assign layer0_outputs[2426] = (inputs[212]) | (inputs[65]);
    assign layer0_outputs[2427] = (inputs[41]) ^ (inputs[80]);
    assign layer0_outputs[2428] = (inputs[51]) & ~(inputs[54]);
    assign layer0_outputs[2429] = ~((inputs[62]) ^ (inputs[228]));
    assign layer0_outputs[2430] = (inputs[205]) | (inputs[228]);
    assign layer0_outputs[2431] = ~(inputs[182]) | (inputs[71]);
    assign layer0_outputs[2432] = 1'b0;
    assign layer0_outputs[2433] = (inputs[74]) & (inputs[33]);
    assign layer0_outputs[2434] = inputs[239];
    assign layer0_outputs[2435] = (inputs[115]) ^ (inputs[129]);
    assign layer0_outputs[2436] = (inputs[77]) & ~(inputs[132]);
    assign layer0_outputs[2437] = ~(inputs[246]);
    assign layer0_outputs[2438] = inputs[19];
    assign layer0_outputs[2439] = 1'b1;
    assign layer0_outputs[2440] = inputs[103];
    assign layer0_outputs[2441] = (inputs[116]) & ~(inputs[178]);
    assign layer0_outputs[2442] = inputs[158];
    assign layer0_outputs[2443] = ~(inputs[115]) | (inputs[180]);
    assign layer0_outputs[2444] = (inputs[183]) ^ (inputs[54]);
    assign layer0_outputs[2445] = ~(inputs[96]);
    assign layer0_outputs[2446] = ~((inputs[175]) ^ (inputs[219]));
    assign layer0_outputs[2447] = inputs[85];
    assign layer0_outputs[2448] = (inputs[12]) | (inputs[34]);
    assign layer0_outputs[2449] = (inputs[160]) | (inputs[208]);
    assign layer0_outputs[2450] = (inputs[170]) | (inputs[144]);
    assign layer0_outputs[2451] = inputs[174];
    assign layer0_outputs[2452] = ~((inputs[252]) ^ (inputs[147]));
    assign layer0_outputs[2453] = (inputs[163]) | (inputs[93]);
    assign layer0_outputs[2454] = (inputs[96]) ^ (inputs[30]);
    assign layer0_outputs[2455] = (inputs[43]) ^ (inputs[28]);
    assign layer0_outputs[2456] = inputs[139];
    assign layer0_outputs[2457] = 1'b0;
    assign layer0_outputs[2458] = inputs[44];
    assign layer0_outputs[2459] = ~(inputs[167]);
    assign layer0_outputs[2460] = (inputs[156]) ^ (inputs[123]);
    assign layer0_outputs[2461] = ~(inputs[234]);
    assign layer0_outputs[2462] = (inputs[114]) ^ (inputs[149]);
    assign layer0_outputs[2463] = ~(inputs[104]);
    assign layer0_outputs[2464] = ~((inputs[189]) | (inputs[174]));
    assign layer0_outputs[2465] = (inputs[16]) & (inputs[239]);
    assign layer0_outputs[2466] = (inputs[245]) & ~(inputs[49]);
    assign layer0_outputs[2467] = ~(inputs[136]);
    assign layer0_outputs[2468] = ~(inputs[202]) | (inputs[70]);
    assign layer0_outputs[2469] = ~(inputs[153]) | (inputs[65]);
    assign layer0_outputs[2470] = ~(inputs[90]) | (inputs[61]);
    assign layer0_outputs[2471] = ~(inputs[73]) | (inputs[158]);
    assign layer0_outputs[2472] = ~(inputs[215]);
    assign layer0_outputs[2473] = ~(inputs[54]);
    assign layer0_outputs[2474] = inputs[68];
    assign layer0_outputs[2475] = ~(inputs[193]);
    assign layer0_outputs[2476] = (inputs[104]) | (inputs[130]);
    assign layer0_outputs[2477] = inputs[36];
    assign layer0_outputs[2478] = (inputs[123]) & ~(inputs[182]);
    assign layer0_outputs[2479] = ~(inputs[186]) | (inputs[33]);
    assign layer0_outputs[2480] = ~(inputs[252]) | (inputs[205]);
    assign layer0_outputs[2481] = ~(inputs[172]);
    assign layer0_outputs[2482] = inputs[215];
    assign layer0_outputs[2483] = (inputs[219]) ^ (inputs[155]);
    assign layer0_outputs[2484] = ~((inputs[123]) & (inputs[249]));
    assign layer0_outputs[2485] = (inputs[89]) ^ (inputs[75]);
    assign layer0_outputs[2486] = ~((inputs[221]) | (inputs[239]));
    assign layer0_outputs[2487] = (inputs[181]) & ~(inputs[130]);
    assign layer0_outputs[2488] = (inputs[237]) ^ (inputs[116]);
    assign layer0_outputs[2489] = inputs[90];
    assign layer0_outputs[2490] = (inputs[47]) | (inputs[61]);
    assign layer0_outputs[2491] = ~(inputs[40]);
    assign layer0_outputs[2492] = (inputs[106]) & (inputs[10]);
    assign layer0_outputs[2493] = ~((inputs[99]) | (inputs[95]));
    assign layer0_outputs[2494] = (inputs[79]) | (inputs[191]);
    assign layer0_outputs[2495] = 1'b1;
    assign layer0_outputs[2496] = (inputs[61]) ^ (inputs[243]);
    assign layer0_outputs[2497] = inputs[73];
    assign layer0_outputs[2498] = (inputs[159]) | (inputs[112]);
    assign layer0_outputs[2499] = ~((inputs[48]) | (inputs[194]));
    assign layer0_outputs[2500] = (inputs[177]) | (inputs[204]);
    assign layer0_outputs[2501] = (inputs[176]) & (inputs[64]);
    assign layer0_outputs[2502] = ~(inputs[116]);
    assign layer0_outputs[2503] = ~((inputs[253]) | (inputs[153]));
    assign layer0_outputs[2504] = 1'b1;
    assign layer0_outputs[2505] = inputs[230];
    assign layer0_outputs[2506] = inputs[239];
    assign layer0_outputs[2507] = ~((inputs[218]) | (inputs[221]));
    assign layer0_outputs[2508] = ~(inputs[66]) | (inputs[172]);
    assign layer0_outputs[2509] = inputs[213];
    assign layer0_outputs[2510] = ~((inputs[11]) | (inputs[26]));
    assign layer0_outputs[2511] = inputs[6];
    assign layer0_outputs[2512] = ~((inputs[217]) ^ (inputs[201]));
    assign layer0_outputs[2513] = (inputs[92]) & ~(inputs[226]);
    assign layer0_outputs[2514] = ~((inputs[157]) ^ (inputs[101]));
    assign layer0_outputs[2515] = ~((inputs[88]) | (inputs[105]));
    assign layer0_outputs[2516] = ~((inputs[220]) | (inputs[231]));
    assign layer0_outputs[2517] = ~(inputs[77]) | (inputs[199]);
    assign layer0_outputs[2518] = ~((inputs[247]) | (inputs[65]));
    assign layer0_outputs[2519] = (inputs[171]) | (inputs[223]);
    assign layer0_outputs[2520] = (inputs[149]) | (inputs[18]);
    assign layer0_outputs[2521] = ~((inputs[111]) ^ (inputs[207]));
    assign layer0_outputs[2522] = inputs[249];
    assign layer0_outputs[2523] = (inputs[43]) | (inputs[164]);
    assign layer0_outputs[2524] = (inputs[121]) & ~(inputs[223]);
    assign layer0_outputs[2525] = ~(inputs[9]);
    assign layer0_outputs[2526] = ~(inputs[188]) | (inputs[107]);
    assign layer0_outputs[2527] = ~((inputs[35]) | (inputs[20]));
    assign layer0_outputs[2528] = ~(inputs[12]);
    assign layer0_outputs[2529] = ~(inputs[96]);
    assign layer0_outputs[2530] = 1'b0;
    assign layer0_outputs[2531] = ~(inputs[214]) | (inputs[21]);
    assign layer0_outputs[2532] = inputs[170];
    assign layer0_outputs[2533] = ~(inputs[92]) | (inputs[215]);
    assign layer0_outputs[2534] = ~(inputs[169]) | (inputs[17]);
    assign layer0_outputs[2535] = (inputs[41]) & (inputs[43]);
    assign layer0_outputs[2536] = (inputs[216]) & ~(inputs[54]);
    assign layer0_outputs[2537] = 1'b0;
    assign layer0_outputs[2538] = ~(inputs[35]) | (inputs[112]);
    assign layer0_outputs[2539] = (inputs[252]) | (inputs[138]);
    assign layer0_outputs[2540] = inputs[215];
    assign layer0_outputs[2541] = ~((inputs[31]) | (inputs[154]));
    assign layer0_outputs[2542] = ~(inputs[63]);
    assign layer0_outputs[2543] = (inputs[210]) & ~(inputs[31]);
    assign layer0_outputs[2544] = ~(inputs[20]) | (inputs[176]);
    assign layer0_outputs[2545] = (inputs[131]) & (inputs[39]);
    assign layer0_outputs[2546] = (inputs[108]) | (inputs[100]);
    assign layer0_outputs[2547] = ~(inputs[123]);
    assign layer0_outputs[2548] = inputs[36];
    assign layer0_outputs[2549] = ~((inputs[130]) | (inputs[190]));
    assign layer0_outputs[2550] = (inputs[97]) ^ (inputs[193]);
    assign layer0_outputs[2551] = (inputs[59]) & ~(inputs[59]);
    assign layer0_outputs[2552] = ~((inputs[76]) | (inputs[173]));
    assign layer0_outputs[2553] = ~(inputs[29]);
    assign layer0_outputs[2554] = ~((inputs[97]) | (inputs[228]));
    assign layer0_outputs[2555] = ~((inputs[15]) & (inputs[238]));
    assign layer0_outputs[2556] = ~(inputs[230]) | (inputs[123]);
    assign layer0_outputs[2557] = inputs[77];
    assign layer0_outputs[2558] = 1'b1;
    assign layer0_outputs[2559] = (inputs[156]) | (inputs[127]);
    assign layer0_outputs[2560] = (inputs[205]) | (inputs[95]);
    assign layer0_outputs[2561] = 1'b1;
    assign layer0_outputs[2562] = inputs[7];
    assign layer0_outputs[2563] = (inputs[207]) | (inputs[136]);
    assign layer0_outputs[2564] = ~(inputs[61]) | (inputs[0]);
    assign layer0_outputs[2565] = ~((inputs[81]) | (inputs[62]));
    assign layer0_outputs[2566] = ~((inputs[194]) ^ (inputs[24]));
    assign layer0_outputs[2567] = (inputs[70]) & ~(inputs[205]);
    assign layer0_outputs[2568] = inputs[38];
    assign layer0_outputs[2569] = (inputs[60]) | (inputs[40]);
    assign layer0_outputs[2570] = (inputs[5]) ^ (inputs[64]);
    assign layer0_outputs[2571] = (inputs[48]) ^ (inputs[103]);
    assign layer0_outputs[2572] = inputs[142];
    assign layer0_outputs[2573] = ~(inputs[23]);
    assign layer0_outputs[2574] = ~(inputs[109]);
    assign layer0_outputs[2575] = inputs[18];
    assign layer0_outputs[2576] = ~(inputs[153]);
    assign layer0_outputs[2577] = inputs[51];
    assign layer0_outputs[2578] = inputs[99];
    assign layer0_outputs[2579] = ~((inputs[245]) | (inputs[221]));
    assign layer0_outputs[2580] = ~((inputs[41]) | (inputs[225]));
    assign layer0_outputs[2581] = ~(inputs[137]) | (inputs[198]);
    assign layer0_outputs[2582] = ~((inputs[142]) ^ (inputs[162]));
    assign layer0_outputs[2583] = ~(inputs[16]);
    assign layer0_outputs[2584] = (inputs[253]) & ~(inputs[31]);
    assign layer0_outputs[2585] = ~(inputs[247]);
    assign layer0_outputs[2586] = ~((inputs[39]) ^ (inputs[223]));
    assign layer0_outputs[2587] = (inputs[235]) ^ (inputs[211]);
    assign layer0_outputs[2588] = ~(inputs[74]);
    assign layer0_outputs[2589] = (inputs[105]) ^ (inputs[163]);
    assign layer0_outputs[2590] = ~(inputs[38]) | (inputs[114]);
    assign layer0_outputs[2591] = (inputs[78]) ^ (inputs[171]);
    assign layer0_outputs[2592] = inputs[153];
    assign layer0_outputs[2593] = (inputs[67]) | (inputs[209]);
    assign layer0_outputs[2594] = ~((inputs[131]) | (inputs[198]));
    assign layer0_outputs[2595] = (inputs[218]) ^ (inputs[182]);
    assign layer0_outputs[2596] = (inputs[157]) ^ (inputs[124]);
    assign layer0_outputs[2597] = ~(inputs[30]) | (inputs[93]);
    assign layer0_outputs[2598] = inputs[197];
    assign layer0_outputs[2599] = ~(inputs[193]);
    assign layer0_outputs[2600] = ~((inputs[3]) | (inputs[125]));
    assign layer0_outputs[2601] = ~(inputs[109]);
    assign layer0_outputs[2602] = (inputs[151]) | (inputs[81]);
    assign layer0_outputs[2603] = ~(inputs[146]);
    assign layer0_outputs[2604] = (inputs[199]) & ~(inputs[10]);
    assign layer0_outputs[2605] = ~((inputs[148]) ^ (inputs[54]));
    assign layer0_outputs[2606] = ~((inputs[96]) ^ (inputs[54]));
    assign layer0_outputs[2607] = ~((inputs[200]) | (inputs[3]));
    assign layer0_outputs[2608] = inputs[179];
    assign layer0_outputs[2609] = ~(inputs[73]);
    assign layer0_outputs[2610] = (inputs[148]) ^ (inputs[195]);
    assign layer0_outputs[2611] = ~((inputs[169]) & (inputs[210]));
    assign layer0_outputs[2612] = (inputs[158]) ^ (inputs[159]);
    assign layer0_outputs[2613] = ~((inputs[195]) | (inputs[76]));
    assign layer0_outputs[2614] = ~(inputs[87]);
    assign layer0_outputs[2615] = (inputs[241]) | (inputs[227]);
    assign layer0_outputs[2616] = (inputs[27]) | (inputs[202]);
    assign layer0_outputs[2617] = ~((inputs[247]) | (inputs[250]));
    assign layer0_outputs[2618] = ~((inputs[231]) ^ (inputs[42]));
    assign layer0_outputs[2619] = ~(inputs[83]) | (inputs[191]);
    assign layer0_outputs[2620] = (inputs[160]) ^ (inputs[37]);
    assign layer0_outputs[2621] = (inputs[15]) | (inputs[52]);
    assign layer0_outputs[2622] = ~(inputs[214]);
    assign layer0_outputs[2623] = inputs[114];
    assign layer0_outputs[2624] = ~(inputs[9]);
    assign layer0_outputs[2625] = ~(inputs[17]) | (inputs[75]);
    assign layer0_outputs[2626] = ~(inputs[238]);
    assign layer0_outputs[2627] = ~(inputs[210]) | (inputs[133]);
    assign layer0_outputs[2628] = (inputs[233]) | (inputs[2]);
    assign layer0_outputs[2629] = ~(inputs[141]) | (inputs[110]);
    assign layer0_outputs[2630] = (inputs[62]) | (inputs[206]);
    assign layer0_outputs[2631] = (inputs[156]) & ~(inputs[225]);
    assign layer0_outputs[2632] = (inputs[160]) | (inputs[251]);
    assign layer0_outputs[2633] = ~((inputs[181]) | (inputs[14]));
    assign layer0_outputs[2634] = (inputs[47]) & ~(inputs[235]);
    assign layer0_outputs[2635] = inputs[182];
    assign layer0_outputs[2636] = ~(inputs[169]);
    assign layer0_outputs[2637] = ~(inputs[132]) | (inputs[226]);
    assign layer0_outputs[2638] = ~(inputs[195]);
    assign layer0_outputs[2639] = (inputs[251]) ^ (inputs[165]);
    assign layer0_outputs[2640] = ~((inputs[96]) | (inputs[49]));
    assign layer0_outputs[2641] = ~(inputs[154]);
    assign layer0_outputs[2642] = (inputs[214]) ^ (inputs[172]);
    assign layer0_outputs[2643] = ~((inputs[200]) | (inputs[141]));
    assign layer0_outputs[2644] = (inputs[6]) ^ (inputs[42]);
    assign layer0_outputs[2645] = inputs[173];
    assign layer0_outputs[2646] = ~((inputs[192]) | (inputs[144]));
    assign layer0_outputs[2647] = inputs[3];
    assign layer0_outputs[2648] = (inputs[188]) ^ (inputs[21]);
    assign layer0_outputs[2649] = ~(inputs[12]);
    assign layer0_outputs[2650] = ~((inputs[244]) | (inputs[103]));
    assign layer0_outputs[2651] = (inputs[51]) ^ (inputs[192]);
    assign layer0_outputs[2652] = (inputs[200]) | (inputs[151]);
    assign layer0_outputs[2653] = ~(inputs[167]);
    assign layer0_outputs[2654] = inputs[33];
    assign layer0_outputs[2655] = ~(inputs[120]) | (inputs[219]);
    assign layer0_outputs[2656] = ~(inputs[109]) | (inputs[115]);
    assign layer0_outputs[2657] = ~((inputs[234]) & (inputs[37]));
    assign layer0_outputs[2658] = (inputs[161]) & ~(inputs[223]);
    assign layer0_outputs[2659] = inputs[101];
    assign layer0_outputs[2660] = ~((inputs[196]) | (inputs[10]));
    assign layer0_outputs[2661] = (inputs[173]) & ~(inputs[76]);
    assign layer0_outputs[2662] = (inputs[101]) & ~(inputs[124]);
    assign layer0_outputs[2663] = (inputs[139]) & (inputs[157]);
    assign layer0_outputs[2664] = (inputs[193]) | (inputs[35]);
    assign layer0_outputs[2665] = (inputs[35]) & (inputs[217]);
    assign layer0_outputs[2666] = ~((inputs[121]) | (inputs[93]));
    assign layer0_outputs[2667] = inputs[59];
    assign layer0_outputs[2668] = ~(inputs[163]) | (inputs[160]);
    assign layer0_outputs[2669] = inputs[122];
    assign layer0_outputs[2670] = ~(inputs[248]);
    assign layer0_outputs[2671] = ~(inputs[197]);
    assign layer0_outputs[2672] = (inputs[3]) ^ (inputs[119]);
    assign layer0_outputs[2673] = ~((inputs[20]) ^ (inputs[140]));
    assign layer0_outputs[2674] = (inputs[245]) | (inputs[19]);
    assign layer0_outputs[2675] = ~((inputs[175]) | (inputs[201]));
    assign layer0_outputs[2676] = ~((inputs[145]) ^ (inputs[173]));
    assign layer0_outputs[2677] = (inputs[123]) ^ (inputs[38]);
    assign layer0_outputs[2678] = ~(inputs[85]);
    assign layer0_outputs[2679] = ~((inputs[152]) ^ (inputs[164]));
    assign layer0_outputs[2680] = ~((inputs[251]) | (inputs[106]));
    assign layer0_outputs[2681] = ~((inputs[211]) | (inputs[212]));
    assign layer0_outputs[2682] = inputs[21];
    assign layer0_outputs[2683] = ~((inputs[156]) | (inputs[126]));
    assign layer0_outputs[2684] = ~(inputs[59]) | (inputs[159]);
    assign layer0_outputs[2685] = ~(inputs[118]);
    assign layer0_outputs[2686] = (inputs[70]) ^ (inputs[64]);
    assign layer0_outputs[2687] = (inputs[173]) & ~(inputs[45]);
    assign layer0_outputs[2688] = ~(inputs[109]);
    assign layer0_outputs[2689] = (inputs[166]) ^ (inputs[146]);
    assign layer0_outputs[2690] = (inputs[220]) & ~(inputs[100]);
    assign layer0_outputs[2691] = ~(inputs[9]) | (inputs[24]);
    assign layer0_outputs[2692] = ~(inputs[23]) | (inputs[11]);
    assign layer0_outputs[2693] = ~(inputs[18]);
    assign layer0_outputs[2694] = ~((inputs[87]) ^ (inputs[69]));
    assign layer0_outputs[2695] = (inputs[247]) & ~(inputs[47]);
    assign layer0_outputs[2696] = ~((inputs[204]) | (inputs[175]));
    assign layer0_outputs[2697] = inputs[154];
    assign layer0_outputs[2698] = ~(inputs[202]) | (inputs[44]);
    assign layer0_outputs[2699] = (inputs[62]) & ~(inputs[105]);
    assign layer0_outputs[2700] = inputs[164];
    assign layer0_outputs[2701] = inputs[24];
    assign layer0_outputs[2702] = ~((inputs[196]) | (inputs[235]));
    assign layer0_outputs[2703] = ~((inputs[38]) | (inputs[169]));
    assign layer0_outputs[2704] = ~(inputs[184]) | (inputs[250]);
    assign layer0_outputs[2705] = ~(inputs[209]) | (inputs[140]);
    assign layer0_outputs[2706] = inputs[104];
    assign layer0_outputs[2707] = ~(inputs[230]);
    assign layer0_outputs[2708] = ~((inputs[161]) ^ (inputs[177]));
    assign layer0_outputs[2709] = ~(inputs[61]) | (inputs[124]);
    assign layer0_outputs[2710] = (inputs[119]) & ~(inputs[142]);
    assign layer0_outputs[2711] = ~(inputs[2]) | (inputs[66]);
    assign layer0_outputs[2712] = (inputs[102]) | (inputs[202]);
    assign layer0_outputs[2713] = ~(inputs[122]) | (inputs[225]);
    assign layer0_outputs[2714] = (inputs[205]) & ~(inputs[222]);
    assign layer0_outputs[2715] = (inputs[20]) ^ (inputs[48]);
    assign layer0_outputs[2716] = (inputs[211]) | (inputs[208]);
    assign layer0_outputs[2717] = (inputs[166]) | (inputs[121]);
    assign layer0_outputs[2718] = ~((inputs[200]) | (inputs[199]));
    assign layer0_outputs[2719] = inputs[6];
    assign layer0_outputs[2720] = ~(inputs[80]) | (inputs[157]);
    assign layer0_outputs[2721] = ~((inputs[169]) | (inputs[216]));
    assign layer0_outputs[2722] = inputs[21];
    assign layer0_outputs[2723] = inputs[58];
    assign layer0_outputs[2724] = inputs[98];
    assign layer0_outputs[2725] = ~(inputs[121]);
    assign layer0_outputs[2726] = ~((inputs[89]) ^ (inputs[18]));
    assign layer0_outputs[2727] = 1'b0;
    assign layer0_outputs[2728] = inputs[72];
    assign layer0_outputs[2729] = (inputs[35]) | (inputs[157]);
    assign layer0_outputs[2730] = ~(inputs[82]) | (inputs[224]);
    assign layer0_outputs[2731] = ~((inputs[85]) | (inputs[66]));
    assign layer0_outputs[2732] = (inputs[112]) | (inputs[21]);
    assign layer0_outputs[2733] = ~(inputs[63]);
    assign layer0_outputs[2734] = inputs[103];
    assign layer0_outputs[2735] = (inputs[202]) & ~(inputs[91]);
    assign layer0_outputs[2736] = ~((inputs[181]) ^ (inputs[211]));
    assign layer0_outputs[2737] = ~(inputs[158]);
    assign layer0_outputs[2738] = ~(inputs[118]) | (inputs[6]);
    assign layer0_outputs[2739] = ~(inputs[251]);
    assign layer0_outputs[2740] = (inputs[230]) & ~(inputs[165]);
    assign layer0_outputs[2741] = ~(inputs[72]);
    assign layer0_outputs[2742] = (inputs[250]) | (inputs[6]);
    assign layer0_outputs[2743] = ~((inputs[186]) ^ (inputs[101]));
    assign layer0_outputs[2744] = ~(inputs[23]) | (inputs[129]);
    assign layer0_outputs[2745] = (inputs[214]) | (inputs[129]);
    assign layer0_outputs[2746] = (inputs[103]) & ~(inputs[108]);
    assign layer0_outputs[2747] = (inputs[115]) ^ (inputs[103]);
    assign layer0_outputs[2748] = ~(inputs[144]);
    assign layer0_outputs[2749] = ~(inputs[132]);
    assign layer0_outputs[2750] = (inputs[35]) & ~(inputs[58]);
    assign layer0_outputs[2751] = (inputs[183]) & ~(inputs[99]);
    assign layer0_outputs[2752] = (inputs[42]) & ~(inputs[16]);
    assign layer0_outputs[2753] = ~(inputs[158]) | (inputs[146]);
    assign layer0_outputs[2754] = ~((inputs[0]) | (inputs[133]));
    assign layer0_outputs[2755] = (inputs[46]) ^ (inputs[18]);
    assign layer0_outputs[2756] = ~(inputs[187]);
    assign layer0_outputs[2757] = ~((inputs[206]) | (inputs[243]));
    assign layer0_outputs[2758] = (inputs[29]) | (inputs[218]);
    assign layer0_outputs[2759] = ~((inputs[148]) ^ (inputs[103]));
    assign layer0_outputs[2760] = ~(inputs[238]);
    assign layer0_outputs[2761] = inputs[164];
    assign layer0_outputs[2762] = inputs[23];
    assign layer0_outputs[2763] = ~((inputs[253]) | (inputs[147]));
    assign layer0_outputs[2764] = ~(inputs[106]);
    assign layer0_outputs[2765] = ~(inputs[235]) | (inputs[93]);
    assign layer0_outputs[2766] = ~((inputs[123]) ^ (inputs[172]));
    assign layer0_outputs[2767] = ~((inputs[202]) ^ (inputs[65]));
    assign layer0_outputs[2768] = (inputs[204]) | (inputs[101]);
    assign layer0_outputs[2769] = (inputs[189]) | (inputs[2]);
    assign layer0_outputs[2770] = (inputs[173]) ^ (inputs[158]);
    assign layer0_outputs[2771] = ~(inputs[7]);
    assign layer0_outputs[2772] = (inputs[238]) & ~(inputs[207]);
    assign layer0_outputs[2773] = (inputs[190]) ^ (inputs[63]);
    assign layer0_outputs[2774] = (inputs[187]) | (inputs[18]);
    assign layer0_outputs[2775] = (inputs[118]) | (inputs[98]);
    assign layer0_outputs[2776] = ~(inputs[53]) | (inputs[102]);
    assign layer0_outputs[2777] = ~(inputs[98]);
    assign layer0_outputs[2778] = (inputs[100]) ^ (inputs[196]);
    assign layer0_outputs[2779] = ~((inputs[209]) ^ (inputs[204]));
    assign layer0_outputs[2780] = ~((inputs[192]) ^ (inputs[204]));
    assign layer0_outputs[2781] = (inputs[31]) | (inputs[18]);
    assign layer0_outputs[2782] = ~(inputs[80]);
    assign layer0_outputs[2783] = (inputs[243]) & ~(inputs[254]);
    assign layer0_outputs[2784] = ~((inputs[213]) ^ (inputs[167]));
    assign layer0_outputs[2785] = inputs[169];
    assign layer0_outputs[2786] = inputs[139];
    assign layer0_outputs[2787] = ~(inputs[115]);
    assign layer0_outputs[2788] = inputs[132];
    assign layer0_outputs[2789] = inputs[219];
    assign layer0_outputs[2790] = ~((inputs[228]) | (inputs[181]));
    assign layer0_outputs[2791] = (inputs[144]) | (inputs[247]);
    assign layer0_outputs[2792] = ~((inputs[58]) & (inputs[71]));
    assign layer0_outputs[2793] = ~((inputs[179]) ^ (inputs[177]));
    assign layer0_outputs[2794] = (inputs[141]) | (inputs[124]);
    assign layer0_outputs[2795] = (inputs[249]) ^ (inputs[71]);
    assign layer0_outputs[2796] = ~((inputs[229]) ^ (inputs[197]));
    assign layer0_outputs[2797] = ~((inputs[47]) | (inputs[219]));
    assign layer0_outputs[2798] = inputs[198];
    assign layer0_outputs[2799] = ~(inputs[100]);
    assign layer0_outputs[2800] = ~((inputs[224]) & (inputs[42]));
    assign layer0_outputs[2801] = ~(inputs[23]) | (inputs[91]);
    assign layer0_outputs[2802] = ~((inputs[26]) | (inputs[67]));
    assign layer0_outputs[2803] = ~(inputs[227]) | (inputs[76]);
    assign layer0_outputs[2804] = ~(inputs[167]) | (inputs[78]);
    assign layer0_outputs[2805] = (inputs[184]) & ~(inputs[103]);
    assign layer0_outputs[2806] = ~(inputs[227]);
    assign layer0_outputs[2807] = (inputs[95]) | (inputs[11]);
    assign layer0_outputs[2808] = inputs[190];
    assign layer0_outputs[2809] = ~(inputs[194]) | (inputs[125]);
    assign layer0_outputs[2810] = ~(inputs[214]) | (inputs[46]);
    assign layer0_outputs[2811] = (inputs[175]) & ~(inputs[1]);
    assign layer0_outputs[2812] = (inputs[16]) | (inputs[255]);
    assign layer0_outputs[2813] = (inputs[151]) & ~(inputs[125]);
    assign layer0_outputs[2814] = (inputs[206]) & ~(inputs[250]);
    assign layer0_outputs[2815] = ~((inputs[212]) ^ (inputs[211]));
    assign layer0_outputs[2816] = ~(inputs[45]);
    assign layer0_outputs[2817] = inputs[58];
    assign layer0_outputs[2818] = ~(inputs[200]);
    assign layer0_outputs[2819] = ~(inputs[51]);
    assign layer0_outputs[2820] = ~(inputs[181]);
    assign layer0_outputs[2821] = ~(inputs[99]) | (inputs[122]);
    assign layer0_outputs[2822] = inputs[60];
    assign layer0_outputs[2823] = ~((inputs[185]) | (inputs[251]));
    assign layer0_outputs[2824] = 1'b0;
    assign layer0_outputs[2825] = (inputs[197]) & ~(inputs[208]);
    assign layer0_outputs[2826] = ~(inputs[45]);
    assign layer0_outputs[2827] = (inputs[198]) ^ (inputs[185]);
    assign layer0_outputs[2828] = ~(inputs[74]);
    assign layer0_outputs[2829] = inputs[37];
    assign layer0_outputs[2830] = ~(inputs[82]);
    assign layer0_outputs[2831] = inputs[43];
    assign layer0_outputs[2832] = ~((inputs[6]) | (inputs[229]));
    assign layer0_outputs[2833] = inputs[74];
    assign layer0_outputs[2834] = ~(inputs[125]) | (inputs[222]);
    assign layer0_outputs[2835] = inputs[111];
    assign layer0_outputs[2836] = ~((inputs[159]) | (inputs[12]));
    assign layer0_outputs[2837] = ~((inputs[5]) ^ (inputs[210]));
    assign layer0_outputs[2838] = ~(inputs[231]) | (inputs[129]);
    assign layer0_outputs[2839] = (inputs[24]) & ~(inputs[237]);
    assign layer0_outputs[2840] = inputs[23];
    assign layer0_outputs[2841] = inputs[57];
    assign layer0_outputs[2842] = (inputs[190]) ^ (inputs[9]);
    assign layer0_outputs[2843] = ~((inputs[80]) | (inputs[128]));
    assign layer0_outputs[2844] = inputs[9];
    assign layer0_outputs[2845] = (inputs[144]) & (inputs[82]);
    assign layer0_outputs[2846] = (inputs[193]) | (inputs[33]);
    assign layer0_outputs[2847] = (inputs[159]) | (inputs[148]);
    assign layer0_outputs[2848] = ~(inputs[118]) | (inputs[95]);
    assign layer0_outputs[2849] = inputs[160];
    assign layer0_outputs[2850] = (inputs[63]) | (inputs[46]);
    assign layer0_outputs[2851] = (inputs[30]) & ~(inputs[110]);
    assign layer0_outputs[2852] = inputs[105];
    assign layer0_outputs[2853] = ~((inputs[129]) | (inputs[219]));
    assign layer0_outputs[2854] = inputs[58];
    assign layer0_outputs[2855] = ~((inputs[100]) ^ (inputs[70]));
    assign layer0_outputs[2856] = ~(inputs[235]) | (inputs[5]);
    assign layer0_outputs[2857] = ~(inputs[180]) | (inputs[112]);
    assign layer0_outputs[2858] = inputs[67];
    assign layer0_outputs[2859] = ~((inputs[217]) & (inputs[182]));
    assign layer0_outputs[2860] = (inputs[246]) | (inputs[148]);
    assign layer0_outputs[2861] = ~((inputs[201]) | (inputs[251]));
    assign layer0_outputs[2862] = (inputs[250]) | (inputs[69]);
    assign layer0_outputs[2863] = (inputs[188]) & ~(inputs[27]);
    assign layer0_outputs[2864] = ~(inputs[151]);
    assign layer0_outputs[2865] = ~(inputs[195]);
    assign layer0_outputs[2866] = (inputs[196]) ^ (inputs[167]);
    assign layer0_outputs[2867] = ~(inputs[65]) | (inputs[252]);
    assign layer0_outputs[2868] = ~(inputs[109]);
    assign layer0_outputs[2869] = ~(inputs[8]) | (inputs[230]);
    assign layer0_outputs[2870] = ~((inputs[151]) | (inputs[1]));
    assign layer0_outputs[2871] = (inputs[25]) & ~(inputs[14]);
    assign layer0_outputs[2872] = ~((inputs[247]) ^ (inputs[175]));
    assign layer0_outputs[2873] = (inputs[85]) & ~(inputs[248]);
    assign layer0_outputs[2874] = (inputs[82]) ^ (inputs[87]);
    assign layer0_outputs[2875] = (inputs[3]) | (inputs[178]);
    assign layer0_outputs[2876] = ~(inputs[14]);
    assign layer0_outputs[2877] = ~(inputs[219]);
    assign layer0_outputs[2878] = (inputs[77]) & ~(inputs[30]);
    assign layer0_outputs[2879] = ~(inputs[66]);
    assign layer0_outputs[2880] = ~((inputs[255]) | (inputs[54]));
    assign layer0_outputs[2881] = (inputs[196]) & ~(inputs[74]);
    assign layer0_outputs[2882] = ~((inputs[42]) | (inputs[169]));
    assign layer0_outputs[2883] = ~(inputs[95]) | (inputs[43]);
    assign layer0_outputs[2884] = ~((inputs[6]) | (inputs[130]));
    assign layer0_outputs[2885] = (inputs[73]) ^ (inputs[117]);
    assign layer0_outputs[2886] = ~(inputs[46]);
    assign layer0_outputs[2887] = (inputs[221]) | (inputs[253]);
    assign layer0_outputs[2888] = ~(inputs[92]);
    assign layer0_outputs[2889] = inputs[141];
    assign layer0_outputs[2890] = (inputs[203]) ^ (inputs[84]);
    assign layer0_outputs[2891] = ~(inputs[76]);
    assign layer0_outputs[2892] = ~(inputs[142]);
    assign layer0_outputs[2893] = (inputs[168]) & (inputs[40]);
    assign layer0_outputs[2894] = ~(inputs[103]) | (inputs[129]);
    assign layer0_outputs[2895] = inputs[193];
    assign layer0_outputs[2896] = ~((inputs[146]) | (inputs[35]));
    assign layer0_outputs[2897] = ~((inputs[241]) ^ (inputs[161]));
    assign layer0_outputs[2898] = ~((inputs[108]) & (inputs[75]));
    assign layer0_outputs[2899] = ~(inputs[69]) | (inputs[194]);
    assign layer0_outputs[2900] = (inputs[222]) | (inputs[55]);
    assign layer0_outputs[2901] = (inputs[18]) | (inputs[166]);
    assign layer0_outputs[2902] = ~((inputs[171]) | (inputs[8]));
    assign layer0_outputs[2903] = (inputs[172]) & ~(inputs[94]);
    assign layer0_outputs[2904] = ~((inputs[172]) & (inputs[236]));
    assign layer0_outputs[2905] = inputs[187];
    assign layer0_outputs[2906] = ~(inputs[209]) | (inputs[138]);
    assign layer0_outputs[2907] = ~((inputs[202]) & (inputs[7]));
    assign layer0_outputs[2908] = (inputs[42]) & ~(inputs[219]);
    assign layer0_outputs[2909] = ~(inputs[188]) | (inputs[110]);
    assign layer0_outputs[2910] = ~((inputs[128]) | (inputs[45]));
    assign layer0_outputs[2911] = inputs[113];
    assign layer0_outputs[2912] = ~(inputs[83]) | (inputs[28]);
    assign layer0_outputs[2913] = ~((inputs[137]) ^ (inputs[156]));
    assign layer0_outputs[2914] = (inputs[231]) & ~(inputs[146]);
    assign layer0_outputs[2915] = ~(inputs[26]) | (inputs[226]);
    assign layer0_outputs[2916] = ~(inputs[19]);
    assign layer0_outputs[2917] = (inputs[192]) ^ (inputs[88]);
    assign layer0_outputs[2918] = inputs[151];
    assign layer0_outputs[2919] = ~(inputs[30]);
    assign layer0_outputs[2920] = ~((inputs[82]) ^ (inputs[177]));
    assign layer0_outputs[2921] = ~(inputs[231]);
    assign layer0_outputs[2922] = (inputs[60]) | (inputs[33]);
    assign layer0_outputs[2923] = ~(inputs[82]) | (inputs[251]);
    assign layer0_outputs[2924] = (inputs[229]) | (inputs[207]);
    assign layer0_outputs[2925] = inputs[193];
    assign layer0_outputs[2926] = ~(inputs[200]) | (inputs[79]);
    assign layer0_outputs[2927] = ~((inputs[52]) | (inputs[160]));
    assign layer0_outputs[2928] = (inputs[165]) ^ (inputs[147]);
    assign layer0_outputs[2929] = ~((inputs[77]) | (inputs[77]));
    assign layer0_outputs[2930] = ~(inputs[161]);
    assign layer0_outputs[2931] = (inputs[51]) | (inputs[146]);
    assign layer0_outputs[2932] = inputs[120];
    assign layer0_outputs[2933] = (inputs[30]) | (inputs[140]);
    assign layer0_outputs[2934] = ~(inputs[43]) | (inputs[227]);
    assign layer0_outputs[2935] = ~((inputs[189]) ^ (inputs[178]));
    assign layer0_outputs[2936] = (inputs[12]) ^ (inputs[71]);
    assign layer0_outputs[2937] = ~(inputs[49]);
    assign layer0_outputs[2938] = ~(inputs[18]);
    assign layer0_outputs[2939] = ~((inputs[124]) ^ (inputs[113]));
    assign layer0_outputs[2940] = ~((inputs[200]) | (inputs[109]));
    assign layer0_outputs[2941] = inputs[58];
    assign layer0_outputs[2942] = (inputs[198]) & (inputs[87]);
    assign layer0_outputs[2943] = ~((inputs[115]) & (inputs[241]));
    assign layer0_outputs[2944] = ~(inputs[89]);
    assign layer0_outputs[2945] = inputs[167];
    assign layer0_outputs[2946] = ~(inputs[123]) | (inputs[205]);
    assign layer0_outputs[2947] = ~(inputs[31]) | (inputs[244]);
    assign layer0_outputs[2948] = (inputs[197]) & ~(inputs[240]);
    assign layer0_outputs[2949] = (inputs[217]) ^ (inputs[93]);
    assign layer0_outputs[2950] = (inputs[77]) | (inputs[164]);
    assign layer0_outputs[2951] = ~((inputs[142]) | (inputs[203]));
    assign layer0_outputs[2952] = (inputs[9]) & ~(inputs[145]);
    assign layer0_outputs[2953] = ~(inputs[3]) | (inputs[241]);
    assign layer0_outputs[2954] = inputs[10];
    assign layer0_outputs[2955] = inputs[119];
    assign layer0_outputs[2956] = ~(inputs[115]);
    assign layer0_outputs[2957] = ~((inputs[162]) ^ (inputs[248]));
    assign layer0_outputs[2958] = (inputs[228]) | (inputs[148]);
    assign layer0_outputs[2959] = (inputs[128]) & ~(inputs[253]);
    assign layer0_outputs[2960] = inputs[103];
    assign layer0_outputs[2961] = (inputs[184]) ^ (inputs[215]);
    assign layer0_outputs[2962] = ~(inputs[131]) | (inputs[13]);
    assign layer0_outputs[2963] = ~(inputs[62]) | (inputs[108]);
    assign layer0_outputs[2964] = 1'b1;
    assign layer0_outputs[2965] = ~((inputs[88]) & (inputs[1]));
    assign layer0_outputs[2966] = ~((inputs[190]) ^ (inputs[42]));
    assign layer0_outputs[2967] = ~(inputs[19]) | (inputs[129]);
    assign layer0_outputs[2968] = (inputs[22]) ^ (inputs[102]);
    assign layer0_outputs[2969] = (inputs[42]) & ~(inputs[146]);
    assign layer0_outputs[2970] = 1'b1;
    assign layer0_outputs[2971] = (inputs[13]) | (inputs[212]);
    assign layer0_outputs[2972] = ~((inputs[70]) | (inputs[73]));
    assign layer0_outputs[2973] = (inputs[18]) | (inputs[238]);
    assign layer0_outputs[2974] = inputs[178];
    assign layer0_outputs[2975] = ~(inputs[209]) | (inputs[5]);
    assign layer0_outputs[2976] = ~(inputs[196]);
    assign layer0_outputs[2977] = (inputs[17]) | (inputs[213]);
    assign layer0_outputs[2978] = (inputs[136]) & ~(inputs[208]);
    assign layer0_outputs[2979] = ~((inputs[224]) ^ (inputs[206]));
    assign layer0_outputs[2980] = (inputs[69]) & ~(inputs[77]);
    assign layer0_outputs[2981] = 1'b0;
    assign layer0_outputs[2982] = inputs[202];
    assign layer0_outputs[2983] = (inputs[208]) ^ (inputs[183]);
    assign layer0_outputs[2984] = (inputs[252]) | (inputs[81]);
    assign layer0_outputs[2985] = ~((inputs[138]) | (inputs[207]));
    assign layer0_outputs[2986] = (inputs[205]) & ~(inputs[31]);
    assign layer0_outputs[2987] = ~((inputs[78]) | (inputs[126]));
    assign layer0_outputs[2988] = ~((inputs[255]) ^ (inputs[56]));
    assign layer0_outputs[2989] = (inputs[25]) | (inputs[155]);
    assign layer0_outputs[2990] = (inputs[197]) & ~(inputs[112]);
    assign layer0_outputs[2991] = (inputs[18]) | (inputs[178]);
    assign layer0_outputs[2992] = (inputs[228]) | (inputs[114]);
    assign layer0_outputs[2993] = (inputs[222]) ^ (inputs[156]);
    assign layer0_outputs[2994] = inputs[211];
    assign layer0_outputs[2995] = (inputs[190]) ^ (inputs[238]);
    assign layer0_outputs[2996] = inputs[162];
    assign layer0_outputs[2997] = (inputs[37]) | (inputs[87]);
    assign layer0_outputs[2998] = 1'b0;
    assign layer0_outputs[2999] = ~((inputs[191]) | (inputs[235]));
    assign layer0_outputs[3000] = (inputs[80]) ^ (inputs[60]);
    assign layer0_outputs[3001] = (inputs[40]) & ~(inputs[243]);
    assign layer0_outputs[3002] = inputs[162];
    assign layer0_outputs[3003] = ~(inputs[37]);
    assign layer0_outputs[3004] = ~((inputs[0]) | (inputs[12]));
    assign layer0_outputs[3005] = (inputs[139]) ^ (inputs[189]);
    assign layer0_outputs[3006] = (inputs[76]) & (inputs[96]);
    assign layer0_outputs[3007] = inputs[157];
    assign layer0_outputs[3008] = ~(inputs[220]) | (inputs[244]);
    assign layer0_outputs[3009] = (inputs[98]) & ~(inputs[94]);
    assign layer0_outputs[3010] = ~(inputs[226]) | (inputs[54]);
    assign layer0_outputs[3011] = ~((inputs[70]) ^ (inputs[53]));
    assign layer0_outputs[3012] = ~((inputs[245]) | (inputs[143]));
    assign layer0_outputs[3013] = inputs[118];
    assign layer0_outputs[3014] = inputs[130];
    assign layer0_outputs[3015] = ~((inputs[24]) | (inputs[191]));
    assign layer0_outputs[3016] = inputs[27];
    assign layer0_outputs[3017] = ~(inputs[173]);
    assign layer0_outputs[3018] = (inputs[205]) ^ (inputs[95]);
    assign layer0_outputs[3019] = ~(inputs[197]);
    assign layer0_outputs[3020] = ~(inputs[26]) | (inputs[241]);
    assign layer0_outputs[3021] = (inputs[185]) & (inputs[31]);
    assign layer0_outputs[3022] = (inputs[85]) & ~(inputs[48]);
    assign layer0_outputs[3023] = ~((inputs[102]) | (inputs[69]));
    assign layer0_outputs[3024] = (inputs[74]) & ~(inputs[197]);
    assign layer0_outputs[3025] = ~((inputs[219]) ^ (inputs[37]));
    assign layer0_outputs[3026] = inputs[180];
    assign layer0_outputs[3027] = ~((inputs[181]) ^ (inputs[138]));
    assign layer0_outputs[3028] = ~((inputs[135]) ^ (inputs[33]));
    assign layer0_outputs[3029] = (inputs[174]) & ~(inputs[94]);
    assign layer0_outputs[3030] = (inputs[150]) & ~(inputs[97]);
    assign layer0_outputs[3031] = inputs[164];
    assign layer0_outputs[3032] = inputs[120];
    assign layer0_outputs[3033] = ~(inputs[84]);
    assign layer0_outputs[3034] = (inputs[118]) | (inputs[234]);
    assign layer0_outputs[3035] = (inputs[102]) & ~(inputs[234]);
    assign layer0_outputs[3036] = inputs[90];
    assign layer0_outputs[3037] = (inputs[32]) & ~(inputs[13]);
    assign layer0_outputs[3038] = inputs[105];
    assign layer0_outputs[3039] = (inputs[137]) & ~(inputs[213]);
    assign layer0_outputs[3040] = inputs[93];
    assign layer0_outputs[3041] = ~((inputs[137]) ^ (inputs[131]));
    assign layer0_outputs[3042] = (inputs[170]) ^ (inputs[136]);
    assign layer0_outputs[3043] = (inputs[26]) ^ (inputs[36]);
    assign layer0_outputs[3044] = ~(inputs[229]);
    assign layer0_outputs[3045] = inputs[197];
    assign layer0_outputs[3046] = inputs[114];
    assign layer0_outputs[3047] = inputs[97];
    assign layer0_outputs[3048] = inputs[203];
    assign layer0_outputs[3049] = ~(inputs[165]) | (inputs[97]);
    assign layer0_outputs[3050] = ~(inputs[41]);
    assign layer0_outputs[3051] = ~((inputs[17]) | (inputs[135]));
    assign layer0_outputs[3052] = ~(inputs[31]);
    assign layer0_outputs[3053] = inputs[50];
    assign layer0_outputs[3054] = ~(inputs[25]);
    assign layer0_outputs[3055] = inputs[125];
    assign layer0_outputs[3056] = ~(inputs[27]);
    assign layer0_outputs[3057] = (inputs[69]) & ~(inputs[239]);
    assign layer0_outputs[3058] = inputs[229];
    assign layer0_outputs[3059] = (inputs[27]) & ~(inputs[254]);
    assign layer0_outputs[3060] = ~((inputs[70]) | (inputs[159]));
    assign layer0_outputs[3061] = ~(inputs[160]);
    assign layer0_outputs[3062] = ~(inputs[75]) | (inputs[176]);
    assign layer0_outputs[3063] = (inputs[168]) | (inputs[49]);
    assign layer0_outputs[3064] = (inputs[247]) & ~(inputs[11]);
    assign layer0_outputs[3065] = ~((inputs[100]) ^ (inputs[76]));
    assign layer0_outputs[3066] = ~(inputs[130]);
    assign layer0_outputs[3067] = ~(inputs[82]);
    assign layer0_outputs[3068] = ~(inputs[208]) | (inputs[174]);
    assign layer0_outputs[3069] = ~((inputs[128]) | (inputs[29]));
    assign layer0_outputs[3070] = (inputs[255]) & (inputs[102]);
    assign layer0_outputs[3071] = ~((inputs[84]) | (inputs[46]));
    assign layer0_outputs[3072] = (inputs[155]) | (inputs[242]);
    assign layer0_outputs[3073] = ~(inputs[215]);
    assign layer0_outputs[3074] = inputs[9];
    assign layer0_outputs[3075] = (inputs[11]) | (inputs[253]);
    assign layer0_outputs[3076] = ~((inputs[82]) & (inputs[243]));
    assign layer0_outputs[3077] = (inputs[3]) | (inputs[219]);
    assign layer0_outputs[3078] = ~(inputs[199]) | (inputs[96]);
    assign layer0_outputs[3079] = inputs[101];
    assign layer0_outputs[3080] = ~((inputs[50]) | (inputs[179]));
    assign layer0_outputs[3081] = inputs[235];
    assign layer0_outputs[3082] = ~((inputs[40]) | (inputs[16]));
    assign layer0_outputs[3083] = ~((inputs[128]) ^ (inputs[148]));
    assign layer0_outputs[3084] = ~(inputs[3]);
    assign layer0_outputs[3085] = (inputs[7]) & (inputs[25]);
    assign layer0_outputs[3086] = ~((inputs[74]) & (inputs[53]));
    assign layer0_outputs[3087] = inputs[178];
    assign layer0_outputs[3088] = ~((inputs[11]) ^ (inputs[46]));
    assign layer0_outputs[3089] = ~((inputs[207]) | (inputs[126]));
    assign layer0_outputs[3090] = ~(inputs[95]) | (inputs[205]);
    assign layer0_outputs[3091] = ~(inputs[108]);
    assign layer0_outputs[3092] = (inputs[60]) & ~(inputs[237]);
    assign layer0_outputs[3093] = (inputs[3]) | (inputs[45]);
    assign layer0_outputs[3094] = inputs[231];
    assign layer0_outputs[3095] = ~(inputs[121]);
    assign layer0_outputs[3096] = (inputs[113]) & ~(inputs[16]);
    assign layer0_outputs[3097] = (inputs[58]) ^ (inputs[86]);
    assign layer0_outputs[3098] = (inputs[246]) ^ (inputs[139]);
    assign layer0_outputs[3099] = ~((inputs[166]) | (inputs[145]));
    assign layer0_outputs[3100] = inputs[233];
    assign layer0_outputs[3101] = ~((inputs[58]) ^ (inputs[10]));
    assign layer0_outputs[3102] = (inputs[241]) & (inputs[79]);
    assign layer0_outputs[3103] = ~((inputs[124]) ^ (inputs[205]));
    assign layer0_outputs[3104] = ~((inputs[243]) | (inputs[217]));
    assign layer0_outputs[3105] = inputs[69];
    assign layer0_outputs[3106] = (inputs[255]) | (inputs[216]);
    assign layer0_outputs[3107] = inputs[23];
    assign layer0_outputs[3108] = (inputs[97]) | (inputs[112]);
    assign layer0_outputs[3109] = ~((inputs[37]) | (inputs[205]));
    assign layer0_outputs[3110] = (inputs[230]) | (inputs[238]);
    assign layer0_outputs[3111] = ~(inputs[83]);
    assign layer0_outputs[3112] = (inputs[56]) | (inputs[16]);
    assign layer0_outputs[3113] = inputs[152];
    assign layer0_outputs[3114] = ~(inputs[29]) | (inputs[176]);
    assign layer0_outputs[3115] = (inputs[117]) & ~(inputs[104]);
    assign layer0_outputs[3116] = inputs[81];
    assign layer0_outputs[3117] = inputs[6];
    assign layer0_outputs[3118] = ~(inputs[93]);
    assign layer0_outputs[3119] = ~((inputs[211]) ^ (inputs[166]));
    assign layer0_outputs[3120] = (inputs[195]) & ~(inputs[175]);
    assign layer0_outputs[3121] = ~(inputs[114]);
    assign layer0_outputs[3122] = ~(inputs[76]) | (inputs[238]);
    assign layer0_outputs[3123] = ~(inputs[94]);
    assign layer0_outputs[3124] = (inputs[74]) & ~(inputs[147]);
    assign layer0_outputs[3125] = (inputs[219]) ^ (inputs[75]);
    assign layer0_outputs[3126] = ~(inputs[203]) | (inputs[251]);
    assign layer0_outputs[3127] = (inputs[98]) | (inputs[154]);
    assign layer0_outputs[3128] = (inputs[142]) ^ (inputs[18]);
    assign layer0_outputs[3129] = inputs[56];
    assign layer0_outputs[3130] = (inputs[236]) | (inputs[147]);
    assign layer0_outputs[3131] = ~(inputs[32]);
    assign layer0_outputs[3132] = (inputs[237]) ^ (inputs[19]);
    assign layer0_outputs[3133] = inputs[208];
    assign layer0_outputs[3134] = ~((inputs[97]) | (inputs[124]));
    assign layer0_outputs[3135] = ~(inputs[148]);
    assign layer0_outputs[3136] = ~(inputs[147]);
    assign layer0_outputs[3137] = ~(inputs[165]);
    assign layer0_outputs[3138] = ~((inputs[195]) ^ (inputs[89]));
    assign layer0_outputs[3139] = (inputs[116]) & ~(inputs[194]);
    assign layer0_outputs[3140] = ~(inputs[57]);
    assign layer0_outputs[3141] = (inputs[151]) & ~(inputs[85]);
    assign layer0_outputs[3142] = ~(inputs[72]) | (inputs[15]);
    assign layer0_outputs[3143] = ~(inputs[235]);
    assign layer0_outputs[3144] = (inputs[234]) | (inputs[158]);
    assign layer0_outputs[3145] = ~(inputs[221]);
    assign layer0_outputs[3146] = inputs[44];
    assign layer0_outputs[3147] = inputs[72];
    assign layer0_outputs[3148] = ~((inputs[17]) | (inputs[124]));
    assign layer0_outputs[3149] = ~(inputs[206]);
    assign layer0_outputs[3150] = inputs[19];
    assign layer0_outputs[3151] = ~((inputs[202]) ^ (inputs[54]));
    assign layer0_outputs[3152] = (inputs[200]) & ~(inputs[67]);
    assign layer0_outputs[3153] = (inputs[224]) & ~(inputs[122]);
    assign layer0_outputs[3154] = inputs[31];
    assign layer0_outputs[3155] = ~((inputs[112]) ^ (inputs[26]));
    assign layer0_outputs[3156] = ~((inputs[194]) ^ (inputs[81]));
    assign layer0_outputs[3157] = ~(inputs[82]) | (inputs[73]);
    assign layer0_outputs[3158] = (inputs[106]) & ~(inputs[18]);
    assign layer0_outputs[3159] = ~((inputs[211]) | (inputs[104]));
    assign layer0_outputs[3160] = (inputs[228]) ^ (inputs[24]);
    assign layer0_outputs[3161] = ~((inputs[71]) & (inputs[161]));
    assign layer0_outputs[3162] = ~(inputs[118]);
    assign layer0_outputs[3163] = ~(inputs[23]);
    assign layer0_outputs[3164] = (inputs[179]) | (inputs[158]);
    assign layer0_outputs[3165] = (inputs[76]) | (inputs[210]);
    assign layer0_outputs[3166] = ~(inputs[4]) | (inputs[84]);
    assign layer0_outputs[3167] = ~((inputs[48]) | (inputs[151]));
    assign layer0_outputs[3168] = inputs[214];
    assign layer0_outputs[3169] = ~(inputs[240]);
    assign layer0_outputs[3170] = (inputs[90]) | (inputs[18]);
    assign layer0_outputs[3171] = ~(inputs[107]);
    assign layer0_outputs[3172] = (inputs[217]) & ~(inputs[90]);
    assign layer0_outputs[3173] = ~(inputs[105]) | (inputs[46]);
    assign layer0_outputs[3174] = (inputs[144]) | (inputs[212]);
    assign layer0_outputs[3175] = (inputs[205]) & ~(inputs[109]);
    assign layer0_outputs[3176] = (inputs[13]) | (inputs[138]);
    assign layer0_outputs[3177] = ~(inputs[90]) | (inputs[192]);
    assign layer0_outputs[3178] = inputs[78];
    assign layer0_outputs[3179] = ~((inputs[51]) | (inputs[129]));
    assign layer0_outputs[3180] = (inputs[106]) ^ (inputs[136]);
    assign layer0_outputs[3181] = (inputs[35]) ^ (inputs[149]);
    assign layer0_outputs[3182] = ~((inputs[40]) | (inputs[171]));
    assign layer0_outputs[3183] = ~(inputs[45]) | (inputs[182]);
    assign layer0_outputs[3184] = ~(inputs[27]) | (inputs[3]);
    assign layer0_outputs[3185] = ~(inputs[174]);
    assign layer0_outputs[3186] = ~(inputs[177]);
    assign layer0_outputs[3187] = (inputs[78]) ^ (inputs[63]);
    assign layer0_outputs[3188] = ~(inputs[20]) | (inputs[178]);
    assign layer0_outputs[3189] = ~(inputs[127]);
    assign layer0_outputs[3190] = ~(inputs[138]) | (inputs[49]);
    assign layer0_outputs[3191] = inputs[20];
    assign layer0_outputs[3192] = inputs[78];
    assign layer0_outputs[3193] = ~(inputs[188]);
    assign layer0_outputs[3194] = ~((inputs[190]) | (inputs[217]));
    assign layer0_outputs[3195] = ~(inputs[224]) | (inputs[49]);
    assign layer0_outputs[3196] = (inputs[175]) | (inputs[229]);
    assign layer0_outputs[3197] = (inputs[200]) & ~(inputs[227]);
    assign layer0_outputs[3198] = (inputs[166]) ^ (inputs[196]);
    assign layer0_outputs[3199] = 1'b1;
    assign layer0_outputs[3200] = (inputs[71]) & ~(inputs[206]);
    assign layer0_outputs[3201] = ~((inputs[111]) ^ (inputs[235]));
    assign layer0_outputs[3202] = (inputs[11]) | (inputs[147]);
    assign layer0_outputs[3203] = ~(inputs[151]) | (inputs[157]);
    assign layer0_outputs[3204] = (inputs[31]) & ~(inputs[136]);
    assign layer0_outputs[3205] = ~(inputs[232]);
    assign layer0_outputs[3206] = (inputs[47]) & ~(inputs[209]);
    assign layer0_outputs[3207] = (inputs[234]) & ~(inputs[143]);
    assign layer0_outputs[3208] = 1'b0;
    assign layer0_outputs[3209] = ~(inputs[111]);
    assign layer0_outputs[3210] = ~(inputs[184]) | (inputs[192]);
    assign layer0_outputs[3211] = ~((inputs[22]) | (inputs[188]));
    assign layer0_outputs[3212] = ~(inputs[210]) | (inputs[247]);
    assign layer0_outputs[3213] = ~(inputs[99]);
    assign layer0_outputs[3214] = ~(inputs[63]);
    assign layer0_outputs[3215] = ~(inputs[164]);
    assign layer0_outputs[3216] = ~((inputs[219]) | (inputs[225]));
    assign layer0_outputs[3217] = inputs[230];
    assign layer0_outputs[3218] = ~(inputs[61]);
    assign layer0_outputs[3219] = (inputs[255]) | (inputs[193]);
    assign layer0_outputs[3220] = (inputs[63]) ^ (inputs[203]);
    assign layer0_outputs[3221] = ~((inputs[214]) | (inputs[97]));
    assign layer0_outputs[3222] = ~(inputs[58]) | (inputs[186]);
    assign layer0_outputs[3223] = ~((inputs[32]) ^ (inputs[132]));
    assign layer0_outputs[3224] = ~((inputs[3]) | (inputs[4]));
    assign layer0_outputs[3225] = ~(inputs[248]);
    assign layer0_outputs[3226] = inputs[37];
    assign layer0_outputs[3227] = (inputs[6]) & ~(inputs[145]);
    assign layer0_outputs[3228] = ~(inputs[21]) | (inputs[99]);
    assign layer0_outputs[3229] = 1'b0;
    assign layer0_outputs[3230] = (inputs[84]) & (inputs[230]);
    assign layer0_outputs[3231] = inputs[148];
    assign layer0_outputs[3232] = ~(inputs[94]);
    assign layer0_outputs[3233] = inputs[164];
    assign layer0_outputs[3234] = ~((inputs[169]) ^ (inputs[22]));
    assign layer0_outputs[3235] = ~(inputs[71]) | (inputs[233]);
    assign layer0_outputs[3236] = ~((inputs[149]) ^ (inputs[252]));
    assign layer0_outputs[3237] = ~((inputs[120]) & (inputs[233]));
    assign layer0_outputs[3238] = (inputs[71]) | (inputs[128]);
    assign layer0_outputs[3239] = inputs[208];
    assign layer0_outputs[3240] = (inputs[121]) ^ (inputs[254]);
    assign layer0_outputs[3241] = (inputs[84]) & ~(inputs[236]);
    assign layer0_outputs[3242] = inputs[94];
    assign layer0_outputs[3243] = inputs[110];
    assign layer0_outputs[3244] = (inputs[154]) & ~(inputs[242]);
    assign layer0_outputs[3245] = ~(inputs[235]);
    assign layer0_outputs[3246] = inputs[56];
    assign layer0_outputs[3247] = ~((inputs[242]) ^ (inputs[167]));
    assign layer0_outputs[3248] = (inputs[187]) | (inputs[172]);
    assign layer0_outputs[3249] = (inputs[107]) & ~(inputs[141]);
    assign layer0_outputs[3250] = (inputs[194]) | (inputs[204]);
    assign layer0_outputs[3251] = ~((inputs[233]) | (inputs[5]));
    assign layer0_outputs[3252] = inputs[71];
    assign layer0_outputs[3253] = ~(inputs[30]);
    assign layer0_outputs[3254] = ~((inputs[182]) | (inputs[147]));
    assign layer0_outputs[3255] = ~((inputs[234]) | (inputs[144]));
    assign layer0_outputs[3256] = ~((inputs[8]) & (inputs[22]));
    assign layer0_outputs[3257] = ~(inputs[210]);
    assign layer0_outputs[3258] = inputs[68];
    assign layer0_outputs[3259] = ~((inputs[124]) | (inputs[26]));
    assign layer0_outputs[3260] = ~(inputs[45]);
    assign layer0_outputs[3261] = ~((inputs[196]) | (inputs[230]));
    assign layer0_outputs[3262] = ~(inputs[88]);
    assign layer0_outputs[3263] = inputs[246];
    assign layer0_outputs[3264] = inputs[118];
    assign layer0_outputs[3265] = ~(inputs[72]);
    assign layer0_outputs[3266] = (inputs[153]) | (inputs[127]);
    assign layer0_outputs[3267] = (inputs[3]) & ~(inputs[255]);
    assign layer0_outputs[3268] = ~((inputs[228]) | (inputs[102]));
    assign layer0_outputs[3269] = (inputs[63]) ^ (inputs[75]);
    assign layer0_outputs[3270] = (inputs[121]) & ~(inputs[164]);
    assign layer0_outputs[3271] = ~((inputs[135]) | (inputs[130]));
    assign layer0_outputs[3272] = inputs[108];
    assign layer0_outputs[3273] = inputs[8];
    assign layer0_outputs[3274] = ~(inputs[221]);
    assign layer0_outputs[3275] = ~(inputs[36]);
    assign layer0_outputs[3276] = ~(inputs[251]);
    assign layer0_outputs[3277] = (inputs[244]) ^ (inputs[22]);
    assign layer0_outputs[3278] = ~(inputs[122]);
    assign layer0_outputs[3279] = ~(inputs[19]);
    assign layer0_outputs[3280] = ~(inputs[33]);
    assign layer0_outputs[3281] = (inputs[10]) & ~(inputs[65]);
    assign layer0_outputs[3282] = ~((inputs[138]) | (inputs[30]));
    assign layer0_outputs[3283] = ~((inputs[177]) | (inputs[67]));
    assign layer0_outputs[3284] = ~(inputs[154]) | (inputs[116]);
    assign layer0_outputs[3285] = (inputs[107]) ^ (inputs[67]);
    assign layer0_outputs[3286] = ~((inputs[6]) ^ (inputs[36]));
    assign layer0_outputs[3287] = ~((inputs[122]) | (inputs[14]));
    assign layer0_outputs[3288] = inputs[157];
    assign layer0_outputs[3289] = ~(inputs[117]);
    assign layer0_outputs[3290] = (inputs[146]) & ~(inputs[80]);
    assign layer0_outputs[3291] = inputs[66];
    assign layer0_outputs[3292] = 1'b0;
    assign layer0_outputs[3293] = inputs[194];
    assign layer0_outputs[3294] = ~(inputs[212]) | (inputs[90]);
    assign layer0_outputs[3295] = inputs[185];
    assign layer0_outputs[3296] = ~((inputs[18]) | (inputs[211]));
    assign layer0_outputs[3297] = ~((inputs[134]) ^ (inputs[101]));
    assign layer0_outputs[3298] = (inputs[219]) ^ (inputs[52]);
    assign layer0_outputs[3299] = (inputs[17]) ^ (inputs[187]);
    assign layer0_outputs[3300] = ~((inputs[1]) | (inputs[170]));
    assign layer0_outputs[3301] = ~((inputs[39]) ^ (inputs[215]));
    assign layer0_outputs[3302] = ~(inputs[125]);
    assign layer0_outputs[3303] = (inputs[158]) | (inputs[100]);
    assign layer0_outputs[3304] = ~((inputs[222]) | (inputs[228]));
    assign layer0_outputs[3305] = (inputs[59]) & ~(inputs[207]);
    assign layer0_outputs[3306] = ~(inputs[83]);
    assign layer0_outputs[3307] = ~((inputs[18]) | (inputs[31]));
    assign layer0_outputs[3308] = ~(inputs[84]);
    assign layer0_outputs[3309] = inputs[145];
    assign layer0_outputs[3310] = (inputs[117]) ^ (inputs[88]);
    assign layer0_outputs[3311] = (inputs[255]) | (inputs[198]);
    assign layer0_outputs[3312] = inputs[115];
    assign layer0_outputs[3313] = ~(inputs[231]);
    assign layer0_outputs[3314] = ~(inputs[103]) | (inputs[94]);
    assign layer0_outputs[3315] = (inputs[155]) | (inputs[145]);
    assign layer0_outputs[3316] = ~((inputs[5]) & (inputs[6]));
    assign layer0_outputs[3317] = ~(inputs[180]) | (inputs[41]);
    assign layer0_outputs[3318] = (inputs[173]) & ~(inputs[169]);
    assign layer0_outputs[3319] = inputs[21];
    assign layer0_outputs[3320] = ~(inputs[137]);
    assign layer0_outputs[3321] = inputs[1];
    assign layer0_outputs[3322] = ~(inputs[83]);
    assign layer0_outputs[3323] = ~(inputs[88]) | (inputs[79]);
    assign layer0_outputs[3324] = inputs[127];
    assign layer0_outputs[3325] = (inputs[193]) & ~(inputs[67]);
    assign layer0_outputs[3326] = (inputs[10]) & ~(inputs[111]);
    assign layer0_outputs[3327] = ~(inputs[58]) | (inputs[183]);
    assign layer0_outputs[3328] = inputs[166];
    assign layer0_outputs[3329] = ~(inputs[138]);
    assign layer0_outputs[3330] = (inputs[179]) | (inputs[109]);
    assign layer0_outputs[3331] = inputs[225];
    assign layer0_outputs[3332] = (inputs[244]) | (inputs[249]);
    assign layer0_outputs[3333] = (inputs[177]) ^ (inputs[216]);
    assign layer0_outputs[3334] = ~(inputs[230]);
    assign layer0_outputs[3335] = ~(inputs[15]) | (inputs[77]);
    assign layer0_outputs[3336] = ~(inputs[233]);
    assign layer0_outputs[3337] = (inputs[99]) & ~(inputs[174]);
    assign layer0_outputs[3338] = ~(inputs[168]);
    assign layer0_outputs[3339] = ~(inputs[163]);
    assign layer0_outputs[3340] = (inputs[219]) ^ (inputs[208]);
    assign layer0_outputs[3341] = (inputs[129]) | (inputs[174]);
    assign layer0_outputs[3342] = (inputs[115]) ^ (inputs[84]);
    assign layer0_outputs[3343] = (inputs[195]) | (inputs[196]);
    assign layer0_outputs[3344] = ~(inputs[61]);
    assign layer0_outputs[3345] = ~((inputs[182]) | (inputs[33]));
    assign layer0_outputs[3346] = ~(inputs[172]) | (inputs[236]);
    assign layer0_outputs[3347] = ~((inputs[93]) ^ (inputs[2]));
    assign layer0_outputs[3348] = ~((inputs[11]) | (inputs[249]));
    assign layer0_outputs[3349] = ~((inputs[138]) | (inputs[251]));
    assign layer0_outputs[3350] = ~(inputs[216]) | (inputs[239]);
    assign layer0_outputs[3351] = ~(inputs[228]) | (inputs[42]);
    assign layer0_outputs[3352] = (inputs[33]) | (inputs[172]);
    assign layer0_outputs[3353] = (inputs[119]) ^ (inputs[159]);
    assign layer0_outputs[3354] = inputs[101];
    assign layer0_outputs[3355] = ~(inputs[243]);
    assign layer0_outputs[3356] = inputs[123];
    assign layer0_outputs[3357] = inputs[102];
    assign layer0_outputs[3358] = (inputs[204]) & ~(inputs[84]);
    assign layer0_outputs[3359] = ~(inputs[15]);
    assign layer0_outputs[3360] = ~(inputs[230]);
    assign layer0_outputs[3361] = ~(inputs[227]);
    assign layer0_outputs[3362] = (inputs[180]) & ~(inputs[165]);
    assign layer0_outputs[3363] = ~((inputs[52]) ^ (inputs[95]));
    assign layer0_outputs[3364] = ~((inputs[219]) ^ (inputs[142]));
    assign layer0_outputs[3365] = ~(inputs[236]) | (inputs[149]);
    assign layer0_outputs[3366] = inputs[120];
    assign layer0_outputs[3367] = ~((inputs[214]) ^ (inputs[46]));
    assign layer0_outputs[3368] = ~(inputs[68]) | (inputs[172]);
    assign layer0_outputs[3369] = inputs[135];
    assign layer0_outputs[3370] = ~((inputs[3]) | (inputs[21]));
    assign layer0_outputs[3371] = ~((inputs[120]) ^ (inputs[187]));
    assign layer0_outputs[3372] = (inputs[39]) & ~(inputs[199]);
    assign layer0_outputs[3373] = ~(inputs[3]);
    assign layer0_outputs[3374] = ~(inputs[79]) | (inputs[78]);
    assign layer0_outputs[3375] = ~((inputs[185]) ^ (inputs[236]));
    assign layer0_outputs[3376] = ~(inputs[207]) | (inputs[191]);
    assign layer0_outputs[3377] = (inputs[226]) & ~(inputs[129]);
    assign layer0_outputs[3378] = ~(inputs[162]);
    assign layer0_outputs[3379] = ~(inputs[22]) | (inputs[193]);
    assign layer0_outputs[3380] = (inputs[132]) & ~(inputs[75]);
    assign layer0_outputs[3381] = (inputs[65]) | (inputs[12]);
    assign layer0_outputs[3382] = (inputs[248]) & ~(inputs[118]);
    assign layer0_outputs[3383] = ~((inputs[224]) | (inputs[232]));
    assign layer0_outputs[3384] = (inputs[90]) | (inputs[4]);
    assign layer0_outputs[3385] = ~(inputs[84]) | (inputs[206]);
    assign layer0_outputs[3386] = ~(inputs[244]);
    assign layer0_outputs[3387] = 1'b1;
    assign layer0_outputs[3388] = ~((inputs[160]) | (inputs[232]));
    assign layer0_outputs[3389] = 1'b1;
    assign layer0_outputs[3390] = inputs[35];
    assign layer0_outputs[3391] = ~((inputs[243]) | (inputs[74]));
    assign layer0_outputs[3392] = (inputs[152]) & ~(inputs[46]);
    assign layer0_outputs[3393] = (inputs[83]) | (inputs[45]);
    assign layer0_outputs[3394] = ~(inputs[83]) | (inputs[136]);
    assign layer0_outputs[3395] = (inputs[123]) & ~(inputs[186]);
    assign layer0_outputs[3396] = ~((inputs[42]) ^ (inputs[143]));
    assign layer0_outputs[3397] = ~(inputs[170]) | (inputs[196]);
    assign layer0_outputs[3398] = ~((inputs[201]) ^ (inputs[234]));
    assign layer0_outputs[3399] = ~(inputs[13]) | (inputs[224]);
    assign layer0_outputs[3400] = ~(inputs[195]);
    assign layer0_outputs[3401] = (inputs[127]) | (inputs[42]);
    assign layer0_outputs[3402] = inputs[59];
    assign layer0_outputs[3403] = ~(inputs[180]);
    assign layer0_outputs[3404] = (inputs[90]) & ~(inputs[170]);
    assign layer0_outputs[3405] = (inputs[223]) & ~(inputs[47]);
    assign layer0_outputs[3406] = ~((inputs[53]) | (inputs[246]));
    assign layer0_outputs[3407] = ~((inputs[236]) ^ (inputs[188]));
    assign layer0_outputs[3408] = ~((inputs[179]) | (inputs[158]));
    assign layer0_outputs[3409] = inputs[230];
    assign layer0_outputs[3410] = inputs[158];
    assign layer0_outputs[3411] = (inputs[101]) & ~(inputs[190]);
    assign layer0_outputs[3412] = ~((inputs[232]) | (inputs[176]));
    assign layer0_outputs[3413] = (inputs[102]) | (inputs[199]);
    assign layer0_outputs[3414] = ~(inputs[93]);
    assign layer0_outputs[3415] = ~(inputs[248]);
    assign layer0_outputs[3416] = ~(inputs[6]);
    assign layer0_outputs[3417] = ~((inputs[9]) | (inputs[171]));
    assign layer0_outputs[3418] = (inputs[149]) & ~(inputs[76]);
    assign layer0_outputs[3419] = (inputs[209]) & ~(inputs[141]);
    assign layer0_outputs[3420] = (inputs[138]) | (inputs[184]);
    assign layer0_outputs[3421] = ~(inputs[195]) | (inputs[112]);
    assign layer0_outputs[3422] = (inputs[2]) | (inputs[225]);
    assign layer0_outputs[3423] = ~((inputs[161]) & (inputs[51]));
    assign layer0_outputs[3424] = (inputs[104]) & ~(inputs[170]);
    assign layer0_outputs[3425] = (inputs[169]) & ~(inputs[79]);
    assign layer0_outputs[3426] = ~(inputs[68]);
    assign layer0_outputs[3427] = (inputs[24]) ^ (inputs[159]);
    assign layer0_outputs[3428] = 1'b0;
    assign layer0_outputs[3429] = inputs[106];
    assign layer0_outputs[3430] = (inputs[195]) & ~(inputs[255]);
    assign layer0_outputs[3431] = ~((inputs[199]) & (inputs[179]));
    assign layer0_outputs[3432] = ~(inputs[93]);
    assign layer0_outputs[3433] = ~(inputs[107]) | (inputs[37]);
    assign layer0_outputs[3434] = (inputs[70]) | (inputs[172]);
    assign layer0_outputs[3435] = inputs[58];
    assign layer0_outputs[3436] = ~((inputs[224]) & (inputs[86]));
    assign layer0_outputs[3437] = ~((inputs[68]) | (inputs[102]));
    assign layer0_outputs[3438] = (inputs[171]) | (inputs[223]);
    assign layer0_outputs[3439] = ~(inputs[134]);
    assign layer0_outputs[3440] = ~(inputs[34]);
    assign layer0_outputs[3441] = ~(inputs[199]) | (inputs[65]);
    assign layer0_outputs[3442] = ~(inputs[101]);
    assign layer0_outputs[3443] = ~(inputs[103]);
    assign layer0_outputs[3444] = ~((inputs[66]) | (inputs[86]));
    assign layer0_outputs[3445] = (inputs[240]) & (inputs[186]);
    assign layer0_outputs[3446] = (inputs[75]) | (inputs[135]);
    assign layer0_outputs[3447] = (inputs[205]) & ~(inputs[126]);
    assign layer0_outputs[3448] = (inputs[8]) & ~(inputs[208]);
    assign layer0_outputs[3449] = inputs[142];
    assign layer0_outputs[3450] = (inputs[17]) | (inputs[60]);
    assign layer0_outputs[3451] = ~(inputs[208]) | (inputs[12]);
    assign layer0_outputs[3452] = ~(inputs[160]) | (inputs[158]);
    assign layer0_outputs[3453] = ~((inputs[152]) | (inputs[219]));
    assign layer0_outputs[3454] = inputs[121];
    assign layer0_outputs[3455] = 1'b1;
    assign layer0_outputs[3456] = ~(inputs[246]);
    assign layer0_outputs[3457] = (inputs[65]) & ~(inputs[209]);
    assign layer0_outputs[3458] = ~((inputs[101]) | (inputs[12]));
    assign layer0_outputs[3459] = ~(inputs[89]) | (inputs[216]);
    assign layer0_outputs[3460] = ~((inputs[203]) ^ (inputs[235]));
    assign layer0_outputs[3461] = (inputs[217]) | (inputs[194]);
    assign layer0_outputs[3462] = ~((inputs[247]) | (inputs[174]));
    assign layer0_outputs[3463] = (inputs[19]) | (inputs[1]);
    assign layer0_outputs[3464] = ~(inputs[11]);
    assign layer0_outputs[3465] = (inputs[78]) | (inputs[199]);
    assign layer0_outputs[3466] = inputs[20];
    assign layer0_outputs[3467] = inputs[208];
    assign layer0_outputs[3468] = inputs[157];
    assign layer0_outputs[3469] = (inputs[169]) & ~(inputs[152]);
    assign layer0_outputs[3470] = inputs[210];
    assign layer0_outputs[3471] = (inputs[207]) | (inputs[251]);
    assign layer0_outputs[3472] = (inputs[224]) ^ (inputs[64]);
    assign layer0_outputs[3473] = (inputs[21]) & ~(inputs[162]);
    assign layer0_outputs[3474] = inputs[87];
    assign layer0_outputs[3475] = (inputs[230]) & ~(inputs[221]);
    assign layer0_outputs[3476] = ~((inputs[211]) ^ (inputs[118]));
    assign layer0_outputs[3477] = (inputs[189]) | (inputs[193]);
    assign layer0_outputs[3478] = inputs[69];
    assign layer0_outputs[3479] = (inputs[219]) | (inputs[185]);
    assign layer0_outputs[3480] = ~(inputs[77]);
    assign layer0_outputs[3481] = ~((inputs[70]) ^ (inputs[89]));
    assign layer0_outputs[3482] = (inputs[180]) ^ (inputs[192]);
    assign layer0_outputs[3483] = ~(inputs[169]) | (inputs[131]);
    assign layer0_outputs[3484] = ~(inputs[231]);
    assign layer0_outputs[3485] = inputs[130];
    assign layer0_outputs[3486] = ~(inputs[100]) | (inputs[178]);
    assign layer0_outputs[3487] = ~((inputs[219]) ^ (inputs[186]));
    assign layer0_outputs[3488] = inputs[214];
    assign layer0_outputs[3489] = (inputs[87]) & ~(inputs[180]);
    assign layer0_outputs[3490] = ~(inputs[186]);
    assign layer0_outputs[3491] = ~(inputs[46]);
    assign layer0_outputs[3492] = ~(inputs[148]);
    assign layer0_outputs[3493] = ~(inputs[237]);
    assign layer0_outputs[3494] = (inputs[198]) ^ (inputs[185]);
    assign layer0_outputs[3495] = inputs[26];
    assign layer0_outputs[3496] = ~((inputs[237]) | (inputs[14]));
    assign layer0_outputs[3497] = (inputs[212]) | (inputs[232]);
    assign layer0_outputs[3498] = ~((inputs[170]) | (inputs[30]));
    assign layer0_outputs[3499] = ~(inputs[223]);
    assign layer0_outputs[3500] = ~((inputs[181]) ^ (inputs[158]));
    assign layer0_outputs[3501] = (inputs[8]) ^ (inputs[109]);
    assign layer0_outputs[3502] = ~(inputs[137]) | (inputs[84]);
    assign layer0_outputs[3503] = (inputs[177]) | (inputs[248]);
    assign layer0_outputs[3504] = ~((inputs[57]) ^ (inputs[76]));
    assign layer0_outputs[3505] = inputs[31];
    assign layer0_outputs[3506] = ~((inputs[53]) ^ (inputs[88]));
    assign layer0_outputs[3507] = ~(inputs[144]);
    assign layer0_outputs[3508] = ~((inputs[217]) | (inputs[38]));
    assign layer0_outputs[3509] = ~(inputs[179]) | (inputs[58]);
    assign layer0_outputs[3510] = (inputs[0]) | (inputs[255]);
    assign layer0_outputs[3511] = (inputs[1]) & ~(inputs[140]);
    assign layer0_outputs[3512] = (inputs[119]) & (inputs[25]);
    assign layer0_outputs[3513] = (inputs[149]) & ~(inputs[201]);
    assign layer0_outputs[3514] = inputs[37];
    assign layer0_outputs[3515] = inputs[182];
    assign layer0_outputs[3516] = (inputs[30]) ^ (inputs[106]);
    assign layer0_outputs[3517] = (inputs[235]) ^ (inputs[16]);
    assign layer0_outputs[3518] = ~((inputs[135]) & (inputs[149]));
    assign layer0_outputs[3519] = inputs[171];
    assign layer0_outputs[3520] = inputs[116];
    assign layer0_outputs[3521] = ~((inputs[59]) | (inputs[135]));
    assign layer0_outputs[3522] = (inputs[89]) | (inputs[6]);
    assign layer0_outputs[3523] = inputs[164];
    assign layer0_outputs[3524] = inputs[164];
    assign layer0_outputs[3525] = (inputs[72]) ^ (inputs[117]);
    assign layer0_outputs[3526] = ~((inputs[38]) & (inputs[214]));
    assign layer0_outputs[3527] = ~(inputs[98]);
    assign layer0_outputs[3528] = (inputs[0]) ^ (inputs[196]);
    assign layer0_outputs[3529] = ~((inputs[29]) | (inputs[71]));
    assign layer0_outputs[3530] = inputs[93];
    assign layer0_outputs[3531] = (inputs[182]) ^ (inputs[212]);
    assign layer0_outputs[3532] = (inputs[196]) ^ (inputs[38]);
    assign layer0_outputs[3533] = inputs[67];
    assign layer0_outputs[3534] = (inputs[159]) ^ (inputs[218]);
    assign layer0_outputs[3535] = inputs[1];
    assign layer0_outputs[3536] = (inputs[44]) | (inputs[65]);
    assign layer0_outputs[3537] = inputs[2];
    assign layer0_outputs[3538] = ~((inputs[194]) | (inputs[208]));
    assign layer0_outputs[3539] = 1'b0;
    assign layer0_outputs[3540] = inputs[150];
    assign layer0_outputs[3541] = ~(inputs[189]);
    assign layer0_outputs[3542] = ~((inputs[18]) | (inputs[182]));
    assign layer0_outputs[3543] = ~(inputs[75]);
    assign layer0_outputs[3544] = (inputs[22]) & ~(inputs[253]);
    assign layer0_outputs[3545] = (inputs[89]) & ~(inputs[201]);
    assign layer0_outputs[3546] = ~((inputs[168]) | (inputs[242]));
    assign layer0_outputs[3547] = ~((inputs[171]) | (inputs[149]));
    assign layer0_outputs[3548] = ~(inputs[250]);
    assign layer0_outputs[3549] = ~((inputs[5]) | (inputs[26]));
    assign layer0_outputs[3550] = (inputs[14]) | (inputs[47]);
    assign layer0_outputs[3551] = (inputs[118]) | (inputs[203]);
    assign layer0_outputs[3552] = inputs[4];
    assign layer0_outputs[3553] = (inputs[57]) & ~(inputs[239]);
    assign layer0_outputs[3554] = (inputs[28]) | (inputs[116]);
    assign layer0_outputs[3555] = ~(inputs[210]) | (inputs[255]);
    assign layer0_outputs[3556] = ~((inputs[113]) | (inputs[192]));
    assign layer0_outputs[3557] = ~((inputs[31]) | (inputs[27]));
    assign layer0_outputs[3558] = (inputs[41]) | (inputs[111]);
    assign layer0_outputs[3559] = ~(inputs[243]) | (inputs[81]);
    assign layer0_outputs[3560] = (inputs[35]) ^ (inputs[24]);
    assign layer0_outputs[3561] = ~(inputs[197]);
    assign layer0_outputs[3562] = ~((inputs[75]) | (inputs[15]));
    assign layer0_outputs[3563] = ~((inputs[52]) | (inputs[101]));
    assign layer0_outputs[3564] = ~(inputs[150]);
    assign layer0_outputs[3565] = (inputs[238]) | (inputs[192]);
    assign layer0_outputs[3566] = ~((inputs[138]) ^ (inputs[152]));
    assign layer0_outputs[3567] = (inputs[183]) & (inputs[198]);
    assign layer0_outputs[3568] = (inputs[246]) & ~(inputs[126]);
    assign layer0_outputs[3569] = ~(inputs[139]) | (inputs[74]);
    assign layer0_outputs[3570] = (inputs[209]) & ~(inputs[208]);
    assign layer0_outputs[3571] = 1'b0;
    assign layer0_outputs[3572] = (inputs[189]) & ~(inputs[221]);
    assign layer0_outputs[3573] = ~(inputs[142]) | (inputs[109]);
    assign layer0_outputs[3574] = (inputs[62]) & ~(inputs[241]);
    assign layer0_outputs[3575] = ~((inputs[235]) & (inputs[107]));
    assign layer0_outputs[3576] = ~((inputs[64]) ^ (inputs[174]));
    assign layer0_outputs[3577] = (inputs[186]) ^ (inputs[197]);
    assign layer0_outputs[3578] = (inputs[69]) & ~(inputs[202]);
    assign layer0_outputs[3579] = ~((inputs[201]) ^ (inputs[89]));
    assign layer0_outputs[3580] = 1'b1;
    assign layer0_outputs[3581] = ~(inputs[6]);
    assign layer0_outputs[3582] = ~((inputs[73]) | (inputs[45]));
    assign layer0_outputs[3583] = ~((inputs[1]) ^ (inputs[105]));
    assign layer0_outputs[3584] = ~(inputs[77]) | (inputs[201]);
    assign layer0_outputs[3585] = (inputs[125]) | (inputs[37]);
    assign layer0_outputs[3586] = (inputs[243]) | (inputs[240]);
    assign layer0_outputs[3587] = inputs[23];
    assign layer0_outputs[3588] = (inputs[111]) | (inputs[182]);
    assign layer0_outputs[3589] = ~(inputs[186]) | (inputs[91]);
    assign layer0_outputs[3590] = 1'b0;
    assign layer0_outputs[3591] = (inputs[197]) & ~(inputs[241]);
    assign layer0_outputs[3592] = ~(inputs[175]);
    assign layer0_outputs[3593] = ~((inputs[217]) | (inputs[163]));
    assign layer0_outputs[3594] = (inputs[76]) & (inputs[120]);
    assign layer0_outputs[3595] = inputs[101];
    assign layer0_outputs[3596] = (inputs[193]) ^ (inputs[181]);
    assign layer0_outputs[3597] = ~(inputs[209]);
    assign layer0_outputs[3598] = inputs[105];
    assign layer0_outputs[3599] = ~(inputs[149]) | (inputs[152]);
    assign layer0_outputs[3600] = (inputs[107]) | (inputs[52]);
    assign layer0_outputs[3601] = (inputs[254]) | (inputs[131]);
    assign layer0_outputs[3602] = (inputs[13]) ^ (inputs[209]);
    assign layer0_outputs[3603] = (inputs[168]) & ~(inputs[27]);
    assign layer0_outputs[3604] = ~(inputs[110]);
    assign layer0_outputs[3605] = ~(inputs[134]) | (inputs[204]);
    assign layer0_outputs[3606] = (inputs[232]) & ~(inputs[115]);
    assign layer0_outputs[3607] = ~(inputs[41]);
    assign layer0_outputs[3608] = ~(inputs[21]);
    assign layer0_outputs[3609] = (inputs[234]) | (inputs[16]);
    assign layer0_outputs[3610] = (inputs[241]) | (inputs[35]);
    assign layer0_outputs[3611] = ~(inputs[70]);
    assign layer0_outputs[3612] = ~(inputs[167]) | (inputs[41]);
    assign layer0_outputs[3613] = (inputs[58]) & ~(inputs[251]);
    assign layer0_outputs[3614] = inputs[234];
    assign layer0_outputs[3615] = inputs[167];
    assign layer0_outputs[3616] = 1'b0;
    assign layer0_outputs[3617] = (inputs[164]) ^ (inputs[111]);
    assign layer0_outputs[3618] = (inputs[9]) | (inputs[63]);
    assign layer0_outputs[3619] = 1'b1;
    assign layer0_outputs[3620] = inputs[134];
    assign layer0_outputs[3621] = (inputs[193]) & ~(inputs[26]);
    assign layer0_outputs[3622] = ~(inputs[252]) | (inputs[64]);
    assign layer0_outputs[3623] = ~((inputs[116]) ^ (inputs[16]));
    assign layer0_outputs[3624] = ~(inputs[243]);
    assign layer0_outputs[3625] = ~(inputs[151]);
    assign layer0_outputs[3626] = inputs[121];
    assign layer0_outputs[3627] = ~((inputs[115]) ^ (inputs[243]));
    assign layer0_outputs[3628] = 1'b1;
    assign layer0_outputs[3629] = (inputs[189]) | (inputs[213]);
    assign layer0_outputs[3630] = ~(inputs[52]) | (inputs[176]);
    assign layer0_outputs[3631] = inputs[146];
    assign layer0_outputs[3632] = ~(inputs[152]);
    assign layer0_outputs[3633] = ~((inputs[174]) & (inputs[189]));
    assign layer0_outputs[3634] = inputs[248];
    assign layer0_outputs[3635] = inputs[150];
    assign layer0_outputs[3636] = (inputs[34]) ^ (inputs[143]);
    assign layer0_outputs[3637] = ~((inputs[76]) | (inputs[105]));
    assign layer0_outputs[3638] = (inputs[33]) | (inputs[219]);
    assign layer0_outputs[3639] = ~(inputs[25]);
    assign layer0_outputs[3640] = (inputs[134]) & ~(inputs[166]);
    assign layer0_outputs[3641] = ~(inputs[19]);
    assign layer0_outputs[3642] = ~((inputs[219]) | (inputs[173]));
    assign layer0_outputs[3643] = ~((inputs[147]) | (inputs[8]));
    assign layer0_outputs[3644] = 1'b0;
    assign layer0_outputs[3645] = (inputs[6]) | (inputs[222]);
    assign layer0_outputs[3646] = (inputs[33]) & ~(inputs[112]);
    assign layer0_outputs[3647] = ~(inputs[17]);
    assign layer0_outputs[3648] = (inputs[27]) & ~(inputs[172]);
    assign layer0_outputs[3649] = ~((inputs[168]) ^ (inputs[242]));
    assign layer0_outputs[3650] = (inputs[123]) & ~(inputs[207]);
    assign layer0_outputs[3651] = (inputs[48]) | (inputs[235]);
    assign layer0_outputs[3652] = inputs[30];
    assign layer0_outputs[3653] = (inputs[103]) & ~(inputs[157]);
    assign layer0_outputs[3654] = (inputs[85]) & ~(inputs[56]);
    assign layer0_outputs[3655] = ~(inputs[253]) | (inputs[78]);
    assign layer0_outputs[3656] = (inputs[209]) & ~(inputs[121]);
    assign layer0_outputs[3657] = (inputs[212]) | (inputs[132]);
    assign layer0_outputs[3658] = (inputs[156]) | (inputs[62]);
    assign layer0_outputs[3659] = ~((inputs[181]) ^ (inputs[229]));
    assign layer0_outputs[3660] = ~((inputs[58]) | (inputs[62]));
    assign layer0_outputs[3661] = ~(inputs[164]) | (inputs[36]);
    assign layer0_outputs[3662] = ~((inputs[48]) | (inputs[1]));
    assign layer0_outputs[3663] = 1'b0;
    assign layer0_outputs[3664] = (inputs[222]) ^ (inputs[2]);
    assign layer0_outputs[3665] = (inputs[190]) ^ (inputs[242]);
    assign layer0_outputs[3666] = ~(inputs[176]);
    assign layer0_outputs[3667] = (inputs[47]) & ~(inputs[236]);
    assign layer0_outputs[3668] = inputs[182];
    assign layer0_outputs[3669] = inputs[84];
    assign layer0_outputs[3670] = (inputs[50]) & ~(inputs[236]);
    assign layer0_outputs[3671] = (inputs[203]) & (inputs[152]);
    assign layer0_outputs[3672] = ~((inputs[160]) | (inputs[214]));
    assign layer0_outputs[3673] = (inputs[122]) & ~(inputs[214]);
    assign layer0_outputs[3674] = inputs[175];
    assign layer0_outputs[3675] = ~(inputs[185]);
    assign layer0_outputs[3676] = (inputs[23]) | (inputs[190]);
    assign layer0_outputs[3677] = ~(inputs[13]);
    assign layer0_outputs[3678] = ~((inputs[176]) | (inputs[164]));
    assign layer0_outputs[3679] = ~(inputs[105]);
    assign layer0_outputs[3680] = (inputs[219]) & ~(inputs[207]);
    assign layer0_outputs[3681] = inputs[232];
    assign layer0_outputs[3682] = ~((inputs[177]) | (inputs[55]));
    assign layer0_outputs[3683] = ~(inputs[9]);
    assign layer0_outputs[3684] = ~((inputs[210]) ^ (inputs[174]));
    assign layer0_outputs[3685] = ~((inputs[169]) | (inputs[254]));
    assign layer0_outputs[3686] = ~(inputs[85]);
    assign layer0_outputs[3687] = (inputs[171]) | (inputs[217]);
    assign layer0_outputs[3688] = (inputs[186]) | (inputs[203]);
    assign layer0_outputs[3689] = ~(inputs[184]);
    assign layer0_outputs[3690] = ~((inputs[72]) ^ (inputs[51]));
    assign layer0_outputs[3691] = ~((inputs[240]) ^ (inputs[127]));
    assign layer0_outputs[3692] = ~(inputs[153]) | (inputs[225]);
    assign layer0_outputs[3693] = ~((inputs[25]) | (inputs[17]));
    assign layer0_outputs[3694] = ~((inputs[254]) ^ (inputs[21]));
    assign layer0_outputs[3695] = ~(inputs[193]);
    assign layer0_outputs[3696] = ~(inputs[231]) | (inputs[90]);
    assign layer0_outputs[3697] = inputs[156];
    assign layer0_outputs[3698] = (inputs[197]) & ~(inputs[28]);
    assign layer0_outputs[3699] = (inputs[98]) & ~(inputs[191]);
    assign layer0_outputs[3700] = ~(inputs[124]);
    assign layer0_outputs[3701] = (inputs[219]) | (inputs[6]);
    assign layer0_outputs[3702] = ~(inputs[102]);
    assign layer0_outputs[3703] = inputs[161];
    assign layer0_outputs[3704] = ~((inputs[140]) ^ (inputs[154]));
    assign layer0_outputs[3705] = inputs[154];
    assign layer0_outputs[3706] = ~((inputs[212]) | (inputs[186]));
    assign layer0_outputs[3707] = ~(inputs[155]) | (inputs[163]);
    assign layer0_outputs[3708] = inputs[61];
    assign layer0_outputs[3709] = inputs[81];
    assign layer0_outputs[3710] = ~(inputs[82]);
    assign layer0_outputs[3711] = (inputs[196]) | (inputs[182]);
    assign layer0_outputs[3712] = (inputs[139]) | (inputs[158]);
    assign layer0_outputs[3713] = ~(inputs[248]);
    assign layer0_outputs[3714] = (inputs[229]) & ~(inputs[3]);
    assign layer0_outputs[3715] = (inputs[206]) ^ (inputs[127]);
    assign layer0_outputs[3716] = ~(inputs[183]) | (inputs[225]);
    assign layer0_outputs[3717] = ~((inputs[34]) & (inputs[142]));
    assign layer0_outputs[3718] = (inputs[85]) & (inputs[85]);
    assign layer0_outputs[3719] = ~(inputs[167]);
    assign layer0_outputs[3720] = ~(inputs[68]);
    assign layer0_outputs[3721] = ~(inputs[125]);
    assign layer0_outputs[3722] = ~(inputs[43]) | (inputs[234]);
    assign layer0_outputs[3723] = (inputs[168]) & (inputs[247]);
    assign layer0_outputs[3724] = (inputs[3]) & ~(inputs[252]);
    assign layer0_outputs[3725] = ~(inputs[9]);
    assign layer0_outputs[3726] = (inputs[160]) ^ (inputs[81]);
    assign layer0_outputs[3727] = ~(inputs[25]);
    assign layer0_outputs[3728] = ~((inputs[65]) | (inputs[7]));
    assign layer0_outputs[3729] = (inputs[20]) ^ (inputs[177]);
    assign layer0_outputs[3730] = (inputs[49]) | (inputs[199]);
    assign layer0_outputs[3731] = (inputs[196]) & ~(inputs[191]);
    assign layer0_outputs[3732] = (inputs[246]) | (inputs[213]);
    assign layer0_outputs[3733] = ~((inputs[9]) ^ (inputs[161]));
    assign layer0_outputs[3734] = (inputs[112]) | (inputs[248]);
    assign layer0_outputs[3735] = (inputs[56]) & (inputs[108]);
    assign layer0_outputs[3736] = (inputs[185]) | (inputs[123]);
    assign layer0_outputs[3737] = (inputs[194]) | (inputs[247]);
    assign layer0_outputs[3738] = (inputs[216]) & ~(inputs[246]);
    assign layer0_outputs[3739] = ~(inputs[44]) | (inputs[252]);
    assign layer0_outputs[3740] = inputs[236];
    assign layer0_outputs[3741] = ~((inputs[254]) | (inputs[62]));
    assign layer0_outputs[3742] = (inputs[138]) ^ (inputs[216]);
    assign layer0_outputs[3743] = ~(inputs[60]) | (inputs[81]);
    assign layer0_outputs[3744] = ~(inputs[112]);
    assign layer0_outputs[3745] = inputs[228];
    assign layer0_outputs[3746] = inputs[15];
    assign layer0_outputs[3747] = ~(inputs[217]);
    assign layer0_outputs[3748] = (inputs[14]) ^ (inputs[126]);
    assign layer0_outputs[3749] = ~(inputs[250]);
    assign layer0_outputs[3750] = ~(inputs[103]);
    assign layer0_outputs[3751] = inputs[129];
    assign layer0_outputs[3752] = (inputs[41]) & ~(inputs[66]);
    assign layer0_outputs[3753] = inputs[2];
    assign layer0_outputs[3754] = (inputs[233]) & ~(inputs[39]);
    assign layer0_outputs[3755] = ~((inputs[38]) | (inputs[21]));
    assign layer0_outputs[3756] = (inputs[149]) & ~(inputs[74]);
    assign layer0_outputs[3757] = ~(inputs[115]) | (inputs[206]);
    assign layer0_outputs[3758] = (inputs[38]) & ~(inputs[145]);
    assign layer0_outputs[3759] = (inputs[28]) & ~(inputs[205]);
    assign layer0_outputs[3760] = ~((inputs[62]) ^ (inputs[24]));
    assign layer0_outputs[3761] = ~((inputs[124]) ^ (inputs[254]));
    assign layer0_outputs[3762] = ~((inputs[162]) | (inputs[191]));
    assign layer0_outputs[3763] = (inputs[64]) | (inputs[174]);
    assign layer0_outputs[3764] = (inputs[229]) & ~(inputs[15]);
    assign layer0_outputs[3765] = ~((inputs[181]) | (inputs[79]));
    assign layer0_outputs[3766] = ~(inputs[49]);
    assign layer0_outputs[3767] = inputs[120];
    assign layer0_outputs[3768] = (inputs[195]) & ~(inputs[12]);
    assign layer0_outputs[3769] = ~((inputs[211]) ^ (inputs[157]));
    assign layer0_outputs[3770] = inputs[168];
    assign layer0_outputs[3771] = ~(inputs[44]);
    assign layer0_outputs[3772] = ~((inputs[255]) | (inputs[49]));
    assign layer0_outputs[3773] = ~((inputs[66]) ^ (inputs[101]));
    assign layer0_outputs[3774] = ~((inputs[179]) | (inputs[98]));
    assign layer0_outputs[3775] = (inputs[175]) | (inputs[79]);
    assign layer0_outputs[3776] = inputs[88];
    assign layer0_outputs[3777] = ~(inputs[102]);
    assign layer0_outputs[3778] = inputs[165];
    assign layer0_outputs[3779] = (inputs[58]) & ~(inputs[47]);
    assign layer0_outputs[3780] = ~(inputs[101]);
    assign layer0_outputs[3781] = ~((inputs[239]) | (inputs[117]));
    assign layer0_outputs[3782] = (inputs[111]) | (inputs[214]);
    assign layer0_outputs[3783] = ~((inputs[198]) | (inputs[243]));
    assign layer0_outputs[3784] = 1'b1;
    assign layer0_outputs[3785] = (inputs[219]) | (inputs[238]);
    assign layer0_outputs[3786] = ~(inputs[101]) | (inputs[6]);
    assign layer0_outputs[3787] = (inputs[56]) | (inputs[209]);
    assign layer0_outputs[3788] = ~(inputs[249]);
    assign layer0_outputs[3789] = inputs[118];
    assign layer0_outputs[3790] = (inputs[209]) | (inputs[217]);
    assign layer0_outputs[3791] = ~((inputs[12]) | (inputs[246]));
    assign layer0_outputs[3792] = ~((inputs[103]) | (inputs[62]));
    assign layer0_outputs[3793] = (inputs[182]) & ~(inputs[143]);
    assign layer0_outputs[3794] = ~(inputs[166]);
    assign layer0_outputs[3795] = 1'b0;
    assign layer0_outputs[3796] = ~((inputs[137]) ^ (inputs[151]));
    assign layer0_outputs[3797] = inputs[204];
    assign layer0_outputs[3798] = inputs[144];
    assign layer0_outputs[3799] = inputs[24];
    assign layer0_outputs[3800] = (inputs[154]) & (inputs[254]);
    assign layer0_outputs[3801] = (inputs[106]) & (inputs[26]);
    assign layer0_outputs[3802] = (inputs[240]) | (inputs[29]);
    assign layer0_outputs[3803] = inputs[86];
    assign layer0_outputs[3804] = (inputs[21]) ^ (inputs[80]);
    assign layer0_outputs[3805] = ~(inputs[186]) | (inputs[168]);
    assign layer0_outputs[3806] = (inputs[58]) | (inputs[194]);
    assign layer0_outputs[3807] = ~(inputs[213]);
    assign layer0_outputs[3808] = (inputs[167]) & ~(inputs[235]);
    assign layer0_outputs[3809] = inputs[107];
    assign layer0_outputs[3810] = ~(inputs[3]) | (inputs[81]);
    assign layer0_outputs[3811] = inputs[142];
    assign layer0_outputs[3812] = 1'b1;
    assign layer0_outputs[3813] = inputs[134];
    assign layer0_outputs[3814] = ~(inputs[98]) | (inputs[169]);
    assign layer0_outputs[3815] = ~(inputs[221]) | (inputs[12]);
    assign layer0_outputs[3816] = inputs[99];
    assign layer0_outputs[3817] = ~((inputs[101]) ^ (inputs[152]));
    assign layer0_outputs[3818] = ~(inputs[75]) | (inputs[112]);
    assign layer0_outputs[3819] = ~(inputs[235]);
    assign layer0_outputs[3820] = ~((inputs[237]) ^ (inputs[64]));
    assign layer0_outputs[3821] = ~(inputs[95]);
    assign layer0_outputs[3822] = (inputs[159]) ^ (inputs[34]);
    assign layer0_outputs[3823] = ~(inputs[156]) | (inputs[137]);
    assign layer0_outputs[3824] = ~((inputs[210]) & (inputs[171]));
    assign layer0_outputs[3825] = ~((inputs[107]) & (inputs[73]));
    assign layer0_outputs[3826] = ~((inputs[234]) | (inputs[143]));
    assign layer0_outputs[3827] = (inputs[93]) & ~(inputs[229]);
    assign layer0_outputs[3828] = inputs[25];
    assign layer0_outputs[3829] = ~(inputs[130]);
    assign layer0_outputs[3830] = ~((inputs[144]) | (inputs[23]));
    assign layer0_outputs[3831] = ~((inputs[51]) ^ (inputs[119]));
    assign layer0_outputs[3832] = (inputs[74]) ^ (inputs[2]);
    assign layer0_outputs[3833] = (inputs[208]) & ~(inputs[162]);
    assign layer0_outputs[3834] = inputs[168];
    assign layer0_outputs[3835] = (inputs[109]) & ~(inputs[137]);
    assign layer0_outputs[3836] = ~(inputs[248]) | (inputs[52]);
    assign layer0_outputs[3837] = inputs[40];
    assign layer0_outputs[3838] = ~(inputs[193]);
    assign layer0_outputs[3839] = (inputs[203]) | (inputs[207]);
    assign layer0_outputs[3840] = ~((inputs[40]) ^ (inputs[70]));
    assign layer0_outputs[3841] = ~((inputs[243]) & (inputs[241]));
    assign layer0_outputs[3842] = ~(inputs[219]) | (inputs[102]);
    assign layer0_outputs[3843] = (inputs[21]) & ~(inputs[157]);
    assign layer0_outputs[3844] = (inputs[142]) & ~(inputs[171]);
    assign layer0_outputs[3845] = (inputs[6]) & ~(inputs[33]);
    assign layer0_outputs[3846] = ~((inputs[255]) | (inputs[169]));
    assign layer0_outputs[3847] = ~((inputs[55]) | (inputs[223]));
    assign layer0_outputs[3848] = ~((inputs[221]) ^ (inputs[236]));
    assign layer0_outputs[3849] = ~((inputs[21]) ^ (inputs[150]));
    assign layer0_outputs[3850] = (inputs[24]) & ~(inputs[225]);
    assign layer0_outputs[3851] = ~((inputs[244]) | (inputs[26]));
    assign layer0_outputs[3852] = (inputs[43]) & ~(inputs[19]);
    assign layer0_outputs[3853] = ~(inputs[147]);
    assign layer0_outputs[3854] = ~((inputs[15]) | (inputs[169]));
    assign layer0_outputs[3855] = ~(inputs[87]);
    assign layer0_outputs[3856] = ~(inputs[248]) | (inputs[87]);
    assign layer0_outputs[3857] = inputs[122];
    assign layer0_outputs[3858] = inputs[90];
    assign layer0_outputs[3859] = ~((inputs[128]) ^ (inputs[22]));
    assign layer0_outputs[3860] = ~(inputs[116]) | (inputs[55]);
    assign layer0_outputs[3861] = ~(inputs[94]);
    assign layer0_outputs[3862] = (inputs[218]) & ~(inputs[32]);
    assign layer0_outputs[3863] = ~(inputs[115]);
    assign layer0_outputs[3864] = ~(inputs[247]) | (inputs[36]);
    assign layer0_outputs[3865] = inputs[194];
    assign layer0_outputs[3866] = ~((inputs[51]) ^ (inputs[207]));
    assign layer0_outputs[3867] = (inputs[150]) ^ (inputs[213]);
    assign layer0_outputs[3868] = (inputs[203]) & ~(inputs[7]);
    assign layer0_outputs[3869] = (inputs[147]) | (inputs[102]);
    assign layer0_outputs[3870] = inputs[0];
    assign layer0_outputs[3871] = ~((inputs[234]) ^ (inputs[161]));
    assign layer0_outputs[3872] = (inputs[92]) & ~(inputs[239]);
    assign layer0_outputs[3873] = (inputs[134]) & (inputs[60]);
    assign layer0_outputs[3874] = ~((inputs[206]) | (inputs[203]));
    assign layer0_outputs[3875] = ~((inputs[124]) ^ (inputs[89]));
    assign layer0_outputs[3876] = ~((inputs[71]) ^ (inputs[254]));
    assign layer0_outputs[3877] = ~((inputs[67]) & (inputs[8]));
    assign layer0_outputs[3878] = inputs[50];
    assign layer0_outputs[3879] = 1'b1;
    assign layer0_outputs[3880] = (inputs[128]) ^ (inputs[172]);
    assign layer0_outputs[3881] = ~((inputs[84]) ^ (inputs[9]));
    assign layer0_outputs[3882] = ~(inputs[137]);
    assign layer0_outputs[3883] = (inputs[152]) & (inputs[74]);
    assign layer0_outputs[3884] = ~((inputs[110]) ^ (inputs[221]));
    assign layer0_outputs[3885] = ~(inputs[233]);
    assign layer0_outputs[3886] = (inputs[93]) | (inputs[51]);
    assign layer0_outputs[3887] = inputs[19];
    assign layer0_outputs[3888] = ~(inputs[163]);
    assign layer0_outputs[3889] = inputs[75];
    assign layer0_outputs[3890] = ~((inputs[131]) | (inputs[203]));
    assign layer0_outputs[3891] = (inputs[205]) | (inputs[252]);
    assign layer0_outputs[3892] = (inputs[67]) | (inputs[185]);
    assign layer0_outputs[3893] = ~(inputs[230]) | (inputs[33]);
    assign layer0_outputs[3894] = ~((inputs[213]) & (inputs[202]));
    assign layer0_outputs[3895] = ~(inputs[8]);
    assign layer0_outputs[3896] = inputs[211];
    assign layer0_outputs[3897] = ~((inputs[52]) | (inputs[37]));
    assign layer0_outputs[3898] = (inputs[92]) & ~(inputs[238]);
    assign layer0_outputs[3899] = inputs[110];
    assign layer0_outputs[3900] = ~(inputs[130]);
    assign layer0_outputs[3901] = ~(inputs[232]) | (inputs[14]);
    assign layer0_outputs[3902] = ~(inputs[68]) | (inputs[16]);
    assign layer0_outputs[3903] = ~((inputs[135]) | (inputs[199]));
    assign layer0_outputs[3904] = ~(inputs[121]);
    assign layer0_outputs[3905] = ~(inputs[102]);
    assign layer0_outputs[3906] = ~(inputs[128]) | (inputs[238]);
    assign layer0_outputs[3907] = inputs[221];
    assign layer0_outputs[3908] = (inputs[171]) ^ (inputs[135]);
    assign layer0_outputs[3909] = (inputs[141]) ^ (inputs[108]);
    assign layer0_outputs[3910] = (inputs[21]) ^ (inputs[175]);
    assign layer0_outputs[3911] = inputs[55];
    assign layer0_outputs[3912] = (inputs[95]) ^ (inputs[135]);
    assign layer0_outputs[3913] = (inputs[130]) | (inputs[34]);
    assign layer0_outputs[3914] = (inputs[91]) & ~(inputs[119]);
    assign layer0_outputs[3915] = ~(inputs[124]);
    assign layer0_outputs[3916] = inputs[224];
    assign layer0_outputs[3917] = (inputs[218]) | (inputs[216]);
    assign layer0_outputs[3918] = inputs[106];
    assign layer0_outputs[3919] = ~((inputs[116]) ^ (inputs[188]));
    assign layer0_outputs[3920] = ~(inputs[19]);
    assign layer0_outputs[3921] = (inputs[194]) & (inputs[138]);
    assign layer0_outputs[3922] = inputs[249];
    assign layer0_outputs[3923] = inputs[166];
    assign layer0_outputs[3924] = (inputs[12]) & ~(inputs[109]);
    assign layer0_outputs[3925] = ~(inputs[103]);
    assign layer0_outputs[3926] = inputs[147];
    assign layer0_outputs[3927] = ~(inputs[69]) | (inputs[116]);
    assign layer0_outputs[3928] = inputs[19];
    assign layer0_outputs[3929] = ~((inputs[196]) | (inputs[166]));
    assign layer0_outputs[3930] = 1'b1;
    assign layer0_outputs[3931] = (inputs[135]) & (inputs[199]);
    assign layer0_outputs[3932] = inputs[52];
    assign layer0_outputs[3933] = ~(inputs[28]) | (inputs[207]);
    assign layer0_outputs[3934] = (inputs[135]) & ~(inputs[185]);
    assign layer0_outputs[3935] = ~(inputs[220]);
    assign layer0_outputs[3936] = (inputs[110]) ^ (inputs[32]);
    assign layer0_outputs[3937] = ~((inputs[226]) | (inputs[146]));
    assign layer0_outputs[3938] = inputs[56];
    assign layer0_outputs[3939] = (inputs[237]) | (inputs[150]);
    assign layer0_outputs[3940] = ~((inputs[122]) | (inputs[163]));
    assign layer0_outputs[3941] = (inputs[95]) & (inputs[37]);
    assign layer0_outputs[3942] = inputs[194];
    assign layer0_outputs[3943] = ~((inputs[65]) ^ (inputs[70]));
    assign layer0_outputs[3944] = (inputs[19]) | (inputs[73]);
    assign layer0_outputs[3945] = (inputs[59]) | (inputs[67]);
    assign layer0_outputs[3946] = ~((inputs[93]) | (inputs[4]));
    assign layer0_outputs[3947] = inputs[52];
    assign layer0_outputs[3948] = ~((inputs[175]) | (inputs[2]));
    assign layer0_outputs[3949] = inputs[63];
    assign layer0_outputs[3950] = (inputs[0]) | (inputs[71]);
    assign layer0_outputs[3951] = inputs[182];
    assign layer0_outputs[3952] = (inputs[16]) | (inputs[173]);
    assign layer0_outputs[3953] = inputs[155];
    assign layer0_outputs[3954] = ~(inputs[61]) | (inputs[149]);
    assign layer0_outputs[3955] = (inputs[100]) | (inputs[141]);
    assign layer0_outputs[3956] = (inputs[39]) | (inputs[221]);
    assign layer0_outputs[3957] = inputs[219];
    assign layer0_outputs[3958] = inputs[225];
    assign layer0_outputs[3959] = ~((inputs[213]) | (inputs[24]));
    assign layer0_outputs[3960] = (inputs[9]) & ~(inputs[128]);
    assign layer0_outputs[3961] = ~(inputs[149]) | (inputs[143]);
    assign layer0_outputs[3962] = (inputs[41]) & ~(inputs[194]);
    assign layer0_outputs[3963] = ~(inputs[174]);
    assign layer0_outputs[3964] = 1'b0;
    assign layer0_outputs[3965] = ~(inputs[168]) | (inputs[241]);
    assign layer0_outputs[3966] = inputs[85];
    assign layer0_outputs[3967] = (inputs[59]) & ~(inputs[193]);
    assign layer0_outputs[3968] = (inputs[22]) | (inputs[55]);
    assign layer0_outputs[3969] = (inputs[164]) ^ (inputs[203]);
    assign layer0_outputs[3970] = 1'b0;
    assign layer0_outputs[3971] = inputs[125];
    assign layer0_outputs[3972] = (inputs[161]) | (inputs[146]);
    assign layer0_outputs[3973] = ~(inputs[178]);
    assign layer0_outputs[3974] = ~(inputs[69]) | (inputs[161]);
    assign layer0_outputs[3975] = (inputs[217]) & ~(inputs[34]);
    assign layer0_outputs[3976] = (inputs[254]) | (inputs[224]);
    assign layer0_outputs[3977] = ~((inputs[24]) | (inputs[33]));
    assign layer0_outputs[3978] = inputs[106];
    assign layer0_outputs[3979] = ~((inputs[238]) | (inputs[109]));
    assign layer0_outputs[3980] = ~((inputs[67]) | (inputs[174]));
    assign layer0_outputs[3981] = ~((inputs[26]) ^ (inputs[60]));
    assign layer0_outputs[3982] = ~((inputs[159]) | (inputs[199]));
    assign layer0_outputs[3983] = inputs[213];
    assign layer0_outputs[3984] = ~((inputs[131]) ^ (inputs[175]));
    assign layer0_outputs[3985] = inputs[173];
    assign layer0_outputs[3986] = (inputs[234]) | (inputs[232]);
    assign layer0_outputs[3987] = ~(inputs[24]);
    assign layer0_outputs[3988] = (inputs[104]) & (inputs[166]);
    assign layer0_outputs[3989] = inputs[39];
    assign layer0_outputs[3990] = ~((inputs[37]) ^ (inputs[0]));
    assign layer0_outputs[3991] = ~(inputs[117]) | (inputs[50]);
    assign layer0_outputs[3992] = (inputs[98]) | (inputs[28]);
    assign layer0_outputs[3993] = inputs[25];
    assign layer0_outputs[3994] = (inputs[6]) & ~(inputs[159]);
    assign layer0_outputs[3995] = (inputs[12]) & (inputs[69]);
    assign layer0_outputs[3996] = (inputs[55]) & ~(inputs[255]);
    assign layer0_outputs[3997] = ~(inputs[74]) | (inputs[169]);
    assign layer0_outputs[3998] = (inputs[131]) ^ (inputs[165]);
    assign layer0_outputs[3999] = inputs[93];
    assign layer0_outputs[4000] = ~((inputs[244]) & (inputs[178]));
    assign layer0_outputs[4001] = ~((inputs[41]) ^ (inputs[234]));
    assign layer0_outputs[4002] = ~((inputs[74]) & (inputs[205]));
    assign layer0_outputs[4003] = ~(inputs[169]);
    assign layer0_outputs[4004] = inputs[99];
    assign layer0_outputs[4005] = ~(inputs[87]);
    assign layer0_outputs[4006] = ~(inputs[115]) | (inputs[46]);
    assign layer0_outputs[4007] = ~((inputs[48]) | (inputs[186]));
    assign layer0_outputs[4008] = (inputs[7]) | (inputs[83]);
    assign layer0_outputs[4009] = (inputs[26]) & ~(inputs[147]);
    assign layer0_outputs[4010] = inputs[211];
    assign layer0_outputs[4011] = inputs[91];
    assign layer0_outputs[4012] = ~(inputs[80]);
    assign layer0_outputs[4013] = ~((inputs[12]) | (inputs[62]));
    assign layer0_outputs[4014] = ~((inputs[231]) | (inputs[191]));
    assign layer0_outputs[4015] = ~((inputs[143]) ^ (inputs[180]));
    assign layer0_outputs[4016] = 1'b1;
    assign layer0_outputs[4017] = ~((inputs[209]) | (inputs[82]));
    assign layer0_outputs[4018] = inputs[223];
    assign layer0_outputs[4019] = ~(inputs[44]);
    assign layer0_outputs[4020] = (inputs[186]) | (inputs[19]);
    assign layer0_outputs[4021] = inputs[46];
    assign layer0_outputs[4022] = inputs[100];
    assign layer0_outputs[4023] = (inputs[53]) & ~(inputs[250]);
    assign layer0_outputs[4024] = ~((inputs[22]) | (inputs[246]));
    assign layer0_outputs[4025] = inputs[98];
    assign layer0_outputs[4026] = inputs[167];
    assign layer0_outputs[4027] = (inputs[159]) | (inputs[235]);
    assign layer0_outputs[4028] = ~(inputs[61]);
    assign layer0_outputs[4029] = ~(inputs[184]);
    assign layer0_outputs[4030] = inputs[151];
    assign layer0_outputs[4031] = inputs[65];
    assign layer0_outputs[4032] = 1'b0;
    assign layer0_outputs[4033] = ~(inputs[241]) | (inputs[78]);
    assign layer0_outputs[4034] = (inputs[5]) | (inputs[131]);
    assign layer0_outputs[4035] = inputs[153];
    assign layer0_outputs[4036] = ~((inputs[165]) ^ (inputs[123]));
    assign layer0_outputs[4037] = inputs[146];
    assign layer0_outputs[4038] = ~((inputs[133]) | (inputs[242]));
    assign layer0_outputs[4039] = (inputs[223]) & (inputs[100]);
    assign layer0_outputs[4040] = ~((inputs[131]) ^ (inputs[20]));
    assign layer0_outputs[4041] = (inputs[69]) ^ (inputs[82]);
    assign layer0_outputs[4042] = (inputs[227]) | (inputs[173]);
    assign layer0_outputs[4043] = inputs[94];
    assign layer0_outputs[4044] = ~(inputs[172]);
    assign layer0_outputs[4045] = (inputs[68]) & ~(inputs[244]);
    assign layer0_outputs[4046] = ~((inputs[188]) & (inputs[94]));
    assign layer0_outputs[4047] = inputs[19];
    assign layer0_outputs[4048] = (inputs[167]) | (inputs[5]);
    assign layer0_outputs[4049] = (inputs[190]) & ~(inputs[26]);
    assign layer0_outputs[4050] = inputs[14];
    assign layer0_outputs[4051] = ~(inputs[133]);
    assign layer0_outputs[4052] = inputs[146];
    assign layer0_outputs[4053] = ~((inputs[11]) | (inputs[50]));
    assign layer0_outputs[4054] = ~((inputs[72]) & (inputs[226]));
    assign layer0_outputs[4055] = inputs[76];
    assign layer0_outputs[4056] = (inputs[248]) ^ (inputs[105]);
    assign layer0_outputs[4057] = (inputs[27]) & ~(inputs[209]);
    assign layer0_outputs[4058] = ~((inputs[201]) & (inputs[227]));
    assign layer0_outputs[4059] = (inputs[249]) | (inputs[150]);
    assign layer0_outputs[4060] = (inputs[9]) | (inputs[172]);
    assign layer0_outputs[4061] = (inputs[20]) ^ (inputs[156]);
    assign layer0_outputs[4062] = (inputs[126]) & ~(inputs[131]);
    assign layer0_outputs[4063] = ~(inputs[141]);
    assign layer0_outputs[4064] = ~((inputs[225]) | (inputs[247]));
    assign layer0_outputs[4065] = ~(inputs[105]);
    assign layer0_outputs[4066] = ~((inputs[135]) & (inputs[85]));
    assign layer0_outputs[4067] = (inputs[104]) ^ (inputs[59]);
    assign layer0_outputs[4068] = (inputs[154]) & ~(inputs[15]);
    assign layer0_outputs[4069] = ~((inputs[140]) & (inputs[12]));
    assign layer0_outputs[4070] = (inputs[52]) ^ (inputs[48]);
    assign layer0_outputs[4071] = ~(inputs[188]);
    assign layer0_outputs[4072] = (inputs[158]) & ~(inputs[255]);
    assign layer0_outputs[4073] = (inputs[20]) | (inputs[226]);
    assign layer0_outputs[4074] = inputs[20];
    assign layer0_outputs[4075] = ~(inputs[22]);
    assign layer0_outputs[4076] = ~((inputs[151]) & (inputs[136]));
    assign layer0_outputs[4077] = ~((inputs[40]) ^ (inputs[69]));
    assign layer0_outputs[4078] = ~(inputs[177]) | (inputs[240]);
    assign layer0_outputs[4079] = ~(inputs[218]);
    assign layer0_outputs[4080] = (inputs[214]) & ~(inputs[203]);
    assign layer0_outputs[4081] = inputs[182];
    assign layer0_outputs[4082] = inputs[147];
    assign layer0_outputs[4083] = ~(inputs[23]);
    assign layer0_outputs[4084] = (inputs[190]) & ~(inputs[65]);
    assign layer0_outputs[4085] = (inputs[103]) ^ (inputs[14]);
    assign layer0_outputs[4086] = ~((inputs[244]) | (inputs[228]));
    assign layer0_outputs[4087] = ~((inputs[19]) | (inputs[78]));
    assign layer0_outputs[4088] = (inputs[38]) & ~(inputs[92]);
    assign layer0_outputs[4089] = ~((inputs[111]) | (inputs[53]));
    assign layer0_outputs[4090] = ~((inputs[72]) ^ (inputs[181]));
    assign layer0_outputs[4091] = ~((inputs[230]) | (inputs[68]));
    assign layer0_outputs[4092] = inputs[148];
    assign layer0_outputs[4093] = ~(inputs[212]);
    assign layer0_outputs[4094] = ~((inputs[47]) | (inputs[73]));
    assign layer0_outputs[4095] = (inputs[216]) & ~(inputs[128]);
    assign layer0_outputs[4096] = ~(inputs[77]);
    assign layer0_outputs[4097] = (inputs[56]) & (inputs[207]);
    assign layer0_outputs[4098] = (inputs[85]) & ~(inputs[47]);
    assign layer0_outputs[4099] = (inputs[186]) & ~(inputs[207]);
    assign layer0_outputs[4100] = (inputs[231]) ^ (inputs[105]);
    assign layer0_outputs[4101] = ~((inputs[135]) ^ (inputs[122]));
    assign layer0_outputs[4102] = ~(inputs[74]) | (inputs[196]);
    assign layer0_outputs[4103] = inputs[57];
    assign layer0_outputs[4104] = (inputs[9]) & (inputs[129]);
    assign layer0_outputs[4105] = ~((inputs[117]) ^ (inputs[34]));
    assign layer0_outputs[4106] = ~(inputs[105]) | (inputs[208]);
    assign layer0_outputs[4107] = ~((inputs[11]) & (inputs[134]));
    assign layer0_outputs[4108] = ~((inputs[193]) | (inputs[9]));
    assign layer0_outputs[4109] = (inputs[114]) & ~(inputs[252]);
    assign layer0_outputs[4110] = ~(inputs[77]);
    assign layer0_outputs[4111] = ~((inputs[119]) ^ (inputs[169]));
    assign layer0_outputs[4112] = ~(inputs[21]);
    assign layer0_outputs[4113] = ~(inputs[39]);
    assign layer0_outputs[4114] = ~(inputs[144]);
    assign layer0_outputs[4115] = ~(inputs[149]);
    assign layer0_outputs[4116] = ~((inputs[35]) | (inputs[210]));
    assign layer0_outputs[4117] = (inputs[51]) | (inputs[37]);
    assign layer0_outputs[4118] = inputs[249];
    assign layer0_outputs[4119] = (inputs[56]) | (inputs[57]);
    assign layer0_outputs[4120] = ~(inputs[220]);
    assign layer0_outputs[4121] = inputs[117];
    assign layer0_outputs[4122] = (inputs[97]) & ~(inputs[175]);
    assign layer0_outputs[4123] = ~(inputs[206]);
    assign layer0_outputs[4124] = ~((inputs[42]) ^ (inputs[17]));
    assign layer0_outputs[4125] = (inputs[217]) & (inputs[0]);
    assign layer0_outputs[4126] = inputs[163];
    assign layer0_outputs[4127] = (inputs[220]) & ~(inputs[110]);
    assign layer0_outputs[4128] = (inputs[183]) | (inputs[32]);
    assign layer0_outputs[4129] = ~(inputs[140]) | (inputs[3]);
    assign layer0_outputs[4130] = inputs[220];
    assign layer0_outputs[4131] = ~((inputs[60]) ^ (inputs[168]));
    assign layer0_outputs[4132] = ~(inputs[119]);
    assign layer0_outputs[4133] = ~(inputs[124]);
    assign layer0_outputs[4134] = ~(inputs[163]);
    assign layer0_outputs[4135] = ~(inputs[74]) | (inputs[203]);
    assign layer0_outputs[4136] = ~(inputs[11]) | (inputs[214]);
    assign layer0_outputs[4137] = (inputs[215]) ^ (inputs[94]);
    assign layer0_outputs[4138] = (inputs[177]) | (inputs[182]);
    assign layer0_outputs[4139] = (inputs[205]) | (inputs[211]);
    assign layer0_outputs[4140] = inputs[26];
    assign layer0_outputs[4141] = ~(inputs[237]);
    assign layer0_outputs[4142] = ~((inputs[155]) ^ (inputs[138]));
    assign layer0_outputs[4143] = (inputs[105]) | (inputs[84]);
    assign layer0_outputs[4144] = (inputs[243]) ^ (inputs[17]);
    assign layer0_outputs[4145] = inputs[230];
    assign layer0_outputs[4146] = ~((inputs[165]) ^ (inputs[189]));
    assign layer0_outputs[4147] = inputs[252];
    assign layer0_outputs[4148] = ~((inputs[16]) | (inputs[122]));
    assign layer0_outputs[4149] = ~(inputs[229]);
    assign layer0_outputs[4150] = inputs[211];
    assign layer0_outputs[4151] = inputs[101];
    assign layer0_outputs[4152] = ~((inputs[114]) ^ (inputs[105]));
    assign layer0_outputs[4153] = (inputs[73]) ^ (inputs[210]);
    assign layer0_outputs[4154] = inputs[34];
    assign layer0_outputs[4155] = ~(inputs[123]) | (inputs[72]);
    assign layer0_outputs[4156] = ~((inputs[90]) | (inputs[47]));
    assign layer0_outputs[4157] = ~(inputs[58]);
    assign layer0_outputs[4158] = ~(inputs[42]) | (inputs[194]);
    assign layer0_outputs[4159] = ~((inputs[128]) & (inputs[93]));
    assign layer0_outputs[4160] = (inputs[121]) | (inputs[20]);
    assign layer0_outputs[4161] = ~((inputs[149]) ^ (inputs[97]));
    assign layer0_outputs[4162] = ~(inputs[195]) | (inputs[30]);
    assign layer0_outputs[4163] = ~(inputs[126]) | (inputs[240]);
    assign layer0_outputs[4164] = inputs[18];
    assign layer0_outputs[4165] = inputs[221];
    assign layer0_outputs[4166] = ~((inputs[195]) | (inputs[194]));
    assign layer0_outputs[4167] = ~(inputs[180]);
    assign layer0_outputs[4168] = ~(inputs[183]);
    assign layer0_outputs[4169] = ~(inputs[46]) | (inputs[223]);
    assign layer0_outputs[4170] = (inputs[77]) ^ (inputs[92]);
    assign layer0_outputs[4171] = ~(inputs[99]) | (inputs[68]);
    assign layer0_outputs[4172] = ~((inputs[139]) | (inputs[63]));
    assign layer0_outputs[4173] = (inputs[52]) | (inputs[241]);
    assign layer0_outputs[4174] = ~(inputs[200]) | (inputs[94]);
    assign layer0_outputs[4175] = ~((inputs[50]) & (inputs[76]));
    assign layer0_outputs[4176] = (inputs[203]) & ~(inputs[186]);
    assign layer0_outputs[4177] = inputs[152];
    assign layer0_outputs[4178] = (inputs[142]) ^ (inputs[102]);
    assign layer0_outputs[4179] = (inputs[175]) | (inputs[66]);
    assign layer0_outputs[4180] = ~((inputs[102]) ^ (inputs[203]));
    assign layer0_outputs[4181] = ~(inputs[211]);
    assign layer0_outputs[4182] = (inputs[78]) | (inputs[42]);
    assign layer0_outputs[4183] = ~(inputs[167]) | (inputs[36]);
    assign layer0_outputs[4184] = ~((inputs[192]) & (inputs[80]));
    assign layer0_outputs[4185] = (inputs[32]) ^ (inputs[53]);
    assign layer0_outputs[4186] = ~((inputs[252]) | (inputs[115]));
    assign layer0_outputs[4187] = inputs[211];
    assign layer0_outputs[4188] = (inputs[136]) & ~(inputs[1]);
    assign layer0_outputs[4189] = ~((inputs[51]) ^ (inputs[90]));
    assign layer0_outputs[4190] = ~(inputs[71]) | (inputs[188]);
    assign layer0_outputs[4191] = ~((inputs[49]) | (inputs[88]));
    assign layer0_outputs[4192] = (inputs[235]) | (inputs[136]);
    assign layer0_outputs[4193] = ~(inputs[76]) | (inputs[195]);
    assign layer0_outputs[4194] = ~(inputs[186]);
    assign layer0_outputs[4195] = ~((inputs[249]) | (inputs[158]));
    assign layer0_outputs[4196] = (inputs[81]) ^ (inputs[5]);
    assign layer0_outputs[4197] = inputs[8];
    assign layer0_outputs[4198] = ~(inputs[203]);
    assign layer0_outputs[4199] = (inputs[116]) ^ (inputs[129]);
    assign layer0_outputs[4200] = ~(inputs[130]);
    assign layer0_outputs[4201] = ~(inputs[221]) | (inputs[120]);
    assign layer0_outputs[4202] = (inputs[172]) & ~(inputs[160]);
    assign layer0_outputs[4203] = ~(inputs[150]);
    assign layer0_outputs[4204] = ~((inputs[82]) | (inputs[8]));
    assign layer0_outputs[4205] = ~((inputs[64]) | (inputs[213]));
    assign layer0_outputs[4206] = ~((inputs[74]) ^ (inputs[64]));
    assign layer0_outputs[4207] = ~(inputs[28]) | (inputs[58]);
    assign layer0_outputs[4208] = inputs[231];
    assign layer0_outputs[4209] = ~(inputs[173]);
    assign layer0_outputs[4210] = (inputs[83]) & ~(inputs[176]);
    assign layer0_outputs[4211] = (inputs[99]) | (inputs[12]);
    assign layer0_outputs[4212] = ~(inputs[204]) | (inputs[34]);
    assign layer0_outputs[4213] = inputs[184];
    assign layer0_outputs[4214] = ~(inputs[241]) | (inputs[179]);
    assign layer0_outputs[4215] = ~((inputs[212]) | (inputs[168]));
    assign layer0_outputs[4216] = ~((inputs[108]) ^ (inputs[104]));
    assign layer0_outputs[4217] = ~((inputs[55]) ^ (inputs[52]));
    assign layer0_outputs[4218] = inputs[95];
    assign layer0_outputs[4219] = inputs[145];
    assign layer0_outputs[4220] = ~((inputs[0]) | (inputs[54]));
    assign layer0_outputs[4221] = ~((inputs[166]) ^ (inputs[205]));
    assign layer0_outputs[4222] = 1'b1;
    assign layer0_outputs[4223] = ~(inputs[2]);
    assign layer0_outputs[4224] = ~((inputs[216]) | (inputs[96]));
    assign layer0_outputs[4225] = inputs[165];
    assign layer0_outputs[4226] = inputs[127];
    assign layer0_outputs[4227] = (inputs[54]) & ~(inputs[166]);
    assign layer0_outputs[4228] = ~(inputs[229]);
    assign layer0_outputs[4229] = ~((inputs[10]) | (inputs[50]));
    assign layer0_outputs[4230] = (inputs[29]) | (inputs[60]);
    assign layer0_outputs[4231] = (inputs[86]) ^ (inputs[130]);
    assign layer0_outputs[4232] = (inputs[17]) ^ (inputs[186]);
    assign layer0_outputs[4233] = inputs[35];
    assign layer0_outputs[4234] = (inputs[215]) ^ (inputs[215]);
    assign layer0_outputs[4235] = ~(inputs[51]);
    assign layer0_outputs[4236] = (inputs[173]) & (inputs[231]);
    assign layer0_outputs[4237] = inputs[219];
    assign layer0_outputs[4238] = (inputs[151]) & ~(inputs[147]);
    assign layer0_outputs[4239] = (inputs[183]) | (inputs[48]);
    assign layer0_outputs[4240] = (inputs[185]) ^ (inputs[65]);
    assign layer0_outputs[4241] = inputs[154];
    assign layer0_outputs[4242] = 1'b1;
    assign layer0_outputs[4243] = ~((inputs[194]) | (inputs[83]));
    assign layer0_outputs[4244] = (inputs[116]) | (inputs[88]);
    assign layer0_outputs[4245] = inputs[132];
    assign layer0_outputs[4246] = ~(inputs[60]);
    assign layer0_outputs[4247] = (inputs[103]) ^ (inputs[229]);
    assign layer0_outputs[4248] = inputs[214];
    assign layer0_outputs[4249] = (inputs[186]) | (inputs[253]);
    assign layer0_outputs[4250] = ~((inputs[178]) | (inputs[78]));
    assign layer0_outputs[4251] = (inputs[249]) & ~(inputs[169]);
    assign layer0_outputs[4252] = (inputs[35]) | (inputs[71]);
    assign layer0_outputs[4253] = (inputs[155]) & ~(inputs[7]);
    assign layer0_outputs[4254] = ~(inputs[100]);
    assign layer0_outputs[4255] = ~((inputs[37]) | (inputs[30]));
    assign layer0_outputs[4256] = ~(inputs[165]);
    assign layer0_outputs[4257] = ~((inputs[15]) ^ (inputs[244]));
    assign layer0_outputs[4258] = (inputs[218]) ^ (inputs[20]);
    assign layer0_outputs[4259] = (inputs[81]) | (inputs[66]);
    assign layer0_outputs[4260] = ~((inputs[45]) & (inputs[24]));
    assign layer0_outputs[4261] = ~((inputs[114]) ^ (inputs[34]));
    assign layer0_outputs[4262] = inputs[119];
    assign layer0_outputs[4263] = ~((inputs[175]) | (inputs[42]));
    assign layer0_outputs[4264] = (inputs[155]) & (inputs[105]);
    assign layer0_outputs[4265] = ~((inputs[106]) | (inputs[23]));
    assign layer0_outputs[4266] = (inputs[226]) | (inputs[84]);
    assign layer0_outputs[4267] = (inputs[7]) & ~(inputs[61]);
    assign layer0_outputs[4268] = (inputs[61]) | (inputs[237]);
    assign layer0_outputs[4269] = (inputs[10]) ^ (inputs[255]);
    assign layer0_outputs[4270] = (inputs[174]) ^ (inputs[239]);
    assign layer0_outputs[4271] = ~((inputs[204]) | (inputs[118]));
    assign layer0_outputs[4272] = ~(inputs[78]);
    assign layer0_outputs[4273] = ~((inputs[135]) ^ (inputs[240]));
    assign layer0_outputs[4274] = ~((inputs[36]) ^ (inputs[0]));
    assign layer0_outputs[4275] = inputs[113];
    assign layer0_outputs[4276] = ~((inputs[137]) | (inputs[10]));
    assign layer0_outputs[4277] = ~((inputs[239]) | (inputs[248]));
    assign layer0_outputs[4278] = ~(inputs[141]);
    assign layer0_outputs[4279] = (inputs[169]) | (inputs[126]);
    assign layer0_outputs[4280] = ~(inputs[233]);
    assign layer0_outputs[4281] = ~(inputs[100]);
    assign layer0_outputs[4282] = ~((inputs[66]) ^ (inputs[139]));
    assign layer0_outputs[4283] = ~((inputs[114]) | (inputs[72]));
    assign layer0_outputs[4284] = ~((inputs[23]) ^ (inputs[55]));
    assign layer0_outputs[4285] = inputs[145];
    assign layer0_outputs[4286] = (inputs[65]) ^ (inputs[198]);
    assign layer0_outputs[4287] = 1'b0;
    assign layer0_outputs[4288] = ~(inputs[66]) | (inputs[253]);
    assign layer0_outputs[4289] = ~((inputs[233]) | (inputs[218]));
    assign layer0_outputs[4290] = (inputs[98]) ^ (inputs[36]);
    assign layer0_outputs[4291] = ~((inputs[128]) ^ (inputs[118]));
    assign layer0_outputs[4292] = ~(inputs[9]) | (inputs[210]);
    assign layer0_outputs[4293] = ~((inputs[196]) | (inputs[97]));
    assign layer0_outputs[4294] = (inputs[133]) & ~(inputs[21]);
    assign layer0_outputs[4295] = inputs[30];
    assign layer0_outputs[4296] = inputs[243];
    assign layer0_outputs[4297] = 1'b1;
    assign layer0_outputs[4298] = (inputs[170]) & ~(inputs[86]);
    assign layer0_outputs[4299] = inputs[24];
    assign layer0_outputs[4300] = ~((inputs[143]) & (inputs[201]));
    assign layer0_outputs[4301] = (inputs[170]) ^ (inputs[107]);
    assign layer0_outputs[4302] = ~(inputs[5]) | (inputs[190]);
    assign layer0_outputs[4303] = ~(inputs[117]);
    assign layer0_outputs[4304] = (inputs[208]) | (inputs[211]);
    assign layer0_outputs[4305] = inputs[51];
    assign layer0_outputs[4306] = ~(inputs[139]) | (inputs[27]);
    assign layer0_outputs[4307] = ~(inputs[233]) | (inputs[56]);
    assign layer0_outputs[4308] = ~((inputs[28]) | (inputs[5]));
    assign layer0_outputs[4309] = (inputs[174]) & ~(inputs[101]);
    assign layer0_outputs[4310] = (inputs[99]) & ~(inputs[2]);
    assign layer0_outputs[4311] = (inputs[17]) | (inputs[147]);
    assign layer0_outputs[4312] = ~((inputs[16]) ^ (inputs[36]));
    assign layer0_outputs[4313] = inputs[195];
    assign layer0_outputs[4314] = ~((inputs[222]) ^ (inputs[116]));
    assign layer0_outputs[4315] = ~((inputs[245]) ^ (inputs[95]));
    assign layer0_outputs[4316] = (inputs[107]) & ~(inputs[233]);
    assign layer0_outputs[4317] = ~((inputs[66]) ^ (inputs[191]));
    assign layer0_outputs[4318] = inputs[167];
    assign layer0_outputs[4319] = ~((inputs[139]) & (inputs[133]));
    assign layer0_outputs[4320] = (inputs[56]) & (inputs[88]);
    assign layer0_outputs[4321] = (inputs[124]) & ~(inputs[22]);
    assign layer0_outputs[4322] = ~((inputs[166]) ^ (inputs[184]));
    assign layer0_outputs[4323] = ~((inputs[168]) ^ (inputs[74]));
    assign layer0_outputs[4324] = (inputs[233]) & ~(inputs[2]);
    assign layer0_outputs[4325] = inputs[166];
    assign layer0_outputs[4326] = (inputs[167]) & ~(inputs[68]);
    assign layer0_outputs[4327] = (inputs[193]) ^ (inputs[196]);
    assign layer0_outputs[4328] = ~(inputs[250]);
    assign layer0_outputs[4329] = (inputs[191]) & (inputs[238]);
    assign layer0_outputs[4330] = ~((inputs[7]) ^ (inputs[237]));
    assign layer0_outputs[4331] = ~((inputs[85]) & (inputs[165]));
    assign layer0_outputs[4332] = ~(inputs[116]);
    assign layer0_outputs[4333] = ~(inputs[228]) | (inputs[83]);
    assign layer0_outputs[4334] = ~(inputs[118]);
    assign layer0_outputs[4335] = ~(inputs[237]);
    assign layer0_outputs[4336] = (inputs[141]) & ~(inputs[31]);
    assign layer0_outputs[4337] = ~((inputs[224]) ^ (inputs[21]));
    assign layer0_outputs[4338] = inputs[104];
    assign layer0_outputs[4339] = (inputs[194]) | (inputs[222]);
    assign layer0_outputs[4340] = ~((inputs[169]) | (inputs[6]));
    assign layer0_outputs[4341] = (inputs[255]) ^ (inputs[114]);
    assign layer0_outputs[4342] = (inputs[107]) ^ (inputs[136]);
    assign layer0_outputs[4343] = ~(inputs[40]);
    assign layer0_outputs[4344] = ~((inputs[84]) | (inputs[29]));
    assign layer0_outputs[4345] = (inputs[25]) & ~(inputs[136]);
    assign layer0_outputs[4346] = (inputs[214]) | (inputs[96]);
    assign layer0_outputs[4347] = ~(inputs[232]);
    assign layer0_outputs[4348] = ~((inputs[222]) ^ (inputs[193]));
    assign layer0_outputs[4349] = inputs[5];
    assign layer0_outputs[4350] = (inputs[190]) | (inputs[192]);
    assign layer0_outputs[4351] = (inputs[191]) | (inputs[251]);
    assign layer0_outputs[4352] = ~(inputs[170]) | (inputs[72]);
    assign layer0_outputs[4353] = inputs[76];
    assign layer0_outputs[4354] = ~((inputs[122]) & (inputs[91]));
    assign layer0_outputs[4355] = ~((inputs[183]) ^ (inputs[28]));
    assign layer0_outputs[4356] = ~(inputs[216]) | (inputs[220]);
    assign layer0_outputs[4357] = ~(inputs[111]) | (inputs[1]);
    assign layer0_outputs[4358] = (inputs[255]) ^ (inputs[173]);
    assign layer0_outputs[4359] = ~((inputs[75]) | (inputs[77]));
    assign layer0_outputs[4360] = ~((inputs[92]) ^ (inputs[255]));
    assign layer0_outputs[4361] = (inputs[21]) & ~(inputs[157]);
    assign layer0_outputs[4362] = ~(inputs[60]);
    assign layer0_outputs[4363] = (inputs[198]) & ~(inputs[183]);
    assign layer0_outputs[4364] = ~((inputs[243]) & (inputs[201]));
    assign layer0_outputs[4365] = ~((inputs[220]) | (inputs[54]));
    assign layer0_outputs[4366] = ~((inputs[249]) | (inputs[142]));
    assign layer0_outputs[4367] = ~(inputs[118]);
    assign layer0_outputs[4368] = (inputs[100]) & ~(inputs[192]);
    assign layer0_outputs[4369] = 1'b0;
    assign layer0_outputs[4370] = inputs[8];
    assign layer0_outputs[4371] = (inputs[85]) & ~(inputs[125]);
    assign layer0_outputs[4372] = (inputs[27]) | (inputs[51]);
    assign layer0_outputs[4373] = ~(inputs[113]);
    assign layer0_outputs[4374] = (inputs[104]) ^ (inputs[48]);
    assign layer0_outputs[4375] = ~(inputs[90]) | (inputs[250]);
    assign layer0_outputs[4376] = ~((inputs[45]) ^ (inputs[87]));
    assign layer0_outputs[4377] = ~((inputs[0]) | (inputs[153]));
    assign layer0_outputs[4378] = inputs[184];
    assign layer0_outputs[4379] = inputs[74];
    assign layer0_outputs[4380] = ~(inputs[183]) | (inputs[191]);
    assign layer0_outputs[4381] = inputs[72];
    assign layer0_outputs[4382] = ~(inputs[59]);
    assign layer0_outputs[4383] = inputs[73];
    assign layer0_outputs[4384] = ~(inputs[118]);
    assign layer0_outputs[4385] = ~(inputs[9]);
    assign layer0_outputs[4386] = ~(inputs[104]);
    assign layer0_outputs[4387] = (inputs[175]) & ~(inputs[54]);
    assign layer0_outputs[4388] = ~((inputs[32]) ^ (inputs[200]));
    assign layer0_outputs[4389] = ~((inputs[206]) | (inputs[98]));
    assign layer0_outputs[4390] = (inputs[60]) ^ (inputs[79]);
    assign layer0_outputs[4391] = ~(inputs[98]);
    assign layer0_outputs[4392] = inputs[134];
    assign layer0_outputs[4393] = ~((inputs[172]) | (inputs[130]));
    assign layer0_outputs[4394] = (inputs[79]) | (inputs[245]);
    assign layer0_outputs[4395] = inputs[16];
    assign layer0_outputs[4396] = ~(inputs[244]);
    assign layer0_outputs[4397] = ~(inputs[176]);
    assign layer0_outputs[4398] = ~((inputs[69]) ^ (inputs[83]));
    assign layer0_outputs[4399] = inputs[35];
    assign layer0_outputs[4400] = (inputs[86]) | (inputs[141]);
    assign layer0_outputs[4401] = ~((inputs[161]) & (inputs[227]));
    assign layer0_outputs[4402] = (inputs[34]) ^ (inputs[123]);
    assign layer0_outputs[4403] = inputs[109];
    assign layer0_outputs[4404] = ~(inputs[98]) | (inputs[94]);
    assign layer0_outputs[4405] = ~((inputs[125]) ^ (inputs[88]));
    assign layer0_outputs[4406] = ~((inputs[230]) ^ (inputs[135]));
    assign layer0_outputs[4407] = 1'b1;
    assign layer0_outputs[4408] = ~(inputs[8]);
    assign layer0_outputs[4409] = ~(inputs[99]);
    assign layer0_outputs[4410] = inputs[104];
    assign layer0_outputs[4411] = (inputs[115]) | (inputs[171]);
    assign layer0_outputs[4412] = ~(inputs[93]);
    assign layer0_outputs[4413] = (inputs[54]) & ~(inputs[113]);
    assign layer0_outputs[4414] = (inputs[32]) ^ (inputs[168]);
    assign layer0_outputs[4415] = ~(inputs[178]);
    assign layer0_outputs[4416] = 1'b0;
    assign layer0_outputs[4417] = ~((inputs[112]) | (inputs[124]));
    assign layer0_outputs[4418] = (inputs[46]) & ~(inputs[76]);
    assign layer0_outputs[4419] = ~((inputs[133]) | (inputs[227]));
    assign layer0_outputs[4420] = (inputs[237]) | (inputs[87]);
    assign layer0_outputs[4421] = (inputs[73]) | (inputs[57]);
    assign layer0_outputs[4422] = ~((inputs[114]) | (inputs[145]));
    assign layer0_outputs[4423] = (inputs[143]) ^ (inputs[212]);
    assign layer0_outputs[4424] = ~(inputs[146]);
    assign layer0_outputs[4425] = (inputs[137]) ^ (inputs[234]);
    assign layer0_outputs[4426] = ~((inputs[87]) ^ (inputs[101]));
    assign layer0_outputs[4427] = (inputs[238]) ^ (inputs[17]);
    assign layer0_outputs[4428] = (inputs[180]) & ~(inputs[128]);
    assign layer0_outputs[4429] = ~((inputs[6]) ^ (inputs[52]));
    assign layer0_outputs[4430] = inputs[167];
    assign layer0_outputs[4431] = (inputs[136]) & ~(inputs[61]);
    assign layer0_outputs[4432] = ~((inputs[220]) | (inputs[255]));
    assign layer0_outputs[4433] = (inputs[205]) ^ (inputs[23]);
    assign layer0_outputs[4434] = 1'b0;
    assign layer0_outputs[4435] = inputs[187];
    assign layer0_outputs[4436] = 1'b1;
    assign layer0_outputs[4437] = (inputs[111]) | (inputs[220]);
    assign layer0_outputs[4438] = ~((inputs[104]) ^ (inputs[59]));
    assign layer0_outputs[4439] = (inputs[35]) ^ (inputs[11]);
    assign layer0_outputs[4440] = ~(inputs[241]);
    assign layer0_outputs[4441] = (inputs[101]) | (inputs[145]);
    assign layer0_outputs[4442] = ~((inputs[131]) & (inputs[159]));
    assign layer0_outputs[4443] = (inputs[61]) & ~(inputs[100]);
    assign layer0_outputs[4444] = ~(inputs[129]) | (inputs[252]);
    assign layer0_outputs[4445] = ~((inputs[45]) ^ (inputs[195]));
    assign layer0_outputs[4446] = (inputs[187]) ^ (inputs[5]);
    assign layer0_outputs[4447] = ~(inputs[70]) | (inputs[194]);
    assign layer0_outputs[4448] = ~(inputs[196]) | (inputs[39]);
    assign layer0_outputs[4449] = (inputs[49]) ^ (inputs[242]);
    assign layer0_outputs[4450] = (inputs[43]) & ~(inputs[221]);
    assign layer0_outputs[4451] = (inputs[112]) | (inputs[234]);
    assign layer0_outputs[4452] = inputs[83];
    assign layer0_outputs[4453] = (inputs[99]) & ~(inputs[79]);
    assign layer0_outputs[4454] = ~(inputs[212]);
    assign layer0_outputs[4455] = ~((inputs[131]) ^ (inputs[199]));
    assign layer0_outputs[4456] = ~(inputs[108]);
    assign layer0_outputs[4457] = ~((inputs[218]) | (inputs[205]));
    assign layer0_outputs[4458] = inputs[134];
    assign layer0_outputs[4459] = ~((inputs[240]) ^ (inputs[63]));
    assign layer0_outputs[4460] = ~((inputs[192]) | (inputs[166]));
    assign layer0_outputs[4461] = (inputs[83]) & ~(inputs[2]);
    assign layer0_outputs[4462] = ~(inputs[7]);
    assign layer0_outputs[4463] = inputs[24];
    assign layer0_outputs[4464] = (inputs[42]) & ~(inputs[211]);
    assign layer0_outputs[4465] = ~(inputs[120]) | (inputs[175]);
    assign layer0_outputs[4466] = ~((inputs[53]) | (inputs[101]));
    assign layer0_outputs[4467] = ~(inputs[28]);
    assign layer0_outputs[4468] = inputs[151];
    assign layer0_outputs[4469] = (inputs[159]) ^ (inputs[224]);
    assign layer0_outputs[4470] = (inputs[229]) | (inputs[245]);
    assign layer0_outputs[4471] = ~(inputs[194]) | (inputs[253]);
    assign layer0_outputs[4472] = ~(inputs[101]);
    assign layer0_outputs[4473] = ~(inputs[150]);
    assign layer0_outputs[4474] = (inputs[102]) ^ (inputs[38]);
    assign layer0_outputs[4475] = (inputs[224]) | (inputs[16]);
    assign layer0_outputs[4476] = inputs[76];
    assign layer0_outputs[4477] = (inputs[165]) ^ (inputs[240]);
    assign layer0_outputs[4478] = ~(inputs[71]);
    assign layer0_outputs[4479] = inputs[93];
    assign layer0_outputs[4480] = inputs[230];
    assign layer0_outputs[4481] = (inputs[194]) | (inputs[171]);
    assign layer0_outputs[4482] = inputs[85];
    assign layer0_outputs[4483] = ~(inputs[107]);
    assign layer0_outputs[4484] = ~(inputs[162]);
    assign layer0_outputs[4485] = inputs[23];
    assign layer0_outputs[4486] = ~(inputs[121]) | (inputs[57]);
    assign layer0_outputs[4487] = (inputs[246]) | (inputs[141]);
    assign layer0_outputs[4488] = ~((inputs[41]) | (inputs[57]));
    assign layer0_outputs[4489] = ~((inputs[82]) ^ (inputs[68]));
    assign layer0_outputs[4490] = inputs[38];
    assign layer0_outputs[4491] = ~(inputs[125]) | (inputs[134]);
    assign layer0_outputs[4492] = inputs[125];
    assign layer0_outputs[4493] = (inputs[149]) ^ (inputs[148]);
    assign layer0_outputs[4494] = ~((inputs[15]) ^ (inputs[69]));
    assign layer0_outputs[4495] = (inputs[173]) & (inputs[122]);
    assign layer0_outputs[4496] = (inputs[56]) & (inputs[119]);
    assign layer0_outputs[4497] = ~(inputs[129]);
    assign layer0_outputs[4498] = ~((inputs[30]) ^ (inputs[218]));
    assign layer0_outputs[4499] = ~(inputs[91]) | (inputs[223]);
    assign layer0_outputs[4500] = ~(inputs[156]);
    assign layer0_outputs[4501] = ~(inputs[60]) | (inputs[104]);
    assign layer0_outputs[4502] = ~((inputs[45]) ^ (inputs[18]));
    assign layer0_outputs[4503] = ~(inputs[105]);
    assign layer0_outputs[4504] = ~((inputs[51]) ^ (inputs[239]));
    assign layer0_outputs[4505] = inputs[130];
    assign layer0_outputs[4506] = ~(inputs[9]);
    assign layer0_outputs[4507] = ~((inputs[233]) | (inputs[213]));
    assign layer0_outputs[4508] = ~(inputs[4]) | (inputs[15]);
    assign layer0_outputs[4509] = ~(inputs[118]);
    assign layer0_outputs[4510] = inputs[214];
    assign layer0_outputs[4511] = ~(inputs[232]);
    assign layer0_outputs[4512] = (inputs[141]) | (inputs[1]);
    assign layer0_outputs[4513] = (inputs[83]) | (inputs[163]);
    assign layer0_outputs[4514] = (inputs[115]) & ~(inputs[17]);
    assign layer0_outputs[4515] = (inputs[165]) ^ (inputs[23]);
    assign layer0_outputs[4516] = ~(inputs[105]) | (inputs[130]);
    assign layer0_outputs[4517] = (inputs[216]) & ~(inputs[8]);
    assign layer0_outputs[4518] = ~(inputs[217]);
    assign layer0_outputs[4519] = (inputs[214]) | (inputs[19]);
    assign layer0_outputs[4520] = (inputs[227]) | (inputs[246]);
    assign layer0_outputs[4521] = (inputs[89]) & ~(inputs[70]);
    assign layer0_outputs[4522] = (inputs[127]) & ~(inputs[88]);
    assign layer0_outputs[4523] = (inputs[89]) ^ (inputs[107]);
    assign layer0_outputs[4524] = ~(inputs[66]);
    assign layer0_outputs[4525] = ~(inputs[163]);
    assign layer0_outputs[4526] = ~(inputs[109]) | (inputs[82]);
    assign layer0_outputs[4527] = ~(inputs[100]);
    assign layer0_outputs[4528] = ~(inputs[200]) | (inputs[63]);
    assign layer0_outputs[4529] = ~(inputs[74]);
    assign layer0_outputs[4530] = ~(inputs[107]);
    assign layer0_outputs[4531] = ~(inputs[3]);
    assign layer0_outputs[4532] = (inputs[96]) | (inputs[183]);
    assign layer0_outputs[4533] = ~(inputs[182]);
    assign layer0_outputs[4534] = (inputs[127]) & ~(inputs[249]);
    assign layer0_outputs[4535] = ~((inputs[52]) | (inputs[128]));
    assign layer0_outputs[4536] = (inputs[52]) | (inputs[94]);
    assign layer0_outputs[4537] = ~(inputs[26]) | (inputs[244]);
    assign layer0_outputs[4538] = (inputs[180]) | (inputs[32]);
    assign layer0_outputs[4539] = ~((inputs[205]) | (inputs[192]));
    assign layer0_outputs[4540] = (inputs[180]) | (inputs[152]);
    assign layer0_outputs[4541] = (inputs[22]) ^ (inputs[147]);
    assign layer0_outputs[4542] = ~((inputs[109]) | (inputs[95]));
    assign layer0_outputs[4543] = (inputs[249]) ^ (inputs[202]);
    assign layer0_outputs[4544] = ~(inputs[75]);
    assign layer0_outputs[4545] = (inputs[32]) | (inputs[197]);
    assign layer0_outputs[4546] = inputs[70];
    assign layer0_outputs[4547] = (inputs[254]) & (inputs[234]);
    assign layer0_outputs[4548] = inputs[224];
    assign layer0_outputs[4549] = ~(inputs[225]) | (inputs[11]);
    assign layer0_outputs[4550] = inputs[30];
    assign layer0_outputs[4551] = (inputs[247]) & ~(inputs[47]);
    assign layer0_outputs[4552] = inputs[10];
    assign layer0_outputs[4553] = ~((inputs[18]) ^ (inputs[94]));
    assign layer0_outputs[4554] = ~(inputs[121]);
    assign layer0_outputs[4555] = inputs[150];
    assign layer0_outputs[4556] = ~((inputs[76]) ^ (inputs[195]));
    assign layer0_outputs[4557] = ~((inputs[7]) & (inputs[223]));
    assign layer0_outputs[4558] = 1'b1;
    assign layer0_outputs[4559] = ~((inputs[122]) | (inputs[106]));
    assign layer0_outputs[4560] = ~((inputs[66]) & (inputs[143]));
    assign layer0_outputs[4561] = ~(inputs[29]);
    assign layer0_outputs[4562] = ~(inputs[109]);
    assign layer0_outputs[4563] = ~((inputs[52]) & (inputs[45]));
    assign layer0_outputs[4564] = (inputs[193]) ^ (inputs[22]);
    assign layer0_outputs[4565] = (inputs[54]) & ~(inputs[34]);
    assign layer0_outputs[4566] = (inputs[123]) ^ (inputs[157]);
    assign layer0_outputs[4567] = inputs[248];
    assign layer0_outputs[4568] = (inputs[95]) | (inputs[55]);
    assign layer0_outputs[4569] = ~(inputs[97]);
    assign layer0_outputs[4570] = ~(inputs[170]) | (inputs[84]);
    assign layer0_outputs[4571] = (inputs[181]) | (inputs[212]);
    assign layer0_outputs[4572] = inputs[192];
    assign layer0_outputs[4573] = ~(inputs[129]);
    assign layer0_outputs[4574] = inputs[29];
    assign layer0_outputs[4575] = ~((inputs[107]) | (inputs[6]));
    assign layer0_outputs[4576] = ~(inputs[102]);
    assign layer0_outputs[4577] = inputs[136];
    assign layer0_outputs[4578] = ~(inputs[108]) | (inputs[31]);
    assign layer0_outputs[4579] = ~(inputs[106]);
    assign layer0_outputs[4580] = (inputs[105]) & ~(inputs[2]);
    assign layer0_outputs[4581] = (inputs[123]) | (inputs[94]);
    assign layer0_outputs[4582] = inputs[98];
    assign layer0_outputs[4583] = (inputs[28]) | (inputs[0]);
    assign layer0_outputs[4584] = (inputs[9]) | (inputs[181]);
    assign layer0_outputs[4585] = ~((inputs[58]) ^ (inputs[72]));
    assign layer0_outputs[4586] = inputs[100];
    assign layer0_outputs[4587] = (inputs[218]) ^ (inputs[171]);
    assign layer0_outputs[4588] = inputs[237];
    assign layer0_outputs[4589] = ~((inputs[102]) ^ (inputs[37]));
    assign layer0_outputs[4590] = inputs[146];
    assign layer0_outputs[4591] = ~((inputs[7]) ^ (inputs[17]));
    assign layer0_outputs[4592] = (inputs[33]) | (inputs[43]);
    assign layer0_outputs[4593] = (inputs[202]) & ~(inputs[143]);
    assign layer0_outputs[4594] = ~((inputs[129]) | (inputs[114]));
    assign layer0_outputs[4595] = inputs[232];
    assign layer0_outputs[4596] = ~((inputs[162]) | (inputs[183]));
    assign layer0_outputs[4597] = (inputs[160]) | (inputs[165]);
    assign layer0_outputs[4598] = ~(inputs[213]) | (inputs[166]);
    assign layer0_outputs[4599] = ~(inputs[113]);
    assign layer0_outputs[4600] = ~(inputs[151]);
    assign layer0_outputs[4601] = (inputs[113]) | (inputs[37]);
    assign layer0_outputs[4602] = (inputs[47]) | (inputs[226]);
    assign layer0_outputs[4603] = (inputs[40]) & ~(inputs[73]);
    assign layer0_outputs[4604] = ~(inputs[130]);
    assign layer0_outputs[4605] = inputs[41];
    assign layer0_outputs[4606] = inputs[162];
    assign layer0_outputs[4607] = ~((inputs[212]) | (inputs[144]));
    assign layer0_outputs[4608] = inputs[94];
    assign layer0_outputs[4609] = (inputs[21]) & ~(inputs[84]);
    assign layer0_outputs[4610] = ~((inputs[68]) ^ (inputs[160]));
    assign layer0_outputs[4611] = ~(inputs[110]) | (inputs[251]);
    assign layer0_outputs[4612] = ~(inputs[40]) | (inputs[242]);
    assign layer0_outputs[4613] = inputs[109];
    assign layer0_outputs[4614] = ~(inputs[140]) | (inputs[177]);
    assign layer0_outputs[4615] = ~((inputs[157]) | (inputs[85]));
    assign layer0_outputs[4616] = (inputs[136]) & ~(inputs[115]);
    assign layer0_outputs[4617] = ~(inputs[27]);
    assign layer0_outputs[4618] = inputs[212];
    assign layer0_outputs[4619] = 1'b0;
    assign layer0_outputs[4620] = inputs[181];
    assign layer0_outputs[4621] = (inputs[91]) & ~(inputs[240]);
    assign layer0_outputs[4622] = (inputs[61]) & (inputs[122]);
    assign layer0_outputs[4623] = (inputs[155]) & ~(inputs[206]);
    assign layer0_outputs[4624] = (inputs[219]) | (inputs[203]);
    assign layer0_outputs[4625] = ~(inputs[92]);
    assign layer0_outputs[4626] = ~(inputs[220]);
    assign layer0_outputs[4627] = ~(inputs[79]);
    assign layer0_outputs[4628] = (inputs[237]) ^ (inputs[106]);
    assign layer0_outputs[4629] = ~((inputs[79]) | (inputs[117]));
    assign layer0_outputs[4630] = ~((inputs[215]) | (inputs[231]));
    assign layer0_outputs[4631] = ~((inputs[69]) | (inputs[63]));
    assign layer0_outputs[4632] = ~(inputs[116]) | (inputs[126]);
    assign layer0_outputs[4633] = inputs[246];
    assign layer0_outputs[4634] = inputs[145];
    assign layer0_outputs[4635] = ~((inputs[39]) & (inputs[40]));
    assign layer0_outputs[4636] = (inputs[150]) & ~(inputs[31]);
    assign layer0_outputs[4637] = inputs[246];
    assign layer0_outputs[4638] = ~(inputs[227]);
    assign layer0_outputs[4639] = ~(inputs[92]);
    assign layer0_outputs[4640] = inputs[246];
    assign layer0_outputs[4641] = ~((inputs[96]) | (inputs[114]));
    assign layer0_outputs[4642] = ~(inputs[229]) | (inputs[166]);
    assign layer0_outputs[4643] = (inputs[69]) & ~(inputs[225]);
    assign layer0_outputs[4644] = ~((inputs[199]) | (inputs[153]));
    assign layer0_outputs[4645] = inputs[109];
    assign layer0_outputs[4646] = (inputs[129]) & (inputs[17]);
    assign layer0_outputs[4647] = ~(inputs[19]) | (inputs[80]);
    assign layer0_outputs[4648] = ~((inputs[143]) ^ (inputs[172]));
    assign layer0_outputs[4649] = ~((inputs[228]) | (inputs[227]));
    assign layer0_outputs[4650] = (inputs[153]) & ~(inputs[18]);
    assign layer0_outputs[4651] = (inputs[123]) & (inputs[91]);
    assign layer0_outputs[4652] = ~((inputs[43]) ^ (inputs[65]));
    assign layer0_outputs[4653] = (inputs[35]) | (inputs[255]);
    assign layer0_outputs[4654] = (inputs[167]) | (inputs[140]);
    assign layer0_outputs[4655] = ~(inputs[201]) | (inputs[35]);
    assign layer0_outputs[4656] = ~((inputs[178]) | (inputs[127]));
    assign layer0_outputs[4657] = inputs[103];
    assign layer0_outputs[4658] = ~(inputs[117]);
    assign layer0_outputs[4659] = ~((inputs[43]) & (inputs[159]));
    assign layer0_outputs[4660] = (inputs[79]) | (inputs[219]);
    assign layer0_outputs[4661] = ~(inputs[99]);
    assign layer0_outputs[4662] = ~((inputs[245]) ^ (inputs[103]));
    assign layer0_outputs[4663] = ~(inputs[85]) | (inputs[250]);
    assign layer0_outputs[4664] = (inputs[160]) ^ (inputs[59]);
    assign layer0_outputs[4665] = ~((inputs[146]) | (inputs[251]));
    assign layer0_outputs[4666] = (inputs[146]) & ~(inputs[66]);
    assign layer0_outputs[4667] = (inputs[255]) & ~(inputs[96]);
    assign layer0_outputs[4668] = ~(inputs[137]) | (inputs[122]);
    assign layer0_outputs[4669] = ~((inputs[38]) & (inputs[104]));
    assign layer0_outputs[4670] = ~((inputs[120]) ^ (inputs[76]));
    assign layer0_outputs[4671] = (inputs[126]) | (inputs[59]);
    assign layer0_outputs[4672] = (inputs[96]) & ~(inputs[250]);
    assign layer0_outputs[4673] = inputs[90];
    assign layer0_outputs[4674] = (inputs[97]) | (inputs[246]);
    assign layer0_outputs[4675] = ~(inputs[164]);
    assign layer0_outputs[4676] = inputs[67];
    assign layer0_outputs[4677] = (inputs[41]) & ~(inputs[253]);
    assign layer0_outputs[4678] = inputs[166];
    assign layer0_outputs[4679] = (inputs[137]) ^ (inputs[213]);
    assign layer0_outputs[4680] = ~(inputs[195]) | (inputs[120]);
    assign layer0_outputs[4681] = ~(inputs[179]) | (inputs[109]);
    assign layer0_outputs[4682] = ~((inputs[202]) ^ (inputs[182]));
    assign layer0_outputs[4683] = ~(inputs[135]);
    assign layer0_outputs[4684] = ~(inputs[199]) | (inputs[62]);
    assign layer0_outputs[4685] = (inputs[36]) & (inputs[246]);
    assign layer0_outputs[4686] = (inputs[178]) | (inputs[185]);
    assign layer0_outputs[4687] = ~(inputs[22]);
    assign layer0_outputs[4688] = ~(inputs[23]) | (inputs[50]);
    assign layer0_outputs[4689] = (inputs[51]) | (inputs[208]);
    assign layer0_outputs[4690] = inputs[255];
    assign layer0_outputs[4691] = inputs[114];
    assign layer0_outputs[4692] = ~(inputs[243]) | (inputs[71]);
    assign layer0_outputs[4693] = (inputs[93]) ^ (inputs[234]);
    assign layer0_outputs[4694] = (inputs[198]) & ~(inputs[87]);
    assign layer0_outputs[4695] = (inputs[130]) | (inputs[78]);
    assign layer0_outputs[4696] = (inputs[198]) & ~(inputs[53]);
    assign layer0_outputs[4697] = ~((inputs[46]) | (inputs[54]));
    assign layer0_outputs[4698] = inputs[75];
    assign layer0_outputs[4699] = ~(inputs[169]);
    assign layer0_outputs[4700] = ~((inputs[234]) | (inputs[25]));
    assign layer0_outputs[4701] = (inputs[191]) | (inputs[233]);
    assign layer0_outputs[4702] = (inputs[181]) | (inputs[96]);
    assign layer0_outputs[4703] = ~(inputs[26]);
    assign layer0_outputs[4704] = (inputs[114]) & ~(inputs[75]);
    assign layer0_outputs[4705] = ~(inputs[136]) | (inputs[238]);
    assign layer0_outputs[4706] = ~(inputs[178]) | (inputs[202]);
    assign layer0_outputs[4707] = ~(inputs[50]);
    assign layer0_outputs[4708] = ~((inputs[163]) | (inputs[220]));
    assign layer0_outputs[4709] = (inputs[8]) & (inputs[105]);
    assign layer0_outputs[4710] = inputs[249];
    assign layer0_outputs[4711] = inputs[9];
    assign layer0_outputs[4712] = (inputs[126]) ^ (inputs[140]);
    assign layer0_outputs[4713] = ~(inputs[177]) | (inputs[249]);
    assign layer0_outputs[4714] = (inputs[161]) & ~(inputs[128]);
    assign layer0_outputs[4715] = inputs[109];
    assign layer0_outputs[4716] = ~(inputs[58]) | (inputs[206]);
    assign layer0_outputs[4717] = (inputs[114]) ^ (inputs[117]);
    assign layer0_outputs[4718] = ~(inputs[183]) | (inputs[57]);
    assign layer0_outputs[4719] = ~(inputs[245]);
    assign layer0_outputs[4720] = inputs[116];
    assign layer0_outputs[4721] = (inputs[154]) & (inputs[7]);
    assign layer0_outputs[4722] = ~((inputs[3]) & (inputs[1]));
    assign layer0_outputs[4723] = (inputs[37]) | (inputs[18]);
    assign layer0_outputs[4724] = ~((inputs[133]) | (inputs[177]));
    assign layer0_outputs[4725] = (inputs[107]) | (inputs[247]);
    assign layer0_outputs[4726] = ~(inputs[85]);
    assign layer0_outputs[4727] = (inputs[119]) & ~(inputs[0]);
    assign layer0_outputs[4728] = ~((inputs[27]) ^ (inputs[238]));
    assign layer0_outputs[4729] = (inputs[137]) & ~(inputs[11]);
    assign layer0_outputs[4730] = ~(inputs[220]);
    assign layer0_outputs[4731] = ~((inputs[96]) & (inputs[58]));
    assign layer0_outputs[4732] = ~(inputs[151]);
    assign layer0_outputs[4733] = ~(inputs[214]) | (inputs[239]);
    assign layer0_outputs[4734] = 1'b0;
    assign layer0_outputs[4735] = inputs[94];
    assign layer0_outputs[4736] = ~(inputs[230]);
    assign layer0_outputs[4737] = ~((inputs[204]) ^ (inputs[89]));
    assign layer0_outputs[4738] = (inputs[190]) & ~(inputs[48]);
    assign layer0_outputs[4739] = ~(inputs[25]);
    assign layer0_outputs[4740] = (inputs[3]) & ~(inputs[190]);
    assign layer0_outputs[4741] = ~(inputs[56]);
    assign layer0_outputs[4742] = (inputs[124]) & ~(inputs[236]);
    assign layer0_outputs[4743] = (inputs[139]) ^ (inputs[158]);
    assign layer0_outputs[4744] = 1'b0;
    assign layer0_outputs[4745] = ~((inputs[227]) | (inputs[250]));
    assign layer0_outputs[4746] = (inputs[146]) | (inputs[145]);
    assign layer0_outputs[4747] = ~(inputs[65]) | (inputs[73]);
    assign layer0_outputs[4748] = inputs[62];
    assign layer0_outputs[4749] = (inputs[236]) ^ (inputs[220]);
    assign layer0_outputs[4750] = inputs[147];
    assign layer0_outputs[4751] = (inputs[191]) | (inputs[212]);
    assign layer0_outputs[4752] = ~(inputs[182]) | (inputs[54]);
    assign layer0_outputs[4753] = (inputs[31]) | (inputs[30]);
    assign layer0_outputs[4754] = ~((inputs[142]) & (inputs[113]));
    assign layer0_outputs[4755] = (inputs[101]) & ~(inputs[61]);
    assign layer0_outputs[4756] = (inputs[85]) & ~(inputs[124]);
    assign layer0_outputs[4757] = (inputs[152]) ^ (inputs[232]);
    assign layer0_outputs[4758] = ~(inputs[231]) | (inputs[205]);
    assign layer0_outputs[4759] = (inputs[248]) | (inputs[34]);
    assign layer0_outputs[4760] = inputs[102];
    assign layer0_outputs[4761] = inputs[201];
    assign layer0_outputs[4762] = ~((inputs[223]) | (inputs[249]));
    assign layer0_outputs[4763] = inputs[88];
    assign layer0_outputs[4764] = (inputs[196]) & ~(inputs[255]);
    assign layer0_outputs[4765] = inputs[188];
    assign layer0_outputs[4766] = (inputs[215]) ^ (inputs[122]);
    assign layer0_outputs[4767] = ~(inputs[245]) | (inputs[151]);
    assign layer0_outputs[4768] = inputs[236];
    assign layer0_outputs[4769] = ~((inputs[158]) & (inputs[37]));
    assign layer0_outputs[4770] = ~(inputs[122]) | (inputs[175]);
    assign layer0_outputs[4771] = ~(inputs[32]) | (inputs[222]);
    assign layer0_outputs[4772] = inputs[210];
    assign layer0_outputs[4773] = ~((inputs[203]) ^ (inputs[169]));
    assign layer0_outputs[4774] = (inputs[102]) ^ (inputs[131]);
    assign layer0_outputs[4775] = ~((inputs[75]) & (inputs[59]));
    assign layer0_outputs[4776] = ~((inputs[251]) & (inputs[46]));
    assign layer0_outputs[4777] = ~(inputs[205]);
    assign layer0_outputs[4778] = ~(inputs[231]) | (inputs[33]);
    assign layer0_outputs[4779] = ~((inputs[57]) & (inputs[6]));
    assign layer0_outputs[4780] = (inputs[157]) ^ (inputs[5]);
    assign layer0_outputs[4781] = (inputs[170]) ^ (inputs[181]);
    assign layer0_outputs[4782] = ~((inputs[48]) | (inputs[89]));
    assign layer0_outputs[4783] = ~((inputs[164]) ^ (inputs[157]));
    assign layer0_outputs[4784] = inputs[218];
    assign layer0_outputs[4785] = ~(inputs[229]);
    assign layer0_outputs[4786] = inputs[234];
    assign layer0_outputs[4787] = (inputs[98]) | (inputs[156]);
    assign layer0_outputs[4788] = ~(inputs[117]);
    assign layer0_outputs[4789] = ~((inputs[2]) | (inputs[4]));
    assign layer0_outputs[4790] = ~(inputs[35]);
    assign layer0_outputs[4791] = (inputs[109]) & ~(inputs[223]);
    assign layer0_outputs[4792] = (inputs[192]) | (inputs[134]);
    assign layer0_outputs[4793] = ~((inputs[177]) | (inputs[100]));
    assign layer0_outputs[4794] = (inputs[236]) & ~(inputs[94]);
    assign layer0_outputs[4795] = ~((inputs[4]) | (inputs[68]));
    assign layer0_outputs[4796] = ~((inputs[212]) | (inputs[128]));
    assign layer0_outputs[4797] = 1'b1;
    assign layer0_outputs[4798] = inputs[63];
    assign layer0_outputs[4799] = (inputs[191]) ^ (inputs[99]);
    assign layer0_outputs[4800] = ~(inputs[217]);
    assign layer0_outputs[4801] = inputs[133];
    assign layer0_outputs[4802] = ~((inputs[64]) ^ (inputs[55]));
    assign layer0_outputs[4803] = ~(inputs[197]) | (inputs[238]);
    assign layer0_outputs[4804] = inputs[134];
    assign layer0_outputs[4805] = (inputs[118]) & (inputs[138]);
    assign layer0_outputs[4806] = 1'b1;
    assign layer0_outputs[4807] = (inputs[227]) | (inputs[97]);
    assign layer0_outputs[4808] = ~((inputs[143]) | (inputs[69]));
    assign layer0_outputs[4809] = ~((inputs[39]) | (inputs[194]));
    assign layer0_outputs[4810] = ~((inputs[128]) & (inputs[79]));
    assign layer0_outputs[4811] = ~((inputs[2]) ^ (inputs[132]));
    assign layer0_outputs[4812] = ~(inputs[54]) | (inputs[12]);
    assign layer0_outputs[4813] = ~(inputs[121]) | (inputs[197]);
    assign layer0_outputs[4814] = (inputs[174]) & ~(inputs[30]);
    assign layer0_outputs[4815] = ~(inputs[211]) | (inputs[57]);
    assign layer0_outputs[4816] = ~(inputs[47]) | (inputs[160]);
    assign layer0_outputs[4817] = (inputs[123]) ^ (inputs[90]);
    assign layer0_outputs[4818] = (inputs[17]) | (inputs[32]);
    assign layer0_outputs[4819] = (inputs[25]) | (inputs[110]);
    assign layer0_outputs[4820] = ~((inputs[13]) | (inputs[16]));
    assign layer0_outputs[4821] = inputs[59];
    assign layer0_outputs[4822] = inputs[109];
    assign layer0_outputs[4823] = ~(inputs[53]);
    assign layer0_outputs[4824] = ~((inputs[225]) | (inputs[37]));
    assign layer0_outputs[4825] = inputs[177];
    assign layer0_outputs[4826] = ~(inputs[31]) | (inputs[198]);
    assign layer0_outputs[4827] = ~(inputs[202]);
    assign layer0_outputs[4828] = ~(inputs[162]);
    assign layer0_outputs[4829] = (inputs[56]) & ~(inputs[208]);
    assign layer0_outputs[4830] = ~(inputs[196]);
    assign layer0_outputs[4831] = (inputs[73]) | (inputs[18]);
    assign layer0_outputs[4832] = 1'b0;
    assign layer0_outputs[4833] = ~(inputs[150]) | (inputs[183]);
    assign layer0_outputs[4834] = ~(inputs[204]);
    assign layer0_outputs[4835] = (inputs[122]) | (inputs[150]);
    assign layer0_outputs[4836] = (inputs[15]) & ~(inputs[157]);
    assign layer0_outputs[4837] = inputs[104];
    assign layer0_outputs[4838] = ~((inputs[111]) | (inputs[104]));
    assign layer0_outputs[4839] = (inputs[85]) ^ (inputs[129]);
    assign layer0_outputs[4840] = inputs[156];
    assign layer0_outputs[4841] = ~((inputs[79]) | (inputs[20]));
    assign layer0_outputs[4842] = (inputs[137]) ^ (inputs[164]);
    assign layer0_outputs[4843] = (inputs[181]) | (inputs[37]);
    assign layer0_outputs[4844] = (inputs[165]) ^ (inputs[29]);
    assign layer0_outputs[4845] = ~(inputs[129]);
    assign layer0_outputs[4846] = 1'b1;
    assign layer0_outputs[4847] = inputs[123];
    assign layer0_outputs[4848] = inputs[91];
    assign layer0_outputs[4849] = (inputs[71]) | (inputs[139]);
    assign layer0_outputs[4850] = (inputs[15]) ^ (inputs[164]);
    assign layer0_outputs[4851] = ~(inputs[109]) | (inputs[222]);
    assign layer0_outputs[4852] = ~((inputs[181]) | (inputs[45]));
    assign layer0_outputs[4853] = inputs[114];
    assign layer0_outputs[4854] = ~((inputs[184]) | (inputs[143]));
    assign layer0_outputs[4855] = (inputs[2]) ^ (inputs[190]);
    assign layer0_outputs[4856] = ~((inputs[135]) ^ (inputs[143]));
    assign layer0_outputs[4857] = ~((inputs[201]) | (inputs[176]));
    assign layer0_outputs[4858] = (inputs[239]) ^ (inputs[84]);
    assign layer0_outputs[4859] = ~(inputs[172]);
    assign layer0_outputs[4860] = ~(inputs[38]);
    assign layer0_outputs[4861] = (inputs[204]) & ~(inputs[110]);
    assign layer0_outputs[4862] = ~(inputs[201]) | (inputs[128]);
    assign layer0_outputs[4863] = (inputs[57]) & ~(inputs[68]);
    assign layer0_outputs[4864] = (inputs[200]) & ~(inputs[10]);
    assign layer0_outputs[4865] = (inputs[106]) & ~(inputs[54]);
    assign layer0_outputs[4866] = (inputs[113]) & (inputs[178]);
    assign layer0_outputs[4867] = ~(inputs[119]);
    assign layer0_outputs[4868] = ~((inputs[86]) | (inputs[220]));
    assign layer0_outputs[4869] = ~(inputs[184]);
    assign layer0_outputs[4870] = inputs[67];
    assign layer0_outputs[4871] = ~((inputs[222]) | (inputs[165]));
    assign layer0_outputs[4872] = ~(inputs[209]);
    assign layer0_outputs[4873] = (inputs[33]) & ~(inputs[97]);
    assign layer0_outputs[4874] = inputs[179];
    assign layer0_outputs[4875] = (inputs[218]) & ~(inputs[110]);
    assign layer0_outputs[4876] = (inputs[207]) | (inputs[249]);
    assign layer0_outputs[4877] = ~(inputs[210]);
    assign layer0_outputs[4878] = (inputs[43]) | (inputs[21]);
    assign layer0_outputs[4879] = inputs[76];
    assign layer0_outputs[4880] = 1'b0;
    assign layer0_outputs[4881] = inputs[108];
    assign layer0_outputs[4882] = ~(inputs[230]);
    assign layer0_outputs[4883] = ~((inputs[232]) ^ (inputs[223]));
    assign layer0_outputs[4884] = (inputs[34]) & ~(inputs[127]);
    assign layer0_outputs[4885] = ~((inputs[38]) ^ (inputs[44]));
    assign layer0_outputs[4886] = ~(inputs[225]);
    assign layer0_outputs[4887] = (inputs[132]) & ~(inputs[205]);
    assign layer0_outputs[4888] = inputs[120];
    assign layer0_outputs[4889] = ~(inputs[105]);
    assign layer0_outputs[4890] = ~((inputs[69]) | (inputs[128]));
    assign layer0_outputs[4891] = (inputs[74]) | (inputs[66]);
    assign layer0_outputs[4892] = ~(inputs[192]) | (inputs[65]);
    assign layer0_outputs[4893] = ~(inputs[19]);
    assign layer0_outputs[4894] = ~(inputs[26]) | (inputs[50]);
    assign layer0_outputs[4895] = ~(inputs[217]) | (inputs[126]);
    assign layer0_outputs[4896] = (inputs[38]) ^ (inputs[229]);
    assign layer0_outputs[4897] = (inputs[155]) ^ (inputs[141]);
    assign layer0_outputs[4898] = ~((inputs[194]) ^ (inputs[9]));
    assign layer0_outputs[4899] = (inputs[173]) | (inputs[83]);
    assign layer0_outputs[4900] = (inputs[16]) | (inputs[185]);
    assign layer0_outputs[4901] = ~(inputs[122]) | (inputs[246]);
    assign layer0_outputs[4902] = ~(inputs[140]);
    assign layer0_outputs[4903] = ~(inputs[220]) | (inputs[114]);
    assign layer0_outputs[4904] = ~((inputs[129]) | (inputs[145]));
    assign layer0_outputs[4905] = (inputs[43]) & ~(inputs[171]);
    assign layer0_outputs[4906] = ~(inputs[182]);
    assign layer0_outputs[4907] = (inputs[220]) ^ (inputs[237]);
    assign layer0_outputs[4908] = (inputs[248]) & ~(inputs[255]);
    assign layer0_outputs[4909] = ~(inputs[253]);
    assign layer0_outputs[4910] = ~(inputs[185]);
    assign layer0_outputs[4911] = ~(inputs[162]) | (inputs[104]);
    assign layer0_outputs[4912] = (inputs[6]) ^ (inputs[239]);
    assign layer0_outputs[4913] = (inputs[215]) & ~(inputs[140]);
    assign layer0_outputs[4914] = ~(inputs[130]);
    assign layer0_outputs[4915] = (inputs[217]) ^ (inputs[205]);
    assign layer0_outputs[4916] = inputs[162];
    assign layer0_outputs[4917] = ~((inputs[1]) | (inputs[55]));
    assign layer0_outputs[4918] = inputs[199];
    assign layer0_outputs[4919] = (inputs[154]) | (inputs[144]);
    assign layer0_outputs[4920] = ~(inputs[81]);
    assign layer0_outputs[4921] = ~((inputs[249]) ^ (inputs[202]));
    assign layer0_outputs[4922] = (inputs[134]) | (inputs[80]);
    assign layer0_outputs[4923] = ~((inputs[77]) | (inputs[43]));
    assign layer0_outputs[4924] = (inputs[116]) & ~(inputs[111]);
    assign layer0_outputs[4925] = ~(inputs[175]);
    assign layer0_outputs[4926] = ~(inputs[215]);
    assign layer0_outputs[4927] = ~(inputs[156]) | (inputs[70]);
    assign layer0_outputs[4928] = ~(inputs[58]);
    assign layer0_outputs[4929] = ~(inputs[100]);
    assign layer0_outputs[4930] = ~(inputs[125]);
    assign layer0_outputs[4931] = ~((inputs[184]) ^ (inputs[174]));
    assign layer0_outputs[4932] = 1'b0;
    assign layer0_outputs[4933] = inputs[150];
    assign layer0_outputs[4934] = (inputs[130]) & ~(inputs[80]);
    assign layer0_outputs[4935] = (inputs[221]) & (inputs[42]);
    assign layer0_outputs[4936] = ~(inputs[204]) | (inputs[103]);
    assign layer0_outputs[4937] = ~((inputs[223]) & (inputs[144]));
    assign layer0_outputs[4938] = (inputs[121]) & ~(inputs[145]);
    assign layer0_outputs[4939] = ~((inputs[195]) | (inputs[175]));
    assign layer0_outputs[4940] = (inputs[241]) | (inputs[120]);
    assign layer0_outputs[4941] = (inputs[86]) ^ (inputs[44]);
    assign layer0_outputs[4942] = (inputs[121]) & ~(inputs[191]);
    assign layer0_outputs[4943] = inputs[209];
    assign layer0_outputs[4944] = (inputs[183]) | (inputs[66]);
    assign layer0_outputs[4945] = inputs[45];
    assign layer0_outputs[4946] = (inputs[166]) & ~(inputs[3]);
    assign layer0_outputs[4947] = ~((inputs[50]) & (inputs[132]));
    assign layer0_outputs[4948] = (inputs[202]) & (inputs[244]);
    assign layer0_outputs[4949] = ~(inputs[129]);
    assign layer0_outputs[4950] = (inputs[79]) & ~(inputs[6]);
    assign layer0_outputs[4951] = (inputs[169]) & ~(inputs[221]);
    assign layer0_outputs[4952] = ~(inputs[91]);
    assign layer0_outputs[4953] = inputs[25];
    assign layer0_outputs[4954] = (inputs[11]) ^ (inputs[72]);
    assign layer0_outputs[4955] = (inputs[244]) & ~(inputs[206]);
    assign layer0_outputs[4956] = ~((inputs[180]) | (inputs[38]));
    assign layer0_outputs[4957] = ~((inputs[38]) | (inputs[158]));
    assign layer0_outputs[4958] = ~(inputs[249]) | (inputs[62]);
    assign layer0_outputs[4959] = ~(inputs[120]) | (inputs[171]);
    assign layer0_outputs[4960] = inputs[24];
    assign layer0_outputs[4961] = ~((inputs[214]) | (inputs[160]));
    assign layer0_outputs[4962] = ~((inputs[158]) | (inputs[77]));
    assign layer0_outputs[4963] = (inputs[104]) & ~(inputs[66]);
    assign layer0_outputs[4964] = (inputs[208]) ^ (inputs[179]);
    assign layer0_outputs[4965] = ~(inputs[208]);
    assign layer0_outputs[4966] = (inputs[90]) | (inputs[51]);
    assign layer0_outputs[4967] = (inputs[177]) | (inputs[192]);
    assign layer0_outputs[4968] = ~(inputs[230]) | (inputs[75]);
    assign layer0_outputs[4969] = ~((inputs[27]) | (inputs[52]));
    assign layer0_outputs[4970] = ~(inputs[91]);
    assign layer0_outputs[4971] = ~(inputs[35]);
    assign layer0_outputs[4972] = ~(inputs[75]) | (inputs[18]);
    assign layer0_outputs[4973] = inputs[20];
    assign layer0_outputs[4974] = (inputs[132]) | (inputs[82]);
    assign layer0_outputs[4975] = (inputs[108]) ^ (inputs[66]);
    assign layer0_outputs[4976] = ~(inputs[236]);
    assign layer0_outputs[4977] = inputs[195];
    assign layer0_outputs[4978] = inputs[45];
    assign layer0_outputs[4979] = (inputs[82]) | (inputs[155]);
    assign layer0_outputs[4980] = (inputs[131]) & (inputs[208]);
    assign layer0_outputs[4981] = ~(inputs[28]);
    assign layer0_outputs[4982] = (inputs[104]) | (inputs[129]);
    assign layer0_outputs[4983] = ~((inputs[251]) | (inputs[118]));
    assign layer0_outputs[4984] = (inputs[86]) & ~(inputs[254]);
    assign layer0_outputs[4985] = (inputs[155]) | (inputs[43]);
    assign layer0_outputs[4986] = inputs[16];
    assign layer0_outputs[4987] = ~((inputs[249]) | (inputs[126]));
    assign layer0_outputs[4988] = ~((inputs[109]) ^ (inputs[106]));
    assign layer0_outputs[4989] = ~(inputs[12]);
    assign layer0_outputs[4990] = (inputs[140]) | (inputs[242]);
    assign layer0_outputs[4991] = (inputs[85]) ^ (inputs[207]);
    assign layer0_outputs[4992] = ~(inputs[53]);
    assign layer0_outputs[4993] = (inputs[229]) & ~(inputs[208]);
    assign layer0_outputs[4994] = ~(inputs[71]) | (inputs[142]);
    assign layer0_outputs[4995] = inputs[36];
    assign layer0_outputs[4996] = (inputs[69]) & ~(inputs[230]);
    assign layer0_outputs[4997] = ~(inputs[69]) | (inputs[196]);
    assign layer0_outputs[4998] = ~((inputs[191]) | (inputs[111]));
    assign layer0_outputs[4999] = ~((inputs[83]) | (inputs[65]));
    assign layer0_outputs[5000] = (inputs[138]) ^ (inputs[153]);
    assign layer0_outputs[5001] = ~(inputs[220]);
    assign layer0_outputs[5002] = (inputs[98]) & ~(inputs[19]);
    assign layer0_outputs[5003] = ~(inputs[104]);
    assign layer0_outputs[5004] = (inputs[88]) & ~(inputs[63]);
    assign layer0_outputs[5005] = (inputs[149]) | (inputs[234]);
    assign layer0_outputs[5006] = (inputs[61]) & ~(inputs[16]);
    assign layer0_outputs[5007] = inputs[209];
    assign layer0_outputs[5008] = inputs[149];
    assign layer0_outputs[5009] = ~(inputs[214]);
    assign layer0_outputs[5010] = ~(inputs[86]);
    assign layer0_outputs[5011] = 1'b1;
    assign layer0_outputs[5012] = (inputs[36]) & ~(inputs[127]);
    assign layer0_outputs[5013] = (inputs[171]) & (inputs[183]);
    assign layer0_outputs[5014] = ~(inputs[179]);
    assign layer0_outputs[5015] = inputs[164];
    assign layer0_outputs[5016] = (inputs[233]) & ~(inputs[28]);
    assign layer0_outputs[5017] = ~((inputs[177]) ^ (inputs[226]));
    assign layer0_outputs[5018] = ~(inputs[103]);
    assign layer0_outputs[5019] = (inputs[82]) & (inputs[114]);
    assign layer0_outputs[5020] = inputs[3];
    assign layer0_outputs[5021] = ~((inputs[130]) ^ (inputs[107]));
    assign layer0_outputs[5022] = (inputs[201]) & (inputs[236]);
    assign layer0_outputs[5023] = ~((inputs[5]) ^ (inputs[15]));
    assign layer0_outputs[5024] = (inputs[234]) & (inputs[229]);
    assign layer0_outputs[5025] = (inputs[4]) | (inputs[227]);
    assign layer0_outputs[5026] = ~((inputs[143]) | (inputs[68]));
    assign layer0_outputs[5027] = ~((inputs[61]) ^ (inputs[28]));
    assign layer0_outputs[5028] = ~(inputs[72]) | (inputs[126]);
    assign layer0_outputs[5029] = ~((inputs[213]) | (inputs[62]));
    assign layer0_outputs[5030] = ~(inputs[196]);
    assign layer0_outputs[5031] = (inputs[185]) & (inputs[188]);
    assign layer0_outputs[5032] = (inputs[242]) ^ (inputs[65]);
    assign layer0_outputs[5033] = ~((inputs[25]) ^ (inputs[43]));
    assign layer0_outputs[5034] = ~(inputs[104]) | (inputs[14]);
    assign layer0_outputs[5035] = ~(inputs[247]) | (inputs[110]);
    assign layer0_outputs[5036] = ~((inputs[102]) | (inputs[133]));
    assign layer0_outputs[5037] = inputs[106];
    assign layer0_outputs[5038] = ~(inputs[205]);
    assign layer0_outputs[5039] = ~(inputs[20]);
    assign layer0_outputs[5040] = inputs[246];
    assign layer0_outputs[5041] = (inputs[186]) & ~(inputs[108]);
    assign layer0_outputs[5042] = inputs[208];
    assign layer0_outputs[5043] = ~(inputs[247]);
    assign layer0_outputs[5044] = (inputs[201]) ^ (inputs[247]);
    assign layer0_outputs[5045] = ~(inputs[243]) | (inputs[105]);
    assign layer0_outputs[5046] = (inputs[167]) & (inputs[160]);
    assign layer0_outputs[5047] = ~(inputs[195]);
    assign layer0_outputs[5048] = inputs[27];
    assign layer0_outputs[5049] = (inputs[75]) ^ (inputs[177]);
    assign layer0_outputs[5050] = ~(inputs[32]);
    assign layer0_outputs[5051] = ~((inputs[234]) ^ (inputs[162]));
    assign layer0_outputs[5052] = ~(inputs[121]) | (inputs[192]);
    assign layer0_outputs[5053] = inputs[100];
    assign layer0_outputs[5054] = (inputs[127]) ^ (inputs[152]);
    assign layer0_outputs[5055] = ~((inputs[13]) ^ (inputs[176]));
    assign layer0_outputs[5056] = ~((inputs[25]) | (inputs[112]));
    assign layer0_outputs[5057] = inputs[229];
    assign layer0_outputs[5058] = ~(inputs[74]);
    assign layer0_outputs[5059] = (inputs[52]) & ~(inputs[32]);
    assign layer0_outputs[5060] = ~((inputs[150]) & (inputs[183]));
    assign layer0_outputs[5061] = (inputs[70]) & ~(inputs[106]);
    assign layer0_outputs[5062] = (inputs[231]) & (inputs[134]);
    assign layer0_outputs[5063] = (inputs[151]) & ~(inputs[100]);
    assign layer0_outputs[5064] = (inputs[215]) ^ (inputs[153]);
    assign layer0_outputs[5065] = ~(inputs[151]) | (inputs[215]);
    assign layer0_outputs[5066] = ~(inputs[35]) | (inputs[128]);
    assign layer0_outputs[5067] = (inputs[113]) & ~(inputs[27]);
    assign layer0_outputs[5068] = inputs[92];
    assign layer0_outputs[5069] = ~(inputs[123]) | (inputs[208]);
    assign layer0_outputs[5070] = ~((inputs[158]) | (inputs[16]));
    assign layer0_outputs[5071] = (inputs[201]) | (inputs[157]);
    assign layer0_outputs[5072] = inputs[210];
    assign layer0_outputs[5073] = ~((inputs[248]) | (inputs[142]));
    assign layer0_outputs[5074] = inputs[55];
    assign layer0_outputs[5075] = (inputs[129]) ^ (inputs[101]);
    assign layer0_outputs[5076] = ~((inputs[6]) ^ (inputs[205]));
    assign layer0_outputs[5077] = (inputs[37]) & ~(inputs[127]);
    assign layer0_outputs[5078] = ~((inputs[50]) | (inputs[122]));
    assign layer0_outputs[5079] = ~((inputs[14]) | (inputs[96]));
    assign layer0_outputs[5080] = (inputs[105]) ^ (inputs[177]);
    assign layer0_outputs[5081] = ~((inputs[186]) | (inputs[115]));
    assign layer0_outputs[5082] = (inputs[66]) & ~(inputs[143]);
    assign layer0_outputs[5083] = inputs[89];
    assign layer0_outputs[5084] = inputs[142];
    assign layer0_outputs[5085] = inputs[169];
    assign layer0_outputs[5086] = (inputs[161]) & ~(inputs[95]);
    assign layer0_outputs[5087] = inputs[128];
    assign layer0_outputs[5088] = inputs[139];
    assign layer0_outputs[5089] = ~((inputs[238]) | (inputs[227]));
    assign layer0_outputs[5090] = ~(inputs[92]);
    assign layer0_outputs[5091] = (inputs[115]) ^ (inputs[64]);
    assign layer0_outputs[5092] = ~(inputs[116]) | (inputs[104]);
    assign layer0_outputs[5093] = (inputs[217]) & (inputs[0]);
    assign layer0_outputs[5094] = ~(inputs[116]) | (inputs[49]);
    assign layer0_outputs[5095] = ~(inputs[156]);
    assign layer0_outputs[5096] = inputs[69];
    assign layer0_outputs[5097] = inputs[151];
    assign layer0_outputs[5098] = (inputs[112]) ^ (inputs[156]);
    assign layer0_outputs[5099] = ~(inputs[133]) | (inputs[252]);
    assign layer0_outputs[5100] = ~((inputs[93]) | (inputs[178]));
    assign layer0_outputs[5101] = ~((inputs[40]) ^ (inputs[8]));
    assign layer0_outputs[5102] = (inputs[133]) ^ (inputs[8]);
    assign layer0_outputs[5103] = ~((inputs[114]) | (inputs[184]));
    assign layer0_outputs[5104] = ~((inputs[89]) ^ (inputs[43]));
    assign layer0_outputs[5105] = inputs[113];
    assign layer0_outputs[5106] = (inputs[116]) & ~(inputs[16]);
    assign layer0_outputs[5107] = ~(inputs[20]) | (inputs[47]);
    assign layer0_outputs[5108] = (inputs[31]) | (inputs[43]);
    assign layer0_outputs[5109] = inputs[153];
    assign layer0_outputs[5110] = inputs[163];
    assign layer0_outputs[5111] = inputs[41];
    assign layer0_outputs[5112] = ~((inputs[164]) | (inputs[226]));
    assign layer0_outputs[5113] = inputs[58];
    assign layer0_outputs[5114] = (inputs[54]) ^ (inputs[64]);
    assign layer0_outputs[5115] = ~(inputs[129]);
    assign layer0_outputs[5116] = ~((inputs[219]) | (inputs[96]));
    assign layer0_outputs[5117] = (inputs[198]) & ~(inputs[88]);
    assign layer0_outputs[5118] = ~(inputs[231]);
    assign layer0_outputs[5119] = ~((inputs[134]) ^ (inputs[182]));
    assign layer0_outputs[5120] = ~(inputs[178]);
    assign layer0_outputs[5121] = (inputs[82]) | (inputs[90]);
    assign layer0_outputs[5122] = ~(inputs[231]);
    assign layer0_outputs[5123] = (inputs[42]) & ~(inputs[0]);
    assign layer0_outputs[5124] = ~(inputs[178]);
    assign layer0_outputs[5125] = (inputs[23]) ^ (inputs[160]);
    assign layer0_outputs[5126] = ~(inputs[152]);
    assign layer0_outputs[5127] = 1'b1;
    assign layer0_outputs[5128] = (inputs[165]) & ~(inputs[96]);
    assign layer0_outputs[5129] = ~(inputs[100]) | (inputs[49]);
    assign layer0_outputs[5130] = inputs[137];
    assign layer0_outputs[5131] = (inputs[9]) | (inputs[179]);
    assign layer0_outputs[5132] = ~((inputs[187]) ^ (inputs[137]));
    assign layer0_outputs[5133] = ~((inputs[58]) & (inputs[245]));
    assign layer0_outputs[5134] = (inputs[66]) | (inputs[164]);
    assign layer0_outputs[5135] = inputs[233];
    assign layer0_outputs[5136] = (inputs[27]) ^ (inputs[131]);
    assign layer0_outputs[5137] = ~(inputs[20]);
    assign layer0_outputs[5138] = 1'b1;
    assign layer0_outputs[5139] = (inputs[98]) ^ (inputs[84]);
    assign layer0_outputs[5140] = ~(inputs[208]);
    assign layer0_outputs[5141] = inputs[153];
    assign layer0_outputs[5142] = inputs[130];
    assign layer0_outputs[5143] = ~(inputs[231]) | (inputs[238]);
    assign layer0_outputs[5144] = (inputs[148]) ^ (inputs[136]);
    assign layer0_outputs[5145] = ~(inputs[103]);
    assign layer0_outputs[5146] = (inputs[77]) | (inputs[23]);
    assign layer0_outputs[5147] = (inputs[166]) & (inputs[187]);
    assign layer0_outputs[5148] = ~(inputs[88]);
    assign layer0_outputs[5149] = (inputs[84]) & ~(inputs[204]);
    assign layer0_outputs[5150] = (inputs[86]) ^ (inputs[99]);
    assign layer0_outputs[5151] = ~(inputs[81]);
    assign layer0_outputs[5152] = ~((inputs[91]) ^ (inputs[164]));
    assign layer0_outputs[5153] = ~(inputs[130]);
    assign layer0_outputs[5154] = inputs[73];
    assign layer0_outputs[5155] = inputs[7];
    assign layer0_outputs[5156] = (inputs[48]) | (inputs[202]);
    assign layer0_outputs[5157] = ~(inputs[25]);
    assign layer0_outputs[5158] = ~(inputs[181]);
    assign layer0_outputs[5159] = ~((inputs[26]) ^ (inputs[41]));
    assign layer0_outputs[5160] = (inputs[137]) ^ (inputs[167]);
    assign layer0_outputs[5161] = ~(inputs[84]) | (inputs[177]);
    assign layer0_outputs[5162] = ~(inputs[148]);
    assign layer0_outputs[5163] = (inputs[135]) & (inputs[235]);
    assign layer0_outputs[5164] = ~((inputs[186]) | (inputs[215]));
    assign layer0_outputs[5165] = inputs[19];
    assign layer0_outputs[5166] = ~(inputs[119]) | (inputs[173]);
    assign layer0_outputs[5167] = ~(inputs[186]) | (inputs[47]);
    assign layer0_outputs[5168] = ~((inputs[160]) | (inputs[170]));
    assign layer0_outputs[5169] = ~(inputs[131]) | (inputs[49]);
    assign layer0_outputs[5170] = (inputs[166]) | (inputs[154]);
    assign layer0_outputs[5171] = (inputs[63]) | (inputs[35]);
    assign layer0_outputs[5172] = ~(inputs[198]) | (inputs[11]);
    assign layer0_outputs[5173] = ~((inputs[206]) | (inputs[213]));
    assign layer0_outputs[5174] = ~(inputs[164]);
    assign layer0_outputs[5175] = ~((inputs[250]) ^ (inputs[55]));
    assign layer0_outputs[5176] = inputs[101];
    assign layer0_outputs[5177] = ~(inputs[230]);
    assign layer0_outputs[5178] = ~((inputs[30]) | (inputs[128]));
    assign layer0_outputs[5179] = inputs[99];
    assign layer0_outputs[5180] = inputs[15];
    assign layer0_outputs[5181] = (inputs[131]) | (inputs[54]);
    assign layer0_outputs[5182] = ~((inputs[243]) ^ (inputs[22]));
    assign layer0_outputs[5183] = inputs[194];
    assign layer0_outputs[5184] = ~(inputs[53]);
    assign layer0_outputs[5185] = ~((inputs[147]) & (inputs[139]));
    assign layer0_outputs[5186] = inputs[196];
    assign layer0_outputs[5187] = (inputs[39]) & ~(inputs[230]);
    assign layer0_outputs[5188] = ~((inputs[182]) | (inputs[245]));
    assign layer0_outputs[5189] = (inputs[104]) ^ (inputs[193]);
    assign layer0_outputs[5190] = 1'b1;
    assign layer0_outputs[5191] = inputs[52];
    assign layer0_outputs[5192] = (inputs[156]) ^ (inputs[4]);
    assign layer0_outputs[5193] = ~(inputs[217]);
    assign layer0_outputs[5194] = ~((inputs[164]) | (inputs[252]));
    assign layer0_outputs[5195] = ~((inputs[247]) | (inputs[174]));
    assign layer0_outputs[5196] = (inputs[189]) & ~(inputs[161]);
    assign layer0_outputs[5197] = ~(inputs[192]);
    assign layer0_outputs[5198] = (inputs[27]) & ~(inputs[166]);
    assign layer0_outputs[5199] = inputs[104];
    assign layer0_outputs[5200] = (inputs[210]) & ~(inputs[96]);
    assign layer0_outputs[5201] = ~(inputs[26]) | (inputs[112]);
    assign layer0_outputs[5202] = ~(inputs[119]);
    assign layer0_outputs[5203] = ~((inputs[36]) | (inputs[91]));
    assign layer0_outputs[5204] = (inputs[59]) ^ (inputs[73]);
    assign layer0_outputs[5205] = (inputs[216]) ^ (inputs[195]);
    assign layer0_outputs[5206] = ~(inputs[249]) | (inputs[54]);
    assign layer0_outputs[5207] = ~(inputs[54]) | (inputs[144]);
    assign layer0_outputs[5208] = inputs[75];
    assign layer0_outputs[5209] = ~(inputs[53]) | (inputs[205]);
    assign layer0_outputs[5210] = ~(inputs[20]);
    assign layer0_outputs[5211] = (inputs[65]) | (inputs[138]);
    assign layer0_outputs[5212] = ~(inputs[105]);
    assign layer0_outputs[5213] = ~(inputs[23]);
    assign layer0_outputs[5214] = ~(inputs[114]);
    assign layer0_outputs[5215] = ~(inputs[154]) | (inputs[27]);
    assign layer0_outputs[5216] = ~(inputs[137]);
    assign layer0_outputs[5217] = ~(inputs[3]) | (inputs[128]);
    assign layer0_outputs[5218] = ~(inputs[7]);
    assign layer0_outputs[5219] = ~(inputs[54]) | (inputs[34]);
    assign layer0_outputs[5220] = ~((inputs[226]) | (inputs[21]));
    assign layer0_outputs[5221] = inputs[129];
    assign layer0_outputs[5222] = ~((inputs[255]) ^ (inputs[163]));
    assign layer0_outputs[5223] = (inputs[209]) | (inputs[118]);
    assign layer0_outputs[5224] = ~(inputs[126]);
    assign layer0_outputs[5225] = ~((inputs[190]) | (inputs[204]));
    assign layer0_outputs[5226] = ~(inputs[145]);
    assign layer0_outputs[5227] = ~(inputs[42]);
    assign layer0_outputs[5228] = (inputs[187]) | (inputs[207]);
    assign layer0_outputs[5229] = ~((inputs[227]) | (inputs[219]));
    assign layer0_outputs[5230] = (inputs[216]) | (inputs[216]);
    assign layer0_outputs[5231] = (inputs[169]) & ~(inputs[50]);
    assign layer0_outputs[5232] = (inputs[209]) | (inputs[237]);
    assign layer0_outputs[5233] = inputs[52];
    assign layer0_outputs[5234] = ~(inputs[207]) | (inputs[223]);
    assign layer0_outputs[5235] = inputs[174];
    assign layer0_outputs[5236] = ~((inputs[204]) ^ (inputs[240]));
    assign layer0_outputs[5237] = 1'b1;
    assign layer0_outputs[5238] = ~((inputs[63]) ^ (inputs[156]));
    assign layer0_outputs[5239] = ~(inputs[152]);
    assign layer0_outputs[5240] = (inputs[231]) & ~(inputs[126]);
    assign layer0_outputs[5241] = ~((inputs[196]) ^ (inputs[27]));
    assign layer0_outputs[5242] = ~((inputs[174]) ^ (inputs[107]));
    assign layer0_outputs[5243] = 1'b1;
    assign layer0_outputs[5244] = ~((inputs[63]) ^ (inputs[199]));
    assign layer0_outputs[5245] = ~(inputs[230]);
    assign layer0_outputs[5246] = ~((inputs[145]) | (inputs[160]));
    assign layer0_outputs[5247] = ~((inputs[204]) ^ (inputs[225]));
    assign layer0_outputs[5248] = ~((inputs[65]) | (inputs[179]));
    assign layer0_outputs[5249] = (inputs[177]) ^ (inputs[144]);
    assign layer0_outputs[5250] = ~(inputs[30]);
    assign layer0_outputs[5251] = ~((inputs[104]) | (inputs[163]));
    assign layer0_outputs[5252] = ~((inputs[196]) ^ (inputs[10]));
    assign layer0_outputs[5253] = ~(inputs[57]) | (inputs[149]);
    assign layer0_outputs[5254] = (inputs[68]) ^ (inputs[133]);
    assign layer0_outputs[5255] = ~((inputs[21]) | (inputs[43]));
    assign layer0_outputs[5256] = (inputs[37]) & ~(inputs[223]);
    assign layer0_outputs[5257] = (inputs[6]) & ~(inputs[199]);
    assign layer0_outputs[5258] = (inputs[247]) | (inputs[88]);
    assign layer0_outputs[5259] = inputs[113];
    assign layer0_outputs[5260] = ~((inputs[63]) | (inputs[247]));
    assign layer0_outputs[5261] = (inputs[176]) ^ (inputs[190]);
    assign layer0_outputs[5262] = ~((inputs[148]) | (inputs[141]));
    assign layer0_outputs[5263] = inputs[205];
    assign layer0_outputs[5264] = (inputs[52]) & ~(inputs[250]);
    assign layer0_outputs[5265] = ~(inputs[194]);
    assign layer0_outputs[5266] = (inputs[4]) ^ (inputs[176]);
    assign layer0_outputs[5267] = (inputs[0]) & ~(inputs[155]);
    assign layer0_outputs[5268] = (inputs[105]) | (inputs[243]);
    assign layer0_outputs[5269] = ~(inputs[176]);
    assign layer0_outputs[5270] = (inputs[169]) | (inputs[237]);
    assign layer0_outputs[5271] = ~((inputs[229]) | (inputs[182]));
    assign layer0_outputs[5272] = ~((inputs[187]) ^ (inputs[149]));
    assign layer0_outputs[5273] = ~(inputs[93]);
    assign layer0_outputs[5274] = inputs[57];
    assign layer0_outputs[5275] = ~(inputs[17]) | (inputs[11]);
    assign layer0_outputs[5276] = (inputs[117]) | (inputs[163]);
    assign layer0_outputs[5277] = ~(inputs[46]) | (inputs[208]);
    assign layer0_outputs[5278] = inputs[39];
    assign layer0_outputs[5279] = ~((inputs[53]) ^ (inputs[114]));
    assign layer0_outputs[5280] = ~(inputs[19]);
    assign layer0_outputs[5281] = inputs[61];
    assign layer0_outputs[5282] = inputs[103];
    assign layer0_outputs[5283] = (inputs[107]) ^ (inputs[90]);
    assign layer0_outputs[5284] = ~((inputs[161]) | (inputs[17]));
    assign layer0_outputs[5285] = ~(inputs[100]) | (inputs[47]);
    assign layer0_outputs[5286] = (inputs[254]) | (inputs[252]);
    assign layer0_outputs[5287] = ~((inputs[196]) | (inputs[80]));
    assign layer0_outputs[5288] = ~((inputs[159]) ^ (inputs[31]));
    assign layer0_outputs[5289] = ~(inputs[138]);
    assign layer0_outputs[5290] = (inputs[68]) & ~(inputs[220]);
    assign layer0_outputs[5291] = ~(inputs[183]);
    assign layer0_outputs[5292] = ~(inputs[181]) | (inputs[237]);
    assign layer0_outputs[5293] = ~(inputs[227]);
    assign layer0_outputs[5294] = (inputs[245]) | (inputs[175]);
    assign layer0_outputs[5295] = (inputs[31]) & (inputs[84]);
    assign layer0_outputs[5296] = ~(inputs[34]);
    assign layer0_outputs[5297] = ~(inputs[175]);
    assign layer0_outputs[5298] = ~((inputs[24]) | (inputs[127]));
    assign layer0_outputs[5299] = ~((inputs[197]) | (inputs[14]));
    assign layer0_outputs[5300] = inputs[98];
    assign layer0_outputs[5301] = (inputs[35]) | (inputs[140]);
    assign layer0_outputs[5302] = inputs[57];
    assign layer0_outputs[5303] = ~(inputs[210]);
    assign layer0_outputs[5304] = ~(inputs[5]) | (inputs[225]);
    assign layer0_outputs[5305] = ~(inputs[139]) | (inputs[248]);
    assign layer0_outputs[5306] = ~(inputs[220]);
    assign layer0_outputs[5307] = (inputs[103]) & ~(inputs[146]);
    assign layer0_outputs[5308] = ~((inputs[177]) & (inputs[210]));
    assign layer0_outputs[5309] = inputs[99];
    assign layer0_outputs[5310] = (inputs[55]) | (inputs[139]);
    assign layer0_outputs[5311] = ~(inputs[152]) | (inputs[55]);
    assign layer0_outputs[5312] = (inputs[230]) & (inputs[170]);
    assign layer0_outputs[5313] = ~((inputs[224]) ^ (inputs[12]));
    assign layer0_outputs[5314] = ~((inputs[141]) | (inputs[144]));
    assign layer0_outputs[5315] = (inputs[62]) | (inputs[42]);
    assign layer0_outputs[5316] = ~(inputs[184]);
    assign layer0_outputs[5317] = ~(inputs[106]);
    assign layer0_outputs[5318] = inputs[209];
    assign layer0_outputs[5319] = ~(inputs[164]) | (inputs[50]);
    assign layer0_outputs[5320] = (inputs[48]) | (inputs[191]);
    assign layer0_outputs[5321] = ~(inputs[90]) | (inputs[95]);
    assign layer0_outputs[5322] = ~(inputs[253]) | (inputs[81]);
    assign layer0_outputs[5323] = (inputs[78]) & ~(inputs[162]);
    assign layer0_outputs[5324] = ~((inputs[144]) | (inputs[83]));
    assign layer0_outputs[5325] = ~((inputs[123]) | (inputs[70]));
    assign layer0_outputs[5326] = (inputs[249]) | (inputs[1]);
    assign layer0_outputs[5327] = ~(inputs[91]);
    assign layer0_outputs[5328] = (inputs[27]) & ~(inputs[149]);
    assign layer0_outputs[5329] = (inputs[68]) ^ (inputs[105]);
    assign layer0_outputs[5330] = inputs[40];
    assign layer0_outputs[5331] = ~(inputs[201]) | (inputs[25]);
    assign layer0_outputs[5332] = ~((inputs[78]) & (inputs[79]));
    assign layer0_outputs[5333] = ~(inputs[38]) | (inputs[139]);
    assign layer0_outputs[5334] = ~(inputs[95]);
    assign layer0_outputs[5335] = ~((inputs[220]) ^ (inputs[161]));
    assign layer0_outputs[5336] = (inputs[77]) & ~(inputs[49]);
    assign layer0_outputs[5337] = inputs[118];
    assign layer0_outputs[5338] = ~(inputs[149]);
    assign layer0_outputs[5339] = inputs[123];
    assign layer0_outputs[5340] = ~(inputs[99]);
    assign layer0_outputs[5341] = inputs[109];
    assign layer0_outputs[5342] = (inputs[201]) | (inputs[137]);
    assign layer0_outputs[5343] = ~(inputs[41]);
    assign layer0_outputs[5344] = ~((inputs[125]) ^ (inputs[240]));
    assign layer0_outputs[5345] = (inputs[42]) | (inputs[2]);
    assign layer0_outputs[5346] = ~((inputs[161]) | (inputs[29]));
    assign layer0_outputs[5347] = ~(inputs[186]) | (inputs[120]);
    assign layer0_outputs[5348] = inputs[86];
    assign layer0_outputs[5349] = inputs[99];
    assign layer0_outputs[5350] = (inputs[88]) | (inputs[194]);
    assign layer0_outputs[5351] = (inputs[185]) | (inputs[235]);
    assign layer0_outputs[5352] = (inputs[7]) & ~(inputs[86]);
    assign layer0_outputs[5353] = (inputs[23]) & ~(inputs[247]);
    assign layer0_outputs[5354] = inputs[137];
    assign layer0_outputs[5355] = (inputs[61]) | (inputs[5]);
    assign layer0_outputs[5356] = ~(inputs[84]) | (inputs[3]);
    assign layer0_outputs[5357] = ~((inputs[96]) | (inputs[30]));
    assign layer0_outputs[5358] = (inputs[139]) & (inputs[139]);
    assign layer0_outputs[5359] = (inputs[79]) & (inputs[31]);
    assign layer0_outputs[5360] = ~(inputs[77]);
    assign layer0_outputs[5361] = (inputs[26]) & ~(inputs[255]);
    assign layer0_outputs[5362] = ~((inputs[175]) | (inputs[147]));
    assign layer0_outputs[5363] = ~((inputs[78]) ^ (inputs[234]));
    assign layer0_outputs[5364] = ~(inputs[139]) | (inputs[234]);
    assign layer0_outputs[5365] = (inputs[136]) | (inputs[148]);
    assign layer0_outputs[5366] = ~(inputs[244]);
    assign layer0_outputs[5367] = ~(inputs[25]);
    assign layer0_outputs[5368] = (inputs[41]) & ~(inputs[48]);
    assign layer0_outputs[5369] = ~(inputs[29]);
    assign layer0_outputs[5370] = ~((inputs[2]) ^ (inputs[141]));
    assign layer0_outputs[5371] = (inputs[102]) | (inputs[215]);
    assign layer0_outputs[5372] = (inputs[217]) ^ (inputs[166]);
    assign layer0_outputs[5373] = (inputs[185]) | (inputs[80]);
    assign layer0_outputs[5374] = (inputs[105]) | (inputs[89]);
    assign layer0_outputs[5375] = ~(inputs[82]);
    assign layer0_outputs[5376] = inputs[111];
    assign layer0_outputs[5377] = inputs[99];
    assign layer0_outputs[5378] = inputs[206];
    assign layer0_outputs[5379] = (inputs[117]) & ~(inputs[205]);
    assign layer0_outputs[5380] = inputs[174];
    assign layer0_outputs[5381] = ~(inputs[94]);
    assign layer0_outputs[5382] = (inputs[56]) & (inputs[244]);
    assign layer0_outputs[5383] = ~(inputs[101]) | (inputs[93]);
    assign layer0_outputs[5384] = ~((inputs[193]) | (inputs[174]));
    assign layer0_outputs[5385] = (inputs[105]) & ~(inputs[49]);
    assign layer0_outputs[5386] = (inputs[161]) | (inputs[146]);
    assign layer0_outputs[5387] = ~(inputs[48]) | (inputs[141]);
    assign layer0_outputs[5388] = ~(inputs[148]);
    assign layer0_outputs[5389] = inputs[178];
    assign layer0_outputs[5390] = ~(inputs[164]);
    assign layer0_outputs[5391] = ~(inputs[85]);
    assign layer0_outputs[5392] = (inputs[141]) & ~(inputs[92]);
    assign layer0_outputs[5393] = (inputs[207]) | (inputs[58]);
    assign layer0_outputs[5394] = inputs[101];
    assign layer0_outputs[5395] = inputs[144];
    assign layer0_outputs[5396] = (inputs[11]) ^ (inputs[51]);
    assign layer0_outputs[5397] = ~(inputs[18]);
    assign layer0_outputs[5398] = ~(inputs[17]) | (inputs[238]);
    assign layer0_outputs[5399] = ~((inputs[229]) | (inputs[191]));
    assign layer0_outputs[5400] = ~((inputs[66]) | (inputs[112]));
    assign layer0_outputs[5401] = ~((inputs[28]) | (inputs[34]));
    assign layer0_outputs[5402] = (inputs[164]) | (inputs[86]);
    assign layer0_outputs[5403] = (inputs[211]) | (inputs[189]);
    assign layer0_outputs[5404] = ~((inputs[95]) | (inputs[84]));
    assign layer0_outputs[5405] = ~(inputs[101]);
    assign layer0_outputs[5406] = inputs[239];
    assign layer0_outputs[5407] = ~((inputs[49]) | (inputs[63]));
    assign layer0_outputs[5408] = (inputs[224]) & ~(inputs[88]);
    assign layer0_outputs[5409] = ~((inputs[83]) ^ (inputs[71]));
    assign layer0_outputs[5410] = (inputs[0]) | (inputs[128]);
    assign layer0_outputs[5411] = (inputs[247]) ^ (inputs[62]);
    assign layer0_outputs[5412] = ~((inputs[226]) & (inputs[95]));
    assign layer0_outputs[5413] = (inputs[163]) & ~(inputs[16]);
    assign layer0_outputs[5414] = ~((inputs[253]) | (inputs[189]));
    assign layer0_outputs[5415] = ~((inputs[64]) | (inputs[255]));
    assign layer0_outputs[5416] = inputs[121];
    assign layer0_outputs[5417] = ~((inputs[53]) ^ (inputs[121]));
    assign layer0_outputs[5418] = inputs[88];
    assign layer0_outputs[5419] = inputs[76];
    assign layer0_outputs[5420] = ~((inputs[20]) ^ (inputs[107]));
    assign layer0_outputs[5421] = ~(inputs[177]) | (inputs[43]);
    assign layer0_outputs[5422] = (inputs[85]) & ~(inputs[156]);
    assign layer0_outputs[5423] = ~(inputs[182]) | (inputs[45]);
    assign layer0_outputs[5424] = (inputs[220]) ^ (inputs[1]);
    assign layer0_outputs[5425] = ~(inputs[75]);
    assign layer0_outputs[5426] = ~((inputs[201]) | (inputs[218]));
    assign layer0_outputs[5427] = inputs[73];
    assign layer0_outputs[5428] = (inputs[237]) | (inputs[149]);
    assign layer0_outputs[5429] = (inputs[141]) & ~(inputs[37]);
    assign layer0_outputs[5430] = (inputs[193]) | (inputs[218]);
    assign layer0_outputs[5431] = (inputs[37]) & ~(inputs[250]);
    assign layer0_outputs[5432] = inputs[105];
    assign layer0_outputs[5433] = inputs[110];
    assign layer0_outputs[5434] = (inputs[61]) & ~(inputs[113]);
    assign layer0_outputs[5435] = ~(inputs[255]) | (inputs[16]);
    assign layer0_outputs[5436] = ~(inputs[246]) | (inputs[127]);
    assign layer0_outputs[5437] = 1'b0;
    assign layer0_outputs[5438] = inputs[180];
    assign layer0_outputs[5439] = ~(inputs[197]);
    assign layer0_outputs[5440] = ~((inputs[208]) | (inputs[103]));
    assign layer0_outputs[5441] = (inputs[138]) & ~(inputs[119]);
    assign layer0_outputs[5442] = (inputs[22]) ^ (inputs[34]);
    assign layer0_outputs[5443] = (inputs[183]) & ~(inputs[238]);
    assign layer0_outputs[5444] = ~(inputs[9]) | (inputs[180]);
    assign layer0_outputs[5445] = inputs[129];
    assign layer0_outputs[5446] = (inputs[231]) ^ (inputs[56]);
    assign layer0_outputs[5447] = ~((inputs[51]) | (inputs[107]));
    assign layer0_outputs[5448] = 1'b1;
    assign layer0_outputs[5449] = ~(inputs[179]);
    assign layer0_outputs[5450] = ~(inputs[169]);
    assign layer0_outputs[5451] = inputs[219];
    assign layer0_outputs[5452] = ~((inputs[49]) | (inputs[184]));
    assign layer0_outputs[5453] = ~(inputs[12]);
    assign layer0_outputs[5454] = (inputs[158]) | (inputs[195]);
    assign layer0_outputs[5455] = (inputs[67]) & ~(inputs[203]);
    assign layer0_outputs[5456] = (inputs[202]) & ~(inputs[113]);
    assign layer0_outputs[5457] = ~(inputs[142]) | (inputs[237]);
    assign layer0_outputs[5458] = inputs[205];
    assign layer0_outputs[5459] = (inputs[0]) ^ (inputs[250]);
    assign layer0_outputs[5460] = (inputs[159]) | (inputs[212]);
    assign layer0_outputs[5461] = ~(inputs[13]) | (inputs[111]);
    assign layer0_outputs[5462] = ~(inputs[86]);
    assign layer0_outputs[5463] = (inputs[32]) | (inputs[55]);
    assign layer0_outputs[5464] = ~(inputs[210]);
    assign layer0_outputs[5465] = (inputs[19]) | (inputs[39]);
    assign layer0_outputs[5466] = ~((inputs[68]) & (inputs[133]));
    assign layer0_outputs[5467] = (inputs[86]) ^ (inputs[20]);
    assign layer0_outputs[5468] = inputs[85];
    assign layer0_outputs[5469] = (inputs[209]) | (inputs[48]);
    assign layer0_outputs[5470] = ~((inputs[24]) & (inputs[194]));
    assign layer0_outputs[5471] = ~((inputs[59]) ^ (inputs[14]));
    assign layer0_outputs[5472] = ~((inputs[3]) ^ (inputs[226]));
    assign layer0_outputs[5473] = inputs[132];
    assign layer0_outputs[5474] = (inputs[243]) & (inputs[240]);
    assign layer0_outputs[5475] = (inputs[76]) & ~(inputs[108]);
    assign layer0_outputs[5476] = ~(inputs[57]);
    assign layer0_outputs[5477] = inputs[229];
    assign layer0_outputs[5478] = ~(inputs[232]);
    assign layer0_outputs[5479] = ~(inputs[219]) | (inputs[109]);
    assign layer0_outputs[5480] = inputs[143];
    assign layer0_outputs[5481] = ~(inputs[116]);
    assign layer0_outputs[5482] = ~((inputs[21]) ^ (inputs[35]));
    assign layer0_outputs[5483] = inputs[86];
    assign layer0_outputs[5484] = (inputs[4]) & ~(inputs[62]);
    assign layer0_outputs[5485] = 1'b1;
    assign layer0_outputs[5486] = inputs[166];
    assign layer0_outputs[5487] = inputs[94];
    assign layer0_outputs[5488] = ~(inputs[40]);
    assign layer0_outputs[5489] = ~(inputs[216]);
    assign layer0_outputs[5490] = (inputs[9]) | (inputs[88]);
    assign layer0_outputs[5491] = (inputs[200]) & ~(inputs[84]);
    assign layer0_outputs[5492] = inputs[225];
    assign layer0_outputs[5493] = (inputs[30]) ^ (inputs[61]);
    assign layer0_outputs[5494] = (inputs[214]) | (inputs[56]);
    assign layer0_outputs[5495] = (inputs[161]) | (inputs[164]);
    assign layer0_outputs[5496] = inputs[138];
    assign layer0_outputs[5497] = ~(inputs[119]);
    assign layer0_outputs[5498] = ~((inputs[67]) | (inputs[65]));
    assign layer0_outputs[5499] = ~((inputs[179]) ^ (inputs[121]));
    assign layer0_outputs[5500] = ~(inputs[132]);
    assign layer0_outputs[5501] = inputs[104];
    assign layer0_outputs[5502] = ~(inputs[120]);
    assign layer0_outputs[5503] = inputs[94];
    assign layer0_outputs[5504] = ~(inputs[183]);
    assign layer0_outputs[5505] = (inputs[143]) | (inputs[61]);
    assign layer0_outputs[5506] = ~(inputs[56]);
    assign layer0_outputs[5507] = ~((inputs[93]) | (inputs[121]));
    assign layer0_outputs[5508] = ~(inputs[105]);
    assign layer0_outputs[5509] = (inputs[42]) | (inputs[92]);
    assign layer0_outputs[5510] = ~(inputs[85]);
    assign layer0_outputs[5511] = (inputs[140]) | (inputs[246]);
    assign layer0_outputs[5512] = ~(inputs[180]);
    assign layer0_outputs[5513] = 1'b0;
    assign layer0_outputs[5514] = ~(inputs[113]);
    assign layer0_outputs[5515] = (inputs[35]) | (inputs[2]);
    assign layer0_outputs[5516] = (inputs[2]) | (inputs[237]);
    assign layer0_outputs[5517] = ~(inputs[45]);
    assign layer0_outputs[5518] = ~(inputs[217]) | (inputs[141]);
    assign layer0_outputs[5519] = (inputs[237]) | (inputs[146]);
    assign layer0_outputs[5520] = ~(inputs[215]) | (inputs[77]);
    assign layer0_outputs[5521] = ~((inputs[115]) | (inputs[156]));
    assign layer0_outputs[5522] = ~(inputs[219]);
    assign layer0_outputs[5523] = inputs[137];
    assign layer0_outputs[5524] = (inputs[229]) | (inputs[118]);
    assign layer0_outputs[5525] = (inputs[242]) & (inputs[228]);
    assign layer0_outputs[5526] = ~((inputs[208]) | (inputs[242]));
    assign layer0_outputs[5527] = (inputs[166]) ^ (inputs[184]);
    assign layer0_outputs[5528] = ~((inputs[34]) ^ (inputs[111]));
    assign layer0_outputs[5529] = ~(inputs[68]) | (inputs[241]);
    assign layer0_outputs[5530] = ~((inputs[92]) | (inputs[77]));
    assign layer0_outputs[5531] = ~(inputs[82]);
    assign layer0_outputs[5532] = ~((inputs[68]) | (inputs[223]));
    assign layer0_outputs[5533] = 1'b0;
    assign layer0_outputs[5534] = (inputs[74]) ^ (inputs[77]);
    assign layer0_outputs[5535] = ~(inputs[19]);
    assign layer0_outputs[5536] = (inputs[209]) | (inputs[216]);
    assign layer0_outputs[5537] = ~((inputs[149]) ^ (inputs[184]));
    assign layer0_outputs[5538] = inputs[169];
    assign layer0_outputs[5539] = ~(inputs[105]);
    assign layer0_outputs[5540] = inputs[25];
    assign layer0_outputs[5541] = ~(inputs[195]);
    assign layer0_outputs[5542] = inputs[236];
    assign layer0_outputs[5543] = (inputs[116]) & ~(inputs[206]);
    assign layer0_outputs[5544] = ~((inputs[236]) ^ (inputs[62]));
    assign layer0_outputs[5545] = (inputs[115]) | (inputs[115]);
    assign layer0_outputs[5546] = inputs[120];
    assign layer0_outputs[5547] = inputs[252];
    assign layer0_outputs[5548] = ~(inputs[245]);
    assign layer0_outputs[5549] = ~(inputs[218]);
    assign layer0_outputs[5550] = ~((inputs[200]) ^ (inputs[174]));
    assign layer0_outputs[5551] = ~(inputs[211]) | (inputs[196]);
    assign layer0_outputs[5552] = inputs[116];
    assign layer0_outputs[5553] = ~(inputs[103]);
    assign layer0_outputs[5554] = inputs[40];
    assign layer0_outputs[5555] = ~(inputs[190]) | (inputs[209]);
    assign layer0_outputs[5556] = (inputs[182]) ^ (inputs[178]);
    assign layer0_outputs[5557] = ~((inputs[28]) | (inputs[14]));
    assign layer0_outputs[5558] = (inputs[190]) & ~(inputs[29]);
    assign layer0_outputs[5559] = ~((inputs[156]) & (inputs[17]));
    assign layer0_outputs[5560] = ~((inputs[7]) | (inputs[20]));
    assign layer0_outputs[5561] = ~(inputs[128]);
    assign layer0_outputs[5562] = ~((inputs[4]) | (inputs[90]));
    assign layer0_outputs[5563] = ~((inputs[171]) & (inputs[134]));
    assign layer0_outputs[5564] = inputs[68];
    assign layer0_outputs[5565] = ~(inputs[156]) | (inputs[237]);
    assign layer0_outputs[5566] = ~(inputs[124]);
    assign layer0_outputs[5567] = ~(inputs[87]) | (inputs[79]);
    assign layer0_outputs[5568] = (inputs[1]) | (inputs[220]);
    assign layer0_outputs[5569] = (inputs[45]) & ~(inputs[96]);
    assign layer0_outputs[5570] = ~(inputs[98]);
    assign layer0_outputs[5571] = (inputs[118]) ^ (inputs[157]);
    assign layer0_outputs[5572] = (inputs[38]) & ~(inputs[167]);
    assign layer0_outputs[5573] = inputs[163];
    assign layer0_outputs[5574] = ~(inputs[228]) | (inputs[118]);
    assign layer0_outputs[5575] = (inputs[242]) & ~(inputs[202]);
    assign layer0_outputs[5576] = ~((inputs[101]) ^ (inputs[99]));
    assign layer0_outputs[5577] = inputs[213];
    assign layer0_outputs[5578] = ~((inputs[221]) | (inputs[181]));
    assign layer0_outputs[5579] = ~(inputs[127]) | (inputs[221]);
    assign layer0_outputs[5580] = (inputs[29]) ^ (inputs[237]);
    assign layer0_outputs[5581] = ~(inputs[180]);
    assign layer0_outputs[5582] = inputs[26];
    assign layer0_outputs[5583] = (inputs[166]) | (inputs[108]);
    assign layer0_outputs[5584] = (inputs[73]) ^ (inputs[132]);
    assign layer0_outputs[5585] = (inputs[171]) | (inputs[33]);
    assign layer0_outputs[5586] = ~(inputs[23]);
    assign layer0_outputs[5587] = ~(inputs[184]) | (inputs[1]);
    assign layer0_outputs[5588] = ~(inputs[30]);
    assign layer0_outputs[5589] = ~(inputs[136]);
    assign layer0_outputs[5590] = ~(inputs[234]);
    assign layer0_outputs[5591] = (inputs[86]) & ~(inputs[111]);
    assign layer0_outputs[5592] = (inputs[122]) ^ (inputs[170]);
    assign layer0_outputs[5593] = ~((inputs[154]) & (inputs[122]));
    assign layer0_outputs[5594] = (inputs[85]) & ~(inputs[224]);
    assign layer0_outputs[5595] = (inputs[62]) & ~(inputs[238]);
    assign layer0_outputs[5596] = (inputs[117]) | (inputs[239]);
    assign layer0_outputs[5597] = ~(inputs[126]);
    assign layer0_outputs[5598] = (inputs[0]) & ~(inputs[12]);
    assign layer0_outputs[5599] = ~((inputs[33]) | (inputs[48]));
    assign layer0_outputs[5600] = ~(inputs[102]) | (inputs[242]);
    assign layer0_outputs[5601] = (inputs[15]) & ~(inputs[61]);
    assign layer0_outputs[5602] = ~(inputs[148]) | (inputs[253]);
    assign layer0_outputs[5603] = (inputs[14]) | (inputs[252]);
    assign layer0_outputs[5604] = ~(inputs[99]) | (inputs[13]);
    assign layer0_outputs[5605] = ~(inputs[142]);
    assign layer0_outputs[5606] = (inputs[174]) | (inputs[188]);
    assign layer0_outputs[5607] = ~(inputs[204]);
    assign layer0_outputs[5608] = inputs[247];
    assign layer0_outputs[5609] = (inputs[229]) & (inputs[165]);
    assign layer0_outputs[5610] = ~((inputs[162]) | (inputs[145]));
    assign layer0_outputs[5611] = ~((inputs[77]) | (inputs[199]));
    assign layer0_outputs[5612] = (inputs[96]) ^ (inputs[104]);
    assign layer0_outputs[5613] = ~(inputs[229]);
    assign layer0_outputs[5614] = ~((inputs[116]) | (inputs[53]));
    assign layer0_outputs[5615] = ~((inputs[50]) | (inputs[83]));
    assign layer0_outputs[5616] = ~(inputs[44]) | (inputs[47]);
    assign layer0_outputs[5617] = ~(inputs[209]) | (inputs[191]);
    assign layer0_outputs[5618] = ~((inputs[97]) | (inputs[53]));
    assign layer0_outputs[5619] = ~((inputs[163]) ^ (inputs[190]));
    assign layer0_outputs[5620] = (inputs[93]) & (inputs[27]);
    assign layer0_outputs[5621] = (inputs[132]) & ~(inputs[224]);
    assign layer0_outputs[5622] = (inputs[5]) & (inputs[181]);
    assign layer0_outputs[5623] = inputs[93];
    assign layer0_outputs[5624] = ~(inputs[82]);
    assign layer0_outputs[5625] = ~(inputs[97]);
    assign layer0_outputs[5626] = (inputs[20]) & ~(inputs[250]);
    assign layer0_outputs[5627] = inputs[185];
    assign layer0_outputs[5628] = ~((inputs[239]) | (inputs[166]));
    assign layer0_outputs[5629] = ~((inputs[233]) | (inputs[209]));
    assign layer0_outputs[5630] = ~((inputs[28]) ^ (inputs[27]));
    assign layer0_outputs[5631] = (inputs[226]) ^ (inputs[96]);
    assign layer0_outputs[5632] = (inputs[9]) & ~(inputs[161]);
    assign layer0_outputs[5633] = inputs[188];
    assign layer0_outputs[5634] = (inputs[185]) | (inputs[4]);
    assign layer0_outputs[5635] = ~((inputs[235]) | (inputs[9]));
    assign layer0_outputs[5636] = ~((inputs[127]) | (inputs[50]));
    assign layer0_outputs[5637] = (inputs[73]) & ~(inputs[109]);
    assign layer0_outputs[5638] = ~(inputs[164]) | (inputs[63]);
    assign layer0_outputs[5639] = (inputs[151]) ^ (inputs[237]);
    assign layer0_outputs[5640] = ~(inputs[148]);
    assign layer0_outputs[5641] = ~(inputs[217]) | (inputs[94]);
    assign layer0_outputs[5642] = (inputs[55]) & ~(inputs[180]);
    assign layer0_outputs[5643] = (inputs[129]) ^ (inputs[48]);
    assign layer0_outputs[5644] = ~((inputs[102]) | (inputs[203]));
    assign layer0_outputs[5645] = ~((inputs[200]) | (inputs[200]));
    assign layer0_outputs[5646] = ~((inputs[254]) | (inputs[199]));
    assign layer0_outputs[5647] = (inputs[171]) & ~(inputs[50]);
    assign layer0_outputs[5648] = (inputs[171]) & ~(inputs[96]);
    assign layer0_outputs[5649] = inputs[117];
    assign layer0_outputs[5650] = inputs[67];
    assign layer0_outputs[5651] = (inputs[254]) ^ (inputs[118]);
    assign layer0_outputs[5652] = inputs[23];
    assign layer0_outputs[5653] = ~((inputs[115]) & (inputs[196]));
    assign layer0_outputs[5654] = (inputs[186]) ^ (inputs[138]);
    assign layer0_outputs[5655] = inputs[250];
    assign layer0_outputs[5656] = inputs[195];
    assign layer0_outputs[5657] = ~((inputs[191]) | (inputs[75]));
    assign layer0_outputs[5658] = 1'b1;
    assign layer0_outputs[5659] = ~(inputs[23]) | (inputs[227]);
    assign layer0_outputs[5660] = ~(inputs[102]);
    assign layer0_outputs[5661] = (inputs[80]) | (inputs[12]);
    assign layer0_outputs[5662] = (inputs[71]) | (inputs[48]);
    assign layer0_outputs[5663] = ~(inputs[185]) | (inputs[133]);
    assign layer0_outputs[5664] = 1'b0;
    assign layer0_outputs[5665] = inputs[41];
    assign layer0_outputs[5666] = ~(inputs[42]);
    assign layer0_outputs[5667] = ~(inputs[21]);
    assign layer0_outputs[5668] = (inputs[209]) | (inputs[101]);
    assign layer0_outputs[5669] = ~(inputs[151]);
    assign layer0_outputs[5670] = ~(inputs[179]) | (inputs[94]);
    assign layer0_outputs[5671] = (inputs[134]) | (inputs[222]);
    assign layer0_outputs[5672] = ~((inputs[156]) ^ (inputs[213]));
    assign layer0_outputs[5673] = (inputs[69]) | (inputs[38]);
    assign layer0_outputs[5674] = ~((inputs[175]) | (inputs[64]));
    assign layer0_outputs[5675] = ~((inputs[56]) & (inputs[109]));
    assign layer0_outputs[5676] = (inputs[14]) | (inputs[239]);
    assign layer0_outputs[5677] = (inputs[216]) ^ (inputs[59]);
    assign layer0_outputs[5678] = inputs[177];
    assign layer0_outputs[5679] = inputs[84];
    assign layer0_outputs[5680] = ~((inputs[226]) ^ (inputs[180]));
    assign layer0_outputs[5681] = ~(inputs[90]);
    assign layer0_outputs[5682] = (inputs[207]) ^ (inputs[236]);
    assign layer0_outputs[5683] = ~(inputs[88]) | (inputs[129]);
    assign layer0_outputs[5684] = (inputs[231]) | (inputs[185]);
    assign layer0_outputs[5685] = ~((inputs[119]) ^ (inputs[232]));
    assign layer0_outputs[5686] = ~((inputs[228]) | (inputs[212]));
    assign layer0_outputs[5687] = inputs[79];
    assign layer0_outputs[5688] = (inputs[138]) & ~(inputs[200]);
    assign layer0_outputs[5689] = (inputs[202]) & ~(inputs[120]);
    assign layer0_outputs[5690] = (inputs[198]) & ~(inputs[118]);
    assign layer0_outputs[5691] = inputs[29];
    assign layer0_outputs[5692] = ~(inputs[69]);
    assign layer0_outputs[5693] = inputs[218];
    assign layer0_outputs[5694] = inputs[216];
    assign layer0_outputs[5695] = 1'b0;
    assign layer0_outputs[5696] = 1'b0;
    assign layer0_outputs[5697] = ~(inputs[233]);
    assign layer0_outputs[5698] = (inputs[86]) | (inputs[149]);
    assign layer0_outputs[5699] = inputs[104];
    assign layer0_outputs[5700] = (inputs[9]) & (inputs[76]);
    assign layer0_outputs[5701] = (inputs[10]) | (inputs[61]);
    assign layer0_outputs[5702] = ~((inputs[45]) ^ (inputs[75]));
    assign layer0_outputs[5703] = inputs[157];
    assign layer0_outputs[5704] = (inputs[139]) | (inputs[178]);
    assign layer0_outputs[5705] = (inputs[110]) | (inputs[3]);
    assign layer0_outputs[5706] = (inputs[238]) & ~(inputs[130]);
    assign layer0_outputs[5707] = inputs[113];
    assign layer0_outputs[5708] = ~(inputs[117]) | (inputs[35]);
    assign layer0_outputs[5709] = (inputs[0]) & ~(inputs[241]);
    assign layer0_outputs[5710] = (inputs[55]) & ~(inputs[204]);
    assign layer0_outputs[5711] = inputs[229];
    assign layer0_outputs[5712] = ~(inputs[97]);
    assign layer0_outputs[5713] = (inputs[22]) | (inputs[228]);
    assign layer0_outputs[5714] = ~((inputs[246]) | (inputs[42]));
    assign layer0_outputs[5715] = (inputs[226]) & (inputs[236]);
    assign layer0_outputs[5716] = ~(inputs[181]);
    assign layer0_outputs[5717] = inputs[24];
    assign layer0_outputs[5718] = (inputs[167]) ^ (inputs[120]);
    assign layer0_outputs[5719] = (inputs[186]) ^ (inputs[185]);
    assign layer0_outputs[5720] = (inputs[163]) & ~(inputs[231]);
    assign layer0_outputs[5721] = ~(inputs[12]) | (inputs[253]);
    assign layer0_outputs[5722] = (inputs[32]) ^ (inputs[6]);
    assign layer0_outputs[5723] = inputs[136];
    assign layer0_outputs[5724] = (inputs[36]) | (inputs[63]);
    assign layer0_outputs[5725] = ~((inputs[106]) ^ (inputs[95]));
    assign layer0_outputs[5726] = ~(inputs[187]) | (inputs[125]);
    assign layer0_outputs[5727] = (inputs[242]) ^ (inputs[53]);
    assign layer0_outputs[5728] = (inputs[111]) & ~(inputs[254]);
    assign layer0_outputs[5729] = ~(inputs[137]) | (inputs[47]);
    assign layer0_outputs[5730] = ~(inputs[35]) | (inputs[129]);
    assign layer0_outputs[5731] = (inputs[204]) | (inputs[20]);
    assign layer0_outputs[5732] = (inputs[7]) ^ (inputs[210]);
    assign layer0_outputs[5733] = inputs[60];
    assign layer0_outputs[5734] = ~(inputs[194]);
    assign layer0_outputs[5735] = (inputs[155]) ^ (inputs[110]);
    assign layer0_outputs[5736] = (inputs[26]) & ~(inputs[222]);
    assign layer0_outputs[5737] = inputs[165];
    assign layer0_outputs[5738] = ~((inputs[79]) | (inputs[36]));
    assign layer0_outputs[5739] = inputs[224];
    assign layer0_outputs[5740] = inputs[168];
    assign layer0_outputs[5741] = (inputs[248]) & ~(inputs[95]);
    assign layer0_outputs[5742] = ~(inputs[29]) | (inputs[180]);
    assign layer0_outputs[5743] = ~((inputs[130]) | (inputs[144]));
    assign layer0_outputs[5744] = 1'b0;
    assign layer0_outputs[5745] = ~((inputs[233]) ^ (inputs[161]));
    assign layer0_outputs[5746] = (inputs[107]) | (inputs[175]);
    assign layer0_outputs[5747] = (inputs[218]) | (inputs[248]);
    assign layer0_outputs[5748] = ~(inputs[87]);
    assign layer0_outputs[5749] = ~(inputs[220]);
    assign layer0_outputs[5750] = (inputs[37]) & ~(inputs[181]);
    assign layer0_outputs[5751] = inputs[210];
    assign layer0_outputs[5752] = ~((inputs[150]) | (inputs[18]));
    assign layer0_outputs[5753] = ~(inputs[82]);
    assign layer0_outputs[5754] = ~(inputs[106]);
    assign layer0_outputs[5755] = inputs[101];
    assign layer0_outputs[5756] = ~(inputs[200]);
    assign layer0_outputs[5757] = (inputs[80]) ^ (inputs[163]);
    assign layer0_outputs[5758] = inputs[164];
    assign layer0_outputs[5759] = ~((inputs[95]) | (inputs[39]));
    assign layer0_outputs[5760] = ~(inputs[120]);
    assign layer0_outputs[5761] = ~((inputs[137]) ^ (inputs[107]));
    assign layer0_outputs[5762] = ~((inputs[196]) | (inputs[141]));
    assign layer0_outputs[5763] = ~((inputs[255]) ^ (inputs[31]));
    assign layer0_outputs[5764] = inputs[115];
    assign layer0_outputs[5765] = 1'b1;
    assign layer0_outputs[5766] = ~(inputs[125]);
    assign layer0_outputs[5767] = inputs[94];
    assign layer0_outputs[5768] = ~((inputs[254]) | (inputs[227]));
    assign layer0_outputs[5769] = inputs[195];
    assign layer0_outputs[5770] = inputs[243];
    assign layer0_outputs[5771] = ~(inputs[185]);
    assign layer0_outputs[5772] = (inputs[117]) | (inputs[114]);
    assign layer0_outputs[5773] = ~((inputs[102]) ^ (inputs[49]));
    assign layer0_outputs[5774] = ~(inputs[99]);
    assign layer0_outputs[5775] = (inputs[188]) | (inputs[107]);
    assign layer0_outputs[5776] = 1'b1;
    assign layer0_outputs[5777] = ~((inputs[239]) ^ (inputs[21]));
    assign layer0_outputs[5778] = inputs[173];
    assign layer0_outputs[5779] = (inputs[65]) | (inputs[134]);
    assign layer0_outputs[5780] = ~(inputs[4]) | (inputs[145]);
    assign layer0_outputs[5781] = (inputs[142]) & ~(inputs[239]);
    assign layer0_outputs[5782] = ~((inputs[146]) ^ (inputs[231]));
    assign layer0_outputs[5783] = ~(inputs[230]);
    assign layer0_outputs[5784] = (inputs[97]) ^ (inputs[255]);
    assign layer0_outputs[5785] = (inputs[216]) & (inputs[30]);
    assign layer0_outputs[5786] = ~(inputs[124]) | (inputs[111]);
    assign layer0_outputs[5787] = ~(inputs[151]);
    assign layer0_outputs[5788] = ~((inputs[0]) ^ (inputs[141]));
    assign layer0_outputs[5789] = (inputs[10]) & ~(inputs[226]);
    assign layer0_outputs[5790] = inputs[166];
    assign layer0_outputs[5791] = ~(inputs[196]) | (inputs[113]);
    assign layer0_outputs[5792] = ~((inputs[62]) ^ (inputs[205]));
    assign layer0_outputs[5793] = (inputs[43]) & ~(inputs[241]);
    assign layer0_outputs[5794] = inputs[6];
    assign layer0_outputs[5795] = ~(inputs[108]);
    assign layer0_outputs[5796] = ~((inputs[108]) | (inputs[58]));
    assign layer0_outputs[5797] = inputs[135];
    assign layer0_outputs[5798] = (inputs[77]) | (inputs[146]);
    assign layer0_outputs[5799] = inputs[26];
    assign layer0_outputs[5800] = inputs[191];
    assign layer0_outputs[5801] = ~(inputs[107]);
    assign layer0_outputs[5802] = ~(inputs[203]) | (inputs[122]);
    assign layer0_outputs[5803] = ~((inputs[69]) ^ (inputs[200]));
    assign layer0_outputs[5804] = (inputs[3]) ^ (inputs[70]);
    assign layer0_outputs[5805] = ~((inputs[216]) | (inputs[17]));
    assign layer0_outputs[5806] = ~(inputs[46]) | (inputs[33]);
    assign layer0_outputs[5807] = (inputs[161]) | (inputs[232]);
    assign layer0_outputs[5808] = ~((inputs[207]) | (inputs[26]));
    assign layer0_outputs[5809] = (inputs[245]) & ~(inputs[166]);
    assign layer0_outputs[5810] = (inputs[72]) | (inputs[232]);
    assign layer0_outputs[5811] = ~((inputs[169]) & (inputs[228]));
    assign layer0_outputs[5812] = (inputs[73]) & ~(inputs[183]);
    assign layer0_outputs[5813] = (inputs[7]) | (inputs[205]);
    assign layer0_outputs[5814] = inputs[102];
    assign layer0_outputs[5815] = inputs[243];
    assign layer0_outputs[5816] = ~(inputs[202]) | (inputs[93]);
    assign layer0_outputs[5817] = ~(inputs[126]);
    assign layer0_outputs[5818] = (inputs[34]) ^ (inputs[80]);
    assign layer0_outputs[5819] = ~(inputs[225]);
    assign layer0_outputs[5820] = ~(inputs[158]) | (inputs[15]);
    assign layer0_outputs[5821] = ~(inputs[154]) | (inputs[254]);
    assign layer0_outputs[5822] = (inputs[23]) ^ (inputs[126]);
    assign layer0_outputs[5823] = inputs[62];
    assign layer0_outputs[5824] = ~((inputs[199]) | (inputs[244]));
    assign layer0_outputs[5825] = ~(inputs[228]);
    assign layer0_outputs[5826] = inputs[114];
    assign layer0_outputs[5827] = ~((inputs[95]) | (inputs[240]));
    assign layer0_outputs[5828] = (inputs[113]) | (inputs[72]);
    assign layer0_outputs[5829] = ~((inputs[250]) ^ (inputs[169]));
    assign layer0_outputs[5830] = ~(inputs[26]) | (inputs[164]);
    assign layer0_outputs[5831] = ~(inputs[167]) | (inputs[39]);
    assign layer0_outputs[5832] = (inputs[14]) & ~(inputs[209]);
    assign layer0_outputs[5833] = inputs[222];
    assign layer0_outputs[5834] = ~(inputs[71]);
    assign layer0_outputs[5835] = inputs[116];
    assign layer0_outputs[5836] = (inputs[46]) & ~(inputs[89]);
    assign layer0_outputs[5837] = inputs[153];
    assign layer0_outputs[5838] = inputs[17];
    assign layer0_outputs[5839] = ~((inputs[191]) ^ (inputs[148]));
    assign layer0_outputs[5840] = inputs[148];
    assign layer0_outputs[5841] = (inputs[142]) | (inputs[222]);
    assign layer0_outputs[5842] = ~(inputs[167]) | (inputs[193]);
    assign layer0_outputs[5843] = ~(inputs[247]) | (inputs[182]);
    assign layer0_outputs[5844] = (inputs[248]) | (inputs[28]);
    assign layer0_outputs[5845] = inputs[140];
    assign layer0_outputs[5846] = (inputs[30]) ^ (inputs[53]);
    assign layer0_outputs[5847] = inputs[55];
    assign layer0_outputs[5848] = (inputs[188]) & ~(inputs[55]);
    assign layer0_outputs[5849] = ~((inputs[143]) & (inputs[96]));
    assign layer0_outputs[5850] = ~((inputs[24]) ^ (inputs[65]));
    assign layer0_outputs[5851] = (inputs[228]) | (inputs[3]);
    assign layer0_outputs[5852] = (inputs[128]) | (inputs[67]);
    assign layer0_outputs[5853] = ~(inputs[130]) | (inputs[11]);
    assign layer0_outputs[5854] = ~((inputs[57]) | (inputs[42]));
    assign layer0_outputs[5855] = ~((inputs[99]) | (inputs[113]));
    assign layer0_outputs[5856] = ~(inputs[149]);
    assign layer0_outputs[5857] = ~(inputs[20]);
    assign layer0_outputs[5858] = (inputs[206]) ^ (inputs[92]);
    assign layer0_outputs[5859] = (inputs[9]) & ~(inputs[210]);
    assign layer0_outputs[5860] = (inputs[173]) & (inputs[216]);
    assign layer0_outputs[5861] = ~(inputs[91]) | (inputs[80]);
    assign layer0_outputs[5862] = (inputs[168]) & ~(inputs[146]);
    assign layer0_outputs[5863] = ~(inputs[145]);
    assign layer0_outputs[5864] = ~(inputs[46]) | (inputs[109]);
    assign layer0_outputs[5865] = (inputs[84]) & ~(inputs[192]);
    assign layer0_outputs[5866] = (inputs[7]) | (inputs[40]);
    assign layer0_outputs[5867] = ~((inputs[106]) & (inputs[90]));
    assign layer0_outputs[5868] = ~(inputs[68]) | (inputs[41]);
    assign layer0_outputs[5869] = ~(inputs[232]);
    assign layer0_outputs[5870] = (inputs[22]) ^ (inputs[69]);
    assign layer0_outputs[5871] = inputs[148];
    assign layer0_outputs[5872] = ~(inputs[114]);
    assign layer0_outputs[5873] = inputs[45];
    assign layer0_outputs[5874] = ~(inputs[24]) | (inputs[163]);
    assign layer0_outputs[5875] = inputs[142];
    assign layer0_outputs[5876] = ~(inputs[251]);
    assign layer0_outputs[5877] = (inputs[90]) & ~(inputs[245]);
    assign layer0_outputs[5878] = (inputs[245]) & ~(inputs[224]);
    assign layer0_outputs[5879] = ~((inputs[254]) ^ (inputs[125]));
    assign layer0_outputs[5880] = inputs[196];
    assign layer0_outputs[5881] = ~(inputs[168]) | (inputs[47]);
    assign layer0_outputs[5882] = ~(inputs[104]);
    assign layer0_outputs[5883] = ~((inputs[151]) ^ (inputs[253]));
    assign layer0_outputs[5884] = (inputs[186]) | (inputs[201]);
    assign layer0_outputs[5885] = 1'b1;
    assign layer0_outputs[5886] = (inputs[25]) ^ (inputs[44]);
    assign layer0_outputs[5887] = ~(inputs[98]);
    assign layer0_outputs[5888] = ~(inputs[75]);
    assign layer0_outputs[5889] = (inputs[207]) ^ (inputs[106]);
    assign layer0_outputs[5890] = inputs[142];
    assign layer0_outputs[5891] = ~(inputs[202]) | (inputs[43]);
    assign layer0_outputs[5892] = ~(inputs[232]);
    assign layer0_outputs[5893] = (inputs[19]) | (inputs[2]);
    assign layer0_outputs[5894] = ~((inputs[28]) | (inputs[14]));
    assign layer0_outputs[5895] = 1'b0;
    assign layer0_outputs[5896] = (inputs[165]) & ~(inputs[66]);
    assign layer0_outputs[5897] = ~(inputs[51]) | (inputs[252]);
    assign layer0_outputs[5898] = ~(inputs[24]) | (inputs[192]);
    assign layer0_outputs[5899] = ~(inputs[71]) | (inputs[45]);
    assign layer0_outputs[5900] = ~((inputs[164]) | (inputs[219]));
    assign layer0_outputs[5901] = (inputs[27]) ^ (inputs[57]);
    assign layer0_outputs[5902] = 1'b1;
    assign layer0_outputs[5903] = inputs[101];
    assign layer0_outputs[5904] = inputs[90];
    assign layer0_outputs[5905] = (inputs[90]) & ~(inputs[187]);
    assign layer0_outputs[5906] = (inputs[101]) & ~(inputs[73]);
    assign layer0_outputs[5907] = ~((inputs[218]) | (inputs[230]));
    assign layer0_outputs[5908] = ~(inputs[162]);
    assign layer0_outputs[5909] = ~(inputs[213]);
    assign layer0_outputs[5910] = (inputs[188]) & (inputs[177]);
    assign layer0_outputs[5911] = (inputs[254]) | (inputs[54]);
    assign layer0_outputs[5912] = ~(inputs[230]) | (inputs[89]);
    assign layer0_outputs[5913] = (inputs[100]) & ~(inputs[80]);
    assign layer0_outputs[5914] = (inputs[172]) ^ (inputs[97]);
    assign layer0_outputs[5915] = (inputs[57]) & (inputs[221]);
    assign layer0_outputs[5916] = (inputs[172]) ^ (inputs[234]);
    assign layer0_outputs[5917] = inputs[103];
    assign layer0_outputs[5918] = ~((inputs[16]) | (inputs[9]));
    assign layer0_outputs[5919] = (inputs[197]) & (inputs[156]);
    assign layer0_outputs[5920] = inputs[94];
    assign layer0_outputs[5921] = inputs[195];
    assign layer0_outputs[5922] = ~(inputs[117]);
    assign layer0_outputs[5923] = ~(inputs[5]);
    assign layer0_outputs[5924] = (inputs[230]) & ~(inputs[107]);
    assign layer0_outputs[5925] = inputs[55];
    assign layer0_outputs[5926] = ~(inputs[80]);
    assign layer0_outputs[5927] = ~((inputs[119]) | (inputs[13]));
    assign layer0_outputs[5928] = (inputs[52]) & ~(inputs[120]);
    assign layer0_outputs[5929] = (inputs[253]) ^ (inputs[75]);
    assign layer0_outputs[5930] = (inputs[91]) & (inputs[25]);
    assign layer0_outputs[5931] = ~(inputs[142]) | (inputs[220]);
    assign layer0_outputs[5932] = (inputs[152]) & ~(inputs[27]);
    assign layer0_outputs[5933] = ~((inputs[222]) | (inputs[138]));
    assign layer0_outputs[5934] = ~(inputs[26]) | (inputs[250]);
    assign layer0_outputs[5935] = ~(inputs[68]) | (inputs[222]);
    assign layer0_outputs[5936] = ~(inputs[186]);
    assign layer0_outputs[5937] = ~(inputs[112]);
    assign layer0_outputs[5938] = (inputs[174]) & (inputs[60]);
    assign layer0_outputs[5939] = (inputs[158]) | (inputs[244]);
    assign layer0_outputs[5940] = (inputs[117]) & (inputs[168]);
    assign layer0_outputs[5941] = inputs[157];
    assign layer0_outputs[5942] = ~(inputs[121]);
    assign layer0_outputs[5943] = inputs[223];
    assign layer0_outputs[5944] = inputs[153];
    assign layer0_outputs[5945] = ~((inputs[54]) ^ (inputs[52]));
    assign layer0_outputs[5946] = ~((inputs[189]) | (inputs[32]));
    assign layer0_outputs[5947] = ~(inputs[110]) | (inputs[123]);
    assign layer0_outputs[5948] = ~(inputs[60]) | (inputs[204]);
    assign layer0_outputs[5949] = inputs[124];
    assign layer0_outputs[5950] = ~((inputs[57]) | (inputs[220]));
    assign layer0_outputs[5951] = ~(inputs[198]) | (inputs[121]);
    assign layer0_outputs[5952] = (inputs[157]) | (inputs[153]);
    assign layer0_outputs[5953] = (inputs[172]) & ~(inputs[65]);
    assign layer0_outputs[5954] = ~(inputs[240]) | (inputs[27]);
    assign layer0_outputs[5955] = ~((inputs[236]) | (inputs[178]));
    assign layer0_outputs[5956] = ~(inputs[23]);
    assign layer0_outputs[5957] = ~((inputs[221]) | (inputs[174]));
    assign layer0_outputs[5958] = ~(inputs[223]) | (inputs[107]);
    assign layer0_outputs[5959] = ~(inputs[78]);
    assign layer0_outputs[5960] = ~(inputs[55]);
    assign layer0_outputs[5961] = ~((inputs[171]) ^ (inputs[125]));
    assign layer0_outputs[5962] = (inputs[122]) & ~(inputs[36]);
    assign layer0_outputs[5963] = ~((inputs[99]) | (inputs[237]));
    assign layer0_outputs[5964] = ~(inputs[8]);
    assign layer0_outputs[5965] = ~(inputs[248]) | (inputs[26]);
    assign layer0_outputs[5966] = ~(inputs[239]);
    assign layer0_outputs[5967] = ~(inputs[250]);
    assign layer0_outputs[5968] = (inputs[237]) & (inputs[158]);
    assign layer0_outputs[5969] = (inputs[130]) & ~(inputs[224]);
    assign layer0_outputs[5970] = (inputs[25]) & (inputs[133]);
    assign layer0_outputs[5971] = ~((inputs[37]) | (inputs[189]));
    assign layer0_outputs[5972] = (inputs[7]) & ~(inputs[15]);
    assign layer0_outputs[5973] = inputs[166];
    assign layer0_outputs[5974] = ~((inputs[59]) | (inputs[111]));
    assign layer0_outputs[5975] = inputs[151];
    assign layer0_outputs[5976] = ~((inputs[64]) | (inputs[133]));
    assign layer0_outputs[5977] = (inputs[21]) & ~(inputs[251]);
    assign layer0_outputs[5978] = (inputs[94]) | (inputs[136]);
    assign layer0_outputs[5979] = inputs[244];
    assign layer0_outputs[5980] = inputs[56];
    assign layer0_outputs[5981] = (inputs[23]) & ~(inputs[19]);
    assign layer0_outputs[5982] = ~(inputs[27]);
    assign layer0_outputs[5983] = ~((inputs[60]) | (inputs[35]));
    assign layer0_outputs[5984] = inputs[42];
    assign layer0_outputs[5985] = ~(inputs[80]);
    assign layer0_outputs[5986] = (inputs[154]) & ~(inputs[33]);
    assign layer0_outputs[5987] = ~((inputs[4]) | (inputs[235]));
    assign layer0_outputs[5988] = ~(inputs[73]);
    assign layer0_outputs[5989] = (inputs[216]) | (inputs[36]);
    assign layer0_outputs[5990] = ~(inputs[227]);
    assign layer0_outputs[5991] = (inputs[169]) & ~(inputs[79]);
    assign layer0_outputs[5992] = inputs[124];
    assign layer0_outputs[5993] = ~(inputs[129]);
    assign layer0_outputs[5994] = (inputs[171]) & ~(inputs[14]);
    assign layer0_outputs[5995] = (inputs[184]) ^ (inputs[26]);
    assign layer0_outputs[5996] = (inputs[138]) & ~(inputs[198]);
    assign layer0_outputs[5997] = ~((inputs[219]) | (inputs[210]));
    assign layer0_outputs[5998] = inputs[92];
    assign layer0_outputs[5999] = (inputs[19]) | (inputs[147]);
    assign layer0_outputs[6000] = ~((inputs[123]) & (inputs[203]));
    assign layer0_outputs[6001] = ~(inputs[124]) | (inputs[78]);
    assign layer0_outputs[6002] = ~((inputs[200]) ^ (inputs[100]));
    assign layer0_outputs[6003] = (inputs[114]) | (inputs[117]);
    assign layer0_outputs[6004] = inputs[145];
    assign layer0_outputs[6005] = ~(inputs[131]);
    assign layer0_outputs[6006] = ~(inputs[245]);
    assign layer0_outputs[6007] = (inputs[75]) & ~(inputs[238]);
    assign layer0_outputs[6008] = (inputs[189]) | (inputs[126]);
    assign layer0_outputs[6009] = (inputs[53]) | (inputs[26]);
    assign layer0_outputs[6010] = ~(inputs[25]);
    assign layer0_outputs[6011] = ~(inputs[116]) | (inputs[173]);
    assign layer0_outputs[6012] = (inputs[131]) & ~(inputs[16]);
    assign layer0_outputs[6013] = ~(inputs[57]);
    assign layer0_outputs[6014] = (inputs[37]) | (inputs[78]);
    assign layer0_outputs[6015] = ~(inputs[99]);
    assign layer0_outputs[6016] = inputs[238];
    assign layer0_outputs[6017] = ~((inputs[165]) | (inputs[24]));
    assign layer0_outputs[6018] = ~(inputs[14]);
    assign layer0_outputs[6019] = ~(inputs[50]) | (inputs[144]);
    assign layer0_outputs[6020] = ~(inputs[172]);
    assign layer0_outputs[6021] = ~(inputs[76]) | (inputs[38]);
    assign layer0_outputs[6022] = (inputs[247]) | (inputs[201]);
    assign layer0_outputs[6023] = (inputs[27]) ^ (inputs[215]);
    assign layer0_outputs[6024] = inputs[95];
    assign layer0_outputs[6025] = ~(inputs[69]);
    assign layer0_outputs[6026] = 1'b0;
    assign layer0_outputs[6027] = (inputs[76]) & (inputs[215]);
    assign layer0_outputs[6028] = (inputs[120]) & ~(inputs[173]);
    assign layer0_outputs[6029] = ~(inputs[88]) | (inputs[192]);
    assign layer0_outputs[6030] = ~(inputs[138]) | (inputs[217]);
    assign layer0_outputs[6031] = ~((inputs[41]) | (inputs[190]));
    assign layer0_outputs[6032] = (inputs[239]) | (inputs[122]);
    assign layer0_outputs[6033] = (inputs[156]) ^ (inputs[32]);
    assign layer0_outputs[6034] = (inputs[125]) & ~(inputs[225]);
    assign layer0_outputs[6035] = ~((inputs[217]) | (inputs[209]));
    assign layer0_outputs[6036] = (inputs[242]) | (inputs[152]);
    assign layer0_outputs[6037] = ~(inputs[79]);
    assign layer0_outputs[6038] = ~((inputs[149]) ^ (inputs[119]));
    assign layer0_outputs[6039] = inputs[82];
    assign layer0_outputs[6040] = (inputs[39]) | (inputs[223]);
    assign layer0_outputs[6041] = ~(inputs[190]);
    assign layer0_outputs[6042] = (inputs[115]) ^ (inputs[96]);
    assign layer0_outputs[6043] = ~(inputs[6]) | (inputs[81]);
    assign layer0_outputs[6044] = (inputs[20]) | (inputs[125]);
    assign layer0_outputs[6045] = (inputs[56]) & ~(inputs[227]);
    assign layer0_outputs[6046] = (inputs[129]) & ~(inputs[190]);
    assign layer0_outputs[6047] = (inputs[67]) | (inputs[116]);
    assign layer0_outputs[6048] = ~((inputs[104]) & (inputs[27]));
    assign layer0_outputs[6049] = 1'b0;
    assign layer0_outputs[6050] = inputs[34];
    assign layer0_outputs[6051] = inputs[87];
    assign layer0_outputs[6052] = inputs[223];
    assign layer0_outputs[6053] = (inputs[123]) & ~(inputs[150]);
    assign layer0_outputs[6054] = ~(inputs[90]);
    assign layer0_outputs[6055] = inputs[60];
    assign layer0_outputs[6056] = (inputs[91]) & ~(inputs[160]);
    assign layer0_outputs[6057] = ~((inputs[186]) ^ (inputs[145]));
    assign layer0_outputs[6058] = ~((inputs[47]) | (inputs[13]));
    assign layer0_outputs[6059] = 1'b1;
    assign layer0_outputs[6060] = ~((inputs[237]) | (inputs[127]));
    assign layer0_outputs[6061] = ~((inputs[51]) | (inputs[184]));
    assign layer0_outputs[6062] = (inputs[22]) & ~(inputs[147]);
    assign layer0_outputs[6063] = ~((inputs[185]) ^ (inputs[218]));
    assign layer0_outputs[6064] = ~((inputs[61]) | (inputs[211]));
    assign layer0_outputs[6065] = ~((inputs[78]) ^ (inputs[175]));
    assign layer0_outputs[6066] = ~(inputs[222]);
    assign layer0_outputs[6067] = ~(inputs[245]);
    assign layer0_outputs[6068] = ~(inputs[219]);
    assign layer0_outputs[6069] = (inputs[125]) ^ (inputs[104]);
    assign layer0_outputs[6070] = inputs[153];
    assign layer0_outputs[6071] = (inputs[78]) | (inputs[93]);
    assign layer0_outputs[6072] = (inputs[139]) & (inputs[125]);
    assign layer0_outputs[6073] = ~((inputs[233]) | (inputs[87]));
    assign layer0_outputs[6074] = (inputs[40]) & ~(inputs[22]);
    assign layer0_outputs[6075] = ~(inputs[7]);
    assign layer0_outputs[6076] = (inputs[191]) | (inputs[145]);
    assign layer0_outputs[6077] = inputs[84];
    assign layer0_outputs[6078] = (inputs[234]) & ~(inputs[112]);
    assign layer0_outputs[6079] = ~(inputs[108]);
    assign layer0_outputs[6080] = (inputs[90]) | (inputs[107]);
    assign layer0_outputs[6081] = (inputs[10]) ^ (inputs[19]);
    assign layer0_outputs[6082] = (inputs[29]) | (inputs[188]);
    assign layer0_outputs[6083] = ~(inputs[120]);
    assign layer0_outputs[6084] = ~(inputs[176]);
    assign layer0_outputs[6085] = ~((inputs[81]) & (inputs[112]));
    assign layer0_outputs[6086] = (inputs[230]) ^ (inputs[4]);
    assign layer0_outputs[6087] = (inputs[240]) ^ (inputs[240]);
    assign layer0_outputs[6088] = ~(inputs[148]);
    assign layer0_outputs[6089] = ~((inputs[139]) & (inputs[200]));
    assign layer0_outputs[6090] = ~(inputs[6]) | (inputs[62]);
    assign layer0_outputs[6091] = ~((inputs[222]) | (inputs[153]));
    assign layer0_outputs[6092] = ~((inputs[101]) | (inputs[222]));
    assign layer0_outputs[6093] = ~(inputs[183]);
    assign layer0_outputs[6094] = ~(inputs[208]) | (inputs[156]);
    assign layer0_outputs[6095] = 1'b0;
    assign layer0_outputs[6096] = ~((inputs[209]) | (inputs[226]));
    assign layer0_outputs[6097] = ~((inputs[49]) & (inputs[188]));
    assign layer0_outputs[6098] = ~(inputs[71]) | (inputs[140]);
    assign layer0_outputs[6099] = inputs[82];
    assign layer0_outputs[6100] = ~((inputs[48]) ^ (inputs[1]));
    assign layer0_outputs[6101] = ~(inputs[86]);
    assign layer0_outputs[6102] = ~(inputs[139]) | (inputs[6]);
    assign layer0_outputs[6103] = ~(inputs[150]) | (inputs[57]);
    assign layer0_outputs[6104] = ~(inputs[93]) | (inputs[130]);
    assign layer0_outputs[6105] = ~(inputs[226]);
    assign layer0_outputs[6106] = ~((inputs[91]) | (inputs[190]));
    assign layer0_outputs[6107] = (inputs[131]) ^ (inputs[80]);
    assign layer0_outputs[6108] = ~((inputs[22]) ^ (inputs[174]));
    assign layer0_outputs[6109] = ~(inputs[91]);
    assign layer0_outputs[6110] = (inputs[142]) & ~(inputs[239]);
    assign layer0_outputs[6111] = (inputs[254]) ^ (inputs[10]);
    assign layer0_outputs[6112] = ~(inputs[201]);
    assign layer0_outputs[6113] = (inputs[121]) | (inputs[97]);
    assign layer0_outputs[6114] = ~((inputs[27]) ^ (inputs[22]));
    assign layer0_outputs[6115] = inputs[19];
    assign layer0_outputs[6116] = (inputs[137]) | (inputs[122]);
    assign layer0_outputs[6117] = ~(inputs[229]);
    assign layer0_outputs[6118] = inputs[120];
    assign layer0_outputs[6119] = ~((inputs[103]) | (inputs[181]));
    assign layer0_outputs[6120] = ~(inputs[103]);
    assign layer0_outputs[6121] = ~(inputs[199]);
    assign layer0_outputs[6122] = 1'b1;
    assign layer0_outputs[6123] = (inputs[240]) | (inputs[1]);
    assign layer0_outputs[6124] = (inputs[163]) & ~(inputs[174]);
    assign layer0_outputs[6125] = ~((inputs[156]) ^ (inputs[103]));
    assign layer0_outputs[6126] = inputs[189];
    assign layer0_outputs[6127] = inputs[90];
    assign layer0_outputs[6128] = (inputs[32]) ^ (inputs[255]);
    assign layer0_outputs[6129] = ~((inputs[80]) | (inputs[46]));
    assign layer0_outputs[6130] = inputs[26];
    assign layer0_outputs[6131] = inputs[68];
    assign layer0_outputs[6132] = inputs[135];
    assign layer0_outputs[6133] = 1'b1;
    assign layer0_outputs[6134] = (inputs[52]) | (inputs[98]);
    assign layer0_outputs[6135] = (inputs[32]) | (inputs[149]);
    assign layer0_outputs[6136] = ~(inputs[87]);
    assign layer0_outputs[6137] = (inputs[213]) & ~(inputs[17]);
    assign layer0_outputs[6138] = ~(inputs[105]);
    assign layer0_outputs[6139] = inputs[103];
    assign layer0_outputs[6140] = ~((inputs[141]) | (inputs[169]));
    assign layer0_outputs[6141] = ~(inputs[21]) | (inputs[5]);
    assign layer0_outputs[6142] = ~((inputs[174]) ^ (inputs[85]));
    assign layer0_outputs[6143] = inputs[101];
    assign layer0_outputs[6144] = ~((inputs[43]) ^ (inputs[55]));
    assign layer0_outputs[6145] = (inputs[4]) | (inputs[13]);
    assign layer0_outputs[6146] = (inputs[69]) | (inputs[68]);
    assign layer0_outputs[6147] = (inputs[195]) | (inputs[220]);
    assign layer0_outputs[6148] = ~(inputs[135]) | (inputs[208]);
    assign layer0_outputs[6149] = ~((inputs[203]) ^ (inputs[195]));
    assign layer0_outputs[6150] = (inputs[13]) | (inputs[224]);
    assign layer0_outputs[6151] = ~((inputs[235]) | (inputs[254]));
    assign layer0_outputs[6152] = (inputs[69]) & ~(inputs[51]);
    assign layer0_outputs[6153] = ~(inputs[195]);
    assign layer0_outputs[6154] = ~((inputs[230]) ^ (inputs[160]));
    assign layer0_outputs[6155] = (inputs[200]) & (inputs[172]);
    assign layer0_outputs[6156] = ~(inputs[246]);
    assign layer0_outputs[6157] = inputs[229];
    assign layer0_outputs[6158] = (inputs[134]) | (inputs[239]);
    assign layer0_outputs[6159] = ~(inputs[189]);
    assign layer0_outputs[6160] = ~(inputs[70]);
    assign layer0_outputs[6161] = ~((inputs[185]) ^ (inputs[201]));
    assign layer0_outputs[6162] = ~(inputs[183]);
    assign layer0_outputs[6163] = inputs[41];
    assign layer0_outputs[6164] = (inputs[148]) & ~(inputs[221]);
    assign layer0_outputs[6165] = (inputs[43]) & ~(inputs[222]);
    assign layer0_outputs[6166] = ~((inputs[222]) & (inputs[236]));
    assign layer0_outputs[6167] = ~(inputs[134]);
    assign layer0_outputs[6168] = (inputs[172]) & ~(inputs[110]);
    assign layer0_outputs[6169] = ~(inputs[215]) | (inputs[93]);
    assign layer0_outputs[6170] = (inputs[82]) ^ (inputs[133]);
    assign layer0_outputs[6171] = ~(inputs[197]) | (inputs[215]);
    assign layer0_outputs[6172] = (inputs[165]) & ~(inputs[242]);
    assign layer0_outputs[6173] = (inputs[228]) & ~(inputs[15]);
    assign layer0_outputs[6174] = (inputs[5]) ^ (inputs[53]);
    assign layer0_outputs[6175] = ~((inputs[176]) | (inputs[169]));
    assign layer0_outputs[6176] = ~(inputs[188]) | (inputs[250]);
    assign layer0_outputs[6177] = inputs[249];
    assign layer0_outputs[6178] = (inputs[132]) | (inputs[248]);
    assign layer0_outputs[6179] = inputs[69];
    assign layer0_outputs[6180] = (inputs[244]) | (inputs[242]);
    assign layer0_outputs[6181] = (inputs[95]) | (inputs[213]);
    assign layer0_outputs[6182] = (inputs[16]) | (inputs[154]);
    assign layer0_outputs[6183] = ~(inputs[161]) | (inputs[15]);
    assign layer0_outputs[6184] = (inputs[100]) | (inputs[10]);
    assign layer0_outputs[6185] = (inputs[246]) ^ (inputs[182]);
    assign layer0_outputs[6186] = ~(inputs[203]) | (inputs[236]);
    assign layer0_outputs[6187] = inputs[176];
    assign layer0_outputs[6188] = ~((inputs[127]) | (inputs[170]));
    assign layer0_outputs[6189] = (inputs[208]) | (inputs[166]);
    assign layer0_outputs[6190] = ~((inputs[23]) | (inputs[63]));
    assign layer0_outputs[6191] = ~(inputs[119]) | (inputs[163]);
    assign layer0_outputs[6192] = ~(inputs[239]);
    assign layer0_outputs[6193] = ~(inputs[148]);
    assign layer0_outputs[6194] = (inputs[154]) ^ (inputs[231]);
    assign layer0_outputs[6195] = (inputs[55]) | (inputs[245]);
    assign layer0_outputs[6196] = (inputs[106]) & ~(inputs[15]);
    assign layer0_outputs[6197] = ~((inputs[138]) ^ (inputs[109]));
    assign layer0_outputs[6198] = ~(inputs[68]);
    assign layer0_outputs[6199] = ~(inputs[126]);
    assign layer0_outputs[6200] = ~(inputs[10]);
    assign layer0_outputs[6201] = (inputs[75]) & (inputs[36]);
    assign layer0_outputs[6202] = inputs[178];
    assign layer0_outputs[6203] = ~((inputs[6]) ^ (inputs[225]));
    assign layer0_outputs[6204] = (inputs[10]) ^ (inputs[138]);
    assign layer0_outputs[6205] = (inputs[223]) | (inputs[7]);
    assign layer0_outputs[6206] = (inputs[65]) & (inputs[45]);
    assign layer0_outputs[6207] = ~(inputs[155]);
    assign layer0_outputs[6208] = ~(inputs[225]) | (inputs[237]);
    assign layer0_outputs[6209] = ~(inputs[40]) | (inputs[190]);
    assign layer0_outputs[6210] = (inputs[30]) & ~(inputs[175]);
    assign layer0_outputs[6211] = inputs[39];
    assign layer0_outputs[6212] = ~(inputs[174]) | (inputs[13]);
    assign layer0_outputs[6213] = ~(inputs[35]);
    assign layer0_outputs[6214] = (inputs[158]) | (inputs[32]);
    assign layer0_outputs[6215] = ~((inputs[89]) ^ (inputs[168]));
    assign layer0_outputs[6216] = (inputs[175]) ^ (inputs[46]);
    assign layer0_outputs[6217] = ~((inputs[161]) ^ (inputs[164]));
    assign layer0_outputs[6218] = (inputs[80]) | (inputs[92]);
    assign layer0_outputs[6219] = ~((inputs[37]) | (inputs[94]));
    assign layer0_outputs[6220] = ~(inputs[167]);
    assign layer0_outputs[6221] = ~((inputs[194]) & (inputs[18]));
    assign layer0_outputs[6222] = 1'b1;
    assign layer0_outputs[6223] = (inputs[219]) & ~(inputs[130]);
    assign layer0_outputs[6224] = ~((inputs[157]) & (inputs[143]));
    assign layer0_outputs[6225] = ~((inputs[88]) ^ (inputs[146]));
    assign layer0_outputs[6226] = ~(inputs[230]) | (inputs[77]);
    assign layer0_outputs[6227] = (inputs[71]) & (inputs[103]);
    assign layer0_outputs[6228] = ~(inputs[131]);
    assign layer0_outputs[6229] = (inputs[197]) ^ (inputs[50]);
    assign layer0_outputs[6230] = ~((inputs[122]) ^ (inputs[61]));
    assign layer0_outputs[6231] = ~(inputs[23]) | (inputs[179]);
    assign layer0_outputs[6232] = ~(inputs[3]);
    assign layer0_outputs[6233] = (inputs[255]) | (inputs[248]);
    assign layer0_outputs[6234] = inputs[192];
    assign layer0_outputs[6235] = ~(inputs[247]);
    assign layer0_outputs[6236] = ~(inputs[119]);
    assign layer0_outputs[6237] = ~((inputs[54]) ^ (inputs[38]));
    assign layer0_outputs[6238] = ~(inputs[166]);
    assign layer0_outputs[6239] = ~((inputs[14]) | (inputs[254]));
    assign layer0_outputs[6240] = ~(inputs[24]);
    assign layer0_outputs[6241] = ~((inputs[222]) | (inputs[72]));
    assign layer0_outputs[6242] = ~((inputs[207]) | (inputs[161]));
    assign layer0_outputs[6243] = ~((inputs[28]) | (inputs[123]));
    assign layer0_outputs[6244] = (inputs[249]) ^ (inputs[86]);
    assign layer0_outputs[6245] = (inputs[68]) | (inputs[32]);
    assign layer0_outputs[6246] = ~(inputs[92]);
    assign layer0_outputs[6247] = inputs[254];
    assign layer0_outputs[6248] = ~(inputs[125]) | (inputs[222]);
    assign layer0_outputs[6249] = ~(inputs[111]);
    assign layer0_outputs[6250] = (inputs[229]) & ~(inputs[42]);
    assign layer0_outputs[6251] = ~(inputs[9]) | (inputs[129]);
    assign layer0_outputs[6252] = inputs[39];
    assign layer0_outputs[6253] = ~((inputs[198]) | (inputs[64]));
    assign layer0_outputs[6254] = inputs[113];
    assign layer0_outputs[6255] = (inputs[119]) & ~(inputs[126]);
    assign layer0_outputs[6256] = ~(inputs[3]);
    assign layer0_outputs[6257] = ~(inputs[61]) | (inputs[129]);
    assign layer0_outputs[6258] = ~(inputs[227]);
    assign layer0_outputs[6259] = ~(inputs[0]) | (inputs[4]);
    assign layer0_outputs[6260] = (inputs[61]) | (inputs[239]);
    assign layer0_outputs[6261] = (inputs[193]) | (inputs[246]);
    assign layer0_outputs[6262] = ~(inputs[172]);
    assign layer0_outputs[6263] = (inputs[203]) & ~(inputs[1]);
    assign layer0_outputs[6264] = inputs[104];
    assign layer0_outputs[6265] = ~((inputs[67]) | (inputs[5]));
    assign layer0_outputs[6266] = (inputs[143]) | (inputs[77]);
    assign layer0_outputs[6267] = inputs[121];
    assign layer0_outputs[6268] = 1'b0;
    assign layer0_outputs[6269] = inputs[183];
    assign layer0_outputs[6270] = ~(inputs[9]);
    assign layer0_outputs[6271] = ~((inputs[44]) ^ (inputs[209]));
    assign layer0_outputs[6272] = (inputs[92]) ^ (inputs[19]);
    assign layer0_outputs[6273] = inputs[55];
    assign layer0_outputs[6274] = ~(inputs[155]);
    assign layer0_outputs[6275] = inputs[141];
    assign layer0_outputs[6276] = ~(inputs[250]);
    assign layer0_outputs[6277] = ~((inputs[221]) | (inputs[20]));
    assign layer0_outputs[6278] = ~(inputs[150]) | (inputs[208]);
    assign layer0_outputs[6279] = inputs[100];
    assign layer0_outputs[6280] = ~(inputs[184]) | (inputs[245]);
    assign layer0_outputs[6281] = (inputs[17]) & (inputs[126]);
    assign layer0_outputs[6282] = ~(inputs[226]);
    assign layer0_outputs[6283] = (inputs[9]) | (inputs[160]);
    assign layer0_outputs[6284] = ~(inputs[77]) | (inputs[80]);
    assign layer0_outputs[6285] = ~(inputs[153]) | (inputs[174]);
    assign layer0_outputs[6286] = ~(inputs[184]) | (inputs[131]);
    assign layer0_outputs[6287] = (inputs[184]) ^ (inputs[176]);
    assign layer0_outputs[6288] = ~((inputs[70]) & (inputs[73]));
    assign layer0_outputs[6289] = inputs[230];
    assign layer0_outputs[6290] = ~(inputs[153]);
    assign layer0_outputs[6291] = ~(inputs[40]);
    assign layer0_outputs[6292] = ~(inputs[216]);
    assign layer0_outputs[6293] = inputs[1];
    assign layer0_outputs[6294] = (inputs[188]) | (inputs[216]);
    assign layer0_outputs[6295] = (inputs[129]) & ~(inputs[10]);
    assign layer0_outputs[6296] = ~((inputs[72]) | (inputs[93]));
    assign layer0_outputs[6297] = inputs[2];
    assign layer0_outputs[6298] = ~((inputs[79]) ^ (inputs[37]));
    assign layer0_outputs[6299] = (inputs[212]) & (inputs[200]);
    assign layer0_outputs[6300] = ~((inputs[49]) ^ (inputs[228]));
    assign layer0_outputs[6301] = (inputs[253]) & ~(inputs[95]);
    assign layer0_outputs[6302] = ~((inputs[206]) ^ (inputs[87]));
    assign layer0_outputs[6303] = 1'b0;
    assign layer0_outputs[6304] = ~(inputs[39]);
    assign layer0_outputs[6305] = (inputs[149]) & ~(inputs[33]);
    assign layer0_outputs[6306] = ~(inputs[41]);
    assign layer0_outputs[6307] = inputs[109];
    assign layer0_outputs[6308] = inputs[202];
    assign layer0_outputs[6309] = ~((inputs[21]) | (inputs[87]));
    assign layer0_outputs[6310] = ~((inputs[171]) ^ (inputs[205]));
    assign layer0_outputs[6311] = ~((inputs[148]) & (inputs[26]));
    assign layer0_outputs[6312] = (inputs[136]) ^ (inputs[21]);
    assign layer0_outputs[6313] = (inputs[63]) | (inputs[55]);
    assign layer0_outputs[6314] = ~((inputs[101]) | (inputs[180]));
    assign layer0_outputs[6315] = ~(inputs[18]) | (inputs[63]);
    assign layer0_outputs[6316] = (inputs[160]) | (inputs[66]);
    assign layer0_outputs[6317] = ~((inputs[173]) ^ (inputs[69]));
    assign layer0_outputs[6318] = inputs[25];
    assign layer0_outputs[6319] = ~((inputs[92]) | (inputs[93]));
    assign layer0_outputs[6320] = (inputs[169]) | (inputs[64]);
    assign layer0_outputs[6321] = ~((inputs[163]) | (inputs[148]));
    assign layer0_outputs[6322] = ~((inputs[4]) ^ (inputs[148]));
    assign layer0_outputs[6323] = ~(inputs[92]) | (inputs[241]);
    assign layer0_outputs[6324] = inputs[89];
    assign layer0_outputs[6325] = (inputs[51]) ^ (inputs[52]);
    assign layer0_outputs[6326] = ~((inputs[171]) & (inputs[198]));
    assign layer0_outputs[6327] = 1'b1;
    assign layer0_outputs[6328] = inputs[157];
    assign layer0_outputs[6329] = (inputs[207]) & ~(inputs[128]);
    assign layer0_outputs[6330] = ~(inputs[100]);
    assign layer0_outputs[6331] = (inputs[52]) & ~(inputs[175]);
    assign layer0_outputs[6332] = ~(inputs[177]) | (inputs[14]);
    assign layer0_outputs[6333] = ~((inputs[103]) ^ (inputs[97]));
    assign layer0_outputs[6334] = ~((inputs[17]) | (inputs[90]));
    assign layer0_outputs[6335] = ~(inputs[24]) | (inputs[241]);
    assign layer0_outputs[6336] = ~(inputs[152]);
    assign layer0_outputs[6337] = (inputs[85]) & ~(inputs[27]);
    assign layer0_outputs[6338] = (inputs[58]) | (inputs[183]);
    assign layer0_outputs[6339] = ~((inputs[10]) | (inputs[127]));
    assign layer0_outputs[6340] = ~((inputs[35]) | (inputs[13]));
    assign layer0_outputs[6341] = ~(inputs[85]) | (inputs[160]);
    assign layer0_outputs[6342] = (inputs[32]) & ~(inputs[25]);
    assign layer0_outputs[6343] = (inputs[28]) ^ (inputs[138]);
    assign layer0_outputs[6344] = (inputs[137]) & ~(inputs[96]);
    assign layer0_outputs[6345] = (inputs[81]) | (inputs[89]);
    assign layer0_outputs[6346] = inputs[123];
    assign layer0_outputs[6347] = ~(inputs[190]);
    assign layer0_outputs[6348] = ~((inputs[88]) ^ (inputs[56]));
    assign layer0_outputs[6349] = ~(inputs[182]);
    assign layer0_outputs[6350] = (inputs[184]) & (inputs[232]);
    assign layer0_outputs[6351] = ~(inputs[170]);
    assign layer0_outputs[6352] = ~(inputs[42]);
    assign layer0_outputs[6353] = ~((inputs[80]) | (inputs[104]));
    assign layer0_outputs[6354] = ~(inputs[235]) | (inputs[15]);
    assign layer0_outputs[6355] = inputs[76];
    assign layer0_outputs[6356] = (inputs[226]) ^ (inputs[65]);
    assign layer0_outputs[6357] = (inputs[38]) ^ (inputs[207]);
    assign layer0_outputs[6358] = ~(inputs[108]) | (inputs[66]);
    assign layer0_outputs[6359] = ~((inputs[127]) | (inputs[131]));
    assign layer0_outputs[6360] = inputs[248];
    assign layer0_outputs[6361] = ~((inputs[179]) | (inputs[208]));
    assign layer0_outputs[6362] = ~(inputs[126]) | (inputs[130]);
    assign layer0_outputs[6363] = (inputs[172]) & ~(inputs[113]);
    assign layer0_outputs[6364] = inputs[121];
    assign layer0_outputs[6365] = ~(inputs[212]) | (inputs[238]);
    assign layer0_outputs[6366] = ~(inputs[114]);
    assign layer0_outputs[6367] = ~((inputs[76]) | (inputs[44]));
    assign layer0_outputs[6368] = ~(inputs[82]);
    assign layer0_outputs[6369] = inputs[193];
    assign layer0_outputs[6370] = inputs[107];
    assign layer0_outputs[6371] = ~(inputs[251]);
    assign layer0_outputs[6372] = (inputs[172]) & ~(inputs[6]);
    assign layer0_outputs[6373] = inputs[124];
    assign layer0_outputs[6374] = ~(inputs[249]);
    assign layer0_outputs[6375] = inputs[164];
    assign layer0_outputs[6376] = ~((inputs[187]) ^ (inputs[105]));
    assign layer0_outputs[6377] = ~((inputs[179]) ^ (inputs[177]));
    assign layer0_outputs[6378] = ~((inputs[216]) ^ (inputs[248]));
    assign layer0_outputs[6379] = (inputs[121]) & ~(inputs[97]);
    assign layer0_outputs[6380] = (inputs[133]) & ~(inputs[218]);
    assign layer0_outputs[6381] = ~((inputs[16]) | (inputs[29]));
    assign layer0_outputs[6382] = ~((inputs[61]) ^ (inputs[37]));
    assign layer0_outputs[6383] = ~(inputs[19]) | (inputs[208]);
    assign layer0_outputs[6384] = (inputs[155]) & ~(inputs[253]);
    assign layer0_outputs[6385] = ~(inputs[166]);
    assign layer0_outputs[6386] = ~(inputs[100]) | (inputs[253]);
    assign layer0_outputs[6387] = (inputs[89]) | (inputs[220]);
    assign layer0_outputs[6388] = (inputs[173]) & ~(inputs[100]);
    assign layer0_outputs[6389] = ~((inputs[158]) ^ (inputs[117]));
    assign layer0_outputs[6390] = ~((inputs[203]) ^ (inputs[65]));
    assign layer0_outputs[6391] = (inputs[231]) ^ (inputs[27]);
    assign layer0_outputs[6392] = (inputs[207]) ^ (inputs[149]);
    assign layer0_outputs[6393] = ~((inputs[246]) & (inputs[195]));
    assign layer0_outputs[6394] = ~(inputs[231]) | (inputs[106]);
    assign layer0_outputs[6395] = ~(inputs[75]);
    assign layer0_outputs[6396] = ~(inputs[53]) | (inputs[243]);
    assign layer0_outputs[6397] = (inputs[48]) | (inputs[149]);
    assign layer0_outputs[6398] = ~(inputs[56]);
    assign layer0_outputs[6399] = ~(inputs[94]);
    assign layer0_outputs[6400] = ~(inputs[110]) | (inputs[182]);
    assign layer0_outputs[6401] = ~(inputs[40]);
    assign layer0_outputs[6402] = (inputs[77]) | (inputs[92]);
    assign layer0_outputs[6403] = ~((inputs[55]) & (inputs[154]));
    assign layer0_outputs[6404] = ~(inputs[72]);
    assign layer0_outputs[6405] = (inputs[36]) ^ (inputs[200]);
    assign layer0_outputs[6406] = (inputs[31]) | (inputs[45]);
    assign layer0_outputs[6407] = ~(inputs[239]);
    assign layer0_outputs[6408] = inputs[72];
    assign layer0_outputs[6409] = ~((inputs[196]) & (inputs[201]));
    assign layer0_outputs[6410] = inputs[100];
    assign layer0_outputs[6411] = (inputs[179]) ^ (inputs[222]);
    assign layer0_outputs[6412] = (inputs[130]) | (inputs[153]);
    assign layer0_outputs[6413] = ~(inputs[39]) | (inputs[178]);
    assign layer0_outputs[6414] = ~((inputs[133]) ^ (inputs[131]));
    assign layer0_outputs[6415] = ~(inputs[59]) | (inputs[239]);
    assign layer0_outputs[6416] = (inputs[155]) ^ (inputs[41]);
    assign layer0_outputs[6417] = (inputs[178]) & ~(inputs[124]);
    assign layer0_outputs[6418] = ~((inputs[5]) | (inputs[43]));
    assign layer0_outputs[6419] = (inputs[171]) & ~(inputs[132]);
    assign layer0_outputs[6420] = ~(inputs[148]) | (inputs[178]);
    assign layer0_outputs[6421] = ~((inputs[250]) | (inputs[229]));
    assign layer0_outputs[6422] = inputs[8];
    assign layer0_outputs[6423] = ~((inputs[5]) ^ (inputs[45]));
    assign layer0_outputs[6424] = ~(inputs[145]);
    assign layer0_outputs[6425] = inputs[76];
    assign layer0_outputs[6426] = ~(inputs[153]) | (inputs[62]);
    assign layer0_outputs[6427] = ~(inputs[23]) | (inputs[190]);
    assign layer0_outputs[6428] = ~(inputs[36]) | (inputs[187]);
    assign layer0_outputs[6429] = ~((inputs[163]) ^ (inputs[198]));
    assign layer0_outputs[6430] = (inputs[36]) & ~(inputs[234]);
    assign layer0_outputs[6431] = ~((inputs[194]) | (inputs[11]));
    assign layer0_outputs[6432] = ~(inputs[222]) | (inputs[31]);
    assign layer0_outputs[6433] = (inputs[61]) ^ (inputs[28]);
    assign layer0_outputs[6434] = ~(inputs[137]) | (inputs[155]);
    assign layer0_outputs[6435] = (inputs[121]) | (inputs[35]);
    assign layer0_outputs[6436] = ~(inputs[62]);
    assign layer0_outputs[6437] = (inputs[203]) & ~(inputs[28]);
    assign layer0_outputs[6438] = ~(inputs[180]);
    assign layer0_outputs[6439] = (inputs[109]) & ~(inputs[12]);
    assign layer0_outputs[6440] = ~(inputs[219]);
    assign layer0_outputs[6441] = (inputs[90]) & ~(inputs[71]);
    assign layer0_outputs[6442] = ~(inputs[246]) | (inputs[14]);
    assign layer0_outputs[6443] = inputs[250];
    assign layer0_outputs[6444] = ~(inputs[171]) | (inputs[223]);
    assign layer0_outputs[6445] = (inputs[64]) & ~(inputs[131]);
    assign layer0_outputs[6446] = (inputs[42]) & (inputs[85]);
    assign layer0_outputs[6447] = ~(inputs[139]);
    assign layer0_outputs[6448] = inputs[113];
    assign layer0_outputs[6449] = ~(inputs[140]);
    assign layer0_outputs[6450] = ~((inputs[132]) ^ (inputs[137]));
    assign layer0_outputs[6451] = (inputs[178]) | (inputs[81]);
    assign layer0_outputs[6452] = ~(inputs[182]);
    assign layer0_outputs[6453] = inputs[95];
    assign layer0_outputs[6454] = ~(inputs[118]) | (inputs[4]);
    assign layer0_outputs[6455] = ~(inputs[31]) | (inputs[52]);
    assign layer0_outputs[6456] = inputs[59];
    assign layer0_outputs[6457] = ~(inputs[1]);
    assign layer0_outputs[6458] = (inputs[18]) | (inputs[56]);
    assign layer0_outputs[6459] = (inputs[254]) ^ (inputs[207]);
    assign layer0_outputs[6460] = (inputs[182]) | (inputs[44]);
    assign layer0_outputs[6461] = (inputs[84]) ^ (inputs[224]);
    assign layer0_outputs[6462] = (inputs[126]) | (inputs[18]);
    assign layer0_outputs[6463] = (inputs[223]) | (inputs[84]);
    assign layer0_outputs[6464] = (inputs[23]) | (inputs[36]);
    assign layer0_outputs[6465] = (inputs[214]) & (inputs[132]);
    assign layer0_outputs[6466] = (inputs[95]) ^ (inputs[57]);
    assign layer0_outputs[6467] = (inputs[199]) & ~(inputs[86]);
    assign layer0_outputs[6468] = (inputs[175]) & ~(inputs[26]);
    assign layer0_outputs[6469] = (inputs[191]) | (inputs[8]);
    assign layer0_outputs[6470] = ~((inputs[249]) ^ (inputs[231]));
    assign layer0_outputs[6471] = inputs[60];
    assign layer0_outputs[6472] = (inputs[2]) ^ (inputs[15]);
    assign layer0_outputs[6473] = (inputs[223]) | (inputs[62]);
    assign layer0_outputs[6474] = (inputs[230]) | (inputs[229]);
    assign layer0_outputs[6475] = inputs[41];
    assign layer0_outputs[6476] = inputs[62];
    assign layer0_outputs[6477] = (inputs[211]) | (inputs[143]);
    assign layer0_outputs[6478] = ~((inputs[143]) ^ (inputs[139]));
    assign layer0_outputs[6479] = (inputs[152]) | (inputs[237]);
    assign layer0_outputs[6480] = ~(inputs[166]);
    assign layer0_outputs[6481] = ~((inputs[12]) | (inputs[94]));
    assign layer0_outputs[6482] = inputs[44];
    assign layer0_outputs[6483] = ~((inputs[175]) ^ (inputs[253]));
    assign layer0_outputs[6484] = 1'b0;
    assign layer0_outputs[6485] = ~(inputs[200]) | (inputs[239]);
    assign layer0_outputs[6486] = (inputs[78]) ^ (inputs[179]);
    assign layer0_outputs[6487] = 1'b1;
    assign layer0_outputs[6488] = (inputs[71]) & ~(inputs[138]);
    assign layer0_outputs[6489] = ~(inputs[117]);
    assign layer0_outputs[6490] = inputs[114];
    assign layer0_outputs[6491] = inputs[229];
    assign layer0_outputs[6492] = ~((inputs[238]) ^ (inputs[47]));
    assign layer0_outputs[6493] = ~(inputs[162]);
    assign layer0_outputs[6494] = ~(inputs[182]);
    assign layer0_outputs[6495] = ~(inputs[5]);
    assign layer0_outputs[6496] = ~(inputs[205]);
    assign layer0_outputs[6497] = ~(inputs[65]);
    assign layer0_outputs[6498] = (inputs[53]) | (inputs[25]);
    assign layer0_outputs[6499] = ~(inputs[97]);
    assign layer0_outputs[6500] = (inputs[165]) & ~(inputs[240]);
    assign layer0_outputs[6501] = ~((inputs[30]) | (inputs[190]));
    assign layer0_outputs[6502] = (inputs[109]) | (inputs[131]);
    assign layer0_outputs[6503] = ~(inputs[162]);
    assign layer0_outputs[6504] = 1'b0;
    assign layer0_outputs[6505] = ~((inputs[189]) & (inputs[5]));
    assign layer0_outputs[6506] = inputs[123];
    assign layer0_outputs[6507] = (inputs[21]) | (inputs[33]);
    assign layer0_outputs[6508] = ~(inputs[119]);
    assign layer0_outputs[6509] = inputs[36];
    assign layer0_outputs[6510] = ~(inputs[68]);
    assign layer0_outputs[6511] = (inputs[209]) & ~(inputs[71]);
    assign layer0_outputs[6512] = ~(inputs[130]);
    assign layer0_outputs[6513] = ~(inputs[248]);
    assign layer0_outputs[6514] = ~(inputs[143]) | (inputs[32]);
    assign layer0_outputs[6515] = (inputs[243]) & (inputs[219]);
    assign layer0_outputs[6516] = ~(inputs[231]);
    assign layer0_outputs[6517] = inputs[197];
    assign layer0_outputs[6518] = ~(inputs[222]) | (inputs[15]);
    assign layer0_outputs[6519] = ~(inputs[200]);
    assign layer0_outputs[6520] = ~(inputs[149]) | (inputs[106]);
    assign layer0_outputs[6521] = (inputs[154]) | (inputs[81]);
    assign layer0_outputs[6522] = (inputs[170]) | (inputs[128]);
    assign layer0_outputs[6523] = ~((inputs[72]) ^ (inputs[15]));
    assign layer0_outputs[6524] = (inputs[142]) | (inputs[11]);
    assign layer0_outputs[6525] = ~(inputs[181]);
    assign layer0_outputs[6526] = ~((inputs[204]) | (inputs[217]));
    assign layer0_outputs[6527] = ~((inputs[126]) ^ (inputs[155]));
    assign layer0_outputs[6528] = (inputs[212]) & (inputs[76]);
    assign layer0_outputs[6529] = ~((inputs[191]) ^ (inputs[110]));
    assign layer0_outputs[6530] = (inputs[36]) & ~(inputs[165]);
    assign layer0_outputs[6531] = ~(inputs[56]) | (inputs[4]);
    assign layer0_outputs[6532] = inputs[123];
    assign layer0_outputs[6533] = (inputs[179]) & (inputs[244]);
    assign layer0_outputs[6534] = (inputs[170]) | (inputs[175]);
    assign layer0_outputs[6535] = inputs[91];
    assign layer0_outputs[6536] = (inputs[248]) | (inputs[125]);
    assign layer0_outputs[6537] = ~((inputs[81]) & (inputs[134]));
    assign layer0_outputs[6538] = inputs[157];
    assign layer0_outputs[6539] = ~(inputs[139]) | (inputs[42]);
    assign layer0_outputs[6540] = ~(inputs[70]);
    assign layer0_outputs[6541] = ~(inputs[209]);
    assign layer0_outputs[6542] = ~(inputs[138]) | (inputs[214]);
    assign layer0_outputs[6543] = ~(inputs[69]);
    assign layer0_outputs[6544] = 1'b1;
    assign layer0_outputs[6545] = ~((inputs[85]) | (inputs[115]));
    assign layer0_outputs[6546] = (inputs[133]) ^ (inputs[98]);
    assign layer0_outputs[6547] = ~(inputs[184]);
    assign layer0_outputs[6548] = ~(inputs[89]);
    assign layer0_outputs[6549] = inputs[113];
    assign layer0_outputs[6550] = ~(inputs[211]) | (inputs[58]);
    assign layer0_outputs[6551] = ~(inputs[242]);
    assign layer0_outputs[6552] = (inputs[40]) | (inputs[62]);
    assign layer0_outputs[6553] = (inputs[87]) ^ (inputs[100]);
    assign layer0_outputs[6554] = (inputs[199]) | (inputs[134]);
    assign layer0_outputs[6555] = inputs[115];
    assign layer0_outputs[6556] = (inputs[141]) | (inputs[188]);
    assign layer0_outputs[6557] = inputs[126];
    assign layer0_outputs[6558] = ~((inputs[2]) | (inputs[1]));
    assign layer0_outputs[6559] = (inputs[211]) | (inputs[160]);
    assign layer0_outputs[6560] = ~(inputs[178]);
    assign layer0_outputs[6561] = inputs[41];
    assign layer0_outputs[6562] = (inputs[195]) & ~(inputs[62]);
    assign layer0_outputs[6563] = ~((inputs[244]) | (inputs[228]));
    assign layer0_outputs[6564] = (inputs[87]) & ~(inputs[185]);
    assign layer0_outputs[6565] = inputs[193];
    assign layer0_outputs[6566] = (inputs[26]) & ~(inputs[133]);
    assign layer0_outputs[6567] = ~((inputs[91]) ^ (inputs[142]));
    assign layer0_outputs[6568] = (inputs[7]) & ~(inputs[174]);
    assign layer0_outputs[6569] = inputs[173];
    assign layer0_outputs[6570] = (inputs[171]) & ~(inputs[53]);
    assign layer0_outputs[6571] = (inputs[22]) | (inputs[33]);
    assign layer0_outputs[6572] = inputs[134];
    assign layer0_outputs[6573] = ~((inputs[80]) | (inputs[99]));
    assign layer0_outputs[6574] = ~((inputs[195]) | (inputs[50]));
    assign layer0_outputs[6575] = (inputs[105]) & ~(inputs[192]);
    assign layer0_outputs[6576] = ~(inputs[136]);
    assign layer0_outputs[6577] = (inputs[2]) | (inputs[231]);
    assign layer0_outputs[6578] = ~(inputs[108]);
    assign layer0_outputs[6579] = (inputs[175]) | (inputs[212]);
    assign layer0_outputs[6580] = (inputs[121]) | (inputs[255]);
    assign layer0_outputs[6581] = ~((inputs[210]) | (inputs[213]));
    assign layer0_outputs[6582] = ~(inputs[98]);
    assign layer0_outputs[6583] = ~((inputs[19]) | (inputs[150]));
    assign layer0_outputs[6584] = (inputs[75]) & (inputs[25]);
    assign layer0_outputs[6585] = ~((inputs[119]) | (inputs[15]));
    assign layer0_outputs[6586] = 1'b0;
    assign layer0_outputs[6587] = (inputs[166]) | (inputs[80]);
    assign layer0_outputs[6588] = (inputs[120]) | (inputs[14]);
    assign layer0_outputs[6589] = ~(inputs[135]);
    assign layer0_outputs[6590] = ~((inputs[156]) | (inputs[216]));
    assign layer0_outputs[6591] = ~(inputs[127]) | (inputs[190]);
    assign layer0_outputs[6592] = ~((inputs[213]) | (inputs[223]));
    assign layer0_outputs[6593] = (inputs[158]) ^ (inputs[118]);
    assign layer0_outputs[6594] = (inputs[62]) ^ (inputs[36]);
    assign layer0_outputs[6595] = inputs[29];
    assign layer0_outputs[6596] = ~((inputs[144]) ^ (inputs[46]));
    assign layer0_outputs[6597] = ~(inputs[77]);
    assign layer0_outputs[6598] = inputs[191];
    assign layer0_outputs[6599] = (inputs[177]) | (inputs[17]);
    assign layer0_outputs[6600] = inputs[91];
    assign layer0_outputs[6601] = ~((inputs[233]) | (inputs[44]));
    assign layer0_outputs[6602] = ~(inputs[245]);
    assign layer0_outputs[6603] = (inputs[221]) & ~(inputs[128]);
    assign layer0_outputs[6604] = ~(inputs[133]);
    assign layer0_outputs[6605] = ~(inputs[158]) | (inputs[254]);
    assign layer0_outputs[6606] = inputs[113];
    assign layer0_outputs[6607] = ~(inputs[8]) | (inputs[212]);
    assign layer0_outputs[6608] = ~(inputs[52]);
    assign layer0_outputs[6609] = (inputs[157]) | (inputs[28]);
    assign layer0_outputs[6610] = (inputs[24]) & ~(inputs[146]);
    assign layer0_outputs[6611] = inputs[69];
    assign layer0_outputs[6612] = inputs[197];
    assign layer0_outputs[6613] = (inputs[205]) ^ (inputs[187]);
    assign layer0_outputs[6614] = ~((inputs[102]) & (inputs[104]));
    assign layer0_outputs[6615] = ~(inputs[245]) | (inputs[3]);
    assign layer0_outputs[6616] = inputs[176];
    assign layer0_outputs[6617] = (inputs[164]) & (inputs[195]);
    assign layer0_outputs[6618] = ~((inputs[89]) ^ (inputs[148]));
    assign layer0_outputs[6619] = (inputs[125]) ^ (inputs[16]);
    assign layer0_outputs[6620] = ~(inputs[161]);
    assign layer0_outputs[6621] = ~((inputs[237]) | (inputs[243]));
    assign layer0_outputs[6622] = ~((inputs[97]) ^ (inputs[47]));
    assign layer0_outputs[6623] = (inputs[141]) | (inputs[198]);
    assign layer0_outputs[6624] = inputs[194];
    assign layer0_outputs[6625] = (inputs[239]) ^ (inputs[224]);
    assign layer0_outputs[6626] = 1'b1;
    assign layer0_outputs[6627] = (inputs[77]) & ~(inputs[18]);
    assign layer0_outputs[6628] = (inputs[20]) ^ (inputs[193]);
    assign layer0_outputs[6629] = ~(inputs[85]);
    assign layer0_outputs[6630] = inputs[176];
    assign layer0_outputs[6631] = ~(inputs[202]);
    assign layer0_outputs[6632] = ~(inputs[232]);
    assign layer0_outputs[6633] = ~((inputs[143]) | (inputs[197]));
    assign layer0_outputs[6634] = ~(inputs[7]);
    assign layer0_outputs[6635] = ~(inputs[14]);
    assign layer0_outputs[6636] = ~((inputs[214]) | (inputs[247]));
    assign layer0_outputs[6637] = inputs[139];
    assign layer0_outputs[6638] = ~((inputs[127]) | (inputs[176]));
    assign layer0_outputs[6639] = ~(inputs[102]);
    assign layer0_outputs[6640] = (inputs[214]) ^ (inputs[246]);
    assign layer0_outputs[6641] = (inputs[66]) | (inputs[232]);
    assign layer0_outputs[6642] = inputs[139];
    assign layer0_outputs[6643] = ~(inputs[180]);
    assign layer0_outputs[6644] = ~(inputs[244]) | (inputs[29]);
    assign layer0_outputs[6645] = ~((inputs[75]) | (inputs[6]));
    assign layer0_outputs[6646] = (inputs[231]) & ~(inputs[30]);
    assign layer0_outputs[6647] = ~(inputs[28]);
    assign layer0_outputs[6648] = inputs[176];
    assign layer0_outputs[6649] = (inputs[174]) & (inputs[250]);
    assign layer0_outputs[6650] = ~((inputs[106]) | (inputs[14]));
    assign layer0_outputs[6651] = ~((inputs[88]) ^ (inputs[124]));
    assign layer0_outputs[6652] = ~(inputs[68]);
    assign layer0_outputs[6653] = ~(inputs[198]);
    assign layer0_outputs[6654] = ~((inputs[19]) | (inputs[127]));
    assign layer0_outputs[6655] = (inputs[141]) & (inputs[105]);
    assign layer0_outputs[6656] = ~((inputs[125]) | (inputs[17]));
    assign layer0_outputs[6657] = inputs[32];
    assign layer0_outputs[6658] = (inputs[24]) & ~(inputs[130]);
    assign layer0_outputs[6659] = (inputs[85]) & ~(inputs[32]);
    assign layer0_outputs[6660] = ~(inputs[85]);
    assign layer0_outputs[6661] = ~((inputs[210]) ^ (inputs[179]));
    assign layer0_outputs[6662] = (inputs[220]) & (inputs[251]);
    assign layer0_outputs[6663] = ~((inputs[126]) | (inputs[197]));
    assign layer0_outputs[6664] = ~((inputs[228]) ^ (inputs[136]));
    assign layer0_outputs[6665] = ~((inputs[245]) | (inputs[239]));
    assign layer0_outputs[6666] = ~(inputs[41]) | (inputs[11]);
    assign layer0_outputs[6667] = inputs[85];
    assign layer0_outputs[6668] = ~((inputs[164]) | (inputs[198]));
    assign layer0_outputs[6669] = ~((inputs[95]) | (inputs[247]));
    assign layer0_outputs[6670] = inputs[196];
    assign layer0_outputs[6671] = ~(inputs[213]) | (inputs[89]);
    assign layer0_outputs[6672] = ~(inputs[142]);
    assign layer0_outputs[6673] = inputs[212];
    assign layer0_outputs[6674] = ~(inputs[164]);
    assign layer0_outputs[6675] = ~((inputs[201]) | (inputs[196]));
    assign layer0_outputs[6676] = (inputs[160]) | (inputs[206]);
    assign layer0_outputs[6677] = (inputs[211]) ^ (inputs[177]);
    assign layer0_outputs[6678] = (inputs[106]) & ~(inputs[31]);
    assign layer0_outputs[6679] = ~(inputs[23]);
    assign layer0_outputs[6680] = ~((inputs[15]) ^ (inputs[168]));
    assign layer0_outputs[6681] = inputs[115];
    assign layer0_outputs[6682] = (inputs[46]) | (inputs[10]);
    assign layer0_outputs[6683] = (inputs[59]) | (inputs[109]);
    assign layer0_outputs[6684] = ~(inputs[124]) | (inputs[243]);
    assign layer0_outputs[6685] = ~((inputs[22]) & (inputs[226]));
    assign layer0_outputs[6686] = (inputs[8]) ^ (inputs[85]);
    assign layer0_outputs[6687] = ~((inputs[232]) & (inputs[91]));
    assign layer0_outputs[6688] = ~(inputs[157]) | (inputs[14]);
    assign layer0_outputs[6689] = (inputs[103]) ^ (inputs[208]);
    assign layer0_outputs[6690] = (inputs[222]) | (inputs[250]);
    assign layer0_outputs[6691] = (inputs[147]) ^ (inputs[234]);
    assign layer0_outputs[6692] = (inputs[1]) ^ (inputs[108]);
    assign layer0_outputs[6693] = inputs[48];
    assign layer0_outputs[6694] = ~((inputs[196]) ^ (inputs[7]));
    assign layer0_outputs[6695] = ~(inputs[199]);
    assign layer0_outputs[6696] = ~(inputs[86]);
    assign layer0_outputs[6697] = (inputs[10]) & ~(inputs[210]);
    assign layer0_outputs[6698] = ~(inputs[253]);
    assign layer0_outputs[6699] = ~((inputs[175]) ^ (inputs[160]));
    assign layer0_outputs[6700] = inputs[125];
    assign layer0_outputs[6701] = ~((inputs[120]) ^ (inputs[69]));
    assign layer0_outputs[6702] = ~(inputs[121]);
    assign layer0_outputs[6703] = inputs[84];
    assign layer0_outputs[6704] = inputs[131];
    assign layer0_outputs[6705] = ~((inputs[9]) ^ (inputs[208]));
    assign layer0_outputs[6706] = ~((inputs[242]) ^ (inputs[170]));
    assign layer0_outputs[6707] = ~(inputs[86]) | (inputs[237]);
    assign layer0_outputs[6708] = inputs[54];
    assign layer0_outputs[6709] = (inputs[14]) & ~(inputs[177]);
    assign layer0_outputs[6710] = inputs[181];
    assign layer0_outputs[6711] = (inputs[199]) & ~(inputs[76]);
    assign layer0_outputs[6712] = ~((inputs[224]) | (inputs[184]));
    assign layer0_outputs[6713] = ~(inputs[22]);
    assign layer0_outputs[6714] = (inputs[4]) | (inputs[94]);
    assign layer0_outputs[6715] = (inputs[135]) & ~(inputs[70]);
    assign layer0_outputs[6716] = ~(inputs[136]) | (inputs[100]);
    assign layer0_outputs[6717] = ~(inputs[58]);
    assign layer0_outputs[6718] = (inputs[20]) & ~(inputs[85]);
    assign layer0_outputs[6719] = (inputs[126]) | (inputs[142]);
    assign layer0_outputs[6720] = ~((inputs[190]) | (inputs[80]));
    assign layer0_outputs[6721] = (inputs[85]) & ~(inputs[78]);
    assign layer0_outputs[6722] = ~((inputs[17]) ^ (inputs[81]));
    assign layer0_outputs[6723] = (inputs[43]) & (inputs[104]);
    assign layer0_outputs[6724] = inputs[69];
    assign layer0_outputs[6725] = ~((inputs[8]) ^ (inputs[159]));
    assign layer0_outputs[6726] = ~(inputs[6]);
    assign layer0_outputs[6727] = ~((inputs[181]) | (inputs[49]));
    assign layer0_outputs[6728] = inputs[212];
    assign layer0_outputs[6729] = inputs[201];
    assign layer0_outputs[6730] = ~(inputs[36]);
    assign layer0_outputs[6731] = ~((inputs[42]) ^ (inputs[31]));
    assign layer0_outputs[6732] = ~((inputs[26]) ^ (inputs[102]));
    assign layer0_outputs[6733] = inputs[233];
    assign layer0_outputs[6734] = inputs[149];
    assign layer0_outputs[6735] = inputs[189];
    assign layer0_outputs[6736] = ~(inputs[58]) | (inputs[233]);
    assign layer0_outputs[6737] = ~(inputs[167]);
    assign layer0_outputs[6738] = ~(inputs[232]);
    assign layer0_outputs[6739] = ~(inputs[44]) | (inputs[135]);
    assign layer0_outputs[6740] = (inputs[34]) ^ (inputs[151]);
    assign layer0_outputs[6741] = (inputs[7]) & ~(inputs[197]);
    assign layer0_outputs[6742] = inputs[207];
    assign layer0_outputs[6743] = inputs[87];
    assign layer0_outputs[6744] = inputs[135];
    assign layer0_outputs[6745] = ~(inputs[243]);
    assign layer0_outputs[6746] = ~(inputs[23]) | (inputs[146]);
    assign layer0_outputs[6747] = (inputs[154]) & ~(inputs[141]);
    assign layer0_outputs[6748] = (inputs[22]) | (inputs[236]);
    assign layer0_outputs[6749] = ~(inputs[99]);
    assign layer0_outputs[6750] = ~(inputs[106]);
    assign layer0_outputs[6751] = ~((inputs[130]) | (inputs[214]));
    assign layer0_outputs[6752] = (inputs[55]) ^ (inputs[71]);
    assign layer0_outputs[6753] = ~(inputs[179]);
    assign layer0_outputs[6754] = (inputs[62]) | (inputs[80]);
    assign layer0_outputs[6755] = ~((inputs[160]) | (inputs[142]));
    assign layer0_outputs[6756] = ~((inputs[0]) ^ (inputs[7]));
    assign layer0_outputs[6757] = ~((inputs[123]) ^ (inputs[89]));
    assign layer0_outputs[6758] = ~(inputs[36]) | (inputs[223]);
    assign layer0_outputs[6759] = ~(inputs[248]);
    assign layer0_outputs[6760] = ~((inputs[97]) & (inputs[30]));
    assign layer0_outputs[6761] = ~(inputs[53]);
    assign layer0_outputs[6762] = ~((inputs[108]) | (inputs[18]));
    assign layer0_outputs[6763] = inputs[69];
    assign layer0_outputs[6764] = ~(inputs[208]);
    assign layer0_outputs[6765] = ~((inputs[88]) & (inputs[172]));
    assign layer0_outputs[6766] = (inputs[245]) | (inputs[249]);
    assign layer0_outputs[6767] = ~((inputs[109]) ^ (inputs[167]));
    assign layer0_outputs[6768] = inputs[254];
    assign layer0_outputs[6769] = (inputs[222]) ^ (inputs[121]);
    assign layer0_outputs[6770] = (inputs[16]) ^ (inputs[52]);
    assign layer0_outputs[6771] = ~(inputs[87]);
    assign layer0_outputs[6772] = ~((inputs[43]) ^ (inputs[70]));
    assign layer0_outputs[6773] = inputs[181];
    assign layer0_outputs[6774] = ~(inputs[229]);
    assign layer0_outputs[6775] = (inputs[51]) | (inputs[31]);
    assign layer0_outputs[6776] = (inputs[36]) ^ (inputs[82]);
    assign layer0_outputs[6777] = inputs[173];
    assign layer0_outputs[6778] = (inputs[205]) & ~(inputs[239]);
    assign layer0_outputs[6779] = (inputs[218]) & ~(inputs[136]);
    assign layer0_outputs[6780] = ~(inputs[187]);
    assign layer0_outputs[6781] = (inputs[88]) & ~(inputs[210]);
    assign layer0_outputs[6782] = (inputs[139]) & ~(inputs[174]);
    assign layer0_outputs[6783] = (inputs[138]) & ~(inputs[75]);
    assign layer0_outputs[6784] = ~((inputs[35]) | (inputs[80]));
    assign layer0_outputs[6785] = ~((inputs[160]) | (inputs[141]));
    assign layer0_outputs[6786] = ~((inputs[132]) | (inputs[62]));
    assign layer0_outputs[6787] = ~(inputs[23]);
    assign layer0_outputs[6788] = ~((inputs[197]) ^ (inputs[96]));
    assign layer0_outputs[6789] = ~((inputs[205]) | (inputs[215]));
    assign layer0_outputs[6790] = inputs[232];
    assign layer0_outputs[6791] = inputs[17];
    assign layer0_outputs[6792] = inputs[215];
    assign layer0_outputs[6793] = (inputs[187]) | (inputs[169]);
    assign layer0_outputs[6794] = ~(inputs[113]);
    assign layer0_outputs[6795] = inputs[89];
    assign layer0_outputs[6796] = (inputs[137]) ^ (inputs[148]);
    assign layer0_outputs[6797] = (inputs[20]) & ~(inputs[159]);
    assign layer0_outputs[6798] = ~((inputs[201]) | (inputs[232]));
    assign layer0_outputs[6799] = ~(inputs[187]) | (inputs[110]);
    assign layer0_outputs[6800] = inputs[34];
    assign layer0_outputs[6801] = ~(inputs[94]) | (inputs[82]);
    assign layer0_outputs[6802] = ~((inputs[119]) | (inputs[219]));
    assign layer0_outputs[6803] = ~(inputs[110]);
    assign layer0_outputs[6804] = ~((inputs[145]) & (inputs[211]));
    assign layer0_outputs[6805] = inputs[69];
    assign layer0_outputs[6806] = (inputs[215]) | (inputs[115]);
    assign layer0_outputs[6807] = (inputs[114]) & ~(inputs[66]);
    assign layer0_outputs[6808] = ~(inputs[109]);
    assign layer0_outputs[6809] = inputs[82];
    assign layer0_outputs[6810] = ~(inputs[66]) | (inputs[250]);
    assign layer0_outputs[6811] = inputs[98];
    assign layer0_outputs[6812] = (inputs[32]) & ~(inputs[225]);
    assign layer0_outputs[6813] = ~((inputs[77]) & (inputs[106]));
    assign layer0_outputs[6814] = (inputs[238]) | (inputs[5]);
    assign layer0_outputs[6815] = (inputs[215]) & ~(inputs[33]);
    assign layer0_outputs[6816] = ~(inputs[67]);
    assign layer0_outputs[6817] = ~(inputs[180]) | (inputs[15]);
    assign layer0_outputs[6818] = ~(inputs[231]) | (inputs[208]);
    assign layer0_outputs[6819] = ~(inputs[60]) | (inputs[194]);
    assign layer0_outputs[6820] = inputs[128];
    assign layer0_outputs[6821] = 1'b0;
    assign layer0_outputs[6822] = (inputs[131]) & ~(inputs[164]);
    assign layer0_outputs[6823] = ~((inputs[54]) & (inputs[175]));
    assign layer0_outputs[6824] = (inputs[49]) & ~(inputs[121]);
    assign layer0_outputs[6825] = ~(inputs[182]);
    assign layer0_outputs[6826] = ~(inputs[204]) | (inputs[168]);
    assign layer0_outputs[6827] = inputs[179];
    assign layer0_outputs[6828] = (inputs[159]) | (inputs[170]);
    assign layer0_outputs[6829] = inputs[48];
    assign layer0_outputs[6830] = (inputs[210]) | (inputs[192]);
    assign layer0_outputs[6831] = ~((inputs[134]) | (inputs[234]));
    assign layer0_outputs[6832] = ~(inputs[255]);
    assign layer0_outputs[6833] = ~(inputs[106]);
    assign layer0_outputs[6834] = ~(inputs[232]) | (inputs[86]);
    assign layer0_outputs[6835] = (inputs[179]) | (inputs[168]);
    assign layer0_outputs[6836] = (inputs[5]) | (inputs[207]);
    assign layer0_outputs[6837] = ~(inputs[216]);
    assign layer0_outputs[6838] = ~(inputs[146]);
    assign layer0_outputs[6839] = ~((inputs[244]) | (inputs[19]));
    assign layer0_outputs[6840] = ~(inputs[154]) | (inputs[147]);
    assign layer0_outputs[6841] = inputs[13];
    assign layer0_outputs[6842] = (inputs[105]) & (inputs[84]);
    assign layer0_outputs[6843] = (inputs[207]) | (inputs[150]);
    assign layer0_outputs[6844] = (inputs[8]) ^ (inputs[130]);
    assign layer0_outputs[6845] = ~((inputs[152]) | (inputs[253]));
    assign layer0_outputs[6846] = ~((inputs[60]) ^ (inputs[49]));
    assign layer0_outputs[6847] = inputs[73];
    assign layer0_outputs[6848] = 1'b0;
    assign layer0_outputs[6849] = inputs[92];
    assign layer0_outputs[6850] = (inputs[144]) | (inputs[155]);
    assign layer0_outputs[6851] = 1'b0;
    assign layer0_outputs[6852] = ~(inputs[19]) | (inputs[175]);
    assign layer0_outputs[6853] = ~((inputs[54]) ^ (inputs[51]));
    assign layer0_outputs[6854] = (inputs[15]) | (inputs[13]);
    assign layer0_outputs[6855] = ~(inputs[201]);
    assign layer0_outputs[6856] = ~((inputs[62]) | (inputs[41]));
    assign layer0_outputs[6857] = (inputs[80]) & (inputs[97]);
    assign layer0_outputs[6858] = inputs[164];
    assign layer0_outputs[6859] = (inputs[81]) | (inputs[173]);
    assign layer0_outputs[6860] = ~(inputs[102]);
    assign layer0_outputs[6861] = inputs[163];
    assign layer0_outputs[6862] = (inputs[99]) ^ (inputs[101]);
    assign layer0_outputs[6863] = ~((inputs[195]) | (inputs[192]));
    assign layer0_outputs[6864] = inputs[225];
    assign layer0_outputs[6865] = (inputs[206]) ^ (inputs[18]);
    assign layer0_outputs[6866] = (inputs[56]) | (inputs[23]);
    assign layer0_outputs[6867] = ~((inputs[134]) | (inputs[251]));
    assign layer0_outputs[6868] = ~(inputs[70]);
    assign layer0_outputs[6869] = ~((inputs[172]) ^ (inputs[146]));
    assign layer0_outputs[6870] = inputs[113];
    assign layer0_outputs[6871] = (inputs[137]) | (inputs[228]);
    assign layer0_outputs[6872] = inputs[218];
    assign layer0_outputs[6873] = inputs[124];
    assign layer0_outputs[6874] = ~(inputs[79]);
    assign layer0_outputs[6875] = (inputs[40]) & ~(inputs[98]);
    assign layer0_outputs[6876] = (inputs[247]) ^ (inputs[184]);
    assign layer0_outputs[6877] = ~(inputs[71]);
    assign layer0_outputs[6878] = (inputs[126]) | (inputs[55]);
    assign layer0_outputs[6879] = ~((inputs[197]) | (inputs[5]));
    assign layer0_outputs[6880] = ~((inputs[219]) | (inputs[223]));
    assign layer0_outputs[6881] = inputs[219];
    assign layer0_outputs[6882] = (inputs[43]) & ~(inputs[5]);
    assign layer0_outputs[6883] = ~(inputs[147]);
    assign layer0_outputs[6884] = (inputs[74]) | (inputs[98]);
    assign layer0_outputs[6885] = inputs[144];
    assign layer0_outputs[6886] = (inputs[251]) | (inputs[74]);
    assign layer0_outputs[6887] = (inputs[56]) | (inputs[84]);
    assign layer0_outputs[6888] = (inputs[149]) | (inputs[193]);
    assign layer0_outputs[6889] = ~(inputs[28]);
    assign layer0_outputs[6890] = ~((inputs[122]) | (inputs[20]));
    assign layer0_outputs[6891] = inputs[186];
    assign layer0_outputs[6892] = ~((inputs[106]) | (inputs[154]));
    assign layer0_outputs[6893] = (inputs[212]) | (inputs[49]);
    assign layer0_outputs[6894] = (inputs[211]) | (inputs[176]);
    assign layer0_outputs[6895] = (inputs[76]) ^ (inputs[90]);
    assign layer0_outputs[6896] = inputs[35];
    assign layer0_outputs[6897] = ~((inputs[228]) ^ (inputs[10]));
    assign layer0_outputs[6898] = (inputs[214]) | (inputs[6]);
    assign layer0_outputs[6899] = ~(inputs[82]);
    assign layer0_outputs[6900] = ~((inputs[87]) | (inputs[187]));
    assign layer0_outputs[6901] = ~(inputs[211]);
    assign layer0_outputs[6902] = ~(inputs[85]);
    assign layer0_outputs[6903] = (inputs[222]) | (inputs[142]);
    assign layer0_outputs[6904] = ~((inputs[92]) | (inputs[209]));
    assign layer0_outputs[6905] = inputs[166];
    assign layer0_outputs[6906] = 1'b1;
    assign layer0_outputs[6907] = (inputs[175]) ^ (inputs[9]);
    assign layer0_outputs[6908] = ~(inputs[187]) | (inputs[31]);
    assign layer0_outputs[6909] = (inputs[15]) ^ (inputs[217]);
    assign layer0_outputs[6910] = ~(inputs[154]);
    assign layer0_outputs[6911] = (inputs[7]) | (inputs[111]);
    assign layer0_outputs[6912] = ~(inputs[131]);
    assign layer0_outputs[6913] = ~((inputs[103]) | (inputs[87]));
    assign layer0_outputs[6914] = ~(inputs[88]);
    assign layer0_outputs[6915] = (inputs[50]) ^ (inputs[238]);
    assign layer0_outputs[6916] = ~(inputs[243]);
    assign layer0_outputs[6917] = ~(inputs[46]);
    assign layer0_outputs[6918] = ~((inputs[197]) | (inputs[82]));
    assign layer0_outputs[6919] = ~((inputs[114]) ^ (inputs[107]));
    assign layer0_outputs[6920] = ~((inputs[223]) & (inputs[224]));
    assign layer0_outputs[6921] = ~(inputs[165]) | (inputs[222]);
    assign layer0_outputs[6922] = ~((inputs[83]) ^ (inputs[16]));
    assign layer0_outputs[6923] = (inputs[94]) ^ (inputs[201]);
    assign layer0_outputs[6924] = ~(inputs[165]);
    assign layer0_outputs[6925] = ~(inputs[71]);
    assign layer0_outputs[6926] = ~((inputs[83]) & (inputs[105]));
    assign layer0_outputs[6927] = 1'b0;
    assign layer0_outputs[6928] = ~(inputs[230]);
    assign layer0_outputs[6929] = ~(inputs[101]) | (inputs[21]);
    assign layer0_outputs[6930] = ~(inputs[113]);
    assign layer0_outputs[6931] = (inputs[25]) ^ (inputs[98]);
    assign layer0_outputs[6932] = (inputs[185]) & ~(inputs[61]);
    assign layer0_outputs[6933] = ~(inputs[86]);
    assign layer0_outputs[6934] = ~(inputs[151]);
    assign layer0_outputs[6935] = 1'b1;
    assign layer0_outputs[6936] = ~((inputs[36]) | (inputs[21]));
    assign layer0_outputs[6937] = ~(inputs[64]);
    assign layer0_outputs[6938] = (inputs[97]) ^ (inputs[76]);
    assign layer0_outputs[6939] = ~(inputs[119]);
    assign layer0_outputs[6940] = ~(inputs[60]);
    assign layer0_outputs[6941] = ~(inputs[36]);
    assign layer0_outputs[6942] = (inputs[210]) & ~(inputs[152]);
    assign layer0_outputs[6943] = ~((inputs[162]) | (inputs[29]));
    assign layer0_outputs[6944] = inputs[99];
    assign layer0_outputs[6945] = ~((inputs[115]) & (inputs[122]));
    assign layer0_outputs[6946] = ~(inputs[87]) | (inputs[239]);
    assign layer0_outputs[6947] = ~(inputs[20]);
    assign layer0_outputs[6948] = ~((inputs[253]) | (inputs[133]));
    assign layer0_outputs[6949] = (inputs[136]) | (inputs[233]);
    assign layer0_outputs[6950] = ~(inputs[167]) | (inputs[16]);
    assign layer0_outputs[6951] = (inputs[157]) & ~(inputs[10]);
    assign layer0_outputs[6952] = (inputs[95]) ^ (inputs[54]);
    assign layer0_outputs[6953] = 1'b1;
    assign layer0_outputs[6954] = (inputs[88]) & ~(inputs[2]);
    assign layer0_outputs[6955] = (inputs[188]) ^ (inputs[185]);
    assign layer0_outputs[6956] = (inputs[48]) | (inputs[28]);
    assign layer0_outputs[6957] = (inputs[99]) ^ (inputs[214]);
    assign layer0_outputs[6958] = ~(inputs[141]);
    assign layer0_outputs[6959] = ~(inputs[35]);
    assign layer0_outputs[6960] = inputs[167];
    assign layer0_outputs[6961] = (inputs[151]) ^ (inputs[197]);
    assign layer0_outputs[6962] = ~(inputs[176]);
    assign layer0_outputs[6963] = ~(inputs[37]);
    assign layer0_outputs[6964] = ~(inputs[81]);
    assign layer0_outputs[6965] = ~(inputs[22]) | (inputs[160]);
    assign layer0_outputs[6966] = ~(inputs[143]);
    assign layer0_outputs[6967] = inputs[147];
    assign layer0_outputs[6968] = ~((inputs[150]) ^ (inputs[103]));
    assign layer0_outputs[6969] = inputs[121];
    assign layer0_outputs[6970] = ~(inputs[117]);
    assign layer0_outputs[6971] = inputs[116];
    assign layer0_outputs[6972] = ~(inputs[98]);
    assign layer0_outputs[6973] = (inputs[202]) & ~(inputs[78]);
    assign layer0_outputs[6974] = (inputs[168]) & ~(inputs[79]);
    assign layer0_outputs[6975] = ~(inputs[165]) | (inputs[90]);
    assign layer0_outputs[6976] = (inputs[79]) | (inputs[106]);
    assign layer0_outputs[6977] = inputs[52];
    assign layer0_outputs[6978] = ~((inputs[59]) | (inputs[111]));
    assign layer0_outputs[6979] = ~(inputs[215]) | (inputs[67]);
    assign layer0_outputs[6980] = inputs[188];
    assign layer0_outputs[6981] = inputs[106];
    assign layer0_outputs[6982] = ~(inputs[99]);
    assign layer0_outputs[6983] = (inputs[242]) & ~(inputs[13]);
    assign layer0_outputs[6984] = (inputs[213]) & (inputs[113]);
    assign layer0_outputs[6985] = (inputs[129]) | (inputs[203]);
    assign layer0_outputs[6986] = inputs[66];
    assign layer0_outputs[6987] = ~(inputs[6]) | (inputs[128]);
    assign layer0_outputs[6988] = (inputs[155]) & (inputs[108]);
    assign layer0_outputs[6989] = (inputs[114]) | (inputs[70]);
    assign layer0_outputs[6990] = ~(inputs[229]);
    assign layer0_outputs[6991] = ~((inputs[239]) & (inputs[13]));
    assign layer0_outputs[6992] = (inputs[86]) & ~(inputs[78]);
    assign layer0_outputs[6993] = inputs[253];
    assign layer0_outputs[6994] = ~(inputs[196]) | (inputs[124]);
    assign layer0_outputs[6995] = (inputs[90]) & ~(inputs[65]);
    assign layer0_outputs[6996] = inputs[237];
    assign layer0_outputs[6997] = (inputs[32]) | (inputs[210]);
    assign layer0_outputs[6998] = (inputs[176]) | (inputs[94]);
    assign layer0_outputs[6999] = (inputs[114]) | (inputs[225]);
    assign layer0_outputs[7000] = inputs[67];
    assign layer0_outputs[7001] = ~(inputs[109]);
    assign layer0_outputs[7002] = ~((inputs[172]) | (inputs[213]));
    assign layer0_outputs[7003] = ~(inputs[103]) | (inputs[114]);
    assign layer0_outputs[7004] = (inputs[188]) | (inputs[2]);
    assign layer0_outputs[7005] = ~(inputs[19]) | (inputs[144]);
    assign layer0_outputs[7006] = inputs[112];
    assign layer0_outputs[7007] = (inputs[83]) & ~(inputs[220]);
    assign layer0_outputs[7008] = inputs[253];
    assign layer0_outputs[7009] = (inputs[38]) & ~(inputs[206]);
    assign layer0_outputs[7010] = inputs[24];
    assign layer0_outputs[7011] = inputs[253];
    assign layer0_outputs[7012] = inputs[146];
    assign layer0_outputs[7013] = ~(inputs[28]);
    assign layer0_outputs[7014] = ~(inputs[171]);
    assign layer0_outputs[7015] = ~((inputs[84]) | (inputs[102]));
    assign layer0_outputs[7016] = (inputs[129]) & ~(inputs[122]);
    assign layer0_outputs[7017] = 1'b1;
    assign layer0_outputs[7018] = ~((inputs[180]) ^ (inputs[178]));
    assign layer0_outputs[7019] = (inputs[95]) & ~(inputs[4]);
    assign layer0_outputs[7020] = inputs[59];
    assign layer0_outputs[7021] = ~(inputs[121]);
    assign layer0_outputs[7022] = ~(inputs[21]) | (inputs[46]);
    assign layer0_outputs[7023] = ~((inputs[205]) | (inputs[43]));
    assign layer0_outputs[7024] = ~(inputs[3]) | (inputs[249]);
    assign layer0_outputs[7025] = (inputs[63]) | (inputs[124]);
    assign layer0_outputs[7026] = ~((inputs[200]) ^ (inputs[133]));
    assign layer0_outputs[7027] = ~((inputs[108]) | (inputs[0]));
    assign layer0_outputs[7028] = ~(inputs[40]);
    assign layer0_outputs[7029] = (inputs[29]) ^ (inputs[11]);
    assign layer0_outputs[7030] = ~((inputs[32]) | (inputs[214]));
    assign layer0_outputs[7031] = inputs[37];
    assign layer0_outputs[7032] = (inputs[34]) | (inputs[75]);
    assign layer0_outputs[7033] = (inputs[72]) ^ (inputs[26]);
    assign layer0_outputs[7034] = (inputs[189]) | (inputs[201]);
    assign layer0_outputs[7035] = ~((inputs[240]) | (inputs[223]));
    assign layer0_outputs[7036] = ~(inputs[99]);
    assign layer0_outputs[7037] = (inputs[80]) | (inputs[65]);
    assign layer0_outputs[7038] = ~(inputs[183]);
    assign layer0_outputs[7039] = (inputs[186]) | (inputs[112]);
    assign layer0_outputs[7040] = (inputs[127]) & ~(inputs[64]);
    assign layer0_outputs[7041] = ~(inputs[245]);
    assign layer0_outputs[7042] = inputs[113];
    assign layer0_outputs[7043] = (inputs[91]) | (inputs[113]);
    assign layer0_outputs[7044] = 1'b0;
    assign layer0_outputs[7045] = ~(inputs[229]);
    assign layer0_outputs[7046] = inputs[124];
    assign layer0_outputs[7047] = (inputs[24]) ^ (inputs[134]);
    assign layer0_outputs[7048] = ~((inputs[213]) | (inputs[213]));
    assign layer0_outputs[7049] = (inputs[217]) ^ (inputs[91]);
    assign layer0_outputs[7050] = ~((inputs[120]) ^ (inputs[88]));
    assign layer0_outputs[7051] = ~(inputs[89]) | (inputs[81]);
    assign layer0_outputs[7052] = (inputs[247]) | (inputs[229]);
    assign layer0_outputs[7053] = inputs[249];
    assign layer0_outputs[7054] = ~((inputs[34]) | (inputs[23]));
    assign layer0_outputs[7055] = ~(inputs[157]);
    assign layer0_outputs[7056] = inputs[34];
    assign layer0_outputs[7057] = (inputs[216]) ^ (inputs[48]);
    assign layer0_outputs[7058] = ~(inputs[22]) | (inputs[249]);
    assign layer0_outputs[7059] = (inputs[38]) ^ (inputs[7]);
    assign layer0_outputs[7060] = ~((inputs[110]) | (inputs[13]));
    assign layer0_outputs[7061] = (inputs[113]) & ~(inputs[115]);
    assign layer0_outputs[7062] = (inputs[14]) ^ (inputs[49]);
    assign layer0_outputs[7063] = (inputs[163]) ^ (inputs[116]);
    assign layer0_outputs[7064] = ~(inputs[89]);
    assign layer0_outputs[7065] = (inputs[199]) & ~(inputs[184]);
    assign layer0_outputs[7066] = 1'b1;
    assign layer0_outputs[7067] = ~(inputs[162]);
    assign layer0_outputs[7068] = ~((inputs[13]) & (inputs[243]));
    assign layer0_outputs[7069] = ~((inputs[35]) | (inputs[95]));
    assign layer0_outputs[7070] = inputs[106];
    assign layer0_outputs[7071] = inputs[61];
    assign layer0_outputs[7072] = ~((inputs[149]) ^ (inputs[209]));
    assign layer0_outputs[7073] = ~((inputs[119]) | (inputs[87]));
    assign layer0_outputs[7074] = (inputs[23]) & ~(inputs[164]);
    assign layer0_outputs[7075] = inputs[202];
    assign layer0_outputs[7076] = (inputs[70]) & ~(inputs[200]);
    assign layer0_outputs[7077] = ~(inputs[3]) | (inputs[190]);
    assign layer0_outputs[7078] = ~(inputs[8]);
    assign layer0_outputs[7079] = (inputs[155]) | (inputs[116]);
    assign layer0_outputs[7080] = ~(inputs[170]) | (inputs[98]);
    assign layer0_outputs[7081] = ~((inputs[214]) | (inputs[184]));
    assign layer0_outputs[7082] = ~(inputs[171]) | (inputs[13]);
    assign layer0_outputs[7083] = inputs[145];
    assign layer0_outputs[7084] = (inputs[56]) ^ (inputs[231]);
    assign layer0_outputs[7085] = (inputs[191]) | (inputs[158]);
    assign layer0_outputs[7086] = ~((inputs[220]) ^ (inputs[87]));
    assign layer0_outputs[7087] = (inputs[81]) | (inputs[133]);
    assign layer0_outputs[7088] = ~((inputs[26]) & (inputs[164]));
    assign layer0_outputs[7089] = ~(inputs[26]) | (inputs[229]);
    assign layer0_outputs[7090] = ~(inputs[246]) | (inputs[61]);
    assign layer0_outputs[7091] = (inputs[179]) & ~(inputs[107]);
    assign layer0_outputs[7092] = (inputs[86]) | (inputs[235]);
    assign layer0_outputs[7093] = (inputs[138]) | (inputs[237]);
    assign layer0_outputs[7094] = ~(inputs[61]) | (inputs[144]);
    assign layer0_outputs[7095] = ~(inputs[45]);
    assign layer0_outputs[7096] = ~((inputs[157]) | (inputs[96]));
    assign layer0_outputs[7097] = (inputs[114]) ^ (inputs[186]);
    assign layer0_outputs[7098] = (inputs[202]) ^ (inputs[61]);
    assign layer0_outputs[7099] = ~((inputs[198]) | (inputs[32]));
    assign layer0_outputs[7100] = inputs[254];
    assign layer0_outputs[7101] = ~(inputs[228]);
    assign layer0_outputs[7102] = inputs[203];
    assign layer0_outputs[7103] = ~(inputs[168]);
    assign layer0_outputs[7104] = ~(inputs[245]);
    assign layer0_outputs[7105] = ~(inputs[29]);
    assign layer0_outputs[7106] = (inputs[155]) ^ (inputs[202]);
    assign layer0_outputs[7107] = ~(inputs[101]) | (inputs[19]);
    assign layer0_outputs[7108] = ~(inputs[213]);
    assign layer0_outputs[7109] = (inputs[167]) & ~(inputs[113]);
    assign layer0_outputs[7110] = (inputs[233]) & ~(inputs[142]);
    assign layer0_outputs[7111] = (inputs[200]) | (inputs[84]);
    assign layer0_outputs[7112] = ~(inputs[251]);
    assign layer0_outputs[7113] = (inputs[116]) | (inputs[102]);
    assign layer0_outputs[7114] = (inputs[149]) & ~(inputs[190]);
    assign layer0_outputs[7115] = ~((inputs[140]) ^ (inputs[15]));
    assign layer0_outputs[7116] = ~((inputs[119]) ^ (inputs[86]));
    assign layer0_outputs[7117] = (inputs[108]) & ~(inputs[31]);
    assign layer0_outputs[7118] = ~(inputs[150]);
    assign layer0_outputs[7119] = (inputs[93]) & (inputs[194]);
    assign layer0_outputs[7120] = inputs[26];
    assign layer0_outputs[7121] = ~(inputs[161]);
    assign layer0_outputs[7122] = (inputs[243]) | (inputs[109]);
    assign layer0_outputs[7123] = (inputs[168]) & ~(inputs[129]);
    assign layer0_outputs[7124] = inputs[151];
    assign layer0_outputs[7125] = (inputs[153]) | (inputs[245]);
    assign layer0_outputs[7126] = (inputs[212]) & ~(inputs[149]);
    assign layer0_outputs[7127] = (inputs[80]) ^ (inputs[48]);
    assign layer0_outputs[7128] = ~((inputs[160]) ^ (inputs[97]));
    assign layer0_outputs[7129] = (inputs[187]) & ~(inputs[1]);
    assign layer0_outputs[7130] = ~(inputs[90]) | (inputs[201]);
    assign layer0_outputs[7131] = ~(inputs[220]) | (inputs[94]);
    assign layer0_outputs[7132] = ~((inputs[79]) ^ (inputs[92]));
    assign layer0_outputs[7133] = inputs[147];
    assign layer0_outputs[7134] = ~(inputs[127]);
    assign layer0_outputs[7135] = inputs[196];
    assign layer0_outputs[7136] = (inputs[14]) & ~(inputs[134]);
    assign layer0_outputs[7137] = (inputs[202]) & ~(inputs[23]);
    assign layer0_outputs[7138] = inputs[177];
    assign layer0_outputs[7139] = inputs[131];
    assign layer0_outputs[7140] = (inputs[75]) | (inputs[54]);
    assign layer0_outputs[7141] = (inputs[111]) | (inputs[131]);
    assign layer0_outputs[7142] = ~(inputs[13]);
    assign layer0_outputs[7143] = ~(inputs[142]);
    assign layer0_outputs[7144] = (inputs[130]) & (inputs[11]);
    assign layer0_outputs[7145] = (inputs[38]) ^ (inputs[143]);
    assign layer0_outputs[7146] = inputs[195];
    assign layer0_outputs[7147] = ~(inputs[230]);
    assign layer0_outputs[7148] = ~((inputs[146]) | (inputs[204]));
    assign layer0_outputs[7149] = 1'b1;
    assign layer0_outputs[7150] = ~(inputs[130]);
    assign layer0_outputs[7151] = (inputs[157]) & ~(inputs[29]);
    assign layer0_outputs[7152] = (inputs[99]) & ~(inputs[47]);
    assign layer0_outputs[7153] = (inputs[177]) | (inputs[160]);
    assign layer0_outputs[7154] = ~((inputs[111]) | (inputs[150]));
    assign layer0_outputs[7155] = ~(inputs[13]) | (inputs[145]);
    assign layer0_outputs[7156] = (inputs[71]) & (inputs[67]);
    assign layer0_outputs[7157] = ~(inputs[117]);
    assign layer0_outputs[7158] = (inputs[198]) ^ (inputs[230]);
    assign layer0_outputs[7159] = ~((inputs[158]) | (inputs[159]));
    assign layer0_outputs[7160] = (inputs[9]) ^ (inputs[127]);
    assign layer0_outputs[7161] = inputs[167];
    assign layer0_outputs[7162] = (inputs[152]) ^ (inputs[90]);
    assign layer0_outputs[7163] = 1'b0;
    assign layer0_outputs[7164] = (inputs[141]) | (inputs[50]);
    assign layer0_outputs[7165] = inputs[131];
    assign layer0_outputs[7166] = inputs[180];
    assign layer0_outputs[7167] = ~((inputs[140]) ^ (inputs[202]));
    assign layer0_outputs[7168] = ~(inputs[106]);
    assign layer0_outputs[7169] = inputs[186];
    assign layer0_outputs[7170] = ~(inputs[160]) | (inputs[72]);
    assign layer0_outputs[7171] = inputs[42];
    assign layer0_outputs[7172] = (inputs[195]) ^ (inputs[224]);
    assign layer0_outputs[7173] = ~(inputs[70]) | (inputs[33]);
    assign layer0_outputs[7174] = (inputs[218]) ^ (inputs[65]);
    assign layer0_outputs[7175] = inputs[22];
    assign layer0_outputs[7176] = inputs[241];
    assign layer0_outputs[7177] = (inputs[73]) & ~(inputs[224]);
    assign layer0_outputs[7178] = (inputs[164]) & ~(inputs[12]);
    assign layer0_outputs[7179] = ~(inputs[228]);
    assign layer0_outputs[7180] = ~(inputs[175]) | (inputs[128]);
    assign layer0_outputs[7181] = ~(inputs[177]);
    assign layer0_outputs[7182] = (inputs[20]) & ~(inputs[146]);
    assign layer0_outputs[7183] = (inputs[245]) & (inputs[199]);
    assign layer0_outputs[7184] = (inputs[55]) | (inputs[176]);
    assign layer0_outputs[7185] = (inputs[112]) | (inputs[29]);
    assign layer0_outputs[7186] = 1'b1;
    assign layer0_outputs[7187] = (inputs[227]) | (inputs[232]);
    assign layer0_outputs[7188] = ~(inputs[71]);
    assign layer0_outputs[7189] = (inputs[138]) | (inputs[239]);
    assign layer0_outputs[7190] = ~(inputs[174]);
    assign layer0_outputs[7191] = (inputs[103]) | (inputs[220]);
    assign layer0_outputs[7192] = (inputs[210]) | (inputs[8]);
    assign layer0_outputs[7193] = ~((inputs[231]) ^ (inputs[184]));
    assign layer0_outputs[7194] = ~(inputs[91]);
    assign layer0_outputs[7195] = (inputs[90]) | (inputs[110]);
    assign layer0_outputs[7196] = ~((inputs[29]) ^ (inputs[12]));
    assign layer0_outputs[7197] = (inputs[40]) & ~(inputs[160]);
    assign layer0_outputs[7198] = ~(inputs[133]);
    assign layer0_outputs[7199] = (inputs[182]) | (inputs[131]);
    assign layer0_outputs[7200] = inputs[116];
    assign layer0_outputs[7201] = (inputs[106]) & ~(inputs[94]);
    assign layer0_outputs[7202] = (inputs[164]) | (inputs[238]);
    assign layer0_outputs[7203] = ~(inputs[228]) | (inputs[125]);
    assign layer0_outputs[7204] = (inputs[249]) & ~(inputs[170]);
    assign layer0_outputs[7205] = (inputs[154]) ^ (inputs[123]);
    assign layer0_outputs[7206] = (inputs[234]) ^ (inputs[96]);
    assign layer0_outputs[7207] = (inputs[243]) & ~(inputs[144]);
    assign layer0_outputs[7208] = ~(inputs[246]) | (inputs[76]);
    assign layer0_outputs[7209] = inputs[23];
    assign layer0_outputs[7210] = ~((inputs[31]) | (inputs[170]));
    assign layer0_outputs[7211] = ~(inputs[28]) | (inputs[252]);
    assign layer0_outputs[7212] = ~(inputs[25]);
    assign layer0_outputs[7213] = ~((inputs[48]) | (inputs[77]));
    assign layer0_outputs[7214] = inputs[122];
    assign layer0_outputs[7215] = (inputs[1]) ^ (inputs[140]);
    assign layer0_outputs[7216] = (inputs[93]) & ~(inputs[81]);
    assign layer0_outputs[7217] = ~(inputs[5]) | (inputs[30]);
    assign layer0_outputs[7218] = (inputs[118]) ^ (inputs[87]);
    assign layer0_outputs[7219] = ~((inputs[221]) | (inputs[216]));
    assign layer0_outputs[7220] = inputs[143];
    assign layer0_outputs[7221] = ~(inputs[74]);
    assign layer0_outputs[7222] = (inputs[135]) & ~(inputs[229]);
    assign layer0_outputs[7223] = ~((inputs[121]) ^ (inputs[169]));
    assign layer0_outputs[7224] = ~((inputs[133]) & (inputs[153]));
    assign layer0_outputs[7225] = ~(inputs[145]);
    assign layer0_outputs[7226] = ~(inputs[146]);
    assign layer0_outputs[7227] = ~((inputs[97]) ^ (inputs[85]));
    assign layer0_outputs[7228] = ~((inputs[206]) & (inputs[2]));
    assign layer0_outputs[7229] = ~((inputs[171]) | (inputs[219]));
    assign layer0_outputs[7230] = ~((inputs[83]) | (inputs[37]));
    assign layer0_outputs[7231] = ~(inputs[230]);
    assign layer0_outputs[7232] = 1'b0;
    assign layer0_outputs[7233] = inputs[178];
    assign layer0_outputs[7234] = ~(inputs[209]) | (inputs[67]);
    assign layer0_outputs[7235] = inputs[47];
    assign layer0_outputs[7236] = ~(inputs[206]) | (inputs[45]);
    assign layer0_outputs[7237] = inputs[91];
    assign layer0_outputs[7238] = ~((inputs[165]) ^ (inputs[192]));
    assign layer0_outputs[7239] = (inputs[131]) ^ (inputs[134]);
    assign layer0_outputs[7240] = (inputs[55]) & ~(inputs[31]);
    assign layer0_outputs[7241] = inputs[95];
    assign layer0_outputs[7242] = ~((inputs[37]) ^ (inputs[21]));
    assign layer0_outputs[7243] = ~(inputs[66]) | (inputs[33]);
    assign layer0_outputs[7244] = ~(inputs[47]) | (inputs[147]);
    assign layer0_outputs[7245] = ~((inputs[133]) | (inputs[132]));
    assign layer0_outputs[7246] = ~((inputs[125]) | (inputs[253]));
    assign layer0_outputs[7247] = ~(inputs[95]) | (inputs[237]);
    assign layer0_outputs[7248] = ~(inputs[123]);
    assign layer0_outputs[7249] = ~(inputs[68]) | (inputs[63]);
    assign layer0_outputs[7250] = ~((inputs[73]) ^ (inputs[91]));
    assign layer0_outputs[7251] = 1'b1;
    assign layer0_outputs[7252] = inputs[128];
    assign layer0_outputs[7253] = (inputs[34]) ^ (inputs[56]);
    assign layer0_outputs[7254] = (inputs[63]) & ~(inputs[14]);
    assign layer0_outputs[7255] = ~(inputs[41]) | (inputs[85]);
    assign layer0_outputs[7256] = (inputs[167]) & (inputs[151]);
    assign layer0_outputs[7257] = (inputs[164]) & (inputs[64]);
    assign layer0_outputs[7258] = ~(inputs[198]);
    assign layer0_outputs[7259] = ~(inputs[74]);
    assign layer0_outputs[7260] = (inputs[180]) ^ (inputs[193]);
    assign layer0_outputs[7261] = ~(inputs[134]) | (inputs[72]);
    assign layer0_outputs[7262] = (inputs[3]) | (inputs[46]);
    assign layer0_outputs[7263] = ~(inputs[130]);
    assign layer0_outputs[7264] = inputs[251];
    assign layer0_outputs[7265] = (inputs[204]) & ~(inputs[16]);
    assign layer0_outputs[7266] = (inputs[217]) ^ (inputs[150]);
    assign layer0_outputs[7267] = inputs[166];
    assign layer0_outputs[7268] = ~((inputs[162]) | (inputs[96]));
    assign layer0_outputs[7269] = (inputs[196]) | (inputs[85]);
    assign layer0_outputs[7270] = ~((inputs[172]) | (inputs[157]));
    assign layer0_outputs[7271] = (inputs[8]) & ~(inputs[220]);
    assign layer0_outputs[7272] = ~(inputs[207]);
    assign layer0_outputs[7273] = (inputs[42]) ^ (inputs[205]);
    assign layer0_outputs[7274] = ~(inputs[142]);
    assign layer0_outputs[7275] = ~((inputs[115]) ^ (inputs[44]));
    assign layer0_outputs[7276] = ~((inputs[141]) | (inputs[132]));
    assign layer0_outputs[7277] = ~(inputs[109]);
    assign layer0_outputs[7278] = inputs[52];
    assign layer0_outputs[7279] = (inputs[100]) & ~(inputs[41]);
    assign layer0_outputs[7280] = (inputs[75]) | (inputs[136]);
    assign layer0_outputs[7281] = (inputs[80]) | (inputs[148]);
    assign layer0_outputs[7282] = (inputs[250]) | (inputs[153]);
    assign layer0_outputs[7283] = ~((inputs[163]) & (inputs[126]));
    assign layer0_outputs[7284] = 1'b0;
    assign layer0_outputs[7285] = ~((inputs[97]) ^ (inputs[81]));
    assign layer0_outputs[7286] = inputs[64];
    assign layer0_outputs[7287] = ~((inputs[37]) | (inputs[95]));
    assign layer0_outputs[7288] = ~((inputs[143]) ^ (inputs[248]));
    assign layer0_outputs[7289] = ~(inputs[181]) | (inputs[188]);
    assign layer0_outputs[7290] = ~(inputs[89]) | (inputs[68]);
    assign layer0_outputs[7291] = ~(inputs[151]);
    assign layer0_outputs[7292] = 1'b0;
    assign layer0_outputs[7293] = ~((inputs[197]) | (inputs[123]));
    assign layer0_outputs[7294] = ~((inputs[209]) | (inputs[182]));
    assign layer0_outputs[7295] = (inputs[171]) ^ (inputs[37]);
    assign layer0_outputs[7296] = (inputs[49]) ^ (inputs[220]);
    assign layer0_outputs[7297] = (inputs[155]) & ~(inputs[197]);
    assign layer0_outputs[7298] = ~(inputs[192]);
    assign layer0_outputs[7299] = ~(inputs[247]) | (inputs[95]);
    assign layer0_outputs[7300] = inputs[65];
    assign layer0_outputs[7301] = ~((inputs[188]) ^ (inputs[246]));
    assign layer0_outputs[7302] = ~((inputs[181]) | (inputs[251]));
    assign layer0_outputs[7303] = ~(inputs[37]) | (inputs[176]);
    assign layer0_outputs[7304] = ~(inputs[130]) | (inputs[71]);
    assign layer0_outputs[7305] = 1'b0;
    assign layer0_outputs[7306] = inputs[54];
    assign layer0_outputs[7307] = ~(inputs[57]);
    assign layer0_outputs[7308] = ~(inputs[69]);
    assign layer0_outputs[7309] = ~((inputs[25]) | (inputs[18]));
    assign layer0_outputs[7310] = inputs[229];
    assign layer0_outputs[7311] = (inputs[95]) | (inputs[33]);
    assign layer0_outputs[7312] = ~((inputs[242]) | (inputs[138]));
    assign layer0_outputs[7313] = ~((inputs[215]) ^ (inputs[207]));
    assign layer0_outputs[7314] = ~(inputs[148]);
    assign layer0_outputs[7315] = (inputs[39]) & ~(inputs[217]);
    assign layer0_outputs[7316] = inputs[190];
    assign layer0_outputs[7317] = 1'b0;
    assign layer0_outputs[7318] = (inputs[148]) & ~(inputs[206]);
    assign layer0_outputs[7319] = (inputs[165]) | (inputs[188]);
    assign layer0_outputs[7320] = ~((inputs[202]) ^ (inputs[144]));
    assign layer0_outputs[7321] = ~(inputs[195]);
    assign layer0_outputs[7322] = ~(inputs[210]);
    assign layer0_outputs[7323] = inputs[53];
    assign layer0_outputs[7324] = inputs[74];
    assign layer0_outputs[7325] = inputs[13];
    assign layer0_outputs[7326] = inputs[99];
    assign layer0_outputs[7327] = ~(inputs[137]) | (inputs[111]);
    assign layer0_outputs[7328] = 1'b0;
    assign layer0_outputs[7329] = inputs[130];
    assign layer0_outputs[7330] = ~(inputs[45]) | (inputs[18]);
    assign layer0_outputs[7331] = ~(inputs[229]);
    assign layer0_outputs[7332] = (inputs[53]) & ~(inputs[126]);
    assign layer0_outputs[7333] = (inputs[196]) ^ (inputs[243]);
    assign layer0_outputs[7334] = ~((inputs[135]) | (inputs[183]));
    assign layer0_outputs[7335] = ~((inputs[8]) ^ (inputs[39]));
    assign layer0_outputs[7336] = ~(inputs[177]);
    assign layer0_outputs[7337] = (inputs[157]) | (inputs[10]);
    assign layer0_outputs[7338] = (inputs[140]) & (inputs[114]);
    assign layer0_outputs[7339] = ~((inputs[74]) | (inputs[73]));
    assign layer0_outputs[7340] = ~(inputs[98]);
    assign layer0_outputs[7341] = (inputs[187]) ^ (inputs[195]);
    assign layer0_outputs[7342] = (inputs[89]) ^ (inputs[97]);
    assign layer0_outputs[7343] = (inputs[24]) & ~(inputs[250]);
    assign layer0_outputs[7344] = ~(inputs[24]) | (inputs[242]);
    assign layer0_outputs[7345] = ~(inputs[46]) | (inputs[187]);
    assign layer0_outputs[7346] = (inputs[53]) ^ (inputs[185]);
    assign layer0_outputs[7347] = (inputs[232]) ^ (inputs[160]);
    assign layer0_outputs[7348] = (inputs[95]) | (inputs[170]);
    assign layer0_outputs[7349] = (inputs[9]) ^ (inputs[217]);
    assign layer0_outputs[7350] = ~(inputs[119]);
    assign layer0_outputs[7351] = (inputs[140]) & (inputs[136]);
    assign layer0_outputs[7352] = (inputs[49]) ^ (inputs[233]);
    assign layer0_outputs[7353] = 1'b0;
    assign layer0_outputs[7354] = (inputs[34]) ^ (inputs[173]);
    assign layer0_outputs[7355] = ~((inputs[65]) | (inputs[165]));
    assign layer0_outputs[7356] = inputs[167];
    assign layer0_outputs[7357] = ~((inputs[104]) | (inputs[238]));
    assign layer0_outputs[7358] = ~((inputs[193]) | (inputs[211]));
    assign layer0_outputs[7359] = inputs[62];
    assign layer0_outputs[7360] = (inputs[182]) | (inputs[231]);
    assign layer0_outputs[7361] = inputs[73];
    assign layer0_outputs[7362] = ~(inputs[131]);
    assign layer0_outputs[7363] = (inputs[105]) & ~(inputs[143]);
    assign layer0_outputs[7364] = ~(inputs[95]);
    assign layer0_outputs[7365] = ~((inputs[135]) | (inputs[75]));
    assign layer0_outputs[7366] = inputs[214];
    assign layer0_outputs[7367] = (inputs[126]) | (inputs[201]);
    assign layer0_outputs[7368] = ~(inputs[0]) | (inputs[179]);
    assign layer0_outputs[7369] = (inputs[119]) & ~(inputs[159]);
    assign layer0_outputs[7370] = ~(inputs[3]) | (inputs[33]);
    assign layer0_outputs[7371] = inputs[53];
    assign layer0_outputs[7372] = ~((inputs[204]) ^ (inputs[197]));
    assign layer0_outputs[7373] = ~(inputs[17]) | (inputs[128]);
    assign layer0_outputs[7374] = ~(inputs[59]) | (inputs[178]);
    assign layer0_outputs[7375] = (inputs[118]) & ~(inputs[149]);
    assign layer0_outputs[7376] = ~(inputs[199]) | (inputs[53]);
    assign layer0_outputs[7377] = ~(inputs[84]);
    assign layer0_outputs[7378] = (inputs[19]) | (inputs[188]);
    assign layer0_outputs[7379] = ~((inputs[141]) & (inputs[158]));
    assign layer0_outputs[7380] = ~(inputs[179]) | (inputs[35]);
    assign layer0_outputs[7381] = (inputs[112]) | (inputs[34]);
    assign layer0_outputs[7382] = (inputs[213]) | (inputs[249]);
    assign layer0_outputs[7383] = (inputs[114]) & ~(inputs[221]);
    assign layer0_outputs[7384] = ~((inputs[234]) & (inputs[140]));
    assign layer0_outputs[7385] = (inputs[158]) & ~(inputs[112]);
    assign layer0_outputs[7386] = ~(inputs[68]);
    assign layer0_outputs[7387] = ~((inputs[125]) | (inputs[47]));
    assign layer0_outputs[7388] = ~((inputs[62]) | (inputs[195]));
    assign layer0_outputs[7389] = (inputs[69]) & (inputs[186]);
    assign layer0_outputs[7390] = inputs[167];
    assign layer0_outputs[7391] = inputs[98];
    assign layer0_outputs[7392] = ~((inputs[234]) ^ (inputs[107]));
    assign layer0_outputs[7393] = inputs[100];
    assign layer0_outputs[7394] = inputs[183];
    assign layer0_outputs[7395] = 1'b1;
    assign layer0_outputs[7396] = (inputs[69]) & ~(inputs[224]);
    assign layer0_outputs[7397] = inputs[168];
    assign layer0_outputs[7398] = ~((inputs[14]) ^ (inputs[56]));
    assign layer0_outputs[7399] = (inputs[157]) | (inputs[9]);
    assign layer0_outputs[7400] = ~(inputs[162]) | (inputs[64]);
    assign layer0_outputs[7401] = ~((inputs[245]) | (inputs[98]));
    assign layer0_outputs[7402] = ~(inputs[75]);
    assign layer0_outputs[7403] = (inputs[185]) ^ (inputs[218]);
    assign layer0_outputs[7404] = inputs[167];
    assign layer0_outputs[7405] = ~((inputs[96]) | (inputs[165]));
    assign layer0_outputs[7406] = (inputs[202]) | (inputs[18]);
    assign layer0_outputs[7407] = (inputs[63]) | (inputs[233]);
    assign layer0_outputs[7408] = ~((inputs[222]) ^ (inputs[180]));
    assign layer0_outputs[7409] = (inputs[77]) | (inputs[3]);
    assign layer0_outputs[7410] = ~((inputs[188]) ^ (inputs[221]));
    assign layer0_outputs[7411] = ~((inputs[188]) ^ (inputs[129]));
    assign layer0_outputs[7412] = ~(inputs[54]);
    assign layer0_outputs[7413] = (inputs[252]) & (inputs[252]);
    assign layer0_outputs[7414] = 1'b1;
    assign layer0_outputs[7415] = (inputs[246]) | (inputs[229]);
    assign layer0_outputs[7416] = ~(inputs[219]);
    assign layer0_outputs[7417] = inputs[105];
    assign layer0_outputs[7418] = ~((inputs[182]) | (inputs[226]));
    assign layer0_outputs[7419] = (inputs[96]) | (inputs[238]);
    assign layer0_outputs[7420] = (inputs[224]) & ~(inputs[30]);
    assign layer0_outputs[7421] = ~(inputs[163]);
    assign layer0_outputs[7422] = ~(inputs[22]);
    assign layer0_outputs[7423] = ~(inputs[94]) | (inputs[153]);
    assign layer0_outputs[7424] = ~((inputs[178]) | (inputs[24]));
    assign layer0_outputs[7425] = ~((inputs[38]) & (inputs[102]));
    assign layer0_outputs[7426] = (inputs[231]) | (inputs[246]);
    assign layer0_outputs[7427] = ~(inputs[100]);
    assign layer0_outputs[7428] = ~((inputs[5]) ^ (inputs[70]));
    assign layer0_outputs[7429] = (inputs[11]) & (inputs[131]);
    assign layer0_outputs[7430] = (inputs[12]) & ~(inputs[79]);
    assign layer0_outputs[7431] = (inputs[7]) | (inputs[204]);
    assign layer0_outputs[7432] = inputs[183];
    assign layer0_outputs[7433] = ~((inputs[216]) | (inputs[226]));
    assign layer0_outputs[7434] = inputs[226];
    assign layer0_outputs[7435] = inputs[121];
    assign layer0_outputs[7436] = (inputs[74]) & ~(inputs[201]);
    assign layer0_outputs[7437] = (inputs[163]) & ~(inputs[222]);
    assign layer0_outputs[7438] = inputs[151];
    assign layer0_outputs[7439] = 1'b0;
    assign layer0_outputs[7440] = ~(inputs[120]);
    assign layer0_outputs[7441] = ~((inputs[102]) ^ (inputs[169]));
    assign layer0_outputs[7442] = inputs[169];
    assign layer0_outputs[7443] = ~(inputs[210]) | (inputs[139]);
    assign layer0_outputs[7444] = ~(inputs[130]);
    assign layer0_outputs[7445] = 1'b1;
    assign layer0_outputs[7446] = ~((inputs[45]) | (inputs[108]));
    assign layer0_outputs[7447] = inputs[179];
    assign layer0_outputs[7448] = ~(inputs[247]);
    assign layer0_outputs[7449] = inputs[140];
    assign layer0_outputs[7450] = ~(inputs[49]);
    assign layer0_outputs[7451] = (inputs[228]) & ~(inputs[86]);
    assign layer0_outputs[7452] = ~((inputs[84]) ^ (inputs[38]));
    assign layer0_outputs[7453] = ~((inputs[223]) | (inputs[206]));
    assign layer0_outputs[7454] = inputs[10];
    assign layer0_outputs[7455] = ~(inputs[91]) | (inputs[159]);
    assign layer0_outputs[7456] = ~(inputs[130]) | (inputs[237]);
    assign layer0_outputs[7457] = inputs[134];
    assign layer0_outputs[7458] = ~(inputs[194]) | (inputs[122]);
    assign layer0_outputs[7459] = inputs[73];
    assign layer0_outputs[7460] = (inputs[113]) ^ (inputs[36]);
    assign layer0_outputs[7461] = (inputs[219]) | (inputs[162]);
    assign layer0_outputs[7462] = ~((inputs[78]) & (inputs[43]));
    assign layer0_outputs[7463] = 1'b0;
    assign layer0_outputs[7464] = ~(inputs[38]);
    assign layer0_outputs[7465] = ~(inputs[53]) | (inputs[13]);
    assign layer0_outputs[7466] = inputs[175];
    assign layer0_outputs[7467] = ~((inputs[71]) ^ (inputs[45]));
    assign layer0_outputs[7468] = (inputs[92]) | (inputs[246]);
    assign layer0_outputs[7469] = ~(inputs[59]) | (inputs[253]);
    assign layer0_outputs[7470] = inputs[112];
    assign layer0_outputs[7471] = (inputs[207]) | (inputs[62]);
    assign layer0_outputs[7472] = (inputs[17]) & (inputs[144]);
    assign layer0_outputs[7473] = ~((inputs[254]) & (inputs[168]));
    assign layer0_outputs[7474] = ~(inputs[222]);
    assign layer0_outputs[7475] = ~((inputs[216]) | (inputs[228]));
    assign layer0_outputs[7476] = inputs[19];
    assign layer0_outputs[7477] = ~(inputs[117]);
    assign layer0_outputs[7478] = ~(inputs[92]);
    assign layer0_outputs[7479] = ~(inputs[53]);
    assign layer0_outputs[7480] = ~(inputs[214]) | (inputs[52]);
    assign layer0_outputs[7481] = (inputs[141]) | (inputs[219]);
    assign layer0_outputs[7482] = inputs[26];
    assign layer0_outputs[7483] = ~((inputs[211]) ^ (inputs[110]));
    assign layer0_outputs[7484] = (inputs[222]) ^ (inputs[251]);
    assign layer0_outputs[7485] = (inputs[45]) & ~(inputs[240]);
    assign layer0_outputs[7486] = ~((inputs[243]) ^ (inputs[197]));
    assign layer0_outputs[7487] = (inputs[97]) | (inputs[109]);
    assign layer0_outputs[7488] = (inputs[212]) ^ (inputs[180]);
    assign layer0_outputs[7489] = ~((inputs[240]) | (inputs[30]));
    assign layer0_outputs[7490] = inputs[134];
    assign layer0_outputs[7491] = ~((inputs[89]) | (inputs[120]));
    assign layer0_outputs[7492] = ~((inputs[136]) ^ (inputs[26]));
    assign layer0_outputs[7493] = ~(inputs[158]);
    assign layer0_outputs[7494] = (inputs[27]) & ~(inputs[209]);
    assign layer0_outputs[7495] = inputs[92];
    assign layer0_outputs[7496] = (inputs[213]) | (inputs[211]);
    assign layer0_outputs[7497] = ~(inputs[175]);
    assign layer0_outputs[7498] = (inputs[114]) | (inputs[99]);
    assign layer0_outputs[7499] = ~(inputs[159]);
    assign layer0_outputs[7500] = inputs[80];
    assign layer0_outputs[7501] = (inputs[154]) & ~(inputs[78]);
    assign layer0_outputs[7502] = ~((inputs[243]) | (inputs[150]));
    assign layer0_outputs[7503] = ~(inputs[232]);
    assign layer0_outputs[7504] = 1'b0;
    assign layer0_outputs[7505] = ~((inputs[105]) ^ (inputs[203]));
    assign layer0_outputs[7506] = (inputs[128]) | (inputs[76]);
    assign layer0_outputs[7507] = ~((inputs[189]) | (inputs[29]));
    assign layer0_outputs[7508] = inputs[77];
    assign layer0_outputs[7509] = 1'b0;
    assign layer0_outputs[7510] = (inputs[80]) | (inputs[82]);
    assign layer0_outputs[7511] = (inputs[116]) | (inputs[149]);
    assign layer0_outputs[7512] = (inputs[9]) & ~(inputs[226]);
    assign layer0_outputs[7513] = ~((inputs[252]) | (inputs[56]));
    assign layer0_outputs[7514] = ~(inputs[120]);
    assign layer0_outputs[7515] = (inputs[132]) & ~(inputs[32]);
    assign layer0_outputs[7516] = ~(inputs[40]) | (inputs[153]);
    assign layer0_outputs[7517] = (inputs[191]) | (inputs[140]);
    assign layer0_outputs[7518] = ~(inputs[9]);
    assign layer0_outputs[7519] = (inputs[228]) & (inputs[116]);
    assign layer0_outputs[7520] = (inputs[180]) | (inputs[66]);
    assign layer0_outputs[7521] = ~((inputs[86]) | (inputs[154]));
    assign layer0_outputs[7522] = (inputs[87]) & ~(inputs[188]);
    assign layer0_outputs[7523] = ~(inputs[45]) | (inputs[191]);
    assign layer0_outputs[7524] = ~((inputs[93]) ^ (inputs[35]));
    assign layer0_outputs[7525] = ~(inputs[161]);
    assign layer0_outputs[7526] = (inputs[211]) & (inputs[45]);
    assign layer0_outputs[7527] = inputs[122];
    assign layer0_outputs[7528] = ~((inputs[97]) | (inputs[92]));
    assign layer0_outputs[7529] = inputs[120];
    assign layer0_outputs[7530] = inputs[162];
    assign layer0_outputs[7531] = ~((inputs[250]) | (inputs[134]));
    assign layer0_outputs[7532] = ~(inputs[104]);
    assign layer0_outputs[7533] = ~((inputs[130]) ^ (inputs[255]));
    assign layer0_outputs[7534] = (inputs[246]) & (inputs[107]);
    assign layer0_outputs[7535] = (inputs[236]) & ~(inputs[50]);
    assign layer0_outputs[7536] = ~(inputs[204]);
    assign layer0_outputs[7537] = ~(inputs[121]) | (inputs[244]);
    assign layer0_outputs[7538] = inputs[130];
    assign layer0_outputs[7539] = (inputs[177]) & ~(inputs[139]);
    assign layer0_outputs[7540] = ~((inputs[172]) & (inputs[196]));
    assign layer0_outputs[7541] = inputs[66];
    assign layer0_outputs[7542] = ~(inputs[167]);
    assign layer0_outputs[7543] = ~(inputs[225]);
    assign layer0_outputs[7544] = inputs[89];
    assign layer0_outputs[7545] = ~(inputs[51]) | (inputs[143]);
    assign layer0_outputs[7546] = ~(inputs[89]);
    assign layer0_outputs[7547] = inputs[211];
    assign layer0_outputs[7548] = ~(inputs[70]);
    assign layer0_outputs[7549] = ~(inputs[125]);
    assign layer0_outputs[7550] = ~(inputs[94]);
    assign layer0_outputs[7551] = inputs[57];
    assign layer0_outputs[7552] = (inputs[219]) & ~(inputs[151]);
    assign layer0_outputs[7553] = inputs[161];
    assign layer0_outputs[7554] = (inputs[21]) ^ (inputs[231]);
    assign layer0_outputs[7555] = ~(inputs[185]) | (inputs[31]);
    assign layer0_outputs[7556] = ~((inputs[217]) | (inputs[184]));
    assign layer0_outputs[7557] = (inputs[72]) & ~(inputs[50]);
    assign layer0_outputs[7558] = ~(inputs[210]);
    assign layer0_outputs[7559] = ~((inputs[143]) | (inputs[224]));
    assign layer0_outputs[7560] = (inputs[126]) | (inputs[131]);
    assign layer0_outputs[7561] = ~(inputs[110]);
    assign layer0_outputs[7562] = ~((inputs[209]) ^ (inputs[96]));
    assign layer0_outputs[7563] = ~((inputs[71]) | (inputs[93]));
    assign layer0_outputs[7564] = 1'b0;
    assign layer0_outputs[7565] = inputs[69];
    assign layer0_outputs[7566] = (inputs[75]) & ~(inputs[158]);
    assign layer0_outputs[7567] = inputs[24];
    assign layer0_outputs[7568] = (inputs[117]) & ~(inputs[57]);
    assign layer0_outputs[7569] = inputs[8];
    assign layer0_outputs[7570] = ~((inputs[44]) ^ (inputs[90]));
    assign layer0_outputs[7571] = ~((inputs[47]) | (inputs[106]));
    assign layer0_outputs[7572] = ~(inputs[100]);
    assign layer0_outputs[7573] = (inputs[227]) ^ (inputs[108]);
    assign layer0_outputs[7574] = ~((inputs[221]) | (inputs[182]));
    assign layer0_outputs[7575] = (inputs[1]) ^ (inputs[183]);
    assign layer0_outputs[7576] = ~(inputs[203]);
    assign layer0_outputs[7577] = inputs[225];
    assign layer0_outputs[7578] = (inputs[227]) | (inputs[71]);
    assign layer0_outputs[7579] = ~((inputs[138]) ^ (inputs[77]));
    assign layer0_outputs[7580] = inputs[210];
    assign layer0_outputs[7581] = (inputs[172]) & (inputs[228]);
    assign layer0_outputs[7582] = 1'b0;
    assign layer0_outputs[7583] = ~((inputs[180]) | (inputs[68]));
    assign layer0_outputs[7584] = (inputs[153]) & ~(inputs[77]);
    assign layer0_outputs[7585] = inputs[231];
    assign layer0_outputs[7586] = inputs[62];
    assign layer0_outputs[7587] = (inputs[61]) | (inputs[20]);
    assign layer0_outputs[7588] = (inputs[111]) ^ (inputs[123]);
    assign layer0_outputs[7589] = ~((inputs[216]) & (inputs[72]));
    assign layer0_outputs[7590] = ~(inputs[231]) | (inputs[237]);
    assign layer0_outputs[7591] = ~(inputs[171]) | (inputs[2]);
    assign layer0_outputs[7592] = (inputs[221]) ^ (inputs[128]);
    assign layer0_outputs[7593] = (inputs[194]) | (inputs[85]);
    assign layer0_outputs[7594] = (inputs[0]) & ~(inputs[55]);
    assign layer0_outputs[7595] = ~((inputs[90]) ^ (inputs[249]));
    assign layer0_outputs[7596] = (inputs[82]) | (inputs[115]);
    assign layer0_outputs[7597] = (inputs[187]) & ~(inputs[149]);
    assign layer0_outputs[7598] = ~(inputs[41]);
    assign layer0_outputs[7599] = (inputs[15]) | (inputs[12]);
    assign layer0_outputs[7600] = (inputs[150]) | (inputs[41]);
    assign layer0_outputs[7601] = (inputs[95]) | (inputs[76]);
    assign layer0_outputs[7602] = ~(inputs[13]);
    assign layer0_outputs[7603] = (inputs[247]) & ~(inputs[69]);
    assign layer0_outputs[7604] = inputs[162];
    assign layer0_outputs[7605] = ~(inputs[29]) | (inputs[43]);
    assign layer0_outputs[7606] = inputs[77];
    assign layer0_outputs[7607] = (inputs[37]) & ~(inputs[83]);
    assign layer0_outputs[7608] = inputs[62];
    assign layer0_outputs[7609] = ~(inputs[136]) | (inputs[238]);
    assign layer0_outputs[7610] = ~(inputs[156]);
    assign layer0_outputs[7611] = inputs[165];
    assign layer0_outputs[7612] = ~(inputs[102]);
    assign layer0_outputs[7613] = ~((inputs[216]) ^ (inputs[232]));
    assign layer0_outputs[7614] = ~((inputs[202]) & (inputs[77]));
    assign layer0_outputs[7615] = (inputs[136]) & ~(inputs[250]);
    assign layer0_outputs[7616] = ~((inputs[123]) | (inputs[51]));
    assign layer0_outputs[7617] = ~(inputs[176]);
    assign layer0_outputs[7618] = inputs[120];
    assign layer0_outputs[7619] = ~((inputs[199]) | (inputs[179]));
    assign layer0_outputs[7620] = inputs[180];
    assign layer0_outputs[7621] = ~(inputs[137]) | (inputs[189]);
    assign layer0_outputs[7622] = ~((inputs[20]) | (inputs[68]));
    assign layer0_outputs[7623] = ~((inputs[45]) ^ (inputs[11]));
    assign layer0_outputs[7624] = ~((inputs[163]) ^ (inputs[137]));
    assign layer0_outputs[7625] = ~((inputs[182]) & (inputs[198]));
    assign layer0_outputs[7626] = ~((inputs[8]) | (inputs[47]));
    assign layer0_outputs[7627] = (inputs[242]) ^ (inputs[215]);
    assign layer0_outputs[7628] = (inputs[4]) ^ (inputs[114]);
    assign layer0_outputs[7629] = ~((inputs[11]) | (inputs[83]));
    assign layer0_outputs[7630] = 1'b1;
    assign layer0_outputs[7631] = (inputs[185]) ^ (inputs[234]);
    assign layer0_outputs[7632] = (inputs[156]) & ~(inputs[255]);
    assign layer0_outputs[7633] = ~(inputs[113]) | (inputs[223]);
    assign layer0_outputs[7634] = ~(inputs[168]) | (inputs[158]);
    assign layer0_outputs[7635] = ~((inputs[45]) | (inputs[7]));
    assign layer0_outputs[7636] = inputs[113];
    assign layer0_outputs[7637] = (inputs[43]) ^ (inputs[46]);
    assign layer0_outputs[7638] = inputs[229];
    assign layer0_outputs[7639] = inputs[33];
    assign layer0_outputs[7640] = inputs[216];
    assign layer0_outputs[7641] = (inputs[45]) ^ (inputs[125]);
    assign layer0_outputs[7642] = (inputs[154]) ^ (inputs[158]);
    assign layer0_outputs[7643] = ~((inputs[154]) ^ (inputs[72]));
    assign layer0_outputs[7644] = (inputs[32]) | (inputs[164]);
    assign layer0_outputs[7645] = inputs[14];
    assign layer0_outputs[7646] = (inputs[220]) | (inputs[197]);
    assign layer0_outputs[7647] = (inputs[189]) | (inputs[2]);
    assign layer0_outputs[7648] = ~(inputs[34]);
    assign layer0_outputs[7649] = ~((inputs[82]) | (inputs[147]));
    assign layer0_outputs[7650] = (inputs[35]) & (inputs[142]);
    assign layer0_outputs[7651] = ~((inputs[208]) | (inputs[223]));
    assign layer0_outputs[7652] = (inputs[21]) | (inputs[219]);
    assign layer0_outputs[7653] = inputs[168];
    assign layer0_outputs[7654] = (inputs[69]) & ~(inputs[243]);
    assign layer0_outputs[7655] = inputs[147];
    assign layer0_outputs[7656] = inputs[162];
    assign layer0_outputs[7657] = ~((inputs[181]) | (inputs[141]));
    assign layer0_outputs[7658] = (inputs[75]) | (inputs[222]);
    assign layer0_outputs[7659] = ~((inputs[23]) & (inputs[134]));
    assign layer0_outputs[7660] = inputs[211];
    assign layer0_outputs[7661] = ~(inputs[25]);
    assign layer0_outputs[7662] = ~((inputs[91]) ^ (inputs[19]));
    assign layer0_outputs[7663] = ~((inputs[220]) ^ (inputs[253]));
    assign layer0_outputs[7664] = ~(inputs[126]);
    assign layer0_outputs[7665] = ~((inputs[160]) ^ (inputs[86]));
    assign layer0_outputs[7666] = inputs[212];
    assign layer0_outputs[7667] = ~(inputs[151]);
    assign layer0_outputs[7668] = inputs[48];
    assign layer0_outputs[7669] = inputs[165];
    assign layer0_outputs[7670] = ~(inputs[186]) | (inputs[246]);
    assign layer0_outputs[7671] = (inputs[42]) & ~(inputs[224]);
    assign layer0_outputs[7672] = (inputs[132]) | (inputs[114]);
    assign layer0_outputs[7673] = (inputs[77]) | (inputs[108]);
    assign layer0_outputs[7674] = (inputs[24]) & ~(inputs[5]);
    assign layer0_outputs[7675] = inputs[202];
    assign layer0_outputs[7676] = (inputs[60]) & ~(inputs[112]);
    assign layer0_outputs[7677] = 1'b1;
    assign layer0_outputs[7678] = ~((inputs[193]) ^ (inputs[238]));
    assign layer0_outputs[7679] = (inputs[202]) | (inputs[159]);
    assign layer0_outputs[7680] = (inputs[82]) | (inputs[240]);
    assign layer0_outputs[7681] = ~((inputs[241]) | (inputs[247]));
    assign layer0_outputs[7682] = inputs[24];
    assign layer0_outputs[7683] = ~(inputs[186]) | (inputs[16]);
    assign layer0_outputs[7684] = inputs[7];
    assign layer0_outputs[7685] = (inputs[180]) | (inputs[168]);
    assign layer0_outputs[7686] = (inputs[225]) | (inputs[145]);
    assign layer0_outputs[7687] = ~((inputs[206]) | (inputs[50]));
    assign layer0_outputs[7688] = (inputs[42]) ^ (inputs[10]);
    assign layer0_outputs[7689] = (inputs[172]) | (inputs[187]);
    assign layer0_outputs[7690] = inputs[225];
    assign layer0_outputs[7691] = ~(inputs[211]) | (inputs[16]);
    assign layer0_outputs[7692] = ~((inputs[24]) | (inputs[247]));
    assign layer0_outputs[7693] = inputs[119];
    assign layer0_outputs[7694] = ~(inputs[27]);
    assign layer0_outputs[7695] = ~(inputs[189]) | (inputs[33]);
    assign layer0_outputs[7696] = inputs[160];
    assign layer0_outputs[7697] = ~(inputs[85]) | (inputs[226]);
    assign layer0_outputs[7698] = ~((inputs[224]) | (inputs[135]));
    assign layer0_outputs[7699] = (inputs[91]) & ~(inputs[160]);
    assign layer0_outputs[7700] = ~((inputs[101]) ^ (inputs[99]));
    assign layer0_outputs[7701] = ~(inputs[241]) | (inputs[66]);
    assign layer0_outputs[7702] = (inputs[21]) & ~(inputs[44]);
    assign layer0_outputs[7703] = ~(inputs[252]);
    assign layer0_outputs[7704] = (inputs[196]) | (inputs[37]);
    assign layer0_outputs[7705] = ~(inputs[183]);
    assign layer0_outputs[7706] = inputs[234];
    assign layer0_outputs[7707] = ~(inputs[229]);
    assign layer0_outputs[7708] = (inputs[70]) | (inputs[183]);
    assign layer0_outputs[7709] = ~(inputs[106]) | (inputs[128]);
    assign layer0_outputs[7710] = (inputs[126]) & ~(inputs[106]);
    assign layer0_outputs[7711] = inputs[245];
    assign layer0_outputs[7712] = ~(inputs[34]);
    assign layer0_outputs[7713] = ~((inputs[94]) | (inputs[8]));
    assign layer0_outputs[7714] = 1'b1;
    assign layer0_outputs[7715] = ~(inputs[219]);
    assign layer0_outputs[7716] = (inputs[101]) | (inputs[228]);
    assign layer0_outputs[7717] = inputs[7];
    assign layer0_outputs[7718] = (inputs[57]) & ~(inputs[252]);
    assign layer0_outputs[7719] = ~((inputs[237]) & (inputs[156]));
    assign layer0_outputs[7720] = ~(inputs[241]);
    assign layer0_outputs[7721] = (inputs[177]) ^ (inputs[246]);
    assign layer0_outputs[7722] = inputs[86];
    assign layer0_outputs[7723] = ~(inputs[216]);
    assign layer0_outputs[7724] = (inputs[39]) | (inputs[223]);
    assign layer0_outputs[7725] = ~(inputs[2]);
    assign layer0_outputs[7726] = (inputs[171]) ^ (inputs[202]);
    assign layer0_outputs[7727] = (inputs[124]) ^ (inputs[63]);
    assign layer0_outputs[7728] = inputs[235];
    assign layer0_outputs[7729] = ~(inputs[86]) | (inputs[93]);
    assign layer0_outputs[7730] = inputs[55];
    assign layer0_outputs[7731] = (inputs[224]) | (inputs[236]);
    assign layer0_outputs[7732] = (inputs[191]) | (inputs[104]);
    assign layer0_outputs[7733] = ~(inputs[147]) | (inputs[50]);
    assign layer0_outputs[7734] = ~((inputs[19]) | (inputs[123]));
    assign layer0_outputs[7735] = ~((inputs[40]) ^ (inputs[111]));
    assign layer0_outputs[7736] = (inputs[190]) | (inputs[176]);
    assign layer0_outputs[7737] = ~((inputs[125]) | (inputs[137]));
    assign layer0_outputs[7738] = ~(inputs[101]) | (inputs[185]);
    assign layer0_outputs[7739] = ~((inputs[71]) | (inputs[159]));
    assign layer0_outputs[7740] = (inputs[135]) & ~(inputs[26]);
    assign layer0_outputs[7741] = ~(inputs[111]) | (inputs[2]);
    assign layer0_outputs[7742] = (inputs[161]) & (inputs[233]);
    assign layer0_outputs[7743] = (inputs[83]) | (inputs[121]);
    assign layer0_outputs[7744] = ~(inputs[53]) | (inputs[27]);
    assign layer0_outputs[7745] = ~(inputs[100]);
    assign layer0_outputs[7746] = (inputs[84]) & ~(inputs[205]);
    assign layer0_outputs[7747] = ~(inputs[64]) | (inputs[249]);
    assign layer0_outputs[7748] = inputs[205];
    assign layer0_outputs[7749] = ~((inputs[146]) & (inputs[130]));
    assign layer0_outputs[7750] = ~((inputs[124]) ^ (inputs[36]));
    assign layer0_outputs[7751] = (inputs[178]) ^ (inputs[116]);
    assign layer0_outputs[7752] = (inputs[16]) & ~(inputs[16]);
    assign layer0_outputs[7753] = inputs[161];
    assign layer0_outputs[7754] = (inputs[13]) | (inputs[236]);
    assign layer0_outputs[7755] = ~(inputs[68]);
    assign layer0_outputs[7756] = (inputs[108]) ^ (inputs[50]);
    assign layer0_outputs[7757] = (inputs[184]) & ~(inputs[116]);
    assign layer0_outputs[7758] = ~(inputs[123]) | (inputs[195]);
    assign layer0_outputs[7759] = (inputs[196]) & ~(inputs[123]);
    assign layer0_outputs[7760] = ~(inputs[65]) | (inputs[141]);
    assign layer0_outputs[7761] = (inputs[172]) & ~(inputs[94]);
    assign layer0_outputs[7762] = (inputs[74]) & ~(inputs[158]);
    assign layer0_outputs[7763] = inputs[73];
    assign layer0_outputs[7764] = ~(inputs[42]);
    assign layer0_outputs[7765] = inputs[78];
    assign layer0_outputs[7766] = inputs[25];
    assign layer0_outputs[7767] = (inputs[170]) ^ (inputs[106]);
    assign layer0_outputs[7768] = (inputs[78]) & ~(inputs[166]);
    assign layer0_outputs[7769] = ~(inputs[228]);
    assign layer0_outputs[7770] = (inputs[234]) ^ (inputs[61]);
    assign layer0_outputs[7771] = ~(inputs[229]) | (inputs[66]);
    assign layer0_outputs[7772] = ~((inputs[54]) | (inputs[193]));
    assign layer0_outputs[7773] = inputs[83];
    assign layer0_outputs[7774] = inputs[102];
    assign layer0_outputs[7775] = (inputs[134]) | (inputs[89]);
    assign layer0_outputs[7776] = ~(inputs[91]);
    assign layer0_outputs[7777] = ~(inputs[246]);
    assign layer0_outputs[7778] = (inputs[43]) & ~(inputs[204]);
    assign layer0_outputs[7779] = (inputs[9]) & ~(inputs[144]);
    assign layer0_outputs[7780] = inputs[161];
    assign layer0_outputs[7781] = inputs[132];
    assign layer0_outputs[7782] = (inputs[174]) | (inputs[204]);
    assign layer0_outputs[7783] = ~(inputs[92]) | (inputs[209]);
    assign layer0_outputs[7784] = (inputs[143]) ^ (inputs[10]);
    assign layer0_outputs[7785] = ~(inputs[146]);
    assign layer0_outputs[7786] = (inputs[71]) ^ (inputs[21]);
    assign layer0_outputs[7787] = (inputs[253]) ^ (inputs[18]);
    assign layer0_outputs[7788] = ~(inputs[76]);
    assign layer0_outputs[7789] = ~((inputs[148]) | (inputs[93]));
    assign layer0_outputs[7790] = (inputs[27]) & ~(inputs[166]);
    assign layer0_outputs[7791] = ~(inputs[24]);
    assign layer0_outputs[7792] = inputs[197];
    assign layer0_outputs[7793] = (inputs[2]) | (inputs[223]);
    assign layer0_outputs[7794] = ~((inputs[142]) | (inputs[84]));
    assign layer0_outputs[7795] = inputs[30];
    assign layer0_outputs[7796] = (inputs[64]) & (inputs[49]);
    assign layer0_outputs[7797] = 1'b0;
    assign layer0_outputs[7798] = (inputs[204]) & ~(inputs[40]);
    assign layer0_outputs[7799] = (inputs[235]) ^ (inputs[150]);
    assign layer0_outputs[7800] = inputs[29];
    assign layer0_outputs[7801] = inputs[57];
    assign layer0_outputs[7802] = ~(inputs[120]);
    assign layer0_outputs[7803] = inputs[123];
    assign layer0_outputs[7804] = ~(inputs[38]);
    assign layer0_outputs[7805] = ~((inputs[212]) | (inputs[238]));
    assign layer0_outputs[7806] = ~(inputs[193]);
    assign layer0_outputs[7807] = (inputs[44]) & ~(inputs[176]);
    assign layer0_outputs[7808] = ~(inputs[60]) | (inputs[118]);
    assign layer0_outputs[7809] = inputs[119];
    assign layer0_outputs[7810] = ~((inputs[67]) | (inputs[218]));
    assign layer0_outputs[7811] = inputs[70];
    assign layer0_outputs[7812] = inputs[29];
    assign layer0_outputs[7813] = ~((inputs[179]) | (inputs[170]));
    assign layer0_outputs[7814] = (inputs[162]) | (inputs[24]);
    assign layer0_outputs[7815] = ~(inputs[210]);
    assign layer0_outputs[7816] = inputs[91];
    assign layer0_outputs[7817] = (inputs[71]) ^ (inputs[218]);
    assign layer0_outputs[7818] = ~(inputs[133]);
    assign layer0_outputs[7819] = (inputs[54]) ^ (inputs[252]);
    assign layer0_outputs[7820] = (inputs[68]) ^ (inputs[51]);
    assign layer0_outputs[7821] = ~((inputs[217]) | (inputs[208]));
    assign layer0_outputs[7822] = inputs[194];
    assign layer0_outputs[7823] = (inputs[188]) | (inputs[86]);
    assign layer0_outputs[7824] = (inputs[182]) | (inputs[83]);
    assign layer0_outputs[7825] = (inputs[54]) & ~(inputs[29]);
    assign layer0_outputs[7826] = ~((inputs[35]) ^ (inputs[192]));
    assign layer0_outputs[7827] = ~(inputs[160]);
    assign layer0_outputs[7828] = ~(inputs[249]);
    assign layer0_outputs[7829] = (inputs[61]) & ~(inputs[132]);
    assign layer0_outputs[7830] = ~(inputs[241]);
    assign layer0_outputs[7831] = ~(inputs[100]);
    assign layer0_outputs[7832] = ~((inputs[171]) & (inputs[178]));
    assign layer0_outputs[7833] = inputs[250];
    assign layer0_outputs[7834] = (inputs[239]) | (inputs[176]);
    assign layer0_outputs[7835] = ~((inputs[231]) | (inputs[94]));
    assign layer0_outputs[7836] = ~(inputs[114]);
    assign layer0_outputs[7837] = ~(inputs[179]);
    assign layer0_outputs[7838] = 1'b0;
    assign layer0_outputs[7839] = ~(inputs[56]);
    assign layer0_outputs[7840] = ~(inputs[227]);
    assign layer0_outputs[7841] = inputs[7];
    assign layer0_outputs[7842] = ~((inputs[26]) ^ (inputs[207]));
    assign layer0_outputs[7843] = (inputs[96]) & (inputs[224]);
    assign layer0_outputs[7844] = (inputs[42]) | (inputs[214]);
    assign layer0_outputs[7845] = (inputs[36]) | (inputs[126]);
    assign layer0_outputs[7846] = ~((inputs[169]) ^ (inputs[149]));
    assign layer0_outputs[7847] = ~((inputs[222]) ^ (inputs[62]));
    assign layer0_outputs[7848] = ~((inputs[23]) | (inputs[6]));
    assign layer0_outputs[7849] = ~(inputs[28]) | (inputs[192]);
    assign layer0_outputs[7850] = (inputs[141]) & ~(inputs[222]);
    assign layer0_outputs[7851] = (inputs[127]) ^ (inputs[27]);
    assign layer0_outputs[7852] = (inputs[143]) | (inputs[3]);
    assign layer0_outputs[7853] = (inputs[202]) ^ (inputs[213]);
    assign layer0_outputs[7854] = ~((inputs[96]) ^ (inputs[130]));
    assign layer0_outputs[7855] = ~(inputs[119]);
    assign layer0_outputs[7856] = (inputs[65]) | (inputs[68]);
    assign layer0_outputs[7857] = (inputs[68]) | (inputs[125]);
    assign layer0_outputs[7858] = ~((inputs[65]) | (inputs[238]));
    assign layer0_outputs[7859] = ~((inputs[23]) | (inputs[225]));
    assign layer0_outputs[7860] = (inputs[155]) | (inputs[18]);
    assign layer0_outputs[7861] = (inputs[204]) | (inputs[174]);
    assign layer0_outputs[7862] = 1'b0;
    assign layer0_outputs[7863] = ~(inputs[80]);
    assign layer0_outputs[7864] = (inputs[101]) & (inputs[198]);
    assign layer0_outputs[7865] = (inputs[121]) & (inputs[212]);
    assign layer0_outputs[7866] = (inputs[4]) & ~(inputs[176]);
    assign layer0_outputs[7867] = ~(inputs[140]);
    assign layer0_outputs[7868] = ~((inputs[110]) | (inputs[3]));
    assign layer0_outputs[7869] = ~(inputs[9]);
    assign layer0_outputs[7870] = 1'b1;
    assign layer0_outputs[7871] = ~(inputs[136]) | (inputs[241]);
    assign layer0_outputs[7872] = inputs[74];
    assign layer0_outputs[7873] = (inputs[244]) & ~(inputs[35]);
    assign layer0_outputs[7874] = ~(inputs[149]);
    assign layer0_outputs[7875] = ~(inputs[8]) | (inputs[83]);
    assign layer0_outputs[7876] = inputs[105];
    assign layer0_outputs[7877] = 1'b0;
    assign layer0_outputs[7878] = ~(inputs[41]);
    assign layer0_outputs[7879] = (inputs[117]) | (inputs[87]);
    assign layer0_outputs[7880] = 1'b0;
    assign layer0_outputs[7881] = inputs[0];
    assign layer0_outputs[7882] = (inputs[204]) & ~(inputs[127]);
    assign layer0_outputs[7883] = ~(inputs[68]) | (inputs[18]);
    assign layer0_outputs[7884] = ~((inputs[103]) ^ (inputs[255]));
    assign layer0_outputs[7885] = ~(inputs[166]);
    assign layer0_outputs[7886] = ~((inputs[196]) | (inputs[53]));
    assign layer0_outputs[7887] = (inputs[248]) | (inputs[192]);
    assign layer0_outputs[7888] = inputs[76];
    assign layer0_outputs[7889] = (inputs[45]) | (inputs[88]);
    assign layer0_outputs[7890] = 1'b1;
    assign layer0_outputs[7891] = (inputs[42]) & ~(inputs[162]);
    assign layer0_outputs[7892] = ~(inputs[22]) | (inputs[81]);
    assign layer0_outputs[7893] = (inputs[180]) | (inputs[23]);
    assign layer0_outputs[7894] = ~((inputs[232]) | (inputs[211]));
    assign layer0_outputs[7895] = (inputs[59]) | (inputs[109]);
    assign layer0_outputs[7896] = ~(inputs[113]);
    assign layer0_outputs[7897] = ~((inputs[190]) ^ (inputs[211]));
    assign layer0_outputs[7898] = ~((inputs[63]) ^ (inputs[18]));
    assign layer0_outputs[7899] = (inputs[249]) | (inputs[100]);
    assign layer0_outputs[7900] = inputs[167];
    assign layer0_outputs[7901] = ~((inputs[1]) | (inputs[55]));
    assign layer0_outputs[7902] = ~(inputs[113]);
    assign layer0_outputs[7903] = ~((inputs[129]) | (inputs[203]));
    assign layer0_outputs[7904] = ~(inputs[199]) | (inputs[13]);
    assign layer0_outputs[7905] = inputs[248];
    assign layer0_outputs[7906] = (inputs[187]) | (inputs[154]);
    assign layer0_outputs[7907] = ~((inputs[54]) & (inputs[112]));
    assign layer0_outputs[7908] = inputs[37];
    assign layer0_outputs[7909] = ~((inputs[41]) | (inputs[35]));
    assign layer0_outputs[7910] = ~((inputs[102]) | (inputs[97]));
    assign layer0_outputs[7911] = ~(inputs[134]);
    assign layer0_outputs[7912] = ~((inputs[14]) | (inputs[151]));
    assign layer0_outputs[7913] = ~((inputs[177]) | (inputs[245]));
    assign layer0_outputs[7914] = ~((inputs[11]) ^ (inputs[98]));
    assign layer0_outputs[7915] = ~(inputs[34]) | (inputs[239]);
    assign layer0_outputs[7916] = inputs[30];
    assign layer0_outputs[7917] = ~(inputs[224]) | (inputs[125]);
    assign layer0_outputs[7918] = ~((inputs[71]) ^ (inputs[101]));
    assign layer0_outputs[7919] = inputs[86];
    assign layer0_outputs[7920] = (inputs[181]) & ~(inputs[108]);
    assign layer0_outputs[7921] = ~(inputs[164]);
    assign layer0_outputs[7922] = (inputs[26]) & ~(inputs[163]);
    assign layer0_outputs[7923] = (inputs[185]) & ~(inputs[52]);
    assign layer0_outputs[7924] = ~(inputs[23]);
    assign layer0_outputs[7925] = ~(inputs[9]);
    assign layer0_outputs[7926] = ~(inputs[146]) | (inputs[138]);
    assign layer0_outputs[7927] = (inputs[64]) & (inputs[208]);
    assign layer0_outputs[7928] = ~((inputs[115]) & (inputs[213]));
    assign layer0_outputs[7929] = inputs[203];
    assign layer0_outputs[7930] = ~(inputs[142]);
    assign layer0_outputs[7931] = ~((inputs[158]) | (inputs[63]));
    assign layer0_outputs[7932] = ~((inputs[38]) ^ (inputs[72]));
    assign layer0_outputs[7933] = inputs[10];
    assign layer0_outputs[7934] = ~((inputs[240]) & (inputs[236]));
    assign layer0_outputs[7935] = (inputs[88]) & ~(inputs[49]);
    assign layer0_outputs[7936] = (inputs[79]) | (inputs[218]);
    assign layer0_outputs[7937] = inputs[123];
    assign layer0_outputs[7938] = ~(inputs[223]);
    assign layer0_outputs[7939] = (inputs[197]) | (inputs[144]);
    assign layer0_outputs[7940] = ~(inputs[25]);
    assign layer0_outputs[7941] = ~((inputs[151]) | (inputs[1]));
    assign layer0_outputs[7942] = ~(inputs[178]);
    assign layer0_outputs[7943] = (inputs[159]) | (inputs[161]);
    assign layer0_outputs[7944] = (inputs[224]) | (inputs[250]);
    assign layer0_outputs[7945] = ~(inputs[91]);
    assign layer0_outputs[7946] = (inputs[231]) & ~(inputs[220]);
    assign layer0_outputs[7947] = ~(inputs[167]);
    assign layer0_outputs[7948] = ~(inputs[48]);
    assign layer0_outputs[7949] = (inputs[229]) & ~(inputs[136]);
    assign layer0_outputs[7950] = (inputs[205]) ^ (inputs[10]);
    assign layer0_outputs[7951] = ~((inputs[144]) | (inputs[49]));
    assign layer0_outputs[7952] = (inputs[74]) | (inputs[110]);
    assign layer0_outputs[7953] = inputs[56];
    assign layer0_outputs[7954] = inputs[114];
    assign layer0_outputs[7955] = ~(inputs[164]);
    assign layer0_outputs[7956] = inputs[211];
    assign layer0_outputs[7957] = ~(inputs[183]) | (inputs[15]);
    assign layer0_outputs[7958] = ~((inputs[228]) | (inputs[148]));
    assign layer0_outputs[7959] = ~((inputs[251]) | (inputs[85]));
    assign layer0_outputs[7960] = (inputs[170]) & ~(inputs[32]);
    assign layer0_outputs[7961] = (inputs[148]) & ~(inputs[178]);
    assign layer0_outputs[7962] = inputs[173];
    assign layer0_outputs[7963] = (inputs[36]) & ~(inputs[148]);
    assign layer0_outputs[7964] = ~(inputs[217]);
    assign layer0_outputs[7965] = inputs[39];
    assign layer0_outputs[7966] = (inputs[1]) ^ (inputs[222]);
    assign layer0_outputs[7967] = inputs[209];
    assign layer0_outputs[7968] = ~(inputs[83]);
    assign layer0_outputs[7969] = ~((inputs[50]) & (inputs[64]));
    assign layer0_outputs[7970] = ~((inputs[198]) ^ (inputs[249]));
    assign layer0_outputs[7971] = ~(inputs[222]);
    assign layer0_outputs[7972] = ~((inputs[171]) ^ (inputs[1]));
    assign layer0_outputs[7973] = (inputs[193]) & ~(inputs[81]);
    assign layer0_outputs[7974] = ~(inputs[22]);
    assign layer0_outputs[7975] = (inputs[248]) & ~(inputs[251]);
    assign layer0_outputs[7976] = ~(inputs[218]);
    assign layer0_outputs[7977] = ~(inputs[139]);
    assign layer0_outputs[7978] = inputs[79];
    assign layer0_outputs[7979] = (inputs[20]) ^ (inputs[176]);
    assign layer0_outputs[7980] = ~(inputs[179]);
    assign layer0_outputs[7981] = (inputs[161]) | (inputs[215]);
    assign layer0_outputs[7982] = (inputs[100]) | (inputs[174]);
    assign layer0_outputs[7983] = inputs[229];
    assign layer0_outputs[7984] = inputs[181];
    assign layer0_outputs[7985] = ~(inputs[150]);
    assign layer0_outputs[7986] = (inputs[193]) & ~(inputs[245]);
    assign layer0_outputs[7987] = (inputs[172]) | (inputs[33]);
    assign layer0_outputs[7988] = (inputs[144]) & ~(inputs[62]);
    assign layer0_outputs[7989] = 1'b1;
    assign layer0_outputs[7990] = (inputs[16]) ^ (inputs[248]);
    assign layer0_outputs[7991] = ~((inputs[10]) | (inputs[141]));
    assign layer0_outputs[7992] = ~((inputs[157]) | (inputs[101]));
    assign layer0_outputs[7993] = (inputs[236]) & ~(inputs[249]);
    assign layer0_outputs[7994] = (inputs[171]) | (inputs[98]);
    assign layer0_outputs[7995] = inputs[91];
    assign layer0_outputs[7996] = (inputs[115]) & ~(inputs[202]);
    assign layer0_outputs[7997] = ~(inputs[195]);
    assign layer0_outputs[7998] = ~((inputs[17]) | (inputs[45]));
    assign layer0_outputs[7999] = ~((inputs[126]) ^ (inputs[48]));
    assign layer0_outputs[8000] = inputs[30];
    assign layer0_outputs[8001] = ~(inputs[169]) | (inputs[15]);
    assign layer0_outputs[8002] = ~(inputs[49]) | (inputs[1]);
    assign layer0_outputs[8003] = ~(inputs[186]) | (inputs[192]);
    assign layer0_outputs[8004] = (inputs[62]) | (inputs[33]);
    assign layer0_outputs[8005] = ~(inputs[59]);
    assign layer0_outputs[8006] = ~(inputs[16]);
    assign layer0_outputs[8007] = (inputs[88]) & ~(inputs[147]);
    assign layer0_outputs[8008] = ~(inputs[41]);
    assign layer0_outputs[8009] = (inputs[255]) | (inputs[147]);
    assign layer0_outputs[8010] = (inputs[184]) & ~(inputs[78]);
    assign layer0_outputs[8011] = (inputs[245]) | (inputs[81]);
    assign layer0_outputs[8012] = ~((inputs[125]) ^ (inputs[86]));
    assign layer0_outputs[8013] = ~(inputs[68]) | (inputs[166]);
    assign layer0_outputs[8014] = (inputs[173]) & ~(inputs[16]);
    assign layer0_outputs[8015] = (inputs[220]) & ~(inputs[91]);
    assign layer0_outputs[8016] = ~((inputs[194]) ^ (inputs[123]));
    assign layer0_outputs[8017] = ~((inputs[61]) | (inputs[95]));
    assign layer0_outputs[8018] = (inputs[75]) & (inputs[79]);
    assign layer0_outputs[8019] = (inputs[248]) | (inputs[208]);
    assign layer0_outputs[8020] = ~((inputs[80]) ^ (inputs[6]));
    assign layer0_outputs[8021] = ~((inputs[102]) ^ (inputs[148]));
    assign layer0_outputs[8022] = inputs[188];
    assign layer0_outputs[8023] = ~(inputs[87]) | (inputs[64]);
    assign layer0_outputs[8024] = (inputs[208]) & ~(inputs[0]);
    assign layer0_outputs[8025] = ~((inputs[190]) | (inputs[95]));
    assign layer0_outputs[8026] = ~(inputs[98]);
    assign layer0_outputs[8027] = ~(inputs[107]) | (inputs[114]);
    assign layer0_outputs[8028] = ~((inputs[206]) ^ (inputs[175]));
    assign layer0_outputs[8029] = ~((inputs[196]) | (inputs[33]));
    assign layer0_outputs[8030] = ~(inputs[24]);
    assign layer0_outputs[8031] = (inputs[179]) & ~(inputs[17]);
    assign layer0_outputs[8032] = ~((inputs[227]) ^ (inputs[1]));
    assign layer0_outputs[8033] = ~((inputs[18]) ^ (inputs[195]));
    assign layer0_outputs[8034] = (inputs[199]) ^ (inputs[181]);
    assign layer0_outputs[8035] = ~((inputs[114]) | (inputs[91]));
    assign layer0_outputs[8036] = inputs[127];
    assign layer0_outputs[8037] = ~((inputs[159]) ^ (inputs[101]));
    assign layer0_outputs[8038] = (inputs[0]) & ~(inputs[255]);
    assign layer0_outputs[8039] = (inputs[36]) ^ (inputs[128]);
    assign layer0_outputs[8040] = inputs[246];
    assign layer0_outputs[8041] = ~((inputs[126]) | (inputs[236]));
    assign layer0_outputs[8042] = ~((inputs[207]) | (inputs[227]));
    assign layer0_outputs[8043] = inputs[25];
    assign layer0_outputs[8044] = ~(inputs[79]);
    assign layer0_outputs[8045] = ~(inputs[45]) | (inputs[55]);
    assign layer0_outputs[8046] = ~((inputs[157]) ^ (inputs[115]));
    assign layer0_outputs[8047] = 1'b0;
    assign layer0_outputs[8048] = ~((inputs[251]) | (inputs[245]));
    assign layer0_outputs[8049] = (inputs[234]) & ~(inputs[165]);
    assign layer0_outputs[8050] = (inputs[23]) ^ (inputs[66]);
    assign layer0_outputs[8051] = ~(inputs[173]) | (inputs[178]);
    assign layer0_outputs[8052] = ~(inputs[221]);
    assign layer0_outputs[8053] = inputs[121];
    assign layer0_outputs[8054] = ~(inputs[59]);
    assign layer0_outputs[8055] = ~(inputs[82]);
    assign layer0_outputs[8056] = (inputs[157]) ^ (inputs[36]);
    assign layer0_outputs[8057] = inputs[180];
    assign layer0_outputs[8058] = (inputs[204]) ^ (inputs[225]);
    assign layer0_outputs[8059] = 1'b0;
    assign layer0_outputs[8060] = ~(inputs[130]) | (inputs[222]);
    assign layer0_outputs[8061] = ~(inputs[142]);
    assign layer0_outputs[8062] = ~(inputs[69]);
    assign layer0_outputs[8063] = inputs[164];
    assign layer0_outputs[8064] = (inputs[194]) ^ (inputs[235]);
    assign layer0_outputs[8065] = ~(inputs[90]);
    assign layer0_outputs[8066] = (inputs[149]) ^ (inputs[189]);
    assign layer0_outputs[8067] = inputs[82];
    assign layer0_outputs[8068] = (inputs[28]) & (inputs[69]);
    assign layer0_outputs[8069] = ~(inputs[41]);
    assign layer0_outputs[8070] = ~(inputs[222]);
    assign layer0_outputs[8071] = ~(inputs[201]);
    assign layer0_outputs[8072] = (inputs[251]) & ~(inputs[241]);
    assign layer0_outputs[8073] = (inputs[65]) | (inputs[83]);
    assign layer0_outputs[8074] = ~((inputs[143]) & (inputs[60]));
    assign layer0_outputs[8075] = (inputs[55]) & ~(inputs[34]);
    assign layer0_outputs[8076] = (inputs[196]) | (inputs[248]);
    assign layer0_outputs[8077] = ~(inputs[220]) | (inputs[87]);
    assign layer0_outputs[8078] = inputs[10];
    assign layer0_outputs[8079] = ~((inputs[13]) | (inputs[144]));
    assign layer0_outputs[8080] = inputs[67];
    assign layer0_outputs[8081] = ~(inputs[67]) | (inputs[73]);
    assign layer0_outputs[8082] = ~((inputs[197]) | (inputs[7]));
    assign layer0_outputs[8083] = ~(inputs[206]) | (inputs[112]);
    assign layer0_outputs[8084] = ~((inputs[255]) | (inputs[143]));
    assign layer0_outputs[8085] = (inputs[123]) & ~(inputs[178]);
    assign layer0_outputs[8086] = ~((inputs[246]) ^ (inputs[169]));
    assign layer0_outputs[8087] = ~(inputs[129]) | (inputs[102]);
    assign layer0_outputs[8088] = ~(inputs[90]);
    assign layer0_outputs[8089] = ~(inputs[214]) | (inputs[123]);
    assign layer0_outputs[8090] = (inputs[123]) | (inputs[20]);
    assign layer0_outputs[8091] = ~(inputs[57]) | (inputs[188]);
    assign layer0_outputs[8092] = inputs[142];
    assign layer0_outputs[8093] = inputs[232];
    assign layer0_outputs[8094] = (inputs[176]) ^ (inputs[171]);
    assign layer0_outputs[8095] = (inputs[63]) | (inputs[48]);
    assign layer0_outputs[8096] = ~(inputs[166]);
    assign layer0_outputs[8097] = ~((inputs[52]) | (inputs[206]));
    assign layer0_outputs[8098] = (inputs[190]) & (inputs[45]);
    assign layer0_outputs[8099] = (inputs[103]) ^ (inputs[73]);
    assign layer0_outputs[8100] = ~((inputs[181]) | (inputs[65]));
    assign layer0_outputs[8101] = (inputs[229]) & ~(inputs[95]);
    assign layer0_outputs[8102] = inputs[40];
    assign layer0_outputs[8103] = ~(inputs[35]) | (inputs[83]);
    assign layer0_outputs[8104] = ~((inputs[193]) | (inputs[2]));
    assign layer0_outputs[8105] = ~(inputs[74]);
    assign layer0_outputs[8106] = ~(inputs[158]);
    assign layer0_outputs[8107] = ~((inputs[104]) | (inputs[174]));
    assign layer0_outputs[8108] = ~(inputs[162]);
    assign layer0_outputs[8109] = ~(inputs[24]) | (inputs[228]);
    assign layer0_outputs[8110] = ~((inputs[125]) ^ (inputs[240]));
    assign layer0_outputs[8111] = ~(inputs[133]) | (inputs[31]);
    assign layer0_outputs[8112] = ~(inputs[223]) | (inputs[200]);
    assign layer0_outputs[8113] = ~(inputs[104]) | (inputs[167]);
    assign layer0_outputs[8114] = (inputs[122]) ^ (inputs[239]);
    assign layer0_outputs[8115] = ~((inputs[137]) & (inputs[209]));
    assign layer0_outputs[8116] = (inputs[117]) & ~(inputs[147]);
    assign layer0_outputs[8117] = (inputs[40]) | (inputs[23]);
    assign layer0_outputs[8118] = ~(inputs[156]);
    assign layer0_outputs[8119] = ~(inputs[163]) | (inputs[83]);
    assign layer0_outputs[8120] = (inputs[169]) ^ (inputs[50]);
    assign layer0_outputs[8121] = (inputs[215]) | (inputs[237]);
    assign layer0_outputs[8122] = ~(inputs[87]) | (inputs[34]);
    assign layer0_outputs[8123] = ~(inputs[1]);
    assign layer0_outputs[8124] = ~((inputs[163]) ^ (inputs[170]));
    assign layer0_outputs[8125] = ~((inputs[121]) ^ (inputs[101]));
    assign layer0_outputs[8126] = inputs[112];
    assign layer0_outputs[8127] = ~((inputs[104]) ^ (inputs[148]));
    assign layer0_outputs[8128] = inputs[177];
    assign layer0_outputs[8129] = inputs[78];
    assign layer0_outputs[8130] = (inputs[69]) | (inputs[208]);
    assign layer0_outputs[8131] = ~(inputs[176]) | (inputs[35]);
    assign layer0_outputs[8132] = inputs[136];
    assign layer0_outputs[8133] = ~((inputs[138]) | (inputs[165]));
    assign layer0_outputs[8134] = (inputs[155]) ^ (inputs[238]);
    assign layer0_outputs[8135] = ~(inputs[206]);
    assign layer0_outputs[8136] = (inputs[240]) ^ (inputs[21]);
    assign layer0_outputs[8137] = ~(inputs[123]);
    assign layer0_outputs[8138] = 1'b1;
    assign layer0_outputs[8139] = ~((inputs[71]) ^ (inputs[227]));
    assign layer0_outputs[8140] = (inputs[231]) & ~(inputs[140]);
    assign layer0_outputs[8141] = inputs[22];
    assign layer0_outputs[8142] = ~(inputs[151]);
    assign layer0_outputs[8143] = (inputs[0]) ^ (inputs[246]);
    assign layer0_outputs[8144] = ~((inputs[19]) ^ (inputs[72]));
    assign layer0_outputs[8145] = inputs[212];
    assign layer0_outputs[8146] = (inputs[124]) & ~(inputs[12]);
    assign layer0_outputs[8147] = (inputs[224]) | (inputs[137]);
    assign layer0_outputs[8148] = ~(inputs[68]) | (inputs[106]);
    assign layer0_outputs[8149] = (inputs[95]) | (inputs[61]);
    assign layer0_outputs[8150] = (inputs[2]) | (inputs[35]);
    assign layer0_outputs[8151] = (inputs[29]) | (inputs[188]);
    assign layer0_outputs[8152] = ~(inputs[111]);
    assign layer0_outputs[8153] = inputs[250];
    assign layer0_outputs[8154] = (inputs[85]) | (inputs[194]);
    assign layer0_outputs[8155] = ~((inputs[51]) | (inputs[112]));
    assign layer0_outputs[8156] = ~(inputs[90]) | (inputs[239]);
    assign layer0_outputs[8157] = ~((inputs[64]) | (inputs[214]));
    assign layer0_outputs[8158] = (inputs[192]) & ~(inputs[251]);
    assign layer0_outputs[8159] = inputs[110];
    assign layer0_outputs[8160] = (inputs[203]) ^ (inputs[171]);
    assign layer0_outputs[8161] = (inputs[178]) & ~(inputs[60]);
    assign layer0_outputs[8162] = ~((inputs[156]) ^ (inputs[157]));
    assign layer0_outputs[8163] = ~((inputs[67]) ^ (inputs[69]));
    assign layer0_outputs[8164] = inputs[206];
    assign layer0_outputs[8165] = (inputs[189]) & ~(inputs[254]);
    assign layer0_outputs[8166] = ~(inputs[142]);
    assign layer0_outputs[8167] = (inputs[7]) & ~(inputs[225]);
    assign layer0_outputs[8168] = ~((inputs[52]) ^ (inputs[33]));
    assign layer0_outputs[8169] = inputs[110];
    assign layer0_outputs[8170] = ~((inputs[140]) & (inputs[131]));
    assign layer0_outputs[8171] = ~(inputs[119]);
    assign layer0_outputs[8172] = (inputs[218]) & ~(inputs[25]);
    assign layer0_outputs[8173] = ~(inputs[22]);
    assign layer0_outputs[8174] = ~((inputs[152]) | (inputs[177]));
    assign layer0_outputs[8175] = ~(inputs[44]);
    assign layer0_outputs[8176] = ~(inputs[14]);
    assign layer0_outputs[8177] = ~(inputs[234]) | (inputs[78]);
    assign layer0_outputs[8178] = ~((inputs[234]) ^ (inputs[62]));
    assign layer0_outputs[8179] = (inputs[197]) & ~(inputs[116]);
    assign layer0_outputs[8180] = ~(inputs[230]) | (inputs[156]);
    assign layer0_outputs[8181] = (inputs[29]) & ~(inputs[32]);
    assign layer0_outputs[8182] = inputs[62];
    assign layer0_outputs[8183] = ~(inputs[129]) | (inputs[223]);
    assign layer0_outputs[8184] = ~(inputs[243]) | (inputs[14]);
    assign layer0_outputs[8185] = (inputs[126]) | (inputs[242]);
    assign layer0_outputs[8186] = ~(inputs[41]) | (inputs[127]);
    assign layer0_outputs[8187] = (inputs[63]) ^ (inputs[248]);
    assign layer0_outputs[8188] = ~((inputs[195]) | (inputs[239]));
    assign layer0_outputs[8189] = ~((inputs[7]) ^ (inputs[74]));
    assign layer0_outputs[8190] = ~(inputs[137]) | (inputs[28]);
    assign layer0_outputs[8191] = (inputs[96]) ^ (inputs[23]);
    assign layer0_outputs[8192] = (inputs[234]) | (inputs[194]);
    assign layer0_outputs[8193] = (inputs[248]) | (inputs[65]);
    assign layer0_outputs[8194] = ~((inputs[58]) | (inputs[59]));
    assign layer0_outputs[8195] = (inputs[86]) & (inputs[176]);
    assign layer0_outputs[8196] = ~((inputs[179]) | (inputs[176]));
    assign layer0_outputs[8197] = inputs[0];
    assign layer0_outputs[8198] = (inputs[202]) | (inputs[241]);
    assign layer0_outputs[8199] = (inputs[247]) & ~(inputs[22]);
    assign layer0_outputs[8200] = (inputs[99]) & (inputs[83]);
    assign layer0_outputs[8201] = ~(inputs[204]) | (inputs[225]);
    assign layer0_outputs[8202] = inputs[118];
    assign layer0_outputs[8203] = ~(inputs[165]) | (inputs[255]);
    assign layer0_outputs[8204] = (inputs[200]) & (inputs[197]);
    assign layer0_outputs[8205] = ~(inputs[213]) | (inputs[206]);
    assign layer0_outputs[8206] = (inputs[159]) ^ (inputs[214]);
    assign layer0_outputs[8207] = (inputs[182]) & ~(inputs[8]);
    assign layer0_outputs[8208] = 1'b1;
    assign layer0_outputs[8209] = (inputs[131]) | (inputs[12]);
    assign layer0_outputs[8210] = ~(inputs[119]) | (inputs[0]);
    assign layer0_outputs[8211] = ~(inputs[210]) | (inputs[254]);
    assign layer0_outputs[8212] = ~(inputs[54]);
    assign layer0_outputs[8213] = ~(inputs[97]) | (inputs[62]);
    assign layer0_outputs[8214] = (inputs[170]) | (inputs[165]);
    assign layer0_outputs[8215] = inputs[196];
    assign layer0_outputs[8216] = (inputs[88]) | (inputs[223]);
    assign layer0_outputs[8217] = inputs[83];
    assign layer0_outputs[8218] = (inputs[178]) | (inputs[92]);
    assign layer0_outputs[8219] = ~(inputs[76]);
    assign layer0_outputs[8220] = ~(inputs[181]);
    assign layer0_outputs[8221] = (inputs[225]) & ~(inputs[63]);
    assign layer0_outputs[8222] = ~(inputs[149]) | (inputs[207]);
    assign layer0_outputs[8223] = ~(inputs[154]);
    assign layer0_outputs[8224] = ~(inputs[66]);
    assign layer0_outputs[8225] = inputs[198];
    assign layer0_outputs[8226] = ~((inputs[13]) ^ (inputs[57]));
    assign layer0_outputs[8227] = ~(inputs[194]);
    assign layer0_outputs[8228] = (inputs[20]) & (inputs[242]);
    assign layer0_outputs[8229] = ~((inputs[111]) | (inputs[13]));
    assign layer0_outputs[8230] = (inputs[39]) & ~(inputs[226]);
    assign layer0_outputs[8231] = (inputs[20]) ^ (inputs[65]);
    assign layer0_outputs[8232] = (inputs[159]) | (inputs[26]);
    assign layer0_outputs[8233] = (inputs[160]) & ~(inputs[137]);
    assign layer0_outputs[8234] = ~(inputs[56]);
    assign layer0_outputs[8235] = ~(inputs[46]);
    assign layer0_outputs[8236] = inputs[119];
    assign layer0_outputs[8237] = (inputs[74]) & ~(inputs[47]);
    assign layer0_outputs[8238] = ~((inputs[149]) ^ (inputs[138]));
    assign layer0_outputs[8239] = inputs[50];
    assign layer0_outputs[8240] = ~(inputs[47]) | (inputs[221]);
    assign layer0_outputs[8241] = ~(inputs[113]);
    assign layer0_outputs[8242] = (inputs[89]) & ~(inputs[209]);
    assign layer0_outputs[8243] = ~((inputs[6]) ^ (inputs[133]));
    assign layer0_outputs[8244] = (inputs[245]) ^ (inputs[213]);
    assign layer0_outputs[8245] = (inputs[195]) ^ (inputs[211]);
    assign layer0_outputs[8246] = (inputs[102]) & ~(inputs[73]);
    assign layer0_outputs[8247] = ~(inputs[44]);
    assign layer0_outputs[8248] = inputs[22];
    assign layer0_outputs[8249] = (inputs[216]) & ~(inputs[44]);
    assign layer0_outputs[8250] = ~(inputs[176]);
    assign layer0_outputs[8251] = ~(inputs[217]);
    assign layer0_outputs[8252] = ~((inputs[22]) | (inputs[36]));
    assign layer0_outputs[8253] = (inputs[162]) & ~(inputs[64]);
    assign layer0_outputs[8254] = ~(inputs[221]) | (inputs[152]);
    assign layer0_outputs[8255] = inputs[91];
    assign layer0_outputs[8256] = ~((inputs[230]) ^ (inputs[195]));
    assign layer0_outputs[8257] = (inputs[50]) | (inputs[115]);
    assign layer0_outputs[8258] = inputs[152];
    assign layer0_outputs[8259] = ~(inputs[93]) | (inputs[79]);
    assign layer0_outputs[8260] = (inputs[10]) ^ (inputs[254]);
    assign layer0_outputs[8261] = (inputs[88]) & (inputs[44]);
    assign layer0_outputs[8262] = (inputs[172]) ^ (inputs[115]);
    assign layer0_outputs[8263] = ~(inputs[116]);
    assign layer0_outputs[8264] = 1'b1;
    assign layer0_outputs[8265] = ~((inputs[135]) & (inputs[5]));
    assign layer0_outputs[8266] = (inputs[118]) | (inputs[234]);
    assign layer0_outputs[8267] = ~((inputs[252]) | (inputs[39]));
    assign layer0_outputs[8268] = inputs[160];
    assign layer0_outputs[8269] = ~(inputs[246]);
    assign layer0_outputs[8270] = ~(inputs[77]);
    assign layer0_outputs[8271] = ~(inputs[45]) | (inputs[138]);
    assign layer0_outputs[8272] = ~((inputs[57]) | (inputs[240]));
    assign layer0_outputs[8273] = (inputs[130]) & (inputs[211]);
    assign layer0_outputs[8274] = ~((inputs[94]) ^ (inputs[219]));
    assign layer0_outputs[8275] = 1'b1;
    assign layer0_outputs[8276] = ~((inputs[197]) ^ (inputs[1]));
    assign layer0_outputs[8277] = (inputs[73]) & ~(inputs[15]);
    assign layer0_outputs[8278] = (inputs[107]) | (inputs[37]);
    assign layer0_outputs[8279] = ~(inputs[55]) | (inputs[132]);
    assign layer0_outputs[8280] = ~(inputs[20]) | (inputs[188]);
    assign layer0_outputs[8281] = inputs[150];
    assign layer0_outputs[8282] = (inputs[27]) ^ (inputs[166]);
    assign layer0_outputs[8283] = ~(inputs[252]);
    assign layer0_outputs[8284] = ~((inputs[193]) | (inputs[161]));
    assign layer0_outputs[8285] = (inputs[89]) ^ (inputs[118]);
    assign layer0_outputs[8286] = inputs[118];
    assign layer0_outputs[8287] = (inputs[122]) & ~(inputs[112]);
    assign layer0_outputs[8288] = ~(inputs[174]);
    assign layer0_outputs[8289] = (inputs[234]) ^ (inputs[221]);
    assign layer0_outputs[8290] = ~(inputs[247]);
    assign layer0_outputs[8291] = inputs[22];
    assign layer0_outputs[8292] = ~(inputs[110]) | (inputs[243]);
    assign layer0_outputs[8293] = inputs[85];
    assign layer0_outputs[8294] = ~(inputs[70]);
    assign layer0_outputs[8295] = (inputs[144]) | (inputs[100]);
    assign layer0_outputs[8296] = (inputs[64]) | (inputs[82]);
    assign layer0_outputs[8297] = ~((inputs[18]) ^ (inputs[4]));
    assign layer0_outputs[8298] = ~((inputs[79]) | (inputs[221]));
    assign layer0_outputs[8299] = ~(inputs[137]) | (inputs[88]);
    assign layer0_outputs[8300] = (inputs[130]) & (inputs[178]);
    assign layer0_outputs[8301] = ~((inputs[117]) | (inputs[48]));
    assign layer0_outputs[8302] = ~((inputs[62]) & (inputs[86]));
    assign layer0_outputs[8303] = (inputs[248]) & ~(inputs[199]);
    assign layer0_outputs[8304] = ~((inputs[129]) | (inputs[83]));
    assign layer0_outputs[8305] = ~((inputs[25]) & (inputs[244]));
    assign layer0_outputs[8306] = (inputs[131]) & ~(inputs[229]);
    assign layer0_outputs[8307] = (inputs[79]) ^ (inputs[125]);
    assign layer0_outputs[8308] = ~(inputs[104]);
    assign layer0_outputs[8309] = (inputs[134]) & ~(inputs[93]);
    assign layer0_outputs[8310] = ~(inputs[51]);
    assign layer0_outputs[8311] = inputs[252];
    assign layer0_outputs[8312] = inputs[181];
    assign layer0_outputs[8313] = inputs[93];
    assign layer0_outputs[8314] = ~((inputs[153]) & (inputs[243]));
    assign layer0_outputs[8315] = (inputs[37]) & ~(inputs[209]);
    assign layer0_outputs[8316] = ~((inputs[213]) | (inputs[19]));
    assign layer0_outputs[8317] = ~(inputs[203]) | (inputs[87]);
    assign layer0_outputs[8318] = (inputs[195]) | (inputs[70]);
    assign layer0_outputs[8319] = (inputs[10]) | (inputs[227]);
    assign layer0_outputs[8320] = inputs[255];
    assign layer0_outputs[8321] = ~(inputs[217]) | (inputs[86]);
    assign layer0_outputs[8322] = (inputs[164]) & ~(inputs[88]);
    assign layer0_outputs[8323] = (inputs[170]) | (inputs[145]);
    assign layer0_outputs[8324] = inputs[91];
    assign layer0_outputs[8325] = ~(inputs[73]) | (inputs[4]);
    assign layer0_outputs[8326] = (inputs[219]) | (inputs[150]);
    assign layer0_outputs[8327] = ~(inputs[97]);
    assign layer0_outputs[8328] = ~((inputs[92]) | (inputs[2]));
    assign layer0_outputs[8329] = ~(inputs[246]);
    assign layer0_outputs[8330] = inputs[233];
    assign layer0_outputs[8331] = ~((inputs[248]) | (inputs[192]));
    assign layer0_outputs[8332] = ~(inputs[62]);
    assign layer0_outputs[8333] = (inputs[27]) ^ (inputs[160]);
    assign layer0_outputs[8334] = ~(inputs[31]);
    assign layer0_outputs[8335] = ~(inputs[115]);
    assign layer0_outputs[8336] = ~(inputs[232]) | (inputs[101]);
    assign layer0_outputs[8337] = ~(inputs[179]);
    assign layer0_outputs[8338] = (inputs[20]) ^ (inputs[80]);
    assign layer0_outputs[8339] = ~((inputs[34]) & (inputs[156]));
    assign layer0_outputs[8340] = inputs[157];
    assign layer0_outputs[8341] = ~(inputs[83]);
    assign layer0_outputs[8342] = (inputs[185]) ^ (inputs[196]);
    assign layer0_outputs[8343] = ~(inputs[121]) | (inputs[174]);
    assign layer0_outputs[8344] = (inputs[14]) | (inputs[83]);
    assign layer0_outputs[8345] = (inputs[77]) & ~(inputs[198]);
    assign layer0_outputs[8346] = (inputs[215]) & (inputs[214]);
    assign layer0_outputs[8347] = inputs[189];
    assign layer0_outputs[8348] = (inputs[214]) | (inputs[232]);
    assign layer0_outputs[8349] = ~((inputs[206]) ^ (inputs[165]));
    assign layer0_outputs[8350] = ~(inputs[78]);
    assign layer0_outputs[8351] = (inputs[253]) | (inputs[75]);
    assign layer0_outputs[8352] = ~((inputs[199]) ^ (inputs[241]));
    assign layer0_outputs[8353] = ~(inputs[166]);
    assign layer0_outputs[8354] = (inputs[121]) | (inputs[82]);
    assign layer0_outputs[8355] = ~(inputs[137]) | (inputs[242]);
    assign layer0_outputs[8356] = inputs[140];
    assign layer0_outputs[8357] = 1'b1;
    assign layer0_outputs[8358] = inputs[197];
    assign layer0_outputs[8359] = ~((inputs[197]) ^ (inputs[58]));
    assign layer0_outputs[8360] = (inputs[219]) & ~(inputs[122]);
    assign layer0_outputs[8361] = inputs[142];
    assign layer0_outputs[8362] = inputs[39];
    assign layer0_outputs[8363] = inputs[25];
    assign layer0_outputs[8364] = inputs[114];
    assign layer0_outputs[8365] = (inputs[73]) ^ (inputs[170]);
    assign layer0_outputs[8366] = ~((inputs[13]) | (inputs[216]));
    assign layer0_outputs[8367] = (inputs[133]) & ~(inputs[253]);
    assign layer0_outputs[8368] = inputs[196];
    assign layer0_outputs[8369] = inputs[184];
    assign layer0_outputs[8370] = ~((inputs[140]) | (inputs[58]));
    assign layer0_outputs[8371] = inputs[139];
    assign layer0_outputs[8372] = inputs[107];
    assign layer0_outputs[8373] = ~(inputs[204]) | (inputs[252]);
    assign layer0_outputs[8374] = ~(inputs[172]) | (inputs[57]);
    assign layer0_outputs[8375] = (inputs[30]) & (inputs[143]);
    assign layer0_outputs[8376] = ~((inputs[247]) | (inputs[124]));
    assign layer0_outputs[8377] = ~(inputs[109]);
    assign layer0_outputs[8378] = ~((inputs[84]) | (inputs[85]));
    assign layer0_outputs[8379] = ~(inputs[70]) | (inputs[127]);
    assign layer0_outputs[8380] = ~((inputs[193]) ^ (inputs[227]));
    assign layer0_outputs[8381] = (inputs[213]) | (inputs[205]);
    assign layer0_outputs[8382] = ~((inputs[192]) | (inputs[177]));
    assign layer0_outputs[8383] = ~(inputs[115]) | (inputs[57]);
    assign layer0_outputs[8384] = ~(inputs[211]) | (inputs[92]);
    assign layer0_outputs[8385] = ~(inputs[82]);
    assign layer0_outputs[8386] = ~(inputs[172]) | (inputs[239]);
    assign layer0_outputs[8387] = inputs[237];
    assign layer0_outputs[8388] = inputs[155];
    assign layer0_outputs[8389] = inputs[76];
    assign layer0_outputs[8390] = inputs[78];
    assign layer0_outputs[8391] = ~(inputs[35]);
    assign layer0_outputs[8392] = (inputs[7]) | (inputs[177]);
    assign layer0_outputs[8393] = ~(inputs[194]);
    assign layer0_outputs[8394] = (inputs[127]) | (inputs[163]);
    assign layer0_outputs[8395] = (inputs[132]) ^ (inputs[168]);
    assign layer0_outputs[8396] = ~(inputs[231]);
    assign layer0_outputs[8397] = ~(inputs[54]);
    assign layer0_outputs[8398] = ~((inputs[74]) | (inputs[4]));
    assign layer0_outputs[8399] = (inputs[109]) & (inputs[56]);
    assign layer0_outputs[8400] = inputs[230];
    assign layer0_outputs[8401] = inputs[40];
    assign layer0_outputs[8402] = (inputs[118]) | (inputs[244]);
    assign layer0_outputs[8403] = ~(inputs[228]);
    assign layer0_outputs[8404] = inputs[74];
    assign layer0_outputs[8405] = ~((inputs[33]) ^ (inputs[121]));
    assign layer0_outputs[8406] = (inputs[218]) | (inputs[236]);
    assign layer0_outputs[8407] = (inputs[132]) | (inputs[163]);
    assign layer0_outputs[8408] = ~(inputs[90]);
    assign layer0_outputs[8409] = (inputs[239]) | (inputs[213]);
    assign layer0_outputs[8410] = (inputs[95]) | (inputs[102]);
    assign layer0_outputs[8411] = ~(inputs[174]) | (inputs[189]);
    assign layer0_outputs[8412] = ~((inputs[232]) | (inputs[87]));
    assign layer0_outputs[8413] = ~(inputs[84]) | (inputs[242]);
    assign layer0_outputs[8414] = (inputs[112]) & ~(inputs[249]);
    assign layer0_outputs[8415] = (inputs[78]) ^ (inputs[149]);
    assign layer0_outputs[8416] = ~(inputs[182]);
    assign layer0_outputs[8417] = (inputs[159]) & ~(inputs[67]);
    assign layer0_outputs[8418] = ~(inputs[13]);
    assign layer0_outputs[8419] = 1'b0;
    assign layer0_outputs[8420] = ~(inputs[214]) | (inputs[33]);
    assign layer0_outputs[8421] = (inputs[20]) & ~(inputs[88]);
    assign layer0_outputs[8422] = inputs[192];
    assign layer0_outputs[8423] = (inputs[116]) ^ (inputs[200]);
    assign layer0_outputs[8424] = ~(inputs[53]) | (inputs[240]);
    assign layer0_outputs[8425] = ~(inputs[13]);
    assign layer0_outputs[8426] = ~(inputs[148]);
    assign layer0_outputs[8427] = (inputs[61]) & ~(inputs[190]);
    assign layer0_outputs[8428] = (inputs[26]) & ~(inputs[250]);
    assign layer0_outputs[8429] = ~((inputs[38]) ^ (inputs[250]));
    assign layer0_outputs[8430] = (inputs[135]) & ~(inputs[18]);
    assign layer0_outputs[8431] = ~(inputs[154]) | (inputs[192]);
    assign layer0_outputs[8432] = ~((inputs[59]) ^ (inputs[168]));
    assign layer0_outputs[8433] = ~((inputs[47]) | (inputs[193]));
    assign layer0_outputs[8434] = ~(inputs[228]) | (inputs[109]);
    assign layer0_outputs[8435] = (inputs[151]) & (inputs[250]);
    assign layer0_outputs[8436] = ~(inputs[58]) | (inputs[184]);
    assign layer0_outputs[8437] = 1'b0;
    assign layer0_outputs[8438] = ~((inputs[157]) ^ (inputs[15]));
    assign layer0_outputs[8439] = ~(inputs[161]) | (inputs[94]);
    assign layer0_outputs[8440] = ~((inputs[249]) ^ (inputs[126]));
    assign layer0_outputs[8441] = ~(inputs[221]);
    assign layer0_outputs[8442] = (inputs[84]) ^ (inputs[112]);
    assign layer0_outputs[8443] = (inputs[24]) & ~(inputs[255]);
    assign layer0_outputs[8444] = ~((inputs[4]) | (inputs[147]));
    assign layer0_outputs[8445] = (inputs[31]) | (inputs[52]);
    assign layer0_outputs[8446] = ~((inputs[141]) | (inputs[179]));
    assign layer0_outputs[8447] = inputs[38];
    assign layer0_outputs[8448] = ~(inputs[237]);
    assign layer0_outputs[8449] = inputs[153];
    assign layer0_outputs[8450] = ~((inputs[234]) | (inputs[201]));
    assign layer0_outputs[8451] = ~(inputs[121]);
    assign layer0_outputs[8452] = 1'b1;
    assign layer0_outputs[8453] = (inputs[131]) ^ (inputs[102]);
    assign layer0_outputs[8454] = inputs[132];
    assign layer0_outputs[8455] = (inputs[239]) | (inputs[181]);
    assign layer0_outputs[8456] = inputs[230];
    assign layer0_outputs[8457] = ~(inputs[59]);
    assign layer0_outputs[8458] = ~((inputs[209]) & (inputs[193]));
    assign layer0_outputs[8459] = (inputs[110]) ^ (inputs[61]);
    assign layer0_outputs[8460] = inputs[230];
    assign layer0_outputs[8461] = (inputs[11]) | (inputs[196]);
    assign layer0_outputs[8462] = ~(inputs[29]);
    assign layer0_outputs[8463] = ~(inputs[189]) | (inputs[184]);
    assign layer0_outputs[8464] = ~(inputs[7]);
    assign layer0_outputs[8465] = ~(inputs[116]);
    assign layer0_outputs[8466] = ~(inputs[113]);
    assign layer0_outputs[8467] = (inputs[173]) & ~(inputs[83]);
    assign layer0_outputs[8468] = inputs[136];
    assign layer0_outputs[8469] = (inputs[204]) & ~(inputs[65]);
    assign layer0_outputs[8470] = (inputs[149]) ^ (inputs[241]);
    assign layer0_outputs[8471] = inputs[55];
    assign layer0_outputs[8472] = (inputs[179]) | (inputs[237]);
    assign layer0_outputs[8473] = (inputs[215]) & ~(inputs[132]);
    assign layer0_outputs[8474] = inputs[203];
    assign layer0_outputs[8475] = ~(inputs[147]) | (inputs[142]);
    assign layer0_outputs[8476] = ~(inputs[166]) | (inputs[209]);
    assign layer0_outputs[8477] = ~(inputs[140]) | (inputs[178]);
    assign layer0_outputs[8478] = ~((inputs[60]) | (inputs[37]));
    assign layer0_outputs[8479] = ~(inputs[81]) | (inputs[169]);
    assign layer0_outputs[8480] = (inputs[235]) & ~(inputs[100]);
    assign layer0_outputs[8481] = ~(inputs[141]);
    assign layer0_outputs[8482] = inputs[146];
    assign layer0_outputs[8483] = (inputs[199]) & ~(inputs[40]);
    assign layer0_outputs[8484] = (inputs[128]) ^ (inputs[246]);
    assign layer0_outputs[8485] = inputs[222];
    assign layer0_outputs[8486] = (inputs[75]) & ~(inputs[209]);
    assign layer0_outputs[8487] = 1'b0;
    assign layer0_outputs[8488] = ~(inputs[183]) | (inputs[208]);
    assign layer0_outputs[8489] = (inputs[239]) | (inputs[228]);
    assign layer0_outputs[8490] = 1'b1;
    assign layer0_outputs[8491] = ~(inputs[40]);
    assign layer0_outputs[8492] = ~((inputs[208]) | (inputs[244]));
    assign layer0_outputs[8493] = ~(inputs[10]);
    assign layer0_outputs[8494] = (inputs[207]) | (inputs[167]);
    assign layer0_outputs[8495] = ~(inputs[223]);
    assign layer0_outputs[8496] = ~((inputs[204]) ^ (inputs[147]));
    assign layer0_outputs[8497] = ~((inputs[204]) & (inputs[39]));
    assign layer0_outputs[8498] = ~(inputs[148]);
    assign layer0_outputs[8499] = (inputs[174]) & ~(inputs[237]);
    assign layer0_outputs[8500] = (inputs[117]) & ~(inputs[251]);
    assign layer0_outputs[8501] = ~(inputs[126]);
    assign layer0_outputs[8502] = ~(inputs[227]);
    assign layer0_outputs[8503] = (inputs[11]) | (inputs[82]);
    assign layer0_outputs[8504] = ~(inputs[100]) | (inputs[223]);
    assign layer0_outputs[8505] = ~((inputs[253]) | (inputs[182]));
    assign layer0_outputs[8506] = ~(inputs[22]);
    assign layer0_outputs[8507] = (inputs[240]) | (inputs[188]);
    assign layer0_outputs[8508] = ~((inputs[61]) ^ (inputs[63]));
    assign layer0_outputs[8509] = (inputs[47]) ^ (inputs[3]);
    assign layer0_outputs[8510] = inputs[110];
    assign layer0_outputs[8511] = ~((inputs[253]) ^ (inputs[52]));
    assign layer0_outputs[8512] = ~((inputs[38]) | (inputs[62]));
    assign layer0_outputs[8513] = (inputs[143]) & ~(inputs[194]);
    assign layer0_outputs[8514] = (inputs[12]) & ~(inputs[221]);
    assign layer0_outputs[8515] = inputs[230];
    assign layer0_outputs[8516] = (inputs[97]) | (inputs[254]);
    assign layer0_outputs[8517] = ~((inputs[170]) | (inputs[230]));
    assign layer0_outputs[8518] = inputs[111];
    assign layer0_outputs[8519] = (inputs[147]) ^ (inputs[184]);
    assign layer0_outputs[8520] = (inputs[46]) | (inputs[232]);
    assign layer0_outputs[8521] = (inputs[151]) | (inputs[77]);
    assign layer0_outputs[8522] = (inputs[72]) & ~(inputs[62]);
    assign layer0_outputs[8523] = inputs[115];
    assign layer0_outputs[8524] = ~((inputs[5]) & (inputs[178]));
    assign layer0_outputs[8525] = ~(inputs[51]) | (inputs[145]);
    assign layer0_outputs[8526] = (inputs[18]) | (inputs[185]);
    assign layer0_outputs[8527] = ~(inputs[100]);
    assign layer0_outputs[8528] = ~(inputs[221]) | (inputs[94]);
    assign layer0_outputs[8529] = ~((inputs[72]) | (inputs[249]));
    assign layer0_outputs[8530] = (inputs[39]) & ~(inputs[173]);
    assign layer0_outputs[8531] = (inputs[100]) | (inputs[249]);
    assign layer0_outputs[8532] = 1'b1;
    assign layer0_outputs[8533] = (inputs[121]) ^ (inputs[251]);
    assign layer0_outputs[8534] = ~(inputs[30]);
    assign layer0_outputs[8535] = ~((inputs[56]) | (inputs[210]));
    assign layer0_outputs[8536] = (inputs[13]) & ~(inputs[239]);
    assign layer0_outputs[8537] = (inputs[8]) ^ (inputs[189]);
    assign layer0_outputs[8538] = (inputs[118]) ^ (inputs[149]);
    assign layer0_outputs[8539] = (inputs[143]) & ~(inputs[239]);
    assign layer0_outputs[8540] = ~((inputs[100]) | (inputs[113]));
    assign layer0_outputs[8541] = ~(inputs[78]);
    assign layer0_outputs[8542] = inputs[193];
    assign layer0_outputs[8543] = ~((inputs[194]) | (inputs[198]));
    assign layer0_outputs[8544] = (inputs[188]) ^ (inputs[136]);
    assign layer0_outputs[8545] = (inputs[100]) ^ (inputs[126]);
    assign layer0_outputs[8546] = (inputs[161]) ^ (inputs[152]);
    assign layer0_outputs[8547] = inputs[26];
    assign layer0_outputs[8548] = (inputs[55]) & ~(inputs[35]);
    assign layer0_outputs[8549] = (inputs[31]) ^ (inputs[67]);
    assign layer0_outputs[8550] = ~((inputs[94]) & (inputs[130]));
    assign layer0_outputs[8551] = (inputs[198]) & ~(inputs[42]);
    assign layer0_outputs[8552] = (inputs[36]) | (inputs[50]);
    assign layer0_outputs[8553] = inputs[130];
    assign layer0_outputs[8554] = (inputs[100]) ^ (inputs[72]);
    assign layer0_outputs[8555] = (inputs[60]) ^ (inputs[143]);
    assign layer0_outputs[8556] = inputs[215];
    assign layer0_outputs[8557] = ~(inputs[254]);
    assign layer0_outputs[8558] = inputs[121];
    assign layer0_outputs[8559] = ~(inputs[95]) | (inputs[129]);
    assign layer0_outputs[8560] = ~(inputs[213]);
    assign layer0_outputs[8561] = (inputs[250]) | (inputs[210]);
    assign layer0_outputs[8562] = ~(inputs[80]);
    assign layer0_outputs[8563] = inputs[17];
    assign layer0_outputs[8564] = (inputs[157]) & ~(inputs[61]);
    assign layer0_outputs[8565] = inputs[215];
    assign layer0_outputs[8566] = 1'b0;
    assign layer0_outputs[8567] = inputs[53];
    assign layer0_outputs[8568] = ~((inputs[202]) | (inputs[218]));
    assign layer0_outputs[8569] = (inputs[48]) & ~(inputs[12]);
    assign layer0_outputs[8570] = 1'b0;
    assign layer0_outputs[8571] = inputs[24];
    assign layer0_outputs[8572] = ~(inputs[168]) | (inputs[34]);
    assign layer0_outputs[8573] = ~((inputs[78]) ^ (inputs[248]));
    assign layer0_outputs[8574] = (inputs[18]) & ~(inputs[199]);
    assign layer0_outputs[8575] = inputs[235];
    assign layer0_outputs[8576] = inputs[211];
    assign layer0_outputs[8577] = ~(inputs[142]) | (inputs[220]);
    assign layer0_outputs[8578] = (inputs[153]) & ~(inputs[38]);
    assign layer0_outputs[8579] = ~((inputs[237]) & (inputs[218]));
    assign layer0_outputs[8580] = ~((inputs[252]) | (inputs[177]));
    assign layer0_outputs[8581] = ~((inputs[119]) | (inputs[121]));
    assign layer0_outputs[8582] = (inputs[211]) | (inputs[84]);
    assign layer0_outputs[8583] = ~((inputs[218]) ^ (inputs[115]));
    assign layer0_outputs[8584] = ~((inputs[27]) ^ (inputs[233]));
    assign layer0_outputs[8585] = (inputs[56]) & ~(inputs[18]);
    assign layer0_outputs[8586] = ~((inputs[230]) | (inputs[223]));
    assign layer0_outputs[8587] = ~(inputs[99]);
    assign layer0_outputs[8588] = inputs[196];
    assign layer0_outputs[8589] = ~((inputs[103]) & (inputs[89]));
    assign layer0_outputs[8590] = inputs[81];
    assign layer0_outputs[8591] = ~((inputs[76]) ^ (inputs[109]));
    assign layer0_outputs[8592] = ~(inputs[120]);
    assign layer0_outputs[8593] = ~((inputs[152]) & (inputs[86]));
    assign layer0_outputs[8594] = ~(inputs[212]) | (inputs[76]);
    assign layer0_outputs[8595] = (inputs[176]) ^ (inputs[138]);
    assign layer0_outputs[8596] = (inputs[133]) & ~(inputs[13]);
    assign layer0_outputs[8597] = ~((inputs[192]) | (inputs[216]));
    assign layer0_outputs[8598] = ~(inputs[132]);
    assign layer0_outputs[8599] = (inputs[2]) | (inputs[156]);
    assign layer0_outputs[8600] = (inputs[186]) | (inputs[163]);
    assign layer0_outputs[8601] = ~(inputs[61]);
    assign layer0_outputs[8602] = (inputs[250]) & ~(inputs[75]);
    assign layer0_outputs[8603] = ~((inputs[214]) | (inputs[188]));
    assign layer0_outputs[8604] = inputs[209];
    assign layer0_outputs[8605] = ~((inputs[59]) ^ (inputs[131]));
    assign layer0_outputs[8606] = (inputs[108]) | (inputs[253]);
    assign layer0_outputs[8607] = ~(inputs[137]) | (inputs[102]);
    assign layer0_outputs[8608] = ~((inputs[222]) | (inputs[5]));
    assign layer0_outputs[8609] = ~(inputs[187]) | (inputs[223]);
    assign layer0_outputs[8610] = (inputs[178]) ^ (inputs[249]);
    assign layer0_outputs[8611] = ~((inputs[146]) ^ (inputs[70]));
    assign layer0_outputs[8612] = ~((inputs[68]) | (inputs[114]));
    assign layer0_outputs[8613] = (inputs[186]) & (inputs[48]);
    assign layer0_outputs[8614] = (inputs[191]) & ~(inputs[14]);
    assign layer0_outputs[8615] = (inputs[25]) & ~(inputs[159]);
    assign layer0_outputs[8616] = (inputs[213]) ^ (inputs[122]);
    assign layer0_outputs[8617] = ~(inputs[151]);
    assign layer0_outputs[8618] = (inputs[131]) & ~(inputs[35]);
    assign layer0_outputs[8619] = (inputs[7]) ^ (inputs[69]);
    assign layer0_outputs[8620] = ~((inputs[212]) & (inputs[215]));
    assign layer0_outputs[8621] = ~((inputs[3]) ^ (inputs[139]));
    assign layer0_outputs[8622] = (inputs[229]) & ~(inputs[143]);
    assign layer0_outputs[8623] = ~((inputs[71]) | (inputs[227]));
    assign layer0_outputs[8624] = ~((inputs[177]) | (inputs[11]));
    assign layer0_outputs[8625] = inputs[184];
    assign layer0_outputs[8626] = ~(inputs[153]);
    assign layer0_outputs[8627] = (inputs[134]) ^ (inputs[87]);
    assign layer0_outputs[8628] = (inputs[98]) & (inputs[134]);
    assign layer0_outputs[8629] = ~(inputs[64]);
    assign layer0_outputs[8630] = inputs[130];
    assign layer0_outputs[8631] = ~(inputs[198]);
    assign layer0_outputs[8632] = ~((inputs[188]) | (inputs[75]));
    assign layer0_outputs[8633] = ~(inputs[182]) | (inputs[97]);
    assign layer0_outputs[8634] = ~(inputs[148]);
    assign layer0_outputs[8635] = inputs[164];
    assign layer0_outputs[8636] = (inputs[237]) | (inputs[145]);
    assign layer0_outputs[8637] = ~((inputs[199]) | (inputs[8]));
    assign layer0_outputs[8638] = inputs[46];
    assign layer0_outputs[8639] = inputs[193];
    assign layer0_outputs[8640] = (inputs[191]) | (inputs[189]);
    assign layer0_outputs[8641] = (inputs[103]) & ~(inputs[163]);
    assign layer0_outputs[8642] = (inputs[64]) & ~(inputs[112]);
    assign layer0_outputs[8643] = ~((inputs[17]) | (inputs[182]));
    assign layer0_outputs[8644] = 1'b0;
    assign layer0_outputs[8645] = (inputs[119]) ^ (inputs[106]);
    assign layer0_outputs[8646] = ~(inputs[128]);
    assign layer0_outputs[8647] = ~((inputs[194]) ^ (inputs[247]));
    assign layer0_outputs[8648] = (inputs[179]) | (inputs[87]);
    assign layer0_outputs[8649] = inputs[22];
    assign layer0_outputs[8650] = ~((inputs[26]) ^ (inputs[64]));
    assign layer0_outputs[8651] = ~((inputs[227]) | (inputs[132]));
    assign layer0_outputs[8652] = inputs[18];
    assign layer0_outputs[8653] = inputs[45];
    assign layer0_outputs[8654] = (inputs[55]) & (inputs[49]);
    assign layer0_outputs[8655] = ~((inputs[202]) | (inputs[233]));
    assign layer0_outputs[8656] = inputs[207];
    assign layer0_outputs[8657] = (inputs[230]) & ~(inputs[56]);
    assign layer0_outputs[8658] = ~(inputs[139]) | (inputs[163]);
    assign layer0_outputs[8659] = (inputs[184]) & ~(inputs[163]);
    assign layer0_outputs[8660] = ~((inputs[207]) ^ (inputs[19]));
    assign layer0_outputs[8661] = inputs[168];
    assign layer0_outputs[8662] = inputs[197];
    assign layer0_outputs[8663] = ~((inputs[240]) ^ (inputs[213]));
    assign layer0_outputs[8664] = (inputs[233]) & ~(inputs[96]);
    assign layer0_outputs[8665] = ~(inputs[118]);
    assign layer0_outputs[8666] = inputs[187];
    assign layer0_outputs[8667] = ~(inputs[253]);
    assign layer0_outputs[8668] = ~(inputs[85]);
    assign layer0_outputs[8669] = (inputs[247]) & ~(inputs[177]);
    assign layer0_outputs[8670] = (inputs[72]) ^ (inputs[46]);
    assign layer0_outputs[8671] = ~(inputs[8]) | (inputs[249]);
    assign layer0_outputs[8672] = (inputs[186]) & ~(inputs[110]);
    assign layer0_outputs[8673] = inputs[211];
    assign layer0_outputs[8674] = (inputs[110]) | (inputs[253]);
    assign layer0_outputs[8675] = inputs[205];
    assign layer0_outputs[8676] = ~(inputs[105]) | (inputs[209]);
    assign layer0_outputs[8677] = (inputs[226]) ^ (inputs[181]);
    assign layer0_outputs[8678] = (inputs[36]) | (inputs[255]);
    assign layer0_outputs[8679] = ~((inputs[75]) | (inputs[154]));
    assign layer0_outputs[8680] = ~(inputs[51]);
    assign layer0_outputs[8681] = ~(inputs[22]);
    assign layer0_outputs[8682] = 1'b1;
    assign layer0_outputs[8683] = inputs[203];
    assign layer0_outputs[8684] = (inputs[174]) | (inputs[245]);
    assign layer0_outputs[8685] = ~(inputs[230]);
    assign layer0_outputs[8686] = ~(inputs[207]);
    assign layer0_outputs[8687] = (inputs[42]) | (inputs[155]);
    assign layer0_outputs[8688] = inputs[85];
    assign layer0_outputs[8689] = ~(inputs[150]);
    assign layer0_outputs[8690] = 1'b1;
    assign layer0_outputs[8691] = ~((inputs[187]) ^ (inputs[183]));
    assign layer0_outputs[8692] = ~((inputs[80]) | (inputs[64]));
    assign layer0_outputs[8693] = ~((inputs[187]) | (inputs[98]));
    assign layer0_outputs[8694] = (inputs[145]) & ~(inputs[79]);
    assign layer0_outputs[8695] = ~(inputs[247]);
    assign layer0_outputs[8696] = inputs[71];
    assign layer0_outputs[8697] = ~((inputs[139]) | (inputs[45]));
    assign layer0_outputs[8698] = inputs[167];
    assign layer0_outputs[8699] = (inputs[96]) | (inputs[150]);
    assign layer0_outputs[8700] = ~(inputs[87]) | (inputs[49]);
    assign layer0_outputs[8701] = (inputs[178]) | (inputs[252]);
    assign layer0_outputs[8702] = ~((inputs[66]) ^ (inputs[25]));
    assign layer0_outputs[8703] = ~((inputs[96]) | (inputs[129]));
    assign layer0_outputs[8704] = ~(inputs[99]);
    assign layer0_outputs[8705] = inputs[162];
    assign layer0_outputs[8706] = inputs[177];
    assign layer0_outputs[8707] = ~(inputs[200]);
    assign layer0_outputs[8708] = (inputs[93]) & ~(inputs[17]);
    assign layer0_outputs[8709] = (inputs[118]) & ~(inputs[133]);
    assign layer0_outputs[8710] = (inputs[71]) & ~(inputs[246]);
    assign layer0_outputs[8711] = ~(inputs[4]);
    assign layer0_outputs[8712] = ~((inputs[124]) & (inputs[44]));
    assign layer0_outputs[8713] = ~((inputs[33]) | (inputs[192]));
    assign layer0_outputs[8714] = (inputs[228]) | (inputs[10]);
    assign layer0_outputs[8715] = ~(inputs[114]);
    assign layer0_outputs[8716] = ~((inputs[157]) ^ (inputs[4]));
    assign layer0_outputs[8717] = ~((inputs[1]) | (inputs[180]));
    assign layer0_outputs[8718] = ~(inputs[40]);
    assign layer0_outputs[8719] = inputs[67];
    assign layer0_outputs[8720] = ~(inputs[20]);
    assign layer0_outputs[8721] = (inputs[228]) | (inputs[230]);
    assign layer0_outputs[8722] = ~(inputs[179]);
    assign layer0_outputs[8723] = ~(inputs[145]);
    assign layer0_outputs[8724] = (inputs[146]) | (inputs[105]);
    assign layer0_outputs[8725] = ~(inputs[18]) | (inputs[14]);
    assign layer0_outputs[8726] = inputs[103];
    assign layer0_outputs[8727] = (inputs[220]) | (inputs[197]);
    assign layer0_outputs[8728] = ~((inputs[189]) & (inputs[122]));
    assign layer0_outputs[8729] = ~((inputs[104]) | (inputs[192]));
    assign layer0_outputs[8730] = (inputs[198]) ^ (inputs[175]);
    assign layer0_outputs[8731] = inputs[43];
    assign layer0_outputs[8732] = ~(inputs[11]);
    assign layer0_outputs[8733] = ~(inputs[156]);
    assign layer0_outputs[8734] = inputs[204];
    assign layer0_outputs[8735] = inputs[188];
    assign layer0_outputs[8736] = (inputs[36]) | (inputs[32]);
    assign layer0_outputs[8737] = ~((inputs[96]) ^ (inputs[83]));
    assign layer0_outputs[8738] = ~(inputs[132]);
    assign layer0_outputs[8739] = (inputs[251]) | (inputs[88]);
    assign layer0_outputs[8740] = inputs[111];
    assign layer0_outputs[8741] = (inputs[28]) & ~(inputs[160]);
    assign layer0_outputs[8742] = inputs[83];
    assign layer0_outputs[8743] = ~(inputs[91]) | (inputs[23]);
    assign layer0_outputs[8744] = (inputs[96]) ^ (inputs[209]);
    assign layer0_outputs[8745] = ~(inputs[202]) | (inputs[59]);
    assign layer0_outputs[8746] = ~((inputs[114]) | (inputs[58]));
    assign layer0_outputs[8747] = (inputs[146]) ^ (inputs[104]);
    assign layer0_outputs[8748] = ~(inputs[230]);
    assign layer0_outputs[8749] = (inputs[203]) & ~(inputs[47]);
    assign layer0_outputs[8750] = (inputs[162]) | (inputs[94]);
    assign layer0_outputs[8751] = ~(inputs[105]);
    assign layer0_outputs[8752] = ~(inputs[152]);
    assign layer0_outputs[8753] = ~(inputs[206]);
    assign layer0_outputs[8754] = ~((inputs[64]) | (inputs[182]));
    assign layer0_outputs[8755] = ~(inputs[173]) | (inputs[158]);
    assign layer0_outputs[8756] = (inputs[0]) | (inputs[247]);
    assign layer0_outputs[8757] = ~((inputs[163]) | (inputs[247]));
    assign layer0_outputs[8758] = (inputs[176]) ^ (inputs[45]);
    assign layer0_outputs[8759] = ~(inputs[25]);
    assign layer0_outputs[8760] = (inputs[185]) ^ (inputs[138]);
    assign layer0_outputs[8761] = (inputs[162]) | (inputs[91]);
    assign layer0_outputs[8762] = ~(inputs[176]);
    assign layer0_outputs[8763] = ~(inputs[246]) | (inputs[126]);
    assign layer0_outputs[8764] = inputs[78];
    assign layer0_outputs[8765] = 1'b1;
    assign layer0_outputs[8766] = inputs[176];
    assign layer0_outputs[8767] = (inputs[224]) & ~(inputs[214]);
    assign layer0_outputs[8768] = ~(inputs[117]);
    assign layer0_outputs[8769] = ~((inputs[91]) | (inputs[240]));
    assign layer0_outputs[8770] = ~(inputs[94]) | (inputs[35]);
    assign layer0_outputs[8771] = ~(inputs[86]);
    assign layer0_outputs[8772] = (inputs[207]) ^ (inputs[142]);
    assign layer0_outputs[8773] = (inputs[233]) & ~(inputs[46]);
    assign layer0_outputs[8774] = ~((inputs[217]) & (inputs[204]));
    assign layer0_outputs[8775] = ~(inputs[59]);
    assign layer0_outputs[8776] = ~(inputs[48]);
    assign layer0_outputs[8777] = ~(inputs[197]) | (inputs[78]);
    assign layer0_outputs[8778] = 1'b0;
    assign layer0_outputs[8779] = (inputs[155]) & ~(inputs[42]);
    assign layer0_outputs[8780] = (inputs[165]) | (inputs[248]);
    assign layer0_outputs[8781] = (inputs[165]) & ~(inputs[59]);
    assign layer0_outputs[8782] = ~(inputs[167]) | (inputs[47]);
    assign layer0_outputs[8783] = (inputs[254]) | (inputs[255]);
    assign layer0_outputs[8784] = (inputs[48]) | (inputs[234]);
    assign layer0_outputs[8785] = (inputs[35]) & ~(inputs[173]);
    assign layer0_outputs[8786] = ~((inputs[163]) | (inputs[134]));
    assign layer0_outputs[8787] = (inputs[92]) ^ (inputs[19]);
    assign layer0_outputs[8788] = ~(inputs[44]);
    assign layer0_outputs[8789] = 1'b0;
    assign layer0_outputs[8790] = (inputs[38]) ^ (inputs[193]);
    assign layer0_outputs[8791] = ~(inputs[32]);
    assign layer0_outputs[8792] = ~((inputs[201]) | (inputs[249]));
    assign layer0_outputs[8793] = inputs[30];
    assign layer0_outputs[8794] = inputs[231];
    assign layer0_outputs[8795] = ~(inputs[133]);
    assign layer0_outputs[8796] = (inputs[148]) & ~(inputs[130]);
    assign layer0_outputs[8797] = (inputs[124]) | (inputs[111]);
    assign layer0_outputs[8798] = (inputs[236]) & (inputs[17]);
    assign layer0_outputs[8799] = (inputs[149]) & ~(inputs[2]);
    assign layer0_outputs[8800] = ~(inputs[232]);
    assign layer0_outputs[8801] = ~((inputs[53]) ^ (inputs[59]));
    assign layer0_outputs[8802] = (inputs[210]) | (inputs[145]);
    assign layer0_outputs[8803] = ~(inputs[88]);
    assign layer0_outputs[8804] = (inputs[198]) | (inputs[149]);
    assign layer0_outputs[8805] = 1'b1;
    assign layer0_outputs[8806] = (inputs[14]) & ~(inputs[5]);
    assign layer0_outputs[8807] = ~(inputs[132]) | (inputs[201]);
    assign layer0_outputs[8808] = (inputs[167]) & ~(inputs[143]);
    assign layer0_outputs[8809] = (inputs[176]) | (inputs[247]);
    assign layer0_outputs[8810] = 1'b1;
    assign layer0_outputs[8811] = ~(inputs[136]);
    assign layer0_outputs[8812] = ~((inputs[73]) ^ (inputs[96]));
    assign layer0_outputs[8813] = (inputs[211]) & ~(inputs[68]);
    assign layer0_outputs[8814] = (inputs[52]) | (inputs[95]);
    assign layer0_outputs[8815] = ~((inputs[145]) | (inputs[171]));
    assign layer0_outputs[8816] = ~(inputs[173]) | (inputs[111]);
    assign layer0_outputs[8817] = 1'b0;
    assign layer0_outputs[8818] = ~((inputs[73]) & (inputs[184]));
    assign layer0_outputs[8819] = ~(inputs[207]);
    assign layer0_outputs[8820] = ~(inputs[165]) | (inputs[192]);
    assign layer0_outputs[8821] = inputs[108];
    assign layer0_outputs[8822] = (inputs[91]) | (inputs[108]);
    assign layer0_outputs[8823] = ~(inputs[74]) | (inputs[145]);
    assign layer0_outputs[8824] = ~(inputs[213]);
    assign layer0_outputs[8825] = (inputs[204]) ^ (inputs[67]);
    assign layer0_outputs[8826] = ~(inputs[245]);
    assign layer0_outputs[8827] = (inputs[86]) | (inputs[91]);
    assign layer0_outputs[8828] = ~((inputs[64]) ^ (inputs[240]));
    assign layer0_outputs[8829] = ~(inputs[14]);
    assign layer0_outputs[8830] = (inputs[248]) | (inputs[157]);
    assign layer0_outputs[8831] = ~(inputs[86]);
    assign layer0_outputs[8832] = ~(inputs[20]);
    assign layer0_outputs[8833] = inputs[240];
    assign layer0_outputs[8834] = ~(inputs[116]) | (inputs[208]);
    assign layer0_outputs[8835] = (inputs[118]) ^ (inputs[51]);
    assign layer0_outputs[8836] = ~((inputs[40]) | (inputs[14]));
    assign layer0_outputs[8837] = ~((inputs[232]) ^ (inputs[70]));
    assign layer0_outputs[8838] = (inputs[135]) & ~(inputs[160]);
    assign layer0_outputs[8839] = (inputs[210]) & ~(inputs[130]);
    assign layer0_outputs[8840] = (inputs[125]) & ~(inputs[254]);
    assign layer0_outputs[8841] = ~(inputs[110]);
    assign layer0_outputs[8842] = ~(inputs[232]);
    assign layer0_outputs[8843] = ~((inputs[145]) | (inputs[42]));
    assign layer0_outputs[8844] = ~((inputs[110]) ^ (inputs[32]));
    assign layer0_outputs[8845] = ~((inputs[90]) ^ (inputs[34]));
    assign layer0_outputs[8846] = ~(inputs[212]);
    assign layer0_outputs[8847] = ~(inputs[6]);
    assign layer0_outputs[8848] = inputs[56];
    assign layer0_outputs[8849] = ~(inputs[141]) | (inputs[157]);
    assign layer0_outputs[8850] = ~(inputs[177]) | (inputs[32]);
    assign layer0_outputs[8851] = (inputs[248]) & ~(inputs[168]);
    assign layer0_outputs[8852] = (inputs[3]) ^ (inputs[33]);
    assign layer0_outputs[8853] = ~((inputs[197]) ^ (inputs[242]));
    assign layer0_outputs[8854] = ~((inputs[97]) | (inputs[192]));
    assign layer0_outputs[8855] = ~(inputs[87]) | (inputs[244]);
    assign layer0_outputs[8856] = ~(inputs[4]);
    assign layer0_outputs[8857] = (inputs[135]) | (inputs[236]);
    assign layer0_outputs[8858] = ~(inputs[217]);
    assign layer0_outputs[8859] = ~(inputs[116]);
    assign layer0_outputs[8860] = ~(inputs[60]);
    assign layer0_outputs[8861] = inputs[193];
    assign layer0_outputs[8862] = inputs[114];
    assign layer0_outputs[8863] = inputs[67];
    assign layer0_outputs[8864] = inputs[108];
    assign layer0_outputs[8865] = (inputs[187]) & ~(inputs[28]);
    assign layer0_outputs[8866] = ~(inputs[253]);
    assign layer0_outputs[8867] = ~(inputs[169]) | (inputs[226]);
    assign layer0_outputs[8868] = ~(inputs[161]) | (inputs[2]);
    assign layer0_outputs[8869] = ~((inputs[188]) | (inputs[189]));
    assign layer0_outputs[8870] = 1'b1;
    assign layer0_outputs[8871] = inputs[117];
    assign layer0_outputs[8872] = inputs[163];
    assign layer0_outputs[8873] = ~(inputs[21]) | (inputs[114]);
    assign layer0_outputs[8874] = ~(inputs[230]);
    assign layer0_outputs[8875] = ~((inputs[187]) | (inputs[111]));
    assign layer0_outputs[8876] = ~(inputs[125]);
    assign layer0_outputs[8877] = ~(inputs[152]) | (inputs[64]);
    assign layer0_outputs[8878] = ~(inputs[102]);
    assign layer0_outputs[8879] = inputs[212];
    assign layer0_outputs[8880] = (inputs[99]) & ~(inputs[250]);
    assign layer0_outputs[8881] = inputs[93];
    assign layer0_outputs[8882] = ~((inputs[115]) ^ (inputs[203]));
    assign layer0_outputs[8883] = ~(inputs[94]);
    assign layer0_outputs[8884] = ~((inputs[106]) ^ (inputs[97]));
    assign layer0_outputs[8885] = ~(inputs[93]);
    assign layer0_outputs[8886] = ~(inputs[34]) | (inputs[145]);
    assign layer0_outputs[8887] = ~((inputs[171]) ^ (inputs[159]));
    assign layer0_outputs[8888] = ~((inputs[119]) & (inputs[178]));
    assign layer0_outputs[8889] = ~((inputs[250]) | (inputs[204]));
    assign layer0_outputs[8890] = ~((inputs[249]) | (inputs[206]));
    assign layer0_outputs[8891] = (inputs[207]) & ~(inputs[97]);
    assign layer0_outputs[8892] = (inputs[145]) | (inputs[229]);
    assign layer0_outputs[8893] = ~(inputs[210]);
    assign layer0_outputs[8894] = ~((inputs[147]) | (inputs[226]));
    assign layer0_outputs[8895] = ~(inputs[81]);
    assign layer0_outputs[8896] = ~(inputs[184]);
    assign layer0_outputs[8897] = ~(inputs[88]) | (inputs[110]);
    assign layer0_outputs[8898] = inputs[57];
    assign layer0_outputs[8899] = inputs[43];
    assign layer0_outputs[8900] = (inputs[64]) | (inputs[222]);
    assign layer0_outputs[8901] = ~((inputs[176]) | (inputs[41]));
    assign layer0_outputs[8902] = ~(inputs[228]) | (inputs[8]);
    assign layer0_outputs[8903] = (inputs[9]) ^ (inputs[63]);
    assign layer0_outputs[8904] = ~((inputs[169]) & (inputs[136]));
    assign layer0_outputs[8905] = ~(inputs[244]) | (inputs[103]);
    assign layer0_outputs[8906] = inputs[110];
    assign layer0_outputs[8907] = (inputs[122]) ^ (inputs[156]);
    assign layer0_outputs[8908] = ~(inputs[218]) | (inputs[90]);
    assign layer0_outputs[8909] = inputs[133];
    assign layer0_outputs[8910] = ~(inputs[93]);
    assign layer0_outputs[8911] = inputs[114];
    assign layer0_outputs[8912] = (inputs[50]) | (inputs[127]);
    assign layer0_outputs[8913] = (inputs[145]) ^ (inputs[116]);
    assign layer0_outputs[8914] = ~((inputs[240]) & (inputs[191]));
    assign layer0_outputs[8915] = ~((inputs[190]) ^ (inputs[10]));
    assign layer0_outputs[8916] = (inputs[200]) ^ (inputs[16]);
    assign layer0_outputs[8917] = ~((inputs[75]) | (inputs[159]));
    assign layer0_outputs[8918] = inputs[147];
    assign layer0_outputs[8919] = ~(inputs[217]) | (inputs[74]);
    assign layer0_outputs[8920] = (inputs[0]) ^ (inputs[193]);
    assign layer0_outputs[8921] = ~(inputs[152]);
    assign layer0_outputs[8922] = (inputs[169]) | (inputs[168]);
    assign layer0_outputs[8923] = ~((inputs[128]) | (inputs[122]));
    assign layer0_outputs[8924] = ~((inputs[40]) ^ (inputs[130]));
    assign layer0_outputs[8925] = inputs[191];
    assign layer0_outputs[8926] = ~(inputs[250]);
    assign layer0_outputs[8927] = (inputs[197]) & ~(inputs[202]);
    assign layer0_outputs[8928] = ~(inputs[95]);
    assign layer0_outputs[8929] = (inputs[221]) & ~(inputs[110]);
    assign layer0_outputs[8930] = inputs[230];
    assign layer0_outputs[8931] = (inputs[229]) & ~(inputs[135]);
    assign layer0_outputs[8932] = ~(inputs[23]);
    assign layer0_outputs[8933] = inputs[84];
    assign layer0_outputs[8934] = inputs[248];
    assign layer0_outputs[8935] = (inputs[215]) & (inputs[115]);
    assign layer0_outputs[8936] = (inputs[84]) & ~(inputs[111]);
    assign layer0_outputs[8937] = ~((inputs[22]) | (inputs[10]));
    assign layer0_outputs[8938] = 1'b0;
    assign layer0_outputs[8939] = ~(inputs[180]) | (inputs[103]);
    assign layer0_outputs[8940] = inputs[131];
    assign layer0_outputs[8941] = ~(inputs[84]);
    assign layer0_outputs[8942] = ~((inputs[162]) ^ (inputs[189]));
    assign layer0_outputs[8943] = inputs[180];
    assign layer0_outputs[8944] = ~(inputs[199]) | (inputs[98]);
    assign layer0_outputs[8945] = ~(inputs[187]) | (inputs[147]);
    assign layer0_outputs[8946] = ~(inputs[0]) | (inputs[156]);
    assign layer0_outputs[8947] = inputs[214];
    assign layer0_outputs[8948] = inputs[114];
    assign layer0_outputs[8949] = ~(inputs[246]);
    assign layer0_outputs[8950] = (inputs[106]) & ~(inputs[195]);
    assign layer0_outputs[8951] = inputs[87];
    assign layer0_outputs[8952] = ~((inputs[11]) & (inputs[93]));
    assign layer0_outputs[8953] = inputs[98];
    assign layer0_outputs[8954] = ~((inputs[30]) & (inputs[56]));
    assign layer0_outputs[8955] = inputs[23];
    assign layer0_outputs[8956] = (inputs[180]) ^ (inputs[183]);
    assign layer0_outputs[8957] = inputs[125];
    assign layer0_outputs[8958] = (inputs[56]) & ~(inputs[6]);
    assign layer0_outputs[8959] = (inputs[83]) ^ (inputs[76]);
    assign layer0_outputs[8960] = (inputs[170]) | (inputs[129]);
    assign layer0_outputs[8961] = ~(inputs[249]);
    assign layer0_outputs[8962] = inputs[97];
    assign layer0_outputs[8963] = ~(inputs[54]) | (inputs[233]);
    assign layer0_outputs[8964] = inputs[234];
    assign layer0_outputs[8965] = (inputs[72]) & ~(inputs[34]);
    assign layer0_outputs[8966] = ~(inputs[146]);
    assign layer0_outputs[8967] = ~(inputs[158]);
    assign layer0_outputs[8968] = ~(inputs[231]);
    assign layer0_outputs[8969] = (inputs[155]) | (inputs[249]);
    assign layer0_outputs[8970] = (inputs[90]) | (inputs[76]);
    assign layer0_outputs[8971] = (inputs[157]) | (inputs[122]);
    assign layer0_outputs[8972] = ~(inputs[139]) | (inputs[145]);
    assign layer0_outputs[8973] = inputs[222];
    assign layer0_outputs[8974] = (inputs[57]) ^ (inputs[110]);
    assign layer0_outputs[8975] = (inputs[63]) | (inputs[58]);
    assign layer0_outputs[8976] = (inputs[123]) & ~(inputs[212]);
    assign layer0_outputs[8977] = ~(inputs[171]);
    assign layer0_outputs[8978] = (inputs[179]) & ~(inputs[96]);
    assign layer0_outputs[8979] = ~((inputs[190]) | (inputs[60]));
    assign layer0_outputs[8980] = (inputs[251]) | (inputs[63]);
    assign layer0_outputs[8981] = ~(inputs[90]);
    assign layer0_outputs[8982] = (inputs[72]) ^ (inputs[44]);
    assign layer0_outputs[8983] = 1'b1;
    assign layer0_outputs[8984] = ~(inputs[0]);
    assign layer0_outputs[8985] = (inputs[212]) | (inputs[81]);
    assign layer0_outputs[8986] = ~((inputs[84]) | (inputs[50]));
    assign layer0_outputs[8987] = (inputs[224]) & ~(inputs[241]);
    assign layer0_outputs[8988] = ~(inputs[103]);
    assign layer0_outputs[8989] = inputs[99];
    assign layer0_outputs[8990] = (inputs[117]) & ~(inputs[2]);
    assign layer0_outputs[8991] = (inputs[43]) & ~(inputs[161]);
    assign layer0_outputs[8992] = ~(inputs[66]);
    assign layer0_outputs[8993] = ~((inputs[32]) | (inputs[63]));
    assign layer0_outputs[8994] = ~(inputs[43]) | (inputs[220]);
    assign layer0_outputs[8995] = (inputs[246]) & ~(inputs[120]);
    assign layer0_outputs[8996] = (inputs[24]) & (inputs[106]);
    assign layer0_outputs[8997] = (inputs[221]) | (inputs[236]);
    assign layer0_outputs[8998] = (inputs[146]) | (inputs[176]);
    assign layer0_outputs[8999] = ~((inputs[118]) | (inputs[199]));
    assign layer0_outputs[9000] = ~(inputs[39]) | (inputs[246]);
    assign layer0_outputs[9001] = inputs[104];
    assign layer0_outputs[9002] = (inputs[67]) | (inputs[113]);
    assign layer0_outputs[9003] = ~((inputs[12]) ^ (inputs[100]));
    assign layer0_outputs[9004] = (inputs[94]) ^ (inputs[126]);
    assign layer0_outputs[9005] = ~(inputs[190]) | (inputs[223]);
    assign layer0_outputs[9006] = (inputs[175]) | (inputs[141]);
    assign layer0_outputs[9007] = (inputs[144]) ^ (inputs[178]);
    assign layer0_outputs[9008] = 1'b0;
    assign layer0_outputs[9009] = ~((inputs[222]) | (inputs[187]));
    assign layer0_outputs[9010] = ~((inputs[64]) ^ (inputs[24]));
    assign layer0_outputs[9011] = ~(inputs[83]);
    assign layer0_outputs[9012] = inputs[96];
    assign layer0_outputs[9013] = ~((inputs[80]) ^ (inputs[77]));
    assign layer0_outputs[9014] = ~((inputs[59]) | (inputs[2]));
    assign layer0_outputs[9015] = ~(inputs[156]) | (inputs[254]);
    assign layer0_outputs[9016] = (inputs[125]) | (inputs[123]);
    assign layer0_outputs[9017] = (inputs[227]) | (inputs[208]);
    assign layer0_outputs[9018] = (inputs[42]) & ~(inputs[133]);
    assign layer0_outputs[9019] = inputs[146];
    assign layer0_outputs[9020] = inputs[232];
    assign layer0_outputs[9021] = inputs[47];
    assign layer0_outputs[9022] = ~(inputs[83]) | (inputs[199]);
    assign layer0_outputs[9023] = ~(inputs[130]);
    assign layer0_outputs[9024] = (inputs[157]) ^ (inputs[78]);
    assign layer0_outputs[9025] = inputs[8];
    assign layer0_outputs[9026] = ~(inputs[66]);
    assign layer0_outputs[9027] = (inputs[23]) & ~(inputs[174]);
    assign layer0_outputs[9028] = (inputs[143]) ^ (inputs[204]);
    assign layer0_outputs[9029] = ~(inputs[81]) | (inputs[178]);
    assign layer0_outputs[9030] = ~((inputs[172]) | (inputs[128]));
    assign layer0_outputs[9031] = ~(inputs[84]);
    assign layer0_outputs[9032] = ~((inputs[132]) | (inputs[146]));
    assign layer0_outputs[9033] = ~((inputs[1]) ^ (inputs[43]));
    assign layer0_outputs[9034] = ~((inputs[82]) ^ (inputs[203]));
    assign layer0_outputs[9035] = ~(inputs[51]) | (inputs[223]);
    assign layer0_outputs[9036] = ~(inputs[66]) | (inputs[156]);
    assign layer0_outputs[9037] = (inputs[87]) ^ (inputs[132]);
    assign layer0_outputs[9038] = (inputs[218]) & ~(inputs[94]);
    assign layer0_outputs[9039] = ~(inputs[75]) | (inputs[150]);
    assign layer0_outputs[9040] = (inputs[169]) | (inputs[70]);
    assign layer0_outputs[9041] = ~((inputs[103]) | (inputs[159]));
    assign layer0_outputs[9042] = (inputs[83]) | (inputs[168]);
    assign layer0_outputs[9043] = inputs[193];
    assign layer0_outputs[9044] = inputs[189];
    assign layer0_outputs[9045] = (inputs[1]) | (inputs[34]);
    assign layer0_outputs[9046] = ~((inputs[219]) | (inputs[192]));
    assign layer0_outputs[9047] = ~(inputs[54]) | (inputs[158]);
    assign layer0_outputs[9048] = ~(inputs[98]);
    assign layer0_outputs[9049] = ~((inputs[134]) | (inputs[171]));
    assign layer0_outputs[9050] = inputs[216];
    assign layer0_outputs[9051] = (inputs[125]) & ~(inputs[186]);
    assign layer0_outputs[9052] = (inputs[132]) & ~(inputs[136]);
    assign layer0_outputs[9053] = inputs[158];
    assign layer0_outputs[9054] = inputs[25];
    assign layer0_outputs[9055] = ~((inputs[219]) | (inputs[192]));
    assign layer0_outputs[9056] = ~((inputs[0]) ^ (inputs[209]));
    assign layer0_outputs[9057] = ~(inputs[178]);
    assign layer0_outputs[9058] = ~(inputs[11]) | (inputs[32]);
    assign layer0_outputs[9059] = ~(inputs[84]);
    assign layer0_outputs[9060] = (inputs[58]) & ~(inputs[37]);
    assign layer0_outputs[9061] = ~(inputs[193]);
    assign layer0_outputs[9062] = (inputs[187]) & ~(inputs[54]);
    assign layer0_outputs[9063] = ~((inputs[212]) | (inputs[208]));
    assign layer0_outputs[9064] = (inputs[98]) | (inputs[160]);
    assign layer0_outputs[9065] = 1'b1;
    assign layer0_outputs[9066] = (inputs[48]) ^ (inputs[254]);
    assign layer0_outputs[9067] = (inputs[168]) | (inputs[233]);
    assign layer0_outputs[9068] = inputs[135];
    assign layer0_outputs[9069] = ~(inputs[80]) | (inputs[159]);
    assign layer0_outputs[9070] = ~((inputs[14]) ^ (inputs[45]));
    assign layer0_outputs[9071] = ~((inputs[205]) | (inputs[44]));
    assign layer0_outputs[9072] = ~(inputs[248]);
    assign layer0_outputs[9073] = ~(inputs[181]);
    assign layer0_outputs[9074] = inputs[118];
    assign layer0_outputs[9075] = (inputs[195]) & (inputs[59]);
    assign layer0_outputs[9076] = (inputs[215]) & ~(inputs[253]);
    assign layer0_outputs[9077] = (inputs[100]) & ~(inputs[202]);
    assign layer0_outputs[9078] = 1'b0;
    assign layer0_outputs[9079] = ~(inputs[43]) | (inputs[179]);
    assign layer0_outputs[9080] = ~((inputs[1]) | (inputs[162]));
    assign layer0_outputs[9081] = (inputs[57]) | (inputs[202]);
    assign layer0_outputs[9082] = (inputs[83]) & ~(inputs[249]);
    assign layer0_outputs[9083] = ~(inputs[229]);
    assign layer0_outputs[9084] = (inputs[246]) ^ (inputs[40]);
    assign layer0_outputs[9085] = (inputs[30]) | (inputs[67]);
    assign layer0_outputs[9086] = (inputs[39]) & (inputs[154]);
    assign layer0_outputs[9087] = ~(inputs[201]);
    assign layer0_outputs[9088] = (inputs[116]) ^ (inputs[129]);
    assign layer0_outputs[9089] = ~((inputs[92]) | (inputs[239]));
    assign layer0_outputs[9090] = ~(inputs[217]);
    assign layer0_outputs[9091] = (inputs[161]) | (inputs[80]);
    assign layer0_outputs[9092] = ~(inputs[241]);
    assign layer0_outputs[9093] = ~(inputs[57]);
    assign layer0_outputs[9094] = ~((inputs[37]) | (inputs[50]));
    assign layer0_outputs[9095] = (inputs[46]) ^ (inputs[18]);
    assign layer0_outputs[9096] = inputs[119];
    assign layer0_outputs[9097] = ~(inputs[92]) | (inputs[4]);
    assign layer0_outputs[9098] = ~(inputs[107]);
    assign layer0_outputs[9099] = ~((inputs[95]) & (inputs[145]));
    assign layer0_outputs[9100] = ~(inputs[170]);
    assign layer0_outputs[9101] = inputs[89];
    assign layer0_outputs[9102] = ~((inputs[249]) & (inputs[135]));
    assign layer0_outputs[9103] = ~(inputs[254]);
    assign layer0_outputs[9104] = inputs[124];
    assign layer0_outputs[9105] = (inputs[242]) | (inputs[221]);
    assign layer0_outputs[9106] = ~((inputs[56]) | (inputs[86]));
    assign layer0_outputs[9107] = ~(inputs[205]) | (inputs[87]);
    assign layer0_outputs[9108] = ~(inputs[67]) | (inputs[235]);
    assign layer0_outputs[9109] = ~((inputs[209]) | (inputs[252]));
    assign layer0_outputs[9110] = inputs[56];
    assign layer0_outputs[9111] = inputs[203];
    assign layer0_outputs[9112] = ~((inputs[25]) ^ (inputs[47]));
    assign layer0_outputs[9113] = ~(inputs[146]) | (inputs[47]);
    assign layer0_outputs[9114] = ~(inputs[89]);
    assign layer0_outputs[9115] = ~((inputs[242]) ^ (inputs[194]));
    assign layer0_outputs[9116] = (inputs[74]) | (inputs[77]);
    assign layer0_outputs[9117] = ~((inputs[177]) | (inputs[85]));
    assign layer0_outputs[9118] = (inputs[32]) & ~(inputs[223]);
    assign layer0_outputs[9119] = ~((inputs[3]) | (inputs[137]));
    assign layer0_outputs[9120] = inputs[103];
    assign layer0_outputs[9121] = ~(inputs[221]);
    assign layer0_outputs[9122] = inputs[178];
    assign layer0_outputs[9123] = inputs[203];
    assign layer0_outputs[9124] = (inputs[142]) ^ (inputs[20]);
    assign layer0_outputs[9125] = ~(inputs[129]);
    assign layer0_outputs[9126] = ~((inputs[135]) | (inputs[78]));
    assign layer0_outputs[9127] = ~(inputs[215]) | (inputs[41]);
    assign layer0_outputs[9128] = inputs[23];
    assign layer0_outputs[9129] = ~(inputs[125]) | (inputs[241]);
    assign layer0_outputs[9130] = (inputs[124]) & (inputs[236]);
    assign layer0_outputs[9131] = (inputs[13]) ^ (inputs[243]);
    assign layer0_outputs[9132] = ~(inputs[105]) | (inputs[149]);
    assign layer0_outputs[9133] = ~(inputs[231]) | (inputs[252]);
    assign layer0_outputs[9134] = (inputs[52]) & ~(inputs[56]);
    assign layer0_outputs[9135] = ~(inputs[54]);
    assign layer0_outputs[9136] = ~(inputs[181]) | (inputs[63]);
    assign layer0_outputs[9137] = inputs[134];
    assign layer0_outputs[9138] = inputs[205];
    assign layer0_outputs[9139] = (inputs[213]) & ~(inputs[165]);
    assign layer0_outputs[9140] = (inputs[14]) | (inputs[97]);
    assign layer0_outputs[9141] = (inputs[204]) ^ (inputs[26]);
    assign layer0_outputs[9142] = ~((inputs[48]) | (inputs[122]));
    assign layer0_outputs[9143] = (inputs[73]) | (inputs[198]);
    assign layer0_outputs[9144] = (inputs[144]) ^ (inputs[53]);
    assign layer0_outputs[9145] = ~(inputs[67]) | (inputs[54]);
    assign layer0_outputs[9146] = (inputs[57]) & ~(inputs[33]);
    assign layer0_outputs[9147] = ~(inputs[91]);
    assign layer0_outputs[9148] = (inputs[0]) & ~(inputs[138]);
    assign layer0_outputs[9149] = ~(inputs[113]);
    assign layer0_outputs[9150] = (inputs[146]) ^ (inputs[183]);
    assign layer0_outputs[9151] = ~((inputs[87]) | (inputs[86]));
    assign layer0_outputs[9152] = inputs[145];
    assign layer0_outputs[9153] = inputs[103];
    assign layer0_outputs[9154] = ~(inputs[39]);
    assign layer0_outputs[9155] = (inputs[244]) & (inputs[215]);
    assign layer0_outputs[9156] = ~((inputs[74]) ^ (inputs[88]));
    assign layer0_outputs[9157] = ~((inputs[168]) ^ (inputs[199]));
    assign layer0_outputs[9158] = (inputs[245]) & ~(inputs[189]);
    assign layer0_outputs[9159] = ~((inputs[27]) ^ (inputs[245]));
    assign layer0_outputs[9160] = (inputs[13]) & ~(inputs[160]);
    assign layer0_outputs[9161] = inputs[36];
    assign layer0_outputs[9162] = ~((inputs[165]) ^ (inputs[61]));
    assign layer0_outputs[9163] = (inputs[149]) & (inputs[244]);
    assign layer0_outputs[9164] = ~((inputs[132]) ^ (inputs[237]));
    assign layer0_outputs[9165] = ~((inputs[123]) | (inputs[29]));
    assign layer0_outputs[9166] = ~(inputs[163]);
    assign layer0_outputs[9167] = (inputs[177]) & ~(inputs[177]);
    assign layer0_outputs[9168] = ~(inputs[56]) | (inputs[140]);
    assign layer0_outputs[9169] = ~(inputs[206]) | (inputs[82]);
    assign layer0_outputs[9170] = ~((inputs[139]) | (inputs[153]));
    assign layer0_outputs[9171] = ~((inputs[160]) & (inputs[193]));
    assign layer0_outputs[9172] = ~((inputs[251]) ^ (inputs[17]));
    assign layer0_outputs[9173] = ~(inputs[230]) | (inputs[147]);
    assign layer0_outputs[9174] = ~((inputs[180]) | (inputs[191]));
    assign layer0_outputs[9175] = (inputs[223]) | (inputs[72]);
    assign layer0_outputs[9176] = (inputs[155]) | (inputs[225]);
    assign layer0_outputs[9177] = inputs[60];
    assign layer0_outputs[9178] = ~(inputs[52]) | (inputs[135]);
    assign layer0_outputs[9179] = (inputs[152]) | (inputs[62]);
    assign layer0_outputs[9180] = (inputs[29]) | (inputs[146]);
    assign layer0_outputs[9181] = ~((inputs[76]) ^ (inputs[57]));
    assign layer0_outputs[9182] = (inputs[167]) & ~(inputs[52]);
    assign layer0_outputs[9183] = ~(inputs[134]) | (inputs[200]);
    assign layer0_outputs[9184] = (inputs[105]) | (inputs[96]);
    assign layer0_outputs[9185] = (inputs[30]) ^ (inputs[188]);
    assign layer0_outputs[9186] = ~(inputs[192]) | (inputs[11]);
    assign layer0_outputs[9187] = ~(inputs[4]);
    assign layer0_outputs[9188] = ~(inputs[142]) | (inputs[6]);
    assign layer0_outputs[9189] = (inputs[5]) & ~(inputs[255]);
    assign layer0_outputs[9190] = ~(inputs[20]);
    assign layer0_outputs[9191] = inputs[77];
    assign layer0_outputs[9192] = ~(inputs[233]) | (inputs[110]);
    assign layer0_outputs[9193] = ~((inputs[245]) & (inputs[21]));
    assign layer0_outputs[9194] = ~((inputs[223]) ^ (inputs[143]));
    assign layer0_outputs[9195] = ~(inputs[248]);
    assign layer0_outputs[9196] = ~(inputs[39]);
    assign layer0_outputs[9197] = ~((inputs[110]) | (inputs[197]));
    assign layer0_outputs[9198] = 1'b0;
    assign layer0_outputs[9199] = (inputs[63]) | (inputs[216]);
    assign layer0_outputs[9200] = inputs[133];
    assign layer0_outputs[9201] = ~((inputs[186]) | (inputs[132]));
    assign layer0_outputs[9202] = (inputs[136]) ^ (inputs[156]);
    assign layer0_outputs[9203] = (inputs[177]) ^ (inputs[75]);
    assign layer0_outputs[9204] = ~(inputs[218]) | (inputs[107]);
    assign layer0_outputs[9205] = 1'b0;
    assign layer0_outputs[9206] = (inputs[167]) | (inputs[157]);
    assign layer0_outputs[9207] = (inputs[129]) & (inputs[158]);
    assign layer0_outputs[9208] = inputs[135];
    assign layer0_outputs[9209] = (inputs[172]) | (inputs[203]);
    assign layer0_outputs[9210] = ~(inputs[145]);
    assign layer0_outputs[9211] = (inputs[233]) ^ (inputs[58]);
    assign layer0_outputs[9212] = ~(inputs[117]);
    assign layer0_outputs[9213] = (inputs[193]) | (inputs[195]);
    assign layer0_outputs[9214] = ~(inputs[151]) | (inputs[109]);
    assign layer0_outputs[9215] = (inputs[119]) ^ (inputs[186]);
    assign layer0_outputs[9216] = (inputs[218]) ^ (inputs[114]);
    assign layer0_outputs[9217] = ~(inputs[228]) | (inputs[49]);
    assign layer0_outputs[9218] = (inputs[249]) & ~(inputs[146]);
    assign layer0_outputs[9219] = (inputs[94]) & ~(inputs[12]);
    assign layer0_outputs[9220] = (inputs[179]) | (inputs[196]);
    assign layer0_outputs[9221] = ~(inputs[166]) | (inputs[4]);
    assign layer0_outputs[9222] = ~(inputs[183]) | (inputs[54]);
    assign layer0_outputs[9223] = (inputs[118]) ^ (inputs[87]);
    assign layer0_outputs[9224] = (inputs[82]) & ~(inputs[242]);
    assign layer0_outputs[9225] = (inputs[130]) ^ (inputs[167]);
    assign layer0_outputs[9226] = ~((inputs[55]) ^ (inputs[11]));
    assign layer0_outputs[9227] = inputs[110];
    assign layer0_outputs[9228] = ~((inputs[116]) | (inputs[157]));
    assign layer0_outputs[9229] = (inputs[176]) ^ (inputs[18]);
    assign layer0_outputs[9230] = (inputs[198]) | (inputs[148]);
    assign layer0_outputs[9231] = ~((inputs[110]) ^ (inputs[16]));
    assign layer0_outputs[9232] = (inputs[48]) & ~(inputs[193]);
    assign layer0_outputs[9233] = (inputs[24]) & (inputs[25]);
    assign layer0_outputs[9234] = ~((inputs[248]) & (inputs[169]));
    assign layer0_outputs[9235] = (inputs[130]) ^ (inputs[22]);
    assign layer0_outputs[9236] = ~(inputs[105]) | (inputs[17]);
    assign layer0_outputs[9237] = ~(inputs[10]);
    assign layer0_outputs[9238] = ~(inputs[129]);
    assign layer0_outputs[9239] = ~(inputs[181]) | (inputs[144]);
    assign layer0_outputs[9240] = inputs[89];
    assign layer0_outputs[9241] = ~((inputs[81]) | (inputs[12]));
    assign layer0_outputs[9242] = (inputs[153]) ^ (inputs[140]);
    assign layer0_outputs[9243] = ~((inputs[12]) | (inputs[134]));
    assign layer0_outputs[9244] = ~((inputs[23]) ^ (inputs[187]));
    assign layer0_outputs[9245] = ~(inputs[157]) | (inputs[17]);
    assign layer0_outputs[9246] = ~(inputs[122]) | (inputs[179]);
    assign layer0_outputs[9247] = (inputs[226]) | (inputs[178]);
    assign layer0_outputs[9248] = ~((inputs[167]) | (inputs[152]));
    assign layer0_outputs[9249] = ~((inputs[74]) | (inputs[128]));
    assign layer0_outputs[9250] = ~((inputs[181]) ^ (inputs[133]));
    assign layer0_outputs[9251] = ~((inputs[64]) ^ (inputs[90]));
    assign layer0_outputs[9252] = (inputs[93]) | (inputs[8]);
    assign layer0_outputs[9253] = ~(inputs[78]);
    assign layer0_outputs[9254] = ~((inputs[211]) ^ (inputs[38]));
    assign layer0_outputs[9255] = (inputs[63]) | (inputs[86]);
    assign layer0_outputs[9256] = inputs[107];
    assign layer0_outputs[9257] = (inputs[45]) | (inputs[185]);
    assign layer0_outputs[9258] = (inputs[95]) & (inputs[189]);
    assign layer0_outputs[9259] = ~((inputs[24]) | (inputs[94]));
    assign layer0_outputs[9260] = (inputs[168]) | (inputs[250]);
    assign layer0_outputs[9261] = (inputs[84]) & ~(inputs[8]);
    assign layer0_outputs[9262] = ~((inputs[51]) | (inputs[31]));
    assign layer0_outputs[9263] = ~(inputs[147]) | (inputs[228]);
    assign layer0_outputs[9264] = (inputs[34]) ^ (inputs[7]);
    assign layer0_outputs[9265] = inputs[155];
    assign layer0_outputs[9266] = ~(inputs[113]);
    assign layer0_outputs[9267] = (inputs[154]) & ~(inputs[76]);
    assign layer0_outputs[9268] = (inputs[176]) & (inputs[219]);
    assign layer0_outputs[9269] = inputs[106];
    assign layer0_outputs[9270] = ~(inputs[128]) | (inputs[238]);
    assign layer0_outputs[9271] = ~(inputs[231]);
    assign layer0_outputs[9272] = ~(inputs[52]);
    assign layer0_outputs[9273] = (inputs[151]) & (inputs[85]);
    assign layer0_outputs[9274] = ~(inputs[149]);
    assign layer0_outputs[9275] = inputs[8];
    assign layer0_outputs[9276] = ~((inputs[223]) | (inputs[229]));
    assign layer0_outputs[9277] = (inputs[67]) | (inputs[185]);
    assign layer0_outputs[9278] = ~(inputs[187]);
    assign layer0_outputs[9279] = (inputs[41]) | (inputs[80]);
    assign layer0_outputs[9280] = ~(inputs[124]);
    assign layer0_outputs[9281] = (inputs[191]) | (inputs[88]);
    assign layer0_outputs[9282] = ~(inputs[96]);
    assign layer0_outputs[9283] = (inputs[242]) & (inputs[70]);
    assign layer0_outputs[9284] = ~((inputs[141]) | (inputs[189]));
    assign layer0_outputs[9285] = inputs[162];
    assign layer0_outputs[9286] = ~(inputs[196]);
    assign layer0_outputs[9287] = (inputs[217]) & ~(inputs[108]);
    assign layer0_outputs[9288] = inputs[131];
    assign layer0_outputs[9289] = ~(inputs[67]);
    assign layer0_outputs[9290] = (inputs[40]) | (inputs[47]);
    assign layer0_outputs[9291] = inputs[247];
    assign layer0_outputs[9292] = inputs[25];
    assign layer0_outputs[9293] = (inputs[217]) & ~(inputs[96]);
    assign layer0_outputs[9294] = (inputs[16]) | (inputs[90]);
    assign layer0_outputs[9295] = inputs[28];
    assign layer0_outputs[9296] = (inputs[73]) ^ (inputs[71]);
    assign layer0_outputs[9297] = inputs[12];
    assign layer0_outputs[9298] = (inputs[5]) ^ (inputs[79]);
    assign layer0_outputs[9299] = ~(inputs[134]) | (inputs[158]);
    assign layer0_outputs[9300] = (inputs[178]) & ~(inputs[47]);
    assign layer0_outputs[9301] = inputs[135];
    assign layer0_outputs[9302] = ~(inputs[140]);
    assign layer0_outputs[9303] = ~(inputs[209]);
    assign layer0_outputs[9304] = inputs[249];
    assign layer0_outputs[9305] = ~(inputs[173]);
    assign layer0_outputs[9306] = ~((inputs[121]) ^ (inputs[180]));
    assign layer0_outputs[9307] = inputs[36];
    assign layer0_outputs[9308] = ~(inputs[249]);
    assign layer0_outputs[9309] = ~(inputs[162]);
    assign layer0_outputs[9310] = ~(inputs[44]);
    assign layer0_outputs[9311] = ~(inputs[165]);
    assign layer0_outputs[9312] = (inputs[173]) ^ (inputs[131]);
    assign layer0_outputs[9313] = ~(inputs[130]);
    assign layer0_outputs[9314] = (inputs[8]) & ~(inputs[74]);
    assign layer0_outputs[9315] = inputs[22];
    assign layer0_outputs[9316] = inputs[109];
    assign layer0_outputs[9317] = (inputs[11]) ^ (inputs[9]);
    assign layer0_outputs[9318] = ~(inputs[69]) | (inputs[48]);
    assign layer0_outputs[9319] = ~(inputs[70]) | (inputs[62]);
    assign layer0_outputs[9320] = (inputs[243]) & (inputs[169]);
    assign layer0_outputs[9321] = (inputs[208]) | (inputs[111]);
    assign layer0_outputs[9322] = ~((inputs[90]) ^ (inputs[29]));
    assign layer0_outputs[9323] = inputs[17];
    assign layer0_outputs[9324] = (inputs[40]) & ~(inputs[81]);
    assign layer0_outputs[9325] = inputs[34];
    assign layer0_outputs[9326] = (inputs[54]) | (inputs[180]);
    assign layer0_outputs[9327] = inputs[126];
    assign layer0_outputs[9328] = (inputs[49]) ^ (inputs[234]);
    assign layer0_outputs[9329] = ~(inputs[76]);
    assign layer0_outputs[9330] = ~((inputs[70]) | (inputs[112]));
    assign layer0_outputs[9331] = 1'b1;
    assign layer0_outputs[9332] = ~((inputs[196]) & (inputs[100]));
    assign layer0_outputs[9333] = (inputs[39]) & ~(inputs[88]);
    assign layer0_outputs[9334] = ~((inputs[74]) ^ (inputs[215]));
    assign layer0_outputs[9335] = ~(inputs[200]) | (inputs[201]);
    assign layer0_outputs[9336] = (inputs[199]) ^ (inputs[185]);
    assign layer0_outputs[9337] = (inputs[42]) | (inputs[14]);
    assign layer0_outputs[9338] = ~((inputs[54]) | (inputs[65]));
    assign layer0_outputs[9339] = (inputs[6]) | (inputs[145]);
    assign layer0_outputs[9340] = (inputs[187]) & ~(inputs[10]);
    assign layer0_outputs[9341] = (inputs[246]) | (inputs[189]);
    assign layer0_outputs[9342] = (inputs[188]) | (inputs[211]);
    assign layer0_outputs[9343] = ~((inputs[37]) | (inputs[192]));
    assign layer0_outputs[9344] = (inputs[219]) ^ (inputs[103]);
    assign layer0_outputs[9345] = (inputs[91]) ^ (inputs[218]);
    assign layer0_outputs[9346] = ~(inputs[51]) | (inputs[225]);
    assign layer0_outputs[9347] = (inputs[225]) ^ (inputs[175]);
    assign layer0_outputs[9348] = ~(inputs[138]);
    assign layer0_outputs[9349] = inputs[39];
    assign layer0_outputs[9350] = ~(inputs[113]);
    assign layer0_outputs[9351] = inputs[146];
    assign layer0_outputs[9352] = 1'b1;
    assign layer0_outputs[9353] = (inputs[121]) & ~(inputs[244]);
    assign layer0_outputs[9354] = (inputs[46]) ^ (inputs[73]);
    assign layer0_outputs[9355] = ~(inputs[40]) | (inputs[193]);
    assign layer0_outputs[9356] = ~(inputs[207]) | (inputs[177]);
    assign layer0_outputs[9357] = inputs[210];
    assign layer0_outputs[9358] = (inputs[225]) | (inputs[162]);
    assign layer0_outputs[9359] = inputs[122];
    assign layer0_outputs[9360] = (inputs[89]) & ~(inputs[160]);
    assign layer0_outputs[9361] = ~((inputs[245]) | (inputs[235]));
    assign layer0_outputs[9362] = ~((inputs[174]) | (inputs[199]));
    assign layer0_outputs[9363] = (inputs[34]) ^ (inputs[235]);
    assign layer0_outputs[9364] = ~(inputs[206]);
    assign layer0_outputs[9365] = inputs[45];
    assign layer0_outputs[9366] = (inputs[51]) | (inputs[207]);
    assign layer0_outputs[9367] = ~((inputs[7]) ^ (inputs[79]));
    assign layer0_outputs[9368] = ~(inputs[160]);
    assign layer0_outputs[9369] = ~(inputs[78]);
    assign layer0_outputs[9370] = inputs[62];
    assign layer0_outputs[9371] = ~((inputs[164]) & (inputs[186]));
    assign layer0_outputs[9372] = ~((inputs[53]) ^ (inputs[51]));
    assign layer0_outputs[9373] = inputs[148];
    assign layer0_outputs[9374] = ~((inputs[126]) | (inputs[1]));
    assign layer0_outputs[9375] = (inputs[132]) & (inputs[72]);
    assign layer0_outputs[9376] = ~(inputs[186]) | (inputs[48]);
    assign layer0_outputs[9377] = ~((inputs[33]) ^ (inputs[49]));
    assign layer0_outputs[9378] = inputs[197];
    assign layer0_outputs[9379] = inputs[230];
    assign layer0_outputs[9380] = ~((inputs[241]) ^ (inputs[46]));
    assign layer0_outputs[9381] = (inputs[142]) | (inputs[112]);
    assign layer0_outputs[9382] = ~(inputs[68]) | (inputs[173]);
    assign layer0_outputs[9383] = ~(inputs[212]);
    assign layer0_outputs[9384] = (inputs[47]) | (inputs[60]);
    assign layer0_outputs[9385] = ~((inputs[13]) & (inputs[12]));
    assign layer0_outputs[9386] = (inputs[18]) & ~(inputs[175]);
    assign layer0_outputs[9387] = (inputs[78]) ^ (inputs[127]);
    assign layer0_outputs[9388] = (inputs[106]) & ~(inputs[232]);
    assign layer0_outputs[9389] = ~((inputs[183]) | (inputs[64]));
    assign layer0_outputs[9390] = inputs[179];
    assign layer0_outputs[9391] = inputs[198];
    assign layer0_outputs[9392] = inputs[14];
    assign layer0_outputs[9393] = (inputs[168]) ^ (inputs[179]);
    assign layer0_outputs[9394] = ~((inputs[11]) | (inputs[104]));
    assign layer0_outputs[9395] = ~((inputs[181]) | (inputs[239]));
    assign layer0_outputs[9396] = (inputs[9]) & ~(inputs[15]);
    assign layer0_outputs[9397] = (inputs[48]) | (inputs[172]);
    assign layer0_outputs[9398] = 1'b1;
    assign layer0_outputs[9399] = 1'b1;
    assign layer0_outputs[9400] = inputs[209];
    assign layer0_outputs[9401] = ~(inputs[245]) | (inputs[20]);
    assign layer0_outputs[9402] = ~((inputs[4]) ^ (inputs[118]));
    assign layer0_outputs[9403] = (inputs[12]) | (inputs[195]);
    assign layer0_outputs[9404] = (inputs[135]) & ~(inputs[110]);
    assign layer0_outputs[9405] = (inputs[46]) | (inputs[190]);
    assign layer0_outputs[9406] = ~((inputs[144]) ^ (inputs[164]));
    assign layer0_outputs[9407] = (inputs[183]) & ~(inputs[117]);
    assign layer0_outputs[9408] = (inputs[131]) & ~(inputs[250]);
    assign layer0_outputs[9409] = ~(inputs[105]);
    assign layer0_outputs[9410] = ~((inputs[6]) ^ (inputs[69]));
    assign layer0_outputs[9411] = inputs[93];
    assign layer0_outputs[9412] = ~((inputs[191]) ^ (inputs[180]));
    assign layer0_outputs[9413] = ~(inputs[145]);
    assign layer0_outputs[9414] = ~(inputs[36]);
    assign layer0_outputs[9415] = ~(inputs[97]);
    assign layer0_outputs[9416] = ~(inputs[183]) | (inputs[140]);
    assign layer0_outputs[9417] = (inputs[242]) ^ (inputs[124]);
    assign layer0_outputs[9418] = (inputs[86]) & ~(inputs[94]);
    assign layer0_outputs[9419] = ~((inputs[6]) | (inputs[17]));
    assign layer0_outputs[9420] = inputs[78];
    assign layer0_outputs[9421] = (inputs[190]) & ~(inputs[191]);
    assign layer0_outputs[9422] = ~(inputs[8]);
    assign layer0_outputs[9423] = ~((inputs[44]) ^ (inputs[59]));
    assign layer0_outputs[9424] = inputs[88];
    assign layer0_outputs[9425] = (inputs[49]) & ~(inputs[138]);
    assign layer0_outputs[9426] = ~(inputs[85]);
    assign layer0_outputs[9427] = ~((inputs[251]) | (inputs[228]));
    assign layer0_outputs[9428] = ~(inputs[110]) | (inputs[32]);
    assign layer0_outputs[9429] = inputs[232];
    assign layer0_outputs[9430] = ~((inputs[98]) ^ (inputs[194]));
    assign layer0_outputs[9431] = ~(inputs[37]) | (inputs[180]);
    assign layer0_outputs[9432] = ~(inputs[123]) | (inputs[151]);
    assign layer0_outputs[9433] = ~((inputs[46]) | (inputs[248]));
    assign layer0_outputs[9434] = ~(inputs[236]);
    assign layer0_outputs[9435] = ~(inputs[110]);
    assign layer0_outputs[9436] = (inputs[207]) | (inputs[79]);
    assign layer0_outputs[9437] = ~((inputs[224]) | (inputs[247]));
    assign layer0_outputs[9438] = (inputs[201]) | (inputs[17]);
    assign layer0_outputs[9439] = (inputs[60]) ^ (inputs[91]);
    assign layer0_outputs[9440] = inputs[34];
    assign layer0_outputs[9441] = (inputs[238]) ^ (inputs[131]);
    assign layer0_outputs[9442] = (inputs[99]) ^ (inputs[227]);
    assign layer0_outputs[9443] = ~((inputs[120]) | (inputs[135]));
    assign layer0_outputs[9444] = ~((inputs[57]) ^ (inputs[173]));
    assign layer0_outputs[9445] = (inputs[36]) & ~(inputs[156]);
    assign layer0_outputs[9446] = ~(inputs[2]) | (inputs[86]);
    assign layer0_outputs[9447] = (inputs[180]) | (inputs[245]);
    assign layer0_outputs[9448] = ~((inputs[113]) ^ (inputs[84]));
    assign layer0_outputs[9449] = ~((inputs[108]) | (inputs[16]));
    assign layer0_outputs[9450] = (inputs[250]) & ~(inputs[11]);
    assign layer0_outputs[9451] = ~(inputs[114]) | (inputs[80]);
    assign layer0_outputs[9452] = ~((inputs[193]) | (inputs[244]));
    assign layer0_outputs[9453] = (inputs[154]) & ~(inputs[5]);
    assign layer0_outputs[9454] = ~(inputs[15]);
    assign layer0_outputs[9455] = ~(inputs[25]);
    assign layer0_outputs[9456] = inputs[88];
    assign layer0_outputs[9457] = ~(inputs[59]);
    assign layer0_outputs[9458] = ~((inputs[171]) | (inputs[27]));
    assign layer0_outputs[9459] = ~((inputs[32]) | (inputs[17]));
    assign layer0_outputs[9460] = inputs[118];
    assign layer0_outputs[9461] = inputs[25];
    assign layer0_outputs[9462] = (inputs[22]) ^ (inputs[9]);
    assign layer0_outputs[9463] = ~(inputs[231]);
    assign layer0_outputs[9464] = (inputs[243]) | (inputs[9]);
    assign layer0_outputs[9465] = inputs[25];
    assign layer0_outputs[9466] = inputs[102];
    assign layer0_outputs[9467] = 1'b1;
    assign layer0_outputs[9468] = inputs[81];
    assign layer0_outputs[9469] = (inputs[156]) & ~(inputs[127]);
    assign layer0_outputs[9470] = ~((inputs[10]) | (inputs[125]));
    assign layer0_outputs[9471] = inputs[53];
    assign layer0_outputs[9472] = ~(inputs[189]);
    assign layer0_outputs[9473] = (inputs[211]) ^ (inputs[198]);
    assign layer0_outputs[9474] = (inputs[235]) & (inputs[5]);
    assign layer0_outputs[9475] = inputs[232];
    assign layer0_outputs[9476] = inputs[84];
    assign layer0_outputs[9477] = ~(inputs[112]);
    assign layer0_outputs[9478] = (inputs[47]) | (inputs[31]);
    assign layer0_outputs[9479] = ~(inputs[89]) | (inputs[115]);
    assign layer0_outputs[9480] = ~(inputs[164]);
    assign layer0_outputs[9481] = ~(inputs[248]);
    assign layer0_outputs[9482] = ~(inputs[128]);
    assign layer0_outputs[9483] = inputs[217];
    assign layer0_outputs[9484] = ~((inputs[113]) ^ (inputs[244]));
    assign layer0_outputs[9485] = ~(inputs[44]) | (inputs[95]);
    assign layer0_outputs[9486] = ~((inputs[44]) & (inputs[159]));
    assign layer0_outputs[9487] = 1'b0;
    assign layer0_outputs[9488] = ~(inputs[250]);
    assign layer0_outputs[9489] = inputs[87];
    assign layer0_outputs[9490] = ~(inputs[124]);
    assign layer0_outputs[9491] = inputs[71];
    assign layer0_outputs[9492] = (inputs[88]) & ~(inputs[36]);
    assign layer0_outputs[9493] = ~((inputs[78]) ^ (inputs[76]));
    assign layer0_outputs[9494] = (inputs[131]) & ~(inputs[192]);
    assign layer0_outputs[9495] = ~(inputs[187]);
    assign layer0_outputs[9496] = ~(inputs[42]) | (inputs[80]);
    assign layer0_outputs[9497] = ~(inputs[122]);
    assign layer0_outputs[9498] = ~((inputs[222]) | (inputs[221]));
    assign layer0_outputs[9499] = ~((inputs[20]) & (inputs[187]));
    assign layer0_outputs[9500] = (inputs[177]) | (inputs[213]);
    assign layer0_outputs[9501] = (inputs[4]) | (inputs[168]);
    assign layer0_outputs[9502] = (inputs[236]) & ~(inputs[32]);
    assign layer0_outputs[9503] = ~(inputs[107]);
    assign layer0_outputs[9504] = (inputs[218]) & ~(inputs[133]);
    assign layer0_outputs[9505] = ~(inputs[120]);
    assign layer0_outputs[9506] = ~((inputs[226]) | (inputs[212]));
    assign layer0_outputs[9507] = (inputs[169]) & ~(inputs[117]);
    assign layer0_outputs[9508] = ~((inputs[72]) | (inputs[170]));
    assign layer0_outputs[9509] = (inputs[93]) ^ (inputs[106]);
    assign layer0_outputs[9510] = inputs[124];
    assign layer0_outputs[9511] = (inputs[27]) ^ (inputs[91]);
    assign layer0_outputs[9512] = (inputs[167]) | (inputs[210]);
    assign layer0_outputs[9513] = ~(inputs[60]) | (inputs[205]);
    assign layer0_outputs[9514] = ~((inputs[233]) | (inputs[88]));
    assign layer0_outputs[9515] = inputs[16];
    assign layer0_outputs[9516] = (inputs[75]) & ~(inputs[159]);
    assign layer0_outputs[9517] = ~((inputs[71]) | (inputs[64]));
    assign layer0_outputs[9518] = ~(inputs[25]);
    assign layer0_outputs[9519] = ~((inputs[104]) | (inputs[218]));
    assign layer0_outputs[9520] = (inputs[139]) & ~(inputs[0]);
    assign layer0_outputs[9521] = 1'b1;
    assign layer0_outputs[9522] = ~((inputs[167]) | (inputs[243]));
    assign layer0_outputs[9523] = 1'b1;
    assign layer0_outputs[9524] = ~((inputs[150]) | (inputs[189]));
    assign layer0_outputs[9525] = ~((inputs[60]) ^ (inputs[145]));
    assign layer0_outputs[9526] = ~(inputs[61]);
    assign layer0_outputs[9527] = ~(inputs[60]) | (inputs[80]);
    assign layer0_outputs[9528] = ~((inputs[228]) & (inputs[226]));
    assign layer0_outputs[9529] = ~(inputs[65]) | (inputs[111]);
    assign layer0_outputs[9530] = ~((inputs[99]) | (inputs[46]));
    assign layer0_outputs[9531] = ~((inputs[23]) ^ (inputs[243]));
    assign layer0_outputs[9532] = ~(inputs[60]) | (inputs[2]);
    assign layer0_outputs[9533] = ~(inputs[159]) | (inputs[12]);
    assign layer0_outputs[9534] = (inputs[208]) | (inputs[248]);
    assign layer0_outputs[9535] = ~(inputs[85]);
    assign layer0_outputs[9536] = (inputs[240]) & ~(inputs[90]);
    assign layer0_outputs[9537] = 1'b1;
    assign layer0_outputs[9538] = (inputs[214]) | (inputs[176]);
    assign layer0_outputs[9539] = (inputs[18]) & ~(inputs[79]);
    assign layer0_outputs[9540] = ~(inputs[99]);
    assign layer0_outputs[9541] = (inputs[76]) & (inputs[10]);
    assign layer0_outputs[9542] = ~(inputs[213]);
    assign layer0_outputs[9543] = ~((inputs[183]) ^ (inputs[69]));
    assign layer0_outputs[9544] = (inputs[177]) ^ (inputs[3]);
    assign layer0_outputs[9545] = ~((inputs[168]) | (inputs[113]));
    assign layer0_outputs[9546] = ~(inputs[4]);
    assign layer0_outputs[9547] = ~(inputs[212]) | (inputs[38]);
    assign layer0_outputs[9548] = ~((inputs[113]) | (inputs[27]));
    assign layer0_outputs[9549] = (inputs[226]) ^ (inputs[243]);
    assign layer0_outputs[9550] = ~(inputs[93]);
    assign layer0_outputs[9551] = ~(inputs[107]);
    assign layer0_outputs[9552] = (inputs[61]) | (inputs[236]);
    assign layer0_outputs[9553] = ~(inputs[13]);
    assign layer0_outputs[9554] = ~(inputs[172]);
    assign layer0_outputs[9555] = inputs[130];
    assign layer0_outputs[9556] = (inputs[102]) & ~(inputs[226]);
    assign layer0_outputs[9557] = inputs[92];
    assign layer0_outputs[9558] = ~(inputs[104]) | (inputs[68]);
    assign layer0_outputs[9559] = ~(inputs[152]);
    assign layer0_outputs[9560] = ~(inputs[235]);
    assign layer0_outputs[9561] = ~(inputs[216]);
    assign layer0_outputs[9562] = ~(inputs[65]);
    assign layer0_outputs[9563] = (inputs[108]) & ~(inputs[225]);
    assign layer0_outputs[9564] = ~(inputs[191]) | (inputs[27]);
    assign layer0_outputs[9565] = ~(inputs[242]);
    assign layer0_outputs[9566] = (inputs[24]) ^ (inputs[55]);
    assign layer0_outputs[9567] = (inputs[116]) | (inputs[119]);
    assign layer0_outputs[9568] = ~((inputs[192]) ^ (inputs[151]));
    assign layer0_outputs[9569] = (inputs[162]) | (inputs[216]);
    assign layer0_outputs[9570] = inputs[102];
    assign layer0_outputs[9571] = ~((inputs[167]) | (inputs[238]));
    assign layer0_outputs[9572] = ~((inputs[158]) ^ (inputs[117]));
    assign layer0_outputs[9573] = 1'b1;
    assign layer0_outputs[9574] = ~((inputs[93]) | (inputs[183]));
    assign layer0_outputs[9575] = ~(inputs[118]);
    assign layer0_outputs[9576] = ~((inputs[190]) | (inputs[63]));
    assign layer0_outputs[9577] = ~((inputs[224]) | (inputs[213]));
    assign layer0_outputs[9578] = ~((inputs[97]) ^ (inputs[147]));
    assign layer0_outputs[9579] = (inputs[121]) | (inputs[239]);
    assign layer0_outputs[9580] = ~((inputs[164]) ^ (inputs[195]));
    assign layer0_outputs[9581] = (inputs[192]) ^ (inputs[174]);
    assign layer0_outputs[9582] = ~((inputs[222]) | (inputs[25]));
    assign layer0_outputs[9583] = ~((inputs[99]) ^ (inputs[121]));
    assign layer0_outputs[9584] = 1'b0;
    assign layer0_outputs[9585] = ~(inputs[7]) | (inputs[71]);
    assign layer0_outputs[9586] = (inputs[73]) & ~(inputs[255]);
    assign layer0_outputs[9587] = ~((inputs[6]) ^ (inputs[133]));
    assign layer0_outputs[9588] = ~((inputs[67]) | (inputs[77]));
    assign layer0_outputs[9589] = ~(inputs[104]) | (inputs[251]);
    assign layer0_outputs[9590] = ~(inputs[210]) | (inputs[163]);
    assign layer0_outputs[9591] = inputs[214];
    assign layer0_outputs[9592] = ~(inputs[146]);
    assign layer0_outputs[9593] = ~(inputs[117]) | (inputs[139]);
    assign layer0_outputs[9594] = ~((inputs[23]) ^ (inputs[231]));
    assign layer0_outputs[9595] = inputs[113];
    assign layer0_outputs[9596] = ~(inputs[22]);
    assign layer0_outputs[9597] = (inputs[195]) ^ (inputs[199]);
    assign layer0_outputs[9598] = 1'b0;
    assign layer0_outputs[9599] = (inputs[121]) ^ (inputs[231]);
    assign layer0_outputs[9600] = ~(inputs[39]);
    assign layer0_outputs[9601] = (inputs[40]) & ~(inputs[222]);
    assign layer0_outputs[9602] = (inputs[138]) & ~(inputs[179]);
    assign layer0_outputs[9603] = (inputs[94]) & ~(inputs[255]);
    assign layer0_outputs[9604] = ~(inputs[86]);
    assign layer0_outputs[9605] = inputs[19];
    assign layer0_outputs[9606] = ~((inputs[105]) | (inputs[62]));
    assign layer0_outputs[9607] = ~((inputs[56]) ^ (inputs[168]));
    assign layer0_outputs[9608] = (inputs[11]) | (inputs[108]);
    assign layer0_outputs[9609] = (inputs[20]) ^ (inputs[78]);
    assign layer0_outputs[9610] = ~(inputs[74]);
    assign layer0_outputs[9611] = ~((inputs[108]) ^ (inputs[6]));
    assign layer0_outputs[9612] = ~(inputs[39]);
    assign layer0_outputs[9613] = inputs[74];
    assign layer0_outputs[9614] = ~(inputs[237]) | (inputs[251]);
    assign layer0_outputs[9615] = (inputs[51]) ^ (inputs[98]);
    assign layer0_outputs[9616] = (inputs[85]) | (inputs[82]);
    assign layer0_outputs[9617] = (inputs[255]) | (inputs[122]);
    assign layer0_outputs[9618] = ~(inputs[163]);
    assign layer0_outputs[9619] = inputs[92];
    assign layer0_outputs[9620] = (inputs[64]) & (inputs[211]);
    assign layer0_outputs[9621] = ~((inputs[92]) ^ (inputs[32]));
    assign layer0_outputs[9622] = inputs[157];
    assign layer0_outputs[9623] = (inputs[162]) & ~(inputs[34]);
    assign layer0_outputs[9624] = ~((inputs[254]) | (inputs[201]));
    assign layer0_outputs[9625] = (inputs[29]) & ~(inputs[117]);
    assign layer0_outputs[9626] = (inputs[183]) & (inputs[185]);
    assign layer0_outputs[9627] = ~((inputs[169]) ^ (inputs[150]));
    assign layer0_outputs[9628] = ~((inputs[80]) ^ (inputs[19]));
    assign layer0_outputs[9629] = ~(inputs[229]);
    assign layer0_outputs[9630] = (inputs[27]) & ~(inputs[200]);
    assign layer0_outputs[9631] = ~(inputs[161]);
    assign layer0_outputs[9632] = ~(inputs[21]) | (inputs[160]);
    assign layer0_outputs[9633] = inputs[57];
    assign layer0_outputs[9634] = ~(inputs[144]);
    assign layer0_outputs[9635] = ~((inputs[87]) | (inputs[105]));
    assign layer0_outputs[9636] = inputs[147];
    assign layer0_outputs[9637] = ~((inputs[147]) | (inputs[208]));
    assign layer0_outputs[9638] = ~(inputs[135]);
    assign layer0_outputs[9639] = (inputs[215]) & ~(inputs[76]);
    assign layer0_outputs[9640] = (inputs[50]) ^ (inputs[238]);
    assign layer0_outputs[9641] = (inputs[16]) | (inputs[59]);
    assign layer0_outputs[9642] = inputs[217];
    assign layer0_outputs[9643] = inputs[68];
    assign layer0_outputs[9644] = ~((inputs[7]) ^ (inputs[88]));
    assign layer0_outputs[9645] = ~((inputs[180]) ^ (inputs[135]));
    assign layer0_outputs[9646] = (inputs[220]) | (inputs[186]);
    assign layer0_outputs[9647] = (inputs[8]) | (inputs[48]);
    assign layer0_outputs[9648] = ~(inputs[161]) | (inputs[47]);
    assign layer0_outputs[9649] = inputs[73];
    assign layer0_outputs[9650] = ~(inputs[119]);
    assign layer0_outputs[9651] = ~((inputs[255]) | (inputs[31]));
    assign layer0_outputs[9652] = ~((inputs[28]) ^ (inputs[251]));
    assign layer0_outputs[9653] = ~(inputs[220]);
    assign layer0_outputs[9654] = inputs[101];
    assign layer0_outputs[9655] = (inputs[112]) | (inputs[183]);
    assign layer0_outputs[9656] = (inputs[3]) & ~(inputs[53]);
    assign layer0_outputs[9657] = ~(inputs[104]) | (inputs[212]);
    assign layer0_outputs[9658] = (inputs[253]) | (inputs[232]);
    assign layer0_outputs[9659] = (inputs[64]) | (inputs[152]);
    assign layer0_outputs[9660] = inputs[44];
    assign layer0_outputs[9661] = ~((inputs[185]) | (inputs[187]));
    assign layer0_outputs[9662] = (inputs[97]) ^ (inputs[74]);
    assign layer0_outputs[9663] = inputs[26];
    assign layer0_outputs[9664] = ~(inputs[117]);
    assign layer0_outputs[9665] = ~((inputs[58]) | (inputs[24]));
    assign layer0_outputs[9666] = (inputs[37]) & ~(inputs[237]);
    assign layer0_outputs[9667] = ~((inputs[251]) | (inputs[252]));
    assign layer0_outputs[9668] = (inputs[159]) & ~(inputs[111]);
    assign layer0_outputs[9669] = ~(inputs[82]) | (inputs[16]);
    assign layer0_outputs[9670] = inputs[37];
    assign layer0_outputs[9671] = (inputs[243]) | (inputs[98]);
    assign layer0_outputs[9672] = ~((inputs[35]) & (inputs[36]));
    assign layer0_outputs[9673] = (inputs[237]) & ~(inputs[143]);
    assign layer0_outputs[9674] = (inputs[231]) & ~(inputs[41]);
    assign layer0_outputs[9675] = inputs[185];
    assign layer0_outputs[9676] = ~((inputs[246]) & (inputs[75]));
    assign layer0_outputs[9677] = ~((inputs[8]) | (inputs[174]));
    assign layer0_outputs[9678] = ~((inputs[207]) | (inputs[200]));
    assign layer0_outputs[9679] = (inputs[249]) | (inputs[114]);
    assign layer0_outputs[9680] = ~((inputs[36]) ^ (inputs[92]));
    assign layer0_outputs[9681] = inputs[23];
    assign layer0_outputs[9682] = (inputs[252]) | (inputs[164]);
    assign layer0_outputs[9683] = ~(inputs[168]) | (inputs[24]);
    assign layer0_outputs[9684] = inputs[124];
    assign layer0_outputs[9685] = (inputs[253]) | (inputs[133]);
    assign layer0_outputs[9686] = ~((inputs[10]) | (inputs[5]));
    assign layer0_outputs[9687] = ~(inputs[162]) | (inputs[96]);
    assign layer0_outputs[9688] = ~(inputs[167]);
    assign layer0_outputs[9689] = inputs[180];
    assign layer0_outputs[9690] = ~(inputs[203]);
    assign layer0_outputs[9691] = ~((inputs[21]) & (inputs[113]));
    assign layer0_outputs[9692] = inputs[107];
    assign layer0_outputs[9693] = inputs[230];
    assign layer0_outputs[9694] = (inputs[5]) & ~(inputs[0]);
    assign layer0_outputs[9695] = (inputs[7]) & ~(inputs[147]);
    assign layer0_outputs[9696] = ~((inputs[137]) ^ (inputs[119]));
    assign layer0_outputs[9697] = inputs[35];
    assign layer0_outputs[9698] = ~(inputs[180]) | (inputs[33]);
    assign layer0_outputs[9699] = ~((inputs[24]) & (inputs[90]));
    assign layer0_outputs[9700] = (inputs[162]) ^ (inputs[147]);
    assign layer0_outputs[9701] = inputs[59];
    assign layer0_outputs[9702] = inputs[44];
    assign layer0_outputs[9703] = ~(inputs[226]);
    assign layer0_outputs[9704] = ~(inputs[183]) | (inputs[133]);
    assign layer0_outputs[9705] = ~((inputs[62]) | (inputs[214]));
    assign layer0_outputs[9706] = (inputs[4]) ^ (inputs[101]);
    assign layer0_outputs[9707] = inputs[166];
    assign layer0_outputs[9708] = ~(inputs[188]) | (inputs[47]);
    assign layer0_outputs[9709] = inputs[9];
    assign layer0_outputs[9710] = (inputs[1]) ^ (inputs[136]);
    assign layer0_outputs[9711] = ~(inputs[17]);
    assign layer0_outputs[9712] = ~(inputs[198]) | (inputs[191]);
    assign layer0_outputs[9713] = ~(inputs[162]);
    assign layer0_outputs[9714] = 1'b1;
    assign layer0_outputs[9715] = (inputs[215]) & ~(inputs[254]);
    assign layer0_outputs[9716] = ~(inputs[79]);
    assign layer0_outputs[9717] = ~(inputs[18]);
    assign layer0_outputs[9718] = ~(inputs[27]);
    assign layer0_outputs[9719] = inputs[117];
    assign layer0_outputs[9720] = inputs[104];
    assign layer0_outputs[9721] = ~(inputs[221]);
    assign layer0_outputs[9722] = ~((inputs[40]) | (inputs[174]));
    assign layer0_outputs[9723] = ~((inputs[2]) & (inputs[109]));
    assign layer0_outputs[9724] = inputs[126];
    assign layer0_outputs[9725] = ~(inputs[141]);
    assign layer0_outputs[9726] = (inputs[38]) | (inputs[212]);
    assign layer0_outputs[9727] = (inputs[49]) | (inputs[231]);
    assign layer0_outputs[9728] = (inputs[92]) & ~(inputs[179]);
    assign layer0_outputs[9729] = ~((inputs[50]) ^ (inputs[47]));
    assign layer0_outputs[9730] = ~(inputs[41]) | (inputs[164]);
    assign layer0_outputs[9731] = (inputs[166]) | (inputs[149]);
    assign layer0_outputs[9732] = ~(inputs[236]);
    assign layer0_outputs[9733] = (inputs[22]) & (inputs[228]);
    assign layer0_outputs[9734] = ~(inputs[182]);
    assign layer0_outputs[9735] = (inputs[89]) ^ (inputs[107]);
    assign layer0_outputs[9736] = (inputs[242]) | (inputs[176]);
    assign layer0_outputs[9737] = (inputs[8]) & ~(inputs[128]);
    assign layer0_outputs[9738] = (inputs[180]) & ~(inputs[159]);
    assign layer0_outputs[9739] = ~(inputs[236]) | (inputs[139]);
    assign layer0_outputs[9740] = ~((inputs[199]) | (inputs[252]));
    assign layer0_outputs[9741] = ~(inputs[200]);
    assign layer0_outputs[9742] = inputs[130];
    assign layer0_outputs[9743] = inputs[158];
    assign layer0_outputs[9744] = ~(inputs[178]);
    assign layer0_outputs[9745] = ~((inputs[118]) | (inputs[225]));
    assign layer0_outputs[9746] = 1'b1;
    assign layer0_outputs[9747] = (inputs[140]) & ~(inputs[237]);
    assign layer0_outputs[9748] = ~(inputs[98]) | (inputs[123]);
    assign layer0_outputs[9749] = (inputs[232]) & ~(inputs[64]);
    assign layer0_outputs[9750] = ~((inputs[185]) ^ (inputs[134]));
    assign layer0_outputs[9751] = (inputs[171]) & ~(inputs[45]);
    assign layer0_outputs[9752] = ~((inputs[173]) ^ (inputs[187]));
    assign layer0_outputs[9753] = (inputs[150]) | (inputs[83]);
    assign layer0_outputs[9754] = (inputs[225]) | (inputs[148]);
    assign layer0_outputs[9755] = inputs[198];
    assign layer0_outputs[9756] = (inputs[7]) | (inputs[204]);
    assign layer0_outputs[9757] = ~((inputs[156]) | (inputs[145]));
    assign layer0_outputs[9758] = ~((inputs[75]) | (inputs[21]));
    assign layer0_outputs[9759] = inputs[163];
    assign layer0_outputs[9760] = inputs[231];
    assign layer0_outputs[9761] = ~((inputs[221]) ^ (inputs[249]));
    assign layer0_outputs[9762] = ~((inputs[62]) | (inputs[48]));
    assign layer0_outputs[9763] = ~(inputs[163]) | (inputs[74]);
    assign layer0_outputs[9764] = ~(inputs[36]) | (inputs[216]);
    assign layer0_outputs[9765] = (inputs[190]) ^ (inputs[32]);
    assign layer0_outputs[9766] = (inputs[235]) | (inputs[251]);
    assign layer0_outputs[9767] = ~((inputs[127]) | (inputs[219]));
    assign layer0_outputs[9768] = inputs[81];
    assign layer0_outputs[9769] = inputs[132];
    assign layer0_outputs[9770] = (inputs[146]) ^ (inputs[238]);
    assign layer0_outputs[9771] = (inputs[18]) | (inputs[181]);
    assign layer0_outputs[9772] = ~((inputs[11]) ^ (inputs[31]));
    assign layer0_outputs[9773] = (inputs[46]) | (inputs[177]);
    assign layer0_outputs[9774] = inputs[59];
    assign layer0_outputs[9775] = inputs[27];
    assign layer0_outputs[9776] = ~(inputs[237]) | (inputs[241]);
    assign layer0_outputs[9777] = ~(inputs[27]) | (inputs[163]);
    assign layer0_outputs[9778] = ~(inputs[226]) | (inputs[120]);
    assign layer0_outputs[9779] = inputs[81];
    assign layer0_outputs[9780] = inputs[88];
    assign layer0_outputs[9781] = (inputs[103]) & ~(inputs[206]);
    assign layer0_outputs[9782] = (inputs[66]) | (inputs[163]);
    assign layer0_outputs[9783] = (inputs[89]) ^ (inputs[222]);
    assign layer0_outputs[9784] = ~(inputs[229]);
    assign layer0_outputs[9785] = (inputs[158]) & (inputs[189]);
    assign layer0_outputs[9786] = (inputs[246]) | (inputs[128]);
    assign layer0_outputs[9787] = (inputs[12]) & ~(inputs[157]);
    assign layer0_outputs[9788] = (inputs[126]) & ~(inputs[219]);
    assign layer0_outputs[9789] = ~((inputs[82]) ^ (inputs[85]));
    assign layer0_outputs[9790] = ~(inputs[105]) | (inputs[22]);
    assign layer0_outputs[9791] = ~(inputs[186]) | (inputs[43]);
    assign layer0_outputs[9792] = inputs[25];
    assign layer0_outputs[9793] = (inputs[132]) | (inputs[246]);
    assign layer0_outputs[9794] = ~(inputs[172]);
    assign layer0_outputs[9795] = ~(inputs[241]);
    assign layer0_outputs[9796] = ~(inputs[173]);
    assign layer0_outputs[9797] = ~(inputs[153]);
    assign layer0_outputs[9798] = (inputs[152]) | (inputs[144]);
    assign layer0_outputs[9799] = ~((inputs[128]) & (inputs[143]));
    assign layer0_outputs[9800] = ~(inputs[248]);
    assign layer0_outputs[9801] = inputs[186];
    assign layer0_outputs[9802] = ~(inputs[63]);
    assign layer0_outputs[9803] = ~(inputs[229]) | (inputs[175]);
    assign layer0_outputs[9804] = ~(inputs[210]) | (inputs[239]);
    assign layer0_outputs[9805] = ~((inputs[121]) | (inputs[106]));
    assign layer0_outputs[9806] = inputs[163];
    assign layer0_outputs[9807] = inputs[231];
    assign layer0_outputs[9808] = ~(inputs[111]);
    assign layer0_outputs[9809] = ~(inputs[74]) | (inputs[164]);
    assign layer0_outputs[9810] = inputs[75];
    assign layer0_outputs[9811] = (inputs[87]) | (inputs[242]);
    assign layer0_outputs[9812] = (inputs[160]) | (inputs[38]);
    assign layer0_outputs[9813] = ~((inputs[216]) ^ (inputs[111]));
    assign layer0_outputs[9814] = ~((inputs[155]) ^ (inputs[198]));
    assign layer0_outputs[9815] = inputs[181];
    assign layer0_outputs[9816] = ~(inputs[165]);
    assign layer0_outputs[9817] = ~(inputs[142]);
    assign layer0_outputs[9818] = ~((inputs[117]) & (inputs[201]));
    assign layer0_outputs[9819] = ~(inputs[227]);
    assign layer0_outputs[9820] = ~((inputs[24]) ^ (inputs[21]));
    assign layer0_outputs[9821] = (inputs[207]) ^ (inputs[77]);
    assign layer0_outputs[9822] = ~((inputs[194]) | (inputs[175]));
    assign layer0_outputs[9823] = ~(inputs[46]);
    assign layer0_outputs[9824] = ~(inputs[39]) | (inputs[26]);
    assign layer0_outputs[9825] = (inputs[141]) & (inputs[235]);
    assign layer0_outputs[9826] = ~((inputs[4]) ^ (inputs[254]));
    assign layer0_outputs[9827] = ~((inputs[102]) ^ (inputs[175]));
    assign layer0_outputs[9828] = (inputs[37]) & ~(inputs[220]);
    assign layer0_outputs[9829] = (inputs[88]) ^ (inputs[23]);
    assign layer0_outputs[9830] = (inputs[110]) & ~(inputs[136]);
    assign layer0_outputs[9831] = ~(inputs[202]);
    assign layer0_outputs[9832] = ~(inputs[86]);
    assign layer0_outputs[9833] = (inputs[164]) | (inputs[80]);
    assign layer0_outputs[9834] = (inputs[177]) | (inputs[81]);
    assign layer0_outputs[9835] = inputs[57];
    assign layer0_outputs[9836] = ~((inputs[70]) & (inputs[214]));
    assign layer0_outputs[9837] = (inputs[63]) | (inputs[226]);
    assign layer0_outputs[9838] = (inputs[141]) & ~(inputs[155]);
    assign layer0_outputs[9839] = ~((inputs[195]) | (inputs[68]));
    assign layer0_outputs[9840] = ~(inputs[75]) | (inputs[34]);
    assign layer0_outputs[9841] = ~(inputs[78]);
    assign layer0_outputs[9842] = inputs[214];
    assign layer0_outputs[9843] = (inputs[228]) ^ (inputs[143]);
    assign layer0_outputs[9844] = inputs[76];
    assign layer0_outputs[9845] = (inputs[228]) & ~(inputs[5]);
    assign layer0_outputs[9846] = inputs[26];
    assign layer0_outputs[9847] = (inputs[108]) | (inputs[9]);
    assign layer0_outputs[9848] = inputs[121];
    assign layer0_outputs[9849] = (inputs[61]) | (inputs[197]);
    assign layer0_outputs[9850] = (inputs[112]) | (inputs[172]);
    assign layer0_outputs[9851] = ~((inputs[195]) & (inputs[10]));
    assign layer0_outputs[9852] = (inputs[176]) & ~(inputs[64]);
    assign layer0_outputs[9853] = ~(inputs[158]);
    assign layer0_outputs[9854] = (inputs[187]) | (inputs[88]);
    assign layer0_outputs[9855] = inputs[22];
    assign layer0_outputs[9856] = ~(inputs[108]);
    assign layer0_outputs[9857] = ~((inputs[150]) | (inputs[10]));
    assign layer0_outputs[9858] = ~((inputs[162]) | (inputs[146]));
    assign layer0_outputs[9859] = inputs[37];
    assign layer0_outputs[9860] = 1'b1;
    assign layer0_outputs[9861] = (inputs[87]) & (inputs[170]);
    assign layer0_outputs[9862] = (inputs[106]) & ~(inputs[158]);
    assign layer0_outputs[9863] = ~(inputs[82]) | (inputs[75]);
    assign layer0_outputs[9864] = ~(inputs[221]);
    assign layer0_outputs[9865] = (inputs[24]) & ~(inputs[236]);
    assign layer0_outputs[9866] = (inputs[242]) ^ (inputs[180]);
    assign layer0_outputs[9867] = ~(inputs[103]);
    assign layer0_outputs[9868] = ~((inputs[221]) | (inputs[192]));
    assign layer0_outputs[9869] = inputs[233];
    assign layer0_outputs[9870] = ~((inputs[129]) ^ (inputs[102]));
    assign layer0_outputs[9871] = ~(inputs[100]);
    assign layer0_outputs[9872] = ~(inputs[218]);
    assign layer0_outputs[9873] = inputs[117];
    assign layer0_outputs[9874] = (inputs[178]) | (inputs[159]);
    assign layer0_outputs[9875] = (inputs[247]) & ~(inputs[106]);
    assign layer0_outputs[9876] = ~(inputs[186]);
    assign layer0_outputs[9877] = ~(inputs[85]);
    assign layer0_outputs[9878] = (inputs[166]) & ~(inputs[176]);
    assign layer0_outputs[9879] = (inputs[86]) ^ (inputs[36]);
    assign layer0_outputs[9880] = ~((inputs[65]) & (inputs[32]));
    assign layer0_outputs[9881] = (inputs[64]) ^ (inputs[161]);
    assign layer0_outputs[9882] = ~(inputs[35]) | (inputs[100]);
    assign layer0_outputs[9883] = (inputs[112]) | (inputs[97]);
    assign layer0_outputs[9884] = ~((inputs[171]) | (inputs[85]));
    assign layer0_outputs[9885] = ~((inputs[187]) ^ (inputs[101]));
    assign layer0_outputs[9886] = ~(inputs[142]);
    assign layer0_outputs[9887] = ~(inputs[119]);
    assign layer0_outputs[9888] = ~(inputs[150]);
    assign layer0_outputs[9889] = 1'b0;
    assign layer0_outputs[9890] = inputs[133];
    assign layer0_outputs[9891] = (inputs[193]) & ~(inputs[2]);
    assign layer0_outputs[9892] = ~(inputs[85]);
    assign layer0_outputs[9893] = ~(inputs[113]) | (inputs[4]);
    assign layer0_outputs[9894] = ~((inputs[191]) | (inputs[182]));
    assign layer0_outputs[9895] = ~((inputs[38]) & (inputs[99]));
    assign layer0_outputs[9896] = ~(inputs[93]) | (inputs[224]);
    assign layer0_outputs[9897] = ~((inputs[112]) & (inputs[128]));
    assign layer0_outputs[9898] = inputs[16];
    assign layer0_outputs[9899] = inputs[8];
    assign layer0_outputs[9900] = (inputs[136]) & ~(inputs[96]);
    assign layer0_outputs[9901] = ~((inputs[237]) | (inputs[23]));
    assign layer0_outputs[9902] = inputs[124];
    assign layer0_outputs[9903] = ~((inputs[92]) ^ (inputs[79]));
    assign layer0_outputs[9904] = (inputs[122]) & ~(inputs[35]);
    assign layer0_outputs[9905] = (inputs[130]) ^ (inputs[103]);
    assign layer0_outputs[9906] = (inputs[63]) | (inputs[250]);
    assign layer0_outputs[9907] = inputs[177];
    assign layer0_outputs[9908] = inputs[59];
    assign layer0_outputs[9909] = (inputs[228]) | (inputs[51]);
    assign layer0_outputs[9910] = (inputs[27]) & ~(inputs[181]);
    assign layer0_outputs[9911] = ~(inputs[84]);
    assign layer0_outputs[9912] = (inputs[174]) ^ (inputs[133]);
    assign layer0_outputs[9913] = inputs[14];
    assign layer0_outputs[9914] = ~(inputs[213]);
    assign layer0_outputs[9915] = inputs[211];
    assign layer0_outputs[9916] = ~((inputs[96]) ^ (inputs[42]));
    assign layer0_outputs[9917] = ~((inputs[242]) | (inputs[248]));
    assign layer0_outputs[9918] = inputs[162];
    assign layer0_outputs[9919] = inputs[196];
    assign layer0_outputs[9920] = ~(inputs[238]) | (inputs[209]);
    assign layer0_outputs[9921] = inputs[248];
    assign layer0_outputs[9922] = ~((inputs[174]) | (inputs[61]));
    assign layer0_outputs[9923] = (inputs[144]) ^ (inputs[1]);
    assign layer0_outputs[9924] = ~(inputs[152]);
    assign layer0_outputs[9925] = ~(inputs[231]);
    assign layer0_outputs[9926] = ~(inputs[246]);
    assign layer0_outputs[9927] = (inputs[230]) & ~(inputs[146]);
    assign layer0_outputs[9928] = ~(inputs[231]);
    assign layer0_outputs[9929] = (inputs[57]) | (inputs[193]);
    assign layer0_outputs[9930] = inputs[143];
    assign layer0_outputs[9931] = (inputs[14]) ^ (inputs[183]);
    assign layer0_outputs[9932] = (inputs[142]) & (inputs[82]);
    assign layer0_outputs[9933] = (inputs[89]) ^ (inputs[209]);
    assign layer0_outputs[9934] = ~(inputs[20]);
    assign layer0_outputs[9935] = ~((inputs[25]) ^ (inputs[80]));
    assign layer0_outputs[9936] = (inputs[95]) & ~(inputs[135]);
    assign layer0_outputs[9937] = ~(inputs[179]) | (inputs[212]);
    assign layer0_outputs[9938] = 1'b0;
    assign layer0_outputs[9939] = ~(inputs[230]);
    assign layer0_outputs[9940] = (inputs[99]) | (inputs[14]);
    assign layer0_outputs[9941] = (inputs[178]) ^ (inputs[188]);
    assign layer0_outputs[9942] = (inputs[91]) & (inputs[30]);
    assign layer0_outputs[9943] = ~((inputs[171]) & (inputs[228]));
    assign layer0_outputs[9944] = (inputs[89]) & ~(inputs[202]);
    assign layer0_outputs[9945] = inputs[174];
    assign layer0_outputs[9946] = ~(inputs[202]);
    assign layer0_outputs[9947] = ~(inputs[153]);
    assign layer0_outputs[9948] = ~(inputs[120]) | (inputs[32]);
    assign layer0_outputs[9949] = (inputs[158]) | (inputs[19]);
    assign layer0_outputs[9950] = (inputs[138]) | (inputs[15]);
    assign layer0_outputs[9951] = ~(inputs[199]) | (inputs[76]);
    assign layer0_outputs[9952] = (inputs[63]) | (inputs[142]);
    assign layer0_outputs[9953] = (inputs[7]) | (inputs[60]);
    assign layer0_outputs[9954] = inputs[10];
    assign layer0_outputs[9955] = inputs[122];
    assign layer0_outputs[9956] = (inputs[196]) & ~(inputs[61]);
    assign layer0_outputs[9957] = (inputs[46]) & ~(inputs[188]);
    assign layer0_outputs[9958] = (inputs[239]) | (inputs[200]);
    assign layer0_outputs[9959] = ~(inputs[43]);
    assign layer0_outputs[9960] = ~(inputs[201]) | (inputs[27]);
    assign layer0_outputs[9961] = (inputs[232]) & ~(inputs[255]);
    assign layer0_outputs[9962] = ~(inputs[30]) | (inputs[254]);
    assign layer0_outputs[9963] = inputs[87];
    assign layer0_outputs[9964] = ~((inputs[93]) ^ (inputs[2]));
    assign layer0_outputs[9965] = inputs[23];
    assign layer0_outputs[9966] = (inputs[34]) | (inputs[255]);
    assign layer0_outputs[9967] = (inputs[216]) ^ (inputs[189]);
    assign layer0_outputs[9968] = (inputs[89]) & ~(inputs[192]);
    assign layer0_outputs[9969] = ~((inputs[160]) ^ (inputs[131]));
    assign layer0_outputs[9970] = ~((inputs[102]) | (inputs[101]));
    assign layer0_outputs[9971] = ~(inputs[2]);
    assign layer0_outputs[9972] = (inputs[111]) ^ (inputs[76]);
    assign layer0_outputs[9973] = ~(inputs[150]) | (inputs[73]);
    assign layer0_outputs[9974] = ~(inputs[33]);
    assign layer0_outputs[9975] = inputs[34];
    assign layer0_outputs[9976] = (inputs[93]) ^ (inputs[233]);
    assign layer0_outputs[9977] = (inputs[180]) ^ (inputs[88]);
    assign layer0_outputs[9978] = inputs[243];
    assign layer0_outputs[9979] = ~(inputs[203]);
    assign layer0_outputs[9980] = ~(inputs[232]);
    assign layer0_outputs[9981] = ~(inputs[68]);
    assign layer0_outputs[9982] = ~((inputs[16]) | (inputs[160]));
    assign layer0_outputs[9983] = ~(inputs[134]) | (inputs[14]);
    assign layer0_outputs[9984] = (inputs[90]) & ~(inputs[118]);
    assign layer0_outputs[9985] = (inputs[32]) ^ (inputs[60]);
    assign layer0_outputs[9986] = inputs[41];
    assign layer0_outputs[9987] = ~(inputs[50]) | (inputs[167]);
    assign layer0_outputs[9988] = ~((inputs[184]) | (inputs[184]));
    assign layer0_outputs[9989] = (inputs[218]) & ~(inputs[63]);
    assign layer0_outputs[9990] = ~((inputs[65]) | (inputs[29]));
    assign layer0_outputs[9991] = ~(inputs[179]) | (inputs[55]);
    assign layer0_outputs[9992] = ~(inputs[104]);
    assign layer0_outputs[9993] = (inputs[147]) ^ (inputs[153]);
    assign layer0_outputs[9994] = ~(inputs[52]) | (inputs[72]);
    assign layer0_outputs[9995] = ~(inputs[89]);
    assign layer0_outputs[9996] = ~(inputs[26]) | (inputs[219]);
    assign layer0_outputs[9997] = ~((inputs[113]) | (inputs[163]));
    assign layer0_outputs[9998] = ~(inputs[6]);
    assign layer0_outputs[9999] = (inputs[239]) & ~(inputs[46]);
    assign layer0_outputs[10000] = ~(inputs[139]) | (inputs[73]);
    assign layer0_outputs[10001] = ~(inputs[71]);
    assign layer0_outputs[10002] = ~(inputs[157]) | (inputs[182]);
    assign layer0_outputs[10003] = ~(inputs[121]) | (inputs[156]);
    assign layer0_outputs[10004] = inputs[18];
    assign layer0_outputs[10005] = ~(inputs[212]);
    assign layer0_outputs[10006] = (inputs[177]) ^ (inputs[92]);
    assign layer0_outputs[10007] = ~(inputs[164]);
    assign layer0_outputs[10008] = (inputs[175]) & ~(inputs[72]);
    assign layer0_outputs[10009] = ~((inputs[21]) ^ (inputs[204]));
    assign layer0_outputs[10010] = ~(inputs[183]);
    assign layer0_outputs[10011] = ~(inputs[36]);
    assign layer0_outputs[10012] = (inputs[10]) | (inputs[1]);
    assign layer0_outputs[10013] = inputs[163];
    assign layer0_outputs[10014] = inputs[44];
    assign layer0_outputs[10015] = inputs[70];
    assign layer0_outputs[10016] = ~(inputs[175]);
    assign layer0_outputs[10017] = (inputs[155]) & ~(inputs[26]);
    assign layer0_outputs[10018] = (inputs[162]) & (inputs[249]);
    assign layer0_outputs[10019] = inputs[100];
    assign layer0_outputs[10020] = inputs[115];
    assign layer0_outputs[10021] = (inputs[94]) & (inputs[92]);
    assign layer0_outputs[10022] = (inputs[150]) | (inputs[204]);
    assign layer0_outputs[10023] = ~(inputs[142]);
    assign layer0_outputs[10024] = ~((inputs[47]) | (inputs[46]));
    assign layer0_outputs[10025] = (inputs[171]) | (inputs[208]);
    assign layer0_outputs[10026] = inputs[194];
    assign layer0_outputs[10027] = ~(inputs[154]);
    assign layer0_outputs[10028] = inputs[165];
    assign layer0_outputs[10029] = inputs[122];
    assign layer0_outputs[10030] = inputs[215];
    assign layer0_outputs[10031] = ~(inputs[114]);
    assign layer0_outputs[10032] = (inputs[187]) & ~(inputs[143]);
    assign layer0_outputs[10033] = ~((inputs[172]) | (inputs[79]));
    assign layer0_outputs[10034] = ~((inputs[109]) | (inputs[93]));
    assign layer0_outputs[10035] = (inputs[116]) & ~(inputs[4]);
    assign layer0_outputs[10036] = (inputs[172]) & ~(inputs[54]);
    assign layer0_outputs[10037] = (inputs[236]) | (inputs[173]);
    assign layer0_outputs[10038] = ~((inputs[22]) ^ (inputs[50]));
    assign layer0_outputs[10039] = (inputs[141]) & ~(inputs[5]);
    assign layer0_outputs[10040] = (inputs[165]) ^ (inputs[76]);
    assign layer0_outputs[10041] = (inputs[70]) ^ (inputs[34]);
    assign layer0_outputs[10042] = (inputs[0]) & ~(inputs[216]);
    assign layer0_outputs[10043] = ~((inputs[56]) ^ (inputs[30]));
    assign layer0_outputs[10044] = (inputs[171]) ^ (inputs[88]);
    assign layer0_outputs[10045] = ~(inputs[114]);
    assign layer0_outputs[10046] = ~(inputs[87]);
    assign layer0_outputs[10047] = ~(inputs[99]) | (inputs[15]);
    assign layer0_outputs[10048] = inputs[191];
    assign layer0_outputs[10049] = ~((inputs[74]) ^ (inputs[72]));
    assign layer0_outputs[10050] = (inputs[42]) ^ (inputs[118]);
    assign layer0_outputs[10051] = inputs[56];
    assign layer0_outputs[10052] = (inputs[239]) & ~(inputs[175]);
    assign layer0_outputs[10053] = inputs[99];
    assign layer0_outputs[10054] = (inputs[142]) | (inputs[217]);
    assign layer0_outputs[10055] = inputs[232];
    assign layer0_outputs[10056] = (inputs[108]) | (inputs[81]);
    assign layer0_outputs[10057] = inputs[5];
    assign layer0_outputs[10058] = (inputs[252]) ^ (inputs[127]);
    assign layer0_outputs[10059] = ~((inputs[127]) | (inputs[201]));
    assign layer0_outputs[10060] = inputs[133];
    assign layer0_outputs[10061] = (inputs[236]) | (inputs[196]);
    assign layer0_outputs[10062] = ~((inputs[4]) | (inputs[51]));
    assign layer0_outputs[10063] = ~(inputs[229]);
    assign layer0_outputs[10064] = (inputs[58]) | (inputs[97]);
    assign layer0_outputs[10065] = ~(inputs[87]) | (inputs[19]);
    assign layer0_outputs[10066] = 1'b1;
    assign layer0_outputs[10067] = ~((inputs[206]) ^ (inputs[7]));
    assign layer0_outputs[10068] = (inputs[210]) | (inputs[220]);
    assign layer0_outputs[10069] = 1'b0;
    assign layer0_outputs[10070] = inputs[216];
    assign layer0_outputs[10071] = (inputs[66]) & ~(inputs[107]);
    assign layer0_outputs[10072] = (inputs[195]) ^ (inputs[189]);
    assign layer0_outputs[10073] = inputs[98];
    assign layer0_outputs[10074] = ~(inputs[88]);
    assign layer0_outputs[10075] = inputs[103];
    assign layer0_outputs[10076] = inputs[151];
    assign layer0_outputs[10077] = (inputs[88]) & (inputs[8]);
    assign layer0_outputs[10078] = inputs[52];
    assign layer0_outputs[10079] = (inputs[66]) | (inputs[38]);
    assign layer0_outputs[10080] = ~((inputs[64]) ^ (inputs[112]));
    assign layer0_outputs[10081] = ~((inputs[192]) ^ (inputs[90]));
    assign layer0_outputs[10082] = inputs[66];
    assign layer0_outputs[10083] = (inputs[234]) & (inputs[41]);
    assign layer0_outputs[10084] = (inputs[74]) ^ (inputs[253]);
    assign layer0_outputs[10085] = (inputs[109]) | (inputs[78]);
    assign layer0_outputs[10086] = ~((inputs[179]) ^ (inputs[128]));
    assign layer0_outputs[10087] = (inputs[176]) | (inputs[141]);
    assign layer0_outputs[10088] = (inputs[42]) & ~(inputs[69]);
    assign layer0_outputs[10089] = ~((inputs[35]) | (inputs[243]));
    assign layer0_outputs[10090] = ~(inputs[12]) | (inputs[154]);
    assign layer0_outputs[10091] = ~((inputs[179]) | (inputs[188]));
    assign layer0_outputs[10092] = (inputs[69]) ^ (inputs[112]);
    assign layer0_outputs[10093] = ~((inputs[118]) | (inputs[205]));
    assign layer0_outputs[10094] = inputs[14];
    assign layer0_outputs[10095] = ~((inputs[86]) | (inputs[78]));
    assign layer0_outputs[10096] = inputs[41];
    assign layer0_outputs[10097] = (inputs[30]) | (inputs[182]);
    assign layer0_outputs[10098] = (inputs[72]) & (inputs[9]);
    assign layer0_outputs[10099] = inputs[102];
    assign layer0_outputs[10100] = ~(inputs[100]);
    assign layer0_outputs[10101] = (inputs[234]) | (inputs[217]);
    assign layer0_outputs[10102] = inputs[77];
    assign layer0_outputs[10103] = ~(inputs[120]);
    assign layer0_outputs[10104] = ~(inputs[162]);
    assign layer0_outputs[10105] = ~(inputs[54]);
    assign layer0_outputs[10106] = ~((inputs[150]) & (inputs[181]));
    assign layer0_outputs[10107] = ~((inputs[173]) ^ (inputs[194]));
    assign layer0_outputs[10108] = ~((inputs[43]) ^ (inputs[11]));
    assign layer0_outputs[10109] = ~((inputs[187]) ^ (inputs[116]));
    assign layer0_outputs[10110] = ~((inputs[197]) | (inputs[158]));
    assign layer0_outputs[10111] = inputs[197];
    assign layer0_outputs[10112] = ~(inputs[235]);
    assign layer0_outputs[10113] = ~(inputs[44]);
    assign layer0_outputs[10114] = ~((inputs[145]) | (inputs[116]));
    assign layer0_outputs[10115] = ~((inputs[196]) ^ (inputs[44]));
    assign layer0_outputs[10116] = ~((inputs[143]) ^ (inputs[139]));
    assign layer0_outputs[10117] = (inputs[204]) & (inputs[233]);
    assign layer0_outputs[10118] = inputs[5];
    assign layer0_outputs[10119] = ~((inputs[252]) ^ (inputs[83]));
    assign layer0_outputs[10120] = ~((inputs[51]) | (inputs[52]));
    assign layer0_outputs[10121] = ~(inputs[131]);
    assign layer0_outputs[10122] = ~((inputs[196]) | (inputs[220]));
    assign layer0_outputs[10123] = inputs[125];
    assign layer0_outputs[10124] = inputs[217];
    assign layer0_outputs[10125] = ~((inputs[81]) | (inputs[225]));
    assign layer0_outputs[10126] = (inputs[72]) ^ (inputs[67]);
    assign layer0_outputs[10127] = (inputs[35]) & (inputs[4]);
    assign layer0_outputs[10128] = ~(inputs[227]);
    assign layer0_outputs[10129] = ~(inputs[25]);
    assign layer0_outputs[10130] = inputs[104];
    assign layer0_outputs[10131] = ~(inputs[28]) | (inputs[193]);
    assign layer0_outputs[10132] = (inputs[57]) | (inputs[37]);
    assign layer0_outputs[10133] = inputs[23];
    assign layer0_outputs[10134] = (inputs[202]) & ~(inputs[37]);
    assign layer0_outputs[10135] = ~((inputs[193]) ^ (inputs[247]));
    assign layer0_outputs[10136] = inputs[144];
    assign layer0_outputs[10137] = (inputs[219]) & (inputs[131]);
    assign layer0_outputs[10138] = (inputs[95]) & ~(inputs[241]);
    assign layer0_outputs[10139] = ~(inputs[29]) | (inputs[144]);
    assign layer0_outputs[10140] = inputs[163];
    assign layer0_outputs[10141] = 1'b0;
    assign layer0_outputs[10142] = ~((inputs[131]) ^ (inputs[161]));
    assign layer0_outputs[10143] = ~(inputs[36]);
    assign layer0_outputs[10144] = (inputs[212]) & (inputs[162]);
    assign layer0_outputs[10145] = ~(inputs[153]);
    assign layer0_outputs[10146] = inputs[198];
    assign layer0_outputs[10147] = inputs[193];
    assign layer0_outputs[10148] = ~((inputs[193]) ^ (inputs[240]));
    assign layer0_outputs[10149] = ~(inputs[147]) | (inputs[208]);
    assign layer0_outputs[10150] = (inputs[204]) & ~(inputs[254]);
    assign layer0_outputs[10151] = (inputs[180]) & ~(inputs[1]);
    assign layer0_outputs[10152] = (inputs[5]) | (inputs[28]);
    assign layer0_outputs[10153] = (inputs[137]) & ~(inputs[18]);
    assign layer0_outputs[10154] = (inputs[132]) ^ (inputs[51]);
    assign layer0_outputs[10155] = inputs[120];
    assign layer0_outputs[10156] = ~((inputs[194]) ^ (inputs[65]));
    assign layer0_outputs[10157] = ~(inputs[26]);
    assign layer0_outputs[10158] = (inputs[131]) | (inputs[78]);
    assign layer0_outputs[10159] = (inputs[171]) ^ (inputs[19]);
    assign layer0_outputs[10160] = ~((inputs[207]) ^ (inputs[23]));
    assign layer0_outputs[10161] = ~((inputs[187]) & (inputs[202]));
    assign layer0_outputs[10162] = inputs[54];
    assign layer0_outputs[10163] = inputs[247];
    assign layer0_outputs[10164] = ~(inputs[7]) | (inputs[86]);
    assign layer0_outputs[10165] = ~((inputs[206]) | (inputs[190]));
    assign layer0_outputs[10166] = inputs[74];
    assign layer0_outputs[10167] = (inputs[248]) & ~(inputs[63]);
    assign layer0_outputs[10168] = (inputs[120]) & ~(inputs[165]);
    assign layer0_outputs[10169] = 1'b1;
    assign layer0_outputs[10170] = inputs[167];
    assign layer0_outputs[10171] = (inputs[46]) ^ (inputs[5]);
    assign layer0_outputs[10172] = ~(inputs[114]) | (inputs[191]);
    assign layer0_outputs[10173] = ~((inputs[38]) | (inputs[239]));
    assign layer0_outputs[10174] = inputs[13];
    assign layer0_outputs[10175] = ~((inputs[29]) | (inputs[225]));
    assign layer0_outputs[10176] = (inputs[42]) & (inputs[133]);
    assign layer0_outputs[10177] = (inputs[152]) | (inputs[124]);
    assign layer0_outputs[10178] = ~(inputs[115]);
    assign layer0_outputs[10179] = inputs[37];
    assign layer0_outputs[10180] = ~(inputs[22]);
    assign layer0_outputs[10181] = ~((inputs[248]) | (inputs[163]));
    assign layer0_outputs[10182] = ~(inputs[240]) | (inputs[78]);
    assign layer0_outputs[10183] = ~(inputs[1]);
    assign layer0_outputs[10184] = ~((inputs[126]) | (inputs[48]));
    assign layer0_outputs[10185] = inputs[25];
    assign layer0_outputs[10186] = inputs[54];
    assign layer0_outputs[10187] = inputs[249];
    assign layer0_outputs[10188] = (inputs[183]) | (inputs[237]);
    assign layer0_outputs[10189] = ~((inputs[140]) ^ (inputs[196]));
    assign layer0_outputs[10190] = (inputs[53]) ^ (inputs[34]);
    assign layer0_outputs[10191] = (inputs[243]) | (inputs[204]);
    assign layer0_outputs[10192] = ~((inputs[169]) ^ (inputs[129]));
    assign layer0_outputs[10193] = inputs[89];
    assign layer0_outputs[10194] = (inputs[172]) & ~(inputs[17]);
    assign layer0_outputs[10195] = inputs[8];
    assign layer0_outputs[10196] = ~((inputs[72]) | (inputs[64]));
    assign layer0_outputs[10197] = (inputs[128]) | (inputs[66]);
    assign layer0_outputs[10198] = ~((inputs[80]) | (inputs[118]));
    assign layer0_outputs[10199] = ~((inputs[236]) & (inputs[35]));
    assign layer0_outputs[10200] = inputs[87];
    assign layer0_outputs[10201] = (inputs[29]) & ~(inputs[226]);
    assign layer0_outputs[10202] = (inputs[186]) | (inputs[17]);
    assign layer0_outputs[10203] = inputs[69];
    assign layer0_outputs[10204] = ~(inputs[9]) | (inputs[143]);
    assign layer0_outputs[10205] = ~(inputs[254]);
    assign layer0_outputs[10206] = 1'b0;
    assign layer0_outputs[10207] = ~((inputs[67]) ^ (inputs[82]));
    assign layer0_outputs[10208] = ~(inputs[67]);
    assign layer0_outputs[10209] = (inputs[184]) | (inputs[165]);
    assign layer0_outputs[10210] = ~((inputs[206]) | (inputs[205]));
    assign layer0_outputs[10211] = (inputs[89]) & ~(inputs[250]);
    assign layer0_outputs[10212] = (inputs[222]) ^ (inputs[78]);
    assign layer0_outputs[10213] = ~(inputs[231]) | (inputs[30]);
    assign layer0_outputs[10214] = ~((inputs[28]) | (inputs[100]));
    assign layer0_outputs[10215] = ~(inputs[131]);
    assign layer0_outputs[10216] = ~(inputs[50]);
    assign layer0_outputs[10217] = inputs[104];
    assign layer0_outputs[10218] = ~((inputs[55]) ^ (inputs[114]));
    assign layer0_outputs[10219] = ~((inputs[4]) | (inputs[34]));
    assign layer0_outputs[10220] = ~(inputs[172]);
    assign layer0_outputs[10221] = ~((inputs[0]) ^ (inputs[50]));
    assign layer0_outputs[10222] = ~((inputs[158]) ^ (inputs[106]));
    assign layer0_outputs[10223] = (inputs[120]) & ~(inputs[9]);
    assign layer0_outputs[10224] = (inputs[105]) & ~(inputs[236]);
    assign layer0_outputs[10225] = (inputs[28]) & ~(inputs[254]);
    assign layer0_outputs[10226] = (inputs[191]) & ~(inputs[166]);
    assign layer0_outputs[10227] = ~(inputs[54]);
    assign layer0_outputs[10228] = ~(inputs[141]);
    assign layer0_outputs[10229] = (inputs[76]) | (inputs[135]);
    assign layer0_outputs[10230] = (inputs[127]) & ~(inputs[252]);
    assign layer0_outputs[10231] = ~((inputs[91]) | (inputs[108]));
    assign layer0_outputs[10232] = (inputs[103]) | (inputs[226]);
    assign layer0_outputs[10233] = ~((inputs[181]) | (inputs[1]));
    assign layer0_outputs[10234] = inputs[30];
    assign layer0_outputs[10235] = inputs[33];
    assign layer0_outputs[10236] = ~(inputs[216]);
    assign layer0_outputs[10237] = ~(inputs[100]);
    assign layer0_outputs[10238] = ~(inputs[79]) | (inputs[190]);
    assign layer0_outputs[10239] = (inputs[113]) & ~(inputs[111]);
    assign outputs[0] = (layer0_outputs[333]) | (layer0_outputs[2974]);
    assign outputs[1] = ~((layer0_outputs[2196]) ^ (layer0_outputs[3350]));
    assign outputs[2] = (layer0_outputs[7747]) & ~(layer0_outputs[509]);
    assign outputs[3] = (layer0_outputs[8588]) ^ (layer0_outputs[7564]);
    assign outputs[4] = (layer0_outputs[3872]) | (layer0_outputs[4473]);
    assign outputs[5] = ~(layer0_outputs[9435]);
    assign outputs[6] = ~(layer0_outputs[9013]);
    assign outputs[7] = ~((layer0_outputs[3640]) ^ (layer0_outputs[2189]));
    assign outputs[8] = ~(layer0_outputs[6306]);
    assign outputs[9] = (layer0_outputs[1357]) & ~(layer0_outputs[4129]);
    assign outputs[10] = ~(layer0_outputs[8901]);
    assign outputs[11] = ~((layer0_outputs[8460]) ^ (layer0_outputs[4558]));
    assign outputs[12] = ~(layer0_outputs[8481]);
    assign outputs[13] = ~((layer0_outputs[7550]) & (layer0_outputs[6540]));
    assign outputs[14] = ~((layer0_outputs[9425]) | (layer0_outputs[3900]));
    assign outputs[15] = layer0_outputs[782];
    assign outputs[16] = (layer0_outputs[7857]) & (layer0_outputs[295]);
    assign outputs[17] = ~(layer0_outputs[4773]);
    assign outputs[18] = layer0_outputs[1423];
    assign outputs[19] = 1'b0;
    assign outputs[20] = layer0_outputs[8422];
    assign outputs[21] = ~((layer0_outputs[2786]) | (layer0_outputs[2517]));
    assign outputs[22] = ~(layer0_outputs[2001]) | (layer0_outputs[8036]);
    assign outputs[23] = (layer0_outputs[231]) ^ (layer0_outputs[7443]);
    assign outputs[24] = ~(layer0_outputs[2970]) | (layer0_outputs[1334]);
    assign outputs[25] = ~(layer0_outputs[2939]);
    assign outputs[26] = (layer0_outputs[2005]) ^ (layer0_outputs[522]);
    assign outputs[27] = layer0_outputs[94];
    assign outputs[28] = ~(layer0_outputs[3334]);
    assign outputs[29] = ~((layer0_outputs[3425]) & (layer0_outputs[9840]));
    assign outputs[30] = layer0_outputs[7195];
    assign outputs[31] = ~(layer0_outputs[1665]) | (layer0_outputs[8291]);
    assign outputs[32] = ~((layer0_outputs[8754]) ^ (layer0_outputs[8451]));
    assign outputs[33] = ~(layer0_outputs[4773]);
    assign outputs[34] = layer0_outputs[4903];
    assign outputs[35] = layer0_outputs[4516];
    assign outputs[36] = ~(layer0_outputs[3773]);
    assign outputs[37] = ~(layer0_outputs[509]);
    assign outputs[38] = (layer0_outputs[4053]) ^ (layer0_outputs[1413]);
    assign outputs[39] = ~(layer0_outputs[9208]);
    assign outputs[40] = (layer0_outputs[9364]) & ~(layer0_outputs[4620]);
    assign outputs[41] = ~((layer0_outputs[1707]) ^ (layer0_outputs[6345]));
    assign outputs[42] = ~((layer0_outputs[3209]) ^ (layer0_outputs[1279]));
    assign outputs[43] = layer0_outputs[4505];
    assign outputs[44] = ~(layer0_outputs[6587]);
    assign outputs[45] = layer0_outputs[2515];
    assign outputs[46] = ~(layer0_outputs[5944]);
    assign outputs[47] = ~(layer0_outputs[1537]);
    assign outputs[48] = ~(layer0_outputs[9371]) | (layer0_outputs[9227]);
    assign outputs[49] = layer0_outputs[2131];
    assign outputs[50] = ~((layer0_outputs[1445]) ^ (layer0_outputs[4328]));
    assign outputs[51] = (layer0_outputs[8993]) & ~(layer0_outputs[4272]);
    assign outputs[52] = (layer0_outputs[9971]) ^ (layer0_outputs[1956]);
    assign outputs[53] = ~(layer0_outputs[9032]);
    assign outputs[54] = (layer0_outputs[1198]) | (layer0_outputs[7892]);
    assign outputs[55] = ~(layer0_outputs[6150]);
    assign outputs[56] = layer0_outputs[3528];
    assign outputs[57] = layer0_outputs[426];
    assign outputs[58] = ~((layer0_outputs[1425]) | (layer0_outputs[3626]));
    assign outputs[59] = ~((layer0_outputs[5377]) ^ (layer0_outputs[837]));
    assign outputs[60] = (layer0_outputs[3616]) | (layer0_outputs[9559]);
    assign outputs[61] = ~(layer0_outputs[6219]);
    assign outputs[62] = ~(layer0_outputs[7298]) | (layer0_outputs[9331]);
    assign outputs[63] = (layer0_outputs[7768]) | (layer0_outputs[3435]);
    assign outputs[64] = ~(layer0_outputs[8659]);
    assign outputs[65] = layer0_outputs[1988];
    assign outputs[66] = (layer0_outputs[7912]) ^ (layer0_outputs[1022]);
    assign outputs[67] = (layer0_outputs[9408]) | (layer0_outputs[7864]);
    assign outputs[68] = (layer0_outputs[6324]) ^ (layer0_outputs[4377]);
    assign outputs[69] = (layer0_outputs[3335]) & ~(layer0_outputs[6783]);
    assign outputs[70] = layer0_outputs[1768];
    assign outputs[71] = ~((layer0_outputs[6070]) & (layer0_outputs[7861]));
    assign outputs[72] = layer0_outputs[6214];
    assign outputs[73] = layer0_outputs[10159];
    assign outputs[74] = (layer0_outputs[5520]) | (layer0_outputs[1967]);
    assign outputs[75] = (layer0_outputs[5067]) | (layer0_outputs[2147]);
    assign outputs[76] = layer0_outputs[7441];
    assign outputs[77] = ~(layer0_outputs[2347]);
    assign outputs[78] = ~(layer0_outputs[6868]);
    assign outputs[79] = (layer0_outputs[8328]) ^ (layer0_outputs[1933]);
    assign outputs[80] = ~(layer0_outputs[4373]);
    assign outputs[81] = ~(layer0_outputs[6199]);
    assign outputs[82] = 1'b1;
    assign outputs[83] = ~(layer0_outputs[7540]);
    assign outputs[84] = (layer0_outputs[969]) & ~(layer0_outputs[368]);
    assign outputs[85] = (layer0_outputs[8749]) ^ (layer0_outputs[672]);
    assign outputs[86] = layer0_outputs[3174];
    assign outputs[87] = ~((layer0_outputs[3744]) ^ (layer0_outputs[8174]));
    assign outputs[88] = layer0_outputs[9443];
    assign outputs[89] = ~(layer0_outputs[3378]);
    assign outputs[90] = layer0_outputs[7644];
    assign outputs[91] = ~(layer0_outputs[9323]) | (layer0_outputs[4880]);
    assign outputs[92] = (layer0_outputs[553]) | (layer0_outputs[7642]);
    assign outputs[93] = layer0_outputs[8070];
    assign outputs[94] = ~(layer0_outputs[2247]);
    assign outputs[95] = layer0_outputs[6178];
    assign outputs[96] = ~((layer0_outputs[3941]) ^ (layer0_outputs[6161]));
    assign outputs[97] = ~(layer0_outputs[7121]) | (layer0_outputs[3926]);
    assign outputs[98] = layer0_outputs[6850];
    assign outputs[99] = (layer0_outputs[3299]) ^ (layer0_outputs[7886]);
    assign outputs[100] = layer0_outputs[10096];
    assign outputs[101] = ~(layer0_outputs[7444]);
    assign outputs[102] = ~((layer0_outputs[2991]) ^ (layer0_outputs[7837]));
    assign outputs[103] = layer0_outputs[1241];
    assign outputs[104] = layer0_outputs[7261];
    assign outputs[105] = ~(layer0_outputs[396]);
    assign outputs[106] = ~(layer0_outputs[5837]);
    assign outputs[107] = layer0_outputs[6110];
    assign outputs[108] = ~((layer0_outputs[2948]) ^ (layer0_outputs[8532]));
    assign outputs[109] = layer0_outputs[4975];
    assign outputs[110] = ~(layer0_outputs[6395]);
    assign outputs[111] = layer0_outputs[542];
    assign outputs[112] = (layer0_outputs[6720]) & (layer0_outputs[4718]);
    assign outputs[113] = layer0_outputs[8761];
    assign outputs[114] = (layer0_outputs[10165]) & ~(layer0_outputs[5990]);
    assign outputs[115] = ~(layer0_outputs[8164]);
    assign outputs[116] = ~(layer0_outputs[2671]);
    assign outputs[117] = ~(layer0_outputs[2165]);
    assign outputs[118] = ~(layer0_outputs[3978]);
    assign outputs[119] = layer0_outputs[6508];
    assign outputs[120] = ~(layer0_outputs[4030]);
    assign outputs[121] = ~((layer0_outputs[9682]) ^ (layer0_outputs[4113]));
    assign outputs[122] = layer0_outputs[9770];
    assign outputs[123] = ~(layer0_outputs[3615]);
    assign outputs[124] = ~(layer0_outputs[9997]);
    assign outputs[125] = layer0_outputs[1686];
    assign outputs[126] = ~(layer0_outputs[5947]);
    assign outputs[127] = ~((layer0_outputs[4754]) & (layer0_outputs[4318]));
    assign outputs[128] = layer0_outputs[9688];
    assign outputs[129] = ~(layer0_outputs[9548]);
    assign outputs[130] = layer0_outputs[6673];
    assign outputs[131] = ~(layer0_outputs[1874]);
    assign outputs[132] = (layer0_outputs[916]) & (layer0_outputs[7753]);
    assign outputs[133] = (layer0_outputs[9505]) & ~(layer0_outputs[8018]);
    assign outputs[134] = (layer0_outputs[9723]) & ~(layer0_outputs[9702]);
    assign outputs[135] = ~((layer0_outputs[4501]) & (layer0_outputs[5565]));
    assign outputs[136] = layer0_outputs[4092];
    assign outputs[137] = ~(layer0_outputs[4817]);
    assign outputs[138] = layer0_outputs[5938];
    assign outputs[139] = ~((layer0_outputs[9129]) & (layer0_outputs[6509]));
    assign outputs[140] = layer0_outputs[3999];
    assign outputs[141] = (layer0_outputs[7406]) ^ (layer0_outputs[2104]);
    assign outputs[142] = (layer0_outputs[9611]) ^ (layer0_outputs[8909]);
    assign outputs[143] = (layer0_outputs[9849]) | (layer0_outputs[7046]);
    assign outputs[144] = ~((layer0_outputs[880]) & (layer0_outputs[8685]));
    assign outputs[145] = (layer0_outputs[7504]) | (layer0_outputs[7315]);
    assign outputs[146] = (layer0_outputs[2841]) & (layer0_outputs[2581]);
    assign outputs[147] = layer0_outputs[690];
    assign outputs[148] = (layer0_outputs[3991]) ^ (layer0_outputs[8479]);
    assign outputs[149] = ~(layer0_outputs[5516]);
    assign outputs[150] = (layer0_outputs[7778]) | (layer0_outputs[9485]);
    assign outputs[151] = (layer0_outputs[1368]) & ~(layer0_outputs[10097]);
    assign outputs[152] = (layer0_outputs[8508]) ^ (layer0_outputs[79]);
    assign outputs[153] = (layer0_outputs[5707]) | (layer0_outputs[4887]);
    assign outputs[154] = (layer0_outputs[2653]) & (layer0_outputs[431]);
    assign outputs[155] = layer0_outputs[7083];
    assign outputs[156] = (layer0_outputs[9804]) ^ (layer0_outputs[157]);
    assign outputs[157] = ~(layer0_outputs[1020]) | (layer0_outputs[7294]);
    assign outputs[158] = ~((layer0_outputs[641]) | (layer0_outputs[3743]));
    assign outputs[159] = ~(layer0_outputs[4507]);
    assign outputs[160] = ~((layer0_outputs[9656]) | (layer0_outputs[6267]));
    assign outputs[161] = ~((layer0_outputs[3978]) | (layer0_outputs[10005]));
    assign outputs[162] = ~(layer0_outputs[5912]);
    assign outputs[163] = (layer0_outputs[9851]) | (layer0_outputs[1593]);
    assign outputs[164] = (layer0_outputs[410]) & ~(layer0_outputs[1853]);
    assign outputs[165] = ~(layer0_outputs[3690]);
    assign outputs[166] = ~((layer0_outputs[3642]) ^ (layer0_outputs[334]));
    assign outputs[167] = layer0_outputs[9341];
    assign outputs[168] = ~(layer0_outputs[9223]);
    assign outputs[169] = (layer0_outputs[1640]) ^ (layer0_outputs[1625]);
    assign outputs[170] = (layer0_outputs[8525]) & ~(layer0_outputs[2851]);
    assign outputs[171] = ~((layer0_outputs[596]) | (layer0_outputs[5130]));
    assign outputs[172] = layer0_outputs[8931];
    assign outputs[173] = ~(layer0_outputs[10121]);
    assign outputs[174] = ~(layer0_outputs[1134]);
    assign outputs[175] = layer0_outputs[358];
    assign outputs[176] = ~(layer0_outputs[8258]);
    assign outputs[177] = ~(layer0_outputs[29]);
    assign outputs[178] = layer0_outputs[4276];
    assign outputs[179] = layer0_outputs[5395];
    assign outputs[180] = ~((layer0_outputs[5616]) & (layer0_outputs[5636]));
    assign outputs[181] = layer0_outputs[6849];
    assign outputs[182] = ~(layer0_outputs[2063]);
    assign outputs[183] = ~(layer0_outputs[8147]);
    assign outputs[184] = ~(layer0_outputs[7590]);
    assign outputs[185] = layer0_outputs[2950];
    assign outputs[186] = (layer0_outputs[6179]) | (layer0_outputs[7703]);
    assign outputs[187] = layer0_outputs[624];
    assign outputs[188] = layer0_outputs[3546];
    assign outputs[189] = (layer0_outputs[3293]) & ~(layer0_outputs[8541]);
    assign outputs[190] = (layer0_outputs[2965]) & ~(layer0_outputs[7568]);
    assign outputs[191] = ~(layer0_outputs[3814]);
    assign outputs[192] = layer0_outputs[6820];
    assign outputs[193] = ~(layer0_outputs[8162]);
    assign outputs[194] = ~(layer0_outputs[8329]);
    assign outputs[195] = (layer0_outputs[8448]) & (layer0_outputs[1594]);
    assign outputs[196] = (layer0_outputs[5884]) ^ (layer0_outputs[1384]);
    assign outputs[197] = ~((layer0_outputs[4443]) ^ (layer0_outputs[5102]));
    assign outputs[198] = ~(layer0_outputs[3044]);
    assign outputs[199] = ~(layer0_outputs[2898]);
    assign outputs[200] = ~(layer0_outputs[4147]);
    assign outputs[201] = ~(layer0_outputs[3122]);
    assign outputs[202] = ~((layer0_outputs[336]) ^ (layer0_outputs[6472]));
    assign outputs[203] = layer0_outputs[8833];
    assign outputs[204] = ~(layer0_outputs[3791]);
    assign outputs[205] = ~((layer0_outputs[7163]) & (layer0_outputs[6768]));
    assign outputs[206] = (layer0_outputs[1464]) ^ (layer0_outputs[2378]);
    assign outputs[207] = layer0_outputs[6290];
    assign outputs[208] = layer0_outputs[4568];
    assign outputs[209] = ~(layer0_outputs[9328]);
    assign outputs[210] = (layer0_outputs[3440]) & (layer0_outputs[47]);
    assign outputs[211] = layer0_outputs[3453];
    assign outputs[212] = layer0_outputs[9638];
    assign outputs[213] = layer0_outputs[2121];
    assign outputs[214] = ~(layer0_outputs[2978]);
    assign outputs[215] = ~((layer0_outputs[1045]) & (layer0_outputs[5743]));
    assign outputs[216] = ~((layer0_outputs[3284]) ^ (layer0_outputs[134]));
    assign outputs[217] = ~(layer0_outputs[6217]);
    assign outputs[218] = ~(layer0_outputs[8060]) | (layer0_outputs[6522]);
    assign outputs[219] = (layer0_outputs[5878]) & ~(layer0_outputs[4963]);
    assign outputs[220] = layer0_outputs[9589];
    assign outputs[221] = (layer0_outputs[3739]) ^ (layer0_outputs[2590]);
    assign outputs[222] = layer0_outputs[6706];
    assign outputs[223] = (layer0_outputs[3761]) ^ (layer0_outputs[9110]);
    assign outputs[224] = ~((layer0_outputs[4659]) ^ (layer0_outputs[6536]));
    assign outputs[225] = ~((layer0_outputs[2694]) | (layer0_outputs[6409]));
    assign outputs[226] = ~(layer0_outputs[6834]);
    assign outputs[227] = layer0_outputs[2267];
    assign outputs[228] = ~(layer0_outputs[3805]);
    assign outputs[229] = ~(layer0_outputs[4885]) | (layer0_outputs[2613]);
    assign outputs[230] = layer0_outputs[4764];
    assign outputs[231] = (layer0_outputs[5621]) & ~(layer0_outputs[791]);
    assign outputs[232] = (layer0_outputs[7828]) ^ (layer0_outputs[9217]);
    assign outputs[233] = ~((layer0_outputs[6237]) ^ (layer0_outputs[5876]));
    assign outputs[234] = (layer0_outputs[4480]) & ~(layer0_outputs[1613]);
    assign outputs[235] = ~((layer0_outputs[5653]) & (layer0_outputs[2709]));
    assign outputs[236] = ~(layer0_outputs[2155]);
    assign outputs[237] = ~((layer0_outputs[4738]) ^ (layer0_outputs[1670]));
    assign outputs[238] = layer0_outputs[4799];
    assign outputs[239] = (layer0_outputs[5254]) & ~(layer0_outputs[6443]);
    assign outputs[240] = ~((layer0_outputs[9172]) ^ (layer0_outputs[5151]));
    assign outputs[241] = ~(layer0_outputs[5932]);
    assign outputs[242] = (layer0_outputs[7514]) & (layer0_outputs[3998]);
    assign outputs[243] = ~(layer0_outputs[7739]);
    assign outputs[244] = (layer0_outputs[3684]) ^ (layer0_outputs[6117]);
    assign outputs[245] = layer0_outputs[1363];
    assign outputs[246] = ~(layer0_outputs[10168]);
    assign outputs[247] = ~(layer0_outputs[2258]);
    assign outputs[248] = (layer0_outputs[7844]) & ~(layer0_outputs[4709]);
    assign outputs[249] = layer0_outputs[3028];
    assign outputs[250] = (layer0_outputs[10146]) ^ (layer0_outputs[6614]);
    assign outputs[251] = layer0_outputs[6261];
    assign outputs[252] = ~((layer0_outputs[10094]) ^ (layer0_outputs[2563]));
    assign outputs[253] = (layer0_outputs[392]) & ~(layer0_outputs[2382]);
    assign outputs[254] = (layer0_outputs[7223]) & ~(layer0_outputs[8628]);
    assign outputs[255] = (layer0_outputs[9246]) & (layer0_outputs[6086]);
    assign outputs[256] = layer0_outputs[5336];
    assign outputs[257] = ~(layer0_outputs[9325]) | (layer0_outputs[5410]);
    assign outputs[258] = layer0_outputs[3806];
    assign outputs[259] = (layer0_outputs[3955]) | (layer0_outputs[1683]);
    assign outputs[260] = ~(layer0_outputs[9244]) | (layer0_outputs[665]);
    assign outputs[261] = ~(layer0_outputs[3550]);
    assign outputs[262] = layer0_outputs[804];
    assign outputs[263] = ~(layer0_outputs[8061]);
    assign outputs[264] = ~(layer0_outputs[694]);
    assign outputs[265] = ~((layer0_outputs[6021]) & (layer0_outputs[9270]));
    assign outputs[266] = ~(layer0_outputs[5199]) | (layer0_outputs[2761]);
    assign outputs[267] = (layer0_outputs[7758]) & ~(layer0_outputs[3319]);
    assign outputs[268] = ~(layer0_outputs[8468]);
    assign outputs[269] = ~((layer0_outputs[9174]) | (layer0_outputs[1895]));
    assign outputs[270] = ~(layer0_outputs[5182]);
    assign outputs[271] = layer0_outputs[2459];
    assign outputs[272] = (layer0_outputs[8799]) ^ (layer0_outputs[3751]);
    assign outputs[273] = ~(layer0_outputs[10124]) | (layer0_outputs[7269]);
    assign outputs[274] = ~(layer0_outputs[519]);
    assign outputs[275] = (layer0_outputs[6464]) ^ (layer0_outputs[5209]);
    assign outputs[276] = layer0_outputs[6047];
    assign outputs[277] = ~((layer0_outputs[9410]) | (layer0_outputs[4427]));
    assign outputs[278] = ~(layer0_outputs[9428]);
    assign outputs[279] = ~((layer0_outputs[7225]) & (layer0_outputs[7423]));
    assign outputs[280] = ~(layer0_outputs[5199]);
    assign outputs[281] = ~(layer0_outputs[6602]);
    assign outputs[282] = layer0_outputs[10167];
    assign outputs[283] = ~((layer0_outputs[770]) | (layer0_outputs[4414]));
    assign outputs[284] = ~(layer0_outputs[5605]);
    assign outputs[285] = (layer0_outputs[3542]) & ~(layer0_outputs[113]);
    assign outputs[286] = (layer0_outputs[7364]) ^ (layer0_outputs[4438]);
    assign outputs[287] = (layer0_outputs[77]) | (layer0_outputs[3685]);
    assign outputs[288] = ~(layer0_outputs[6687]);
    assign outputs[289] = (layer0_outputs[7350]) & ~(layer0_outputs[4164]);
    assign outputs[290] = ~(layer0_outputs[8801]);
    assign outputs[291] = layer0_outputs[4608];
    assign outputs[292] = ~(layer0_outputs[9523]) | (layer0_outputs[3806]);
    assign outputs[293] = (layer0_outputs[3798]) & ~(layer0_outputs[3970]);
    assign outputs[294] = layer0_outputs[624];
    assign outputs[295] = layer0_outputs[7291];
    assign outputs[296] = layer0_outputs[5389];
    assign outputs[297] = ~(layer0_outputs[8876]);
    assign outputs[298] = ~(layer0_outputs[4711]);
    assign outputs[299] = layer0_outputs[517];
    assign outputs[300] = ~(layer0_outputs[8430]);
    assign outputs[301] = ~(layer0_outputs[6503]);
    assign outputs[302] = ~(layer0_outputs[9363]);
    assign outputs[303] = ~(layer0_outputs[2524]);
    assign outputs[304] = ~(layer0_outputs[3456]);
    assign outputs[305] = layer0_outputs[8355];
    assign outputs[306] = (layer0_outputs[370]) ^ (layer0_outputs[7302]);
    assign outputs[307] = ~((layer0_outputs[9468]) & (layer0_outputs[2953]));
    assign outputs[308] = ~(layer0_outputs[8132]);
    assign outputs[309] = layer0_outputs[9907];
    assign outputs[310] = layer0_outputs[438];
    assign outputs[311] = layer0_outputs[5728];
    assign outputs[312] = ~(layer0_outputs[8900]);
    assign outputs[313] = ~((layer0_outputs[3862]) ^ (layer0_outputs[10236]));
    assign outputs[314] = (layer0_outputs[3338]) & (layer0_outputs[6860]);
    assign outputs[315] = ~(layer0_outputs[3506]);
    assign outputs[316] = layer0_outputs[5433];
    assign outputs[317] = ~(layer0_outputs[531]) | (layer0_outputs[8154]);
    assign outputs[318] = layer0_outputs[9619];
    assign outputs[319] = ~(layer0_outputs[337]) | (layer0_outputs[2686]);
    assign outputs[320] = (layer0_outputs[6296]) ^ (layer0_outputs[4921]);
    assign outputs[321] = (layer0_outputs[3085]) | (layer0_outputs[7166]);
    assign outputs[322] = ~(layer0_outputs[4678]);
    assign outputs[323] = (layer0_outputs[2680]) & (layer0_outputs[3345]);
    assign outputs[324] = layer0_outputs[8308];
    assign outputs[325] = ~((layer0_outputs[1732]) & (layer0_outputs[9208]));
    assign outputs[326] = ~(layer0_outputs[9401]);
    assign outputs[327] = (layer0_outputs[3435]) & ~(layer0_outputs[4945]);
    assign outputs[328] = ~((layer0_outputs[8436]) ^ (layer0_outputs[6627]));
    assign outputs[329] = ~((layer0_outputs[498]) | (layer0_outputs[4892]));
    assign outputs[330] = layer0_outputs[1366];
    assign outputs[331] = ~((layer0_outputs[4914]) & (layer0_outputs[3374]));
    assign outputs[332] = (layer0_outputs[2084]) & ~(layer0_outputs[9839]);
    assign outputs[333] = (layer0_outputs[837]) | (layer0_outputs[8511]);
    assign outputs[334] = ~(layer0_outputs[5664]) | (layer0_outputs[9795]);
    assign outputs[335] = ~((layer0_outputs[4652]) & (layer0_outputs[3123]));
    assign outputs[336] = (layer0_outputs[7302]) | (layer0_outputs[467]);
    assign outputs[337] = ~(layer0_outputs[2620]);
    assign outputs[338] = ~(layer0_outputs[4631]) | (layer0_outputs[6494]);
    assign outputs[339] = ~(layer0_outputs[5196]);
    assign outputs[340] = ~((layer0_outputs[1895]) & (layer0_outputs[4382]));
    assign outputs[341] = ~(layer0_outputs[1502]) | (layer0_outputs[2847]);
    assign outputs[342] = ~(layer0_outputs[6883]);
    assign outputs[343] = ~((layer0_outputs[9187]) & (layer0_outputs[9438]));
    assign outputs[344] = ~(layer0_outputs[58]);
    assign outputs[345] = layer0_outputs[7588];
    assign outputs[346] = layer0_outputs[639];
    assign outputs[347] = layer0_outputs[7441];
    assign outputs[348] = ~((layer0_outputs[3414]) & (layer0_outputs[4970]));
    assign outputs[349] = ~((layer0_outputs[2783]) & (layer0_outputs[8885]));
    assign outputs[350] = (layer0_outputs[8940]) & ~(layer0_outputs[2058]);
    assign outputs[351] = ~((layer0_outputs[1641]) ^ (layer0_outputs[7114]));
    assign outputs[352] = ~(layer0_outputs[177]);
    assign outputs[353] = (layer0_outputs[3459]) & ~(layer0_outputs[7767]);
    assign outputs[354] = ~(layer0_outputs[2100]);
    assign outputs[355] = ~((layer0_outputs[2451]) ^ (layer0_outputs[1351]));
    assign outputs[356] = ~(layer0_outputs[3473]);
    assign outputs[357] = (layer0_outputs[8443]) & ~(layer0_outputs[6821]);
    assign outputs[358] = layer0_outputs[3904];
    assign outputs[359] = ~(layer0_outputs[4972]);
    assign outputs[360] = ~(layer0_outputs[6032]);
    assign outputs[361] = (layer0_outputs[409]) ^ (layer0_outputs[1151]);
    assign outputs[362] = layer0_outputs[8626];
    assign outputs[363] = (layer0_outputs[3357]) ^ (layer0_outputs[9311]);
    assign outputs[364] = layer0_outputs[8907];
    assign outputs[365] = ~((layer0_outputs[2495]) ^ (layer0_outputs[8688]));
    assign outputs[366] = layer0_outputs[9248];
    assign outputs[367] = layer0_outputs[606];
    assign outputs[368] = ~(layer0_outputs[8326]);
    assign outputs[369] = layer0_outputs[5942];
    assign outputs[370] = layer0_outputs[7857];
    assign outputs[371] = ~((layer0_outputs[10170]) | (layer0_outputs[3789]));
    assign outputs[372] = ~((layer0_outputs[7397]) | (layer0_outputs[1696]));
    assign outputs[373] = layer0_outputs[3094];
    assign outputs[374] = ~(layer0_outputs[8086]);
    assign outputs[375] = (layer0_outputs[6215]) & (layer0_outputs[1466]);
    assign outputs[376] = (layer0_outputs[1312]) & (layer0_outputs[627]);
    assign outputs[377] = ~((layer0_outputs[6206]) | (layer0_outputs[4972]));
    assign outputs[378] = ~(layer0_outputs[4949]);
    assign outputs[379] = ~(layer0_outputs[5530]) | (layer0_outputs[1876]);
    assign outputs[380] = layer0_outputs[2567];
    assign outputs[381] = ~((layer0_outputs[3991]) ^ (layer0_outputs[7012]));
    assign outputs[382] = ~((layer0_outputs[1476]) & (layer0_outputs[9307]));
    assign outputs[383] = ~((layer0_outputs[5671]) & (layer0_outputs[3019]));
    assign outputs[384] = layer0_outputs[7918];
    assign outputs[385] = layer0_outputs[4955];
    assign outputs[386] = (layer0_outputs[8671]) & ~(layer0_outputs[3570]);
    assign outputs[387] = layer0_outputs[6955];
    assign outputs[388] = layer0_outputs[3904];
    assign outputs[389] = ~(layer0_outputs[9309]) | (layer0_outputs[7736]);
    assign outputs[390] = ~(layer0_outputs[5790]);
    assign outputs[391] = ~((layer0_outputs[169]) ^ (layer0_outputs[3546]));
    assign outputs[392] = (layer0_outputs[385]) ^ (layer0_outputs[8878]);
    assign outputs[393] = (layer0_outputs[8786]) ^ (layer0_outputs[8821]);
    assign outputs[394] = ~(layer0_outputs[6838]);
    assign outputs[395] = (layer0_outputs[8851]) ^ (layer0_outputs[8197]);
    assign outputs[396] = layer0_outputs[6702];
    assign outputs[397] = layer0_outputs[296];
    assign outputs[398] = layer0_outputs[9603];
    assign outputs[399] = ~(layer0_outputs[6620]) | (layer0_outputs[3698]);
    assign outputs[400] = (layer0_outputs[7696]) | (layer0_outputs[2460]);
    assign outputs[401] = ~(layer0_outputs[580]);
    assign outputs[402] = ~(layer0_outputs[9808]) | (layer0_outputs[643]);
    assign outputs[403] = ~((layer0_outputs[6079]) | (layer0_outputs[7249]));
    assign outputs[404] = ~((layer0_outputs[3513]) | (layer0_outputs[999]));
    assign outputs[405] = (layer0_outputs[6655]) ^ (layer0_outputs[1175]);
    assign outputs[406] = layer0_outputs[10000];
    assign outputs[407] = layer0_outputs[3496];
    assign outputs[408] = layer0_outputs[8947];
    assign outputs[409] = ~(layer0_outputs[1143]);
    assign outputs[410] = (layer0_outputs[3850]) ^ (layer0_outputs[2560]);
    assign outputs[411] = ~(layer0_outputs[5550]);
    assign outputs[412] = (layer0_outputs[6836]) ^ (layer0_outputs[4229]);
    assign outputs[413] = ~(layer0_outputs[7029]);
    assign outputs[414] = ~(layer0_outputs[6228]);
    assign outputs[415] = layer0_outputs[3679];
    assign outputs[416] = ~(layer0_outputs[5431]);
    assign outputs[417] = (layer0_outputs[8745]) & ~(layer0_outputs[2603]);
    assign outputs[418] = ~(layer0_outputs[7561]);
    assign outputs[419] = (layer0_outputs[1362]) & (layer0_outputs[7468]);
    assign outputs[420] = layer0_outputs[5807];
    assign outputs[421] = ~(layer0_outputs[2000]);
    assign outputs[422] = layer0_outputs[6557];
    assign outputs[423] = layer0_outputs[4735];
    assign outputs[424] = (layer0_outputs[628]) ^ (layer0_outputs[3925]);
    assign outputs[425] = layer0_outputs[845];
    assign outputs[426] = ~(layer0_outputs[9579]);
    assign outputs[427] = ~(layer0_outputs[8033]) | (layer0_outputs[9874]);
    assign outputs[428] = layer0_outputs[5746];
    assign outputs[429] = layer0_outputs[6938];
    assign outputs[430] = ~((layer0_outputs[475]) & (layer0_outputs[3567]));
    assign outputs[431] = ~(layer0_outputs[4357]);
    assign outputs[432] = ~(layer0_outputs[9406]);
    assign outputs[433] = ~((layer0_outputs[8641]) ^ (layer0_outputs[8661]));
    assign outputs[434] = ~((layer0_outputs[2643]) & (layer0_outputs[9422]));
    assign outputs[435] = ~((layer0_outputs[2815]) & (layer0_outputs[6364]));
    assign outputs[436] = (layer0_outputs[967]) ^ (layer0_outputs[10202]);
    assign outputs[437] = layer0_outputs[6465];
    assign outputs[438] = ~((layer0_outputs[4533]) ^ (layer0_outputs[4327]));
    assign outputs[439] = ~((layer0_outputs[3842]) & (layer0_outputs[2364]));
    assign outputs[440] = layer0_outputs[61];
    assign outputs[441] = ~(layer0_outputs[1795]) | (layer0_outputs[6889]);
    assign outputs[442] = layer0_outputs[3882];
    assign outputs[443] = layer0_outputs[9555];
    assign outputs[444] = (layer0_outputs[6975]) ^ (layer0_outputs[6350]);
    assign outputs[445] = (layer0_outputs[4492]) & ~(layer0_outputs[8846]);
    assign outputs[446] = ~(layer0_outputs[5130]);
    assign outputs[447] = ~(layer0_outputs[6264]);
    assign outputs[448] = (layer0_outputs[4474]) & ~(layer0_outputs[7254]);
    assign outputs[449] = ~(layer0_outputs[9318]) | (layer0_outputs[4003]);
    assign outputs[450] = layer0_outputs[1322];
    assign outputs[451] = ~(layer0_outputs[357]);
    assign outputs[452] = layer0_outputs[2958];
    assign outputs[453] = (layer0_outputs[6613]) & (layer0_outputs[8713]);
    assign outputs[454] = ~(layer0_outputs[2317]);
    assign outputs[455] = (layer0_outputs[3318]) & ~(layer0_outputs[8625]);
    assign outputs[456] = ~((layer0_outputs[9094]) ^ (layer0_outputs[6682]));
    assign outputs[457] = (layer0_outputs[1907]) & ~(layer0_outputs[3921]);
    assign outputs[458] = ~((layer0_outputs[1391]) ^ (layer0_outputs[4051]));
    assign outputs[459] = ~(layer0_outputs[8793]);
    assign outputs[460] = layer0_outputs[2210];
    assign outputs[461] = layer0_outputs[344];
    assign outputs[462] = ~(layer0_outputs[7824]) | (layer0_outputs[3892]);
    assign outputs[463] = layer0_outputs[266];
    assign outputs[464] = ~(layer0_outputs[9531]) | (layer0_outputs[688]);
    assign outputs[465] = layer0_outputs[2157];
    assign outputs[466] = ~(layer0_outputs[5783]);
    assign outputs[467] = layer0_outputs[6533];
    assign outputs[468] = ~((layer0_outputs[877]) & (layer0_outputs[121]));
    assign outputs[469] = layer0_outputs[2062];
    assign outputs[470] = (layer0_outputs[5681]) ^ (layer0_outputs[9596]);
    assign outputs[471] = ~((layer0_outputs[6328]) ^ (layer0_outputs[6102]));
    assign outputs[472] = ~(layer0_outputs[5561]);
    assign outputs[473] = layer0_outputs[4509];
    assign outputs[474] = (layer0_outputs[5587]) | (layer0_outputs[2631]);
    assign outputs[475] = (layer0_outputs[3178]) ^ (layer0_outputs[1928]);
    assign outputs[476] = (layer0_outputs[8456]) & ~(layer0_outputs[3404]);
    assign outputs[477] = ~(layer0_outputs[2808]) | (layer0_outputs[1488]);
    assign outputs[478] = layer0_outputs[1163];
    assign outputs[479] = (layer0_outputs[2297]) ^ (layer0_outputs[8951]);
    assign outputs[480] = ~((layer0_outputs[2376]) ^ (layer0_outputs[1004]));
    assign outputs[481] = ~(layer0_outputs[3730]);
    assign outputs[482] = ~(layer0_outputs[1176]) | (layer0_outputs[6177]);
    assign outputs[483] = ~(layer0_outputs[593]);
    assign outputs[484] = ~((layer0_outputs[2994]) ^ (layer0_outputs[7571]));
    assign outputs[485] = (layer0_outputs[10013]) & (layer0_outputs[2904]);
    assign outputs[486] = ~(layer0_outputs[6399]);
    assign outputs[487] = ~(layer0_outputs[2595]) | (layer0_outputs[8732]);
    assign outputs[488] = ~(layer0_outputs[6228]);
    assign outputs[489] = ~(layer0_outputs[9916]);
    assign outputs[490] = (layer0_outputs[3382]) & ~(layer0_outputs[2734]);
    assign outputs[491] = ~(layer0_outputs[8550]);
    assign outputs[492] = ~(layer0_outputs[3232]);
    assign outputs[493] = (layer0_outputs[3913]) ^ (layer0_outputs[9288]);
    assign outputs[494] = layer0_outputs[7721];
    assign outputs[495] = ~(layer0_outputs[7660]) | (layer0_outputs[7506]);
    assign outputs[496] = ~(layer0_outputs[7584]);
    assign outputs[497] = layer0_outputs[10103];
    assign outputs[498] = ~((layer0_outputs[6320]) ^ (layer0_outputs[7430]));
    assign outputs[499] = ~((layer0_outputs[6400]) & (layer0_outputs[9896]));
    assign outputs[500] = ~((layer0_outputs[6192]) ^ (layer0_outputs[2503]));
    assign outputs[501] = layer0_outputs[8714];
    assign outputs[502] = (layer0_outputs[4506]) & ~(layer0_outputs[37]);
    assign outputs[503] = ~(layer0_outputs[387]);
    assign outputs[504] = ~((layer0_outputs[9640]) | (layer0_outputs[7777]));
    assign outputs[505] = (layer0_outputs[4517]) ^ (layer0_outputs[5562]);
    assign outputs[506] = layer0_outputs[5066];
    assign outputs[507] = (layer0_outputs[438]) & (layer0_outputs[7026]);
    assign outputs[508] = (layer0_outputs[6926]) & ~(layer0_outputs[1436]);
    assign outputs[509] = layer0_outputs[977];
    assign outputs[510] = ~(layer0_outputs[2369]) | (layer0_outputs[974]);
    assign outputs[511] = ~(layer0_outputs[3471]) | (layer0_outputs[5784]);
    assign outputs[512] = layer0_outputs[1053];
    assign outputs[513] = ~(layer0_outputs[9096]);
    assign outputs[514] = (layer0_outputs[1448]) & ~(layer0_outputs[1067]);
    assign outputs[515] = layer0_outputs[10145];
    assign outputs[516] = layer0_outputs[8218];
    assign outputs[517] = layer0_outputs[7672];
    assign outputs[518] = (layer0_outputs[2527]) & ~(layer0_outputs[2034]);
    assign outputs[519] = ~((layer0_outputs[1544]) ^ (layer0_outputs[6164]));
    assign outputs[520] = layer0_outputs[9285];
    assign outputs[521] = ~((layer0_outputs[3030]) ^ (layer0_outputs[705]));
    assign outputs[522] = ~((layer0_outputs[3184]) | (layer0_outputs[2502]));
    assign outputs[523] = layer0_outputs[3634];
    assign outputs[524] = ~(layer0_outputs[418]) | (layer0_outputs[4790]);
    assign outputs[525] = ~((layer0_outputs[619]) & (layer0_outputs[7826]));
    assign outputs[526] = (layer0_outputs[1046]) & ~(layer0_outputs[5862]);
    assign outputs[527] = ~(layer0_outputs[4059]) | (layer0_outputs[4683]);
    assign outputs[528] = layer0_outputs[9473];
    assign outputs[529] = layer0_outputs[1146];
    assign outputs[530] = (layer0_outputs[6410]) & (layer0_outputs[1288]);
    assign outputs[531] = layer0_outputs[5809];
    assign outputs[532] = ~(layer0_outputs[9245]) | (layer0_outputs[9633]);
    assign outputs[533] = ~(layer0_outputs[2579]);
    assign outputs[534] = ~(layer0_outputs[5541]);
    assign outputs[535] = (layer0_outputs[3903]) ^ (layer0_outputs[4763]);
    assign outputs[536] = layer0_outputs[960];
    assign outputs[537] = layer0_outputs[4321];
    assign outputs[538] = ~(layer0_outputs[9368]);
    assign outputs[539] = layer0_outputs[796];
    assign outputs[540] = (layer0_outputs[7011]) ^ (layer0_outputs[6750]);
    assign outputs[541] = layer0_outputs[8293];
    assign outputs[542] = ~(layer0_outputs[1767]);
    assign outputs[543] = ~(layer0_outputs[9893]) | (layer0_outputs[2419]);
    assign outputs[544] = (layer0_outputs[3945]) | (layer0_outputs[219]);
    assign outputs[545] = ~(layer0_outputs[579]);
    assign outputs[546] = layer0_outputs[5044];
    assign outputs[547] = ~(layer0_outputs[1655]);
    assign outputs[548] = ~((layer0_outputs[1864]) | (layer0_outputs[9068]));
    assign outputs[549] = ~((layer0_outputs[10219]) ^ (layer0_outputs[2486]));
    assign outputs[550] = layer0_outputs[182];
    assign outputs[551] = ~(layer0_outputs[8746]);
    assign outputs[552] = (layer0_outputs[9408]) & ~(layer0_outputs[205]);
    assign outputs[553] = ~(layer0_outputs[8733]);
    assign outputs[554] = (layer0_outputs[3384]) ^ (layer0_outputs[47]);
    assign outputs[555] = (layer0_outputs[9776]) & ~(layer0_outputs[1820]);
    assign outputs[556] = layer0_outputs[3320];
    assign outputs[557] = layer0_outputs[481];
    assign outputs[558] = layer0_outputs[7327];
    assign outputs[559] = 1'b1;
    assign outputs[560] = layer0_outputs[1772];
    assign outputs[561] = ~(layer0_outputs[9484]) | (layer0_outputs[8865]);
    assign outputs[562] = (layer0_outputs[5985]) & (layer0_outputs[5039]);
    assign outputs[563] = (layer0_outputs[10030]) | (layer0_outputs[2543]);
    assign outputs[564] = ~(layer0_outputs[6512]);
    assign outputs[565] = layer0_outputs[7141];
    assign outputs[566] = ~(layer0_outputs[4804]);
    assign outputs[567] = layer0_outputs[4285];
    assign outputs[568] = ~(layer0_outputs[3934]);
    assign outputs[569] = ~(layer0_outputs[3537]);
    assign outputs[570] = ~((layer0_outputs[7580]) ^ (layer0_outputs[9169]));
    assign outputs[571] = ~(layer0_outputs[8521]);
    assign outputs[572] = (layer0_outputs[3086]) ^ (layer0_outputs[7211]);
    assign outputs[573] = (layer0_outputs[7712]) & (layer0_outputs[7605]);
    assign outputs[574] = ~(layer0_outputs[3360]);
    assign outputs[575] = (layer0_outputs[5068]) | (layer0_outputs[1727]);
    assign outputs[576] = layer0_outputs[4320];
    assign outputs[577] = ~((layer0_outputs[5385]) | (layer0_outputs[203]));
    assign outputs[578] = ~(layer0_outputs[9131]) | (layer0_outputs[1738]);
    assign outputs[579] = layer0_outputs[9627];
    assign outputs[580] = ~(layer0_outputs[6776]);
    assign outputs[581] = ~(layer0_outputs[7733]);
    assign outputs[582] = layer0_outputs[1106];
    assign outputs[583] = ~(layer0_outputs[2439]) | (layer0_outputs[4867]);
    assign outputs[584] = ~(layer0_outputs[8722]) | (layer0_outputs[263]);
    assign outputs[585] = ~(layer0_outputs[1425]);
    assign outputs[586] = (layer0_outputs[5313]) & ~(layer0_outputs[6919]);
    assign outputs[587] = layer0_outputs[2300];
    assign outputs[588] = ~((layer0_outputs[318]) ^ (layer0_outputs[9405]));
    assign outputs[589] = ~(layer0_outputs[4026]);
    assign outputs[590] = ~(layer0_outputs[96]);
    assign outputs[591] = (layer0_outputs[9785]) | (layer0_outputs[3372]);
    assign outputs[592] = (layer0_outputs[7705]) & (layer0_outputs[1658]);
    assign outputs[593] = ~(layer0_outputs[7664]);
    assign outputs[594] = (layer0_outputs[1595]) & ~(layer0_outputs[5718]);
    assign outputs[595] = ~((layer0_outputs[8007]) ^ (layer0_outputs[7325]));
    assign outputs[596] = (layer0_outputs[4205]) ^ (layer0_outputs[3705]);
    assign outputs[597] = layer0_outputs[6434];
    assign outputs[598] = layer0_outputs[7520];
    assign outputs[599] = layer0_outputs[143];
    assign outputs[600] = layer0_outputs[4683];
    assign outputs[601] = (layer0_outputs[1917]) ^ (layer0_outputs[7719]);
    assign outputs[602] = ~(layer0_outputs[8494]);
    assign outputs[603] = ~((layer0_outputs[4919]) ^ (layer0_outputs[10002]));
    assign outputs[604] = ~(layer0_outputs[8838]);
    assign outputs[605] = (layer0_outputs[5811]) ^ (layer0_outputs[5479]);
    assign outputs[606] = ~(layer0_outputs[7854]) | (layer0_outputs[1477]);
    assign outputs[607] = (layer0_outputs[10179]) ^ (layer0_outputs[9498]);
    assign outputs[608] = layer0_outputs[7083];
    assign outputs[609] = ~((layer0_outputs[1061]) ^ (layer0_outputs[3040]));
    assign outputs[610] = ~((layer0_outputs[4196]) & (layer0_outputs[5219]));
    assign outputs[611] = ~(layer0_outputs[1696]);
    assign outputs[612] = ~((layer0_outputs[7800]) ^ (layer0_outputs[2571]));
    assign outputs[613] = ~((layer0_outputs[1329]) ^ (layer0_outputs[6826]));
    assign outputs[614] = ~(layer0_outputs[2987]);
    assign outputs[615] = layer0_outputs[7334];
    assign outputs[616] = layer0_outputs[419];
    assign outputs[617] = layer0_outputs[8921];
    assign outputs[618] = ~(layer0_outputs[5734]);
    assign outputs[619] = ~((layer0_outputs[5840]) ^ (layer0_outputs[9035]));
    assign outputs[620] = (layer0_outputs[4820]) & ~(layer0_outputs[9501]);
    assign outputs[621] = (layer0_outputs[7483]) ^ (layer0_outputs[3508]);
    assign outputs[622] = layer0_outputs[5317];
    assign outputs[623] = ~(layer0_outputs[6398]) | (layer0_outputs[6165]);
    assign outputs[624] = (layer0_outputs[1857]) | (layer0_outputs[2402]);
    assign outputs[625] = (layer0_outputs[4065]) | (layer0_outputs[2510]);
    assign outputs[626] = ~(layer0_outputs[9037]);
    assign outputs[627] = ~(layer0_outputs[10076]);
    assign outputs[628] = ~(layer0_outputs[4580]);
    assign outputs[629] = layer0_outputs[4148];
    assign outputs[630] = ~(layer0_outputs[614]);
    assign outputs[631] = layer0_outputs[1353];
    assign outputs[632] = ~((layer0_outputs[9937]) ^ (layer0_outputs[8926]));
    assign outputs[633] = ~(layer0_outputs[7143]) | (layer0_outputs[6882]);
    assign outputs[634] = ~(layer0_outputs[1033]);
    assign outputs[635] = layer0_outputs[7016];
    assign outputs[636] = ~(layer0_outputs[1576]);
    assign outputs[637] = ~(layer0_outputs[881]);
    assign outputs[638] = ~(layer0_outputs[1190]);
    assign outputs[639] = ~(layer0_outputs[1392]);
    assign outputs[640] = ~((layer0_outputs[1631]) ^ (layer0_outputs[4436]));
    assign outputs[641] = layer0_outputs[9122];
    assign outputs[642] = ~(layer0_outputs[6310]);
    assign outputs[643] = layer0_outputs[4717];
    assign outputs[644] = layer0_outputs[2515];
    assign outputs[645] = ~(layer0_outputs[7704]) | (layer0_outputs[9852]);
    assign outputs[646] = layer0_outputs[3025];
    assign outputs[647] = ~((layer0_outputs[9493]) | (layer0_outputs[3808]));
    assign outputs[648] = ~((layer0_outputs[1352]) ^ (layer0_outputs[2042]));
    assign outputs[649] = layer0_outputs[6892];
    assign outputs[650] = (layer0_outputs[7236]) & ~(layer0_outputs[4117]);
    assign outputs[651] = layer0_outputs[781];
    assign outputs[652] = ~((layer0_outputs[1799]) & (layer0_outputs[9744]));
    assign outputs[653] = layer0_outputs[9700];
    assign outputs[654] = layer0_outputs[3238];
    assign outputs[655] = (layer0_outputs[5472]) ^ (layer0_outputs[2448]);
    assign outputs[656] = ~((layer0_outputs[7740]) | (layer0_outputs[6118]));
    assign outputs[657] = (layer0_outputs[1574]) ^ (layer0_outputs[7901]);
    assign outputs[658] = ~(layer0_outputs[4]);
    assign outputs[659] = layer0_outputs[6648];
    assign outputs[660] = ~(layer0_outputs[750]);
    assign outputs[661] = layer0_outputs[8787];
    assign outputs[662] = layer0_outputs[6486];
    assign outputs[663] = ~((layer0_outputs[4947]) ^ (layer0_outputs[7918]));
    assign outputs[664] = layer0_outputs[6125];
    assign outputs[665] = ~((layer0_outputs[5455]) ^ (layer0_outputs[8406]));
    assign outputs[666] = ~(layer0_outputs[4333]) | (layer0_outputs[6007]);
    assign outputs[667] = ~((layer0_outputs[7358]) | (layer0_outputs[6572]));
    assign outputs[668] = ~(layer0_outputs[6377]);
    assign outputs[669] = ~(layer0_outputs[4325]);
    assign outputs[670] = ~(layer0_outputs[8016]);
    assign outputs[671] = (layer0_outputs[3165]) & ~(layer0_outputs[6116]);
    assign outputs[672] = ~((layer0_outputs[7190]) ^ (layer0_outputs[7581]));
    assign outputs[673] = ~((layer0_outputs[8449]) | (layer0_outputs[348]));
    assign outputs[674] = layer0_outputs[3287];
    assign outputs[675] = ~((layer0_outputs[7400]) & (layer0_outputs[7048]));
    assign outputs[676] = ~(layer0_outputs[129]);
    assign outputs[677] = ~((layer0_outputs[2872]) | (layer0_outputs[8194]));
    assign outputs[678] = layer0_outputs[6480];
    assign outputs[679] = (layer0_outputs[6027]) & (layer0_outputs[4337]);
    assign outputs[680] = ~(layer0_outputs[9432]) | (layer0_outputs[9985]);
    assign outputs[681] = layer0_outputs[1206];
    assign outputs[682] = ~((layer0_outputs[3107]) ^ (layer0_outputs[213]));
    assign outputs[683] = ~((layer0_outputs[9691]) & (layer0_outputs[4713]));
    assign outputs[684] = ~(layer0_outputs[9836]);
    assign outputs[685] = ~(layer0_outputs[2834]);
    assign outputs[686] = ~((layer0_outputs[4164]) | (layer0_outputs[10225]));
    assign outputs[687] = (layer0_outputs[1384]) ^ (layer0_outputs[7388]);
    assign outputs[688] = ~(layer0_outputs[9451]);
    assign outputs[689] = (layer0_outputs[9544]) | (layer0_outputs[8031]);
    assign outputs[690] = (layer0_outputs[8387]) ^ (layer0_outputs[4687]);
    assign outputs[691] = layer0_outputs[5075];
    assign outputs[692] = (layer0_outputs[3104]) & ~(layer0_outputs[5308]);
    assign outputs[693] = (layer0_outputs[8575]) ^ (layer0_outputs[6066]);
    assign outputs[694] = ~((layer0_outputs[3505]) | (layer0_outputs[3366]));
    assign outputs[695] = (layer0_outputs[10117]) ^ (layer0_outputs[6165]);
    assign outputs[696] = ~(layer0_outputs[1884]);
    assign outputs[697] = ~((layer0_outputs[7744]) & (layer0_outputs[7421]));
    assign outputs[698] = layer0_outputs[403];
    assign outputs[699] = layer0_outputs[5554];
    assign outputs[700] = layer0_outputs[3779];
    assign outputs[701] = ~(layer0_outputs[7529]);
    assign outputs[702] = (layer0_outputs[3485]) ^ (layer0_outputs[846]);
    assign outputs[703] = ~(layer0_outputs[7836]) | (layer0_outputs[2959]);
    assign outputs[704] = ~((layer0_outputs[458]) ^ (layer0_outputs[1864]));
    assign outputs[705] = (layer0_outputs[9151]) ^ (layer0_outputs[1226]);
    assign outputs[706] = ~(layer0_outputs[9392]);
    assign outputs[707] = ~(layer0_outputs[7577]);
    assign outputs[708] = (layer0_outputs[2598]) | (layer0_outputs[3450]);
    assign outputs[709] = layer0_outputs[599];
    assign outputs[710] = ~(layer0_outputs[3207]);
    assign outputs[711] = layer0_outputs[1495];
    assign outputs[712] = ~((layer0_outputs[545]) ^ (layer0_outputs[2137]));
    assign outputs[713] = ~(layer0_outputs[9171]);
    assign outputs[714] = (layer0_outputs[3364]) ^ (layer0_outputs[1267]);
    assign outputs[715] = layer0_outputs[2415];
    assign outputs[716] = ~((layer0_outputs[2618]) ^ (layer0_outputs[3401]));
    assign outputs[717] = ~((layer0_outputs[6635]) ^ (layer0_outputs[1840]));
    assign outputs[718] = ~(layer0_outputs[4966]) | (layer0_outputs[1793]);
    assign outputs[719] = ~(layer0_outputs[6144]);
    assign outputs[720] = ~(layer0_outputs[3342]);
    assign outputs[721] = layer0_outputs[7802];
    assign outputs[722] = ~(layer0_outputs[5319]);
    assign outputs[723] = ~(layer0_outputs[7072]);
    assign outputs[724] = ~(layer0_outputs[8651]);
    assign outputs[725] = ~((layer0_outputs[9073]) ^ (layer0_outputs[8998]));
    assign outputs[726] = ~(layer0_outputs[2812]) | (layer0_outputs[4197]);
    assign outputs[727] = ~((layer0_outputs[8044]) ^ (layer0_outputs[3711]));
    assign outputs[728] = ~(layer0_outputs[9728]);
    assign outputs[729] = (layer0_outputs[9416]) ^ (layer0_outputs[1707]);
    assign outputs[730] = ~(layer0_outputs[4283]);
    assign outputs[731] = ~(layer0_outputs[5618]);
    assign outputs[732] = ~((layer0_outputs[1054]) | (layer0_outputs[473]));
    assign outputs[733] = ~(layer0_outputs[711]);
    assign outputs[734] = ~(layer0_outputs[7499]);
    assign outputs[735] = ~(layer0_outputs[5723]);
    assign outputs[736] = layer0_outputs[6107];
    assign outputs[737] = ~(layer0_outputs[82]);
    assign outputs[738] = ~(layer0_outputs[7456]);
    assign outputs[739] = layer0_outputs[3564];
    assign outputs[740] = ~(layer0_outputs[3660]);
    assign outputs[741] = layer0_outputs[1195];
    assign outputs[742] = ~((layer0_outputs[5794]) ^ (layer0_outputs[3824]));
    assign outputs[743] = layer0_outputs[8298];
    assign outputs[744] = ~(layer0_outputs[4391]);
    assign outputs[745] = ~(layer0_outputs[4444]);
    assign outputs[746] = layer0_outputs[484];
    assign outputs[747] = ~(layer0_outputs[3661]) | (layer0_outputs[7073]);
    assign outputs[748] = layer0_outputs[3143];
    assign outputs[749] = ~((layer0_outputs[840]) ^ (layer0_outputs[1471]));
    assign outputs[750] = ~(layer0_outputs[8373]) | (layer0_outputs[4022]);
    assign outputs[751] = layer0_outputs[7098];
    assign outputs[752] = layer0_outputs[2928];
    assign outputs[753] = ~(layer0_outputs[2036]);
    assign outputs[754] = (layer0_outputs[7119]) | (layer0_outputs[1150]);
    assign outputs[755] = ~(layer0_outputs[8396]);
    assign outputs[756] = ~(layer0_outputs[6212]);
    assign outputs[757] = layer0_outputs[4199];
    assign outputs[758] = ~(layer0_outputs[6669]) | (layer0_outputs[402]);
    assign outputs[759] = (layer0_outputs[7365]) & ~(layer0_outputs[7336]);
    assign outputs[760] = 1'b1;
    assign outputs[761] = ~((layer0_outputs[5654]) ^ (layer0_outputs[5001]));
    assign outputs[762] = ~(layer0_outputs[5653]);
    assign outputs[763] = layer0_outputs[9553];
    assign outputs[764] = ~((layer0_outputs[6420]) ^ (layer0_outputs[2911]));
    assign outputs[765] = ~(layer0_outputs[4162]);
    assign outputs[766] = ~(layer0_outputs[7999]);
    assign outputs[767] = (layer0_outputs[2713]) & ~(layer0_outputs[2060]);
    assign outputs[768] = ~(layer0_outputs[1217]) | (layer0_outputs[10064]);
    assign outputs[769] = layer0_outputs[120];
    assign outputs[770] = ~((layer0_outputs[9308]) ^ (layer0_outputs[7722]));
    assign outputs[771] = ~(layer0_outputs[7749]);
    assign outputs[772] = ~((layer0_outputs[3534]) ^ (layer0_outputs[6721]));
    assign outputs[773] = ~(layer0_outputs[9781]);
    assign outputs[774] = layer0_outputs[3397];
    assign outputs[775] = (layer0_outputs[2172]) & (layer0_outputs[5732]);
    assign outputs[776] = (layer0_outputs[10132]) & (layer0_outputs[2216]);
    assign outputs[777] = layer0_outputs[4036];
    assign outputs[778] = ~((layer0_outputs[4968]) ^ (layer0_outputs[1835]));
    assign outputs[779] = layer0_outputs[4226];
    assign outputs[780] = (layer0_outputs[6380]) ^ (layer0_outputs[9851]);
    assign outputs[781] = ~(layer0_outputs[6958]);
    assign outputs[782] = ~(layer0_outputs[3298]) | (layer0_outputs[5727]);
    assign outputs[783] = layer0_outputs[4712];
    assign outputs[784] = (layer0_outputs[6286]) & ~(layer0_outputs[5523]);
    assign outputs[785] = layer0_outputs[6589];
    assign outputs[786] = ~(layer0_outputs[7926]);
    assign outputs[787] = ~(layer0_outputs[3476]);
    assign outputs[788] = ~(layer0_outputs[5353]);
    assign outputs[789] = ~(layer0_outputs[1896]);
    assign outputs[790] = ~(layer0_outputs[9259]);
    assign outputs[791] = (layer0_outputs[726]) & ~(layer0_outputs[2338]);
    assign outputs[792] = ~((layer0_outputs[1688]) ^ (layer0_outputs[3749]));
    assign outputs[793] = (layer0_outputs[1738]) | (layer0_outputs[8882]);
    assign outputs[794] = ~((layer0_outputs[8032]) ^ (layer0_outputs[799]));
    assign outputs[795] = layer0_outputs[6164];
    assign outputs[796] = (layer0_outputs[3707]) & ~(layer0_outputs[9182]);
    assign outputs[797] = 1'b1;
    assign outputs[798] = (layer0_outputs[5842]) & ~(layer0_outputs[2592]);
    assign outputs[799] = ~(layer0_outputs[2381]);
    assign outputs[800] = ~(layer0_outputs[6242]);
    assign outputs[801] = layer0_outputs[2817];
    assign outputs[802] = (layer0_outputs[7814]) & ~(layer0_outputs[1828]);
    assign outputs[803] = ~((layer0_outputs[7859]) ^ (layer0_outputs[5001]));
    assign outputs[804] = ~(layer0_outputs[356]);
    assign outputs[805] = ~(layer0_outputs[6479]);
    assign outputs[806] = layer0_outputs[388];
    assign outputs[807] = layer0_outputs[2847];
    assign outputs[808] = ~((layer0_outputs[5315]) ^ (layer0_outputs[9355]));
    assign outputs[809] = ~(layer0_outputs[8812]);
    assign outputs[810] = ~((layer0_outputs[7490]) ^ (layer0_outputs[6543]));
    assign outputs[811] = (layer0_outputs[4465]) & ~(layer0_outputs[7484]);
    assign outputs[812] = layer0_outputs[5467];
    assign outputs[813] = (layer0_outputs[3899]) | (layer0_outputs[7220]);
    assign outputs[814] = ~(layer0_outputs[5899]);
    assign outputs[815] = layer0_outputs[4273];
    assign outputs[816] = (layer0_outputs[6197]) ^ (layer0_outputs[1121]);
    assign outputs[817] = ~(layer0_outputs[6435]);
    assign outputs[818] = layer0_outputs[1833];
    assign outputs[819] = ~(layer0_outputs[10201]);
    assign outputs[820] = ~((layer0_outputs[2992]) ^ (layer0_outputs[6480]));
    assign outputs[821] = ~(layer0_outputs[8466]);
    assign outputs[822] = ~(layer0_outputs[4627]) | (layer0_outputs[277]);
    assign outputs[823] = ~((layer0_outputs[1898]) & (layer0_outputs[4548]));
    assign outputs[824] = (layer0_outputs[5400]) & (layer0_outputs[4915]);
    assign outputs[825] = ~(layer0_outputs[3067]) | (layer0_outputs[5749]);
    assign outputs[826] = (layer0_outputs[2977]) | (layer0_outputs[3055]);
    assign outputs[827] = layer0_outputs[9894];
    assign outputs[828] = ~((layer0_outputs[5675]) & (layer0_outputs[4675]));
    assign outputs[829] = ~((layer0_outputs[910]) | (layer0_outputs[5346]));
    assign outputs[830] = (layer0_outputs[9420]) ^ (layer0_outputs[4981]);
    assign outputs[831] = layer0_outputs[3196];
    assign outputs[832] = ~(layer0_outputs[8634]) | (layer0_outputs[2146]);
    assign outputs[833] = ~((layer0_outputs[9228]) | (layer0_outputs[5118]));
    assign outputs[834] = layer0_outputs[5274];
    assign outputs[835] = (layer0_outputs[1357]) & ~(layer0_outputs[6078]);
    assign outputs[836] = ~(layer0_outputs[8857]);
    assign outputs[837] = ~((layer0_outputs[5488]) & (layer0_outputs[4007]));
    assign outputs[838] = ~(layer0_outputs[2122]);
    assign outputs[839] = ~(layer0_outputs[7741]);
    assign outputs[840] = ~(layer0_outputs[8723]);
    assign outputs[841] = ~(layer0_outputs[3255]) | (layer0_outputs[1816]);
    assign outputs[842] = layer0_outputs[2699];
    assign outputs[843] = ~((layer0_outputs[3358]) | (layer0_outputs[3353]));
    assign outputs[844] = ~(layer0_outputs[9413]);
    assign outputs[845] = (layer0_outputs[6119]) & ~(layer0_outputs[5604]);
    assign outputs[846] = ~(layer0_outputs[1154]) | (layer0_outputs[9389]);
    assign outputs[847] = ~(layer0_outputs[1650]);
    assign outputs[848] = layer0_outputs[7239];
    assign outputs[849] = (layer0_outputs[1266]) & (layer0_outputs[9052]);
    assign outputs[850] = layer0_outputs[3523];
    assign outputs[851] = layer0_outputs[359];
    assign outputs[852] = layer0_outputs[8774];
    assign outputs[853] = ~((layer0_outputs[699]) ^ (layer0_outputs[1196]));
    assign outputs[854] = ~(layer0_outputs[5047]);
    assign outputs[855] = ~(layer0_outputs[1997]);
    assign outputs[856] = ~(layer0_outputs[4392]);
    assign outputs[857] = ~((layer0_outputs[5406]) & (layer0_outputs[4612]));
    assign outputs[858] = ~(layer0_outputs[4406]);
    assign outputs[859] = ~(layer0_outputs[6916]);
    assign outputs[860] = ~((layer0_outputs[7397]) | (layer0_outputs[4154]));
    assign outputs[861] = layer0_outputs[5508];
    assign outputs[862] = ~(layer0_outputs[9648]);
    assign outputs[863] = ~(layer0_outputs[6804]);
    assign outputs[864] = layer0_outputs[6840];
    assign outputs[865] = ~((layer0_outputs[10071]) ^ (layer0_outputs[9445]));
    assign outputs[866] = layer0_outputs[9830];
    assign outputs[867] = layer0_outputs[4980];
    assign outputs[868] = layer0_outputs[259];
    assign outputs[869] = layer0_outputs[9575];
    assign outputs[870] = ~(layer0_outputs[4593]);
    assign outputs[871] = (layer0_outputs[4685]) & (layer0_outputs[5902]);
    assign outputs[872] = ~((layer0_outputs[1305]) | (layer0_outputs[6658]));
    assign outputs[873] = layer0_outputs[4556];
    assign outputs[874] = layer0_outputs[6528];
    assign outputs[875] = ~((layer0_outputs[622]) ^ (layer0_outputs[5089]));
    assign outputs[876] = (layer0_outputs[7576]) & ~(layer0_outputs[7544]);
    assign outputs[877] = ~((layer0_outputs[3586]) ^ (layer0_outputs[6643]));
    assign outputs[878] = (layer0_outputs[1688]) & ~(layer0_outputs[152]);
    assign outputs[879] = ~(layer0_outputs[1672]) | (layer0_outputs[616]);
    assign outputs[880] = (layer0_outputs[6932]) | (layer0_outputs[5631]);
    assign outputs[881] = ~(layer0_outputs[139]) | (layer0_outputs[6884]);
    assign outputs[882] = ~(layer0_outputs[1402]);
    assign outputs[883] = layer0_outputs[2908];
    assign outputs[884] = layer0_outputs[8728];
    assign outputs[885] = ~(layer0_outputs[5561]) | (layer0_outputs[6611]);
    assign outputs[886] = ~(layer0_outputs[160]);
    assign outputs[887] = layer0_outputs[3337];
    assign outputs[888] = ~(layer0_outputs[9383]);
    assign outputs[889] = (layer0_outputs[7242]) & (layer0_outputs[9389]);
    assign outputs[890] = ~(layer0_outputs[8887]);
    assign outputs[891] = ~(layer0_outputs[5381]);
    assign outputs[892] = ~((layer0_outputs[4364]) ^ (layer0_outputs[3799]));
    assign outputs[893] = layer0_outputs[4522];
    assign outputs[894] = layer0_outputs[155];
    assign outputs[895] = ~((layer0_outputs[3215]) & (layer0_outputs[1763]));
    assign outputs[896] = layer0_outputs[5882];
    assign outputs[897] = layer0_outputs[9569];
    assign outputs[898] = layer0_outputs[7178];
    assign outputs[899] = ~(layer0_outputs[2209]);
    assign outputs[900] = (layer0_outputs[3841]) ^ (layer0_outputs[340]);
    assign outputs[901] = ~((layer0_outputs[7897]) | (layer0_outputs[478]));
    assign outputs[902] = ~(layer0_outputs[6248]);
    assign outputs[903] = ~((layer0_outputs[10189]) ^ (layer0_outputs[180]));
    assign outputs[904] = (layer0_outputs[6744]) ^ (layer0_outputs[2368]);
    assign outputs[905] = (layer0_outputs[2857]) ^ (layer0_outputs[4000]);
    assign outputs[906] = ~((layer0_outputs[9712]) ^ (layer0_outputs[5389]));
    assign outputs[907] = layer0_outputs[4321];
    assign outputs[908] = (layer0_outputs[2222]) ^ (layer0_outputs[6387]);
    assign outputs[909] = ~((layer0_outputs[3073]) & (layer0_outputs[6470]));
    assign outputs[910] = layer0_outputs[9019];
    assign outputs[911] = ~(layer0_outputs[7410]);
    assign outputs[912] = (layer0_outputs[4636]) ^ (layer0_outputs[3583]);
    assign outputs[913] = ~(layer0_outputs[3825]) | (layer0_outputs[7006]);
    assign outputs[914] = layer0_outputs[8811];
    assign outputs[915] = (layer0_outputs[5078]) & ~(layer0_outputs[7862]);
    assign outputs[916] = (layer0_outputs[7275]) & (layer0_outputs[2693]);
    assign outputs[917] = layer0_outputs[4284];
    assign outputs[918] = ~(layer0_outputs[2420]) | (layer0_outputs[2457]);
    assign outputs[919] = (layer0_outputs[3572]) ^ (layer0_outputs[6506]);
    assign outputs[920] = layer0_outputs[1113];
    assign outputs[921] = ~(layer0_outputs[7225]);
    assign outputs[922] = layer0_outputs[331];
    assign outputs[923] = ~(layer0_outputs[4578]);
    assign outputs[924] = ~(layer0_outputs[7568]);
    assign outputs[925] = layer0_outputs[317];
    assign outputs[926] = (layer0_outputs[2870]) & ~(layer0_outputs[8114]);
    assign outputs[927] = 1'b1;
    assign outputs[928] = layer0_outputs[2017];
    assign outputs[929] = ~((layer0_outputs[6514]) & (layer0_outputs[1722]));
    assign outputs[930] = ~(layer0_outputs[8365]);
    assign outputs[931] = ~(layer0_outputs[3864]);
    assign outputs[932] = ~(layer0_outputs[8642]);
    assign outputs[933] = ~(layer0_outputs[3221]);
    assign outputs[934] = (layer0_outputs[3877]) ^ (layer0_outputs[6590]);
    assign outputs[935] = ~((layer0_outputs[5363]) & (layer0_outputs[941]));
    assign outputs[936] = ~((layer0_outputs[9301]) | (layer0_outputs[3958]));
    assign outputs[937] = ~(layer0_outputs[336]);
    assign outputs[938] = (layer0_outputs[4388]) & ~(layer0_outputs[1487]);
    assign outputs[939] = ~(layer0_outputs[3089]);
    assign outputs[940] = ~((layer0_outputs[7966]) | (layer0_outputs[6879]));
    assign outputs[941] = (layer0_outputs[7137]) | (layer0_outputs[9152]);
    assign outputs[942] = ~((layer0_outputs[4228]) | (layer0_outputs[1695]));
    assign outputs[943] = (layer0_outputs[2075]) ^ (layer0_outputs[5088]);
    assign outputs[944] = (layer0_outputs[1210]) ^ (layer0_outputs[6727]);
    assign outputs[945] = ~(layer0_outputs[2694]);
    assign outputs[946] = (layer0_outputs[8617]) & ~(layer0_outputs[3208]);
    assign outputs[947] = (layer0_outputs[9616]) & (layer0_outputs[6283]);
    assign outputs[948] = (layer0_outputs[3075]) ^ (layer0_outputs[1664]);
    assign outputs[949] = layer0_outputs[6562];
    assign outputs[950] = ~(layer0_outputs[2531]) | (layer0_outputs[721]);
    assign outputs[951] = ~(layer0_outputs[6935]) | (layer0_outputs[140]);
    assign outputs[952] = (layer0_outputs[604]) ^ (layer0_outputs[9361]);
    assign outputs[953] = layer0_outputs[1434];
    assign outputs[954] = layer0_outputs[3243];
    assign outputs[955] = ~(layer0_outputs[395]);
    assign outputs[956] = layer0_outputs[3320];
    assign outputs[957] = ~((layer0_outputs[3322]) ^ (layer0_outputs[3035]));
    assign outputs[958] = ~(layer0_outputs[6057]);
    assign outputs[959] = (layer0_outputs[806]) & ~(layer0_outputs[2671]);
    assign outputs[960] = layer0_outputs[4170];
    assign outputs[961] = layer0_outputs[3488];
    assign outputs[962] = (layer0_outputs[2824]) | (layer0_outputs[6027]);
    assign outputs[963] = layer0_outputs[9524];
    assign outputs[964] = ~(layer0_outputs[6203]) | (layer0_outputs[3332]);
    assign outputs[965] = ~((layer0_outputs[725]) ^ (layer0_outputs[4529]));
    assign outputs[966] = layer0_outputs[328];
    assign outputs[967] = (layer0_outputs[3997]) & ~(layer0_outputs[3206]);
    assign outputs[968] = ~((layer0_outputs[5538]) | (layer0_outputs[2179]));
    assign outputs[969] = ~(layer0_outputs[5109]);
    assign outputs[970] = ~((layer0_outputs[6422]) ^ (layer0_outputs[8188]));
    assign outputs[971] = ~(layer0_outputs[971]);
    assign outputs[972] = (layer0_outputs[7787]) ^ (layer0_outputs[9429]);
    assign outputs[973] = ~((layer0_outputs[7449]) ^ (layer0_outputs[8020]));
    assign outputs[974] = layer0_outputs[9764];
    assign outputs[975] = (layer0_outputs[3210]) & ~(layer0_outputs[1516]);
    assign outputs[976] = ~((layer0_outputs[1538]) | (layer0_outputs[6319]));
    assign outputs[977] = ~(layer0_outputs[4835]) | (layer0_outputs[1869]);
    assign outputs[978] = ~((layer0_outputs[2779]) ^ (layer0_outputs[9027]));
    assign outputs[979] = layer0_outputs[4698];
    assign outputs[980] = layer0_outputs[5152];
    assign outputs[981] = (layer0_outputs[8448]) & (layer0_outputs[1687]);
    assign outputs[982] = (layer0_outputs[1882]) | (layer0_outputs[5828]);
    assign outputs[983] = ~(layer0_outputs[1995]) | (layer0_outputs[7849]);
    assign outputs[984] = ~(layer0_outputs[874]);
    assign outputs[985] = ~(layer0_outputs[9426]) | (layer0_outputs[6304]);
    assign outputs[986] = (layer0_outputs[8595]) ^ (layer0_outputs[9821]);
    assign outputs[987] = layer0_outputs[3449];
    assign outputs[988] = ~(layer0_outputs[7465]);
    assign outputs[989] = ~(layer0_outputs[8698]);
    assign outputs[990] = ~((layer0_outputs[445]) | (layer0_outputs[4338]));
    assign outputs[991] = (layer0_outputs[4707]) & ~(layer0_outputs[1181]);
    assign outputs[992] = ~(layer0_outputs[5222]);
    assign outputs[993] = ~((layer0_outputs[1410]) ^ (layer0_outputs[810]));
    assign outputs[994] = ~(layer0_outputs[4096]);
    assign outputs[995] = layer0_outputs[5382];
    assign outputs[996] = layer0_outputs[5902];
    assign outputs[997] = (layer0_outputs[3196]) & (layer0_outputs[7437]);
    assign outputs[998] = ~(layer0_outputs[4598]);
    assign outputs[999] = ~((layer0_outputs[1186]) | (layer0_outputs[2734]));
    assign outputs[1000] = (layer0_outputs[1731]) & ~(layer0_outputs[6978]);
    assign outputs[1001] = (layer0_outputs[5678]) ^ (layer0_outputs[9390]);
    assign outputs[1002] = layer0_outputs[311];
    assign outputs[1003] = layer0_outputs[7975];
    assign outputs[1004] = ~(layer0_outputs[5174]);
    assign outputs[1005] = ~(layer0_outputs[7263]);
    assign outputs[1006] = layer0_outputs[1042];
    assign outputs[1007] = layer0_outputs[408];
    assign outputs[1008] = ~(layer0_outputs[429]) | (layer0_outputs[7846]);
    assign outputs[1009] = (layer0_outputs[4400]) | (layer0_outputs[8129]);
    assign outputs[1010] = ~((layer0_outputs[6745]) & (layer0_outputs[4936]));
    assign outputs[1011] = ~(layer0_outputs[4599]) | (layer0_outputs[570]);
    assign outputs[1012] = ~((layer0_outputs[4628]) | (layer0_outputs[7419]));
    assign outputs[1013] = (layer0_outputs[1099]) ^ (layer0_outputs[4770]);
    assign outputs[1014] = ~((layer0_outputs[7678]) & (layer0_outputs[6800]));
    assign outputs[1015] = layer0_outputs[9761];
    assign outputs[1016] = ~(layer0_outputs[5425]);
    assign outputs[1017] = (layer0_outputs[2505]) & ~(layer0_outputs[10155]);
    assign outputs[1018] = ~(layer0_outputs[3494]);
    assign outputs[1019] = ~(layer0_outputs[7161]);
    assign outputs[1020] = layer0_outputs[471];
    assign outputs[1021] = layer0_outputs[10191];
    assign outputs[1022] = layer0_outputs[1741];
    assign outputs[1023] = ~(layer0_outputs[6929]);
    assign outputs[1024] = layer0_outputs[7757];
    assign outputs[1025] = (layer0_outputs[7207]) & ~(layer0_outputs[1618]);
    assign outputs[1026] = (layer0_outputs[9268]) & ~(layer0_outputs[1400]);
    assign outputs[1027] = (layer0_outputs[3370]) & (layer0_outputs[4192]);
    assign outputs[1028] = ~(layer0_outputs[9277]);
    assign outputs[1029] = (layer0_outputs[4271]) & (layer0_outputs[5262]);
    assign outputs[1030] = ~((layer0_outputs[1491]) | (layer0_outputs[5373]));
    assign outputs[1031] = (layer0_outputs[10115]) & ~(layer0_outputs[4060]);
    assign outputs[1032] = (layer0_outputs[6852]) & ~(layer0_outputs[9793]);
    assign outputs[1033] = ~((layer0_outputs[7354]) | (layer0_outputs[5110]));
    assign outputs[1034] = (layer0_outputs[3920]) & ~(layer0_outputs[310]);
    assign outputs[1035] = ~((layer0_outputs[3688]) | (layer0_outputs[4536]));
    assign outputs[1036] = (layer0_outputs[5936]) & (layer0_outputs[10120]);
    assign outputs[1037] = ~((layer0_outputs[59]) ^ (layer0_outputs[7110]));
    assign outputs[1038] = (layer0_outputs[10224]) & ~(layer0_outputs[6034]);
    assign outputs[1039] = (layer0_outputs[5968]) & ~(layer0_outputs[5757]);
    assign outputs[1040] = ~((layer0_outputs[9706]) | (layer0_outputs[6530]));
    assign outputs[1041] = (layer0_outputs[7853]) & ~(layer0_outputs[3142]);
    assign outputs[1042] = (layer0_outputs[7635]) & (layer0_outputs[7267]);
    assign outputs[1043] = (layer0_outputs[5360]) & (layer0_outputs[1193]);
    assign outputs[1044] = layer0_outputs[4320];
    assign outputs[1045] = (layer0_outputs[9475]) & (layer0_outputs[6094]);
    assign outputs[1046] = layer0_outputs[4546];
    assign outputs[1047] = (layer0_outputs[6344]) & ~(layer0_outputs[6518]);
    assign outputs[1048] = layer0_outputs[843];
    assign outputs[1049] = (layer0_outputs[2173]) & ~(layer0_outputs[8418]);
    assign outputs[1050] = ~((layer0_outputs[3226]) ^ (layer0_outputs[5223]));
    assign outputs[1051] = (layer0_outputs[6537]) & ~(layer0_outputs[9953]);
    assign outputs[1052] = (layer0_outputs[4261]) ^ (layer0_outputs[3340]);
    assign outputs[1053] = (layer0_outputs[6470]) ^ (layer0_outputs[6867]);
    assign outputs[1054] = (layer0_outputs[3000]) ^ (layer0_outputs[8965]);
    assign outputs[1055] = (layer0_outputs[1747]) & (layer0_outputs[9112]);
    assign outputs[1056] = ~(layer0_outputs[6184]);
    assign outputs[1057] = ~((layer0_outputs[762]) | (layer0_outputs[3145]));
    assign outputs[1058] = ~((layer0_outputs[2548]) | (layer0_outputs[879]));
    assign outputs[1059] = 1'b0;
    assign outputs[1060] = ~((layer0_outputs[4796]) ^ (layer0_outputs[7293]));
    assign outputs[1061] = layer0_outputs[9431];
    assign outputs[1062] = (layer0_outputs[10213]) & ~(layer0_outputs[6903]);
    assign outputs[1063] = ~((layer0_outputs[6371]) & (layer0_outputs[3479]));
    assign outputs[1064] = 1'b0;
    assign outputs[1065] = (layer0_outputs[2122]) | (layer0_outputs[2355]);
    assign outputs[1066] = ~((layer0_outputs[3323]) | (layer0_outputs[5379]));
    assign outputs[1067] = (layer0_outputs[10067]) & (layer0_outputs[1246]);
    assign outputs[1068] = (layer0_outputs[6004]) ^ (layer0_outputs[6660]);
    assign outputs[1069] = (layer0_outputs[936]) & ~(layer0_outputs[2732]);
    assign outputs[1070] = (layer0_outputs[9165]) ^ (layer0_outputs[8902]);
    assign outputs[1071] = 1'b0;
    assign outputs[1072] = (layer0_outputs[4053]) & (layer0_outputs[6358]);
    assign outputs[1073] = (layer0_outputs[939]) & (layer0_outputs[9725]);
    assign outputs[1074] = (layer0_outputs[3234]) & ~(layer0_outputs[7962]);
    assign outputs[1075] = (layer0_outputs[5976]) & (layer0_outputs[3662]);
    assign outputs[1076] = layer0_outputs[2731];
    assign outputs[1077] = layer0_outputs[9162];
    assign outputs[1078] = (layer0_outputs[9147]) ^ (layer0_outputs[2193]);
    assign outputs[1079] = ~(layer0_outputs[7346]);
    assign outputs[1080] = (layer0_outputs[2551]) ^ (layer0_outputs[1176]);
    assign outputs[1081] = (layer0_outputs[3131]) & ~(layer0_outputs[5253]);
    assign outputs[1082] = ~((layer0_outputs[9605]) | (layer0_outputs[568]));
    assign outputs[1083] = ~((layer0_outputs[4819]) | (layer0_outputs[5941]));
    assign outputs[1084] = (layer0_outputs[5307]) & ~(layer0_outputs[102]);
    assign outputs[1085] = (layer0_outputs[2672]) & (layer0_outputs[6442]);
    assign outputs[1086] = ~((layer0_outputs[888]) | (layer0_outputs[2860]));
    assign outputs[1087] = (layer0_outputs[8659]) & (layer0_outputs[1030]);
    assign outputs[1088] = (layer0_outputs[8087]) & (layer0_outputs[789]);
    assign outputs[1089] = layer0_outputs[8201];
    assign outputs[1090] = (layer0_outputs[2164]) & (layer0_outputs[1749]);
    assign outputs[1091] = (layer0_outputs[6025]) & (layer0_outputs[9870]);
    assign outputs[1092] = layer0_outputs[4524];
    assign outputs[1093] = ~((layer0_outputs[4732]) ^ (layer0_outputs[9453]));
    assign outputs[1094] = ~(layer0_outputs[7704]);
    assign outputs[1095] = ~((layer0_outputs[5103]) | (layer0_outputs[3393]));
    assign outputs[1096] = (layer0_outputs[1932]) & (layer0_outputs[5140]);
    assign outputs[1097] = layer0_outputs[1394];
    assign outputs[1098] = (layer0_outputs[4088]) & ~(layer0_outputs[1723]);
    assign outputs[1099] = ~((layer0_outputs[1261]) | (layer0_outputs[7802]));
    assign outputs[1100] = layer0_outputs[4087];
    assign outputs[1101] = (layer0_outputs[8016]) & (layer0_outputs[1822]);
    assign outputs[1102] = ~(layer0_outputs[2293]);
    assign outputs[1103] = (layer0_outputs[9976]) ^ (layer0_outputs[4993]);
    assign outputs[1104] = ~((layer0_outputs[176]) | (layer0_outputs[4437]));
    assign outputs[1105] = layer0_outputs[5372];
    assign outputs[1106] = ~(layer0_outputs[4737]);
    assign outputs[1107] = (layer0_outputs[8612]) & ~(layer0_outputs[4889]);
    assign outputs[1108] = ~((layer0_outputs[4522]) | (layer0_outputs[3995]));
    assign outputs[1109] = layer0_outputs[6227];
    assign outputs[1110] = (layer0_outputs[1294]) & ~(layer0_outputs[3699]);
    assign outputs[1111] = layer0_outputs[8767];
    assign outputs[1112] = ~(layer0_outputs[1969]);
    assign outputs[1113] = (layer0_outputs[8029]) & ~(layer0_outputs[6121]);
    assign outputs[1114] = ~(layer0_outputs[6343]);
    assign outputs[1115] = (layer0_outputs[2351]) & ~(layer0_outputs[3258]);
    assign outputs[1116] = ~((layer0_outputs[6174]) | (layer0_outputs[1815]));
    assign outputs[1117] = ~((layer0_outputs[2103]) ^ (layer0_outputs[4377]));
    assign outputs[1118] = ~((layer0_outputs[2520]) ^ (layer0_outputs[1184]));
    assign outputs[1119] = layer0_outputs[5340];
    assign outputs[1120] = (layer0_outputs[9146]) & ~(layer0_outputs[6071]);
    assign outputs[1121] = (layer0_outputs[9237]) & ~(layer0_outputs[4538]);
    assign outputs[1122] = layer0_outputs[8097];
    assign outputs[1123] = (layer0_outputs[7571]) & (layer0_outputs[8792]);
    assign outputs[1124] = (layer0_outputs[210]) & ~(layer0_outputs[1906]);
    assign outputs[1125] = ~((layer0_outputs[6412]) ^ (layer0_outputs[6585]));
    assign outputs[1126] = ~((layer0_outputs[611]) | (layer0_outputs[10037]));
    assign outputs[1127] = (layer0_outputs[2814]) ^ (layer0_outputs[670]);
    assign outputs[1128] = ~(layer0_outputs[2033]);
    assign outputs[1129] = (layer0_outputs[4739]) ^ (layer0_outputs[2065]);
    assign outputs[1130] = (layer0_outputs[3317]) & ~(layer0_outputs[3712]);
    assign outputs[1131] = (layer0_outputs[730]) & ~(layer0_outputs[1531]);
    assign outputs[1132] = (layer0_outputs[9980]) ^ (layer0_outputs[3603]);
    assign outputs[1133] = (layer0_outputs[1121]) & ~(layer0_outputs[1453]);
    assign outputs[1134] = ~((layer0_outputs[4844]) | (layer0_outputs[724]));
    assign outputs[1135] = ~(layer0_outputs[7631]);
    assign outputs[1136] = (layer0_outputs[3915]) & ~(layer0_outputs[5468]);
    assign outputs[1137] = ~((layer0_outputs[8165]) | (layer0_outputs[8897]));
    assign outputs[1138] = (layer0_outputs[5028]) & ~(layer0_outputs[6519]);
    assign outputs[1139] = layer0_outputs[3182];
    assign outputs[1140] = ~(layer0_outputs[7164]);
    assign outputs[1141] = (layer0_outputs[3738]) | (layer0_outputs[7428]);
    assign outputs[1142] = ~(layer0_outputs[4008]);
    assign outputs[1143] = (layer0_outputs[4542]) & (layer0_outputs[7629]);
    assign outputs[1144] = ~((layer0_outputs[3867]) | (layer0_outputs[7658]));
    assign outputs[1145] = ~((layer0_outputs[7442]) ^ (layer0_outputs[350]));
    assign outputs[1146] = (layer0_outputs[8541]) & (layer0_outputs[7439]);
    assign outputs[1147] = ~(layer0_outputs[239]) | (layer0_outputs[1532]);
    assign outputs[1148] = ~((layer0_outputs[1792]) ^ (layer0_outputs[2581]));
    assign outputs[1149] = (layer0_outputs[6798]) & (layer0_outputs[5438]);
    assign outputs[1150] = (layer0_outputs[6588]) & ~(layer0_outputs[3816]);
    assign outputs[1151] = (layer0_outputs[9533]) & ~(layer0_outputs[3910]);
    assign outputs[1152] = (layer0_outputs[2345]) & ~(layer0_outputs[5301]);
    assign outputs[1153] = ~(layer0_outputs[3504]);
    assign outputs[1154] = ~(layer0_outputs[7498]);
    assign outputs[1155] = ~((layer0_outputs[8375]) | (layer0_outputs[1716]));
    assign outputs[1156] = (layer0_outputs[5334]) & ~(layer0_outputs[1492]);
    assign outputs[1157] = ~(layer0_outputs[2233]);
    assign outputs[1158] = (layer0_outputs[7430]) ^ (layer0_outputs[5465]);
    assign outputs[1159] = (layer0_outputs[3052]) & ~(layer0_outputs[3926]);
    assign outputs[1160] = layer0_outputs[6372];
    assign outputs[1161] = ~((layer0_outputs[3473]) | (layer0_outputs[6894]));
    assign outputs[1162] = (layer0_outputs[5971]) & (layer0_outputs[3406]);
    assign outputs[1163] = (layer0_outputs[9529]) & (layer0_outputs[4611]);
    assign outputs[1164] = (layer0_outputs[5409]) & ~(layer0_outputs[717]);
    assign outputs[1165] = ~((layer0_outputs[1010]) | (layer0_outputs[306]));
    assign outputs[1166] = ~(layer0_outputs[2664]);
    assign outputs[1167] = (layer0_outputs[3984]) & (layer0_outputs[10051]);
    assign outputs[1168] = (layer0_outputs[3750]) & ~(layer0_outputs[4775]);
    assign outputs[1169] = ~(layer0_outputs[8615]);
    assign outputs[1170] = (layer0_outputs[6441]) & (layer0_outputs[8103]);
    assign outputs[1171] = (layer0_outputs[2516]) & ~(layer0_outputs[6812]);
    assign outputs[1172] = ~(layer0_outputs[10001]);
    assign outputs[1173] = ~((layer0_outputs[7351]) | (layer0_outputs[9275]));
    assign outputs[1174] = ~(layer0_outputs[7727]);
    assign outputs[1175] = (layer0_outputs[8837]) & ~(layer0_outputs[2072]);
    assign outputs[1176] = layer0_outputs[9354];
    assign outputs[1177] = ~(layer0_outputs[6880]);
    assign outputs[1178] = (layer0_outputs[6259]) ^ (layer0_outputs[2164]);
    assign outputs[1179] = (layer0_outputs[2493]) & ~(layer0_outputs[9552]);
    assign outputs[1180] = ~((layer0_outputs[3442]) ^ (layer0_outputs[3830]));
    assign outputs[1181] = (layer0_outputs[4929]) & ~(layer0_outputs[7218]);
    assign outputs[1182] = layer0_outputs[9858];
    assign outputs[1183] = ~(layer0_outputs[449]);
    assign outputs[1184] = ~((layer0_outputs[8189]) | (layer0_outputs[9793]));
    assign outputs[1185] = ~(layer0_outputs[2768]);
    assign outputs[1186] = ~((layer0_outputs[1684]) ^ (layer0_outputs[188]));
    assign outputs[1187] = (layer0_outputs[6252]) ^ (layer0_outputs[1733]);
    assign outputs[1188] = layer0_outputs[1067];
    assign outputs[1189] = ~((layer0_outputs[601]) ^ (layer0_outputs[3361]));
    assign outputs[1190] = layer0_outputs[2604];
    assign outputs[1191] = ~(layer0_outputs[7343]);
    assign outputs[1192] = (layer0_outputs[8648]) & ~(layer0_outputs[3636]);
    assign outputs[1193] = layer0_outputs[10215];
    assign outputs[1194] = (layer0_outputs[1514]) & (layer0_outputs[7835]);
    assign outputs[1195] = (layer0_outputs[1103]) & ~(layer0_outputs[510]);
    assign outputs[1196] = (layer0_outputs[6949]) & ~(layer0_outputs[2370]);
    assign outputs[1197] = (layer0_outputs[1170]) & (layer0_outputs[5299]);
    assign outputs[1198] = ~((layer0_outputs[1921]) | (layer0_outputs[6147]));
    assign outputs[1199] = (layer0_outputs[5773]) & ~(layer0_outputs[7064]);
    assign outputs[1200] = (layer0_outputs[2061]) & ~(layer0_outputs[3873]);
    assign outputs[1201] = (layer0_outputs[1108]) & (layer0_outputs[4904]);
    assign outputs[1202] = ~((layer0_outputs[8936]) | (layer0_outputs[1560]));
    assign outputs[1203] = (layer0_outputs[4081]) ^ (layer0_outputs[9502]);
    assign outputs[1204] = layer0_outputs[9026];
    assign outputs[1205] = (layer0_outputs[5054]) | (layer0_outputs[7590]);
    assign outputs[1206] = (layer0_outputs[8723]) & (layer0_outputs[5213]);
    assign outputs[1207] = 1'b0;
    assign outputs[1208] = (layer0_outputs[4850]) & ~(layer0_outputs[4434]);
    assign outputs[1209] = (layer0_outputs[6647]) ^ (layer0_outputs[3384]);
    assign outputs[1210] = (layer0_outputs[918]) ^ (layer0_outputs[8122]);
    assign outputs[1211] = ~(layer0_outputs[5537]);
    assign outputs[1212] = (layer0_outputs[7579]) & ~(layer0_outputs[2144]);
    assign outputs[1213] = layer0_outputs[5159];
    assign outputs[1214] = (layer0_outputs[1284]) ^ (layer0_outputs[4365]);
    assign outputs[1215] = ~((layer0_outputs[2757]) ^ (layer0_outputs[1712]));
    assign outputs[1216] = (layer0_outputs[575]) & ~(layer0_outputs[1962]);
    assign outputs[1217] = (layer0_outputs[3017]) & ~(layer0_outputs[9918]);
    assign outputs[1218] = layer0_outputs[10167];
    assign outputs[1219] = (layer0_outputs[10108]) & ~(layer0_outputs[5729]);
    assign outputs[1220] = (layer0_outputs[3451]) & ~(layer0_outputs[2096]);
    assign outputs[1221] = ~(layer0_outputs[1589]);
    assign outputs[1222] = ~(layer0_outputs[8453]);
    assign outputs[1223] = (layer0_outputs[878]) & ~(layer0_outputs[70]);
    assign outputs[1224] = layer0_outputs[4876];
    assign outputs[1225] = ~((layer0_outputs[3160]) ^ (layer0_outputs[6440]));
    assign outputs[1226] = (layer0_outputs[7886]) & (layer0_outputs[2128]);
    assign outputs[1227] = (layer0_outputs[6324]) & ~(layer0_outputs[6290]);
    assign outputs[1228] = ~((layer0_outputs[2134]) ^ (layer0_outputs[4669]));
    assign outputs[1229] = ~(layer0_outputs[8902]) | (layer0_outputs[9201]);
    assign outputs[1230] = ~(layer0_outputs[2991]);
    assign outputs[1231] = (layer0_outputs[504]) & ~(layer0_outputs[9517]);
    assign outputs[1232] = ~((layer0_outputs[6354]) ^ (layer0_outputs[1629]));
    assign outputs[1233] = (layer0_outputs[3367]) ^ (layer0_outputs[4238]);
    assign outputs[1234] = ~((layer0_outputs[9583]) ^ (layer0_outputs[7002]));
    assign outputs[1235] = ~((layer0_outputs[6730]) ^ (layer0_outputs[8254]));
    assign outputs[1236] = ~((layer0_outputs[2288]) ^ (layer0_outputs[4295]));
    assign outputs[1237] = layer0_outputs[9063];
    assign outputs[1238] = (layer0_outputs[3173]) ^ (layer0_outputs[8898]);
    assign outputs[1239] = (layer0_outputs[6970]) & ~(layer0_outputs[3952]);
    assign outputs[1240] = ~(layer0_outputs[9514]);
    assign outputs[1241] = (layer0_outputs[5904]) & ~(layer0_outputs[4541]);
    assign outputs[1242] = ~(layer0_outputs[2716]);
    assign outputs[1243] = ~((layer0_outputs[10]) | (layer0_outputs[9312]));
    assign outputs[1244] = ~((layer0_outputs[6686]) | (layer0_outputs[618]));
    assign outputs[1245] = ~((layer0_outputs[3724]) | (layer0_outputs[1107]));
    assign outputs[1246] = (layer0_outputs[1186]) ^ (layer0_outputs[9062]);
    assign outputs[1247] = (layer0_outputs[3148]) & (layer0_outputs[7924]);
    assign outputs[1248] = ~((layer0_outputs[2033]) | (layer0_outputs[1285]));
    assign outputs[1249] = ~(layer0_outputs[6244]);
    assign outputs[1250] = (layer0_outputs[5027]) & ~(layer0_outputs[8501]);
    assign outputs[1251] = (layer0_outputs[1104]) & ~(layer0_outputs[586]);
    assign outputs[1252] = (layer0_outputs[1972]) ^ (layer0_outputs[9284]);
    assign outputs[1253] = ~((layer0_outputs[5941]) | (layer0_outputs[4145]));
    assign outputs[1254] = ~(layer0_outputs[1096]);
    assign outputs[1255] = (layer0_outputs[5644]) & (layer0_outputs[5692]);
    assign outputs[1256] = (layer0_outputs[7529]) & (layer0_outputs[7243]);
    assign outputs[1257] = (layer0_outputs[493]) & ~(layer0_outputs[7117]);
    assign outputs[1258] = ~(layer0_outputs[3502]);
    assign outputs[1259] = (layer0_outputs[5407]) & ~(layer0_outputs[6482]);
    assign outputs[1260] = (layer0_outputs[2795]) ^ (layer0_outputs[8243]);
    assign outputs[1261] = ~((layer0_outputs[8398]) ^ (layer0_outputs[1782]));
    assign outputs[1262] = ~(layer0_outputs[228]);
    assign outputs[1263] = (layer0_outputs[6145]) ^ (layer0_outputs[9344]);
    assign outputs[1264] = (layer0_outputs[4859]) & ~(layer0_outputs[275]);
    assign outputs[1265] = ~(layer0_outputs[4211]);
    assign outputs[1266] = ~(layer0_outputs[6446]);
    assign outputs[1267] = layer0_outputs[1558];
    assign outputs[1268] = (layer0_outputs[6699]) & ~(layer0_outputs[7679]);
    assign outputs[1269] = (layer0_outputs[8248]) ^ (layer0_outputs[1356]);
    assign outputs[1270] = layer0_outputs[9594];
    assign outputs[1271] = ~(layer0_outputs[5731]);
    assign outputs[1272] = (layer0_outputs[7450]) & ~(layer0_outputs[8352]);
    assign outputs[1273] = ~((layer0_outputs[2219]) | (layer0_outputs[4885]));
    assign outputs[1274] = (layer0_outputs[6675]) & ~(layer0_outputs[9065]);
    assign outputs[1275] = (layer0_outputs[4726]) & ~(layer0_outputs[5883]);
    assign outputs[1276] = ~(layer0_outputs[7814]);
    assign outputs[1277] = (layer0_outputs[2923]) & ~(layer0_outputs[9397]);
    assign outputs[1278] = (layer0_outputs[6727]) & (layer0_outputs[9993]);
    assign outputs[1279] = (layer0_outputs[3541]) & (layer0_outputs[7266]);
    assign outputs[1280] = (layer0_outputs[5269]) & ~(layer0_outputs[777]);
    assign outputs[1281] = (layer0_outputs[6756]) & ~(layer0_outputs[3035]);
    assign outputs[1282] = (layer0_outputs[4429]) & (layer0_outputs[7082]);
    assign outputs[1283] = (layer0_outputs[5329]) & ~(layer0_outputs[1513]);
    assign outputs[1284] = ~(layer0_outputs[8154]);
    assign outputs[1285] = (layer0_outputs[4016]) & ~(layer0_outputs[6985]);
    assign outputs[1286] = ~(layer0_outputs[932]);
    assign outputs[1287] = ~((layer0_outputs[4613]) | (layer0_outputs[3299]));
    assign outputs[1288] = (layer0_outputs[4188]) & ~(layer0_outputs[10016]);
    assign outputs[1289] = (layer0_outputs[1671]) & ~(layer0_outputs[7139]);
    assign outputs[1290] = (layer0_outputs[8070]) & (layer0_outputs[4494]);
    assign outputs[1291] = ~(layer0_outputs[10043]);
    assign outputs[1292] = ~((layer0_outputs[9514]) | (layer0_outputs[8957]));
    assign outputs[1293] = (layer0_outputs[2759]) & ~(layer0_outputs[8581]);
    assign outputs[1294] = (layer0_outputs[2927]) & (layer0_outputs[7066]);
    assign outputs[1295] = ~((layer0_outputs[9486]) | (layer0_outputs[4911]));
    assign outputs[1296] = layer0_outputs[9618];
    assign outputs[1297] = ~(layer0_outputs[6410]);
    assign outputs[1298] = (layer0_outputs[5662]) & ~(layer0_outputs[7492]);
    assign outputs[1299] = layer0_outputs[9628];
    assign outputs[1300] = layer0_outputs[4040];
    assign outputs[1301] = (layer0_outputs[662]) ^ (layer0_outputs[4206]);
    assign outputs[1302] = ~((layer0_outputs[8027]) | (layer0_outputs[3756]));
    assign outputs[1303] = (layer0_outputs[4675]) & ~(layer0_outputs[1385]);
    assign outputs[1304] = ~((layer0_outputs[4012]) ^ (layer0_outputs[2749]));
    assign outputs[1305] = (layer0_outputs[9117]) & ~(layer0_outputs[8654]);
    assign outputs[1306] = ~((layer0_outputs[9721]) & (layer0_outputs[4026]));
    assign outputs[1307] = ~((layer0_outputs[9456]) ^ (layer0_outputs[2544]));
    assign outputs[1308] = (layer0_outputs[1617]) & ~(layer0_outputs[1314]);
    assign outputs[1309] = (layer0_outputs[9637]) & ~(layer0_outputs[3516]);
    assign outputs[1310] = ~(layer0_outputs[10040]);
    assign outputs[1311] = (layer0_outputs[856]) & ~(layer0_outputs[3697]);
    assign outputs[1312] = layer0_outputs[3301];
    assign outputs[1313] = (layer0_outputs[6853]) & (layer0_outputs[8578]);
    assign outputs[1314] = 1'b0;
    assign outputs[1315] = (layer0_outputs[9885]) & (layer0_outputs[5560]);
    assign outputs[1316] = (layer0_outputs[9398]) & (layer0_outputs[6713]);
    assign outputs[1317] = (layer0_outputs[9344]) & ~(layer0_outputs[9124]);
    assign outputs[1318] = ~((layer0_outputs[6187]) | (layer0_outputs[207]));
    assign outputs[1319] = ~((layer0_outputs[1544]) ^ (layer0_outputs[32]));
    assign outputs[1320] = (layer0_outputs[9092]) ^ (layer0_outputs[205]);
    assign outputs[1321] = (layer0_outputs[9459]) & ~(layer0_outputs[2022]);
    assign outputs[1322] = (layer0_outputs[184]) & ~(layer0_outputs[3245]);
    assign outputs[1323] = (layer0_outputs[5743]) & ~(layer0_outputs[1937]);
    assign outputs[1324] = (layer0_outputs[10095]) ^ (layer0_outputs[7652]);
    assign outputs[1325] = (layer0_outputs[8030]) ^ (layer0_outputs[8974]);
    assign outputs[1326] = (layer0_outputs[6645]) & ~(layer0_outputs[42]);
    assign outputs[1327] = (layer0_outputs[2481]) & ~(layer0_outputs[9118]);
    assign outputs[1328] = ~((layer0_outputs[4463]) | (layer0_outputs[175]));
    assign outputs[1329] = ~((layer0_outputs[8234]) ^ (layer0_outputs[7070]));
    assign outputs[1330] = (layer0_outputs[9497]) & ~(layer0_outputs[2807]);
    assign outputs[1331] = layer0_outputs[2398];
    assign outputs[1332] = (layer0_outputs[250]) & (layer0_outputs[1490]);
    assign outputs[1333] = ~((layer0_outputs[9336]) ^ (layer0_outputs[9299]));
    assign outputs[1334] = (layer0_outputs[4228]) & ~(layer0_outputs[2428]);
    assign outputs[1335] = (layer0_outputs[8224]) & (layer0_outputs[6736]);
    assign outputs[1336] = (layer0_outputs[8725]) & (layer0_outputs[6550]);
    assign outputs[1337] = (layer0_outputs[8377]) & ~(layer0_outputs[4662]);
    assign outputs[1338] = ~(layer0_outputs[6498]);
    assign outputs[1339] = (layer0_outputs[659]) & (layer0_outputs[2212]);
    assign outputs[1340] = (layer0_outputs[1482]) ^ (layer0_outputs[3602]);
    assign outputs[1341] = (layer0_outputs[6066]) & ~(layer0_outputs[2485]);
    assign outputs[1342] = (layer0_outputs[6073]) ^ (layer0_outputs[5911]);
    assign outputs[1343] = (layer0_outputs[4864]) & ~(layer0_outputs[3887]);
    assign outputs[1344] = ~((layer0_outputs[2804]) ^ (layer0_outputs[9801]));
    assign outputs[1345] = (layer0_outputs[7557]) & ~(layer0_outputs[8039]);
    assign outputs[1346] = ~(layer0_outputs[2077]);
    assign outputs[1347] = ~((layer0_outputs[8436]) | (layer0_outputs[7067]));
    assign outputs[1348] = (layer0_outputs[1938]) & (layer0_outputs[342]);
    assign outputs[1349] = (layer0_outputs[8810]) & ~(layer0_outputs[2427]);
    assign outputs[1350] = (layer0_outputs[4648]) & (layer0_outputs[4646]);
    assign outputs[1351] = (layer0_outputs[8041]) ^ (layer0_outputs[3612]);
    assign outputs[1352] = ~((layer0_outputs[6392]) | (layer0_outputs[2456]));
    assign outputs[1353] = (layer0_outputs[3497]) & ~(layer0_outputs[398]);
    assign outputs[1354] = ~((layer0_outputs[5261]) | (layer0_outputs[5291]));
    assign outputs[1355] = (layer0_outputs[4642]) & ~(layer0_outputs[3420]);
    assign outputs[1356] = (layer0_outputs[2765]) ^ (layer0_outputs[2097]);
    assign outputs[1357] = layer0_outputs[5907];
    assign outputs[1358] = layer0_outputs[8522];
    assign outputs[1359] = ~(layer0_outputs[8139]);
    assign outputs[1360] = (layer0_outputs[8008]) & ~(layer0_outputs[4356]);
    assign outputs[1361] = ~(layer0_outputs[5736]);
    assign outputs[1362] = (layer0_outputs[362]) & ~(layer0_outputs[7510]);
    assign outputs[1363] = (layer0_outputs[7942]) & (layer0_outputs[1926]);
    assign outputs[1364] = (layer0_outputs[6478]) & (layer0_outputs[7222]);
    assign outputs[1365] = ~(layer0_outputs[6548]);
    assign outputs[1366] = (layer0_outputs[7384]) & ~(layer0_outputs[10025]);
    assign outputs[1367] = (layer0_outputs[3118]) & ~(layer0_outputs[2456]);
    assign outputs[1368] = (layer0_outputs[5093]) & ~(layer0_outputs[7517]);
    assign outputs[1369] = (layer0_outputs[901]) & ~(layer0_outputs[8484]);
    assign outputs[1370] = (layer0_outputs[6383]) & ~(layer0_outputs[2450]);
    assign outputs[1371] = (layer0_outputs[7646]) & ~(layer0_outputs[9213]);
    assign outputs[1372] = (layer0_outputs[1426]) & ~(layer0_outputs[8805]);
    assign outputs[1373] = (layer0_outputs[8234]) ^ (layer0_outputs[3587]);
    assign outputs[1374] = ~((layer0_outputs[2899]) ^ (layer0_outputs[3900]));
    assign outputs[1375] = (layer0_outputs[5100]) & ~(layer0_outputs[3305]);
    assign outputs[1376] = ~((layer0_outputs[9966]) | (layer0_outputs[5760]));
    assign outputs[1377] = (layer0_outputs[6140]) & ~(layer0_outputs[8257]);
    assign outputs[1378] = ~((layer0_outputs[7233]) | (layer0_outputs[5493]));
    assign outputs[1379] = ~((layer0_outputs[8014]) | (layer0_outputs[6204]));
    assign outputs[1380] = (layer0_outputs[1695]) & ~(layer0_outputs[1429]);
    assign outputs[1381] = (layer0_outputs[4445]) & ~(layer0_outputs[655]);
    assign outputs[1382] = ~(layer0_outputs[6384]);
    assign outputs[1383] = (layer0_outputs[9391]) & (layer0_outputs[8901]);
    assign outputs[1384] = ~((layer0_outputs[1076]) ^ (layer0_outputs[7166]));
    assign outputs[1385] = (layer0_outputs[2689]) & (layer0_outputs[8716]);
    assign outputs[1386] = layer0_outputs[3589];
    assign outputs[1387] = (layer0_outputs[5302]) ^ (layer0_outputs[9016]);
    assign outputs[1388] = ~((layer0_outputs[8714]) | (layer0_outputs[638]));
    assign outputs[1389] = (layer0_outputs[3183]) ^ (layer0_outputs[2794]);
    assign outputs[1390] = (layer0_outputs[5119]) & ~(layer0_outputs[10035]);
    assign outputs[1391] = ~((layer0_outputs[9922]) ^ (layer0_outputs[5638]));
    assign outputs[1392] = ~((layer0_outputs[9950]) ^ (layer0_outputs[6191]));
    assign outputs[1393] = (layer0_outputs[1201]) ^ (layer0_outputs[3241]);
    assign outputs[1394] = (layer0_outputs[6823]) & ~(layer0_outputs[975]);
    assign outputs[1395] = (layer0_outputs[2939]) & (layer0_outputs[6274]);
    assign outputs[1396] = (layer0_outputs[4326]) & (layer0_outputs[4663]);
    assign outputs[1397] = (layer0_outputs[8730]) & ~(layer0_outputs[7292]);
    assign outputs[1398] = (layer0_outputs[6854]) & ~(layer0_outputs[913]);
    assign outputs[1399] = (layer0_outputs[7222]) | (layer0_outputs[1981]);
    assign outputs[1400] = (layer0_outputs[4589]) & (layer0_outputs[3604]);
    assign outputs[1401] = ~((layer0_outputs[1936]) ^ (layer0_outputs[1297]));
    assign outputs[1402] = ~(layer0_outputs[8226]);
    assign outputs[1403] = ~(layer0_outputs[8529]);
    assign outputs[1404] = ~(layer0_outputs[9640]);
    assign outputs[1405] = (layer0_outputs[6495]) & ~(layer0_outputs[3352]);
    assign outputs[1406] = (layer0_outputs[6023]) & (layer0_outputs[7251]);
    assign outputs[1407] = (layer0_outputs[6158]) & ~(layer0_outputs[5778]);
    assign outputs[1408] = ~(layer0_outputs[9703]);
    assign outputs[1409] = ~(layer0_outputs[5967]);
    assign outputs[1410] = ~((layer0_outputs[5222]) ^ (layer0_outputs[3033]));
    assign outputs[1411] = (layer0_outputs[719]) & ~(layer0_outputs[10085]);
    assign outputs[1412] = ~(layer0_outputs[5923]) | (layer0_outputs[3912]);
    assign outputs[1413] = (layer0_outputs[6396]) & ~(layer0_outputs[4430]);
    assign outputs[1414] = ~((layer0_outputs[7929]) | (layer0_outputs[2620]));
    assign outputs[1415] = (layer0_outputs[6918]) & (layer0_outputs[3122]);
    assign outputs[1416] = (layer0_outputs[4059]) & (layer0_outputs[904]);
    assign outputs[1417] = ~((layer0_outputs[1347]) | (layer0_outputs[2989]));
    assign outputs[1418] = (layer0_outputs[8438]) & ~(layer0_outputs[8890]);
    assign outputs[1419] = ~((layer0_outputs[3816]) | (layer0_outputs[8920]));
    assign outputs[1420] = ~((layer0_outputs[8687]) | (layer0_outputs[4735]));
    assign outputs[1421] = ~((layer0_outputs[8352]) | (layer0_outputs[1040]));
    assign outputs[1422] = (layer0_outputs[45]) & ~(layer0_outputs[4101]);
    assign outputs[1423] = (layer0_outputs[2865]) & (layer0_outputs[4114]);
    assign outputs[1424] = ~((layer0_outputs[5509]) ^ (layer0_outputs[71]));
    assign outputs[1425] = (layer0_outputs[4971]) & (layer0_outputs[7931]);
    assign outputs[1426] = ~((layer0_outputs[9334]) ^ (layer0_outputs[312]));
    assign outputs[1427] = ~(layer0_outputs[8892]);
    assign outputs[1428] = ~((layer0_outputs[3771]) ^ (layer0_outputs[6943]));
    assign outputs[1429] = ~((layer0_outputs[9951]) | (layer0_outputs[5937]));
    assign outputs[1430] = (layer0_outputs[8318]) ^ (layer0_outputs[5482]);
    assign outputs[1431] = ~(layer0_outputs[8552]);
    assign outputs[1432] = (layer0_outputs[8747]) & (layer0_outputs[8945]);
    assign outputs[1433] = layer0_outputs[6803];
    assign outputs[1434] = ~((layer0_outputs[403]) | (layer0_outputs[2227]));
    assign outputs[1435] = (layer0_outputs[5517]) ^ (layer0_outputs[5237]);
    assign outputs[1436] = (layer0_outputs[3809]) ^ (layer0_outputs[6382]);
    assign outputs[1437] = (layer0_outputs[2612]) & ~(layer0_outputs[6260]);
    assign outputs[1438] = (layer0_outputs[1133]) & ~(layer0_outputs[7087]);
    assign outputs[1439] = ~((layer0_outputs[4960]) | (layer0_outputs[2260]));
    assign outputs[1440] = (layer0_outputs[4180]) & ~(layer0_outputs[2559]);
    assign outputs[1441] = (layer0_outputs[7025]) ^ (layer0_outputs[4560]);
    assign outputs[1442] = (layer0_outputs[3458]) & (layer0_outputs[4963]);
    assign outputs[1443] = layer0_outputs[3103];
    assign outputs[1444] = ~((layer0_outputs[2985]) ^ (layer0_outputs[8601]));
    assign outputs[1445] = (layer0_outputs[4330]) & ~(layer0_outputs[6993]);
    assign outputs[1446] = (layer0_outputs[3575]) & (layer0_outputs[4707]);
    assign outputs[1447] = layer0_outputs[4078];
    assign outputs[1448] = (layer0_outputs[2766]) & ~(layer0_outputs[2265]);
    assign outputs[1449] = (layer0_outputs[9585]) & ~(layer0_outputs[5585]);
    assign outputs[1450] = ~((layer0_outputs[7917]) ^ (layer0_outputs[95]));
    assign outputs[1451] = layer0_outputs[8221];
    assign outputs[1452] = layer0_outputs[8832];
    assign outputs[1453] = layer0_outputs[4243];
    assign outputs[1454] = ~(layer0_outputs[7494]);
    assign outputs[1455] = (layer0_outputs[1098]) & (layer0_outputs[174]);
    assign outputs[1456] = 1'b0;
    assign outputs[1457] = (layer0_outputs[1083]) & ~(layer0_outputs[794]);
    assign outputs[1458] = ~(layer0_outputs[10012]);
    assign outputs[1459] = (layer0_outputs[8029]) & ~(layer0_outputs[4673]);
    assign outputs[1460] = (layer0_outputs[1011]) & (layer0_outputs[2380]);
    assign outputs[1461] = 1'b0;
    assign outputs[1462] = (layer0_outputs[7932]) & ~(layer0_outputs[9002]);
    assign outputs[1463] = ~(layer0_outputs[5096]);
    assign outputs[1464] = ~((layer0_outputs[7679]) | (layer0_outputs[9650]));
    assign outputs[1465] = (layer0_outputs[9031]) & ~(layer0_outputs[1478]);
    assign outputs[1466] = (layer0_outputs[9343]) & ~(layer0_outputs[7689]);
    assign outputs[1467] = ~((layer0_outputs[9450]) ^ (layer0_outputs[5634]));
    assign outputs[1468] = (layer0_outputs[3567]) & ~(layer0_outputs[3971]);
    assign outputs[1469] = ~((layer0_outputs[3954]) ^ (layer0_outputs[3346]));
    assign outputs[1470] = (layer0_outputs[1611]) & (layer0_outputs[354]);
    assign outputs[1471] = (layer0_outputs[7558]) & (layer0_outputs[4046]);
    assign outputs[1472] = layer0_outputs[3988];
    assign outputs[1473] = ~((layer0_outputs[848]) | (layer0_outputs[9134]));
    assign outputs[1474] = (layer0_outputs[1903]) ^ (layer0_outputs[3650]);
    assign outputs[1475] = (layer0_outputs[5273]) & (layer0_outputs[5517]);
    assign outputs[1476] = ~((layer0_outputs[7667]) ^ (layer0_outputs[8407]));
    assign outputs[1477] = (layer0_outputs[1800]) & ~(layer0_outputs[3315]);
    assign outputs[1478] = ~(layer0_outputs[9387]);
    assign outputs[1479] = ~((layer0_outputs[2616]) | (layer0_outputs[3670]));
    assign outputs[1480] = (layer0_outputs[1651]) & ~(layer0_outputs[5621]);
    assign outputs[1481] = layer0_outputs[7578];
    assign outputs[1482] = ~((layer0_outputs[10139]) | (layer0_outputs[579]));
    assign outputs[1483] = layer0_outputs[6262];
    assign outputs[1484] = layer0_outputs[4969];
    assign outputs[1485] = ~(layer0_outputs[1582]);
    assign outputs[1486] = ~((layer0_outputs[5234]) | (layer0_outputs[6807]));
    assign outputs[1487] = (layer0_outputs[456]) & (layer0_outputs[3101]);
    assign outputs[1488] = (layer0_outputs[6922]) & ~(layer0_outputs[4380]);
    assign outputs[1489] = (layer0_outputs[1818]) & ~(layer0_outputs[9544]);
    assign outputs[1490] = layer0_outputs[7992];
    assign outputs[1491] = (layer0_outputs[1178]) ^ (layer0_outputs[9337]);
    assign outputs[1492] = ~((layer0_outputs[6778]) ^ (layer0_outputs[3960]));
    assign outputs[1493] = (layer0_outputs[5029]) & ~(layer0_outputs[721]);
    assign outputs[1494] = (layer0_outputs[6005]) & ~(layer0_outputs[2968]);
    assign outputs[1495] = ~((layer0_outputs[10010]) | (layer0_outputs[7476]));
    assign outputs[1496] = ~(layer0_outputs[559]);
    assign outputs[1497] = ~((layer0_outputs[5882]) | (layer0_outputs[6353]));
    assign outputs[1498] = layer0_outputs[4317];
    assign outputs[1499] = layer0_outputs[7078];
    assign outputs[1500] = (layer0_outputs[1151]) & (layer0_outputs[3931]);
    assign outputs[1501] = layer0_outputs[2008];
    assign outputs[1502] = ~((layer0_outputs[10233]) ^ (layer0_outputs[2161]));
    assign outputs[1503] = layer0_outputs[9878];
    assign outputs[1504] = (layer0_outputs[6367]) & (layer0_outputs[7559]);
    assign outputs[1505] = (layer0_outputs[2644]) & ~(layer0_outputs[6845]);
    assign outputs[1506] = (layer0_outputs[8612]) & ~(layer0_outputs[7716]);
    assign outputs[1507] = (layer0_outputs[7900]) & ~(layer0_outputs[2344]);
    assign outputs[1508] = (layer0_outputs[2276]) & ~(layer0_outputs[2829]);
    assign outputs[1509] = ~((layer0_outputs[8657]) | (layer0_outputs[7075]));
    assign outputs[1510] = (layer0_outputs[4115]) & (layer0_outputs[2748]);
    assign outputs[1511] = ~((layer0_outputs[4721]) ^ (layer0_outputs[4051]));
    assign outputs[1512] = ~(layer0_outputs[5417]);
    assign outputs[1513] = (layer0_outputs[5140]) & (layer0_outputs[2912]);
    assign outputs[1514] = (layer0_outputs[3858]) | (layer0_outputs[5004]);
    assign outputs[1515] = ~((layer0_outputs[5919]) | (layer0_outputs[43]));
    assign outputs[1516] = (layer0_outputs[1808]) ^ (layer0_outputs[2681]);
    assign outputs[1517] = (layer0_outputs[309]) ^ (layer0_outputs[10231]);
    assign outputs[1518] = ~(layer0_outputs[9461]);
    assign outputs[1519] = (layer0_outputs[8315]) ^ (layer0_outputs[3398]);
    assign outputs[1520] = (layer0_outputs[5947]) & ~(layer0_outputs[1095]);
    assign outputs[1521] = layer0_outputs[6361];
    assign outputs[1522] = ~((layer0_outputs[3810]) ^ (layer0_outputs[9981]));
    assign outputs[1523] = (layer0_outputs[5863]) & ~(layer0_outputs[1993]);
    assign outputs[1524] = ~((layer0_outputs[8353]) ^ (layer0_outputs[3605]));
    assign outputs[1525] = (layer0_outputs[1879]) & ~(layer0_outputs[8095]);
    assign outputs[1526] = (layer0_outputs[5383]) & (layer0_outputs[4390]);
    assign outputs[1527] = ~((layer0_outputs[4919]) ^ (layer0_outputs[8988]));
    assign outputs[1528] = ~(layer0_outputs[8139]);
    assign outputs[1529] = ~(layer0_outputs[5885]);
    assign outputs[1530] = ~(layer0_outputs[8890]);
    assign outputs[1531] = layer0_outputs[5104];
    assign outputs[1532] = ~((layer0_outputs[1870]) ^ (layer0_outputs[4033]));
    assign outputs[1533] = (layer0_outputs[8527]) & ~(layer0_outputs[3262]);
    assign outputs[1534] = ~((layer0_outputs[8779]) | (layer0_outputs[9307]));
    assign outputs[1535] = ~((layer0_outputs[4380]) ^ (layer0_outputs[965]));
    assign outputs[1536] = (layer0_outputs[6060]) & (layer0_outputs[3614]);
    assign outputs[1537] = ~(layer0_outputs[7295]);
    assign outputs[1538] = ~((layer0_outputs[4206]) | (layer0_outputs[5476]));
    assign outputs[1539] = (layer0_outputs[1674]) & ~(layer0_outputs[4294]);
    assign outputs[1540] = (layer0_outputs[5365]) ^ (layer0_outputs[2677]);
    assign outputs[1541] = (layer0_outputs[8142]) ^ (layer0_outputs[9150]);
    assign outputs[1542] = (layer0_outputs[5588]) & ~(layer0_outputs[8157]);
    assign outputs[1543] = (layer0_outputs[5710]) & ~(layer0_outputs[6777]);
    assign outputs[1544] = ~((layer0_outputs[2801]) ^ (layer0_outputs[7952]));
    assign outputs[1545] = (layer0_outputs[1944]) & (layer0_outputs[4250]);
    assign outputs[1546] = (layer0_outputs[6940]) ^ (layer0_outputs[3265]);
    assign outputs[1547] = layer0_outputs[8522];
    assign outputs[1548] = ~((layer0_outputs[724]) ^ (layer0_outputs[688]));
    assign outputs[1549] = ~((layer0_outputs[10195]) | (layer0_outputs[5836]));
    assign outputs[1550] = (layer0_outputs[241]) & (layer0_outputs[468]);
    assign outputs[1551] = ~(layer0_outputs[3520]);
    assign outputs[1552] = (layer0_outputs[7122]) & ~(layer0_outputs[2895]);
    assign outputs[1553] = ~(layer0_outputs[707]);
    assign outputs[1554] = (layer0_outputs[6199]) ^ (layer0_outputs[676]);
    assign outputs[1555] = layer0_outputs[4914];
    assign outputs[1556] = layer0_outputs[3151];
    assign outputs[1557] = (layer0_outputs[7902]) & ~(layer0_outputs[4731]);
    assign outputs[1558] = (layer0_outputs[9661]) & ~(layer0_outputs[9765]);
    assign outputs[1559] = (layer0_outputs[264]) & ~(layer0_outputs[2989]);
    assign outputs[1560] = ~((layer0_outputs[3519]) | (layer0_outputs[9788]));
    assign outputs[1561] = (layer0_outputs[1022]) & ~(layer0_outputs[2409]);
    assign outputs[1562] = ~(layer0_outputs[9325]);
    assign outputs[1563] = (layer0_outputs[4629]) & ~(layer0_outputs[7076]);
    assign outputs[1564] = (layer0_outputs[7097]) ^ (layer0_outputs[5692]);
    assign outputs[1565] = layer0_outputs[7799];
    assign outputs[1566] = ~((layer0_outputs[6731]) ^ (layer0_outputs[4178]));
    assign outputs[1567] = (layer0_outputs[8784]) & ~(layer0_outputs[4931]);
    assign outputs[1568] = ~((layer0_outputs[9975]) | (layer0_outputs[1407]));
    assign outputs[1569] = (layer0_outputs[4056]) & ~(layer0_outputs[3341]);
    assign outputs[1570] = (layer0_outputs[7935]) ^ (layer0_outputs[170]);
    assign outputs[1571] = (layer0_outputs[7187]) & ~(layer0_outputs[3266]);
    assign outputs[1572] = (layer0_outputs[6089]) & (layer0_outputs[4243]);
    assign outputs[1573] = (layer0_outputs[6743]) | (layer0_outputs[9182]);
    assign outputs[1574] = ~((layer0_outputs[5799]) | (layer0_outputs[4805]));
    assign outputs[1575] = (layer0_outputs[945]) & ~(layer0_outputs[4679]);
    assign outputs[1576] = (layer0_outputs[8223]) & ~(layer0_outputs[2570]);
    assign outputs[1577] = (layer0_outputs[8822]) ^ (layer0_outputs[3771]);
    assign outputs[1578] = (layer0_outputs[105]) & (layer0_outputs[9482]);
    assign outputs[1579] = ~(layer0_outputs[9566]);
    assign outputs[1580] = layer0_outputs[1797];
    assign outputs[1581] = (layer0_outputs[5786]) & (layer0_outputs[1529]);
    assign outputs[1582] = layer0_outputs[9942];
    assign outputs[1583] = (layer0_outputs[7818]) & (layer0_outputs[10221]);
    assign outputs[1584] = ~(layer0_outputs[5460]);
    assign outputs[1585] = ~((layer0_outputs[4060]) ^ (layer0_outputs[7383]));
    assign outputs[1586] = (layer0_outputs[7651]) & ~(layer0_outputs[8790]);
    assign outputs[1587] = (layer0_outputs[5614]) & (layer0_outputs[1659]);
    assign outputs[1588] = (layer0_outputs[4288]) & ~(layer0_outputs[9077]);
    assign outputs[1589] = (layer0_outputs[959]) & (layer0_outputs[7997]);
    assign outputs[1590] = ~(layer0_outputs[1224]);
    assign outputs[1591] = layer0_outputs[6690];
    assign outputs[1592] = (layer0_outputs[3728]) & ~(layer0_outputs[7632]);
    assign outputs[1593] = (layer0_outputs[6092]) & ~(layer0_outputs[9082]);
    assign outputs[1594] = (layer0_outputs[8155]) & ~(layer0_outputs[1064]);
    assign outputs[1595] = (layer0_outputs[5223]) ^ (layer0_outputs[7093]);
    assign outputs[1596] = 1'b0;
    assign outputs[1597] = (layer0_outputs[3660]) & ~(layer0_outputs[5387]);
    assign outputs[1598] = (layer0_outputs[1692]) & (layer0_outputs[9921]);
    assign outputs[1599] = ~((layer0_outputs[8454]) | (layer0_outputs[7097]));
    assign outputs[1600] = (layer0_outputs[8021]) & ~(layer0_outputs[7986]);
    assign outputs[1601] = layer0_outputs[4728];
    assign outputs[1602] = ~((layer0_outputs[3355]) | (layer0_outputs[8729]));
    assign outputs[1603] = (layer0_outputs[8949]) & (layer0_outputs[2639]);
    assign outputs[1604] = ~((layer0_outputs[8640]) | (layer0_outputs[1429]));
    assign outputs[1605] = (layer0_outputs[8965]) & (layer0_outputs[8501]);
    assign outputs[1606] = ~((layer0_outputs[6181]) | (layer0_outputs[9168]));
    assign outputs[1607] = (layer0_outputs[9573]) & ~(layer0_outputs[5798]);
    assign outputs[1608] = 1'b0;
    assign outputs[1609] = ~((layer0_outputs[4660]) | (layer0_outputs[3503]));
    assign outputs[1610] = (layer0_outputs[1917]) & ~(layer0_outputs[73]);
    assign outputs[1611] = layer0_outputs[8148];
    assign outputs[1612] = (layer0_outputs[1276]) & ~(layer0_outputs[9999]);
    assign outputs[1613] = (layer0_outputs[3893]) & ~(layer0_outputs[9091]);
    assign outputs[1614] = ~((layer0_outputs[10087]) | (layer0_outputs[4995]));
    assign outputs[1615] = ~((layer0_outputs[7709]) ^ (layer0_outputs[6227]));
    assign outputs[1616] = layer0_outputs[7974];
    assign outputs[1617] = (layer0_outputs[6163]) ^ (layer0_outputs[4678]);
    assign outputs[1618] = (layer0_outputs[8638]) & ~(layer0_outputs[8752]);
    assign outputs[1619] = (layer0_outputs[6375]) ^ (layer0_outputs[35]);
    assign outputs[1620] = (layer0_outputs[6574]) & ~(layer0_outputs[3501]);
    assign outputs[1621] = (layer0_outputs[2705]) & ~(layer0_outputs[1240]);
    assign outputs[1622] = (layer0_outputs[8875]) ^ (layer0_outputs[172]);
    assign outputs[1623] = (layer0_outputs[165]) ^ (layer0_outputs[10042]);
    assign outputs[1624] = ~(layer0_outputs[4912]);
    assign outputs[1625] = ~(layer0_outputs[1694]);
    assign outputs[1626] = (layer0_outputs[1010]) & (layer0_outputs[8580]);
    assign outputs[1627] = ~((layer0_outputs[1691]) ^ (layer0_outputs[9695]));
    assign outputs[1628] = (layer0_outputs[8042]) ^ (layer0_outputs[4194]);
    assign outputs[1629] = (layer0_outputs[10156]) & ~(layer0_outputs[2781]);
    assign outputs[1630] = layer0_outputs[8378];
    assign outputs[1631] = (layer0_outputs[3490]) & (layer0_outputs[1795]);
    assign outputs[1632] = (layer0_outputs[4254]) & (layer0_outputs[3589]);
    assign outputs[1633] = ~(layer0_outputs[6701]);
    assign outputs[1634] = 1'b0;
    assign outputs[1635] = (layer0_outputs[9963]) & ~(layer0_outputs[9604]);
    assign outputs[1636] = (layer0_outputs[3695]) & (layer0_outputs[10189]);
    assign outputs[1637] = (layer0_outputs[10062]) & ~(layer0_outputs[3715]);
    assign outputs[1638] = (layer0_outputs[3653]) & ~(layer0_outputs[6130]);
    assign outputs[1639] = (layer0_outputs[8021]) & (layer0_outputs[1555]);
    assign outputs[1640] = layer0_outputs[3259];
    assign outputs[1641] = (layer0_outputs[9909]) ^ (layer0_outputs[5366]);
    assign outputs[1642] = (layer0_outputs[1981]) & ~(layer0_outputs[8754]);
    assign outputs[1643] = ~((layer0_outputs[7471]) | (layer0_outputs[8822]));
    assign outputs[1644] = (layer0_outputs[9713]) & (layer0_outputs[3424]);
    assign outputs[1645] = layer0_outputs[9509];
    assign outputs[1646] = layer0_outputs[6759];
    assign outputs[1647] = (layer0_outputs[9074]) ^ (layer0_outputs[6322]);
    assign outputs[1648] = ~(layer0_outputs[69]);
    assign outputs[1649] = (layer0_outputs[3598]) & (layer0_outputs[8301]);
    assign outputs[1650] = (layer0_outputs[1385]) ^ (layer0_outputs[5472]);
    assign outputs[1651] = (layer0_outputs[8047]) & ~(layer0_outputs[4993]);
    assign outputs[1652] = (layer0_outputs[4902]) & ~(layer0_outputs[5986]);
    assign outputs[1653] = (layer0_outputs[6981]) ^ (layer0_outputs[9249]);
    assign outputs[1654] = ~(layer0_outputs[4801]);
    assign outputs[1655] = ~((layer0_outputs[992]) & (layer0_outputs[2088]));
    assign outputs[1656] = (layer0_outputs[3710]) & ~(layer0_outputs[8256]);
    assign outputs[1657] = (layer0_outputs[2041]) & (layer0_outputs[5857]);
    assign outputs[1658] = layer0_outputs[9266];
    assign outputs[1659] = ~((layer0_outputs[781]) ^ (layer0_outputs[1343]));
    assign outputs[1660] = ~((layer0_outputs[4549]) | (layer0_outputs[2832]));
    assign outputs[1661] = ~((layer0_outputs[1101]) | (layer0_outputs[2038]));
    assign outputs[1662] = ~((layer0_outputs[5895]) ^ (layer0_outputs[8771]));
    assign outputs[1663] = ~((layer0_outputs[10089]) ^ (layer0_outputs[30]));
    assign outputs[1664] = (layer0_outputs[10219]) & (layer0_outputs[2308]);
    assign outputs[1665] = ~(layer0_outputs[4474]);
    assign outputs[1666] = layer0_outputs[2326];
    assign outputs[1667] = (layer0_outputs[7521]) ^ (layer0_outputs[863]);
    assign outputs[1668] = (layer0_outputs[198]) & ~(layer0_outputs[2248]);
    assign outputs[1669] = (layer0_outputs[1952]) & ~(layer0_outputs[1486]);
    assign outputs[1670] = ~(layer0_outputs[8212]) | (layer0_outputs[3931]);
    assign outputs[1671] = (layer0_outputs[6688]) & (layer0_outputs[10038]);
    assign outputs[1672] = (layer0_outputs[2857]) & ~(layer0_outputs[8855]);
    assign outputs[1673] = layer0_outputs[2527];
    assign outputs[1674] = ~((layer0_outputs[7317]) | (layer0_outputs[9114]));
    assign outputs[1675] = layer0_outputs[2230];
    assign outputs[1676] = ~(layer0_outputs[6148]) | (layer0_outputs[6052]);
    assign outputs[1677] = ~(layer0_outputs[5553]) | (layer0_outputs[1209]);
    assign outputs[1678] = ~((layer0_outputs[6893]) | (layer0_outputs[8567]));
    assign outputs[1679] = layer0_outputs[9322];
    assign outputs[1680] = (layer0_outputs[5217]) & ~(layer0_outputs[9235]);
    assign outputs[1681] = layer0_outputs[8759];
    assign outputs[1682] = layer0_outputs[7640];
    assign outputs[1683] = (layer0_outputs[5427]) ^ (layer0_outputs[9038]);
    assign outputs[1684] = (layer0_outputs[10002]) & ~(layer0_outputs[6822]);
    assign outputs[1685] = (layer0_outputs[2106]) & (layer0_outputs[1580]);
    assign outputs[1686] = ~(layer0_outputs[4221]);
    assign outputs[1687] = (layer0_outputs[9417]) & ~(layer0_outputs[7155]);
    assign outputs[1688] = ~(layer0_outputs[4023]);
    assign outputs[1689] = layer0_outputs[6762];
    assign outputs[1690] = layer0_outputs[4489];
    assign outputs[1691] = ~((layer0_outputs[4111]) | (layer0_outputs[1025]));
    assign outputs[1692] = layer0_outputs[2902];
    assign outputs[1693] = ~(layer0_outputs[9643]);
    assign outputs[1694] = (layer0_outputs[1397]) & (layer0_outputs[1556]);
    assign outputs[1695] = ~(layer0_outputs[8547]);
    assign outputs[1696] = (layer0_outputs[6230]) & ~(layer0_outputs[249]);
    assign outputs[1697] = (layer0_outputs[4896]) & (layer0_outputs[9423]);
    assign outputs[1698] = (layer0_outputs[10034]) & (layer0_outputs[2823]);
    assign outputs[1699] = (layer0_outputs[2002]) & ~(layer0_outputs[3330]);
    assign outputs[1700] = (layer0_outputs[2361]) & ~(layer0_outputs[8925]);
    assign outputs[1701] = ~((layer0_outputs[8980]) | (layer0_outputs[8962]));
    assign outputs[1702] = 1'b0;
    assign outputs[1703] = (layer0_outputs[2880]) & ~(layer0_outputs[5685]);
    assign outputs[1704] = (layer0_outputs[8966]) & ~(layer0_outputs[8134]);
    assign outputs[1705] = (layer0_outputs[1828]) & ~(layer0_outputs[5852]);
    assign outputs[1706] = ~((layer0_outputs[8784]) ^ (layer0_outputs[9505]));
    assign outputs[1707] = ~(layer0_outputs[814]);
    assign outputs[1708] = ~((layer0_outputs[8607]) | (layer0_outputs[8785]));
    assign outputs[1709] = ~((layer0_outputs[484]) ^ (layer0_outputs[6292]));
    assign outputs[1710] = (layer0_outputs[4466]) & (layer0_outputs[2676]);
    assign outputs[1711] = (layer0_outputs[7964]) ^ (layer0_outputs[1041]);
    assign outputs[1712] = (layer0_outputs[9458]) & ~(layer0_outputs[2786]);
    assign outputs[1713] = ~((layer0_outputs[6323]) ^ (layer0_outputs[928]));
    assign outputs[1714] = (layer0_outputs[375]) & ~(layer0_outputs[9357]);
    assign outputs[1715] = (layer0_outputs[3163]) & ~(layer0_outputs[6851]);
    assign outputs[1716] = (layer0_outputs[3080]) & ~(layer0_outputs[246]);
    assign outputs[1717] = (layer0_outputs[7089]) & ~(layer0_outputs[2322]);
    assign outputs[1718] = (layer0_outputs[973]) & (layer0_outputs[3541]);
    assign outputs[1719] = (layer0_outputs[4014]) & ~(layer0_outputs[380]);
    assign outputs[1720] = ~((layer0_outputs[9233]) | (layer0_outputs[3891]));
    assign outputs[1721] = (layer0_outputs[2235]) & ~(layer0_outputs[7628]);
    assign outputs[1722] = (layer0_outputs[8702]) & ~(layer0_outputs[5378]);
    assign outputs[1723] = ~(layer0_outputs[4241]);
    assign outputs[1724] = layer0_outputs[4941];
    assign outputs[1725] = (layer0_outputs[4743]) & (layer0_outputs[5603]);
    assign outputs[1726] = (layer0_outputs[3623]) & (layer0_outputs[8]);
    assign outputs[1727] = layer0_outputs[2105];
    assign outputs[1728] = (layer0_outputs[7386]) & (layer0_outputs[1044]);
    assign outputs[1729] = (layer0_outputs[963]) & ~(layer0_outputs[6797]);
    assign outputs[1730] = ~(layer0_outputs[1372]);
    assign outputs[1731] = ~(layer0_outputs[2203]);
    assign outputs[1732] = ~((layer0_outputs[2940]) ^ (layer0_outputs[9437]));
    assign outputs[1733] = ~((layer0_outputs[9085]) ^ (layer0_outputs[7348]));
    assign outputs[1734] = (layer0_outputs[3930]) & ~(layer0_outputs[4259]);
    assign outputs[1735] = ~(layer0_outputs[6181]);
    assign outputs[1736] = ~((layer0_outputs[4298]) ^ (layer0_outputs[1713]));
    assign outputs[1737] = 1'b0;
    assign outputs[1738] = ~(layer0_outputs[6916]);
    assign outputs[1739] = layer0_outputs[7927];
    assign outputs[1740] = layer0_outputs[8483];
    assign outputs[1741] = ~((layer0_outputs[8164]) | (layer0_outputs[7514]));
    assign outputs[1742] = (layer0_outputs[8133]) & ~(layer0_outputs[9929]);
    assign outputs[1743] = (layer0_outputs[7369]) & ~(layer0_outputs[3408]);
    assign outputs[1744] = ~((layer0_outputs[2535]) | (layer0_outputs[1765]));
    assign outputs[1745] = (layer0_outputs[139]) & (layer0_outputs[5922]);
    assign outputs[1746] = ~((layer0_outputs[6782]) | (layer0_outputs[1450]));
    assign outputs[1747] = (layer0_outputs[8378]) & (layer0_outputs[9629]);
    assign outputs[1748] = (layer0_outputs[2990]) & (layer0_outputs[8414]);
    assign outputs[1749] = (layer0_outputs[4255]) & ~(layer0_outputs[1908]);
    assign outputs[1750] = ~((layer0_outputs[8159]) | (layer0_outputs[4358]));
    assign outputs[1751] = ~(layer0_outputs[4310]);
    assign outputs[1752] = ~(layer0_outputs[4090]);
    assign outputs[1753] = (layer0_outputs[3884]) & ~(layer0_outputs[1503]);
    assign outputs[1754] = ~(layer0_outputs[5606]);
    assign outputs[1755] = (layer0_outputs[3609]) ^ (layer0_outputs[7317]);
    assign outputs[1756] = ~(layer0_outputs[1216]);
    assign outputs[1757] = (layer0_outputs[1092]) & ~(layer0_outputs[7667]);
    assign outputs[1758] = (layer0_outputs[5849]) & ~(layer0_outputs[5819]);
    assign outputs[1759] = (layer0_outputs[8777]) & ~(layer0_outputs[8959]);
    assign outputs[1760] = layer0_outputs[8680];
    assign outputs[1761] = (layer0_outputs[2549]) & (layer0_outputs[1262]);
    assign outputs[1762] = 1'b0;
    assign outputs[1763] = layer0_outputs[9884];
    assign outputs[1764] = ~((layer0_outputs[4923]) ^ (layer0_outputs[1868]));
    assign outputs[1765] = (layer0_outputs[8243]) & ~(layer0_outputs[9792]);
    assign outputs[1766] = ~((layer0_outputs[9577]) | (layer0_outputs[6279]));
    assign outputs[1767] = (layer0_outputs[3186]) & ~(layer0_outputs[7357]);
    assign outputs[1768] = (layer0_outputs[5872]) & (layer0_outputs[3439]);
    assign outputs[1769] = (layer0_outputs[81]) & ~(layer0_outputs[3000]);
    assign outputs[1770] = (layer0_outputs[9435]) & ~(layer0_outputs[7798]);
    assign outputs[1771] = (layer0_outputs[4957]) & ~(layer0_outputs[9684]);
    assign outputs[1772] = layer0_outputs[8645];
    assign outputs[1773] = (layer0_outputs[8675]) ^ (layer0_outputs[7436]);
    assign outputs[1774] = (layer0_outputs[2179]) & (layer0_outputs[8807]);
    assign outputs[1775] = (layer0_outputs[2901]) ^ (layer0_outputs[5099]);
    assign outputs[1776] = (layer0_outputs[9463]) & (layer0_outputs[10080]);
    assign outputs[1777] = ~((layer0_outputs[2846]) | (layer0_outputs[7501]));
    assign outputs[1778] = (layer0_outputs[8018]) ^ (layer0_outputs[2156]);
    assign outputs[1779] = (layer0_outputs[4828]) & (layer0_outputs[3256]);
    assign outputs[1780] = layer0_outputs[1699];
    assign outputs[1781] = (layer0_outputs[5570]) & (layer0_outputs[9587]);
    assign outputs[1782] = (layer0_outputs[7712]) & ~(layer0_outputs[3248]);
    assign outputs[1783] = (layer0_outputs[5076]) & ~(layer0_outputs[7759]);
    assign outputs[1784] = ~((layer0_outputs[4459]) ^ (layer0_outputs[8048]));
    assign outputs[1785] = (layer0_outputs[9686]) & ~(layer0_outputs[2718]);
    assign outputs[1786] = ~((layer0_outputs[4067]) | (layer0_outputs[5091]));
    assign outputs[1787] = ~((layer0_outputs[5833]) | (layer0_outputs[3178]));
    assign outputs[1788] = (layer0_outputs[233]) & ~(layer0_outputs[6450]);
    assign outputs[1789] = (layer0_outputs[6945]) & ~(layer0_outputs[1809]);
    assign outputs[1790] = ~((layer0_outputs[6430]) | (layer0_outputs[699]));
    assign outputs[1791] = (layer0_outputs[7707]) & (layer0_outputs[6314]);
    assign outputs[1792] = (layer0_outputs[4063]) & (layer0_outputs[9103]);
    assign outputs[1793] = (layer0_outputs[6936]) & (layer0_outputs[9250]);
    assign outputs[1794] = (layer0_outputs[3499]) & ~(layer0_outputs[6316]);
    assign outputs[1795] = (layer0_outputs[10217]) & ~(layer0_outputs[976]);
    assign outputs[1796] = (layer0_outputs[7075]) ^ (layer0_outputs[2220]);
    assign outputs[1797] = (layer0_outputs[5909]) & ~(layer0_outputs[4355]);
    assign outputs[1798] = layer0_outputs[9935];
    assign outputs[1799] = (layer0_outputs[74]) & ~(layer0_outputs[4279]);
    assign outputs[1800] = ~((layer0_outputs[8599]) | (layer0_outputs[7007]));
    assign outputs[1801] = ~((layer0_outputs[465]) | (layer0_outputs[6640]));
    assign outputs[1802] = ~((layer0_outputs[8613]) | (layer0_outputs[4297]));
    assign outputs[1803] = ~((layer0_outputs[8690]) | (layer0_outputs[3254]));
    assign outputs[1804] = ~((layer0_outputs[5036]) ^ (layer0_outputs[3109]));
    assign outputs[1805] = (layer0_outputs[9003]) & ~(layer0_outputs[2788]);
    assign outputs[1806] = (layer0_outputs[1345]) ^ (layer0_outputs[1908]);
    assign outputs[1807] = (layer0_outputs[2552]) & ~(layer0_outputs[215]);
    assign outputs[1808] = ~(layer0_outputs[1380]);
    assign outputs[1809] = ~((layer0_outputs[3315]) | (layer0_outputs[2808]));
    assign outputs[1810] = layer0_outputs[6210];
    assign outputs[1811] = (layer0_outputs[387]) & ~(layer0_outputs[8700]);
    assign outputs[1812] = ~((layer0_outputs[7383]) | (layer0_outputs[8441]));
    assign outputs[1813] = (layer0_outputs[5428]) & ~(layer0_outputs[8256]);
    assign outputs[1814] = (layer0_outputs[7217]) & ~(layer0_outputs[5859]);
    assign outputs[1815] = (layer0_outputs[741]) & ~(layer0_outputs[8231]);
    assign outputs[1816] = ~((layer0_outputs[1018]) | (layer0_outputs[3028]));
    assign outputs[1817] = (layer0_outputs[9783]) & ~(layer0_outputs[4257]);
    assign outputs[1818] = ~(layer0_outputs[7112]);
    assign outputs[1819] = (layer0_outputs[3373]) & ~(layer0_outputs[6474]);
    assign outputs[1820] = ~((layer0_outputs[7808]) | (layer0_outputs[6044]));
    assign outputs[1821] = ~(layer0_outputs[3]);
    assign outputs[1822] = ~(layer0_outputs[791]);
    assign outputs[1823] = layer0_outputs[9424];
    assign outputs[1824] = ~((layer0_outputs[3645]) | (layer0_outputs[5977]));
    assign outputs[1825] = (layer0_outputs[417]) & ~(layer0_outputs[7970]);
    assign outputs[1826] = ~((layer0_outputs[1403]) ^ (layer0_outputs[908]));
    assign outputs[1827] = ~(layer0_outputs[8635]) | (layer0_outputs[7737]);
    assign outputs[1828] = ~((layer0_outputs[9995]) | (layer0_outputs[1794]));
    assign outputs[1829] = layer0_outputs[9083];
    assign outputs[1830] = ~((layer0_outputs[7104]) | (layer0_outputs[7811]));
    assign outputs[1831] = (layer0_outputs[3728]) & (layer0_outputs[2059]);
    assign outputs[1832] = ~(layer0_outputs[7652]);
    assign outputs[1833] = 1'b0;
    assign outputs[1834] = layer0_outputs[587];
    assign outputs[1835] = (layer0_outputs[6278]) ^ (layer0_outputs[7211]);
    assign outputs[1836] = (layer0_outputs[5197]) & (layer0_outputs[6065]);
    assign outputs[1837] = ~((layer0_outputs[1198]) | (layer0_outputs[2411]));
    assign outputs[1838] = layer0_outputs[4710];
    assign outputs[1839] = layer0_outputs[630];
    assign outputs[1840] = ~((layer0_outputs[6119]) ^ (layer0_outputs[5230]));
    assign outputs[1841] = (layer0_outputs[8710]) & ~(layer0_outputs[2294]);
    assign outputs[1842] = (layer0_outputs[3637]) ^ (layer0_outputs[10173]);
    assign outputs[1843] = (layer0_outputs[2859]) & ~(layer0_outputs[3016]);
    assign outputs[1844] = ~((layer0_outputs[803]) | (layer0_outputs[3648]));
    assign outputs[1845] = ~(layer0_outputs[9084]);
    assign outputs[1846] = (layer0_outputs[8278]) & ~(layer0_outputs[7585]);
    assign outputs[1847] = (layer0_outputs[307]) & (layer0_outputs[6138]);
    assign outputs[1848] = (layer0_outputs[5225]) & ~(layer0_outputs[5623]);
    assign outputs[1849] = (layer0_outputs[3375]) & ~(layer0_outputs[5240]);
    assign outputs[1850] = (layer0_outputs[7747]) & ~(layer0_outputs[5807]);
    assign outputs[1851] = (layer0_outputs[5796]) & ~(layer0_outputs[5736]);
    assign outputs[1852] = ~((layer0_outputs[2755]) | (layer0_outputs[2070]));
    assign outputs[1853] = ~((layer0_outputs[5669]) & (layer0_outputs[7981]));
    assign outputs[1854] = (layer0_outputs[3206]) & (layer0_outputs[1132]);
    assign outputs[1855] = ~((layer0_outputs[9213]) | (layer0_outputs[3822]));
    assign outputs[1856] = 1'b0;
    assign outputs[1857] = ~((layer0_outputs[6182]) | (layer0_outputs[6754]));
    assign outputs[1858] = (layer0_outputs[86]) & ~(layer0_outputs[8958]);
    assign outputs[1859] = (layer0_outputs[8002]) & ~(layer0_outputs[1511]);
    assign outputs[1860] = (layer0_outputs[3008]) & ~(layer0_outputs[1760]);
    assign outputs[1861] = (layer0_outputs[6271]) ^ (layer0_outputs[5123]);
    assign outputs[1862] = ~((layer0_outputs[3612]) | (layer0_outputs[9923]));
    assign outputs[1863] = (layer0_outputs[9934]) & (layer0_outputs[8939]);
    assign outputs[1864] = (layer0_outputs[974]) ^ (layer0_outputs[6197]);
    assign outputs[1865] = layer0_outputs[5039];
    assign outputs[1866] = ~((layer0_outputs[657]) ^ (layer0_outputs[4909]));
    assign outputs[1867] = ~((layer0_outputs[9478]) | (layer0_outputs[4780]));
    assign outputs[1868] = (layer0_outputs[7789]) & ~(layer0_outputs[9255]);
    assign outputs[1869] = (layer0_outputs[3702]) ^ (layer0_outputs[6239]);
    assign outputs[1870] = (layer0_outputs[400]) & (layer0_outputs[5314]);
    assign outputs[1871] = (layer0_outputs[4172]) & ~(layer0_outputs[696]);
    assign outputs[1872] = layer0_outputs[5157];
    assign outputs[1873] = ~((layer0_outputs[6082]) ^ (layer0_outputs[3314]));
    assign outputs[1874] = ~(layer0_outputs[806]);
    assign outputs[1875] = ~((layer0_outputs[8499]) | (layer0_outputs[4695]));
    assign outputs[1876] = (layer0_outputs[8732]) & ~(layer0_outputs[1307]);
    assign outputs[1877] = ~(layer0_outputs[3524]) | (layer0_outputs[4708]);
    assign outputs[1878] = (layer0_outputs[328]) ^ (layer0_outputs[8410]);
    assign outputs[1879] = ~((layer0_outputs[6388]) | (layer0_outputs[3782]));
    assign outputs[1880] = (layer0_outputs[4329]) & (layer0_outputs[23]);
    assign outputs[1881] = (layer0_outputs[864]) & ~(layer0_outputs[871]);
    assign outputs[1882] = ~((layer0_outputs[3671]) | (layer0_outputs[642]));
    assign outputs[1883] = (layer0_outputs[712]) & ~(layer0_outputs[3226]);
    assign outputs[1884] = (layer0_outputs[4359]) & (layer0_outputs[4971]);
    assign outputs[1885] = (layer0_outputs[9599]) & ~(layer0_outputs[9835]);
    assign outputs[1886] = (layer0_outputs[8299]) ^ (layer0_outputs[7658]);
    assign outputs[1887] = ~((layer0_outputs[6262]) ^ (layer0_outputs[3091]));
    assign outputs[1888] = (layer0_outputs[1185]) & (layer0_outputs[4852]);
    assign outputs[1889] = ~((layer0_outputs[1252]) | (layer0_outputs[2523]));
    assign outputs[1890] = ~(layer0_outputs[6793]);
    assign outputs[1891] = ~((layer0_outputs[9366]) | (layer0_outputs[6599]));
    assign outputs[1892] = ~((layer0_outputs[1774]) | (layer0_outputs[8539]));
    assign outputs[1893] = (layer0_outputs[7826]) & (layer0_outputs[5918]);
    assign outputs[1894] = layer0_outputs[7335];
    assign outputs[1895] = ~((layer0_outputs[9725]) ^ (layer0_outputs[700]));
    assign outputs[1896] = (layer0_outputs[7245]) & ~(layer0_outputs[2257]);
    assign outputs[1897] = (layer0_outputs[18]) & ~(layer0_outputs[4953]);
    assign outputs[1898] = ~(layer0_outputs[2174]);
    assign outputs[1899] = ~(layer0_outputs[5960]);
    assign outputs[1900] = (layer0_outputs[5079]) & (layer0_outputs[7944]);
    assign outputs[1901] = ~((layer0_outputs[6369]) | (layer0_outputs[6490]));
    assign outputs[1902] = ~(layer0_outputs[3885]);
    assign outputs[1903] = (layer0_outputs[7758]) & ~(layer0_outputs[7416]);
    assign outputs[1904] = ~(layer0_outputs[569]) | (layer0_outputs[7109]);
    assign outputs[1905] = (layer0_outputs[4498]) & ~(layer0_outputs[9139]);
    assign outputs[1906] = ~((layer0_outputs[1393]) | (layer0_outputs[7589]));
    assign outputs[1907] = ~((layer0_outputs[8392]) | (layer0_outputs[1109]));
    assign outputs[1908] = ~(layer0_outputs[6891]);
    assign outputs[1909] = ~((layer0_outputs[1779]) | (layer0_outputs[9736]));
    assign outputs[1910] = (layer0_outputs[441]) & ~(layer0_outputs[486]);
    assign outputs[1911] = ~((layer0_outputs[562]) | (layer0_outputs[2575]));
    assign outputs[1912] = ~((layer0_outputs[5948]) ^ (layer0_outputs[206]));
    assign outputs[1913] = (layer0_outputs[6408]) & (layer0_outputs[5022]);
    assign outputs[1914] = (layer0_outputs[3084]) & ~(layer0_outputs[6297]);
    assign outputs[1915] = ~(layer0_outputs[2723]);
    assign outputs[1916] = ~((layer0_outputs[21]) | (layer0_outputs[8823]));
    assign outputs[1917] = (layer0_outputs[7413]) & ~(layer0_outputs[8957]);
    assign outputs[1918] = ~((layer0_outputs[1079]) | (layer0_outputs[7289]));
    assign outputs[1919] = (layer0_outputs[4722]) & (layer0_outputs[9160]);
    assign outputs[1920] = (layer0_outputs[9803]) & ~(layer0_outputs[4031]);
    assign outputs[1921] = (layer0_outputs[2655]) & ~(layer0_outputs[4125]);
    assign outputs[1922] = layer0_outputs[5056];
    assign outputs[1923] = (layer0_outputs[6740]) & ~(layer0_outputs[9134]);
    assign outputs[1924] = (layer0_outputs[5637]) & (layer0_outputs[5144]);
    assign outputs[1925] = layer0_outputs[6510];
    assign outputs[1926] = ~((layer0_outputs[9279]) & (layer0_outputs[470]));
    assign outputs[1927] = (layer0_outputs[4782]) ^ (layer0_outputs[9447]);
    assign outputs[1928] = ~((layer0_outputs[3255]) ^ (layer0_outputs[4138]));
    assign outputs[1929] = (layer0_outputs[4235]) & (layer0_outputs[6063]);
    assign outputs[1930] = ~((layer0_outputs[951]) ^ (layer0_outputs[1901]));
    assign outputs[1931] = ~((layer0_outputs[426]) | (layer0_outputs[1258]));
    assign outputs[1932] = (layer0_outputs[8155]) & ~(layer0_outputs[3191]);
    assign outputs[1933] = layer0_outputs[6348];
    assign outputs[1934] = ~(layer0_outputs[5858]);
    assign outputs[1935] = (layer0_outputs[7298]) & (layer0_outputs[2416]);
    assign outputs[1936] = (layer0_outputs[6638]) & (layer0_outputs[1609]);
    assign outputs[1937] = (layer0_outputs[8302]) & ~(layer0_outputs[4752]);
    assign outputs[1938] = ~((layer0_outputs[5410]) | (layer0_outputs[8447]));
    assign outputs[1939] = (layer0_outputs[5777]) & (layer0_outputs[299]);
    assign outputs[1940] = (layer0_outputs[1850]) ^ (layer0_outputs[9177]);
    assign outputs[1941] = layer0_outputs[6636];
    assign outputs[1942] = (layer0_outputs[2998]) & ~(layer0_outputs[940]);
    assign outputs[1943] = (layer0_outputs[2852]) & (layer0_outputs[5677]);
    assign outputs[1944] = ~((layer0_outputs[1170]) ^ (layer0_outputs[2]));
    assign outputs[1945] = (layer0_outputs[760]) & ~(layer0_outputs[655]);
    assign outputs[1946] = (layer0_outputs[9625]) & (layer0_outputs[6588]);
    assign outputs[1947] = (layer0_outputs[1570]) & (layer0_outputs[1044]);
    assign outputs[1948] = ~(layer0_outputs[50]);
    assign outputs[1949] = (layer0_outputs[1424]) & ~(layer0_outputs[7870]);
    assign outputs[1950] = ~(layer0_outputs[8760]);
    assign outputs[1951] = (layer0_outputs[8181]) & (layer0_outputs[2314]);
    assign outputs[1952] = (layer0_outputs[4431]) & ~(layer0_outputs[4329]);
    assign outputs[1953] = (layer0_outputs[7401]) & ~(layer0_outputs[4298]);
    assign outputs[1954] = (layer0_outputs[8951]) & ~(layer0_outputs[191]);
    assign outputs[1955] = ~((layer0_outputs[2422]) ^ (layer0_outputs[10105]));
    assign outputs[1956] = (layer0_outputs[5982]) & (layer0_outputs[5527]);
    assign outputs[1957] = (layer0_outputs[3221]) & (layer0_outputs[2594]);
    assign outputs[1958] = (layer0_outputs[1633]) & (layer0_outputs[6582]);
    assign outputs[1959] = (layer0_outputs[1973]) & ~(layer0_outputs[9140]);
    assign outputs[1960] = (layer0_outputs[445]) & ~(layer0_outputs[6331]);
    assign outputs[1961] = (layer0_outputs[853]) ^ (layer0_outputs[7982]);
    assign outputs[1962] = ~((layer0_outputs[7022]) ^ (layer0_outputs[2057]));
    assign outputs[1963] = ~(layer0_outputs[3788]);
    assign outputs[1964] = layer0_outputs[2068];
    assign outputs[1965] = layer0_outputs[7486];
    assign outputs[1966] = (layer0_outputs[6167]) ^ (layer0_outputs[9843]);
    assign outputs[1967] = (layer0_outputs[6960]) & (layer0_outputs[136]);
    assign outputs[1968] = (layer0_outputs[4864]) & ~(layer0_outputs[3817]);
    assign outputs[1969] = ~((layer0_outputs[6107]) | (layer0_outputs[2430]));
    assign outputs[1970] = (layer0_outputs[9729]) & ~(layer0_outputs[8830]);
    assign outputs[1971] = (layer0_outputs[7240]) & (layer0_outputs[8049]);
    assign outputs[1972] = layer0_outputs[3650];
    assign outputs[1973] = (layer0_outputs[6057]) & ~(layer0_outputs[4609]);
    assign outputs[1974] = ~((layer0_outputs[1698]) | (layer0_outputs[8160]));
    assign outputs[1975] = (layer0_outputs[9356]) & ~(layer0_outputs[598]);
    assign outputs[1976] = (layer0_outputs[9211]) & ~(layer0_outputs[9062]);
    assign outputs[1977] = (layer0_outputs[1785]) & (layer0_outputs[3604]);
    assign outputs[1978] = ~((layer0_outputs[4791]) ^ (layer0_outputs[4433]));
    assign outputs[1979] = ~((layer0_outputs[1530]) ^ (layer0_outputs[4663]));
    assign outputs[1980] = (layer0_outputs[6622]) & ~(layer0_outputs[639]);
    assign outputs[1981] = ~((layer0_outputs[9033]) ^ (layer0_outputs[892]));
    assign outputs[1982] = (layer0_outputs[2885]) & ~(layer0_outputs[8589]);
    assign outputs[1983] = ~((layer0_outputs[3676]) | (layer0_outputs[9425]));
    assign outputs[1984] = ~(layer0_outputs[10182]);
    assign outputs[1985] = (layer0_outputs[755]) & ~(layer0_outputs[5495]);
    assign outputs[1986] = ~((layer0_outputs[294]) ^ (layer0_outputs[8309]));
    assign outputs[1987] = ~((layer0_outputs[5266]) | (layer0_outputs[179]));
    assign outputs[1988] = 1'b0;
    assign outputs[1989] = ~(layer0_outputs[3048]);
    assign outputs[1990] = ~((layer0_outputs[4870]) | (layer0_outputs[2091]));
    assign outputs[1991] = (layer0_outputs[4246]) & ~(layer0_outputs[4979]);
    assign outputs[1992] = layer0_outputs[6198];
    assign outputs[1993] = 1'b0;
    assign outputs[1994] = ~((layer0_outputs[9773]) | (layer0_outputs[8531]));
    assign outputs[1995] = (layer0_outputs[6069]) & ~(layer0_outputs[4441]);
    assign outputs[1996] = (layer0_outputs[2627]) & (layer0_outputs[99]);
    assign outputs[1997] = ~(layer0_outputs[1669]);
    assign outputs[1998] = ~((layer0_outputs[3619]) | (layer0_outputs[4907]));
    assign outputs[1999] = ~(layer0_outputs[8476]);
    assign outputs[2000] = layer0_outputs[1781];
    assign outputs[2001] = (layer0_outputs[7575]) & ~(layer0_outputs[2995]);
    assign outputs[2002] = ~((layer0_outputs[10029]) ^ (layer0_outputs[521]));
    assign outputs[2003] = (layer0_outputs[2127]) & (layer0_outputs[3154]);
    assign outputs[2004] = layer0_outputs[211];
    assign outputs[2005] = (layer0_outputs[5471]) & ~(layer0_outputs[10004]);
    assign outputs[2006] = (layer0_outputs[9708]) & ~(layer0_outputs[1430]);
    assign outputs[2007] = ~(layer0_outputs[808]);
    assign outputs[2008] = layer0_outputs[1528];
    assign outputs[2009] = ~((layer0_outputs[6531]) | (layer0_outputs[6818]));
    assign outputs[2010] = 1'b0;
    assign outputs[2011] = (layer0_outputs[1481]) & ~(layer0_outputs[6980]);
    assign outputs[2012] = 1'b0;
    assign outputs[2013] = (layer0_outputs[4851]) & ~(layer0_outputs[5007]);
    assign outputs[2014] = (layer0_outputs[4703]) & ~(layer0_outputs[1771]);
    assign outputs[2015] = (layer0_outputs[4826]) & ~(layer0_outputs[2550]);
    assign outputs[2016] = ~((layer0_outputs[2426]) | (layer0_outputs[8073]));
    assign outputs[2017] = (layer0_outputs[9106]) & ~(layer0_outputs[8050]);
    assign outputs[2018] = (layer0_outputs[9495]) & ~(layer0_outputs[6719]);
    assign outputs[2019] = ~((layer0_outputs[4844]) | (layer0_outputs[8863]));
    assign outputs[2020] = layer0_outputs[1126];
    assign outputs[2021] = (layer0_outputs[5287]) & ~(layer0_outputs[8987]);
    assign outputs[2022] = layer0_outputs[5586];
    assign outputs[2023] = (layer0_outputs[104]) & ~(layer0_outputs[330]);
    assign outputs[2024] = ~(layer0_outputs[2022]);
    assign outputs[2025] = (layer0_outputs[5026]) & ~(layer0_outputs[7409]);
    assign outputs[2026] = ~(layer0_outputs[6770]) | (layer0_outputs[2291]);
    assign outputs[2027] = (layer0_outputs[5521]) & ~(layer0_outputs[5136]);
    assign outputs[2028] = (layer0_outputs[1299]) ^ (layer0_outputs[6121]);
    assign outputs[2029] = ~(layer0_outputs[1451]);
    assign outputs[2030] = layer0_outputs[998];
    assign outputs[2031] = (layer0_outputs[7874]) & (layer0_outputs[897]);
    assign outputs[2032] = layer0_outputs[333];
    assign outputs[2033] = (layer0_outputs[7812]) & ~(layer0_outputs[6103]);
    assign outputs[2034] = (layer0_outputs[6312]) & ~(layer0_outputs[4109]);
    assign outputs[2035] = layer0_outputs[8162];
    assign outputs[2036] = (layer0_outputs[7914]) & ~(layer0_outputs[5098]);
    assign outputs[2037] = (layer0_outputs[8370]) & ~(layer0_outputs[4179]);
    assign outputs[2038] = ~(layer0_outputs[4959]) | (layer0_outputs[4646]);
    assign outputs[2039] = (layer0_outputs[9015]) & (layer0_outputs[1157]);
    assign outputs[2040] = (layer0_outputs[3347]) & (layer0_outputs[6124]);
    assign outputs[2041] = (layer0_outputs[5933]) ^ (layer0_outputs[8970]);
    assign outputs[2042] = ~((layer0_outputs[5518]) | (layer0_outputs[6648]));
    assign outputs[2043] = ~((layer0_outputs[9436]) | (layer0_outputs[6952]));
    assign outputs[2044] = (layer0_outputs[6633]) & (layer0_outputs[1411]);
    assign outputs[2045] = (layer0_outputs[3194]) & ~(layer0_outputs[5651]);
    assign outputs[2046] = ~(layer0_outputs[6704]);
    assign outputs[2047] = (layer0_outputs[8757]) ^ (layer0_outputs[4073]);
    assign outputs[2048] = ~(layer0_outputs[8502]);
    assign outputs[2049] = ~(layer0_outputs[9561]) | (layer0_outputs[2242]);
    assign outputs[2050] = ~(layer0_outputs[8939]);
    assign outputs[2051] = (layer0_outputs[5758]) | (layer0_outputs[3720]);
    assign outputs[2052] = ~(layer0_outputs[3594]);
    assign outputs[2053] = ~(layer0_outputs[2870]) | (layer0_outputs[6320]);
    assign outputs[2054] = ~(layer0_outputs[9109]);
    assign outputs[2055] = ~(layer0_outputs[6811]);
    assign outputs[2056] = layer0_outputs[7107];
    assign outputs[2057] = (layer0_outputs[1816]) ^ (layer0_outputs[9656]);
    assign outputs[2058] = ~(layer0_outputs[1185]);
    assign outputs[2059] = ~((layer0_outputs[1750]) ^ (layer0_outputs[3885]));
    assign outputs[2060] = ~(layer0_outputs[1589]);
    assign outputs[2061] = layer0_outputs[7125];
    assign outputs[2062] = layer0_outputs[638];
    assign outputs[2063] = layer0_outputs[7427];
    assign outputs[2064] = ~(layer0_outputs[6651]) | (layer0_outputs[1129]);
    assign outputs[2065] = ~(layer0_outputs[316]) | (layer0_outputs[4617]);
    assign outputs[2066] = layer0_outputs[4889];
    assign outputs[2067] = ~(layer0_outputs[8200]);
    assign outputs[2068] = (layer0_outputs[2636]) ^ (layer0_outputs[9546]);
    assign outputs[2069] = ~(layer0_outputs[8071]);
    assign outputs[2070] = ~((layer0_outputs[4202]) | (layer0_outputs[3760]));
    assign outputs[2071] = layer0_outputs[54];
    assign outputs[2072] = (layer0_outputs[6595]) ^ (layer0_outputs[10023]);
    assign outputs[2073] = (layer0_outputs[9697]) ^ (layer0_outputs[6138]);
    assign outputs[2074] = ~(layer0_outputs[6019]) | (layer0_outputs[903]);
    assign outputs[2075] = ~((layer0_outputs[4962]) ^ (layer0_outputs[8462]));
    assign outputs[2076] = ~(layer0_outputs[7418]);
    assign outputs[2077] = (layer0_outputs[6462]) ^ (layer0_outputs[2557]);
    assign outputs[2078] = ~(layer0_outputs[2125]);
    assign outputs[2079] = (layer0_outputs[8253]) & ~(layer0_outputs[3326]);
    assign outputs[2080] = ~((layer0_outputs[9185]) ^ (layer0_outputs[5380]));
    assign outputs[2081] = ~((layer0_outputs[4432]) & (layer0_outputs[5674]));
    assign outputs[2082] = layer0_outputs[8704];
    assign outputs[2083] = ~((layer0_outputs[4558]) ^ (layer0_outputs[9125]));
    assign outputs[2084] = ~(layer0_outputs[5574]);
    assign outputs[2085] = ~(layer0_outputs[7485]);
    assign outputs[2086] = (layer0_outputs[1592]) & ~(layer0_outputs[7650]);
    assign outputs[2087] = ~(layer0_outputs[21]);
    assign outputs[2088] = (layer0_outputs[6397]) ^ (layer0_outputs[2545]);
    assign outputs[2089] = ~((layer0_outputs[5652]) ^ (layer0_outputs[2473]));
    assign outputs[2090] = (layer0_outputs[4068]) | (layer0_outputs[9165]);
    assign outputs[2091] = ~(layer0_outputs[3145]);
    assign outputs[2092] = (layer0_outputs[1381]) ^ (layer0_outputs[9257]);
    assign outputs[2093] = ~(layer0_outputs[1141]);
    assign outputs[2094] = ~(layer0_outputs[2054]);
    assign outputs[2095] = layer0_outputs[5129];
    assign outputs[2096] = ~(layer0_outputs[9740]);
    assign outputs[2097] = ~(layer0_outputs[5608]) | (layer0_outputs[4218]);
    assign outputs[2098] = ~(layer0_outputs[1936]);
    assign outputs[2099] = ~((layer0_outputs[4868]) | (layer0_outputs[1740]));
    assign outputs[2100] = (layer0_outputs[5667]) ^ (layer0_outputs[5766]);
    assign outputs[2101] = ~(layer0_outputs[5000]);
    assign outputs[2102] = layer0_outputs[9150];
    assign outputs[2103] = (layer0_outputs[3031]) | (layer0_outputs[7756]);
    assign outputs[2104] = ~((layer0_outputs[2905]) ^ (layer0_outputs[991]));
    assign outputs[2105] = ~(layer0_outputs[816]);
    assign outputs[2106] = layer0_outputs[9512];
    assign outputs[2107] = ~(layer0_outputs[8933]);
    assign outputs[2108] = (layer0_outputs[3041]) & (layer0_outputs[9897]);
    assign outputs[2109] = ~(layer0_outputs[5452]);
    assign outputs[2110] = layer0_outputs[3045];
    assign outputs[2111] = (layer0_outputs[2300]) & ~(layer0_outputs[8344]);
    assign outputs[2112] = ~((layer0_outputs[6116]) & (layer0_outputs[6361]));
    assign outputs[2113] = (layer0_outputs[4535]) & ~(layer0_outputs[5045]);
    assign outputs[2114] = ~((layer0_outputs[9758]) ^ (layer0_outputs[5825]));
    assign outputs[2115] = ~(layer0_outputs[7683]);
    assign outputs[2116] = layer0_outputs[5277];
    assign outputs[2117] = layer0_outputs[1449];
    assign outputs[2118] = ~((layer0_outputs[9876]) & (layer0_outputs[1868]));
    assign outputs[2119] = ~(layer0_outputs[4988]);
    assign outputs[2120] = ~(layer0_outputs[9901]);
    assign outputs[2121] = (layer0_outputs[276]) ^ (layer0_outputs[3113]);
    assign outputs[2122] = ~((layer0_outputs[9057]) & (layer0_outputs[8002]));
    assign outputs[2123] = layer0_outputs[615];
    assign outputs[2124] = ~((layer0_outputs[3590]) ^ (layer0_outputs[324]));
    assign outputs[2125] = layer0_outputs[9407];
    assign outputs[2126] = layer0_outputs[6011];
    assign outputs[2127] = layer0_outputs[1066];
    assign outputs[2128] = layer0_outputs[2642];
    assign outputs[2129] = ~((layer0_outputs[8116]) | (layer0_outputs[584]));
    assign outputs[2130] = ~((layer0_outputs[5194]) & (layer0_outputs[1703]));
    assign outputs[2131] = ~(layer0_outputs[226]) | (layer0_outputs[4900]);
    assign outputs[2132] = (layer0_outputs[5046]) ^ (layer0_outputs[9989]);
    assign outputs[2133] = ~(layer0_outputs[1596]);
    assign outputs[2134] = ~((layer0_outputs[4021]) ^ (layer0_outputs[3775]));
    assign outputs[2135] = ~(layer0_outputs[3820]);
    assign outputs[2136] = layer0_outputs[10028];
    assign outputs[2137] = ~((layer0_outputs[272]) ^ (layer0_outputs[4563]));
    assign outputs[2138] = ~((layer0_outputs[1311]) & (layer0_outputs[7806]));
    assign outputs[2139] = ~(layer0_outputs[3455]) | (layer0_outputs[3839]);
    assign outputs[2140] = ~(layer0_outputs[7525]) | (layer0_outputs[6342]);
    assign outputs[2141] = (layer0_outputs[2554]) ^ (layer0_outputs[9116]);
    assign outputs[2142] = layer0_outputs[9289];
    assign outputs[2143] = layer0_outputs[194];
    assign outputs[2144] = layer0_outputs[7984];
    assign outputs[2145] = layer0_outputs[7106];
    assign outputs[2146] = (layer0_outputs[2738]) & (layer0_outputs[8339]);
    assign outputs[2147] = ~((layer0_outputs[2040]) ^ (layer0_outputs[3421]));
    assign outputs[2148] = layer0_outputs[4845];
    assign outputs[2149] = ~((layer0_outputs[8316]) ^ (layer0_outputs[57]));
    assign outputs[2150] = (layer0_outputs[5605]) & ~(layer0_outputs[7743]);
    assign outputs[2151] = layer0_outputs[2887];
    assign outputs[2152] = ~((layer0_outputs[7778]) ^ (layer0_outputs[2695]));
    assign outputs[2153] = ~((layer0_outputs[4693]) ^ (layer0_outputs[4324]));
    assign outputs[2154] = layer0_outputs[7015];
    assign outputs[2155] = ~(layer0_outputs[258]) | (layer0_outputs[3430]);
    assign outputs[2156] = ~(layer0_outputs[3492]);
    assign outputs[2157] = layer0_outputs[6202];
    assign outputs[2158] = (layer0_outputs[1211]) ^ (layer0_outputs[939]);
    assign outputs[2159] = ~(layer0_outputs[8835]);
    assign outputs[2160] = layer0_outputs[7469];
    assign outputs[2161] = ~((layer0_outputs[5354]) ^ (layer0_outputs[9939]));
    assign outputs[2162] = layer0_outputs[1081];
    assign outputs[2163] = ~(layer0_outputs[3695]);
    assign outputs[2164] = ~(layer0_outputs[6723]);
    assign outputs[2165] = ~(layer0_outputs[5850]);
    assign outputs[2166] = ~(layer0_outputs[4526]) | (layer0_outputs[2449]);
    assign outputs[2167] = ~((layer0_outputs[4839]) ^ (layer0_outputs[9492]));
    assign outputs[2168] = layer0_outputs[5033];
    assign outputs[2169] = ~(layer0_outputs[6965]) | (layer0_outputs[2171]);
    assign outputs[2170] = ~(layer0_outputs[4982]);
    assign outputs[2171] = ~(layer0_outputs[4897]);
    assign outputs[2172] = ~((layer0_outputs[6127]) & (layer0_outputs[8681]));
    assign outputs[2173] = ~((layer0_outputs[3189]) ^ (layer0_outputs[6917]));
    assign outputs[2174] = ~(layer0_outputs[5826]);
    assign outputs[2175] = ~(layer0_outputs[2019]) | (layer0_outputs[5722]);
    assign outputs[2176] = layer0_outputs[668];
    assign outputs[2177] = layer0_outputs[1680];
    assign outputs[2178] = ~(layer0_outputs[9732]);
    assign outputs[2179] = ~((layer0_outputs[1928]) | (layer0_outputs[2784]));
    assign outputs[2180] = layer0_outputs[2614];
    assign outputs[2181] = ~(layer0_outputs[2185]) | (layer0_outputs[2346]);
    assign outputs[2182] = ~((layer0_outputs[3794]) ^ (layer0_outputs[7318]));
    assign outputs[2183] = layer0_outputs[5462];
    assign outputs[2184] = ~((layer0_outputs[4367]) ^ (layer0_outputs[10031]));
    assign outputs[2185] = ~(layer0_outputs[6551]);
    assign outputs[2186] = layer0_outputs[8408];
    assign outputs[2187] = (layer0_outputs[9438]) & ~(layer0_outputs[9240]);
    assign outputs[2188] = ~(layer0_outputs[2319]);
    assign outputs[2189] = layer0_outputs[2670];
    assign outputs[2190] = (layer0_outputs[1939]) | (layer0_outputs[6676]);
    assign outputs[2191] = (layer0_outputs[4423]) & ~(layer0_outputs[10053]);
    assign outputs[2192] = ~(layer0_outputs[816]);
    assign outputs[2193] = ~((layer0_outputs[1804]) ^ (layer0_outputs[10134]));
    assign outputs[2194] = 1'b1;
    assign outputs[2195] = (layer0_outputs[2757]) ^ (layer0_outputs[8667]);
    assign outputs[2196] = ~(layer0_outputs[3421]);
    assign outputs[2197] = ~(layer0_outputs[5174]);
    assign outputs[2198] = (layer0_outputs[954]) ^ (layer0_outputs[9680]);
    assign outputs[2199] = ~(layer0_outputs[9244]);
    assign outputs[2200] = layer0_outputs[503];
    assign outputs[2201] = ~(layer0_outputs[6080]);
    assign outputs[2202] = ~(layer0_outputs[2957]);
    assign outputs[2203] = ~(layer0_outputs[7774]);
    assign outputs[2204] = ~(layer0_outputs[6440]);
    assign outputs[2205] = ~(layer0_outputs[1653]) | (layer0_outputs[7575]);
    assign outputs[2206] = layer0_outputs[5453];
    assign outputs[2207] = ~((layer0_outputs[1439]) & (layer0_outputs[7827]));
    assign outputs[2208] = layer0_outputs[2855];
    assign outputs[2209] = ~(layer0_outputs[833]);
    assign outputs[2210] = (layer0_outputs[2410]) ^ (layer0_outputs[2465]);
    assign outputs[2211] = ~(layer0_outputs[1248]);
    assign outputs[2212] = (layer0_outputs[3136]) ^ (layer0_outputs[9803]);
    assign outputs[2213] = (layer0_outputs[9823]) & ~(layer0_outputs[9074]);
    assign outputs[2214] = layer0_outputs[2398];
    assign outputs[2215] = (layer0_outputs[2103]) ^ (layer0_outputs[10089]);
    assign outputs[2216] = ~(layer0_outputs[10098]);
    assign outputs[2217] = ~(layer0_outputs[1552]);
    assign outputs[2218] = ~(layer0_outputs[3079]);
    assign outputs[2219] = (layer0_outputs[5405]) & ~(layer0_outputs[7599]);
    assign outputs[2220] = layer0_outputs[8576];
    assign outputs[2221] = ~(layer0_outputs[4720]);
    assign outputs[2222] = (layer0_outputs[2324]) | (layer0_outputs[7017]);
    assign outputs[2223] = ~(layer0_outputs[2659]);
    assign outputs[2224] = layer0_outputs[1123];
    assign outputs[2225] = ~(layer0_outputs[4256]);
    assign outputs[2226] = ~(layer0_outputs[1027]) | (layer0_outputs[5856]);
    assign outputs[2227] = ~((layer0_outputs[6904]) & (layer0_outputs[7382]));
    assign outputs[2228] = ~(layer0_outputs[6345]);
    assign outputs[2229] = ~(layer0_outputs[4695]);
    assign outputs[2230] = (layer0_outputs[2684]) ^ (layer0_outputs[4386]);
    assign outputs[2231] = (layer0_outputs[9125]) & ~(layer0_outputs[3014]);
    assign outputs[2232] = ~(layer0_outputs[9734]);
    assign outputs[2233] = (layer0_outputs[8527]) & ~(layer0_outputs[906]);
    assign outputs[2234] = ~(layer0_outputs[2442]);
    assign outputs[2235] = ~(layer0_outputs[9838]);
    assign outputs[2236] = (layer0_outputs[685]) & (layer0_outputs[6129]);
    assign outputs[2237] = ~((layer0_outputs[6288]) ^ (layer0_outputs[9236]));
    assign outputs[2238] = layer0_outputs[2196];
    assign outputs[2239] = (layer0_outputs[4503]) | (layer0_outputs[1138]);
    assign outputs[2240] = ~(layer0_outputs[4052]) | (layer0_outputs[1436]);
    assign outputs[2241] = layer0_outputs[5921];
    assign outputs[2242] = (layer0_outputs[1422]) ^ (layer0_outputs[312]);
    assign outputs[2243] = (layer0_outputs[6386]) & (layer0_outputs[7602]);
    assign outputs[2244] = (layer0_outputs[3625]) ^ (layer0_outputs[7786]);
    assign outputs[2245] = (layer0_outputs[34]) ^ (layer0_outputs[847]);
    assign outputs[2246] = layer0_outputs[9948];
    assign outputs[2247] = layer0_outputs[8163];
    assign outputs[2248] = layer0_outputs[8584];
    assign outputs[2249] = ~(layer0_outputs[7885]);
    assign outputs[2250] = ~(layer0_outputs[5300]);
    assign outputs[2251] = layer0_outputs[9431];
    assign outputs[2252] = ~((layer0_outputs[8937]) ^ (layer0_outputs[9819]));
    assign outputs[2253] = ~((layer0_outputs[3182]) ^ (layer0_outputs[7708]));
    assign outputs[2254] = ~(layer0_outputs[3838]);
    assign outputs[2255] = layer0_outputs[5438];
    assign outputs[2256] = ~(layer0_outputs[9187]) | (layer0_outputs[520]);
    assign outputs[2257] = ~(layer0_outputs[397]) | (layer0_outputs[260]);
    assign outputs[2258] = ~(layer0_outputs[4727]);
    assign outputs[2259] = layer0_outputs[7206];
    assign outputs[2260] = ~(layer0_outputs[6432]);
    assign outputs[2261] = layer0_outputs[4061];
    assign outputs[2262] = ~((layer0_outputs[2020]) & (layer0_outputs[5782]));
    assign outputs[2263] = ~(layer0_outputs[2403]);
    assign outputs[2264] = (layer0_outputs[3271]) & (layer0_outputs[6327]);
    assign outputs[2265] = ~((layer0_outputs[6152]) ^ (layer0_outputs[9468]));
    assign outputs[2266] = layer0_outputs[6489];
    assign outputs[2267] = ~(layer0_outputs[6012]);
    assign outputs[2268] = ~((layer0_outputs[9622]) | (layer0_outputs[6954]));
    assign outputs[2269] = ~(layer0_outputs[8894]);
    assign outputs[2270] = layer0_outputs[8768];
    assign outputs[2271] = (layer0_outputs[1039]) | (layer0_outputs[9759]);
    assign outputs[2272] = ~(layer0_outputs[2339]);
    assign outputs[2273] = ~((layer0_outputs[6624]) ^ (layer0_outputs[731]));
    assign outputs[2274] = ~(layer0_outputs[8660]) | (layer0_outputs[7757]);
    assign outputs[2275] = ~(layer0_outputs[1363]);
    assign outputs[2276] = layer0_outputs[8843];
    assign outputs[2277] = (layer0_outputs[10164]) ^ (layer0_outputs[472]);
    assign outputs[2278] = (layer0_outputs[4082]) | (layer0_outputs[7270]);
    assign outputs[2279] = ~(layer0_outputs[7899]);
    assign outputs[2280] = ~(layer0_outputs[564]);
    assign outputs[2281] = (layer0_outputs[7773]) ^ (layer0_outputs[1371]);
    assign outputs[2282] = ~(layer0_outputs[1344]);
    assign outputs[2283] = ~(layer0_outputs[75]) | (layer0_outputs[6748]);
    assign outputs[2284] = ~((layer0_outputs[8602]) ^ (layer0_outputs[5612]));
    assign outputs[2285] = (layer0_outputs[4107]) ^ (layer0_outputs[4493]);
    assign outputs[2286] = layer0_outputs[3688];
    assign outputs[2287] = ~((layer0_outputs[8579]) & (layer0_outputs[1916]));
    assign outputs[2288] = ~(layer0_outputs[6560]);
    assign outputs[2289] = (layer0_outputs[7745]) & (layer0_outputs[1861]);
    assign outputs[2290] = layer0_outputs[3175];
    assign outputs[2291] = ~(layer0_outputs[6452]) | (layer0_outputs[1976]);
    assign outputs[2292] = layer0_outputs[5128];
    assign outputs[2293] = (layer0_outputs[6040]) ^ (layer0_outputs[1069]);
    assign outputs[2294] = layer0_outputs[3207];
    assign outputs[2295] = ~(layer0_outputs[3286]);
    assign outputs[2296] = ~(layer0_outputs[7342]) | (layer0_outputs[6848]);
    assign outputs[2297] = (layer0_outputs[6414]) & ~(layer0_outputs[2703]);
    assign outputs[2298] = layer0_outputs[8145];
    assign outputs[2299] = ~((layer0_outputs[9381]) | (layer0_outputs[10224]));
    assign outputs[2300] = layer0_outputs[2787];
    assign outputs[2301] = layer0_outputs[2956];
    assign outputs[2302] = layer0_outputs[9415];
    assign outputs[2303] = ~((layer0_outputs[217]) & (layer0_outputs[8321]));
    assign outputs[2304] = (layer0_outputs[1905]) ^ (layer0_outputs[3443]);
    assign outputs[2305] = ~(layer0_outputs[4004]);
    assign outputs[2306] = ~(layer0_outputs[3955]);
    assign outputs[2307] = layer0_outputs[4714];
    assign outputs[2308] = (layer0_outputs[8272]) ^ (layer0_outputs[2089]);
    assign outputs[2309] = ~((layer0_outputs[5281]) ^ (layer0_outputs[10187]));
    assign outputs[2310] = layer0_outputs[8189];
    assign outputs[2311] = (layer0_outputs[1848]) & ~(layer0_outputs[8364]);
    assign outputs[2312] = ~(layer0_outputs[3622]) | (layer0_outputs[2690]);
    assign outputs[2313] = (layer0_outputs[379]) & (layer0_outputs[3717]);
    assign outputs[2314] = ~(layer0_outputs[8502]);
    assign outputs[2315] = layer0_outputs[8808];
    assign outputs[2316] = (layer0_outputs[3335]) & (layer0_outputs[9324]);
    assign outputs[2317] = layer0_outputs[7488];
    assign outputs[2318] = layer0_outputs[8474];
    assign outputs[2319] = layer0_outputs[4254];
    assign outputs[2320] = ~((layer0_outputs[9216]) ^ (layer0_outputs[4463]));
    assign outputs[2321] = (layer0_outputs[1244]) ^ (layer0_outputs[9653]);
    assign outputs[2322] = ~(layer0_outputs[7975]);
    assign outputs[2323] = ~(layer0_outputs[9864]) | (layer0_outputs[3645]);
    assign outputs[2324] = ~(layer0_outputs[658]);
    assign outputs[2325] = ~(layer0_outputs[1266]);
    assign outputs[2326] = (layer0_outputs[6544]) ^ (layer0_outputs[8903]);
    assign outputs[2327] = ~(layer0_outputs[3803]);
    assign outputs[2328] = ~(layer0_outputs[8497]);
    assign outputs[2329] = layer0_outputs[6696];
    assign outputs[2330] = layer0_outputs[376];
    assign outputs[2331] = layer0_outputs[1419];
    assign outputs[2332] = ~((layer0_outputs[1489]) ^ (layer0_outputs[5387]));
    assign outputs[2333] = ~((layer0_outputs[5886]) ^ (layer0_outputs[6568]));
    assign outputs[2334] = ~(layer0_outputs[3212]) | (layer0_outputs[4880]);
    assign outputs[2335] = (layer0_outputs[7264]) ^ (layer0_outputs[8338]);
    assign outputs[2336] = layer0_outputs[1106];
    assign outputs[2337] = layer0_outputs[2918];
    assign outputs[2338] = (layer0_outputs[8025]) ^ (layer0_outputs[3641]);
    assign outputs[2339] = ~((layer0_outputs[7879]) | (layer0_outputs[8514]));
    assign outputs[2340] = layer0_outputs[9530];
    assign outputs[2341] = ~(layer0_outputs[5574]);
    assign outputs[2342] = (layer0_outputs[3883]) ^ (layer0_outputs[9096]);
    assign outputs[2343] = layer0_outputs[3213];
    assign outputs[2344] = layer0_outputs[5753];
    assign outputs[2345] = ~((layer0_outputs[2796]) | (layer0_outputs[9768]));
    assign outputs[2346] = layer0_outputs[7442];
    assign outputs[2347] = layer0_outputs[3563];
    assign outputs[2348] = ~((layer0_outputs[6925]) ^ (layer0_outputs[6340]));
    assign outputs[2349] = layer0_outputs[5790];
    assign outputs[2350] = ~(layer0_outputs[3762]);
    assign outputs[2351] = ~((layer0_outputs[15]) | (layer0_outputs[5971]));
    assign outputs[2352] = ~(layer0_outputs[1726]);
    assign outputs[2353] = layer0_outputs[7304];
    assign outputs[2354] = ~((layer0_outputs[6535]) & (layer0_outputs[1583]));
    assign outputs[2355] = ~(layer0_outputs[2285]);
    assign outputs[2356] = layer0_outputs[1505];
    assign outputs[2357] = (layer0_outputs[5625]) & (layer0_outputs[8138]);
    assign outputs[2358] = ~(layer0_outputs[7014]);
    assign outputs[2359] = (layer0_outputs[349]) ^ (layer0_outputs[7055]);
    assign outputs[2360] = ~(layer0_outputs[9879]);
    assign outputs[2361] = layer0_outputs[4126];
    assign outputs[2362] = ~(layer0_outputs[7905]);
    assign outputs[2363] = layer0_outputs[10237];
    assign outputs[2364] = layer0_outputs[2232];
    assign outputs[2365] = (layer0_outputs[8734]) & ~(layer0_outputs[5808]);
    assign outputs[2366] = ~((layer0_outputs[2212]) ^ (layer0_outputs[2656]));
    assign outputs[2367] = ~(layer0_outputs[6407]) | (layer0_outputs[1958]);
    assign outputs[2368] = layer0_outputs[9754];
    assign outputs[2369] = layer0_outputs[3577];
    assign outputs[2370] = ~(layer0_outputs[8553]);
    assign outputs[2371] = ~(layer0_outputs[6699]) | (layer0_outputs[76]);
    assign outputs[2372] = layer0_outputs[4204];
    assign outputs[2373] = layer0_outputs[2200];
    assign outputs[2374] = layer0_outputs[2761];
    assign outputs[2375] = ~(layer0_outputs[1610]) | (layer0_outputs[3565]);
    assign outputs[2376] = ~((layer0_outputs[2868]) | (layer0_outputs[7574]));
    assign outputs[2377] = ~((layer0_outputs[5167]) & (layer0_outputs[835]));
    assign outputs[2378] = ~((layer0_outputs[8948]) | (layer0_outputs[9624]));
    assign outputs[2379] = ~((layer0_outputs[569]) ^ (layer0_outputs[8563]));
    assign outputs[2380] = ~(layer0_outputs[5432]);
    assign outputs[2381] = ~(layer0_outputs[543]);
    assign outputs[2382] = ~(layer0_outputs[4364]) | (layer0_outputs[2117]);
    assign outputs[2383] = ~(layer0_outputs[7946]) | (layer0_outputs[994]);
    assign outputs[2384] = layer0_outputs[5813];
    assign outputs[2385] = layer0_outputs[2543];
    assign outputs[2386] = layer0_outputs[6565];
    assign outputs[2387] = ~((layer0_outputs[2395]) ^ (layer0_outputs[2035]));
    assign outputs[2388] = (layer0_outputs[5240]) | (layer0_outputs[8024]);
    assign outputs[2389] = layer0_outputs[1179];
    assign outputs[2390] = ~(layer0_outputs[2325]) | (layer0_outputs[5627]);
    assign outputs[2391] = layer0_outputs[3506];
    assign outputs[2392] = ~(layer0_outputs[6782]);
    assign outputs[2393] = ~((layer0_outputs[8992]) ^ (layer0_outputs[6937]));
    assign outputs[2394] = ~(layer0_outputs[9955]) | (layer0_outputs[5441]);
    assign outputs[2395] = ~(layer0_outputs[116]);
    assign outputs[2396] = ~(layer0_outputs[2476]);
    assign outputs[2397] = ~(layer0_outputs[257]);
    assign outputs[2398] = ~(layer0_outputs[8948]);
    assign outputs[2399] = ~((layer0_outputs[6652]) ^ (layer0_outputs[4080]));
    assign outputs[2400] = layer0_outputs[2915];
    assign outputs[2401] = (layer0_outputs[526]) ^ (layer0_outputs[612]);
    assign outputs[2402] = layer0_outputs[6794];
    assign outputs[2403] = ~((layer0_outputs[4208]) ^ (layer0_outputs[7706]));
    assign outputs[2404] = (layer0_outputs[8493]) ^ (layer0_outputs[6476]);
    assign outputs[2405] = ~(layer0_outputs[5608]);
    assign outputs[2406] = ~(layer0_outputs[9120]);
    assign outputs[2407] = ~(layer0_outputs[3820]);
    assign outputs[2408] = layer0_outputs[7580];
    assign outputs[2409] = (layer0_outputs[7551]) ^ (layer0_outputs[3326]);
    assign outputs[2410] = ~(layer0_outputs[4455]);
    assign outputs[2411] = ~(layer0_outputs[10014]);
    assign outputs[2412] = ~(layer0_outputs[5829]);
    assign outputs[2413] = (layer0_outputs[5145]) | (layer0_outputs[5134]);
    assign outputs[2414] = ~(layer0_outputs[7586]);
    assign outputs[2415] = layer0_outputs[9482];
    assign outputs[2416] = ~(layer0_outputs[335]);
    assign outputs[2417] = ~(layer0_outputs[93]);
    assign outputs[2418] = ~(layer0_outputs[415]);
    assign outputs[2419] = (layer0_outputs[6349]) ^ (layer0_outputs[6604]);
    assign outputs[2420] = (layer0_outputs[10176]) ^ (layer0_outputs[6259]);
    assign outputs[2421] = layer0_outputs[6356];
    assign outputs[2422] = ~(layer0_outputs[1813]);
    assign outputs[2423] = (layer0_outputs[2484]) & ~(layer0_outputs[7812]);
    assign outputs[2424] = layer0_outputs[3855];
    assign outputs[2425] = ~(layer0_outputs[8962]);
    assign outputs[2426] = layer0_outputs[930];
    assign outputs[2427] = ~(layer0_outputs[1877]);
    assign outputs[2428] = ~(layer0_outputs[5549]);
    assign outputs[2429] = layer0_outputs[9970];
    assign outputs[2430] = layer0_outputs[6389];
    assign outputs[2431] = ~((layer0_outputs[2672]) | (layer0_outputs[8934]));
    assign outputs[2432] = layer0_outputs[6892];
    assign outputs[2433] = ~((layer0_outputs[367]) ^ (layer0_outputs[2854]));
    assign outputs[2434] = (layer0_outputs[5573]) | (layer0_outputs[4784]);
    assign outputs[2435] = (layer0_outputs[3385]) & ~(layer0_outputs[7522]);
    assign outputs[2436] = layer0_outputs[5186];
    assign outputs[2437] = layer0_outputs[1638];
    assign outputs[2438] = ~(layer0_outputs[6664]);
    assign outputs[2439] = ~((layer0_outputs[5494]) ^ (layer0_outputs[4090]));
    assign outputs[2440] = ~((layer0_outputs[8267]) ^ (layer0_outputs[1182]));
    assign outputs[2441] = layer0_outputs[2335];
    assign outputs[2442] = ~(layer0_outputs[8242]);
    assign outputs[2443] = ~(layer0_outputs[4681]);
    assign outputs[2444] = (layer0_outputs[6281]) ^ (layer0_outputs[6874]);
    assign outputs[2445] = ~((layer0_outputs[16]) ^ (layer0_outputs[5043]));
    assign outputs[2446] = (layer0_outputs[2748]) & (layer0_outputs[2106]);
    assign outputs[2447] = ~(layer0_outputs[6108]);
    assign outputs[2448] = layer0_outputs[2323];
    assign outputs[2449] = layer0_outputs[4943];
    assign outputs[2450] = layer0_outputs[7973];
    assign outputs[2451] = (layer0_outputs[8839]) & ~(layer0_outputs[6277]);
    assign outputs[2452] = (layer0_outputs[3081]) | (layer0_outputs[2812]);
    assign outputs[2453] = layer0_outputs[9509];
    assign outputs[2454] = ~(layer0_outputs[227]) | (layer0_outputs[159]);
    assign outputs[2455] = ~((layer0_outputs[3211]) ^ (layer0_outputs[4787]));
    assign outputs[2456] = layer0_outputs[5351];
    assign outputs[2457] = ~(layer0_outputs[4877]);
    assign outputs[2458] = layer0_outputs[1863];
    assign outputs[2459] = layer0_outputs[499];
    assign outputs[2460] = ~(layer0_outputs[1700]) | (layer0_outputs[3586]);
    assign outputs[2461] = layer0_outputs[961];
    assign outputs[2462] = layer0_outputs[3260];
    assign outputs[2463] = ~(layer0_outputs[3803]) | (layer0_outputs[9132]);
    assign outputs[2464] = ~((layer0_outputs[4]) ^ (layer0_outputs[4676]));
    assign outputs[2465] = (layer0_outputs[383]) ^ (layer0_outputs[9310]);
    assign outputs[2466] = ~((layer0_outputs[9961]) & (layer0_outputs[2498]));
    assign outputs[2467] = layer0_outputs[566];
    assign outputs[2468] = layer0_outputs[9731];
    assign outputs[2469] = (layer0_outputs[2785]) & ~(layer0_outputs[5144]);
    assign outputs[2470] = ~(layer0_outputs[5307]);
    assign outputs[2471] = layer0_outputs[8376];
    assign outputs[2472] = ~(layer0_outputs[7985]);
    assign outputs[2473] = ~(layer0_outputs[9781]) | (layer0_outputs[8636]);
    assign outputs[2474] = layer0_outputs[7135];
    assign outputs[2475] = (layer0_outputs[4604]) & ~(layer0_outputs[3230]);
    assign outputs[2476] = (layer0_outputs[3205]) ^ (layer0_outputs[4539]);
    assign outputs[2477] = ~(layer0_outputs[7971]) | (layer0_outputs[3656]);
    assign outputs[2478] = layer0_outputs[6876];
    assign outputs[2479] = ~(layer0_outputs[1251]) | (layer0_outputs[5373]);
    assign outputs[2480] = ~((layer0_outputs[6090]) & (layer0_outputs[8028]));
    assign outputs[2481] = ~(layer0_outputs[147]);
    assign outputs[2482] = (layer0_outputs[301]) | (layer0_outputs[6677]);
    assign outputs[2483] = ~(layer0_outputs[4903]);
    assign outputs[2484] = layer0_outputs[4417];
    assign outputs[2485] = ~(layer0_outputs[4141]);
    assign outputs[2486] = (layer0_outputs[3214]) ^ (layer0_outputs[9136]);
    assign outputs[2487] = layer0_outputs[1371];
    assign outputs[2488] = (layer0_outputs[3114]) ^ (layer0_outputs[890]);
    assign outputs[2489] = layer0_outputs[7230];
    assign outputs[2490] = ~(layer0_outputs[6438]);
    assign outputs[2491] = ~(layer0_outputs[1114]);
    assign outputs[2492] = ~(layer0_outputs[5512]);
    assign outputs[2493] = ~((layer0_outputs[6685]) & (layer0_outputs[2599]));
    assign outputs[2494] = ~(layer0_outputs[4181]);
    assign outputs[2495] = layer0_outputs[128];
    assign outputs[2496] = (layer0_outputs[9253]) & ~(layer0_outputs[5109]);
    assign outputs[2497] = ~((layer0_outputs[2073]) ^ (layer0_outputs[284]));
    assign outputs[2498] = (layer0_outputs[5231]) | (layer0_outputs[4428]);
    assign outputs[2499] = (layer0_outputs[818]) ^ (layer0_outputs[2567]);
    assign outputs[2500] = layer0_outputs[5720];
    assign outputs[2501] = (layer0_outputs[8941]) & ~(layer0_outputs[4457]);
    assign outputs[2502] = ~(layer0_outputs[3201]);
    assign outputs[2503] = ~(layer0_outputs[7329]);
    assign outputs[2504] = ~(layer0_outputs[1871]);
    assign outputs[2505] = ~(layer0_outputs[6798]);
    assign outputs[2506] = (layer0_outputs[9772]) | (layer0_outputs[4953]);
    assign outputs[2507] = ~(layer0_outputs[5108]) | (layer0_outputs[6180]);
    assign outputs[2508] = ~((layer0_outputs[7495]) ^ (layer0_outputs[5088]));
    assign outputs[2509] = (layer0_outputs[2049]) ^ (layer0_outputs[2978]);
    assign outputs[2510] = layer0_outputs[441];
    assign outputs[2511] = (layer0_outputs[9380]) & (layer0_outputs[9372]);
    assign outputs[2512] = layer0_outputs[5624];
    assign outputs[2513] = ~(layer0_outputs[4871]);
    assign outputs[2514] = ~(layer0_outputs[2476]);
    assign outputs[2515] = ~((layer0_outputs[6067]) ^ (layer0_outputs[8627]));
    assign outputs[2516] = ~(layer0_outputs[2148]) | (layer0_outputs[6773]);
    assign outputs[2517] = layer0_outputs[6048];
    assign outputs[2518] = layer0_outputs[5870];
    assign outputs[2519] = layer0_outputs[10028];
    assign outputs[2520] = (layer0_outputs[7010]) ^ (layer0_outputs[6632]);
    assign outputs[2521] = (layer0_outputs[2025]) ^ (layer0_outputs[6746]);
    assign outputs[2522] = layer0_outputs[2789];
    assign outputs[2523] = layer0_outputs[1418];
    assign outputs[2524] = ~(layer0_outputs[4022]);
    assign outputs[2525] = ~(layer0_outputs[366]);
    assign outputs[2526] = ~((layer0_outputs[6755]) ^ (layer0_outputs[1258]));
    assign outputs[2527] = ~(layer0_outputs[4077]) | (layer0_outputs[6996]);
    assign outputs[2528] = ~(layer0_outputs[250]);
    assign outputs[2529] = ~(layer0_outputs[7636]);
    assign outputs[2530] = layer0_outputs[5993];
    assign outputs[2531] = (layer0_outputs[152]) ^ (layer0_outputs[1335]);
    assign outputs[2532] = ~(layer0_outputs[5445]);
    assign outputs[2533] = (layer0_outputs[7217]) & ~(layer0_outputs[6772]);
    assign outputs[2534] = layer0_outputs[2010];
    assign outputs[2535] = ~((layer0_outputs[4024]) ^ (layer0_outputs[6839]));
    assign outputs[2536] = layer0_outputs[4291];
    assign outputs[2537] = ~(layer0_outputs[5791]);
    assign outputs[2538] = (layer0_outputs[1434]) ^ (layer0_outputs[3631]);
    assign outputs[2539] = ~((layer0_outputs[1547]) & (layer0_outputs[7543]));
    assign outputs[2540] = ~(layer0_outputs[4077]);
    assign outputs[2541] = ~(layer0_outputs[3789]);
    assign outputs[2542] = (layer0_outputs[9350]) & (layer0_outputs[7612]);
    assign outputs[2543] = (layer0_outputs[66]) | (layer0_outputs[3939]);
    assign outputs[2544] = (layer0_outputs[628]) | (layer0_outputs[9069]);
    assign outputs[2545] = (layer0_outputs[4996]) ^ (layer0_outputs[369]);
    assign outputs[2546] = ~((layer0_outputs[46]) & (layer0_outputs[6426]));
    assign outputs[2547] = ~((layer0_outputs[5859]) | (layer0_outputs[7976]));
    assign outputs[2548] = ~((layer0_outputs[5755]) | (layer0_outputs[9741]));
    assign outputs[2549] = ~(layer0_outputs[2775]);
    assign outputs[2550] = layer0_outputs[4339];
    assign outputs[2551] = layer0_outputs[8878];
    assign outputs[2552] = (layer0_outputs[9532]) ^ (layer0_outputs[3356]);
    assign outputs[2553] = (layer0_outputs[5238]) & ~(layer0_outputs[2194]);
    assign outputs[2554] = layer0_outputs[1838];
    assign outputs[2555] = (layer0_outputs[2181]) ^ (layer0_outputs[9201]);
    assign outputs[2556] = ~(layer0_outputs[4862]);
    assign outputs[2557] = ~(layer0_outputs[4978]);
    assign outputs[2558] = ~(layer0_outputs[6448]);
    assign outputs[2559] = (layer0_outputs[5023]) | (layer0_outputs[4480]);
    assign outputs[2560] = ~(layer0_outputs[8143]);
    assign outputs[2561] = ~((layer0_outputs[2920]) | (layer0_outputs[5598]));
    assign outputs[2562] = layer0_outputs[5064];
    assign outputs[2563] = ~(layer0_outputs[5306]);
    assign outputs[2564] = ~(layer0_outputs[6764]);
    assign outputs[2565] = ~(layer0_outputs[6099]);
    assign outputs[2566] = ~(layer0_outputs[1200]);
    assign outputs[2567] = ~(layer0_outputs[8741]) | (layer0_outputs[1606]);
    assign outputs[2568] = (layer0_outputs[9481]) & (layer0_outputs[6607]);
    assign outputs[2569] = (layer0_outputs[2749]) & ~(layer0_outputs[8146]);
    assign outputs[2570] = ~(layer0_outputs[8104]);
    assign outputs[2571] = ~((layer0_outputs[339]) ^ (layer0_outputs[9368]));
    assign outputs[2572] = layer0_outputs[9569];
    assign outputs[2573] = layer0_outputs[212];
    assign outputs[2574] = layer0_outputs[7296];
    assign outputs[2575] = layer0_outputs[501];
    assign outputs[2576] = layer0_outputs[8037];
    assign outputs[2577] = ~(layer0_outputs[9197]);
    assign outputs[2578] = ~(layer0_outputs[4210]);
    assign outputs[2579] = (layer0_outputs[3069]) & (layer0_outputs[4627]);
    assign outputs[2580] = ~(layer0_outputs[2446]);
    assign outputs[2581] = layer0_outputs[5510];
    assign outputs[2582] = layer0_outputs[1790];
    assign outputs[2583] = ~((layer0_outputs[512]) & (layer0_outputs[560]));
    assign outputs[2584] = ~(layer0_outputs[6544]) | (layer0_outputs[4477]);
    assign outputs[2585] = ~((layer0_outputs[6661]) & (layer0_outputs[4634]));
    assign outputs[2586] = ~(layer0_outputs[6971]);
    assign outputs[2587] = (layer0_outputs[7793]) | (layer0_outputs[2982]);
    assign outputs[2588] = ~(layer0_outputs[7868]);
    assign outputs[2589] = layer0_outputs[9433];
    assign outputs[2590] = layer0_outputs[9215];
    assign outputs[2591] = ~(layer0_outputs[5089]);
    assign outputs[2592] = ~((layer0_outputs[2291]) ^ (layer0_outputs[1714]));
    assign outputs[2593] = layer0_outputs[8335];
    assign outputs[2594] = (layer0_outputs[3348]) ^ (layer0_outputs[4479]);
    assign outputs[2595] = ~(layer0_outputs[9722]) | (layer0_outputs[3405]);
    assign outputs[2596] = ~((layer0_outputs[2601]) ^ (layer0_outputs[5264]));
    assign outputs[2597] = ~((layer0_outputs[8089]) | (layer0_outputs[1023]));
    assign outputs[2598] = (layer0_outputs[5332]) & ~(layer0_outputs[7954]);
    assign outputs[2599] = ~(layer0_outputs[5734]);
    assign outputs[2600] = (layer0_outputs[2239]) & (layer0_outputs[7096]);
    assign outputs[2601] = ~(layer0_outputs[3526]);
    assign outputs[2602] = (layer0_outputs[5588]) | (layer0_outputs[3087]);
    assign outputs[2603] = ~(layer0_outputs[10038]);
    assign outputs[2604] = ~(layer0_outputs[9571]);
    assign outputs[2605] = layer0_outputs[1364];
    assign outputs[2606] = layer0_outputs[5708];
    assign outputs[2607] = (layer0_outputs[3763]) | (layer0_outputs[3976]);
    assign outputs[2608] = layer0_outputs[9966];
    assign outputs[2609] = (layer0_outputs[2519]) & ~(layer0_outputs[4744]);
    assign outputs[2610] = ~(layer0_outputs[5322]) | (layer0_outputs[8698]);
    assign outputs[2611] = ~(layer0_outputs[3748]);
    assign outputs[2612] = ~((layer0_outputs[4118]) ^ (layer0_outputs[3897]));
    assign outputs[2613] = (layer0_outputs[156]) & (layer0_outputs[9048]);
    assign outputs[2614] = layer0_outputs[1938];
    assign outputs[2615] = ~(layer0_outputs[1591]) | (layer0_outputs[6997]);
    assign outputs[2616] = ~(layer0_outputs[1053]);
    assign outputs[2617] = ~((layer0_outputs[9581]) ^ (layer0_outputs[3050]));
    assign outputs[2618] = ~(layer0_outputs[277]) | (layer0_outputs[5577]);
    assign outputs[2619] = layer0_outputs[8179];
    assign outputs[2620] = ~(layer0_outputs[103]);
    assign outputs[2621] = ~(layer0_outputs[1870]);
    assign outputs[2622] = layer0_outputs[236];
    assign outputs[2623] = ~(layer0_outputs[3202]) | (layer0_outputs[616]);
    assign outputs[2624] = layer0_outputs[6136];
    assign outputs[2625] = (layer0_outputs[4812]) ^ (layer0_outputs[6270]);
    assign outputs[2626] = ~(layer0_outputs[2638]);
    assign outputs[2627] = ~(layer0_outputs[5571]);
    assign outputs[2628] = layer0_outputs[2528];
    assign outputs[2629] = ~(layer0_outputs[9630]) | (layer0_outputs[8311]);
    assign outputs[2630] = (layer0_outputs[5690]) | (layer0_outputs[4950]);
    assign outputs[2631] = layer0_outputs[9328];
    assign outputs[2632] = ~(layer0_outputs[9912]);
    assign outputs[2633] = ~((layer0_outputs[3582]) ^ (layer0_outputs[6808]));
    assign outputs[2634] = ~((layer0_outputs[1095]) ^ (layer0_outputs[1187]));
    assign outputs[2635] = ~((layer0_outputs[8755]) & (layer0_outputs[8866]));
    assign outputs[2636] = (layer0_outputs[6363]) ^ (layer0_outputs[2017]);
    assign outputs[2637] = ~((layer0_outputs[6761]) ^ (layer0_outputs[8050]));
    assign outputs[2638] = layer0_outputs[7377];
    assign outputs[2639] = ~((layer0_outputs[829]) ^ (layer0_outputs[9466]));
    assign outputs[2640] = ~((layer0_outputs[2009]) | (layer0_outputs[2663]));
    assign outputs[2641] = layer0_outputs[7347];
    assign outputs[2642] = (layer0_outputs[2539]) ^ (layer0_outputs[286]);
    assign outputs[2643] = (layer0_outputs[3511]) | (layer0_outputs[5125]);
    assign outputs[2644] = ~((layer0_outputs[3060]) ^ (layer0_outputs[5930]));
    assign outputs[2645] = ~((layer0_outputs[9506]) & (layer0_outputs[5526]));
    assign outputs[2646] = ~((layer0_outputs[2090]) ^ (layer0_outputs[9747]));
    assign outputs[2647] = (layer0_outputs[3698]) | (layer0_outputs[5320]);
    assign outputs[2648] = layer0_outputs[5887];
    assign outputs[2649] = ~(layer0_outputs[189]);
    assign outputs[2650] = ~((layer0_outputs[6158]) ^ (layer0_outputs[1365]));
    assign outputs[2651] = ~((layer0_outputs[3082]) ^ (layer0_outputs[8205]));
    assign outputs[2652] = (layer0_outputs[478]) ^ (layer0_outputs[442]);
    assign outputs[2653] = ~(layer0_outputs[8544]);
    assign outputs[2654] = layer0_outputs[3686];
    assign outputs[2655] = ~(layer0_outputs[8976]);
    assign outputs[2656] = layer0_outputs[6814];
    assign outputs[2657] = ~(layer0_outputs[6354]) | (layer0_outputs[1976]);
    assign outputs[2658] = ~((layer0_outputs[6322]) ^ (layer0_outputs[8510]));
    assign outputs[2659] = ~((layer0_outputs[4601]) & (layer0_outputs[1983]));
    assign outputs[2660] = ~(layer0_outputs[1881]);
    assign outputs[2661] = ~(layer0_outputs[3395]);
    assign outputs[2662] = ~(layer0_outputs[1679]);
    assign outputs[2663] = ~(layer0_outputs[6254]);
    assign outputs[2664] = ~(layer0_outputs[3644]);
    assign outputs[2665] = ~(layer0_outputs[8523]);
    assign outputs[2666] = layer0_outputs[8263];
    assign outputs[2667] = ~(layer0_outputs[9510]);
    assign outputs[2668] = ~((layer0_outputs[4760]) | (layer0_outputs[5826]));
    assign outputs[2669] = (layer0_outputs[583]) & ~(layer0_outputs[7555]);
    assign outputs[2670] = layer0_outputs[6317];
    assign outputs[2671] = (layer0_outputs[2994]) & ~(layer0_outputs[6809]);
    assign outputs[2672] = (layer0_outputs[736]) ^ (layer0_outputs[4075]);
    assign outputs[2673] = ~(layer0_outputs[549]);
    assign outputs[2674] = ~(layer0_outputs[7904]);
    assign outputs[2675] = layer0_outputs[8587];
    assign outputs[2676] = layer0_outputs[3615];
    assign outputs[2677] = (layer0_outputs[8697]) & ~(layer0_outputs[2394]);
    assign outputs[2678] = layer0_outputs[5862];
    assign outputs[2679] = ~(layer0_outputs[800]) | (layer0_outputs[9067]);
    assign outputs[2680] = ~(layer0_outputs[2442]);
    assign outputs[2681] = ~(layer0_outputs[4869]);
    assign outputs[2682] = ~(layer0_outputs[6220]) | (layer0_outputs[2700]);
    assign outputs[2683] = ~(layer0_outputs[5179]);
    assign outputs[2684] = layer0_outputs[5945];
    assign outputs[2685] = (layer0_outputs[5890]) ^ (layer0_outputs[6148]);
    assign outputs[2686] = layer0_outputs[1632];
    assign outputs[2687] = layer0_outputs[2197];
    assign outputs[2688] = ~(layer0_outputs[1832]) | (layer0_outputs[1507]);
    assign outputs[2689] = ~(layer0_outputs[9767]);
    assign outputs[2690] = ~(layer0_outputs[6547]);
    assign outputs[2691] = ~((layer0_outputs[1622]) ^ (layer0_outputs[1055]));
    assign outputs[2692] = ~(layer0_outputs[2524]);
    assign outputs[2693] = layer0_outputs[1130];
    assign outputs[2694] = layer0_outputs[757];
    assign outputs[2695] = layer0_outputs[4599];
    assign outputs[2696] = layer0_outputs[65];
    assign outputs[2697] = layer0_outputs[8290];
    assign outputs[2698] = layer0_outputs[2899];
    assign outputs[2699] = ~(layer0_outputs[4340]) | (layer0_outputs[5682]);
    assign outputs[2700] = ~(layer0_outputs[5236]);
    assign outputs[2701] = layer0_outputs[6630];
    assign outputs[2702] = layer0_outputs[780];
    assign outputs[2703] = ~(layer0_outputs[1924]);
    assign outputs[2704] = ~((layer0_outputs[8909]) & (layer0_outputs[2125]));
    assign outputs[2705] = (layer0_outputs[3327]) & ~(layer0_outputs[4924]);
    assign outputs[2706] = ~((layer0_outputs[389]) & (layer0_outputs[8586]));
    assign outputs[2707] = ~(layer0_outputs[9905]);
    assign outputs[2708] = (layer0_outputs[4952]) | (layer0_outputs[1221]);
    assign outputs[2709] = (layer0_outputs[7728]) & (layer0_outputs[7664]);
    assign outputs[2710] = layer0_outputs[72];
    assign outputs[2711] = (layer0_outputs[6151]) ^ (layer0_outputs[7426]);
    assign outputs[2712] = layer0_outputs[3011];
    assign outputs[2713] = ~((layer0_outputs[48]) & (layer0_outputs[3937]));
    assign outputs[2714] = layer0_outputs[5858];
    assign outputs[2715] = ~(layer0_outputs[4514]);
    assign outputs[2716] = (layer0_outputs[2739]) ^ (layer0_outputs[5851]);
    assign outputs[2717] = ~((layer0_outputs[1612]) ^ (layer0_outputs[1670]));
    assign outputs[2718] = (layer0_outputs[3860]) & ~(layer0_outputs[801]);
    assign outputs[2719] = layer0_outputs[0];
    assign outputs[2720] = ~((layer0_outputs[3046]) & (layer0_outputs[6991]));
    assign outputs[2721] = (layer0_outputs[10016]) ^ (layer0_outputs[9046]);
    assign outputs[2722] = (layer0_outputs[8228]) | (layer0_outputs[8198]);
    assign outputs[2723] = ~((layer0_outputs[8153]) | (layer0_outputs[1036]));
    assign outputs[2724] = (layer0_outputs[4716]) | (layer0_outputs[1305]);
    assign outputs[2725] = (layer0_outputs[1680]) & ~(layer0_outputs[970]);
    assign outputs[2726] = ~((layer0_outputs[2306]) & (layer0_outputs[2392]));
    assign outputs[2727] = layer0_outputs[273];
    assign outputs[2728] = ~(layer0_outputs[677]);
    assign outputs[2729] = ~(layer0_outputs[1252]) | (layer0_outputs[3293]);
    assign outputs[2730] = (layer0_outputs[5026]) ^ (layer0_outputs[8670]);
    assign outputs[2731] = layer0_outputs[2990];
    assign outputs[2732] = (layer0_outputs[798]) & ~(layer0_outputs[5797]);
    assign outputs[2733] = layer0_outputs[8412];
    assign outputs[2734] = ~(layer0_outputs[7815]);
    assign outputs[2735] = layer0_outputs[2905];
    assign outputs[2736] = ~(layer0_outputs[9883]);
    assign outputs[2737] = ~((layer0_outputs[2007]) ^ (layer0_outputs[4458]));
    assign outputs[2738] = ~((layer0_outputs[242]) ^ (layer0_outputs[922]));
    assign outputs[2739] = layer0_outputs[1220];
    assign outputs[2740] = ~((layer0_outputs[1538]) | (layer0_outputs[8536]));
    assign outputs[2741] = ~((layer0_outputs[9876]) & (layer0_outputs[9850]));
    assign outputs[2742] = (layer0_outputs[828]) ^ (layer0_outputs[992]);
    assign outputs[2743] = ~(layer0_outputs[2960]);
    assign outputs[2744] = layer0_outputs[1897];
    assign outputs[2745] = ~(layer0_outputs[1427]) | (layer0_outputs[3377]);
    assign outputs[2746] = ~((layer0_outputs[10116]) ^ (layer0_outputs[5557]));
    assign outputs[2747] = layer0_outputs[5456];
    assign outputs[2748] = layer0_outputs[756];
    assign outputs[2749] = ~(layer0_outputs[5505]);
    assign outputs[2750] = (layer0_outputs[8537]) ^ (layer0_outputs[2053]);
    assign outputs[2751] = ~((layer0_outputs[7598]) ^ (layer0_outputs[7121]));
    assign outputs[2752] = layer0_outputs[4334];
    assign outputs[2753] = ~((layer0_outputs[2450]) ^ (layer0_outputs[6502]));
    assign outputs[2754] = layer0_outputs[6356];
    assign outputs[2755] = (layer0_outputs[4560]) & ~(layer0_outputs[3124]);
    assign outputs[2756] = layer0_outputs[7920];
    assign outputs[2757] = (layer0_outputs[1007]) ^ (layer0_outputs[9653]);
    assign outputs[2758] = layer0_outputs[31];
    assign outputs[2759] = ~(layer0_outputs[8307]);
    assign outputs[2760] = ~(layer0_outputs[1324]) | (layer0_outputs[641]);
    assign outputs[2761] = layer0_outputs[3588];
    assign outputs[2762] = ~((layer0_outputs[9496]) ^ (layer0_outputs[2692]));
    assign outputs[2763] = ~((layer0_outputs[6975]) & (layer0_outputs[8184]));
    assign outputs[2764] = layer0_outputs[6079];
    assign outputs[2765] = ~(layer0_outputs[9395]);
    assign outputs[2766] = (layer0_outputs[10045]) & (layer0_outputs[4061]);
    assign outputs[2767] = ~(layer0_outputs[5956]);
    assign outputs[2768] = layer0_outputs[581];
    assign outputs[2769] = ~(layer0_outputs[2270]) | (layer0_outputs[8179]);
    assign outputs[2770] = ~(layer0_outputs[7671]) | (layer0_outputs[7440]);
    assign outputs[2771] = layer0_outputs[3088];
    assign outputs[2772] = layer0_outputs[10214];
    assign outputs[2773] = (layer0_outputs[5012]) ^ (layer0_outputs[825]);
    assign outputs[2774] = ~((layer0_outputs[10021]) | (layer0_outputs[3590]));
    assign outputs[2775] = ~(layer0_outputs[2906]);
    assign outputs[2776] = ~(layer0_outputs[9190]);
    assign outputs[2777] = ~(layer0_outputs[3852]);
    assign outputs[2778] = layer0_outputs[4249];
    assign outputs[2779] = layer0_outputs[9131];
    assign outputs[2780] = layer0_outputs[8895];
    assign outputs[2781] = layer0_outputs[7447];
    assign outputs[2782] = ~((layer0_outputs[10073]) | (layer0_outputs[9574]));
    assign outputs[2783] = layer0_outputs[9022];
    assign outputs[2784] = layer0_outputs[10006];
    assign outputs[2785] = (layer0_outputs[5917]) ^ (layer0_outputs[4447]);
    assign outputs[2786] = ~(layer0_outputs[1096]) | (layer0_outputs[9298]);
    assign outputs[2787] = layer0_outputs[7736];
    assign outputs[2788] = ~(layer0_outputs[8543]);
    assign outputs[2789] = layer0_outputs[2329];
    assign outputs[2790] = ~(layer0_outputs[3125]);
    assign outputs[2791] = ~(layer0_outputs[3303]);
    assign outputs[2792] = layer0_outputs[2370];
    assign outputs[2793] = layer0_outputs[6922];
    assign outputs[2794] = ~(layer0_outputs[8089]) | (layer0_outputs[10188]);
    assign outputs[2795] = ~(layer0_outputs[294]);
    assign outputs[2796] = ~(layer0_outputs[794]);
    assign outputs[2797] = layer0_outputs[29];
    assign outputs[2798] = ~((layer0_outputs[4421]) ^ (layer0_outputs[2977]));
    assign outputs[2799] = ~(layer0_outputs[4440]) | (layer0_outputs[8507]);
    assign outputs[2800] = layer0_outputs[1825];
    assign outputs[2801] = (layer0_outputs[9877]) & ~(layer0_outputs[4945]);
    assign outputs[2802] = ~((layer0_outputs[2340]) & (layer0_outputs[8261]));
    assign outputs[2803] = (layer0_outputs[8489]) & ~(layer0_outputs[4050]);
    assign outputs[2804] = ~(layer0_outputs[4205]) | (layer0_outputs[10021]);
    assign outputs[2805] = (layer0_outputs[6982]) & ~(layer0_outputs[8630]);
    assign outputs[2806] = layer0_outputs[7825];
    assign outputs[2807] = (layer0_outputs[4644]) ^ (layer0_outputs[8265]);
    assign outputs[2808] = ~(layer0_outputs[6659]);
    assign outputs[2809] = ~(layer0_outputs[7522]);
    assign outputs[2810] = layer0_outputs[1328];
    assign outputs[2811] = (layer0_outputs[6639]) & ~(layer0_outputs[5594]);
    assign outputs[2812] = ~(layer0_outputs[3595]);
    assign outputs[2813] = layer0_outputs[6414];
    assign outputs[2814] = layer0_outputs[3289];
    assign outputs[2815] = layer0_outputs[8455];
    assign outputs[2816] = (layer0_outputs[5885]) & ~(layer0_outputs[2245]);
    assign outputs[2817] = (layer0_outputs[3467]) | (layer0_outputs[5117]);
    assign outputs[2818] = ~(layer0_outputs[2270]) | (layer0_outputs[2242]);
    assign outputs[2819] = ~(layer0_outputs[6112]);
    assign outputs[2820] = (layer0_outputs[4114]) ^ (layer0_outputs[10174]);
    assign outputs[2821] = ~(layer0_outputs[7957]);
    assign outputs[2822] = ~(layer0_outputs[4275]);
    assign outputs[2823] = layer0_outputs[9970];
    assign outputs[2824] = layer0_outputs[1569];
    assign outputs[2825] = ~(layer0_outputs[10200]);
    assign outputs[2826] = (layer0_outputs[1177]) | (layer0_outputs[2111]);
    assign outputs[2827] = ~(layer0_outputs[7641]);
    assign outputs[2828] = ~(layer0_outputs[944]);
    assign outputs[2829] = ~((layer0_outputs[4485]) ^ (layer0_outputs[8930]));
    assign outputs[2830] = layer0_outputs[1502];
    assign outputs[2831] = layer0_outputs[49];
    assign outputs[2832] = ~(layer0_outputs[3848]);
    assign outputs[2833] = ~((layer0_outputs[1137]) ^ (layer0_outputs[3726]));
    assign outputs[2834] = (layer0_outputs[2434]) | (layer0_outputs[210]);
    assign outputs[2835] = ~(layer0_outputs[6407]) | (layer0_outputs[10151]);
    assign outputs[2836] = ~(layer0_outputs[3131]) | (layer0_outputs[7353]);
    assign outputs[2837] = ~((layer0_outputs[8190]) & (layer0_outputs[5489]));
    assign outputs[2838] = ~(layer0_outputs[4607]) | (layer0_outputs[5363]);
    assign outputs[2839] = (layer0_outputs[8282]) | (layer0_outputs[811]);
    assign outputs[2840] = ~(layer0_outputs[6541]) | (layer0_outputs[9334]);
    assign outputs[2841] = ~((layer0_outputs[3136]) ^ (layer0_outputs[230]));
    assign outputs[2842] = ~(layer0_outputs[3821]) | (layer0_outputs[6933]);
    assign outputs[2843] = layer0_outputs[5357];
    assign outputs[2844] = ~((layer0_outputs[5522]) ^ (layer0_outputs[1500]));
    assign outputs[2845] = layer0_outputs[2560];
    assign outputs[2846] = ~(layer0_outputs[5629]) | (layer0_outputs[1682]);
    assign outputs[2847] = ~(layer0_outputs[3884]);
    assign outputs[2848] = layer0_outputs[4332];
    assign outputs[2849] = layer0_outputs[8715];
    assign outputs[2850] = layer0_outputs[9597];
    assign outputs[2851] = ~(layer0_outputs[7744]) | (layer0_outputs[8592]);
    assign outputs[2852] = ~((layer0_outputs[9604]) ^ (layer0_outputs[3399]));
    assign outputs[2853] = layer0_outputs[0];
    assign outputs[2854] = ~(layer0_outputs[7723]) | (layer0_outputs[4232]);
    assign outputs[2855] = ~(layer0_outputs[6649]) | (layer0_outputs[2547]);
    assign outputs[2856] = ~(layer0_outputs[3296]);
    assign outputs[2857] = ~(layer0_outputs[541]);
    assign outputs[2858] = ~(layer0_outputs[9184]);
    assign outputs[2859] = ~(layer0_outputs[6863]);
    assign outputs[2860] = layer0_outputs[8504];
    assign outputs[2861] = ~((layer0_outputs[1675]) & (layer0_outputs[6563]));
    assign outputs[2862] = ~(layer0_outputs[5752]);
    assign outputs[2863] = ~(layer0_outputs[1535]);
    assign outputs[2864] = (layer0_outputs[5362]) ^ (layer0_outputs[8801]);
    assign outputs[2865] = (layer0_outputs[3529]) & ~(layer0_outputs[3078]);
    assign outputs[2866] = (layer0_outputs[3552]) ^ (layer0_outputs[1292]);
    assign outputs[2867] = ~(layer0_outputs[5107]) | (layer0_outputs[7102]);
    assign outputs[2868] = layer0_outputs[8600];
    assign outputs[2869] = ~(layer0_outputs[8838]);
    assign outputs[2870] = layer0_outputs[8973];
    assign outputs[2871] = (layer0_outputs[6749]) & (layer0_outputs[1999]);
    assign outputs[2872] = ~(layer0_outputs[2267]);
    assign outputs[2873] = ~(layer0_outputs[3490]) | (layer0_outputs[7644]);
    assign outputs[2874] = ~((layer0_outputs[9952]) | (layer0_outputs[4236]));
    assign outputs[2875] = layer0_outputs[5660];
    assign outputs[2876] = ~(layer0_outputs[185]);
    assign outputs[2877] = ~(layer0_outputs[9740]) | (layer0_outputs[4065]);
    assign outputs[2878] = ~(layer0_outputs[5271]);
    assign outputs[2879] = (layer0_outputs[3722]) & ~(layer0_outputs[7391]);
    assign outputs[2880] = ~((layer0_outputs[2461]) ^ (layer0_outputs[6126]));
    assign outputs[2881] = ~(layer0_outputs[9511]);
    assign outputs[2882] = ~((layer0_outputs[8497]) & (layer0_outputs[1164]));
    assign outputs[2883] = ~(layer0_outputs[9239]);
    assign outputs[2884] = ~(layer0_outputs[8403]);
    assign outputs[2885] = ~(layer0_outputs[4626]) | (layer0_outputs[772]);
    assign outputs[2886] = (layer0_outputs[7392]) ^ (layer0_outputs[2723]);
    assign outputs[2887] = (layer0_outputs[735]) & ~(layer0_outputs[8078]);
    assign outputs[2888] = ~(layer0_outputs[8707]);
    assign outputs[2889] = layer0_outputs[4005];
    assign outputs[2890] = layer0_outputs[4304];
    assign outputs[2891] = (layer0_outputs[4278]) | (layer0_outputs[2204]);
    assign outputs[2892] = (layer0_outputs[6272]) & (layer0_outputs[5927]);
    assign outputs[2893] = layer0_outputs[930];
    assign outputs[2894] = (layer0_outputs[2842]) ^ (layer0_outputs[3055]);
    assign outputs[2895] = layer0_outputs[4291];
    assign outputs[2896] = ~((layer0_outputs[8339]) ^ (layer0_outputs[5324]));
    assign outputs[2897] = layer0_outputs[3077];
    assign outputs[2898] = ~((layer0_outputs[1169]) ^ (layer0_outputs[8232]));
    assign outputs[2899] = ~((layer0_outputs[7022]) ^ (layer0_outputs[7278]));
    assign outputs[2900] = (layer0_outputs[4107]) & (layer0_outputs[6813]);
    assign outputs[2901] = ~((layer0_outputs[2418]) ^ (layer0_outputs[3388]));
    assign outputs[2902] = (layer0_outputs[5340]) & ~(layer0_outputs[6074]);
    assign outputs[2903] = (layer0_outputs[4466]) ^ (layer0_outputs[4449]);
    assign outputs[2904] = ~(layer0_outputs[1085]) | (layer0_outputs[1839]);
    assign outputs[2905] = ~((layer0_outputs[8611]) ^ (layer0_outputs[9812]));
    assign outputs[2906] = (layer0_outputs[4587]) & (layer0_outputs[3730]);
    assign outputs[2907] = (layer0_outputs[7724]) | (layer0_outputs[2843]);
    assign outputs[2908] = ~(layer0_outputs[198]);
    assign outputs[2909] = ~(layer0_outputs[7435]);
    assign outputs[2910] = layer0_outputs[460];
    assign outputs[2911] = layer0_outputs[2608];
    assign outputs[2912] = ~((layer0_outputs[8917]) ^ (layer0_outputs[5239]));
    assign outputs[2913] = ~(layer0_outputs[462]);
    assign outputs[2914] = ~(layer0_outputs[1199]);
    assign outputs[2915] = ~(layer0_outputs[4056]);
    assign outputs[2916] = (layer0_outputs[1918]) & ~(layer0_outputs[2157]);
    assign outputs[2917] = ~(layer0_outputs[761]);
    assign outputs[2918] = ~(layer0_outputs[6072]);
    assign outputs[2919] = (layer0_outputs[8802]) & (layer0_outputs[2830]);
    assign outputs[2920] = ~((layer0_outputs[3697]) ^ (layer0_outputs[3281]));
    assign outputs[2921] = (layer0_outputs[7103]) ^ (layer0_outputs[4736]);
    assign outputs[2922] = (layer0_outputs[5473]) ^ (layer0_outputs[9576]);
    assign outputs[2923] = ~(layer0_outputs[7200]);
    assign outputs[2924] = (layer0_outputs[1315]) ^ (layer0_outputs[2728]);
    assign outputs[2925] = ~(layer0_outputs[548]);
    assign outputs[2926] = (layer0_outputs[6226]) ^ (layer0_outputs[6205]);
    assign outputs[2927] = (layer0_outputs[1910]) | (layer0_outputs[5156]);
    assign outputs[2928] = layer0_outputs[4426];
    assign outputs[2929] = (layer0_outputs[275]) ^ (layer0_outputs[8223]);
    assign outputs[2930] = ~(layer0_outputs[9261]);
    assign outputs[2931] = layer0_outputs[4350];
    assign outputs[2932] = ~(layer0_outputs[3364]) | (layer0_outputs[8392]);
    assign outputs[2933] = (layer0_outputs[1954]) & ~(layer0_outputs[4215]);
    assign outputs[2934] = (layer0_outputs[2051]) | (layer0_outputs[10235]);
    assign outputs[2935] = ~(layer0_outputs[7617]) | (layer0_outputs[2616]);
    assign outputs[2936] = ~(layer0_outputs[9024]) | (layer0_outputs[4623]);
    assign outputs[2937] = (layer0_outputs[156]) & (layer0_outputs[3491]);
    assign outputs[2938] = (layer0_outputs[7692]) ^ (layer0_outputs[9749]);
    assign outputs[2939] = layer0_outputs[9504];
    assign outputs[2940] = ~((layer0_outputs[6626]) ^ (layer0_outputs[9348]));
    assign outputs[2941] = ~(layer0_outputs[4586]);
    assign outputs[2942] = layer0_outputs[871];
    assign outputs[2943] = (layer0_outputs[7010]) & (layer0_outputs[14]);
    assign outputs[2944] = (layer0_outputs[9226]) & (layer0_outputs[3963]);
    assign outputs[2945] = layer0_outputs[3358];
    assign outputs[2946] = ~(layer0_outputs[2076]);
    assign outputs[2947] = layer0_outputs[9771];
    assign outputs[2948] = layer0_outputs[3843];
    assign outputs[2949] = (layer0_outputs[9606]) & ~(layer0_outputs[9700]);
    assign outputs[2950] = layer0_outputs[4001];
    assign outputs[2951] = layer0_outputs[2281];
    assign outputs[2952] = layer0_outputs[6750];
    assign outputs[2953] = ~((layer0_outputs[6169]) | (layer0_outputs[7375]));
    assign outputs[2954] = layer0_outputs[3831];
    assign outputs[2955] = ~(layer0_outputs[341]);
    assign outputs[2956] = ~((layer0_outputs[7673]) & (layer0_outputs[3559]));
    assign outputs[2957] = ~(layer0_outputs[3494]);
    assign outputs[2958] = ~(layer0_outputs[8580]);
    assign outputs[2959] = ~(layer0_outputs[3247]);
    assign outputs[2960] = ~((layer0_outputs[6483]) & (layer0_outputs[3927]));
    assign outputs[2961] = (layer0_outputs[3362]) ^ (layer0_outputs[3447]);
    assign outputs[2962] = layer0_outputs[9958];
    assign outputs[2963] = ~(layer0_outputs[9286]);
    assign outputs[2964] = layer0_outputs[2848];
    assign outputs[2965] = (layer0_outputs[5288]) & ~(layer0_outputs[8620]);
    assign outputs[2966] = ~(layer0_outputs[4976]);
    assign outputs[2967] = layer0_outputs[4132];
    assign outputs[2968] = ~(layer0_outputs[8643]);
    assign outputs[2969] = ~(layer0_outputs[9163]) | (layer0_outputs[7339]);
    assign outputs[2970] = ~(layer0_outputs[3580]) | (layer0_outputs[228]);
    assign outputs[2971] = layer0_outputs[5049];
    assign outputs[2972] = ~(layer0_outputs[7772]) | (layer0_outputs[5230]);
    assign outputs[2973] = (layer0_outputs[199]) ^ (layer0_outputs[1985]);
    assign outputs[2974] = ~(layer0_outputs[5160]);
    assign outputs[2975] = ~(layer0_outputs[5803]) | (layer0_outputs[5320]);
    assign outputs[2976] = (layer0_outputs[5446]) & ~(layer0_outputs[3844]);
    assign outputs[2977] = layer0_outputs[8836];
    assign outputs[2978] = ~((layer0_outputs[4732]) & (layer0_outputs[1454]));
    assign outputs[2979] = ~((layer0_outputs[9665]) ^ (layer0_outputs[7775]));
    assign outputs[2980] = layer0_outputs[2141];
    assign outputs[2981] = (layer0_outputs[6572]) | (layer0_outputs[8369]);
    assign outputs[2982] = (layer0_outputs[5951]) ^ (layer0_outputs[7947]);
    assign outputs[2983] = (layer0_outputs[1521]) & (layer0_outputs[8192]);
    assign outputs[2984] = layer0_outputs[5033];
    assign outputs[2985] = ~(layer0_outputs[1713]);
    assign outputs[2986] = layer0_outputs[3981];
    assign outputs[2987] = ~(layer0_outputs[7519]);
    assign outputs[2988] = layer0_outputs[9895];
    assign outputs[2989] = (layer0_outputs[4010]) & (layer0_outputs[2348]);
    assign outputs[2990] = (layer0_outputs[5615]) ^ (layer0_outputs[1133]);
    assign outputs[2991] = ~((layer0_outputs[5258]) ^ (layer0_outputs[5352]));
    assign outputs[2992] = layer0_outputs[1588];
    assign outputs[2993] = ~(layer0_outputs[9560]) | (layer0_outputs[4019]);
    assign outputs[2994] = layer0_outputs[3087];
    assign outputs[2995] = ~(layer0_outputs[1312]);
    assign outputs[2996] = ~(layer0_outputs[820]);
    assign outputs[2997] = ~(layer0_outputs[6908]);
    assign outputs[2998] = ~(layer0_outputs[7670]);
    assign outputs[2999] = ~((layer0_outputs[9434]) ^ (layer0_outputs[10071]));
    assign outputs[3000] = ~(layer0_outputs[5835]);
    assign outputs[3001] = ~((layer0_outputs[3847]) & (layer0_outputs[2693]));
    assign outputs[3002] = layer0_outputs[4576];
    assign outputs[3003] = layer0_outputs[3750];
    assign outputs[3004] = ~((layer0_outputs[5702]) & (layer0_outputs[3257]));
    assign outputs[3005] = ~((layer0_outputs[2203]) & (layer0_outputs[4333]));
    assign outputs[3006] = ~((layer0_outputs[41]) ^ (layer0_outputs[9564]));
    assign outputs[3007] = ~(layer0_outputs[4942]);
    assign outputs[3008] = (layer0_outputs[10197]) ^ (layer0_outputs[3481]);
    assign outputs[3009] = layer0_outputs[3610];
    assign outputs[3010] = ~((layer0_outputs[9180]) | (layer0_outputs[8618]));
    assign outputs[3011] = ~(layer0_outputs[3796]) | (layer0_outputs[10083]);
    assign outputs[3012] = (layer0_outputs[5774]) & (layer0_outputs[4920]);
    assign outputs[3013] = ~((layer0_outputs[9913]) | (layer0_outputs[162]));
    assign outputs[3014] = ~(layer0_outputs[6550]);
    assign outputs[3015] = ~(layer0_outputs[7393]);
    assign outputs[3016] = ~(layer0_outputs[5699]);
    assign outputs[3017] = ~((layer0_outputs[1899]) ^ (layer0_outputs[7132]));
    assign outputs[3018] = ~((layer0_outputs[6323]) ^ (layer0_outputs[2412]));
    assign outputs[3019] = ~(layer0_outputs[5810]) | (layer0_outputs[2277]);
    assign outputs[3020] = (layer0_outputs[5436]) & ~(layer0_outputs[2394]);
    assign outputs[3021] = layer0_outputs[2295];
    assign outputs[3022] = ~(layer0_outputs[3992]);
    assign outputs[3023] = ~((layer0_outputs[7153]) ^ (layer0_outputs[852]));
    assign outputs[3024] = ~(layer0_outputs[2526]) | (layer0_outputs[7684]);
    assign outputs[3025] = layer0_outputs[5553];
    assign outputs[3026] = ~((layer0_outputs[9085]) ^ (layer0_outputs[381]));
    assign outputs[3027] = ~((layer0_outputs[9020]) ^ (layer0_outputs[6447]));
    assign outputs[3028] = ~((layer0_outputs[8629]) & (layer0_outputs[7605]));
    assign outputs[3029] = (layer0_outputs[8017]) | (layer0_outputs[2666]);
    assign outputs[3030] = layer0_outputs[961];
    assign outputs[3031] = layer0_outputs[8831];
    assign outputs[3032] = ~(layer0_outputs[9051]);
    assign outputs[3033] = layer0_outputs[2329];
    assign outputs[3034] = ~((layer0_outputs[1190]) | (layer0_outputs[267]));
    assign outputs[3035] = (layer0_outputs[7655]) ^ (layer0_outputs[5099]);
    assign outputs[3036] = ~(layer0_outputs[656]);
    assign outputs[3037] = ~((layer0_outputs[6712]) | (layer0_outputs[5087]));
    assign outputs[3038] = (layer0_outputs[6330]) & ~(layer0_outputs[6951]);
    assign outputs[3039] = layer0_outputs[1217];
    assign outputs[3040] = (layer0_outputs[10124]) | (layer0_outputs[9393]);
    assign outputs[3041] = ~(layer0_outputs[5105]);
    assign outputs[3042] = (layer0_outputs[4303]) ^ (layer0_outputs[1421]);
    assign outputs[3043] = (layer0_outputs[386]) & (layer0_outputs[5508]);
    assign outputs[3044] = ~(layer0_outputs[10092]) | (layer0_outputs[5031]);
    assign outputs[3045] = ~((layer0_outputs[404]) ^ (layer0_outputs[8972]));
    assign outputs[3046] = ~(layer0_outputs[7181]);
    assign outputs[3047] = ~(layer0_outputs[1205]);
    assign outputs[3048] = layer0_outputs[7731];
    assign outputs[3049] = layer0_outputs[1622];
    assign outputs[3050] = (layer0_outputs[9925]) ^ (layer0_outputs[8012]);
    assign outputs[3051] = ~(layer0_outputs[609]);
    assign outputs[3052] = ~(layer0_outputs[4151]);
    assign outputs[3053] = layer0_outputs[5063];
    assign outputs[3054] = ~(layer0_outputs[6664]);
    assign outputs[3055] = ~(layer0_outputs[3139]);
    assign outputs[3056] = ~(layer0_outputs[7942]) | (layer0_outputs[6173]);
    assign outputs[3057] = ~(layer0_outputs[1528]) | (layer0_outputs[4311]);
    assign outputs[3058] = layer0_outputs[2169];
    assign outputs[3059] = ~(layer0_outputs[6720]) | (layer0_outputs[7793]);
    assign outputs[3060] = ~(layer0_outputs[2763]) | (layer0_outputs[4948]);
    assign outputs[3061] = layer0_outputs[3923];
    assign outputs[3062] = layer0_outputs[7595];
    assign outputs[3063] = ~(layer0_outputs[8345]);
    assign outputs[3064] = ~(layer0_outputs[1278]);
    assign outputs[3065] = ~(layer0_outputs[3353]);
    assign outputs[3066] = layer0_outputs[9501];
    assign outputs[3067] = (layer0_outputs[6624]) & (layer0_outputs[2568]);
    assign outputs[3068] = ~(layer0_outputs[9088]);
    assign outputs[3069] = layer0_outputs[1390];
    assign outputs[3070] = ~((layer0_outputs[1479]) ^ (layer0_outputs[9713]));
    assign outputs[3071] = ~(layer0_outputs[5211]);
    assign outputs[3072] = ~(layer0_outputs[9804]) | (layer0_outputs[2728]);
    assign outputs[3073] = ~(layer0_outputs[6236]);
    assign outputs[3074] = layer0_outputs[5652];
    assign outputs[3075] = ~(layer0_outputs[2485]);
    assign outputs[3076] = ~((layer0_outputs[4741]) ^ (layer0_outputs[5368]));
    assign outputs[3077] = ~(layer0_outputs[7536]);
    assign outputs[3078] = layer0_outputs[9026];
    assign outputs[3079] = layer0_outputs[7597];
    assign outputs[3080] = ~(layer0_outputs[7759]);
    assign outputs[3081] = ~((layer0_outputs[3517]) ^ (layer0_outputs[6952]));
    assign outputs[3082] = ~(layer0_outputs[3411]);
    assign outputs[3083] = (layer0_outputs[5157]) ^ (layer0_outputs[243]);
    assign outputs[3084] = ~(layer0_outputs[8860]) | (layer0_outputs[4202]);
    assign outputs[3085] = (layer0_outputs[9423]) & (layer0_outputs[7537]);
    assign outputs[3086] = ~(layer0_outputs[5497]);
    assign outputs[3087] = ~(layer0_outputs[5015]);
    assign outputs[3088] = layer0_outputs[8675];
    assign outputs[3089] = layer0_outputs[2961];
    assign outputs[3090] = ~(layer0_outputs[2276]) | (layer0_outputs[9601]);
    assign outputs[3091] = ~((layer0_outputs[2468]) & (layer0_outputs[6347]));
    assign outputs[3092] = layer0_outputs[2138];
    assign outputs[3093] = ~(layer0_outputs[1325]) | (layer0_outputs[9025]);
    assign outputs[3094] = ~(layer0_outputs[5689]);
    assign outputs[3095] = (layer0_outputs[1863]) ^ (layer0_outputs[3186]);
    assign outputs[3096] = layer0_outputs[7405];
    assign outputs[3097] = layer0_outputs[2111];
    assign outputs[3098] = ~((layer0_outputs[2393]) ^ (layer0_outputs[111]));
    assign outputs[3099] = (layer0_outputs[3480]) ^ (layer0_outputs[10196]);
    assign outputs[3100] = ~(layer0_outputs[4902]);
    assign outputs[3101] = ~(layer0_outputs[4376]);
    assign outputs[3102] = (layer0_outputs[1605]) & ~(layer0_outputs[3043]);
    assign outputs[3103] = layer0_outputs[595];
    assign outputs[3104] = ~(layer0_outputs[8589]);
    assign outputs[3105] = ~(layer0_outputs[7524]) | (layer0_outputs[9938]);
    assign outputs[3106] = layer0_outputs[5953];
    assign outputs[3107] = (layer0_outputs[8129]) | (layer0_outputs[7434]);
    assign outputs[3108] = (layer0_outputs[68]) & ~(layer0_outputs[3268]);
    assign outputs[3109] = ~(layer0_outputs[7847]);
    assign outputs[3110] = layer0_outputs[6689];
    assign outputs[3111] = ~(layer0_outputs[5270]);
    assign outputs[3112] = (layer0_outputs[245]) & ~(layer0_outputs[468]);
    assign outputs[3113] = ~((layer0_outputs[6605]) & (layer0_outputs[4428]));
    assign outputs[3114] = ~((layer0_outputs[471]) ^ (layer0_outputs[7751]));
    assign outputs[3115] = ~((layer0_outputs[3474]) ^ (layer0_outputs[7788]));
    assign outputs[3116] = layer0_outputs[8389];
    assign outputs[3117] = layer0_outputs[8245];
    assign outputs[3118] = layer0_outputs[9191];
    assign outputs[3119] = ~((layer0_outputs[4399]) ^ (layer0_outputs[6075]));
    assign outputs[3120] = ~((layer0_outputs[3947]) ^ (layer0_outputs[549]));
    assign outputs[3121] = ~(layer0_outputs[8554]);
    assign outputs[3122] = layer0_outputs[644];
    assign outputs[3123] = ~(layer0_outputs[2656]) | (layer0_outputs[9994]);
    assign outputs[3124] = ~((layer0_outputs[10018]) ^ (layer0_outputs[263]));
    assign outputs[3125] = layer0_outputs[168];
    assign outputs[3126] = ~(layer0_outputs[10190]);
    assign outputs[3127] = ~(layer0_outputs[9995]);
    assign outputs[3128] = (layer0_outputs[2920]) & ~(layer0_outputs[576]);
    assign outputs[3129] = ~((layer0_outputs[2685]) ^ (layer0_outputs[6599]));
    assign outputs[3130] = ~(layer0_outputs[693]);
    assign outputs[3131] = ~(layer0_outputs[5502]);
    assign outputs[3132] = (layer0_outputs[600]) ^ (layer0_outputs[4039]);
    assign outputs[3133] = ~(layer0_outputs[6257]);
    assign outputs[3134] = ~(layer0_outputs[7530]);
    assign outputs[3135] = (layer0_outputs[9059]) & ~(layer0_outputs[5539]);
    assign outputs[3136] = (layer0_outputs[4236]) | (layer0_outputs[10153]);
    assign outputs[3137] = (layer0_outputs[1901]) ^ (layer0_outputs[6277]);
    assign outputs[3138] = ~(layer0_outputs[2444]);
    assign outputs[3139] = (layer0_outputs[9149]) & ~(layer0_outputs[6967]);
    assign outputs[3140] = (layer0_outputs[1563]) ^ (layer0_outputs[7897]);
    assign outputs[3141] = ~(layer0_outputs[3654]);
    assign outputs[3142] = ~(layer0_outputs[5737]);
    assign outputs[3143] = (layer0_outputs[9990]) ^ (layer0_outputs[3296]);
    assign outputs[3144] = ~((layer0_outputs[8156]) | (layer0_outputs[3057]));
    assign outputs[3145] = (layer0_outputs[4009]) & ~(layer0_outputs[2982]);
    assign outputs[3146] = layer0_outputs[2231];
    assign outputs[3147] = (layer0_outputs[2316]) & (layer0_outputs[9011]);
    assign outputs[3148] = ~(layer0_outputs[9555]);
    assign outputs[3149] = ~(layer0_outputs[5818]);
    assign outputs[3150] = ~((layer0_outputs[2716]) ^ (layer0_outputs[9983]));
    assign outputs[3151] = (layer0_outputs[7215]) & ~(layer0_outputs[7440]);
    assign outputs[3152] = (layer0_outputs[3837]) & (layer0_outputs[3611]);
    assign outputs[3153] = ~(layer0_outputs[8621]);
    assign outputs[3154] = (layer0_outputs[3500]) & ~(layer0_outputs[986]);
    assign outputs[3155] = layer0_outputs[1821];
    assign outputs[3156] = ~((layer0_outputs[6067]) & (layer0_outputs[9962]));
    assign outputs[3157] = layer0_outputs[8222];
    assign outputs[3158] = ~(layer0_outputs[4375]);
    assign outputs[3159] = (layer0_outputs[1191]) & ~(layer0_outputs[8113]);
    assign outputs[3160] = layer0_outputs[5703];
    assign outputs[3161] = ~(layer0_outputs[5264]);
    assign outputs[3162] = (layer0_outputs[2439]) & ~(layer0_outputs[3392]);
    assign outputs[3163] = ~((layer0_outputs[2627]) ^ (layer0_outputs[8467]));
    assign outputs[3164] = (layer0_outputs[3849]) ^ (layer0_outputs[2919]);
    assign outputs[3165] = (layer0_outputs[7947]) ^ (layer0_outputs[1006]);
    assign outputs[3166] = (layer0_outputs[8304]) & (layer0_outputs[4684]);
    assign outputs[3167] = layer0_outputs[2917];
    assign outputs[3168] = ~((layer0_outputs[1758]) & (layer0_outputs[1267]));
    assign outputs[3169] = layer0_outputs[6491];
    assign outputs[3170] = ~(layer0_outputs[6587]);
    assign outputs[3171] = ~(layer0_outputs[2101]);
    assign outputs[3172] = layer0_outputs[9241];
    assign outputs[3173] = ~(layer0_outputs[6703]);
    assign outputs[3174] = ~(layer0_outputs[3528]);
    assign outputs[3175] = layer0_outputs[4394];
    assign outputs[3176] = (layer0_outputs[2311]) ^ (layer0_outputs[5801]);
    assign outputs[3177] = layer0_outputs[9627];
    assign outputs[3178] = ~((layer0_outputs[7381]) | (layer0_outputs[3482]));
    assign outputs[3179] = layer0_outputs[1873];
    assign outputs[3180] = (layer0_outputs[5375]) & (layer0_outputs[5718]);
    assign outputs[3181] = ~((layer0_outputs[5847]) ^ (layer0_outputs[4728]));
    assign outputs[3182] = layer0_outputs[8413];
    assign outputs[3183] = ~((layer0_outputs[7560]) | (layer0_outputs[8386]));
    assign outputs[3184] = ~(layer0_outputs[2145]);
    assign outputs[3185] = layer0_outputs[6223];
    assign outputs[3186] = ~(layer0_outputs[3120]);
    assign outputs[3187] = ~((layer0_outputs[8303]) ^ (layer0_outputs[8532]));
    assign outputs[3188] = (layer0_outputs[7444]) & ~(layer0_outputs[3588]);
    assign outputs[3189] = ~((layer0_outputs[5557]) ^ (layer0_outputs[3840]));
    assign outputs[3190] = layer0_outputs[5778];
    assign outputs[3191] = ~((layer0_outputs[3064]) ^ (layer0_outputs[2892]));
    assign outputs[3192] = ~(layer0_outputs[4816]);
    assign outputs[3193] = layer0_outputs[4622];
    assign outputs[3194] = ~((layer0_outputs[1912]) ^ (layer0_outputs[7766]));
    assign outputs[3195] = ~(layer0_outputs[6398]) | (layer0_outputs[4455]);
    assign outputs[3196] = layer0_outputs[2483];
    assign outputs[3197] = ~(layer0_outputs[4705]);
    assign outputs[3198] = ~((layer0_outputs[1780]) | (layer0_outputs[4280]));
    assign outputs[3199] = ~(layer0_outputs[7248]) | (layer0_outputs[6376]);
    assign outputs[3200] = ~((layer0_outputs[9775]) | (layer0_outputs[5843]));
    assign outputs[3201] = (layer0_outputs[5663]) ^ (layer0_outputs[4511]);
    assign outputs[3202] = ~(layer0_outputs[9823]) | (layer0_outputs[7702]);
    assign outputs[3203] = (layer0_outputs[2987]) ^ (layer0_outputs[7477]);
    assign outputs[3204] = ~(layer0_outputs[5973]);
    assign outputs[3205] = ~((layer0_outputs[544]) ^ (layer0_outputs[8847]));
    assign outputs[3206] = layer0_outputs[2202];
    assign outputs[3207] = ~(layer0_outputs[2228]);
    assign outputs[3208] = layer0_outputs[8324];
    assign outputs[3209] = (layer0_outputs[9454]) & (layer0_outputs[2360]);
    assign outputs[3210] = ~(layer0_outputs[1767]);
    assign outputs[3211] = (layer0_outputs[9434]) ^ (layer0_outputs[9278]);
    assign outputs[3212] = ~(layer0_outputs[6463]);
    assign outputs[3213] = ~(layer0_outputs[9597]);
    assign outputs[3214] = ~(layer0_outputs[9121]);
    assign outputs[3215] = layer0_outputs[5524];
    assign outputs[3216] = ~(layer0_outputs[831]) | (layer0_outputs[9117]);
    assign outputs[3217] = layer0_outputs[9018];
    assign outputs[3218] = ~((layer0_outputs[5700]) ^ (layer0_outputs[3946]));
    assign outputs[3219] = layer0_outputs[3426];
    assign outputs[3220] = layer0_outputs[7921];
    assign outputs[3221] = layer0_outputs[9644];
    assign outputs[3222] = ~((layer0_outputs[148]) ^ (layer0_outputs[2582]));
    assign outputs[3223] = layer0_outputs[3752];
    assign outputs[3224] = layer0_outputs[8848];
    assign outputs[3225] = layer0_outputs[1038];
    assign outputs[3226] = (layer0_outputs[5492]) ^ (layer0_outputs[7146]);
    assign outputs[3227] = (layer0_outputs[1562]) ^ (layer0_outputs[5894]);
    assign outputs[3228] = ~(layer0_outputs[7411]);
    assign outputs[3229] = ~(layer0_outputs[3481]);
    assign outputs[3230] = ~(layer0_outputs[3443]) | (layer0_outputs[2896]);
    assign outputs[3231] = ~(layer0_outputs[4002]) | (layer0_outputs[2353]);
    assign outputs[3232] = layer0_outputs[2708];
    assign outputs[3233] = (layer0_outputs[7632]) & ~(layer0_outputs[10060]);
    assign outputs[3234] = (layer0_outputs[8245]) & ~(layer0_outputs[2501]);
    assign outputs[3235] = (layer0_outputs[9536]) ^ (layer0_outputs[10212]);
    assign outputs[3236] = layer0_outputs[2258];
    assign outputs[3237] = (layer0_outputs[720]) ^ (layer0_outputs[9491]);
    assign outputs[3238] = ~(layer0_outputs[4513]);
    assign outputs[3239] = (layer0_outputs[2762]) & ~(layer0_outputs[4704]);
    assign outputs[3240] = layer0_outputs[8216];
    assign outputs[3241] = layer0_outputs[4577];
    assign outputs[3242] = layer0_outputs[7729];
    assign outputs[3243] = ~(layer0_outputs[8591]);
    assign outputs[3244] = (layer0_outputs[5312]) ^ (layer0_outputs[6735]);
    assign outputs[3245] = layer0_outputs[8982];
    assign outputs[3246] = ~(layer0_outputs[8285]);
    assign outputs[3247] = ~(layer0_outputs[9285]);
    assign outputs[3248] = (layer0_outputs[8738]) & ~(layer0_outputs[7424]);
    assign outputs[3249] = (layer0_outputs[1719]) & ~(layer0_outputs[3873]);
    assign outputs[3250] = layer0_outputs[3943];
    assign outputs[3251] = ~((layer0_outputs[5950]) & (layer0_outputs[6296]));
    assign outputs[3252] = ~((layer0_outputs[7394]) | (layer0_outputs[656]));
    assign outputs[3253] = ~(layer0_outputs[9471]);
    assign outputs[3254] = (layer0_outputs[2081]) & ~(layer0_outputs[4393]);
    assign outputs[3255] = ~((layer0_outputs[1773]) ^ (layer0_outputs[5364]));
    assign outputs[3256] = (layer0_outputs[778]) & ~(layer0_outputs[4037]);
    assign outputs[3257] = ~((layer0_outputs[3508]) ^ (layer0_outputs[1074]));
    assign outputs[3258] = layer0_outputs[4831];
    assign outputs[3259] = ~(layer0_outputs[6257]);
    assign outputs[3260] = layer0_outputs[1158];
    assign outputs[3261] = layer0_outputs[7846];
    assign outputs[3262] = ~((layer0_outputs[342]) ^ (layer0_outputs[3072]));
    assign outputs[3263] = ~((layer0_outputs[8340]) ^ (layer0_outputs[10148]));
    assign outputs[3264] = ~((layer0_outputs[6698]) ^ (layer0_outputs[1942]));
    assign outputs[3265] = layer0_outputs[3902];
    assign outputs[3266] = (layer0_outputs[2971]) ^ (layer0_outputs[3538]);
    assign outputs[3267] = ~(layer0_outputs[2838]);
    assign outputs[3268] = layer0_outputs[1245];
    assign outputs[3269] = ~(layer0_outputs[5758]);
    assign outputs[3270] = (layer0_outputs[5452]) & ~(layer0_outputs[7141]);
    assign outputs[3271] = ~(layer0_outputs[4777]);
    assign outputs[3272] = (layer0_outputs[42]) & ~(layer0_outputs[8685]);
    assign outputs[3273] = layer0_outputs[1798];
    assign outputs[3274] = ~(layer0_outputs[293]) | (layer0_outputs[9990]);
    assign outputs[3275] = (layer0_outputs[4174]) & (layer0_outputs[10226]);
    assign outputs[3276] = ~((layer0_outputs[1991]) ^ (layer0_outputs[4581]));
    assign outputs[3277] = (layer0_outputs[3242]) | (layer0_outputs[1387]);
    assign outputs[3278] = layer0_outputs[8372];
    assign outputs[3279] = layer0_outputs[4814];
    assign outputs[3280] = ~((layer0_outputs[5706]) | (layer0_outputs[7094]));
    assign outputs[3281] = ~(layer0_outputs[491]);
    assign outputs[3282] = ~((layer0_outputs[8393]) ^ (layer0_outputs[538]));
    assign outputs[3283] = ~(layer0_outputs[5247]);
    assign outputs[3284] = ~(layer0_outputs[3065]);
    assign outputs[3285] = ~(layer0_outputs[1970]);
    assign outputs[3286] = ~(layer0_outputs[1446]);
    assign outputs[3287] = ~((layer0_outputs[6665]) ^ (layer0_outputs[2021]));
    assign outputs[3288] = ~((layer0_outputs[335]) ^ (layer0_outputs[1001]));
    assign outputs[3289] = ~((layer0_outputs[1045]) & (layer0_outputs[8720]));
    assign outputs[3290] = layer0_outputs[1420];
    assign outputs[3291] = (layer0_outputs[6230]) & (layer0_outputs[2615]);
    assign outputs[3292] = layer0_outputs[3527];
    assign outputs[3293] = layer0_outputs[4495];
    assign outputs[3294] = ~((layer0_outputs[8728]) | (layer0_outputs[6301]));
    assign outputs[3295] = ~(layer0_outputs[1736]);
    assign outputs[3296] = layer0_outputs[10075];
    assign outputs[3297] = ~((layer0_outputs[3311]) | (layer0_outputs[10138]));
    assign outputs[3298] = layer0_outputs[9360];
    assign outputs[3299] = (layer0_outputs[3710]) & (layer0_outputs[942]);
    assign outputs[3300] = ~((layer0_outputs[9655]) | (layer0_outputs[8200]));
    assign outputs[3301] = layer0_outputs[3444];
    assign outputs[3302] = (layer0_outputs[8331]) ^ (layer0_outputs[4998]);
    assign outputs[3303] = ~(layer0_outputs[5297]);
    assign outputs[3304] = ~(layer0_outputs[9181]);
    assign outputs[3305] = ~((layer0_outputs[4462]) & (layer0_outputs[8032]));
    assign outputs[3306] = (layer0_outputs[122]) ^ (layer0_outputs[1950]);
    assign outputs[3307] = (layer0_outputs[7492]) & ~(layer0_outputs[3009]);
    assign outputs[3308] = (layer0_outputs[150]) ^ (layer0_outputs[9813]);
    assign outputs[3309] = (layer0_outputs[3853]) & ~(layer0_outputs[5715]);
    assign outputs[3310] = ~(layer0_outputs[8932]);
    assign outputs[3311] = layer0_outputs[2057];
    assign outputs[3312] = layer0_outputs[4167];
    assign outputs[3313] = ~((layer0_outputs[1852]) | (layer0_outputs[5910]));
    assign outputs[3314] = (layer0_outputs[1803]) & (layer0_outputs[2555]);
    assign outputs[3315] = ~((layer0_outputs[4182]) ^ (layer0_outputs[3611]));
    assign outputs[3316] = (layer0_outputs[9818]) ^ (layer0_outputs[5749]);
    assign outputs[3317] = layer0_outputs[4424];
    assign outputs[3318] = ~(layer0_outputs[2189]);
    assign outputs[3319] = layer0_outputs[6528];
    assign outputs[3320] = ~(layer0_outputs[4553]);
    assign outputs[3321] = (layer0_outputs[9352]) & ~(layer0_outputs[4151]);
    assign outputs[3322] = ~(layer0_outputs[8869]);
    assign outputs[3323] = layer0_outputs[9888];
    assign outputs[3324] = layer0_outputs[3501];
    assign outputs[3325] = 1'b0;
    assign outputs[3326] = (layer0_outputs[1824]) & ~(layer0_outputs[8783]);
    assign outputs[3327] = layer0_outputs[6543];
    assign outputs[3328] = ~(layer0_outputs[10137]);
    assign outputs[3329] = ~(layer0_outputs[8872]);
    assign outputs[3330] = layer0_outputs[2591];
    assign outputs[3331] = (layer0_outputs[3492]) & ~(layer0_outputs[2052]);
    assign outputs[3332] = ~(layer0_outputs[8796]);
    assign outputs[3333] = layer0_outputs[5330];
    assign outputs[3334] = ~((layer0_outputs[7220]) ^ (layer0_outputs[6927]));
    assign outputs[3335] = ~((layer0_outputs[1120]) ^ (layer0_outputs[2387]));
    assign outputs[3336] = ~(layer0_outputs[94]);
    assign outputs[3337] = ~((layer0_outputs[8273]) | (layer0_outputs[5874]));
    assign outputs[3338] = layer0_outputs[6314];
    assign outputs[3339] = (layer0_outputs[6995]) | (layer0_outputs[6342]);
    assign outputs[3340] = layer0_outputs[10114];
    assign outputs[3341] = layer0_outputs[832];
    assign outputs[3342] = ~(layer0_outputs[7023]);
    assign outputs[3343] = ~(layer0_outputs[4378]);
    assign outputs[3344] = layer0_outputs[129];
    assign outputs[3345] = ~(layer0_outputs[60]) | (layer0_outputs[9568]);
    assign outputs[3346] = ~(layer0_outputs[3365]);
    assign outputs[3347] = ~(layer0_outputs[3375]) | (layer0_outputs[7466]);
    assign outputs[3348] = layer0_outputs[4338];
    assign outputs[3349] = ~(layer0_outputs[3583]);
    assign outputs[3350] = (layer0_outputs[6496]) ^ (layer0_outputs[3498]);
    assign outputs[3351] = ~(layer0_outputs[900]);
    assign outputs[3352] = ~((layer0_outputs[3577]) | (layer0_outputs[3723]));
    assign outputs[3353] = ~(layer0_outputs[6551]) | (layer0_outputs[6061]);
    assign outputs[3354] = ~(layer0_outputs[163]);
    assign outputs[3355] = layer0_outputs[2328];
    assign outputs[3356] = layer0_outputs[7015];
    assign outputs[3357] = ~(layer0_outputs[3015]);
    assign outputs[3358] = (layer0_outputs[2275]) | (layer0_outputs[7026]);
    assign outputs[3359] = ~(layer0_outputs[2945]);
    assign outputs[3360] = (layer0_outputs[1149]) ^ (layer0_outputs[1926]);
    assign outputs[3361] = (layer0_outputs[1031]) & (layer0_outputs[4940]);
    assign outputs[3362] = layer0_outputs[9199];
    assign outputs[3363] = ~(layer0_outputs[8506]) | (layer0_outputs[7033]);
    assign outputs[3364] = layer0_outputs[1592];
    assign outputs[3365] = layer0_outputs[2636];
    assign outputs[3366] = layer0_outputs[9715];
    assign outputs[3367] = layer0_outputs[5281];
    assign outputs[3368] = ~(layer0_outputs[6553]);
    assign outputs[3369] = layer0_outputs[2667];
    assign outputs[3370] = layer0_outputs[4941];
    assign outputs[3371] = layer0_outputs[320];
    assign outputs[3372] = ~((layer0_outputs[6054]) ^ (layer0_outputs[3150]));
    assign outputs[3373] = (layer0_outputs[6556]) & ~(layer0_outputs[4544]);
    assign outputs[3374] = (layer0_outputs[2153]) & (layer0_outputs[9848]);
    assign outputs[3375] = ~(layer0_outputs[9007]);
    assign outputs[3376] = ~((layer0_outputs[5257]) ^ (layer0_outputs[4860]));
    assign outputs[3377] = layer0_outputs[8735];
    assign outputs[3378] = layer0_outputs[476];
    assign outputs[3379] = ~(layer0_outputs[1737]);
    assign outputs[3380] = ~((layer0_outputs[5831]) ^ (layer0_outputs[3308]));
    assign outputs[3381] = layer0_outputs[9235];
    assign outputs[3382] = ~(layer0_outputs[6006]);
    assign outputs[3383] = ~(layer0_outputs[8943]);
    assign outputs[3384] = layer0_outputs[2679];
    assign outputs[3385] = ~(layer0_outputs[459]);
    assign outputs[3386] = layer0_outputs[8144];
    assign outputs[3387] = ~(layer0_outputs[8226]);
    assign outputs[3388] = (layer0_outputs[3029]) & (layer0_outputs[8227]);
    assign outputs[3389] = ~(layer0_outputs[5384]);
    assign outputs[3390] = ~(layer0_outputs[6617]);
    assign outputs[3391] = layer0_outputs[4293];
    assign outputs[3392] = ~((layer0_outputs[677]) ^ (layer0_outputs[4657]));
    assign outputs[3393] = ~((layer0_outputs[735]) & (layer0_outputs[5190]));
    assign outputs[3394] = layer0_outputs[1949];
    assign outputs[3395] = ~(layer0_outputs[8590]);
    assign outputs[3396] = (layer0_outputs[7407]) | (layer0_outputs[3007]);
    assign outputs[3397] = (layer0_outputs[1082]) ^ (layer0_outputs[6547]);
    assign outputs[3398] = ~((layer0_outputs[2950]) ^ (layer0_outputs[262]));
    assign outputs[3399] = ~(layer0_outputs[1149]) | (layer0_outputs[2355]);
    assign outputs[3400] = ~(layer0_outputs[7396]);
    assign outputs[3401] = layer0_outputs[9274];
    assign outputs[3402] = (layer0_outputs[8992]) & ~(layer0_outputs[6974]);
    assign outputs[3403] = ~(layer0_outputs[10203]);
    assign outputs[3404] = (layer0_outputs[8579]) & ~(layer0_outputs[9931]);
    assign outputs[3405] = ~((layer0_outputs[3026]) | (layer0_outputs[5973]));
    assign outputs[3406] = layer0_outputs[4699];
    assign outputs[3407] = layer0_outputs[5047];
    assign outputs[3408] = ~((layer0_outputs[6694]) & (layer0_outputs[4272]));
    assign outputs[3409] = ~(layer0_outputs[6190]);
    assign outputs[3410] = layer0_outputs[8404];
    assign outputs[3411] = (layer0_outputs[6834]) ^ (layer0_outputs[9971]);
    assign outputs[3412] = ~(layer0_outputs[6000]);
    assign outputs[3413] = ~(layer0_outputs[8592]);
    assign outputs[3414] = ~(layer0_outputs[9722]);
    assign outputs[3415] = ~(layer0_outputs[4094]);
    assign outputs[3416] = layer0_outputs[10150];
    assign outputs[3417] = ~(layer0_outputs[9225]);
    assign outputs[3418] = layer0_outputs[8475];
    assign outputs[3419] = ~(layer0_outputs[2287]);
    assign outputs[3420] = ~((layer0_outputs[4822]) ^ (layer0_outputs[1947]));
    assign outputs[3421] = layer0_outputs[3128];
    assign outputs[3422] = (layer0_outputs[4803]) & ~(layer0_outputs[8059]);
    assign outputs[3423] = ~(layer0_outputs[9193]);
    assign outputs[3424] = layer0_outputs[4264];
    assign outputs[3425] = (layer0_outputs[6359]) & ~(layer0_outputs[5805]);
    assign outputs[3426] = ~(layer0_outputs[101]);
    assign outputs[3427] = layer0_outputs[3426];
    assign outputs[3428] = (layer0_outputs[1667]) ^ (layer0_outputs[9095]);
    assign outputs[3429] = ~(layer0_outputs[7272]);
    assign outputs[3430] = ~(layer0_outputs[5440]);
    assign outputs[3431] = layer0_outputs[2955];
    assign outputs[3432] = layer0_outputs[9480];
    assign outputs[3433] = ~(layer0_outputs[9767]);
    assign outputs[3434] = (layer0_outputs[4391]) & ~(layer0_outputs[3515]);
    assign outputs[3435] = layer0_outputs[8670];
    assign outputs[3436] = ~(layer0_outputs[7133]);
    assign outputs[3437] = layer0_outputs[9053];
    assign outputs[3438] = (layer0_outputs[4594]) & ~(layer0_outputs[596]);
    assign outputs[3439] = ~(layer0_outputs[6611]);
    assign outputs[3440] = ~((layer0_outputs[8881]) ^ (layer0_outputs[8979]));
    assign outputs[3441] = layer0_outputs[6776];
    assign outputs[3442] = (layer0_outputs[2827]) ^ (layer0_outputs[309]);
    assign outputs[3443] = ~((layer0_outputs[2578]) ^ (layer0_outputs[2506]));
    assign outputs[3444] = layer0_outputs[3736];
    assign outputs[3445] = ~((layer0_outputs[2012]) & (layer0_outputs[8803]));
    assign outputs[3446] = ~(layer0_outputs[6247]) | (layer0_outputs[4656]);
    assign outputs[3447] = layer0_outputs[8787];
    assign outputs[3448] = ~(layer0_outputs[8295]);
    assign outputs[3449] = ~(layer0_outputs[5683]);
    assign outputs[3450] = ~(layer0_outputs[8816]);
    assign outputs[3451] = (layer0_outputs[7360]) ^ (layer0_outputs[682]);
    assign outputs[3452] = (layer0_outputs[6943]) & ~(layer0_outputs[100]);
    assign outputs[3453] = layer0_outputs[6980];
    assign outputs[3454] = ~((layer0_outputs[4344]) ^ (layer0_outputs[8854]));
    assign outputs[3455] = layer0_outputs[7289];
    assign outputs[3456] = ~(layer0_outputs[6106]);
    assign outputs[3457] = ~(layer0_outputs[491]);
    assign outputs[3458] = ~(layer0_outputs[2931]);
    assign outputs[3459] = ~(layer0_outputs[7050]);
    assign outputs[3460] = layer0_outputs[5338];
    assign outputs[3461] = ~(layer0_outputs[1941]);
    assign outputs[3462] = layer0_outputs[664];
    assign outputs[3463] = ~(layer0_outputs[3216]) | (layer0_outputs[8653]);
    assign outputs[3464] = (layer0_outputs[9745]) & ~(layer0_outputs[764]);
    assign outputs[3465] = (layer0_outputs[6253]) ^ (layer0_outputs[676]);
    assign outputs[3466] = (layer0_outputs[6370]) & (layer0_outputs[8703]);
    assign outputs[3467] = ~(layer0_outputs[7546]) | (layer0_outputs[4296]);
    assign outputs[3468] = ~(layer0_outputs[8463]);
    assign outputs[3469] = layer0_outputs[3332];
    assign outputs[3470] = layer0_outputs[3985];
    assign outputs[3471] = ~((layer0_outputs[347]) ^ (layer0_outputs[1374]));
    assign outputs[3472] = ~((layer0_outputs[9539]) ^ (layer0_outputs[1820]));
    assign outputs[3473] = (layer0_outputs[5434]) ^ (layer0_outputs[2440]);
    assign outputs[3474] = (layer0_outputs[8196]) & (layer0_outputs[9710]);
    assign outputs[3475] = (layer0_outputs[3110]) | (layer0_outputs[4174]);
    assign outputs[3476] = ~((layer0_outputs[1443]) ^ (layer0_outputs[34]));
    assign outputs[3477] = layer0_outputs[5339];
    assign outputs[3478] = ~((layer0_outputs[3964]) | (layer0_outputs[1229]));
    assign outputs[3479] = (layer0_outputs[8277]) & ~(layer0_outputs[283]);
    assign outputs[3480] = (layer0_outputs[4614]) ^ (layer0_outputs[6207]);
    assign outputs[3481] = ~(layer0_outputs[3075]);
    assign outputs[3482] = ~(layer0_outputs[1032]);
    assign outputs[3483] = (layer0_outputs[9906]) & (layer0_outputs[5614]);
    assign outputs[3484] = (layer0_outputs[716]) & ~(layer0_outputs[3748]);
    assign outputs[3485] = ~(layer0_outputs[1238]) | (layer0_outputs[7783]);
    assign outputs[3486] = layer0_outputs[9735];
    assign outputs[3487] = ~(layer0_outputs[8052]) | (layer0_outputs[1793]);
    assign outputs[3488] = layer0_outputs[7755];
    assign outputs[3489] = layer0_outputs[1404];
    assign outputs[3490] = (layer0_outputs[417]) ^ (layer0_outputs[8588]);
    assign outputs[3491] = ~(layer0_outputs[4306]) | (layer0_outputs[7079]);
    assign outputs[3492] = layer0_outputs[7682];
    assign outputs[3493] = ~(layer0_outputs[1962]);
    assign outputs[3494] = layer0_outputs[1937];
    assign outputs[3495] = ~(layer0_outputs[1506]) | (layer0_outputs[8473]);
    assign outputs[3496] = ~(layer0_outputs[5969]);
    assign outputs[3497] = layer0_outputs[432];
    assign outputs[3498] = layer0_outputs[4134];
    assign outputs[3499] = ~((layer0_outputs[2996]) | (layer0_outputs[5740]));
    assign outputs[3500] = layer0_outputs[5812];
    assign outputs[3501] = layer0_outputs[396];
    assign outputs[3502] = ~(layer0_outputs[377]);
    assign outputs[3503] = layer0_outputs[6493];
    assign outputs[3504] = ~(layer0_outputs[8545]);
    assign outputs[3505] = layer0_outputs[10130];
    assign outputs[3506] = layer0_outputs[6171];
    assign outputs[3507] = layer0_outputs[3036];
    assign outputs[3508] = (layer0_outputs[3306]) & ~(layer0_outputs[7988]);
    assign outputs[3509] = (layer0_outputs[1374]) ^ (layer0_outputs[2452]);
    assign outputs[3510] = ~(layer0_outputs[163]);
    assign outputs[3511] = ~(layer0_outputs[4895]);
    assign outputs[3512] = ~((layer0_outputs[2512]) ^ (layer0_outputs[8778]));
    assign outputs[3513] = layer0_outputs[3965];
    assign outputs[3514] = ~(layer0_outputs[8173]);
    assign outputs[3515] = layer0_outputs[9581];
    assign outputs[3516] = (layer0_outputs[2733]) ^ (layer0_outputs[3370]);
    assign outputs[3517] = ~(layer0_outputs[7199]);
    assign outputs[3518] = (layer0_outputs[3468]) & (layer0_outputs[6871]);
    assign outputs[3519] = layer0_outputs[4487];
    assign outputs[3520] = ~((layer0_outputs[9159]) ^ (layer0_outputs[4033]));
    assign outputs[3521] = ~((layer0_outputs[26]) | (layer0_outputs[5551]));
    assign outputs[3522] = ~(layer0_outputs[3770]);
    assign outputs[3523] = (layer0_outputs[6598]) | (layer0_outputs[5016]);
    assign outputs[3524] = (layer0_outputs[1118]) & ~(layer0_outputs[5143]);
    assign outputs[3525] = ~(layer0_outputs[4318]);
    assign outputs[3526] = layer0_outputs[6280];
    assign outputs[3527] = ~(layer0_outputs[8695]);
    assign outputs[3528] = (layer0_outputs[5388]) ^ (layer0_outputs[896]);
    assign outputs[3529] = (layer0_outputs[6491]) & ~(layer0_outputs[8330]);
    assign outputs[3530] = layer0_outputs[1011];
    assign outputs[3531] = layer0_outputs[1602];
    assign outputs[3532] = (layer0_outputs[7282]) ^ (layer0_outputs[8748]);
    assign outputs[3533] = ~((layer0_outputs[8340]) | (layer0_outputs[8696]));
    assign outputs[3534] = ~((layer0_outputs[3716]) ^ (layer0_outputs[3786]));
    assign outputs[3535] = ~((layer0_outputs[112]) ^ (layer0_outputs[7491]));
    assign outputs[3536] = layer0_outputs[795];
    assign outputs[3537] = layer0_outputs[1289];
    assign outputs[3538] = layer0_outputs[2880];
    assign outputs[3539] = layer0_outputs[2633];
    assign outputs[3540] = (layer0_outputs[4156]) ^ (layer0_outputs[1940]);
    assign outputs[3541] = (layer0_outputs[8983]) & ~(layer0_outputs[1102]);
    assign outputs[3542] = ~(layer0_outputs[7239]);
    assign outputs[3543] = (layer0_outputs[7071]) & ~(layer0_outputs[2078]);
    assign outputs[3544] = (layer0_outputs[9826]) ^ (layer0_outputs[4108]);
    assign outputs[3545] = ~((layer0_outputs[5022]) ^ (layer0_outputs[8804]));
    assign outputs[3546] = ~(layer0_outputs[2692]);
    assign outputs[3547] = ~(layer0_outputs[1851]);
    assign outputs[3548] = ~(layer0_outputs[7041]);
    assign outputs[3549] = (layer0_outputs[3121]) & ~(layer0_outputs[7663]);
    assign outputs[3550] = ~(layer0_outputs[2229]);
    assign outputs[3551] = ~(layer0_outputs[5780]);
    assign outputs[3552] = (layer0_outputs[9831]) ^ (layer0_outputs[8140]);
    assign outputs[3553] = (layer0_outputs[9667]) ^ (layer0_outputs[225]);
    assign outputs[3554] = ~(layer0_outputs[7710]) | (layer0_outputs[2665]);
    assign outputs[3555] = (layer0_outputs[2589]) & ~(layer0_outputs[4185]);
    assign outputs[3556] = ~(layer0_outputs[1393]);
    assign outputs[3557] = (layer0_outputs[6406]) ^ (layer0_outputs[8696]);
    assign outputs[3558] = 1'b1;
    assign outputs[3559] = (layer0_outputs[10199]) & ~(layer0_outputs[3731]);
    assign outputs[3560] = (layer0_outputs[44]) ^ (layer0_outputs[7939]);
    assign outputs[3561] = ~(layer0_outputs[5142]);
    assign outputs[3562] = ~((layer0_outputs[6026]) ^ (layer0_outputs[5966]));
    assign outputs[3563] = ~(layer0_outputs[1509]);
    assign outputs[3564] = (layer0_outputs[9871]) & (layer0_outputs[9937]);
    assign outputs[3565] = layer0_outputs[1515];
    assign outputs[3566] = ~(layer0_outputs[2366]);
    assign outputs[3567] = layer0_outputs[8372];
    assign outputs[3568] = layer0_outputs[8303];
    assign outputs[3569] = ~((layer0_outputs[6358]) & (layer0_outputs[1899]));
    assign outputs[3570] = ~(layer0_outputs[1308]);
    assign outputs[3571] = ~(layer0_outputs[4758]);
    assign outputs[3572] = ~(layer0_outputs[8314]) | (layer0_outputs[2674]);
    assign outputs[3573] = layer0_outputs[2630];
    assign outputs[3574] = layer0_outputs[8058];
    assign outputs[3575] = (layer0_outputs[7889]) & ~(layer0_outputs[3603]);
    assign outputs[3576] = layer0_outputs[10150];
    assign outputs[3577] = (layer0_outputs[5276]) ^ (layer0_outputs[2669]);
    assign outputs[3578] = layer0_outputs[782];
    assign outputs[3579] = (layer0_outputs[7803]) & ~(layer0_outputs[5906]);
    assign outputs[3580] = ~(layer0_outputs[457]);
    assign outputs[3581] = (layer0_outputs[2758]) & (layer0_outputs[6950]);
    assign outputs[3582] = (layer0_outputs[7198]) & (layer0_outputs[4992]);
    assign outputs[3583] = ~((layer0_outputs[8526]) ^ (layer0_outputs[6706]));
    assign outputs[3584] = ~(layer0_outputs[5609]);
    assign outputs[3585] = ~(layer0_outputs[9071]);
    assign outputs[3586] = ~(layer0_outputs[7161]);
    assign outputs[3587] = layer0_outputs[7829];
    assign outputs[3588] = layer0_outputs[7657];
    assign outputs[3589] = ~(layer0_outputs[7875]);
    assign outputs[3590] = ~((layer0_outputs[4591]) & (layer0_outputs[6096]));
    assign outputs[3591] = ~(layer0_outputs[4081]) | (layer0_outputs[6627]);
    assign outputs[3592] = layer0_outputs[4596];
    assign outputs[3593] = layer0_outputs[4139];
    assign outputs[3594] = ~(layer0_outputs[2753]);
    assign outputs[3595] = ~((layer0_outputs[5003]) & (layer0_outputs[3538]));
    assign outputs[3596] = ~(layer0_outputs[1634]);
    assign outputs[3597] = (layer0_outputs[8955]) | (layer0_outputs[1224]);
    assign outputs[3598] = (layer0_outputs[7809]) & ~(layer0_outputs[7312]);
    assign outputs[3599] = ~(layer0_outputs[9558]);
    assign outputs[3600] = ~((layer0_outputs[7610]) ^ (layer0_outputs[5289]));
    assign outputs[3601] = ~(layer0_outputs[8429]) | (layer0_outputs[7129]);
    assign outputs[3602] = ~((layer0_outputs[8792]) | (layer0_outputs[8581]));
    assign outputs[3603] = ~((layer0_outputs[1065]) ^ (layer0_outputs[9321]));
    assign outputs[3604] = (layer0_outputs[3244]) ^ (layer0_outputs[4379]);
    assign outputs[3605] = ~((layer0_outputs[738]) ^ (layer0_outputs[1677]));
    assign outputs[3606] = (layer0_outputs[4479]) | (layer0_outputs[1197]);
    assign outputs[3607] = layer0_outputs[6168];
    assign outputs[3608] = (layer0_outputs[4938]) & ~(layer0_outputs[1961]);
    assign outputs[3609] = (layer0_outputs[3657]) ^ (layer0_outputs[6362]);
    assign outputs[3610] = ~(layer0_outputs[977]);
    assign outputs[3611] = layer0_outputs[5442];
    assign outputs[3612] = ~(layer0_outputs[3669]);
    assign outputs[3613] = layer0_outputs[3135];
    assign outputs[3614] = ~(layer0_outputs[6378]);
    assign outputs[3615] = ~(layer0_outputs[8613]);
    assign outputs[3616] = layer0_outputs[364];
    assign outputs[3617] = ~(layer0_outputs[8067]);
    assign outputs[3618] = ~(layer0_outputs[6068]);
    assign outputs[3619] = layer0_outputs[6180];
    assign outputs[3620] = (layer0_outputs[5686]) ^ (layer0_outputs[6514]);
    assign outputs[3621] = ~((layer0_outputs[3334]) ^ (layer0_outputs[1069]));
    assign outputs[3622] = layer0_outputs[1161];
    assign outputs[3623] = ~((layer0_outputs[1048]) | (layer0_outputs[3287]));
    assign outputs[3624] = ~(layer0_outputs[7511]);
    assign outputs[3625] = ~(layer0_outputs[10033]);
    assign outputs[3626] = (layer0_outputs[7673]) & (layer0_outputs[5536]);
    assign outputs[3627] = (layer0_outputs[7738]) ^ (layer0_outputs[3913]);
    assign outputs[3628] = ~(layer0_outputs[7193]);
    assign outputs[3629] = layer0_outputs[4215];
    assign outputs[3630] = (layer0_outputs[4091]) ^ (layer0_outputs[5315]);
    assign outputs[3631] = ~((layer0_outputs[4843]) & (layer0_outputs[6666]));
    assign outputs[3632] = ~(layer0_outputs[3951]);
    assign outputs[3633] = (layer0_outputs[7748]) & (layer0_outputs[6078]);
    assign outputs[3634] = ~(layer0_outputs[4286]);
    assign outputs[3635] = layer0_outputs[6655];
    assign outputs[3636] = layer0_outputs[6127];
    assign outputs[3637] = ~(layer0_outputs[7253]);
    assign outputs[3638] = layer0_outputs[1894];
    assign outputs[3639] = (layer0_outputs[4497]) & ~(layer0_outputs[1400]);
    assign outputs[3640] = (layer0_outputs[3888]) & (layer0_outputs[7603]);
    assign outputs[3641] = layer0_outputs[743];
    assign outputs[3642] = ~(layer0_outputs[1029]) | (layer0_outputs[4624]);
    assign outputs[3643] = (layer0_outputs[3776]) | (layer0_outputs[7468]);
    assign outputs[3644] = (layer0_outputs[4163]) ^ (layer0_outputs[8225]);
    assign outputs[3645] = layer0_outputs[6388];
    assign outputs[3646] = layer0_outputs[9927];
    assign outputs[3647] = ~(layer0_outputs[429]);
    assign outputs[3648] = layer0_outputs[3729];
    assign outputs[3649] = ~((layer0_outputs[8782]) ^ (layer0_outputs[901]));
    assign outputs[3650] = layer0_outputs[6693];
    assign outputs[3651] = (layer0_outputs[6819]) ^ (layer0_outputs[6726]);
    assign outputs[3652] = (layer0_outputs[6093]) & (layer0_outputs[8479]);
    assign outputs[3653] = ~((layer0_outputs[3999]) ^ (layer0_outputs[1250]));
    assign outputs[3654] = (layer0_outputs[5615]) & (layer0_outputs[2597]);
    assign outputs[3655] = layer0_outputs[2722];
    assign outputs[3656] = layer0_outputs[1919];
    assign outputs[3657] = ~((layer0_outputs[7936]) ^ (layer0_outputs[4557]));
    assign outputs[3658] = (layer0_outputs[9808]) & ~(layer0_outputs[2587]);
    assign outputs[3659] = ~(layer0_outputs[6763]);
    assign outputs[3660] = ~((layer0_outputs[773]) ^ (layer0_outputs[6483]));
    assign outputs[3661] = layer0_outputs[1590];
    assign outputs[3662] = ~(layer0_outputs[899]) | (layer0_outputs[5972]);
    assign outputs[3663] = (layer0_outputs[3774]) ^ (layer0_outputs[4534]);
    assign outputs[3664] = (layer0_outputs[8622]) & ~(layer0_outputs[6612]);
    assign outputs[3665] = layer0_outputs[6594];
    assign outputs[3666] = ~((layer0_outputs[8274]) ^ (layer0_outputs[5163]));
    assign outputs[3667] = ~((layer0_outputs[578]) & (layer0_outputs[4054]));
    assign outputs[3668] = ~(layer0_outputs[5181]);
    assign outputs[3669] = layer0_outputs[8062];
    assign outputs[3670] = ~(layer0_outputs[8239]);
    assign outputs[3671] = (layer0_outputs[4494]) & (layer0_outputs[9446]);
    assign outputs[3672] = ~(layer0_outputs[6442]);
    assign outputs[3673] = ~(layer0_outputs[10220]);
    assign outputs[3674] = ~((layer0_outputs[6947]) ^ (layer0_outputs[7566]));
    assign outputs[3675] = ~((layer0_outputs[5635]) | (layer0_outputs[10093]));
    assign outputs[3676] = (layer0_outputs[8474]) & ~(layer0_outputs[1737]);
    assign outputs[3677] = (layer0_outputs[6930]) & ~(layer0_outputs[9753]);
    assign outputs[3678] = (layer0_outputs[2919]) & ~(layer0_outputs[3282]);
    assign outputs[3679] = ~((layer0_outputs[1061]) & (layer0_outputs[1253]));
    assign outputs[3680] = ~(layer0_outputs[4025]);
    assign outputs[3681] = ~(layer0_outputs[4630]);
    assign outputs[3682] = ~(layer0_outputs[9998]) | (layer0_outputs[149]);
    assign outputs[3683] = layer0_outputs[5856];
    assign outputs[3684] = ~(layer0_outputs[8445]);
    assign outputs[3685] = (layer0_outputs[4198]) ^ (layer0_outputs[4207]);
    assign outputs[3686] = layer0_outputs[9405];
    assign outputs[3687] = (layer0_outputs[894]) & ~(layer0_outputs[623]);
    assign outputs[3688] = ~(layer0_outputs[9707]);
    assign outputs[3689] = ~((layer0_outputs[1097]) ^ (layer0_outputs[4160]));
    assign outputs[3690] = ~((layer0_outputs[1031]) ^ (layer0_outputs[4733]));
    assign outputs[3691] = (layer0_outputs[3187]) ^ (layer0_outputs[1229]);
    assign outputs[3692] = ~(layer0_outputs[4741]) | (layer0_outputs[8861]);
    assign outputs[3693] = layer0_outputs[7625];
    assign outputs[3694] = layer0_outputs[6552];
    assign outputs[3695] = ~(layer0_outputs[3262]) | (layer0_outputs[4475]);
    assign outputs[3696] = layer0_outputs[8327];
    assign outputs[3697] = (layer0_outputs[6276]) ^ (layer0_outputs[7095]);
    assign outputs[3698] = ~(layer0_outputs[7662]);
    assign outputs[3699] = (layer0_outputs[7745]) & ~(layer0_outputs[6351]);
    assign outputs[3700] = ~((layer0_outputs[3433]) ^ (layer0_outputs[8552]));
    assign outputs[3701] = (layer0_outputs[9001]) & ~(layer0_outputs[7016]);
    assign outputs[3702] = layer0_outputs[6753];
    assign outputs[3703] = ~(layer0_outputs[9042]);
    assign outputs[3704] = layer0_outputs[9239];
    assign outputs[3705] = ~((layer0_outputs[9489]) ^ (layer0_outputs[8624]));
    assign outputs[3706] = ~(layer0_outputs[5203]);
    assign outputs[3707] = ~(layer0_outputs[2474]);
    assign outputs[3708] = layer0_outputs[9113];
    assign outputs[3709] = (layer0_outputs[4653]) ^ (layer0_outputs[559]);
    assign outputs[3710] = ~((layer0_outputs[4351]) ^ (layer0_outputs[1543]));
    assign outputs[3711] = (layer0_outputs[1340]) & ~(layer0_outputs[6423]);
    assign outputs[3712] = ~((layer0_outputs[4994]) ^ (layer0_outputs[1123]));
    assign outputs[3713] = ~(layer0_outputs[8394]);
    assign outputs[3714] = ~(layer0_outputs[1872]);
    assign outputs[3715] = layer0_outputs[2244];
    assign outputs[3716] = ~(layer0_outputs[5804]);
    assign outputs[3717] = ~(layer0_outputs[7180]) | (layer0_outputs[4416]);
    assign outputs[3718] = layer0_outputs[8347];
    assign outputs[3719] = ~(layer0_outputs[5467]);
    assign outputs[3720] = ~(layer0_outputs[4779]);
    assign outputs[3721] = layer0_outputs[5929];
    assign outputs[3722] = layer0_outputs[8737];
    assign outputs[3723] = ~(layer0_outputs[4002]);
    assign outputs[3724] = (layer0_outputs[5030]) ^ (layer0_outputs[4086]);
    assign outputs[3725] = ~(layer0_outputs[6284]);
    assign outputs[3726] = ~(layer0_outputs[480]);
    assign outputs[3727] = layer0_outputs[27];
    assign outputs[3728] = layer0_outputs[1282];
    assign outputs[3729] = layer0_outputs[1581];
    assign outputs[3730] = (layer0_outputs[902]) & (layer0_outputs[8841]);
    assign outputs[3731] = ~(layer0_outputs[7023]);
    assign outputs[3732] = (layer0_outputs[5515]) ^ (layer0_outputs[7420]);
    assign outputs[3733] = layer0_outputs[6696];
    assign outputs[3734] = (layer0_outputs[6385]) & ~(layer0_outputs[38]);
    assign outputs[3735] = ~(layer0_outputs[9129]) | (layer0_outputs[536]);
    assign outputs[3736] = (layer0_outputs[8667]) & ~(layer0_outputs[3608]);
    assign outputs[3737] = layer0_outputs[748];
    assign outputs[3738] = (layer0_outputs[10133]) & ~(layer0_outputs[9271]);
    assign outputs[3739] = layer0_outputs[3410];
    assign outputs[3740] = (layer0_outputs[7972]) & ~(layer0_outputs[2088]);
    assign outputs[3741] = layer0_outputs[6055];
    assign outputs[3742] = layer0_outputs[6603];
    assign outputs[3743] = ~((layer0_outputs[6304]) ^ (layer0_outputs[8894]));
    assign outputs[3744] = layer0_outputs[9618];
    assign outputs[3745] = layer0_outputs[5711];
    assign outputs[3746] = ~(layer0_outputs[84]);
    assign outputs[3747] = ~(layer0_outputs[4330]);
    assign outputs[3748] = (layer0_outputs[6419]) ^ (layer0_outputs[1985]);
    assign outputs[3749] = ~((layer0_outputs[9943]) | (layer0_outputs[1338]));
    assign outputs[3750] = layer0_outputs[9578];
    assign outputs[3751] = ~((layer0_outputs[2010]) ^ (layer0_outputs[8320]));
    assign outputs[3752] = ~(layer0_outputs[5486]);
    assign outputs[3753] = (layer0_outputs[5080]) & (layer0_outputs[3544]);
    assign outputs[3754] = ~((layer0_outputs[7890]) & (layer0_outputs[5034]));
    assign outputs[3755] = ~((layer0_outputs[7479]) ^ (layer0_outputs[4528]));
    assign outputs[3756] = ~(layer0_outputs[2658]);
    assign outputs[3757] = (layer0_outputs[5435]) ^ (layer0_outputs[2725]);
    assign outputs[3758] = layer0_outputs[7085];
    assign outputs[3759] = layer0_outputs[9469];
    assign outputs[3760] = ~((layer0_outputs[4748]) ^ (layer0_outputs[5297]));
    assign outputs[3761] = (layer0_outputs[5233]) ^ (layer0_outputs[249]);
    assign outputs[3762] = layer0_outputs[1456];
    assign outputs[3763] = (layer0_outputs[9335]) & ~(layer0_outputs[5463]);
    assign outputs[3764] = layer0_outputs[9006];
    assign outputs[3765] = (layer0_outputs[5873]) ^ (layer0_outputs[6741]);
    assign outputs[3766] = layer0_outputs[10088];
    assign outputs[3767] = layer0_outputs[2093];
    assign outputs[3768] = ~(layer0_outputs[3514]) | (layer0_outputs[7668]);
    assign outputs[3769] = ~((layer0_outputs[8236]) ^ (layer0_outputs[4892]));
    assign outputs[3770] = ~((layer0_outputs[3386]) & (layer0_outputs[2321]));
    assign outputs[3771] = ~(layer0_outputs[7202]);
    assign outputs[3772] = (layer0_outputs[5415]) | (layer0_outputs[62]);
    assign outputs[3773] = ~(layer0_outputs[1416]) | (layer0_outputs[2645]);
    assign outputs[3774] = (layer0_outputs[413]) & (layer0_outputs[3099]);
    assign outputs[3775] = (layer0_outputs[632]) & (layer0_outputs[7603]);
    assign outputs[3776] = (layer0_outputs[8483]) ^ (layer0_outputs[7955]);
    assign outputs[3777] = ~((layer0_outputs[3396]) ^ (layer0_outputs[1896]));
    assign outputs[3778] = (layer0_outputs[3780]) & (layer0_outputs[9330]);
    assign outputs[3779] = ~((layer0_outputs[8806]) ^ (layer0_outputs[5583]));
    assign outputs[3780] = ~((layer0_outputs[8764]) ^ (layer0_outputs[9739]));
    assign outputs[3781] = (layer0_outputs[8027]) ^ (layer0_outputs[7071]);
    assign outputs[3782] = ~((layer0_outputs[7299]) & (layer0_outputs[2564]));
    assign outputs[3783] = (layer0_outputs[5992]) ^ (layer0_outputs[8116]);
    assign outputs[3784] = (layer0_outputs[1287]) & ~(layer0_outputs[1643]);
    assign outputs[3785] = layer0_outputs[4353];
    assign outputs[3786] = ~(layer0_outputs[8368]);
    assign outputs[3787] = ~(layer0_outputs[6809]);
    assign outputs[3788] = ~((layer0_outputs[6124]) | (layer0_outputs[5309]));
    assign outputs[3789] = (layer0_outputs[3861]) ^ (layer0_outputs[1467]);
    assign outputs[3790] = (layer0_outputs[1866]) & ~(layer0_outputs[9809]);
    assign outputs[3791] = ~((layer0_outputs[4781]) & (layer0_outputs[9964]));
    assign outputs[3792] = (layer0_outputs[9592]) & ~(layer0_outputs[9225]);
    assign outputs[3793] = (layer0_outputs[295]) & (layer0_outputs[8348]);
    assign outputs[3794] = ~((layer0_outputs[3208]) | (layer0_outputs[5216]));
    assign outputs[3795] = layer0_outputs[4999];
    assign outputs[3796] = (layer0_outputs[6015]) & ~(layer0_outputs[3313]);
    assign outputs[3797] = (layer0_outputs[4153]) | (layer0_outputs[1724]);
    assign outputs[3798] = layer0_outputs[6918];
    assign outputs[3799] = (layer0_outputs[5391]) & ~(layer0_outputs[3418]);
    assign outputs[3800] = ~(layer0_outputs[1336]);
    assign outputs[3801] = ~((layer0_outputs[3304]) | (layer0_outputs[6888]));
    assign outputs[3802] = layer0_outputs[7570];
    assign outputs[3803] = layer0_outputs[934];
    assign outputs[3804] = ~(layer0_outputs[8549]);
    assign outputs[3805] = ~((layer0_outputs[5746]) ^ (layer0_outputs[4508]));
    assign outputs[3806] = ~(layer0_outputs[2468]);
    assign outputs[3807] = (layer0_outputs[10121]) & ~(layer0_outputs[8616]);
    assign outputs[3808] = layer0_outputs[6969];
    assign outputs[3809] = (layer0_outputs[9538]) ^ (layer0_outputs[7670]);
    assign outputs[3810] = layer0_outputs[6875];
    assign outputs[3811] = ~((layer0_outputs[1796]) ^ (layer0_outputs[7419]));
    assign outputs[3812] = layer0_outputs[6883];
    assign outputs[3813] = ~((layer0_outputs[542]) ^ (layer0_outputs[2741]));
    assign outputs[3814] = (layer0_outputs[5622]) & ~(layer0_outputs[1513]);
    assign outputs[3815] = (layer0_outputs[3470]) & (layer0_outputs[5785]);
    assign outputs[3816] = ~(layer0_outputs[7984]);
    assign outputs[3817] = (layer0_outputs[6080]) & ~(layer0_outputs[5591]);
    assign outputs[3818] = ~(layer0_outputs[7746]);
    assign outputs[3819] = ~((layer0_outputs[6458]) ^ (layer0_outputs[3391]));
    assign outputs[3820] = layer0_outputs[785];
    assign outputs[3821] = (layer0_outputs[4840]) ^ (layer0_outputs[3550]);
    assign outputs[3822] = layer0_outputs[224];
    assign outputs[3823] = ~(layer0_outputs[771]);
    assign outputs[3824] = layer0_outputs[7334];
    assign outputs[3825] = ~(layer0_outputs[8034]);
    assign outputs[3826] = ~(layer0_outputs[1625]);
    assign outputs[3827] = ~(layer0_outputs[5871]);
    assign outputs[3828] = layer0_outputs[9395];
    assign outputs[3829] = layer0_outputs[5040];
    assign outputs[3830] = (layer0_outputs[5775]) & (layer0_outputs[8081]);
    assign outputs[3831] = layer0_outputs[6767];
    assign outputs[3832] = ~(layer0_outputs[8305]);
    assign outputs[3833] = ~(layer0_outputs[8686]) | (layer0_outputs[2811]);
    assign outputs[3834] = ~((layer0_outputs[6362]) ^ (layer0_outputs[6419]));
    assign outputs[3835] = ~((layer0_outputs[9582]) ^ (layer0_outputs[8471]));
    assign outputs[3836] = layer0_outputs[9786];
    assign outputs[3837] = ~((layer0_outputs[1867]) ^ (layer0_outputs[4699]));
    assign outputs[3838] = ~((layer0_outputs[1794]) ^ (layer0_outputs[4638]));
    assign outputs[3839] = layer0_outputs[715];
    assign outputs[3840] = ~(layer0_outputs[3328]);
    assign outputs[3841] = ~(layer0_outputs[8927]);
    assign outputs[3842] = layer0_outputs[3067];
    assign outputs[3843] = ~((layer0_outputs[6773]) | (layer0_outputs[551]));
    assign outputs[3844] = ~(layer0_outputs[2148]) | (layer0_outputs[5361]);
    assign outputs[3845] = (layer0_outputs[4875]) | (layer0_outputs[9023]);
    assign outputs[3846] = layer0_outputs[8505];
    assign outputs[3847] = ~(layer0_outputs[9010]);
    assign outputs[3848] = ~((layer0_outputs[8171]) & (layer0_outputs[8535]));
    assign outputs[3849] = ~(layer0_outputs[1635]);
    assign outputs[3850] = (layer0_outputs[5422]) ^ (layer0_outputs[3762]);
    assign outputs[3851] = layer0_outputs[8735];
    assign outputs[3852] = ~((layer0_outputs[5097]) ^ (layer0_outputs[7655]));
    assign outputs[3853] = ~((layer0_outputs[883]) | (layer0_outputs[713]));
    assign outputs[3854] = layer0_outputs[933];
    assign outputs[3855] = ~(layer0_outputs[2700]);
    assign outputs[3856] = layer0_outputs[8341];
    assign outputs[3857] = layer0_outputs[7386];
    assign outputs[3858] = ~(layer0_outputs[3901]);
    assign outputs[3859] = ~(layer0_outputs[4858]);
    assign outputs[3860] = ~((layer0_outputs[547]) ^ (layer0_outputs[4605]));
    assign outputs[3861] = (layer0_outputs[8385]) ^ (layer0_outputs[10052]);
    assign outputs[3862] = layer0_outputs[8012];
    assign outputs[3863] = layer0_outputs[9221];
    assign outputs[3864] = ~(layer0_outputs[503]);
    assign outputs[3865] = (layer0_outputs[2268]) ^ (layer0_outputs[7460]);
    assign outputs[3866] = (layer0_outputs[7156]) ^ (layer0_outputs[5672]);
    assign outputs[3867] = (layer0_outputs[2182]) | (layer0_outputs[11]);
    assign outputs[3868] = ~((layer0_outputs[8516]) | (layer0_outputs[1173]));
    assign outputs[3869] = ~(layer0_outputs[634]);
    assign outputs[3870] = layer0_outputs[88];
    assign outputs[3871] = (layer0_outputs[8168]) ^ (layer0_outputs[7708]);
    assign outputs[3872] = (layer0_outputs[7154]) | (layer0_outputs[8969]);
    assign outputs[3873] = (layer0_outputs[7352]) | (layer0_outputs[8986]);
    assign outputs[3874] = layer0_outputs[5374];
    assign outputs[3875] = ~(layer0_outputs[3834]);
    assign outputs[3876] = ~(layer0_outputs[6710]);
    assign outputs[3877] = (layer0_outputs[5214]) & ~(layer0_outputs[5556]);
    assign outputs[3878] = layer0_outputs[7885];
    assign outputs[3879] = ~((layer0_outputs[4685]) ^ (layer0_outputs[5218]));
    assign outputs[3880] = ~((layer0_outputs[2334]) | (layer0_outputs[4275]));
    assign outputs[3881] = ~(layer0_outputs[8788]);
    assign outputs[3882] = layer0_outputs[4595];
    assign outputs[3883] = ~(layer0_outputs[8106]) | (layer0_outputs[2405]);
    assign outputs[3884] = ~(layer0_outputs[3635]);
    assign outputs[3885] = ~(layer0_outputs[3581]);
    assign outputs[3886] = ~((layer0_outputs[9591]) ^ (layer0_outputs[1343]));
    assign outputs[3887] = ~(layer0_outputs[9260]) | (layer0_outputs[4684]);
    assign outputs[3888] = layer0_outputs[908];
    assign outputs[3889] = layer0_outputs[4890];
    assign outputs[3890] = ~(layer0_outputs[9738]);
    assign outputs[3891] = layer0_outputs[9978];
    assign outputs[3892] = ~(layer0_outputs[3894]);
    assign outputs[3893] = ~(layer0_outputs[6109]) | (layer0_outputs[3147]);
    assign outputs[3894] = ~(layer0_outputs[9706]);
    assign outputs[3895] = ~(layer0_outputs[5959]);
    assign outputs[3896] = (layer0_outputs[4308]) ^ (layer0_outputs[8660]);
    assign outputs[3897] = layer0_outputs[7637];
    assign outputs[3898] = (layer0_outputs[4969]) ^ (layer0_outputs[5198]);
    assign outputs[3899] = (layer0_outputs[507]) & ~(layer0_outputs[4794]);
    assign outputs[3900] = layer0_outputs[6744];
    assign outputs[3901] = (layer0_outputs[5926]) & ~(layer0_outputs[7996]);
    assign outputs[3902] = layer0_outputs[4460];
    assign outputs[3903] = (layer0_outputs[3692]) ^ (layer0_outputs[1907]);
    assign outputs[3904] = (layer0_outputs[6238]) & ~(layer0_outputs[7771]);
    assign outputs[3905] = ~(layer0_outputs[10073]);
    assign outputs[3906] = (layer0_outputs[6877]) ^ (layer0_outputs[9616]);
    assign outputs[3907] = (layer0_outputs[2361]) ^ (layer0_outputs[9526]);
    assign outputs[3908] = (layer0_outputs[345]) | (layer0_outputs[1202]);
    assign outputs[3909] = layer0_outputs[5523];
    assign outputs[3910] = (layer0_outputs[7227]) & ~(layer0_outputs[8699]);
    assign outputs[3911] = (layer0_outputs[8776]) ^ (layer0_outputs[6505]);
    assign outputs[3912] = ~(layer0_outputs[8318]);
    assign outputs[3913] = layer0_outputs[2913];
    assign outputs[3914] = layer0_outputs[107];
    assign outputs[3915] = (layer0_outputs[9911]) ^ (layer0_outputs[6458]);
    assign outputs[3916] = layer0_outputs[1799];
    assign outputs[3917] = ~(layer0_outputs[8210]);
    assign outputs[3918] = layer0_outputs[374];
    assign outputs[3919] = (layer0_outputs[6379]) ^ (layer0_outputs[7256]);
    assign outputs[3920] = ~((layer0_outputs[5483]) ^ (layer0_outputs[6915]));
    assign outputs[3921] = (layer0_outputs[444]) ^ (layer0_outputs[5177]);
    assign outputs[3922] = ~((layer0_outputs[7358]) ^ (layer0_outputs[2791]));
    assign outputs[3923] = (layer0_outputs[199]) & ~(layer0_outputs[7391]);
    assign outputs[3924] = (layer0_outputs[7775]) & ~(layer0_outputs[3407]);
    assign outputs[3925] = (layer0_outputs[835]) ^ (layer0_outputs[9513]);
    assign outputs[3926] = ~(layer0_outputs[9828]);
    assign outputs[3927] = (layer0_outputs[5484]) & ~(layer0_outputs[3777]);
    assign outputs[3928] = ~(layer0_outputs[1834]);
    assign outputs[3929] = layer0_outputs[3918];
    assign outputs[3930] = ~(layer0_outputs[5792]);
    assign outputs[3931] = (layer0_outputs[3990]) ^ (layer0_outputs[5114]);
    assign outputs[3932] = layer0_outputs[7896];
    assign outputs[3933] = ~(layer0_outputs[633]);
    assign outputs[3934] = (layer0_outputs[5016]) & (layer0_outputs[6510]);
    assign outputs[3935] = layer0_outputs[7342];
    assign outputs[3936] = (layer0_outputs[1774]) & (layer0_outputs[4186]);
    assign outputs[3937] = layer0_outputs[6657];
    assign outputs[3938] = ~(layer0_outputs[9336]);
    assign outputs[3939] = (layer0_outputs[214]) & (layer0_outputs[7174]);
    assign outputs[3940] = ~(layer0_outputs[1728]) | (layer0_outputs[530]);
    assign outputs[3941] = layer0_outputs[4290];
    assign outputs[3942] = (layer0_outputs[9771]) ^ (layer0_outputs[3365]);
    assign outputs[3943] = ~(layer0_outputs[4502]);
    assign outputs[3944] = ~(layer0_outputs[2629]);
    assign outputs[3945] = ~((layer0_outputs[5628]) ^ (layer0_outputs[9592]));
    assign outputs[3946] = (layer0_outputs[5010]) & ~(layer0_outputs[8396]);
    assign outputs[3947] = (layer0_outputs[415]) ^ (layer0_outputs[8235]);
    assign outputs[3948] = ~(layer0_outputs[5447]) | (layer0_outputs[75]);
    assign outputs[3949] = ~(layer0_outputs[12]) | (layer0_outputs[7876]);
    assign outputs[3950] = ~(layer0_outputs[2269]);
    assign outputs[3951] = layer0_outputs[5980];
    assign outputs[3952] = (layer0_outputs[702]) ^ (layer0_outputs[1932]);
    assign outputs[3953] = ~(layer0_outputs[4098]);
    assign outputs[3954] = layer0_outputs[5595];
    assign outputs[3955] = (layer0_outputs[1279]) | (layer0_outputs[1399]);
    assign outputs[3956] = ~(layer0_outputs[297]);
    assign outputs[3957] = ~(layer0_outputs[4260]);
    assign outputs[3958] = (layer0_outputs[4237]) & (layer0_outputs[4168]);
    assign outputs[3959] = layer0_outputs[718];
    assign outputs[3960] = layer0_outputs[2409];
    assign outputs[3961] = ~(layer0_outputs[9635]);
    assign outputs[3962] = ~(layer0_outputs[7554]);
    assign outputs[3963] = ~((layer0_outputs[7374]) | (layer0_outputs[7295]));
    assign outputs[3964] = ~(layer0_outputs[10041]);
    assign outputs[3965] = layer0_outputs[3339];
    assign outputs[3966] = (layer0_outputs[8188]) & ~(layer0_outputs[6050]);
    assign outputs[3967] = (layer0_outputs[5662]) ^ (layer0_outputs[5582]);
    assign outputs[3968] = layer0_outputs[7623];
    assign outputs[3969] = ~(layer0_outputs[6492]);
    assign outputs[3970] = ~(layer0_outputs[4944]);
    assign outputs[3971] = ~(layer0_outputs[4642]);
    assign outputs[3972] = ~(layer0_outputs[2467]);
    assign outputs[3973] = layer0_outputs[4725];
    assign outputs[3974] = (layer0_outputs[865]) & ~(layer0_outputs[883]);
    assign outputs[3975] = layer0_outputs[10171];
    assign outputs[3976] = (layer0_outputs[3860]) & (layer0_outputs[9178]);
    assign outputs[3977] = layer0_outputs[2115];
    assign outputs[3978] = (layer0_outputs[4668]) ^ (layer0_outputs[7493]);
    assign outputs[3979] = ~((layer0_outputs[896]) ^ (layer0_outputs[3230]));
    assign outputs[3980] = (layer0_outputs[8694]) ^ (layer0_outputs[10007]);
    assign outputs[3981] = (layer0_outputs[6898]) & (layer0_outputs[4409]);
    assign outputs[3982] = ~((layer0_outputs[407]) ^ (layer0_outputs[6370]));
    assign outputs[3983] = (layer0_outputs[8337]) & (layer0_outputs[3024]);
    assign outputs[3984] = (layer0_outputs[4822]) ^ (layer0_outputs[4831]);
    assign outputs[3985] = (layer0_outputs[3223]) & ~(layer0_outputs[7879]);
    assign outputs[3986] = (layer0_outputs[5658]) ^ (layer0_outputs[8186]);
    assign outputs[3987] = layer0_outputs[1887];
    assign outputs[3988] = layer0_outputs[8898];
    assign outputs[3989] = ~(layer0_outputs[2491]);
    assign outputs[3990] = ~(layer0_outputs[3778]);
    assign outputs[3991] = ~(layer0_outputs[594]);
    assign outputs[3992] = (layer0_outputs[8666]) & ~(layer0_outputs[10058]);
    assign outputs[3993] = ~(layer0_outputs[9829]);
    assign outputs[3994] = (layer0_outputs[5845]) | (layer0_outputs[3512]);
    assign outputs[3995] = ~(layer0_outputs[8635]);
    assign outputs[3996] = layer0_outputs[9973];
    assign outputs[3997] = ~((layer0_outputs[8186]) | (layer0_outputs[141]));
    assign outputs[3998] = ~((layer0_outputs[8344]) | (layer0_outputs[9373]));
    assign outputs[3999] = (layer0_outputs[7987]) & ~(layer0_outputs[5639]);
    assign outputs[4000] = layer0_outputs[1939];
    assign outputs[4001] = (layer0_outputs[1398]) & ~(layer0_outputs[1837]);
    assign outputs[4002] = (layer0_outputs[414]) ^ (layer0_outputs[8011]);
    assign outputs[4003] = ~((layer0_outputs[2512]) | (layer0_outputs[1383]));
    assign outputs[4004] = (layer0_outputs[1382]) | (layer0_outputs[9087]);
    assign outputs[4005] = layer0_outputs[5162];
    assign outputs[4006] = ~((layer0_outputs[8953]) | (layer0_outputs[8551]));
    assign outputs[4007] = ~(layer0_outputs[1547]);
    assign outputs[4008] = (layer0_outputs[4504]) & ~(layer0_outputs[554]);
    assign outputs[4009] = ~(layer0_outputs[6020]);
    assign outputs[4010] = (layer0_outputs[6906]) & ~(layer0_outputs[751]);
    assign outputs[4011] = layer0_outputs[8287];
    assign outputs[4012] = layer0_outputs[7314];
    assign outputs[4013] = (layer0_outputs[6229]) ^ (layer0_outputs[5303]);
    assign outputs[4014] = (layer0_outputs[2626]) & ~(layer0_outputs[8478]);
    assign outputs[4015] = ~((layer0_outputs[5788]) ^ (layer0_outputs[1616]));
    assign outputs[4016] = ~(layer0_outputs[9040]);
    assign outputs[4017] = layer0_outputs[8053];
    assign outputs[4018] = ~((layer0_outputs[9824]) ^ (layer0_outputs[3402]));
    assign outputs[4019] = ~(layer0_outputs[60]);
    assign outputs[4020] = ~(layer0_outputs[523]);
    assign outputs[4021] = layer0_outputs[3665];
    assign outputs[4022] = ~(layer0_outputs[4688]);
    assign outputs[4023] = (layer0_outputs[1805]) ^ (layer0_outputs[5690]);
    assign outputs[4024] = ~(layer0_outputs[4540]);
    assign outputs[4025] = ~(layer0_outputs[5245]);
    assign outputs[4026] = layer0_outputs[5546];
    assign outputs[4027] = ~((layer0_outputs[4746]) | (layer0_outputs[5413]));
    assign outputs[4028] = layer0_outputs[7162];
    assign outputs[4029] = layer0_outputs[8117];
    assign outputs[4030] = layer0_outputs[2719];
    assign outputs[4031] = ~(layer0_outputs[8199]) | (layer0_outputs[10054]);
    assign outputs[4032] = layer0_outputs[3099];
    assign outputs[4033] = layer0_outputs[5418];
    assign outputs[4034] = ~((layer0_outputs[3085]) ^ (layer0_outputs[5021]));
    assign outputs[4035] = ~(layer0_outputs[6209]) | (layer0_outputs[1945]);
    assign outputs[4036] = (layer0_outputs[5841]) | (layer0_outputs[7479]);
    assign outputs[4037] = layer0_outputs[187];
    assign outputs[4038] = layer0_outputs[7294];
    assign outputs[4039] = layer0_outputs[2497];
    assign outputs[4040] = ~(layer0_outputs[9119]);
    assign outputs[4041] = ~(layer0_outputs[9885]);
    assign outputs[4042] = ~((layer0_outputs[4372]) & (layer0_outputs[8107]));
    assign outputs[4043] = layer0_outputs[8687];
    assign outputs[4044] = (layer0_outputs[10143]) ^ (layer0_outputs[9367]);
    assign outputs[4045] = ~((layer0_outputs[1110]) ^ (layer0_outputs[4295]));
    assign outputs[4046] = (layer0_outputs[8807]) ^ (layer0_outputs[6235]);
    assign outputs[4047] = layer0_outputs[9379];
    assign outputs[4048] = ~(layer0_outputs[4500]);
    assign outputs[4049] = layer0_outputs[2285];
    assign outputs[4050] = (layer0_outputs[1577]) ^ (layer0_outputs[2252]);
    assign outputs[4051] = ~(layer0_outputs[752]);
    assign outputs[4052] = (layer0_outputs[7072]) & ~(layer0_outputs[2308]);
    assign outputs[4053] = ~(layer0_outputs[4219]);
    assign outputs[4054] = layer0_outputs[7352];
    assign outputs[4055] = (layer0_outputs[7763]) | (layer0_outputs[8538]);
    assign outputs[4056] = layer0_outputs[4616];
    assign outputs[4057] = layer0_outputs[5160];
    assign outputs[4058] = ~(layer0_outputs[3171]);
    assign outputs[4059] = ~((layer0_outputs[8172]) ^ (layer0_outputs[8981]));
    assign outputs[4060] = (layer0_outputs[2746]) & (layer0_outputs[10205]);
    assign outputs[4061] = ~(layer0_outputs[3707]);
    assign outputs[4062] = ~(layer0_outputs[1634]);
    assign outputs[4063] = layer0_outputs[9059];
    assign outputs[4064] = ~(layer0_outputs[1506]);
    assign outputs[4065] = ~((layer0_outputs[7737]) ^ (layer0_outputs[2454]));
    assign outputs[4066] = layer0_outputs[4073];
    assign outputs[4067] = (layer0_outputs[7415]) & (layer0_outputs[914]);
    assign outputs[4068] = (layer0_outputs[24]) & (layer0_outputs[8771]);
    assign outputs[4069] = ~((layer0_outputs[151]) ^ (layer0_outputs[4482]));
    assign outputs[4070] = ~(layer0_outputs[3963]) | (layer0_outputs[9420]);
    assign outputs[4071] = ~(layer0_outputs[9611]);
    assign outputs[4072] = layer0_outputs[1534];
    assign outputs[4073] = (layer0_outputs[7229]) ^ (layer0_outputs[291]);
    assign outputs[4074] = (layer0_outputs[6368]) & (layer0_outputs[5421]);
    assign outputs[4075] = layer0_outputs[2436];
    assign outputs[4076] = ~(layer0_outputs[2336]);
    assign outputs[4077] = layer0_outputs[9609];
    assign outputs[4078] = (layer0_outputs[6806]) ^ (layer0_outputs[8929]);
    assign outputs[4079] = layer0_outputs[8498];
    assign outputs[4080] = (layer0_outputs[1759]) ^ (layer0_outputs[4014]);
    assign outputs[4081] = layer0_outputs[6723];
    assign outputs[4082] = ~(layer0_outputs[1192]) | (layer0_outputs[674]);
    assign outputs[4083] = ~(layer0_outputs[1814]);
    assign outputs[4084] = (layer0_outputs[2964]) & ~(layer0_outputs[1152]);
    assign outputs[4085] = ~(layer0_outputs[5349]);
    assign outputs[4086] = (layer0_outputs[5265]) & ~(layer0_outputs[6870]);
    assign outputs[4087] = (layer0_outputs[6697]) ^ (layer0_outputs[2782]);
    assign outputs[4088] = ~(layer0_outputs[4425]) | (layer0_outputs[2494]);
    assign outputs[4089] = layer0_outputs[4476];
    assign outputs[4090] = ~((layer0_outputs[9917]) & (layer0_outputs[9102]));
    assign outputs[4091] = layer0_outputs[197];
    assign outputs[4092] = ~((layer0_outputs[8850]) ^ (layer0_outputs[3294]));
    assign outputs[4093] = (layer0_outputs[7129]) & (layer0_outputs[3349]);
    assign outputs[4094] = layer0_outputs[6005];
    assign outputs[4095] = (layer0_outputs[1236]) ^ (layer0_outputs[8679]);
    assign outputs[4096] = layer0_outputs[797];
    assign outputs[4097] = layer0_outputs[5252];
    assign outputs[4098] = ~(layer0_outputs[9647]);
    assign outputs[4099] = (layer0_outputs[931]) | (layer0_outputs[2235]);
    assign outputs[4100] = (layer0_outputs[8533]) & (layer0_outputs[444]);
    assign outputs[4101] = layer0_outputs[7964];
    assign outputs[4102] = (layer0_outputs[10039]) | (layer0_outputs[6662]);
    assign outputs[4103] = ~(layer0_outputs[4358]);
    assign outputs[4104] = ~(layer0_outputs[5897]) | (layer0_outputs[2966]);
    assign outputs[4105] = ~(layer0_outputs[3497]);
    assign outputs[4106] = layer0_outputs[8623];
    assign outputs[4107] = ~(layer0_outputs[5131]);
    assign outputs[4108] = layer0_outputs[4177];
    assign outputs[4109] = ~((layer0_outputs[7472]) & (layer0_outputs[5771]));
    assign outputs[4110] = ~(layer0_outputs[7337]);
    assign outputs[4111] = (layer0_outputs[8269]) & ~(layer0_outputs[8137]);
    assign outputs[4112] = ~(layer0_outputs[9429]);
    assign outputs[4113] = ~(layer0_outputs[6081]);
    assign outputs[4114] = ~(layer0_outputs[1490]) | (layer0_outputs[696]);
    assign outputs[4115] = ~(layer0_outputs[8693]);
    assign outputs[4116] = ~(layer0_outputs[273]);
    assign outputs[4117] = ~(layer0_outputs[10055]);
    assign outputs[4118] = ~(layer0_outputs[10061]);
    assign outputs[4119] = layer0_outputs[5358];
    assign outputs[4120] = ~((layer0_outputs[829]) | (layer0_outputs[9535]));
    assign outputs[4121] = ~(layer0_outputs[2900]);
    assign outputs[4122] = ~(layer0_outputs[7883]);
    assign outputs[4123] = ~((layer0_outputs[9622]) ^ (layer0_outputs[989]));
    assign outputs[4124] = layer0_outputs[5377];
    assign outputs[4125] = ~((layer0_outputs[4759]) ^ (layer0_outputs[6827]));
    assign outputs[4126] = layer0_outputs[7108];
    assign outputs[4127] = ~(layer0_outputs[686]);
    assign outputs[4128] = layer0_outputs[5182];
    assign outputs[4129] = ~(layer0_outputs[4596]) | (layer0_outputs[572]);
    assign outputs[4130] = layer0_outputs[10128];
    assign outputs[4131] = ~((layer0_outputs[5602]) ^ (layer0_outputs[10092]));
    assign outputs[4132] = ~(layer0_outputs[9183]) | (layer0_outputs[5848]);
    assign outputs[4133] = layer0_outputs[1281];
    assign outputs[4134] = layer0_outputs[269];
    assign outputs[4135] = layer0_outputs[752];
    assign outputs[4136] = (layer0_outputs[935]) & ~(layer0_outputs[9049]);
    assign outputs[4137] = ~(layer0_outputs[6752]);
    assign outputs[4138] = layer0_outputs[7424];
    assign outputs[4139] = ~(layer0_outputs[4370]) | (layer0_outputs[5402]);
    assign outputs[4140] = ~(layer0_outputs[9551]);
    assign outputs[4141] = ~(layer0_outputs[6195]);
    assign outputs[4142] = ~(layer0_outputs[3676]);
    assign outputs[4143] = layer0_outputs[9083];
    assign outputs[4144] = ~(layer0_outputs[1529]);
    assign outputs[4145] = (layer0_outputs[6100]) & (layer0_outputs[9716]);
    assign outputs[4146] = (layer0_outputs[9540]) ^ (layer0_outputs[6221]);
    assign outputs[4147] = (layer0_outputs[2068]) & ~(layer0_outputs[7021]);
    assign outputs[4148] = ~(layer0_outputs[9465]);
    assign outputs[4149] = ~(layer0_outputs[4145]);
    assign outputs[4150] = (layer0_outputs[7840]) & (layer0_outputs[1242]);
    assign outputs[4151] = layer0_outputs[10135];
    assign outputs[4152] = layer0_outputs[7388];
    assign outputs[4153] = (layer0_outputs[2810]) & ~(layer0_outputs[5979]);
    assign outputs[4154] = (layer0_outputs[785]) & (layer0_outputs[5136]);
    assign outputs[4155] = ~((layer0_outputs[10230]) | (layer0_outputs[9773]));
    assign outputs[4156] = (layer0_outputs[8883]) & ~(layer0_outputs[4465]);
    assign outputs[4157] = ~(layer0_outputs[3782]);
    assign outputs[4158] = ~(layer0_outputs[4661]);
    assign outputs[4159] = (layer0_outputs[3517]) ^ (layer0_outputs[2698]);
    assign outputs[4160] = layer0_outputs[52];
    assign outputs[4161] = layer0_outputs[7069];
    assign outputs[4162] = (layer0_outputs[5569]) ^ (layer0_outputs[1442]);
    assign outputs[4163] = ~(layer0_outputs[7750]);
    assign outputs[4164] = ~(layer0_outputs[1559]);
    assign outputs[4165] = ~(layer0_outputs[355]);
    assign outputs[4166] = ~(layer0_outputs[3498]);
    assign outputs[4167] = ~(layer0_outputs[5125]);
    assign outputs[4168] = ~(layer0_outputs[3120]);
    assign outputs[4169] = ~(layer0_outputs[3168]);
    assign outputs[4170] = ~(layer0_outputs[10]);
    assign outputs[4171] = ~(layer0_outputs[4543]);
    assign outputs[4172] = ~(layer0_outputs[3496]);
    assign outputs[4173] = ~(layer0_outputs[461]);
    assign outputs[4174] = ~(layer0_outputs[3243]) | (layer0_outputs[2255]);
    assign outputs[4175] = (layer0_outputs[1732]) & ~(layer0_outputs[9041]);
    assign outputs[4176] = ~((layer0_outputs[2541]) & (layer0_outputs[1998]));
    assign outputs[4177] = ~(layer0_outputs[4702]) | (layer0_outputs[947]);
    assign outputs[4178] = ~(layer0_outputs[8818]) | (layer0_outputs[7433]);
    assign outputs[4179] = (layer0_outputs[2660]) & ~(layer0_outputs[6469]);
    assign outputs[4180] = layer0_outputs[7971];
    assign outputs[4181] = ~(layer0_outputs[5369]);
    assign outputs[4182] = ~(layer0_outputs[2129]);
    assign outputs[4183] = layer0_outputs[7969];
    assign outputs[4184] = ~(layer0_outputs[6330]);
    assign outputs[4185] = layer0_outputs[764];
    assign outputs[4186] = (layer0_outputs[8793]) ^ (layer0_outputs[3229]);
    assign outputs[4187] = layer0_outputs[1996];
    assign outputs[4188] = (layer0_outputs[5416]) & ~(layer0_outputs[6248]);
    assign outputs[4189] = ~((layer0_outputs[8819]) ^ (layer0_outputs[5677]));
    assign outputs[4190] = layer0_outputs[9338];
    assign outputs[4191] = layer0_outputs[2109];
    assign outputs[4192] = layer0_outputs[5030];
    assign outputs[4193] = (layer0_outputs[10207]) & (layer0_outputs[8770]);
    assign outputs[4194] = ~(layer0_outputs[6038]);
    assign outputs[4195] = layer0_outputs[1050];
    assign outputs[4196] = (layer0_outputs[6377]) & (layer0_outputs[5149]);
    assign outputs[4197] = ~((layer0_outputs[2416]) ^ (layer0_outputs[8770]));
    assign outputs[4198] = ~((layer0_outputs[3898]) ^ (layer0_outputs[10234]));
    assign outputs[4199] = ~(layer0_outputs[7572]);
    assign outputs[4200] = ~(layer0_outputs[9465]);
    assign outputs[4201] = ~((layer0_outputs[768]) | (layer0_outputs[8782]));
    assign outputs[4202] = ~(layer0_outputs[7688]);
    assign outputs[4203] = layer0_outputs[3578];
    assign outputs[4204] = (layer0_outputs[7174]) ^ (layer0_outputs[5421]);
    assign outputs[4205] = layer0_outputs[2780];
    assign outputs[4206] = layer0_outputs[4817];
    assign outputs[4207] = ~(layer0_outputs[3757]);
    assign outputs[4208] = (layer0_outputs[2578]) | (layer0_outputs[2124]);
    assign outputs[4209] = ~((layer0_outputs[3980]) ^ (layer0_outputs[7565]));
    assign outputs[4210] = (layer0_outputs[9848]) & ~(layer0_outputs[1419]);
    assign outputs[4211] = layer0_outputs[5399];
    assign outputs[4212] = ~((layer0_outputs[5077]) | (layer0_outputs[119]));
    assign outputs[4213] = ~(layer0_outputs[3764]);
    assign outputs[4214] = layer0_outputs[215];
    assign outputs[4215] = (layer0_outputs[3713]) & (layer0_outputs[8250]);
    assign outputs[4216] = (layer0_outputs[5834]) ^ (layer0_outputs[9128]);
    assign outputs[4217] = layer0_outputs[4586];
    assign outputs[4218] = layer0_outputs[7048];
    assign outputs[4219] = layer0_outputs[9629];
    assign outputs[4220] = ~((layer0_outputs[3547]) & (layer0_outputs[7400]));
    assign outputs[4221] = (layer0_outputs[3396]) & (layer0_outputs[3766]);
    assign outputs[4222] = ~(layer0_outputs[5728]);
    assign outputs[4223] = ~((layer0_outputs[5935]) | (layer0_outputs[1567]));
    assign outputs[4224] = (layer0_outputs[2136]) & ~(layer0_outputs[10230]);
    assign outputs[4225] = (layer0_outputs[8323]) & ~(layer0_outputs[8228]);
    assign outputs[4226] = (layer0_outputs[4745]) & (layer0_outputs[8112]);
    assign outputs[4227] = ~(layer0_outputs[4592]) | (layer0_outputs[3116]);
    assign outputs[4228] = layer0_outputs[9130];
    assign outputs[4229] = layer0_outputs[7344];
    assign outputs[4230] = ~(layer0_outputs[612]);
    assign outputs[4231] = ~(layer0_outputs[5870]);
    assign outputs[4232] = ~(layer0_outputs[5318]);
    assign outputs[4233] = layer0_outputs[10217];
    assign outputs[4234] = (layer0_outputs[1493]) & ~(layer0_outputs[7990]);
    assign outputs[4235] = layer0_outputs[6992];
    assign outputs[4236] = ~(layer0_outputs[10100]);
    assign outputs[4237] = layer0_outputs[1213];
    assign outputs[4238] = layer0_outputs[2648];
    assign outputs[4239] = ~(layer0_outputs[1466]);
    assign outputs[4240] = ~(layer0_outputs[3059]);
    assign outputs[4241] = layer0_outputs[4397];
    assign outputs[4242] = ~(layer0_outputs[8183]) | (layer0_outputs[6337]);
    assign outputs[4243] = layer0_outputs[9296];
    assign outputs[4244] = layer0_outputs[4315];
    assign outputs[4245] = layer0_outputs[9196];
    assign outputs[4246] = ~(layer0_outputs[6289]);
    assign outputs[4247] = ~((layer0_outputs[6250]) | (layer0_outputs[1165]));
    assign outputs[4248] = layer0_outputs[2332];
    assign outputs[4249] = layer0_outputs[2499];
    assign outputs[4250] = ~((layer0_outputs[2458]) & (layer0_outputs[6906]));
    assign outputs[4251] = layer0_outputs[2140];
    assign outputs[4252] = (layer0_outputs[738]) & ~(layer0_outputs[3729]);
    assign outputs[4253] = layer0_outputs[5201];
    assign outputs[4254] = layer0_outputs[5176];
    assign outputs[4255] = ~(layer0_outputs[651]);
    assign outputs[4256] = ~(layer0_outputs[6455]) | (layer0_outputs[6046]);
    assign outputs[4257] = layer0_outputs[4294];
    assign outputs[4258] = (layer0_outputs[4540]) & ~(layer0_outputs[1265]);
    assign outputs[4259] = (layer0_outputs[10075]) | (layer0_outputs[8683]);
    assign outputs[4260] = ~((layer0_outputs[9280]) ^ (layer0_outputs[7201]));
    assign outputs[4261] = layer0_outputs[1205];
    assign outputs[4262] = layer0_outputs[7028];
    assign outputs[4263] = layer0_outputs[8681];
    assign outputs[4264] = ~((layer0_outputs[8202]) ^ (layer0_outputs[3829]));
    assign outputs[4265] = (layer0_outputs[4282]) ^ (layer0_outputs[448]);
    assign outputs[4266] = ~((layer0_outputs[4062]) | (layer0_outputs[125]));
    assign outputs[4267] = ~(layer0_outputs[9493]);
    assign outputs[4268] = (layer0_outputs[6846]) | (layer0_outputs[1927]);
    assign outputs[4269] = ~((layer0_outputs[3685]) | (layer0_outputs[4496]));
    assign outputs[4270] = (layer0_outputs[3561]) & (layer0_outputs[4277]);
    assign outputs[4271] = (layer0_outputs[3108]) ^ (layer0_outputs[5495]);
    assign outputs[4272] = (layer0_outputs[9303]) & ~(layer0_outputs[1227]);
    assign outputs[4273] = ~((layer0_outputs[4183]) | (layer0_outputs[4203]));
    assign outputs[4274] = ~((layer0_outputs[760]) | (layer0_outputs[5052]));
    assign outputs[4275] = layer0_outputs[4086];
    assign outputs[4276] = ~(layer0_outputs[10100]);
    assign outputs[4277] = layer0_outputs[7735];
    assign outputs[4278] = layer0_outputs[3908];
    assign outputs[4279] = ~(layer0_outputs[3692]);
    assign outputs[4280] = ~((layer0_outputs[6096]) ^ (layer0_outputs[3592]));
    assign outputs[4281] = layer0_outputs[3966];
    assign outputs[4282] = (layer0_outputs[7043]) & ~(layer0_outputs[1550]);
    assign outputs[4283] = (layer0_outputs[8724]) & ~(layer0_outputs[795]);
    assign outputs[4284] = (layer0_outputs[7251]) ^ (layer0_outputs[3011]);
    assign outputs[4285] = ~((layer0_outputs[406]) & (layer0_outputs[9621]));
    assign outputs[4286] = ~(layer0_outputs[45]) | (layer0_outputs[337]);
    assign outputs[4287] = ~((layer0_outputs[5178]) & (layer0_outputs[4135]));
    assign outputs[4288] = layer0_outputs[2369];
    assign outputs[4289] = ~(layer0_outputs[2237]);
    assign outputs[4290] = ~((layer0_outputs[7027]) & (layer0_outputs[3661]));
    assign outputs[4291] = ~(layer0_outputs[3129]);
    assign outputs[4292] = layer0_outputs[821];
    assign outputs[4293] = (layer0_outputs[2374]) & ~(layer0_outputs[9790]);
    assign outputs[4294] = layer0_outputs[8178];
    assign outputs[4295] = 1'b0;
    assign outputs[4296] = ~(layer0_outputs[2949]) | (layer0_outputs[1539]);
    assign outputs[4297] = ~(layer0_outputs[4118]);
    assign outputs[4298] = ~(layer0_outputs[822]) | (layer0_outputs[8932]);
    assign outputs[4299] = layer0_outputs[5255];
    assign outputs[4300] = ~((layer0_outputs[10074]) ^ (layer0_outputs[9861]));
    assign outputs[4301] = layer0_outputs[584];
    assign outputs[4302] = layer0_outputs[1627];
    assign outputs[4303] = layer0_outputs[9010];
    assign outputs[4304] = layer0_outputs[7739];
    assign outputs[4305] = ~(layer0_outputs[6294]) | (layer0_outputs[5532]);
    assign outputs[4306] = layer0_outputs[6769];
    assign outputs[4307] = ~(layer0_outputs[8895]) | (layer0_outputs[5455]);
    assign outputs[4308] = layer0_outputs[5220];
    assign outputs[4309] = layer0_outputs[4729];
    assign outputs[4310] = ~(layer0_outputs[3319]);
    assign outputs[4311] = ~((layer0_outputs[9483]) ^ (layer0_outputs[9519]));
    assign outputs[4312] = ~(layer0_outputs[9474]);
    assign outputs[4313] = ~((layer0_outputs[6839]) ^ (layer0_outputs[8692]));
    assign outputs[4314] = (layer0_outputs[1341]) ^ (layer0_outputs[695]);
    assign outputs[4315] = ~(layer0_outputs[4486]);
    assign outputs[4316] = layer0_outputs[4461];
    assign outputs[4317] = layer0_outputs[1240];
    assign outputs[4318] = ~(layer0_outputs[6024]);
    assign outputs[4319] = ~(layer0_outputs[5095]) | (layer0_outputs[247]);
    assign outputs[4320] = ~(layer0_outputs[6921]);
    assign outputs[4321] = ~(layer0_outputs[2844]);
    assign outputs[4322] = (layer0_outputs[8683]) ^ (layer0_outputs[4730]);
    assign outputs[4323] = (layer0_outputs[5426]) & ~(layer0_outputs[3371]);
    assign outputs[4324] = ~((layer0_outputs[800]) ^ (layer0_outputs[1337]));
    assign outputs[4325] = ~(layer0_outputs[3023]);
    assign outputs[4326] = (layer0_outputs[1920]) | (layer0_outputs[3738]);
    assign outputs[4327] = ~((layer0_outputs[282]) & (layer0_outputs[3235]));
    assign outputs[4328] = (layer0_outputs[9528]) & ~(layer0_outputs[8839]);
    assign outputs[4329] = ~(layer0_outputs[499]) | (layer0_outputs[3309]);
    assign outputs[4330] = layer0_outputs[1302];
    assign outputs[4331] = ~(layer0_outputs[3177]) | (layer0_outputs[4512]);
    assign outputs[4332] = ~((layer0_outputs[7943]) ^ (layer0_outputs[6055]));
    assign outputs[4333] = ~(layer0_outputs[9114]) | (layer0_outputs[7694]);
    assign outputs[4334] = (layer0_outputs[64]) & (layer0_outputs[5394]);
    assign outputs[4335] = ~((layer0_outputs[3630]) ^ (layer0_outputs[2774]));
    assign outputs[4336] = ~((layer0_outputs[5469]) | (layer0_outputs[4370]));
    assign outputs[4337] = (layer0_outputs[6638]) & (layer0_outputs[9520]);
    assign outputs[4338] = (layer0_outputs[3908]) & (layer0_outputs[10199]);
    assign outputs[4339] = ~(layer0_outputs[10172]);
    assign outputs[4340] = layer0_outputs[3959];
    assign outputs[4341] = layer0_outputs[1321];
    assign outputs[4342] = ~(layer0_outputs[8435]);
    assign outputs[4343] = ~(layer0_outputs[6411]);
    assign outputs[4344] = ~(layer0_outputs[5769]);
    assign outputs[4345] = layer0_outputs[2488];
    assign outputs[4346] = layer0_outputs[3520];
    assign outputs[4347] = (layer0_outputs[10076]) & ~(layer0_outputs[5787]);
    assign outputs[4348] = (layer0_outputs[8942]) | (layer0_outputs[1598]);
    assign outputs[4349] = ~(layer0_outputs[4314]);
    assign outputs[4350] = layer0_outputs[6401];
    assign outputs[4351] = layer0_outputs[4004];
    assign outputs[4352] = layer0_outputs[8217];
    assign outputs[4353] = ~(layer0_outputs[3732]) | (layer0_outputs[8618]);
    assign outputs[4354] = layer0_outputs[9705];
    assign outputs[4355] = ~(layer0_outputs[6317]);
    assign outputs[4356] = ~(layer0_outputs[2240]) | (layer0_outputs[2780]);
    assign outputs[4357] = ~(layer0_outputs[2773]);
    assign outputs[4358] = ~(layer0_outputs[8804]) | (layer0_outputs[2945]);
    assign outputs[4359] = (layer0_outputs[1411]) ^ (layer0_outputs[9638]);
    assign outputs[4360] = ~(layer0_outputs[3324]) | (layer0_outputs[2727]);
    assign outputs[4361] = layer0_outputs[1840];
    assign outputs[4362] = layer0_outputs[7913];
    assign outputs[4363] = ~(layer0_outputs[7145]);
    assign outputs[4364] = ~(layer0_outputs[10096]);
    assign outputs[4365] = ~(layer0_outputs[2406]);
    assign outputs[4366] = (layer0_outputs[8653]) & ~(layer0_outputs[3331]);
    assign outputs[4367] = (layer0_outputs[8080]) ^ (layer0_outputs[6521]);
    assign outputs[4368] = ~(layer0_outputs[933]);
    assign outputs[4369] = layer0_outputs[9742];
    assign outputs[4370] = ~(layer0_outputs[8117]);
    assign outputs[4371] = ~((layer0_outputs[4040]) | (layer0_outputs[9645]));
    assign outputs[4372] = (layer0_outputs[2564]) & (layer0_outputs[1624]);
    assign outputs[4373] = (layer0_outputs[8274]) & ~(layer0_outputs[6970]);
    assign outputs[4374] = ~(layer0_outputs[5630]) | (layer0_outputs[681]);
    assign outputs[4375] = (layer0_outputs[8212]) & ~(layer0_outputs[6910]);
    assign outputs[4376] = layer0_outputs[6861];
    assign outputs[4377] = ~(layer0_outputs[3558]);
    assign outputs[4378] = ~((layer0_outputs[3174]) | (layer0_outputs[8426]));
    assign outputs[4379] = ~(layer0_outputs[1969]);
    assign outputs[4380] = layer0_outputs[9813];
    assign outputs[4381] = layer0_outputs[4654];
    assign outputs[4382] = ~(layer0_outputs[1406]);
    assign outputs[4383] = ~(layer0_outputs[2048]);
    assign outputs[4384] = (layer0_outputs[854]) ^ (layer0_outputs[2046]);
    assign outputs[4385] = ~((layer0_outputs[5235]) | (layer0_outputs[6001]));
    assign outputs[4386] = (layer0_outputs[2638]) & ~(layer0_outputs[4251]);
    assign outputs[4387] = (layer0_outputs[1880]) ^ (layer0_outputs[430]);
    assign outputs[4388] = layer0_outputs[5439];
    assign outputs[4389] = (layer0_outputs[9194]) ^ (layer0_outputs[2037]);
    assign outputs[4390] = (layer0_outputs[9206]) & ~(layer0_outputs[159]);
    assign outputs[4391] = layer0_outputs[6433];
    assign outputs[4392] = (layer0_outputs[9043]) & ~(layer0_outputs[8299]);
    assign outputs[4393] = ~((layer0_outputs[9024]) ^ (layer0_outputs[3740]));
    assign outputs[4394] = ~(layer0_outputs[5481]);
    assign outputs[4395] = layer0_outputs[4342];
    assign outputs[4396] = layer0_outputs[4316];
    assign outputs[4397] = layer0_outputs[805];
    assign outputs[4398] = ~((layer0_outputs[6794]) | (layer0_outputs[2981]));
    assign outputs[4399] = (layer0_outputs[6928]) & ~(layer0_outputs[5631]);
    assign outputs[4400] = layer0_outputs[8630];
    assign outputs[4401] = ~(layer0_outputs[813]);
    assign outputs[4402] = ~(layer0_outputs[3043]);
    assign outputs[4403] = layer0_outputs[3412];
    assign outputs[4404] = (layer0_outputs[5248]) ^ (layer0_outputs[2027]);
    assign outputs[4405] = ~((layer0_outputs[8573]) ^ (layer0_outputs[4998]));
    assign outputs[4406] = layer0_outputs[5528];
    assign outputs[4407] = (layer0_outputs[1020]) & (layer0_outputs[1244]);
    assign outputs[4408] = (layer0_outputs[1839]) & ~(layer0_outputs[9842]);
    assign outputs[4409] = (layer0_outputs[290]) & ~(layer0_outputs[799]);
    assign outputs[4410] = (layer0_outputs[2717]) & ~(layer0_outputs[117]);
    assign outputs[4411] = layer0_outputs[7000];
    assign outputs[4412] = layer0_outputs[300];
    assign outputs[4413] = layer0_outputs[1109];
    assign outputs[4414] = layer0_outputs[6596];
    assign outputs[4415] = ~((layer0_outputs[8707]) ^ (layer0_outputs[5191]));
    assign outputs[4416] = layer0_outputs[1326];
    assign outputs[4417] = ~(layer0_outputs[8689]);
    assign outputs[4418] = ~(layer0_outputs[1643]);
    assign outputs[4419] = ~((layer0_outputs[10079]) & (layer0_outputs[5540]));
    assign outputs[4420] = ~(layer0_outputs[9]);
    assign outputs[4421] = (layer0_outputs[4635]) & ~(layer0_outputs[7616]);
    assign outputs[4422] = ~(layer0_outputs[5924]);
    assign outputs[4423] = ~(layer0_outputs[9292]);
    assign outputs[4424] = ~(layer0_outputs[41]);
    assign outputs[4425] = (layer0_outputs[3918]) | (layer0_outputs[6033]);
    assign outputs[4426] = ~(layer0_outputs[2418]);
    assign outputs[4427] = (layer0_outputs[7483]) & ~(layer0_outputs[4798]);
    assign outputs[4428] = ~(layer0_outputs[3430]);
    assign outputs[4429] = layer0_outputs[5043];
    assign outputs[4430] = ~(layer0_outputs[3799]);
    assign outputs[4431] = ~((layer0_outputs[3282]) ^ (layer0_outputs[5648]));
    assign outputs[4432] = (layer0_outputs[3290]) | (layer0_outputs[402]);
    assign outputs[4433] = (layer0_outputs[7450]) & ~(layer0_outputs[5129]);
    assign outputs[4434] = ~((layer0_outputs[9988]) | (layer0_outputs[3092]));
    assign outputs[4435] = ~(layer0_outputs[3121]);
    assign outputs[4436] = (layer0_outputs[8656]) ^ (layer0_outputs[2877]);
    assign outputs[4437] = ~(layer0_outputs[1572]);
    assign outputs[4438] = ~(layer0_outputs[1994]);
    assign outputs[4439] = ~(layer0_outputs[875]) | (layer0_outputs[6995]);
    assign outputs[4440] = (layer0_outputs[10001]) & ~(layer0_outputs[3111]);
    assign outputs[4441] = ~(layer0_outputs[131]) | (layer0_outputs[2903]);
    assign outputs[4442] = layer0_outputs[3462];
    assign outputs[4443] = layer0_outputs[3042];
    assign outputs[4444] = layer0_outputs[5772];
    assign outputs[4445] = ~((layer0_outputs[7893]) ^ (layer0_outputs[5860]));
    assign outputs[4446] = (layer0_outputs[7614]) ^ (layer0_outputs[6341]);
    assign outputs[4447] = ~((layer0_outputs[8132]) ^ (layer0_outputs[7396]));
    assign outputs[4448] = ~(layer0_outputs[2704]) | (layer0_outputs[2342]);
    assign outputs[4449] = ~((layer0_outputs[6820]) ^ (layer0_outputs[6015]));
    assign outputs[4450] = ~(layer0_outputs[4252]);
    assign outputs[4451] = (layer0_outputs[4122]) & (layer0_outputs[5579]);
    assign outputs[4452] = (layer0_outputs[6162]) ^ (layer0_outputs[5849]);
    assign outputs[4453] = ~(layer0_outputs[926]);
    assign outputs[4454] = ~((layer0_outputs[1139]) ^ (layer0_outputs[229]));
    assign outputs[4455] = (layer0_outputs[4925]) & (layer0_outputs[9752]);
    assign outputs[4456] = (layer0_outputs[7720]) & (layer0_outputs[1953]);
    assign outputs[4457] = ~(layer0_outputs[9805]);
    assign outputs[4458] = ~((layer0_outputs[1049]) | (layer0_outputs[1637]));
    assign outputs[4459] = (layer0_outputs[6592]) & (layer0_outputs[8135]);
    assign outputs[4460] = (layer0_outputs[5342]) & ~(layer0_outputs[7451]);
    assign outputs[4461] = ~(layer0_outputs[3107]);
    assign outputs[4462] = layer0_outputs[3127];
    assign outputs[4463] = ~(layer0_outputs[1807]);
    assign outputs[4464] = ~(layer0_outputs[3940]);
    assign outputs[4465] = (layer0_outputs[582]) ^ (layer0_outputs[9295]);
    assign outputs[4466] = layer0_outputs[4785];
    assign outputs[4467] = ~((layer0_outputs[1608]) ^ (layer0_outputs[1090]));
    assign outputs[4468] = ~(layer0_outputs[256]) | (layer0_outputs[1179]);
    assign outputs[4469] = ~(layer0_outputs[2534]);
    assign outputs[4470] = ~(layer0_outputs[3074]);
    assign outputs[4471] = layer0_outputs[483];
    assign outputs[4472] = ~((layer0_outputs[3896]) | (layer0_outputs[3117]));
    assign outputs[4473] = layer0_outputs[2778];
    assign outputs[4474] = layer0_outputs[5122];
    assign outputs[4475] = (layer0_outputs[3437]) ^ (layer0_outputs[3871]);
    assign outputs[4476] = ~(layer0_outputs[10068]);
    assign outputs[4477] = layer0_outputs[2190];
    assign outputs[4478] = ~((layer0_outputs[1665]) ^ (layer0_outputs[1088]));
    assign outputs[4479] = layer0_outputs[8759];
    assign outputs[4480] = layer0_outputs[6258];
    assign outputs[4481] = ~((layer0_outputs[4604]) & (layer0_outputs[5839]));
    assign outputs[4482] = ~(layer0_outputs[5729]) | (layer0_outputs[7394]);
    assign outputs[4483] = ~((layer0_outputs[3532]) | (layer0_outputs[353]));
    assign outputs[4484] = (layer0_outputs[1264]) & ~(layer0_outputs[8485]);
    assign outputs[4485] = ~((layer0_outputs[9576]) ^ (layer0_outputs[1704]));
    assign outputs[4486] = ~(layer0_outputs[1160]);
    assign outputs[4487] = ~(layer0_outputs[8465]);
    assign outputs[4488] = ~(layer0_outputs[2085]);
    assign outputs[4489] = layer0_outputs[6700];
    assign outputs[4490] = ~((layer0_outputs[7324]) ^ (layer0_outputs[5610]));
    assign outputs[4491] = ~(layer0_outputs[6698]) | (layer0_outputs[4753]);
    assign outputs[4492] = ~(layer0_outputs[9844]);
    assign outputs[4493] = (layer0_outputs[4706]) & ~(layer0_outputs[9709]);
    assign outputs[4494] = (layer0_outputs[3920]) & (layer0_outputs[9900]);
    assign outputs[4495] = ~(layer0_outputs[969]);
    assign outputs[4496] = (layer0_outputs[6431]) & (layer0_outputs[9282]);
    assign outputs[4497] = ~(layer0_outputs[5065]) | (layer0_outputs[6023]);
    assign outputs[4498] = (layer0_outputs[9364]) & ~(layer0_outputs[8930]);
    assign outputs[4499] = layer0_outputs[3407];
    assign outputs[4500] = ~(layer0_outputs[8292]);
    assign outputs[4501] = ~((layer0_outputs[5487]) | (layer0_outputs[5261]));
    assign outputs[4502] = ~(layer0_outputs[3865]) | (layer0_outputs[3584]);
    assign outputs[4503] = layer0_outputs[4824];
    assign outputs[4504] = ~(layer0_outputs[3378]);
    assign outputs[4505] = (layer0_outputs[6788]) & ~(layer0_outputs[6733]);
    assign outputs[4506] = layer0_outputs[3857];
    assign outputs[4507] = layer0_outputs[9517];
    assign outputs[4508] = layer0_outputs[3549];
    assign outputs[4509] = ~(layer0_outputs[1601]);
    assign outputs[4510] = layer0_outputs[9369];
    assign outputs[4511] = ~(layer0_outputs[7949]);
    assign outputs[4512] = ~((layer0_outputs[1568]) ^ (layer0_outputs[4607]));
    assign outputs[4513] = ~((layer0_outputs[9402]) | (layer0_outputs[4042]));
    assign outputs[4514] = ~((layer0_outputs[932]) ^ (layer0_outputs[1230]));
    assign outputs[4515] = (layer0_outputs[4414]) & ~(layer0_outputs[960]);
    assign outputs[4516] = layer0_outputs[2303];
    assign outputs[4517] = ~((layer0_outputs[2313]) ^ (layer0_outputs[3350]));
    assign outputs[4518] = ~((layer0_outputs[6236]) ^ (layer0_outputs[6652]));
    assign outputs[4519] = (layer0_outputs[5780]) & ~(layer0_outputs[8859]);
    assign outputs[4520] = (layer0_outputs[5533]) ^ (layer0_outputs[5986]);
    assign outputs[4521] = (layer0_outputs[2963]) & ~(layer0_outputs[4327]);
    assign outputs[4522] = (layer0_outputs[7681]) & (layer0_outputs[2631]);
    assign outputs[4523] = ~(layer0_outputs[4510]);
    assign outputs[4524] = layer0_outputs[4506];
    assign outputs[4525] = layer0_outputs[8284];
    assign outputs[4526] = (layer0_outputs[8478]) | (layer0_outputs[6270]);
    assign outputs[4527] = layer0_outputs[2058];
    assign outputs[4528] = layer0_outputs[6549];
    assign outputs[4529] = (layer0_outputs[3185]) ^ (layer0_outputs[6605]);
    assign outputs[4530] = ~(layer0_outputs[5321]);
    assign outputs[4531] = ~((layer0_outputs[2831]) ^ (layer0_outputs[3675]));
    assign outputs[4532] = (layer0_outputs[3464]) & (layer0_outputs[8606]);
    assign outputs[4533] = ~((layer0_outputs[4854]) ^ (layer0_outputs[5480]));
    assign outputs[4534] = ~((layer0_outputs[1542]) | (layer0_outputs[6762]));
    assign outputs[4535] = (layer0_outputs[329]) ^ (layer0_outputs[7939]);
    assign outputs[4536] = (layer0_outputs[7507]) & (layer0_outputs[7189]);
    assign outputs[4537] = (layer0_outputs[4918]) ^ (layer0_outputs[6223]);
    assign outputs[4538] = ~(layer0_outputs[3622]);
    assign outputs[4539] = layer0_outputs[9582];
    assign outputs[4540] = layer0_outputs[9009];
    assign outputs[4541] = ~(layer0_outputs[1215]);
    assign outputs[4542] = ~(layer0_outputs[6283]);
    assign outputs[4543] = layer0_outputs[443];
    assign outputs[4544] = ~(layer0_outputs[7585]);
    assign outputs[4545] = (layer0_outputs[5814]) | (layer0_outputs[9104]);
    assign outputs[4546] = ~(layer0_outputs[7378]);
    assign outputs[4547] = ~(layer0_outputs[3162]);
    assign outputs[4548] = layer0_outputs[7596];
    assign outputs[4549] = ~((layer0_outputs[9326]) | (layer0_outputs[7192]));
    assign outputs[4550] = ~(layer0_outputs[164]);
    assign outputs[4551] = (layer0_outputs[761]) & ~(layer0_outputs[4616]);
    assign outputs[4552] = layer0_outputs[5372];
    assign outputs[4553] = layer0_outputs[6675];
    assign outputs[4554] = layer0_outputs[1119];
    assign outputs[4555] = ~((layer0_outputs[9821]) | (layer0_outputs[793]));
    assign outputs[4556] = ~((layer0_outputs[8001]) ^ (layer0_outputs[8858]));
    assign outputs[4557] = ~(layer0_outputs[2823]) | (layer0_outputs[1700]);
    assign outputs[4558] = ~((layer0_outputs[10034]) ^ (layer0_outputs[8281]));
    assign outputs[4559] = ~(layer0_outputs[2231]);
    assign outputs[4560] = ~(layer0_outputs[4267]);
    assign outputs[4561] = layer0_outputs[343];
    assign outputs[4562] = ~(layer0_outputs[111]);
    assign outputs[4563] = (layer0_outputs[1181]) ^ (layer0_outputs[7476]);
    assign outputs[4564] = ~(layer0_outputs[5404]) | (layer0_outputs[7781]);
    assign outputs[4565] = ~(layer0_outputs[2004]);
    assign outputs[4566] = ~(layer0_outputs[4270]);
    assign outputs[4567] = ~(layer0_outputs[790]);
    assign outputs[4568] = layer0_outputs[6401];
    assign outputs[4569] = ~((layer0_outputs[9045]) | (layer0_outputs[3331]));
    assign outputs[4570] = (layer0_outputs[7323]) & ~(layer0_outputs[6025]);
    assign outputs[4571] = layer0_outputs[5444];
    assign outputs[4572] = layer0_outputs[9612];
    assign outputs[4573] = (layer0_outputs[7567]) ^ (layer0_outputs[2542]);
    assign outputs[4574] = ~(layer0_outputs[2795]);
    assign outputs[4575] = (layer0_outputs[716]) ^ (layer0_outputs[8124]);
    assign outputs[4576] = ~((layer0_outputs[4200]) & (layer0_outputs[2726]));
    assign outputs[4577] = ~(layer0_outputs[3679]);
    assign outputs[4578] = layer0_outputs[5385];
    assign outputs[4579] = ~(layer0_outputs[984]);
    assign outputs[4580] = ~(layer0_outputs[5632]);
    assign outputs[4581] = (layer0_outputs[307]) & (layer0_outputs[2583]);
    assign outputs[4582] = (layer0_outputs[9917]) | (layer0_outputs[535]);
    assign outputs[4583] = layer0_outputs[7588];
    assign outputs[4584] = ~(layer0_outputs[5713]);
    assign outputs[4585] = layer0_outputs[5721];
    assign outputs[4586] = ~(layer0_outputs[7248]);
    assign outputs[4587] = ~(layer0_outputs[1633]);
    assign outputs[4588] = ~(layer0_outputs[3837]);
    assign outputs[4589] = (layer0_outputs[6097]) & ~(layer0_outputs[9859]);
    assign outputs[4590] = ~(layer0_outputs[2071]) | (layer0_outputs[3851]);
    assign outputs[4591] = ~(layer0_outputs[10228]);
    assign outputs[4592] = layer0_outputs[3672];
    assign outputs[4593] = ~(layer0_outputs[2762]);
    assign outputs[4594] = ~(layer0_outputs[3981]);
    assign outputs[4595] = ~((layer0_outputs[9775]) ^ (layer0_outputs[8247]));
    assign outputs[4596] = (layer0_outputs[306]) ^ (layer0_outputs[7715]);
    assign outputs[4597] = (layer0_outputs[6113]) & ~(layer0_outputs[3989]);
    assign outputs[4598] = ~((layer0_outputs[1435]) ^ (layer0_outputs[5704]));
    assign outputs[4599] = (layer0_outputs[9719]) & ~(layer0_outputs[1571]);
    assign outputs[4600] = (layer0_outputs[8434]) & (layer0_outputs[9256]);
    assign outputs[4601] = ~((layer0_outputs[5640]) ^ (layer0_outputs[7877]));
    assign outputs[4602] = ~((layer0_outputs[5155]) ^ (layer0_outputs[1549]));
    assign outputs[4603] = ~((layer0_outputs[8204]) ^ (layer0_outputs[2421]));
    assign outputs[4604] = (layer0_outputs[8051]) & ~(layer0_outputs[8137]);
    assign outputs[4605] = ~(layer0_outputs[4527]);
    assign outputs[4606] = layer0_outputs[2589];
    assign outputs[4607] = (layer0_outputs[988]) & (layer0_outputs[2354]);
    assign outputs[4608] = ~(layer0_outputs[4140]);
    assign outputs[4609] = ~(layer0_outputs[5460]);
    assign outputs[4610] = ~(layer0_outputs[10079]) | (layer0_outputs[8943]);
    assign outputs[4611] = ~(layer0_outputs[9451]);
    assign outputs[4612] = (layer0_outputs[6200]) & ~(layer0_outputs[4901]);
    assign outputs[4613] = ~(layer0_outputs[2174]);
    assign outputs[4614] = ~(layer0_outputs[7817]);
    assign outputs[4615] = ~(layer0_outputs[1238]);
    assign outputs[4616] = ~(layer0_outputs[4772]);
    assign outputs[4617] = (layer0_outputs[7974]) & ~(layer0_outputs[5475]);
    assign outputs[4618] = ~((layer0_outputs[10106]) ^ (layer0_outputs[6310]));
    assign outputs[4619] = layer0_outputs[5170];
    assign outputs[4620] = layer0_outputs[8825];
    assign outputs[4621] = (layer0_outputs[9677]) & (layer0_outputs[3973]);
    assign outputs[4622] = ~(layer0_outputs[5475]);
    assign outputs[4623] = (layer0_outputs[9542]) & ~(layer0_outputs[4038]);
    assign outputs[4624] = ~(layer0_outputs[748]);
    assign outputs[4625] = layer0_outputs[7637];
    assign outputs[4626] = (layer0_outputs[9265]) ^ (layer0_outputs[4643]);
    assign outputs[4627] = ~((layer0_outputs[274]) | (layer0_outputs[2986]));
    assign outputs[4628] = (layer0_outputs[5757]) ^ (layer0_outputs[762]);
    assign outputs[4629] = ~(layer0_outputs[8923]);
    assign outputs[4630] = ~((layer0_outputs[5135]) | (layer0_outputs[3648]));
    assign outputs[4631] = layer0_outputs[7898];
    assign outputs[4632] = layer0_outputs[7203];
    assign outputs[4633] = (layer0_outputs[6075]) & (layer0_outputs[2796]);
    assign outputs[4634] = ~((layer0_outputs[9251]) | (layer0_outputs[2690]));
    assign outputs[4635] = ~(layer0_outputs[6336]);
    assign outputs[4636] = (layer0_outputs[5228]) ^ (layer0_outputs[4468]);
    assign outputs[4637] = (layer0_outputs[3240]) & (layer0_outputs[1543]);
    assign outputs[4638] = ~(layer0_outputs[6426]);
    assign outputs[4639] = ~(layer0_outputs[7624]);
    assign outputs[4640] = ~((layer0_outputs[9220]) | (layer0_outputs[2925]));
    assign outputs[4641] = ~(layer0_outputs[2562]);
    assign outputs[4642] = ~(layer0_outputs[6545]) | (layer0_outputs[8293]);
    assign outputs[4643] = layer0_outputs[3545];
    assign outputs[4644] = (layer0_outputs[990]) & (layer0_outputs[2302]);
    assign outputs[4645] = layer0_outputs[1743];
    assign outputs[4646] = ~(layer0_outputs[1878]);
    assign outputs[4647] = ~(layer0_outputs[10072]);
    assign outputs[4648] = (layer0_outputs[6161]) & (layer0_outputs[7948]);
    assign outputs[4649] = (layer0_outputs[9847]) ^ (layer0_outputs[9634]);
    assign outputs[4650] = ~(layer0_outputs[7250]);
    assign outputs[4651] = ~(layer0_outputs[4200]) | (layer0_outputs[2428]);
    assign outputs[4652] = ~((layer0_outputs[9787]) & (layer0_outputs[6941]));
    assign outputs[4653] = (layer0_outputs[8682]) ^ (layer0_outputs[5853]);
    assign outputs[4654] = ~(layer0_outputs[7983]);
    assign outputs[4655] = (layer0_outputs[4093]) | (layer0_outputs[535]);
    assign outputs[4656] = ~((layer0_outputs[5813]) ^ (layer0_outputs[414]));
    assign outputs[4657] = (layer0_outputs[3369]) & ~(layer0_outputs[6030]);
    assign outputs[4658] = (layer0_outputs[455]) & (layer0_outputs[8847]);
    assign outputs[4659] = ~(layer0_outputs[8093]);
    assign outputs[4660] = (layer0_outputs[6987]) ^ (layer0_outputs[2487]);
    assign outputs[4661] = ~(layer0_outputs[6539]);
    assign outputs[4662] = ~(layer0_outputs[6998]);
    assign outputs[4663] = (layer0_outputs[2028]) & (layer0_outputs[7906]);
    assign outputs[4664] = (layer0_outputs[3766]) & ~(layer0_outputs[7311]);
    assign outputs[4665] = ~(layer0_outputs[4644]);
    assign outputs[4666] = layer0_outputs[8056];
    assign outputs[4667] = ~(layer0_outputs[6366]);
    assign outputs[4668] = ~(layer0_outputs[9992]);
    assign outputs[4669] = ~(layer0_outputs[9031]);
    assign outputs[4670] = (layer0_outputs[490]) & ~(layer0_outputs[9736]);
    assign outputs[4671] = layer0_outputs[9672];
    assign outputs[4672] = ~((layer0_outputs[143]) & (layer0_outputs[5065]));
    assign outputs[4673] = ~((layer0_outputs[6059]) | (layer0_outputs[4534]));
    assign outputs[4674] = ~(layer0_outputs[8078]);
    assign outputs[4675] = layer0_outputs[2386];
    assign outputs[4676] = ~(layer0_outputs[7150]);
    assign outputs[4677] = layer0_outputs[3549];
    assign outputs[4678] = ~((layer0_outputs[6329]) | (layer0_outputs[2864]));
    assign outputs[4679] = ~(layer0_outputs[3974]);
    assign outputs[4680] = (layer0_outputs[9895]) & ~(layer0_outputs[1729]);
    assign outputs[4681] = layer0_outputs[10160];
    assign outputs[4682] = layer0_outputs[1078];
    assign outputs[4683] = ~(layer0_outputs[9313]);
    assign outputs[4684] = ~(layer0_outputs[859]) | (layer0_outputs[5676]);
    assign outputs[4685] = ~(layer0_outputs[6838]) | (layer0_outputs[4657]);
    assign outputs[4686] = ~(layer0_outputs[1006]);
    assign outputs[4687] = ~(layer0_outputs[5770]);
    assign outputs[4688] = ~(layer0_outputs[8431]);
    assign outputs[4689] = ~((layer0_outputs[4079]) ^ (layer0_outputs[1788]));
    assign outputs[4690] = ~(layer0_outputs[882]);
    assign outputs[4691] = ~((layer0_outputs[7331]) ^ (layer0_outputs[1154]));
    assign outputs[4692] = layer0_outputs[706];
    assign outputs[4693] = ~(layer0_outputs[1881]);
    assign outputs[4694] = (layer0_outputs[5792]) & (layer0_outputs[904]);
    assign outputs[4695] = ~(layer0_outputs[4131]);
    assign outputs[4696] = layer0_outputs[7562];
    assign outputs[4697] = (layer0_outputs[4688]) & (layer0_outputs[8491]);
    assign outputs[4698] = layer0_outputs[8742];
    assign outputs[4699] = ~((layer0_outputs[927]) & (layer0_outputs[8248]));
    assign outputs[4700] = (layer0_outputs[6581]) & (layer0_outputs[8134]);
    assign outputs[4701] = ~(layer0_outputs[9967]) | (layer0_outputs[6300]);
    assign outputs[4702] = ~(layer0_outputs[8565]);
    assign outputs[4703] = layer0_outputs[7309];
    assign outputs[4704] = (layer0_outputs[3039]) ^ (layer0_outputs[9978]);
    assign outputs[4705] = layer0_outputs[1316];
    assign outputs[4706] = ~(layer0_outputs[6369]);
    assign outputs[4707] = ~((layer0_outputs[3056]) ^ (layer0_outputs[6518]));
    assign outputs[4708] = (layer0_outputs[893]) & ~(layer0_outputs[1361]);
    assign outputs[4709] = ~(layer0_outputs[3173]) | (layer0_outputs[6870]);
    assign outputs[4710] = ~(layer0_outputs[8665]);
    assign outputs[4711] = (layer0_outputs[5173]) & ~(layer0_outputs[1463]);
    assign outputs[4712] = layer0_outputs[4840];
    assign outputs[4713] = ~(layer0_outputs[4197]);
    assign outputs[4714] = (layer0_outputs[5282]) ^ (layer0_outputs[7004]);
    assign outputs[4715] = ~(layer0_outputs[5266]);
    assign outputs[4716] = ~(layer0_outputs[8649]);
    assign outputs[4717] = (layer0_outputs[6996]) | (layer0_outputs[2652]);
    assign outputs[4718] = (layer0_outputs[70]) & ~(layer0_outputs[8867]);
    assign outputs[4719] = ~(layer0_outputs[8319]);
    assign outputs[4720] = layer0_outputs[4951];
    assign outputs[4721] = ~((layer0_outputs[207]) ^ (layer0_outputs[6831]));
    assign outputs[4722] = ~(layer0_outputs[5405]) | (layer0_outputs[5714]);
    assign outputs[4723] = layer0_outputs[5337];
    assign outputs[4724] = (layer0_outputs[9494]) | (layer0_outputs[8863]);
    assign outputs[4725] = (layer0_outputs[6186]) & ~(layer0_outputs[4988]);
    assign outputs[4726] = ~(layer0_outputs[6420]);
    assign outputs[4727] = ~(layer0_outputs[5153]);
    assign outputs[4728] = layer0_outputs[7114];
    assign outputs[4729] = ~(layer0_outputs[5773]);
    assign outputs[4730] = ~(layer0_outputs[3854]);
    assign outputs[4731] = ~(layer0_outputs[9349]);
    assign outputs[4732] = layer0_outputs[1935];
    assign outputs[4733] = (layer0_outputs[3699]) & (layer0_outputs[6421]);
    assign outputs[4734] = ~(layer0_outputs[7922]);
    assign outputs[4735] = ~(layer0_outputs[2777]) | (layer0_outputs[1817]);
    assign outputs[4736] = layer0_outputs[4917];
    assign outputs[4737] = ~(layer0_outputs[1983]);
    assign outputs[4738] = ~((layer0_outputs[9997]) & (layer0_outputs[8308]));
    assign outputs[4739] = ~(layer0_outputs[7606]);
    assign outputs[4740] = ~((layer0_outputs[10164]) ^ (layer0_outputs[3452]));
    assign outputs[4741] = (layer0_outputs[9649]) ^ (layer0_outputs[3383]);
    assign outputs[4742] = layer0_outputs[6701];
    assign outputs[4743] = ~(layer0_outputs[10010]);
    assign outputs[4744] = ~(layer0_outputs[7697]);
    assign outputs[4745] = layer0_outputs[4454];
    assign outputs[4746] = layer0_outputs[9692];
    assign outputs[4747] = ~(layer0_outputs[9119]);
    assign outputs[4748] = layer0_outputs[8650];
    assign outputs[4749] = ~(layer0_outputs[5810]);
    assign outputs[4750] = layer0_outputs[5104];
    assign outputs[4751] = (layer0_outputs[1536]) & ~(layer0_outputs[3220]);
    assign outputs[4752] = layer0_outputs[9104];
    assign outputs[4753] = ~(layer0_outputs[5463]);
    assign outputs[4754] = (layer0_outputs[1140]) ^ (layer0_outputs[5100]);
    assign outputs[4755] = ~(layer0_outputs[4393]);
    assign outputs[4756] = (layer0_outputs[7869]) & ~(layer0_outputs[7624]);
    assign outputs[4757] = (layer0_outputs[1119]) & ~(layer0_outputs[4217]);
    assign outputs[4758] = layer0_outputs[3420];
    assign outputs[4759] = ~(layer0_outputs[7107]);
    assign outputs[4760] = ~(layer0_outputs[9415]);
    assign outputs[4761] = layer0_outputs[5037];
    assign outputs[4762] = layer0_outputs[2869];
    assign outputs[4763] = ~((layer0_outputs[10095]) ^ (layer0_outputs[3899]));
    assign outputs[4764] = layer0_outputs[1554];
    assign outputs[4765] = (layer0_outputs[7224]) ^ (layer0_outputs[6097]);
    assign outputs[4766] = layer0_outputs[6154];
    assign outputs[4767] = ~(layer0_outputs[3433]);
    assign outputs[4768] = ~((layer0_outputs[5784]) ^ (layer0_outputs[2678]));
    assign outputs[4769] = (layer0_outputs[5983]) | (layer0_outputs[8889]);
    assign outputs[4770] = ~((layer0_outputs[4672]) ^ (layer0_outputs[2208]));
    assign outputs[4771] = layer0_outputs[2234];
    assign outputs[4772] = (layer0_outputs[1199]) & (layer0_outputs[3061]);
    assign outputs[4773] = layer0_outputs[1660];
    assign outputs[4774] = ~((layer0_outputs[6799]) ^ (layer0_outputs[4122]));
    assign outputs[4775] = layer0_outputs[6373];
    assign outputs[4776] = (layer0_outputs[5217]) ^ (layer0_outputs[4023]);
    assign outputs[4777] = ~(layer0_outputs[4319]);
    assign outputs[4778] = ~((layer0_outputs[6540]) ^ (layer0_outputs[2883]));
    assign outputs[4779] = (layer0_outputs[3515]) ^ (layer0_outputs[9602]);
    assign outputs[4780] = (layer0_outputs[5850]) & ~(layer0_outputs[965]);
    assign outputs[4781] = layer0_outputs[6895];
    assign outputs[4782] = ~(layer0_outputs[1373]);
    assign outputs[4783] = ~(layer0_outputs[5712]) | (layer0_outputs[5585]);
    assign outputs[4784] = layer0_outputs[7661];
    assign outputs[4785] = (layer0_outputs[864]) & ~(layer0_outputs[4954]);
    assign outputs[4786] = (layer0_outputs[1661]) & (layer0_outputs[8880]);
    assign outputs[4787] = (layer0_outputs[8326]) & (layer0_outputs[915]);
    assign outputs[4788] = ~((layer0_outputs[3558]) ^ (layer0_outputs[9396]));
    assign outputs[4789] = ~(layer0_outputs[4584]);
    assign outputs[4790] = layer0_outputs[2573];
    assign outputs[4791] = ~(layer0_outputs[8610]) | (layer0_outputs[3108]);
    assign outputs[4792] = layer0_outputs[4924];
    assign outputs[4793] = layer0_outputs[7923];
    assign outputs[4794] = (layer0_outputs[788]) & ~(layer0_outputs[895]);
    assign outputs[4795] = ~((layer0_outputs[319]) & (layer0_outputs[4483]));
    assign outputs[4796] = (layer0_outputs[1632]) ^ (layer0_outputs[6084]);
    assign outputs[4797] = (layer0_outputs[9905]) & (layer0_outputs[2907]);
    assign outputs[4798] = ~(layer0_outputs[563]);
    assign outputs[4799] = (layer0_outputs[3416]) & (layer0_outputs[561]);
    assign outputs[4800] = ~((layer0_outputs[4450]) | (layer0_outputs[9155]));
    assign outputs[4801] = ~(layer0_outputs[9976]);
    assign outputs[4802] = (layer0_outputs[6708]) ^ (layer0_outputs[8503]);
    assign outputs[4803] = ~((layer0_outputs[6189]) ^ (layer0_outputs[3617]));
    assign outputs[4804] = layer0_outputs[3857];
    assign outputs[4805] = ~(layer0_outputs[7533]);
    assign outputs[4806] = ~(layer0_outputs[6910]);
    assign outputs[4807] = layer0_outputs[949];
    assign outputs[4808] = (layer0_outputs[1271]) & ~(layer0_outputs[884]);
    assign outputs[4809] = ~((layer0_outputs[9028]) | (layer0_outputs[8795]));
    assign outputs[4810] = ~(layer0_outputs[2048]);
    assign outputs[4811] = ~((layer0_outputs[3745]) | (layer0_outputs[5454]));
    assign outputs[4812] = layer0_outputs[10148];
    assign outputs[4813] = ~(layer0_outputs[2799]);
    assign outputs[4814] = (layer0_outputs[9200]) | (layer0_outputs[2249]);
    assign outputs[4815] = layer0_outputs[10213];
    assign outputs[4816] = ~((layer0_outputs[8921]) | (layer0_outputs[6130]));
    assign outputs[4817] = ~(layer0_outputs[8049]);
    assign outputs[4818] = ~(layer0_outputs[4660]);
    assign outputs[4819] = ~(layer0_outputs[7965]);
    assign outputs[4820] = ~(layer0_outputs[6629]);
    assign outputs[4821] = ~(layer0_outputs[5822]);
    assign outputs[4822] = (layer0_outputs[1681]) & ~(layer0_outputs[8499]);
    assign outputs[4823] = layer0_outputs[8251];
    assign outputs[4824] = ~(layer0_outputs[8191]);
    assign outputs[4825] = ~(layer0_outputs[4845]);
    assign outputs[4826] = ~(layer0_outputs[1739]);
    assign outputs[4827] = layer0_outputs[948];
    assign outputs[4828] = layer0_outputs[4939];
    assign outputs[4829] = ~(layer0_outputs[8362]);
    assign outputs[4830] = ~((layer0_outputs[5949]) ^ (layer0_outputs[2944]));
    assign outputs[4831] = (layer0_outputs[6017]) & (layer0_outputs[3139]);
    assign outputs[4832] = ~(layer0_outputs[4594]);
    assign outputs[4833] = ~(layer0_outputs[8834]);
    assign outputs[4834] = layer0_outputs[10177];
    assign outputs[4835] = (layer0_outputs[6553]) & ~(layer0_outputs[5403]);
    assign outputs[4836] = ~(layer0_outputs[5311]);
    assign outputs[4837] = ~((layer0_outputs[1620]) ^ (layer0_outputs[1715]));
    assign outputs[4838] = (layer0_outputs[3593]) ^ (layer0_outputs[1668]);
    assign outputs[4839] = layer0_outputs[3901];
    assign outputs[4840] = layer0_outputs[5764];
    assign outputs[4841] = layer0_outputs[5204];
    assign outputs[4842] = ~(layer0_outputs[3427]);
    assign outputs[4843] = ~((layer0_outputs[1809]) ^ (layer0_outputs[8461]));
    assign outputs[4844] = layer0_outputs[187];
    assign outputs[4845] = (layer0_outputs[9173]) & ~(layer0_outputs[6468]);
    assign outputs[4846] = layer0_outputs[5548];
    assign outputs[4847] = (layer0_outputs[6492]) | (layer0_outputs[9224]);
    assign outputs[4848] = layer0_outputs[6282];
    assign outputs[4849] = ~((layer0_outputs[3631]) ^ (layer0_outputs[8795]));
    assign outputs[4850] = ~(layer0_outputs[7382]);
    assign outputs[4851] = (layer0_outputs[954]) & (layer0_outputs[6962]);
    assign outputs[4852] = (layer0_outputs[4311]) ^ (layer0_outputs[3267]);
    assign outputs[4853] = ~((layer0_outputs[787]) | (layer0_outputs[7843]));
    assign outputs[4854] = (layer0_outputs[3209]) & ~(layer0_outputs[9212]);
    assign outputs[4855] = ~(layer0_outputs[9633]);
    assign outputs[4856] = ~(layer0_outputs[2743]);
    assign outputs[4857] = (layer0_outputs[7834]) ^ (layer0_outputs[10108]);
    assign outputs[4858] = ~(layer0_outputs[5278]);
    assign outputs[4859] = ~(layer0_outputs[327]);
    assign outputs[4860] = layer0_outputs[9595];
    assign outputs[4861] = ~(layer0_outputs[8108]);
    assign outputs[4862] = ~((layer0_outputs[9377]) ^ (layer0_outputs[1915]));
    assign outputs[4863] = ~((layer0_outputs[1719]) ^ (layer0_outputs[2480]));
    assign outputs[4864] = ~(layer0_outputs[2956]) | (layer0_outputs[5994]);
    assign outputs[4865] = ~(layer0_outputs[2180]);
    assign outputs[4866] = (layer0_outputs[10151]) ^ (layer0_outputs[6689]);
    assign outputs[4867] = (layer0_outputs[885]) ^ (layer0_outputs[6041]);
    assign outputs[4868] = ~(layer0_outputs[284]);
    assign outputs[4869] = layer0_outputs[2771];
    assign outputs[4870] = ~(layer0_outputs[3333]);
    assign outputs[4871] = layer0_outputs[8637];
    assign outputs[4872] = ~(layer0_outputs[6622]) | (layer0_outputs[2333]);
    assign outputs[4873] = ~(layer0_outputs[5935]);
    assign outputs[4874] = ~((layer0_outputs[4738]) ^ (layer0_outputs[3363]));
    assign outputs[4875] = (layer0_outputs[7941]) ^ (layer0_outputs[9527]);
    assign outputs[4876] = (layer0_outputs[2892]) & ~(layer0_outputs[909]);
    assign outputs[4877] = layer0_outputs[3487];
    assign outputs[4878] = ~(layer0_outputs[7175]);
    assign outputs[4879] = ~(layer0_outputs[6830]);
    assign outputs[4880] = ~(layer0_outputs[882]);
    assign outputs[4881] = ~((layer0_outputs[3416]) ^ (layer0_outputs[1392]));
    assign outputs[4882] = (layer0_outputs[4270]) ^ (layer0_outputs[8928]);
    assign outputs[4883] = (layer0_outputs[2112]) & ~(layer0_outputs[6912]);
    assign outputs[4884] = (layer0_outputs[6241]) & ~(layer0_outputs[8141]);
    assign outputs[4885] = ~(layer0_outputs[10057]);
    assign outputs[4886] = (layer0_outputs[3684]) & ~(layer0_outputs[10145]);
    assign outputs[4887] = layer0_outputs[6003];
    assign outputs[4888] = (layer0_outputs[3847]) & ~(layer0_outputs[9139]);
    assign outputs[4889] = ~(layer0_outputs[6707]);
    assign outputs[4890] = ~(layer0_outputs[246]);
    assign outputs[4891] = (layer0_outputs[3718]) & (layer0_outputs[6436]);
    assign outputs[4892] = layer0_outputs[7212];
    assign outputs[4893] = layer0_outputs[4703];
    assign outputs[4894] = ~(layer0_outputs[4186]);
    assign outputs[4895] = ~((layer0_outputs[7466]) ^ (layer0_outputs[5684]));
    assign outputs[4896] = layer0_outputs[8578];
    assign outputs[4897] = ~((layer0_outputs[4328]) ^ (layer0_outputs[4445]));
    assign outputs[4898] = (layer0_outputs[6309]) | (layer0_outputs[1649]);
    assign outputs[4899] = (layer0_outputs[4755]) | (layer0_outputs[647]);
    assign outputs[4900] = layer0_outputs[4411];
    assign outputs[4901] = (layer0_outputs[5798]) & (layer0_outputs[9013]);
    assign outputs[4902] = ~((layer0_outputs[7024]) ^ (layer0_outputs[3601]));
    assign outputs[4903] = ~(layer0_outputs[7340]);
    assign outputs[4904] = layer0_outputs[572];
    assign outputs[4905] = layer0_outputs[7372];
    assign outputs[4906] = ~(layer0_outputs[7157]);
    assign outputs[4907] = (layer0_outputs[231]) ^ (layer0_outputs[7924]);
    assign outputs[4908] = layer0_outputs[681];
    assign outputs[4909] = ~(layer0_outputs[7873]);
    assign outputs[4910] = layer0_outputs[3460];
    assign outputs[4911] = layer0_outputs[3156];
    assign outputs[4912] = layer0_outputs[7791];
    assign outputs[4913] = layer0_outputs[2162];
    assign outputs[4914] = ~(layer0_outputs[3033]);
    assign outputs[4915] = layer0_outputs[5000];
    assign outputs[4916] = ~(layer0_outputs[9054]);
    assign outputs[4917] = layer0_outputs[2832];
    assign outputs[4918] = ~(layer0_outputs[2094]);
    assign outputs[4919] = ~((layer0_outputs[6517]) | (layer0_outputs[1459]));
    assign outputs[4920] = ~(layer0_outputs[1599]);
    assign outputs[4921] = layer0_outputs[1769];
    assign outputs[4922] = ~((layer0_outputs[7908]) & (layer0_outputs[2226]));
    assign outputs[4923] = layer0_outputs[10044];
    assign outputs[4924] = (layer0_outputs[5449]) ^ (layer0_outputs[10070]);
    assign outputs[4925] = ~(layer0_outputs[4930]) | (layer0_outputs[2845]);
    assign outputs[4926] = (layer0_outputs[2577]) & ~(layer0_outputs[9840]);
    assign outputs[4927] = ~(layer0_outputs[7845]);
    assign outputs[4928] = ~(layer0_outputs[9960]) | (layer0_outputs[1956]);
    assign outputs[4929] = (layer0_outputs[2793]) & ~(layer0_outputs[9884]);
    assign outputs[4930] = (layer0_outputs[6895]) | (layer0_outputs[1771]);
    assign outputs[4931] = layer0_outputs[1548];
    assign outputs[4932] = layer0_outputs[4397];
    assign outputs[4933] = (layer0_outputs[10154]) & ~(layer0_outputs[4935]);
    assign outputs[4934] = ~((layer0_outputs[1100]) | (layer0_outputs[6234]));
    assign outputs[4935] = (layer0_outputs[5844]) ^ (layer0_outputs[7951]);
    assign outputs[4936] = ~((layer0_outputs[9004]) | (layer0_outputs[4381]));
    assign outputs[4937] = ~(layer0_outputs[4472]);
    assign outputs[4938] = ~(layer0_outputs[4111]);
    assign outputs[4939] = ~(layer0_outputs[9947]);
    assign outputs[4940] = (layer0_outputs[5543]) ^ (layer0_outputs[8789]);
    assign outputs[4941] = ~(layer0_outputs[9853]) | (layer0_outputs[4231]);
    assign outputs[4942] = ~(layer0_outputs[8102]);
    assign outputs[4943] = ~((layer0_outputs[3093]) ^ (layer0_outputs[8160]));
    assign outputs[4944] = ~(layer0_outputs[6287]);
    assign outputs[4945] = (layer0_outputs[10184]) & ~(layer0_outputs[9834]);
    assign outputs[4946] = (layer0_outputs[2805]) ^ (layer0_outputs[1810]);
    assign outputs[4947] = layer0_outputs[5534];
    assign outputs[4948] = ~((layer0_outputs[5609]) ^ (layer0_outputs[5558]));
    assign outputs[4949] = ~((layer0_outputs[4775]) ^ (layer0_outputs[6046]));
    assign outputs[4950] = layer0_outputs[6863];
    assign outputs[4951] = layer0_outputs[5964];
    assign outputs[4952] = ~(layer0_outputs[2281]);
    assign outputs[4953] = ~(layer0_outputs[6899]);
    assign outputs[4954] = ~(layer0_outputs[9805]);
    assign outputs[4955] = ~(layer0_outputs[6576]);
    assign outputs[4956] = ~(layer0_outputs[2914]);
    assign outputs[4957] = (layer0_outputs[1299]) & ~(layer0_outputs[8809]);
    assign outputs[4958] = (layer0_outputs[2599]) & ~(layer0_outputs[1278]);
    assign outputs[4959] = layer0_outputs[5720];
    assign outputs[4960] = layer0_outputs[1055];
    assign outputs[4961] = layer0_outputs[4113];
    assign outputs[4962] = ~((layer0_outputs[8407]) ^ (layer0_outputs[8870]));
    assign outputs[4963] = ~(layer0_outputs[4632]);
    assign outputs[4964] = (layer0_outputs[5967]) & (layer0_outputs[5811]);
    assign outputs[4965] = ~((layer0_outputs[4723]) ^ (layer0_outputs[9091]));
    assign outputs[4966] = layer0_outputs[6721];
    assign outputs[4967] = ~(layer0_outputs[3854]);
    assign outputs[4968] = layer0_outputs[6099];
    assign outputs[4969] = (layer0_outputs[6332]) & ~(layer0_outputs[6938]);
    assign outputs[4970] = ~((layer0_outputs[6351]) ^ (layer0_outputs[7371]));
    assign outputs[4971] = ~(layer0_outputs[897]);
    assign outputs[4972] = layer0_outputs[8285];
    assign outputs[4973] = ~(layer0_outputs[5205]);
    assign outputs[4974] = (layer0_outputs[6634]) ^ (layer0_outputs[703]);
    assign outputs[4975] = layer0_outputs[3809];
    assign outputs[4976] = ~(layer0_outputs[1404]);
    assign outputs[4977] = ~(layer0_outputs[7033]);
    assign outputs[4978] = layer0_outputs[3303];
    assign outputs[4979] = ~((layer0_outputs[7447]) | (layer0_outputs[6610]));
    assign outputs[4980] = layer0_outputs[8276];
    assign outputs[4981] = (layer0_outputs[2551]) ^ (layer0_outputs[4017]);
    assign outputs[4982] = (layer0_outputs[5122]) & (layer0_outputs[3452]);
    assign outputs[4983] = (layer0_outputs[4453]) & ~(layer0_outputs[5705]);
    assign outputs[4984] = ~(layer0_outputs[7649]);
    assign outputs[4985] = ~(layer0_outputs[405]);
    assign outputs[4986] = layer0_outputs[2310];
    assign outputs[4987] = (layer0_outputs[2711]) & ~(layer0_outputs[9263]);
    assign outputs[4988] = (layer0_outputs[9617]) & (layer0_outputs[1088]);
    assign outputs[4989] = (layer0_outputs[2453]) | (layer0_outputs[7787]);
    assign outputs[4990] = ~((layer0_outputs[2327]) & (layer0_outputs[488]));
    assign outputs[4991] = layer0_outputs[8905];
    assign outputs[4992] = ~(layer0_outputs[8421]);
    assign outputs[4993] = ~((layer0_outputs[7985]) | (layer0_outputs[3866]));
    assign outputs[4994] = ~(layer0_outputs[7682]);
    assign outputs[4995] = (layer0_outputs[7824]) & (layer0_outputs[4224]);
    assign outputs[4996] = layer0_outputs[876];
    assign outputs[4997] = ~(layer0_outputs[6018]) | (layer0_outputs[6522]);
    assign outputs[4998] = ~((layer0_outputs[5120]) ^ (layer0_outputs[7469]));
    assign outputs[4999] = (layer0_outputs[4598]) & ~(layer0_outputs[2952]);
    assign outputs[5000] = layer0_outputs[4124];
    assign outputs[5001] = ~(layer0_outputs[9664]) | (layer0_outputs[7498]);
    assign outputs[5002] = layer0_outputs[7165];
    assign outputs[5003] = layer0_outputs[232];
    assign outputs[5004] = layer0_outputs[4939];
    assign outputs[5005] = layer0_outputs[9261];
    assign outputs[5006] = layer0_outputs[6154];
    assign outputs[5007] = ~(layer0_outputs[5161]);
    assign outputs[5008] = ~((layer0_outputs[4946]) ^ (layer0_outputs[8712]));
    assign outputs[5009] = layer0_outputs[439];
    assign outputs[5010] = ~((layer0_outputs[6357]) | (layer0_outputs[9156]));
    assign outputs[5011] = ~((layer0_outputs[7531]) ^ (layer0_outputs[5424]));
    assign outputs[5012] = (layer0_outputs[617]) ^ (layer0_outputs[6575]);
    assign outputs[5013] = ~((layer0_outputs[847]) ^ (layer0_outputs[2327]));
    assign outputs[5014] = layer0_outputs[4093];
    assign outputs[5015] = (layer0_outputs[1262]) ^ (layer0_outputs[7216]);
    assign outputs[5016] = layer0_outputs[2635];
    assign outputs[5017] = layer0_outputs[4719];
    assign outputs[5018] = layer0_outputs[6258];
    assign outputs[5019] = ~((layer0_outputs[5197]) ^ (layer0_outputs[9686]));
    assign outputs[5020] = ~(layer0_outputs[3027]);
    assign outputs[5021] = (layer0_outputs[8562]) & ~(layer0_outputs[1973]);
    assign outputs[5022] = layer0_outputs[5832];
    assign outputs[5023] = (layer0_outputs[6502]) & ~(layer0_outputs[5061]);
    assign outputs[5024] = ~((layer0_outputs[6650]) & (layer0_outputs[6088]));
    assign outputs[5025] = ~(layer0_outputs[7688]);
    assign outputs[5026] = (layer0_outputs[666]) ^ (layer0_outputs[9160]);
    assign outputs[5027] = layer0_outputs[3733];
    assign outputs[5028] = ~(layer0_outputs[1201]) | (layer0_outputs[1447]);
    assign outputs[5029] = ~(layer0_outputs[5185]);
    assign outputs[5030] = ~(layer0_outputs[6499]);
    assign outputs[5031] = ~(layer0_outputs[6187]);
    assign outputs[5032] = (layer0_outputs[1606]) | (layer0_outputs[6560]);
    assign outputs[5033] = ~((layer0_outputs[1755]) & (layer0_outputs[1395]));
    assign outputs[5034] = ~((layer0_outputs[5620]) | (layer0_outputs[4983]));
    assign outputs[5035] = ~(layer0_outputs[1805]);
    assign outputs[5036] = ~(layer0_outputs[2240]) | (layer0_outputs[6275]);
    assign outputs[5037] = ~((layer0_outputs[4262]) ^ (layer0_outputs[1930]));
    assign outputs[5038] = ~(layer0_outputs[1510]);
    assign outputs[5039] = layer0_outputs[10223];
    assign outputs[5040] = (layer0_outputs[7422]) & ~(layer0_outputs[8530]);
    assign outputs[5041] = ~(layer0_outputs[4332]);
    assign outputs[5042] = ~(layer0_outputs[1189]);
    assign outputs[5043] = ~(layer0_outputs[1223]);
    assign outputs[5044] = ~(layer0_outputs[10072]);
    assign outputs[5045] = ~(layer0_outputs[5034]) | (layer0_outputs[9950]);
    assign outputs[5046] = ~(layer0_outputs[4303]) | (layer0_outputs[2584]);
    assign outputs[5047] = ~((layer0_outputs[6860]) ^ (layer0_outputs[8935]));
    assign outputs[5048] = (layer0_outputs[3982]) ^ (layer0_outputs[4987]);
    assign outputs[5049] = ~((layer0_outputs[2587]) | (layer0_outputs[4855]));
    assign outputs[5050] = ~(layer0_outputs[7434]);
    assign outputs[5051] = (layer0_outputs[6905]) & ~(layer0_outputs[8218]);
    assign outputs[5052] = layer0_outputs[4037];
    assign outputs[5053] = ~(layer0_outputs[326]) | (layer0_outputs[3404]);
    assign outputs[5054] = ~((layer0_outputs[8385]) ^ (layer0_outputs[6045]));
    assign outputs[5055] = ~((layer0_outputs[3423]) ^ (layer0_outputs[2112]));
    assign outputs[5056] = ~((layer0_outputs[6151]) ^ (layer0_outputs[8828]));
    assign outputs[5057] = (layer0_outputs[8663]) & ~(layer0_outputs[7702]);
    assign outputs[5058] = (layer0_outputs[5201]) ^ (layer0_outputs[4572]);
    assign outputs[5059] = ~(layer0_outputs[2011]) | (layer0_outputs[1412]);
    assign outputs[5060] = layer0_outputs[7596];
    assign outputs[5061] = (layer0_outputs[123]) ^ (layer0_outputs[5326]);
    assign outputs[5062] = layer0_outputs[774];
    assign outputs[5063] = (layer0_outputs[8862]) & (layer0_outputs[7188]);
    assign outputs[5064] = layer0_outputs[2707];
    assign outputs[5065] = ~(layer0_outputs[872]);
    assign outputs[5066] = layer0_outputs[5221];
    assign outputs[5067] = (layer0_outputs[8949]) & ~(layer0_outputs[380]);
    assign outputs[5068] = ~(layer0_outputs[2413]);
    assign outputs[5069] = ~((layer0_outputs[2232]) | (layer0_outputs[7254]));
    assign outputs[5070] = ~((layer0_outputs[9835]) | (layer0_outputs[9147]));
    assign outputs[5071] = ~((layer0_outputs[532]) | (layer0_outputs[5597]));
    assign outputs[5072] = ~(layer0_outputs[2482]) | (layer0_outputs[6601]);
    assign outputs[5073] = ~(layer0_outputs[10015]);
    assign outputs[5074] = ~(layer0_outputs[4564]);
    assign outputs[5075] = ~((layer0_outputs[9992]) | (layer0_outputs[7008]));
    assign outputs[5076] = ~(layer0_outputs[7640]);
    assign outputs[5077] = layer0_outputs[2724];
    assign outputs[5078] = layer0_outputs[5877];
    assign outputs[5079] = ~(layer0_outputs[2625]) | (layer0_outputs[5366]);
    assign outputs[5080] = ~(layer0_outputs[5103]);
    assign outputs[5081] = (layer0_outputs[1877]) | (layer0_outputs[9636]);
    assign outputs[5082] = (layer0_outputs[6432]) ^ (layer0_outputs[10055]);
    assign outputs[5083] = ~(layer0_outputs[6907]);
    assign outputs[5084] = ~((layer0_outputs[6210]) ^ (layer0_outputs[3677]));
    assign outputs[5085] = ~((layer0_outputs[8374]) & (layer0_outputs[4313]));
    assign outputs[5086] = ~((layer0_outputs[4783]) ^ (layer0_outputs[8971]));
    assign outputs[5087] = ~(layer0_outputs[5754]);
    assign outputs[5088] = (layer0_outputs[8544]) & ~(layer0_outputs[9474]);
    assign outputs[5089] = ~((layer0_outputs[1283]) | (layer0_outputs[8619]));
    assign outputs[5090] = ~(layer0_outputs[9530]);
    assign outputs[5091] = layer0_outputs[1272];
    assign outputs[5092] = layer0_outputs[3639];
    assign outputs[5093] = ~(layer0_outputs[2514]);
    assign outputs[5094] = (layer0_outputs[1012]) ^ (layer0_outputs[4977]);
    assign outputs[5095] = layer0_outputs[7029];
    assign outputs[5096] = (layer0_outputs[1500]) & ~(layer0_outputs[5915]);
    assign outputs[5097] = ~((layer0_outputs[165]) ^ (layer0_outputs[920]));
    assign outputs[5098] = layer0_outputs[9518];
    assign outputs[5099] = layer0_outputs[2623];
    assign outputs[5100] = layer0_outputs[7068];
    assign outputs[5101] = ~(layer0_outputs[7271]);
    assign outputs[5102] = layer0_outputs[5913];
    assign outputs[5103] = layer0_outputs[7195];
    assign outputs[5104] = 1'b1;
    assign outputs[5105] = layer0_outputs[7279];
    assign outputs[5106] = ~(layer0_outputs[135]);
    assign outputs[5107] = ~(layer0_outputs[9164]);
    assign outputs[5108] = layer0_outputs[3233];
    assign outputs[5109] = layer0_outputs[4415];
    assign outputs[5110] = (layer0_outputs[3666]) & ~(layer0_outputs[4624]);
    assign outputs[5111] = (layer0_outputs[9729]) ^ (layer0_outputs[466]);
    assign outputs[5112] = (layer0_outputs[338]) & ~(layer0_outputs[7607]);
    assign outputs[5113] = (layer0_outputs[6094]) & (layer0_outputs[1320]);
    assign outputs[5114] = layer0_outputs[4881];
    assign outputs[5115] = ~((layer0_outputs[5269]) ^ (layer0_outputs[4733]));
    assign outputs[5116] = ~((layer0_outputs[292]) | (layer0_outputs[1153]));
    assign outputs[5117] = (layer0_outputs[8800]) | (layer0_outputs[2060]);
    assign outputs[5118] = layer0_outputs[3127];
    assign outputs[5119] = layer0_outputs[10155];
    assign outputs[5120] = ~(layer0_outputs[6365]);
    assign outputs[5121] = (layer0_outputs[127]) ^ (layer0_outputs[7810]);
    assign outputs[5122] = ~((layer0_outputs[9584]) | (layer0_outputs[850]));
    assign outputs[5123] = ~((layer0_outputs[1115]) | (layer0_outputs[8540]));
    assign outputs[5124] = ~((layer0_outputs[8240]) | (layer0_outputs[6719]));
    assign outputs[5125] = layer0_outputs[1564];
    assign outputs[5126] = ~(layer0_outputs[6149]);
    assign outputs[5127] = ~((layer0_outputs[726]) ^ (layer0_outputs[2173]));
    assign outputs[5128] = (layer0_outputs[7560]) ^ (layer0_outputs[2740]);
    assign outputs[5129] = ~(layer0_outputs[8214]);
    assign outputs[5130] = layer0_outputs[7001];
    assign outputs[5131] = (layer0_outputs[5166]) & ~(layer0_outputs[5855]);
    assign outputs[5132] = (layer0_outputs[3518]) & ~(layer0_outputs[4018]);
    assign outputs[5133] = ~((layer0_outputs[6818]) ^ (layer0_outputs[7616]));
    assign outputs[5134] = (layer0_outputs[440]) | (layer0_outputs[8756]);
    assign outputs[5135] = ~((layer0_outputs[1941]) | (layer0_outputs[812]));
    assign outputs[5136] = (layer0_outputs[8152]) & ~(layer0_outputs[8603]);
    assign outputs[5137] = ~((layer0_outputs[39]) ^ (layer0_outputs[1360]));
    assign outputs[5138] = ~((layer0_outputs[2609]) ^ (layer0_outputs[4160]));
    assign outputs[5139] = ~(layer0_outputs[5654]);
    assign outputs[5140] = ~(layer0_outputs[5241]);
    assign outputs[5141] = layer0_outputs[4737];
    assign outputs[5142] = (layer0_outputs[8343]) ^ (layer0_outputs[5571]);
    assign outputs[5143] = layer0_outputs[7407];
    assign outputs[5144] = (layer0_outputs[6775]) & ~(layer0_outputs[8881]);
    assign outputs[5145] = ~(layer0_outputs[5753]) | (layer0_outputs[3022]);
    assign outputs[5146] = ~(layer0_outputs[7910]);
    assign outputs[5147] = ~(layer0_outputs[5997]);
    assign outputs[5148] = (layer0_outputs[1515]) ^ (layer0_outputs[7321]);
    assign outputs[5149] = (layer0_outputs[2049]) & ~(layer0_outputs[6660]);
    assign outputs[5150] = layer0_outputs[3472];
    assign outputs[5151] = ~((layer0_outputs[2649]) ^ (layer0_outputs[2202]));
    assign outputs[5152] = ~((layer0_outputs[8312]) ^ (layer0_outputs[768]));
    assign outputs[5153] = ~((layer0_outputs[4312]) | (layer0_outputs[3686]));
    assign outputs[5154] = ~((layer0_outputs[9663]) ^ (layer0_outputs[1830]));
    assign outputs[5155] = (layer0_outputs[56]) ^ (layer0_outputs[4454]);
    assign outputs[5156] = ~((layer0_outputs[4043]) | (layer0_outputs[5519]));
    assign outputs[5157] = ~(layer0_outputs[1977]);
    assign outputs[5158] = (layer0_outputs[4857]) ^ (layer0_outputs[7821]);
    assign outputs[5159] = (layer0_outputs[2510]) ^ (layer0_outputs[4157]);
    assign outputs[5160] = layer0_outputs[775];
    assign outputs[5161] = ~((layer0_outputs[2102]) ^ (layer0_outputs[6221]));
    assign outputs[5162] = (layer0_outputs[2073]) & (layer0_outputs[9525]);
    assign outputs[5163] = (layer0_outputs[8505]) | (layer0_outputs[304]);
    assign outputs[5164] = layer0_outputs[5888];
    assign outputs[5165] = ~((layer0_outputs[9079]) ^ (layer0_outputs[8896]));
    assign outputs[5166] = layer0_outputs[7205];
    assign outputs[5167] = ~((layer0_outputs[6609]) ^ (layer0_outputs[2041]));
    assign outputs[5168] = (layer0_outputs[270]) ^ (layer0_outputs[1639]);
    assign outputs[5169] = (layer0_outputs[4382]) & ~(layer0_outputs[1415]);
    assign outputs[5170] = (layer0_outputs[9500]) & (layer0_outputs[4797]);
    assign outputs[5171] = ~(layer0_outputs[1178]);
    assign outputs[5172] = ~(layer0_outputs[1931]);
    assign outputs[5173] = layer0_outputs[479];
    assign outputs[5174] = ~(layer0_outputs[756]) | (layer0_outputs[2637]);
    assign outputs[5175] = (layer0_outputs[4858]) & ~(layer0_outputs[57]);
    assign outputs[5176] = layer0_outputs[4148];
    assign outputs[5177] = (layer0_outputs[7435]) ^ (layer0_outputs[3696]);
    assign outputs[5178] = layer0_outputs[9021];
    assign outputs[5179] = layer0_outputs[3434];
    assign outputs[5180] = ~((layer0_outputs[1846]) ^ (layer0_outputs[1757]));
    assign outputs[5181] = (layer0_outputs[8446]) & ~(layer0_outputs[8038]);
    assign outputs[5182] = layer0_outputs[9963];
    assign outputs[5183] = ~(layer0_outputs[5017]);
    assign outputs[5184] = (layer0_outputs[6934]) & ~(layer0_outputs[9543]);
    assign outputs[5185] = layer0_outputs[5411];
    assign outputs[5186] = (layer0_outputs[1838]) | (layer0_outputs[9362]);
    assign outputs[5187] = layer0_outputs[3278];
    assign outputs[5188] = ~((layer0_outputs[8537]) | (layer0_outputs[1600]));
    assign outputs[5189] = ~((layer0_outputs[3071]) | (layer0_outputs[990]));
    assign outputs[5190] = layer0_outputs[6956];
    assign outputs[5191] = ~(layer0_outputs[2871]);
    assign outputs[5192] = (layer0_outputs[8376]) & ~(layer0_outputs[2886]);
    assign outputs[5193] = (layer0_outputs[2833]) ^ (layer0_outputs[6436]);
    assign outputs[5194] = (layer0_outputs[4680]) & ~(layer0_outputs[8546]);
    assign outputs[5195] = ~(layer0_outputs[4105]);
    assign outputs[5196] = (layer0_outputs[3581]) & ~(layer0_outputs[7742]);
    assign outputs[5197] = ~(layer0_outputs[2759]);
    assign outputs[5198] = ~(layer0_outputs[8954]);
    assign outputs[5199] = layer0_outputs[8453];
    assign outputs[5200] = (layer0_outputs[314]) ^ (layer0_outputs[443]);
    assign outputs[5201] = (layer0_outputs[4212]) & (layer0_outputs[8265]);
    assign outputs[5202] = ~((layer0_outputs[2126]) ^ (layer0_outputs[1959]));
    assign outputs[5203] = ~(layer0_outputs[2462]);
    assign outputs[5204] = ~(layer0_outputs[1790]);
    assign outputs[5205] = ~(layer0_outputs[6960]);
    assign outputs[5206] = ~(layer0_outputs[3527]);
    assign outputs[5207] = ~((layer0_outputs[1139]) ^ (layer0_outputs[3464]));
    assign outputs[5208] = (layer0_outputs[7508]) ^ (layer0_outputs[5158]);
    assign outputs[5209] = ~(layer0_outputs[6141]);
    assign outputs[5210] = ~(layer0_outputs[9411]);
    assign outputs[5211] = (layer0_outputs[722]) ^ (layer0_outputs[8181]);
    assign outputs[5212] = layer0_outputs[7657];
    assign outputs[5213] = ~(layer0_outputs[5063]);
    assign outputs[5214] = (layer0_outputs[3628]) ^ (layer0_outputs[9540]);
    assign outputs[5215] = ~(layer0_outputs[9430]);
    assign outputs[5216] = (layer0_outputs[7555]) & ~(layer0_outputs[4720]);
    assign outputs[5217] = (layer0_outputs[8702]) & (layer0_outputs[4244]);
    assign outputs[5218] = (layer0_outputs[6705]) | (layer0_outputs[6409]);
    assign outputs[5219] = 1'b1;
    assign outputs[5220] = ~(layer0_outputs[9644]) | (layer0_outputs[4574]);
    assign outputs[5221] = ~(layer0_outputs[9832]);
    assign outputs[5222] = ~(layer0_outputs[5700]) | (layer0_outputs[7551]);
    assign outputs[5223] = ~((layer0_outputs[497]) | (layer0_outputs[3038]));
    assign outputs[5224] = (layer0_outputs[7409]) ^ (layer0_outputs[2858]);
    assign outputs[5225] = layer0_outputs[3339];
    assign outputs[5226] = ~(layer0_outputs[10045]);
    assign outputs[5227] = ~(layer0_outputs[4610]);
    assign outputs[5228] = ~(layer0_outputs[1752]) | (layer0_outputs[6805]);
    assign outputs[5229] = ~(layer0_outputs[1173]);
    assign outputs[5230] = ~((layer0_outputs[7330]) ^ (layer0_outputs[5202]));
    assign outputs[5231] = layer0_outputs[2005];
    assign outputs[5232] = ~(layer0_outputs[3909]);
    assign outputs[5233] = layer0_outputs[9480];
    assign outputs[5234] = ~((layer0_outputs[9841]) ^ (layer0_outputs[5423]));
    assign outputs[5235] = ~(layer0_outputs[6614]);
    assign outputs[5236] = layer0_outputs[3254];
    assign outputs[5237] = ~(layer0_outputs[4796]) | (layer0_outputs[2714]);
    assign outputs[5238] = ~((layer0_outputs[9590]) & (layer0_outputs[2733]));
    assign outputs[5239] = ~((layer0_outputs[2639]) ^ (layer0_outputs[1756]));
    assign outputs[5240] = ~((layer0_outputs[5092]) ^ (layer0_outputs[6951]));
    assign outputs[5241] = layer0_outputs[9820];
    assign outputs[5242] = layer0_outputs[2023];
    assign outputs[5243] = layer0_outputs[8099];
    assign outputs[5244] = ~(layer0_outputs[6534]);
    assign outputs[5245] = (layer0_outputs[7730]) ^ (layer0_outputs[8425]);
    assign outputs[5246] = ~(layer0_outputs[5189]);
    assign outputs[5247] = (layer0_outputs[5763]) ^ (layer0_outputs[4448]);
    assign outputs[5248] = (layer0_outputs[6529]) & (layer0_outputs[7269]);
    assign outputs[5249] = (layer0_outputs[7205]) ^ (layer0_outputs[1029]);
    assign outputs[5250] = (layer0_outputs[6525]) & ~(layer0_outputs[8518]);
    assign outputs[5251] = ~((layer0_outputs[4420]) ^ (layer0_outputs[4789]));
    assign outputs[5252] = ~(layer0_outputs[6036]);
    assign outputs[5253] = layer0_outputs[8262];
    assign outputs[5254] = layer0_outputs[4499];
    assign outputs[5255] = ~(layer0_outputs[9705]);
    assign outputs[5256] = (layer0_outputs[149]) ^ (layer0_outputs[4071]);
    assign outputs[5257] = ~(layer0_outputs[4749]);
    assign outputs[5258] = ~((layer0_outputs[7582]) ^ (layer0_outputs[1122]));
    assign outputs[5259] = ~((layer0_outputs[90]) ^ (layer0_outputs[10223]));
    assign outputs[5260] = ~(layer0_outputs[2436]);
    assign outputs[5261] = (layer0_outputs[3274]) ^ (layer0_outputs[2742]);
    assign outputs[5262] = (layer0_outputs[2413]) ^ (layer0_outputs[8574]);
    assign outputs[5263] = ~((layer0_outputs[6644]) ^ (layer0_outputs[2274]));
    assign outputs[5264] = ~(layer0_outputs[7260]);
    assign outputs[5265] = ~(layer0_outputs[4379]);
    assign outputs[5266] = ~(layer0_outputs[8418]);
    assign outputs[5267] = layer0_outputs[8582];
    assign outputs[5268] = (layer0_outputs[9099]) & (layer0_outputs[7493]);
    assign outputs[5269] = ~((layer0_outputs[8131]) & (layer0_outputs[784]));
    assign outputs[5270] = layer0_outputs[2610];
    assign outputs[5271] = (layer0_outputs[2362]) & (layer0_outputs[1091]);
    assign outputs[5272] = (layer0_outputs[4625]) ^ (layer0_outputs[5622]);
    assign outputs[5273] = ~((layer0_outputs[8440]) ^ (layer0_outputs[9394]));
    assign outputs[5274] = ~(layer0_outputs[3493]) | (layer0_outputs[7051]);
    assign outputs[5275] = (layer0_outputs[9693]) & ~(layer0_outputs[9022]);
    assign outputs[5276] = (layer0_outputs[5058]) & ~(layer0_outputs[33]);
    assign outputs[5277] = layer0_outputs[5305];
    assign outputs[5278] = (layer0_outputs[6463]) & (layer0_outputs[272]);
    assign outputs[5279] = layer0_outputs[3180];
    assign outputs[5280] = (layer0_outputs[8858]) ^ (layer0_outputs[6308]);
    assign outputs[5281] = ~(layer0_outputs[7952]);
    assign outputs[5282] = (layer0_outputs[7421]) & (layer0_outputs[9197]);
    assign outputs[5283] = layer0_outputs[8736];
    assign outputs[5284] = ~(layer0_outputs[5094]);
    assign outputs[5285] = layer0_outputs[1298];
    assign outputs[5286] = ~((layer0_outputs[119]) ^ (layer0_outputs[5908]));
    assign outputs[5287] = ~(layer0_outputs[8780]);
    assign outputs[5288] = ~((layer0_outputs[3314]) ^ (layer0_outputs[4343]));
    assign outputs[5289] = (layer0_outputs[859]) & (layer0_outputs[660]);
    assign outputs[5290] = ~((layer0_outputs[3164]) | (layer0_outputs[1699]));
    assign outputs[5291] = ~((layer0_outputs[1723]) ^ (layer0_outputs[9907]));
    assign outputs[5292] = ~(layer0_outputs[9659]) | (layer0_outputs[9283]);
    assign outputs[5293] = layer0_outputs[1256];
    assign outputs[5294] = ~(layer0_outputs[4777]);
    assign outputs[5295] = ~(layer0_outputs[3906]) | (layer0_outputs[9442]);
    assign outputs[5296] = ~((layer0_outputs[6880]) ^ (layer0_outputs[4133]));
    assign outputs[5297] = layer0_outputs[3010];
    assign outputs[5298] = ~(layer0_outputs[5998]);
    assign outputs[5299] = ~((layer0_outputs[4900]) ^ (layer0_outputs[5169]));
    assign outputs[5300] = ~((layer0_outputs[7372]) & (layer0_outputs[3307]));
    assign outputs[5301] = layer0_outputs[2146];
    assign outputs[5302] = layer0_outputs[776];
    assign outputs[5303] = layer0_outputs[2591];
    assign outputs[5304] = ~((layer0_outputs[873]) ^ (layer0_outputs[7829]));
    assign outputs[5305] = ~(layer0_outputs[5503]);
    assign outputs[5306] = layer0_outputs[2360];
    assign outputs[5307] = (layer0_outputs[3667]) ^ (layer0_outputs[9954]);
    assign outputs[5308] = (layer0_outputs[4767]) ^ (layer0_outputs[10044]);
    assign outputs[5309] = layer0_outputs[6242];
    assign outputs[5310] = (layer0_outputs[1678]) ^ (layer0_outputs[2013]);
    assign outputs[5311] = ~(layer0_outputs[5761]);
    assign outputs[5312] = (layer0_outputs[5268]) ^ (layer0_outputs[10009]);
    assign outputs[5313] = layer0_outputs[9478];
    assign outputs[5314] = (layer0_outputs[935]) ^ (layer0_outputs[613]);
    assign outputs[5315] = layer0_outputs[4031];
    assign outputs[5316] = ~(layer0_outputs[8289]);
    assign outputs[5317] = ~((layer0_outputs[6271]) ^ (layer0_outputs[3224]));
    assign outputs[5318] = ~((layer0_outputs[1902]) ^ (layer0_outputs[7429]));
    assign outputs[5319] = layer0_outputs[4015];
    assign outputs[5320] = layer0_outputs[5328];
    assign outputs[5321] = ~(layer0_outputs[2854]);
    assign outputs[5322] = ~(layer0_outputs[9892]);
    assign outputs[5323] = layer0_outputs[8835];
    assign outputs[5324] = ~((layer0_outputs[5704]) | (layer0_outputs[8310]));
    assign outputs[5325] = layer0_outputs[9314];
    assign outputs[5326] = (layer0_outputs[43]) ^ (layer0_outputs[5085]);
    assign outputs[5327] = (layer0_outputs[7901]) ^ (layer0_outputs[2246]);
    assign outputs[5328] = layer0_outputs[5867];
    assign outputs[5329] = (layer0_outputs[6917]) ^ (layer0_outputs[9369]);
    assign outputs[5330] = (layer0_outputs[7629]) ^ (layer0_outputs[2914]);
    assign outputs[5331] = ~((layer0_outputs[539]) & (layer0_outputs[5442]));
    assign outputs[5332] = ~(layer0_outputs[3704]);
    assign outputs[5333] = ~((layer0_outputs[4472]) & (layer0_outputs[5506]));
    assign outputs[5334] = ~((layer0_outputs[5989]) ^ (layer0_outputs[5866]));
    assign outputs[5335] = (layer0_outputs[1600]) ^ (layer0_outputs[1028]);
    assign outputs[5336] = (layer0_outputs[2666]) & ~(layer0_outputs[9450]);
    assign outputs[5337] = ~((layer0_outputs[701]) | (layer0_outputs[7639]));
    assign outputs[5338] = (layer0_outputs[8028]) & (layer0_outputs[7518]);
    assign outputs[5339] = layer0_outputs[2420];
    assign outputs[5340] = ~(layer0_outputs[809]);
    assign outputs[5341] = ~(layer0_outputs[2714]);
    assign outputs[5342] = ~(layer0_outputs[5187]);
    assign outputs[5343] = layer0_outputs[5900];
    assign outputs[5344] = (layer0_outputs[2385]) ^ (layer0_outputs[80]);
    assign outputs[5345] = ~(layer0_outputs[7237]);
    assign outputs[5346] = ~(layer0_outputs[5110]);
    assign outputs[5347] = layer0_outputs[7645];
    assign outputs[5348] = ~(layer0_outputs[7267]);
    assign outputs[5349] = (layer0_outputs[7856]) & ~(layer0_outputs[2983]);
    assign outputs[5350] = layer0_outputs[9447];
    assign outputs[5351] = layer0_outputs[8928];
    assign outputs[5352] = ~(layer0_outputs[7615]);
    assign outputs[5353] = ~((layer0_outputs[5419]) ^ (layer0_outputs[4763]));
    assign outputs[5354] = layer0_outputs[6674];
    assign outputs[5355] = ~((layer0_outputs[3693]) | (layer0_outputs[8644]));
    assign outputs[5356] = (layer0_outputs[9218]) & ~(layer0_outputs[8323]);
    assign outputs[5357] = (layer0_outputs[4201]) ^ (layer0_outputs[4992]);
    assign outputs[5358] = layer0_outputs[8633];
    assign outputs[5359] = layer0_outputs[5242];
    assign outputs[5360] = ~((layer0_outputs[5424]) ^ (layer0_outputs[6064]));
    assign outputs[5361] = (layer0_outputs[2884]) ^ (layer0_outputs[8729]);
    assign outputs[5362] = ~(layer0_outputs[4847]);
    assign outputs[5363] = ~((layer0_outputs[7950]) | (layer0_outputs[3048]));
    assign outputs[5364] = ~((layer0_outputs[6240]) ^ (layer0_outputs[5164]));
    assign outputs[5365] = layer0_outputs[7680];
    assign outputs[5366] = (layer0_outputs[9262]) ^ (layer0_outputs[1779]);
    assign outputs[5367] = ~((layer0_outputs[9317]) & (layer0_outputs[8668]));
    assign outputs[5368] = (layer0_outputs[3462]) & ~(layer0_outputs[2162]);
    assign outputs[5369] = layer0_outputs[6745];
    assign outputs[5370] = layer0_outputs[1988];
    assign outputs[5371] = ~(layer0_outputs[4404]);
    assign outputs[5372] = ~((layer0_outputs[9737]) ^ (layer0_outputs[8994]));
    assign outputs[5373] = (layer0_outputs[8007]) | (layer0_outputs[9258]);
    assign outputs[5374] = ~((layer0_outputs[5531]) & (layer0_outputs[9203]));
    assign outputs[5375] = ~(layer0_outputs[8519]);
    assign outputs[5376] = ~((layer0_outputs[9636]) ^ (layer0_outputs[5464]));
    assign outputs[5377] = (layer0_outputs[9945]) ^ (layer0_outputs[4579]);
    assign outputs[5378] = (layer0_outputs[8350]) & (layer0_outputs[7891]);
    assign outputs[5379] = ~((layer0_outputs[5741]) ^ (layer0_outputs[7863]));
    assign outputs[5380] = ~(layer0_outputs[9839]);
    assign outputs[5381] = ~((layer0_outputs[7160]) & (layer0_outputs[3306]));
    assign outputs[5382] = ~(layer0_outputs[9141]);
    assign outputs[5383] = (layer0_outputs[2688]) & ~(layer0_outputs[2871]);
    assign outputs[5384] = ~((layer0_outputs[8128]) ^ (layer0_outputs[6117]));
    assign outputs[5385] = ~(layer0_outputs[631]) | (layer0_outputs[1247]);
    assign outputs[5386] = layer0_outputs[4036];
    assign outputs[5387] = (layer0_outputs[6886]) ^ (layer0_outputs[9061]);
    assign outputs[5388] = ~((layer0_outputs[6167]) ^ (layer0_outputs[3514]));
    assign outputs[5389] = layer0_outputs[6955];
    assign outputs[5390] = ~(layer0_outputs[435]) | (layer0_outputs[3602]);
    assign outputs[5391] = ~((layer0_outputs[6064]) | (layer0_outputs[7517]));
    assign outputs[5392] = ~(layer0_outputs[3394]);
    assign outputs[5393] = ~(layer0_outputs[5432]);
    assign outputs[5394] = ~((layer0_outputs[2130]) ^ (layer0_outputs[437]));
    assign outputs[5395] = ~(layer0_outputs[3003]) | (layer0_outputs[9297]);
    assign outputs[5396] = ~(layer0_outputs[9143]);
    assign outputs[5397] = ~((layer0_outputs[5579]) ^ (layer0_outputs[2092]));
    assign outputs[5398] = layer0_outputs[1832];
    assign outputs[5399] = layer0_outputs[3059];
    assign outputs[5400] = (layer0_outputs[6503]) & ~(layer0_outputs[9167]);
    assign outputs[5401] = (layer0_outputs[7550]) & (layer0_outputs[4242]);
    assign outputs[5402] = layer0_outputs[1596];
    assign outputs[5403] = layer0_outputs[140];
    assign outputs[5404] = ~(layer0_outputs[1586]);
    assign outputs[5405] = ~(layer0_outputs[4658]) | (layer0_outputs[2575]);
    assign outputs[5406] = ~(layer0_outputs[7]);
    assign outputs[5407] = layer0_outputs[2452];
    assign outputs[5408] = (layer0_outputs[8151]) ^ (layer0_outputs[10157]);
    assign outputs[5409] = (layer0_outputs[9946]) ^ (layer0_outputs[8090]);
    assign outputs[5410] = layer0_outputs[7347];
    assign outputs[5411] = ~(layer0_outputs[3560]);
    assign outputs[5412] = (layer0_outputs[4846]) ^ (layer0_outputs[9462]);
    assign outputs[5413] = ~(layer0_outputs[2320]);
    assign outputs[5414] = ~((layer0_outputs[9817]) ^ (layer0_outputs[8476]));
    assign outputs[5415] = ~(layer0_outputs[8148]);
    assign outputs[5416] = (layer0_outputs[7252]) ^ (layer0_outputs[7979]);
    assign outputs[5417] = ~(layer0_outputs[8711]) | (layer0_outputs[1132]);
    assign outputs[5418] = (layer0_outputs[3694]) & (layer0_outputs[7113]);
    assign outputs[5419] = ~((layer0_outputs[457]) ^ (layer0_outputs[7604]));
    assign outputs[5420] = ~(layer0_outputs[2801]);
    assign outputs[5421] = ~((layer0_outputs[7004]) ^ (layer0_outputs[204]));
    assign outputs[5422] = layer0_outputs[10049];
    assign outputs[5423] = ~((layer0_outputs[4501]) ^ (layer0_outputs[2029]));
    assign outputs[5424] = ~(layer0_outputs[289]);
    assign outputs[5425] = ~(layer0_outputs[1819]);
    assign outputs[5426] = (layer0_outputs[8142]) | (layer0_outputs[1087]);
    assign outputs[5427] = ~(layer0_outputs[9863]) | (layer0_outputs[2550]);
    assign outputs[5428] = (layer0_outputs[1705]) ^ (layer0_outputs[8214]);
    assign outputs[5429] = ~((layer0_outputs[9484]) ^ (layer0_outputs[8500]));
    assign outputs[5430] = ~(layer0_outputs[7803]);
    assign outputs[5431] = (layer0_outputs[9776]) ^ (layer0_outputs[8294]);
    assign outputs[5432] = ~(layer0_outputs[7653]);
    assign outputs[5433] = (layer0_outputs[3864]) & ~(layer0_outputs[3720]);
    assign outputs[5434] = ~(layer0_outputs[3596]) | (layer0_outputs[2683]);
    assign outputs[5435] = layer0_outputs[4585];
    assign outputs[5436] = (layer0_outputs[4456]) ^ (layer0_outputs[6903]);
    assign outputs[5437] = ~(layer0_outputs[5747]);
    assign outputs[5438] = ~(layer0_outputs[1859]);
    assign outputs[5439] = (layer0_outputs[8411]) ^ (layer0_outputs[5378]);
    assign outputs[5440] = (layer0_outputs[1082]) ^ (layer0_outputs[2261]);
    assign outputs[5441] = (layer0_outputs[5349]) & (layer0_outputs[4718]);
    assign outputs[5442] = (layer0_outputs[3606]) ^ (layer0_outputs[9012]);
    assign outputs[5443] = layer0_outputs[8547];
    assign outputs[5444] = layer0_outputs[1854];
    assign outputs[5445] = ~(layer0_outputs[9557]);
    assign outputs[5446] = (layer0_outputs[3696]) ^ (layer0_outputs[5581]);
    assign outputs[5447] = layer0_outputs[1430];
    assign outputs[5448] = ~((layer0_outputs[2807]) ^ (layer0_outputs[9899]));
    assign outputs[5449] = (layer0_outputs[7779]) & ~(layer0_outputs[5997]);
    assign outputs[5450] = ~(layer0_outputs[6714]);
    assign outputs[5451] = ~(layer0_outputs[9944]);
    assign outputs[5452] = layer0_outputs[4088];
    assign outputs[5453] = (layer0_outputs[7422]) & ~(layer0_outputs[4961]);
    assign outputs[5454] = ~(layer0_outputs[6135]);
    assign outputs[5455] = layer0_outputs[1086];
    assign outputs[5456] = ~(layer0_outputs[10198]);
    assign outputs[5457] = layer0_outputs[2882];
    assign outputs[5458] = ~((layer0_outputs[4633]) ^ (layer0_outputs[4372]));
    assign outputs[5459] = ~(layer0_outputs[1473]);
    assign outputs[5460] = ~((layer0_outputs[5400]) & (layer0_outputs[436]));
    assign outputs[5461] = layer0_outputs[551];
    assign outputs[5462] = ~(layer0_outputs[9462]);
    assign outputs[5463] = ~(layer0_outputs[6575]) | (layer0_outputs[4115]);
    assign outputs[5464] = layer0_outputs[8538];
    assign outputs[5465] = ~((layer0_outputs[4239]) ^ (layer0_outputs[9557]));
    assign outputs[5466] = ~(layer0_outputs[3040]);
    assign outputs[5467] = ~((layer0_outputs[4348]) ^ (layer0_outputs[7552]));
    assign outputs[5468] = ~((layer0_outputs[8057]) ^ (layer0_outputs[6378]));
    assign outputs[5469] = (layer0_outputs[6726]) & ~(layer0_outputs[3052]);
    assign outputs[5470] = ~(layer0_outputs[365]);
    assign outputs[5471] = (layer0_outputs[9090]) ^ (layer0_outputs[425]);
    assign outputs[5472] = layer0_outputs[1107];
    assign outputs[5473] = ~(layer0_outputs[3566]);
    assign outputs[5474] = ~((layer0_outputs[1810]) ^ (layer0_outputs[1269]));
    assign outputs[5475] = (layer0_outputs[1845]) & ~(layer0_outputs[1572]);
    assign outputs[5476] = (layer0_outputs[2199]) & ~(layer0_outputs[1763]);
    assign outputs[5477] = ~((layer0_outputs[378]) ^ (layer0_outputs[4429]));
    assign outputs[5478] = (layer0_outputs[4674]) ^ (layer0_outputs[4268]);
    assign outputs[5479] = ~((layer0_outputs[8908]) ^ (layer0_outputs[8915]));
    assign outputs[5480] = ~((layer0_outputs[863]) ^ (layer0_outputs[10156]));
    assign outputs[5481] = ~((layer0_outputs[10211]) | (layer0_outputs[6861]));
    assign outputs[5482] = ~((layer0_outputs[2086]) ^ (layer0_outputs[3318]));
    assign outputs[5483] = layer0_outputs[9797];
    assign outputs[5484] = layer0_outputs[6238];
    assign outputs[5485] = layer0_outputs[423];
    assign outputs[5486] = layer0_outputs[7811];
    assign outputs[5487] = ~((layer0_outputs[5808]) ^ (layer0_outputs[1930]));
    assign outputs[5488] = ~((layer0_outputs[3101]) ^ (layer0_outputs[4464]));
    assign outputs[5489] = (layer0_outputs[7185]) ^ (layer0_outputs[4476]);
    assign outputs[5490] = ~(layer0_outputs[888]);
    assign outputs[5491] = ~(layer0_outputs[4439]);
    assign outputs[5492] = (layer0_outputs[5931]) & ~(layer0_outputs[2863]);
    assign outputs[5493] = ~(layer0_outputs[3796]);
    assign outputs[5494] = ~(layer0_outputs[1910]);
    assign outputs[5495] = (layer0_outputs[8330]) ^ (layer0_outputs[9191]);
    assign outputs[5496] = ~(layer0_outputs[6814]);
    assign outputs[5497] = (layer0_outputs[5226]) & ~(layer0_outputs[6196]);
    assign outputs[5498] = layer0_outputs[5846];
    assign outputs[5499] = (layer0_outputs[5114]) | (layer0_outputs[1998]);
    assign outputs[5500] = ~((layer0_outputs[5055]) & (layer0_outputs[271]));
    assign outputs[5501] = ~(layer0_outputs[1748]);
    assign outputs[5502] = (layer0_outputs[6424]) & ~(layer0_outputs[3002]);
    assign outputs[5503] = (layer0_outputs[10024]) ^ (layer0_outputs[810]);
    assign outputs[5504] = ~((layer0_outputs[4649]) ^ (layer0_outputs[755]));
    assign outputs[5505] = (layer0_outputs[1409]) ^ (layer0_outputs[8824]);
    assign outputs[5506] = ~((layer0_outputs[9264]) | (layer0_outputs[6016]));
    assign outputs[5507] = ~(layer0_outputs[4092]);
    assign outputs[5508] = layer0_outputs[1008];
    assign outputs[5509] = ~(layer0_outputs[3673]);
    assign outputs[5510] = (layer0_outputs[3432]) & ~(layer0_outputs[6072]);
    assign outputs[5511] = layer0_outputs[5499];
    assign outputs[5512] = layer0_outputs[1446];
    assign outputs[5513] = (layer0_outputs[3441]) | (layer0_outputs[8758]);
    assign outputs[5514] = (layer0_outputs[6924]) & ~(layer0_outputs[1171]);
    assign outputs[5515] = layer0_outputs[5537];
    assign outputs[5516] = (layer0_outputs[133]) ^ (layer0_outputs[7482]);
    assign outputs[5517] = ~((layer0_outputs[6279]) ^ (layer0_outputs[2377]));
    assign outputs[5518] = ~((layer0_outputs[9810]) | (layer0_outputs[9380]));
    assign outputs[5519] = ~((layer0_outputs[8701]) ^ (layer0_outputs[1984]));
    assign outputs[5520] = layer0_outputs[1334];
    assign outputs[5521] = ~((layer0_outputs[8193]) ^ (layer0_outputs[8896]));
    assign outputs[5522] = ~((layer0_outputs[2580]) ^ (layer0_outputs[9036]));
    assign outputs[5523] = layer0_outputs[1120];
    assign outputs[5524] = ~((layer0_outputs[9198]) | (layer0_outputs[2979]));
    assign outputs[5525] = ~(layer0_outputs[6760]) | (layer0_outputs[9654]);
    assign outputs[5526] = layer0_outputs[10239];
    assign outputs[5527] = (layer0_outputs[1235]) ^ (layer0_outputs[8706]);
    assign outputs[5528] = (layer0_outputs[1235]) ^ (layer0_outputs[4853]);
    assign outputs[5529] = (layer0_outputs[488]) ^ (layer0_outputs[6476]);
    assign outputs[5530] = (layer0_outputs[377]) ^ (layer0_outputs[3272]);
    assign outputs[5531] = ~(layer0_outputs[9070]);
    assign outputs[5532] = ~(layer0_outputs[9393]);
    assign outputs[5533] = layer0_outputs[7776];
    assign outputs[5534] = layer0_outputs[9374];
    assign outputs[5535] = ~(layer0_outputs[3098]);
    assign outputs[5536] = ~(layer0_outputs[9115]);
    assign outputs[5537] = ~(layer0_outputs[1311]) | (layer0_outputs[1581]);
    assign outputs[5538] = ~(layer0_outputs[921]) | (layer0_outputs[3153]);
    assign outputs[5539] = ~(layer0_outputs[7280]);
    assign outputs[5540] = (layer0_outputs[7809]) ^ (layer0_outputs[485]);
    assign outputs[5541] = ~((layer0_outputs[9207]) | (layer0_outputs[9922]));
    assign outputs[5542] = ~(layer0_outputs[10214]);
    assign outputs[5543] = (layer0_outputs[3066]) ^ (layer0_outputs[907]);
    assign outputs[5544] = layer0_outputs[7751];
    assign outputs[5545] = (layer0_outputs[4378]) ^ (layer0_outputs[6940]);
    assign outputs[5546] = ~(layer0_outputs[5080]) | (layer0_outputs[9941]);
    assign outputs[5547] = ~((layer0_outputs[1577]) ^ (layer0_outputs[6936]));
    assign outputs[5548] = ~((layer0_outputs[5929]) | (layer0_outputs[2357]));
    assign outputs[5549] = (layer0_outputs[5152]) & ~(layer0_outputs[675]);
    assign outputs[5550] = (layer0_outputs[1453]) & ~(layer0_outputs[8705]);
    assign outputs[5551] = ~(layer0_outputs[339]) | (layer0_outputs[6471]);
    assign outputs[5552] = ~(layer0_outputs[8241]);
    assign outputs[5553] = ~(layer0_outputs[5623]);
    assign outputs[5554] = ~(layer0_outputs[5342]);
    assign outputs[5555] = (layer0_outputs[8333]) & ~(layer0_outputs[3524]);
    assign outputs[5556] = ~((layer0_outputs[7361]) ^ (layer0_outputs[2822]));
    assign outputs[5557] = ~((layer0_outputs[3312]) ^ (layer0_outputs[7087]));
    assign outputs[5558] = ~(layer0_outputs[3912]);
    assign outputs[5559] = layer0_outputs[7113];
    assign outputs[5560] = ~((layer0_outputs[5566]) ^ (layer0_outputs[6232]));
    assign outputs[5561] = layer0_outputs[2331];
    assign outputs[5562] = (layer0_outputs[146]) ^ (layer0_outputs[8515]);
    assign outputs[5563] = layer0_outputs[8641];
    assign outputs[5564] = ~(layer0_outputs[6968]);
    assign outputs[5565] = ~(layer0_outputs[9444]);
    assign outputs[5566] = layer0_outputs[7578];
    assign outputs[5567] = ~(layer0_outputs[5092]);
    assign outputs[5568] = ~(layer0_outputs[9202]);
    assign outputs[5569] = (layer0_outputs[7510]) & ~(layer0_outputs[1585]);
    assign outputs[5570] = ~((layer0_outputs[3060]) | (layer0_outputs[1366]));
    assign outputs[5571] = layer0_outputs[6185];
    assign outputs[5572] = ~((layer0_outputs[8005]) ^ (layer0_outputs[3632]));
    assign outputs[5573] = (layer0_outputs[7589]) & (layer0_outputs[3091]);
    assign outputs[5574] = ~((layer0_outputs[9186]) ^ (layer0_outputs[1462]));
    assign outputs[5575] = layer0_outputs[2980];
    assign outputs[5576] = ~((layer0_outputs[609]) ^ (layer0_outputs[5717]));
    assign outputs[5577] = ~((layer0_outputs[3400]) ^ (layer0_outputs[8082]));
    assign outputs[5578] = ~(layer0_outputs[7356]);
    assign outputs[5579] = ~(layer0_outputs[4848]);
    assign outputs[5580] = layer0_outputs[3504];
    assign outputs[5581] = (layer0_outputs[1245]) & ~(layer0_outputs[9209]);
    assign outputs[5582] = (layer0_outputs[7456]) & (layer0_outputs[1940]);
    assign outputs[5583] = ~(layer0_outputs[252]) | (layer0_outputs[4853]);
    assign outputs[5584] = layer0_outputs[8645];
    assign outputs[5585] = (layer0_outputs[8400]) ^ (layer0_outputs[7515]);
    assign outputs[5586] = (layer0_outputs[2571]) & ~(layer0_outputs[8781]);
    assign outputs[5587] = (layer0_outputs[6233]) ^ (layer0_outputs[3259]);
    assign outputs[5588] = layer0_outputs[1997];
    assign outputs[5589] = ~(layer0_outputs[2866]);
    assign outputs[5590] = (layer0_outputs[5661]) & ~(layer0_outputs[364]);
    assign outputs[5591] = (layer0_outputs[466]) & (layer0_outputs[5691]);
    assign outputs[5592] = ~((layer0_outputs[4369]) ^ (layer0_outputs[6460]));
    assign outputs[5593] = ~((layer0_outputs[844]) ^ (layer0_outputs[9329]));
    assign outputs[5594] = (layer0_outputs[8507]) ^ (layer0_outputs[1850]);
    assign outputs[5595] = (layer0_outputs[182]) ^ (layer0_outputs[3457]);
    assign outputs[5596] = ~((layer0_outputs[1265]) ^ (layer0_outputs[2167]));
    assign outputs[5597] = (layer0_outputs[6739]) & ~(layer0_outputs[5626]);
    assign outputs[5598] = layer0_outputs[9089];
    assign outputs[5599] = layer0_outputs[1518];
    assign outputs[5600] = ~(layer0_outputs[6391]);
    assign outputs[5601] = (layer0_outputs[1968]) | (layer0_outputs[3167]);
    assign outputs[5602] = layer0_outputs[5801];
    assign outputs[5603] = ~(layer0_outputs[6953]) | (layer0_outputs[9492]);
    assign outputs[5604] = (layer0_outputs[5059]) | (layer0_outputs[5740]);
    assign outputs[5605] = ~((layer0_outputs[3896]) ^ (layer0_outputs[9864]));
    assign outputs[5606] = layer0_outputs[1296];
    assign outputs[5607] = ~(layer0_outputs[6925]) | (layer0_outputs[6039]);
    assign outputs[5608] = layer0_outputs[9940];
    assign outputs[5609] = ~((layer0_outputs[3038]) ^ (layer0_outputs[606]));
    assign outputs[5610] = layer0_outputs[2101];
    assign outputs[5611] = ~((layer0_outputs[22]) & (layer0_outputs[697]));
    assign outputs[5612] = ~((layer0_outputs[10137]) & (layer0_outputs[6844]));
    assign outputs[5613] = ~((layer0_outputs[4767]) ^ (layer0_outputs[754]));
    assign outputs[5614] = layer0_outputs[5425];
    assign outputs[5615] = ~((layer0_outputs[5643]) ^ (layer0_outputs[4116]));
    assign outputs[5616] = layer0_outputs[4076];
    assign outputs[5617] = layer0_outputs[6763];
    assign outputs[5618] = ~((layer0_outputs[9535]) | (layer0_outputs[2118]));
    assign outputs[5619] = ~(layer0_outputs[4606]);
    assign outputs[5620] = ~(layer0_outputs[5904]);
    assign outputs[5621] = (layer0_outputs[2835]) ^ (layer0_outputs[3049]);
    assign outputs[5622] = (layer0_outputs[4371]) & ~(layer0_outputs[8146]);
    assign outputs[5623] = (layer0_outputs[6325]) | (layer0_outputs[4070]);
    assign outputs[5624] = layer0_outputs[9891];
    assign outputs[5625] = ~(layer0_outputs[2553]) | (layer0_outputs[7645]);
    assign outputs[5626] = layer0_outputs[6594];
    assign outputs[5627] = ~(layer0_outputs[8351]) | (layer0_outputs[1432]);
    assign outputs[5628] = layer0_outputs[1330];
    assign outputs[5629] = ~(layer0_outputs[9296]);
    assign outputs[5630] = ~(layer0_outputs[2425]);
    assign outputs[5631] = ~((layer0_outputs[5560]) ^ (layer0_outputs[3109]));
    assign outputs[5632] = ~((layer0_outputs[5864]) ^ (layer0_outputs[4165]));
    assign outputs[5633] = ~((layer0_outputs[8272]) ^ (layer0_outputs[1174]));
    assign outputs[5634] = (layer0_outputs[704]) ^ (layer0_outputs[6194]);
    assign outputs[5635] = ~((layer0_outputs[10158]) ^ (layer0_outputs[4561]));
    assign outputs[5636] = ~((layer0_outputs[5934]) ^ (layer0_outputs[6111]));
    assign outputs[5637] = ~((layer0_outputs[4258]) & (layer0_outputs[4879]));
    assign outputs[5638] = ~((layer0_outputs[4261]) ^ (layer0_outputs[5881]));
    assign outputs[5639] = ~(layer0_outputs[2067]);
    assign outputs[5640] = ~(layer0_outputs[1673]) | (layer0_outputs[73]);
    assign outputs[5641] = ~((layer0_outputs[8167]) ^ (layer0_outputs[6619]));
    assign outputs[5642] = layer0_outputs[5112];
    assign outputs[5643] = ~((layer0_outputs[64]) ^ (layer0_outputs[6193]));
    assign outputs[5644] = (layer0_outputs[2015]) | (layer0_outputs[39]);
    assign outputs[5645] = (layer0_outputs[5427]) ^ (layer0_outputs[3568]);
    assign outputs[5646] = (layer0_outputs[4385]) ^ (layer0_outputs[9016]);
    assign outputs[5647] = ~(layer0_outputs[6911]);
    assign outputs[5648] = ~(layer0_outputs[2963]) | (layer0_outputs[8989]);
    assign outputs[5649] = ~(layer0_outputs[5592]);
    assign outputs[5650] = ~(layer0_outputs[10013]);
    assign outputs[5651] = (layer0_outputs[7364]) & ~(layer0_outputs[5715]);
    assign outputs[5652] = ~((layer0_outputs[565]) ^ (layer0_outputs[3682]));
    assign outputs[5653] = ~(layer0_outputs[9186]);
    assign outputs[5654] = ~((layer0_outputs[8371]) | (layer0_outputs[2069]));
    assign outputs[5655] = (layer0_outputs[3745]) ^ (layer0_outputs[9458]);
    assign outputs[5656] = ~(layer0_outputs[4384]);
    assign outputs[5657] = (layer0_outputs[7270]) ^ (layer0_outputs[4551]);
    assign outputs[5658] = ~(layer0_outputs[7273]);
    assign outputs[5659] = (layer0_outputs[5397]) & ~(layer0_outputs[5117]);
    assign outputs[5660] = ~(layer0_outputs[5375]) | (layer0_outputs[1220]);
    assign outputs[5661] = ~(layer0_outputs[2821]);
    assign outputs[5662] = (layer0_outputs[3236]) & ~(layer0_outputs[133]);
    assign outputs[5663] = ~(layer0_outputs[2192]);
    assign outputs[5664] = ~(layer0_outputs[6056]);
    assign outputs[5665] = (layer0_outputs[9144]) ^ (layer0_outputs[2248]);
    assign outputs[5666] = ~(layer0_outputs[244]);
    assign outputs[5667] = layer0_outputs[9511];
    assign outputs[5668] = layer0_outputs[206];
    assign outputs[5669] = ~((layer0_outputs[7833]) & (layer0_outputs[6390]));
    assign outputs[5670] = ~(layer0_outputs[2935]);
    assign outputs[5671] = (layer0_outputs[3787]) | (layer0_outputs[4786]);
    assign outputs[5672] = ~((layer0_outputs[8432]) ^ (layer0_outputs[9193]));
    assign outputs[5673] = ~(layer0_outputs[3530]);
    assign outputs[5674] = ~(layer0_outputs[8831]);
    assign outputs[5675] = ~(layer0_outputs[6533]);
    assign outputs[5676] = layer0_outputs[6725];
    assign outputs[5677] = (layer0_outputs[4125]) ^ (layer0_outputs[1200]);
    assign outputs[5678] = layer0_outputs[7168];
    assign outputs[5679] = ~(layer0_outputs[1074]);
    assign outputs[5680] = (layer0_outputs[2774]) ^ (layer0_outputs[5073]);
    assign outputs[5681] = (layer0_outputs[6821]) | (layer0_outputs[7314]);
    assign outputs[5682] = ~(layer0_outputs[8185]);
    assign outputs[5683] = (layer0_outputs[9401]) ^ (layer0_outputs[7618]);
    assign outputs[5684] = ~(layer0_outputs[7890]) | (layer0_outputs[7892]);
    assign outputs[5685] = (layer0_outputs[4371]) & (layer0_outputs[4242]);
    assign outputs[5686] = (layer0_outputs[3996]) & ~(layer0_outputs[9173]);
    assign outputs[5687] = ~((layer0_outputs[8913]) ^ (layer0_outputs[9133]));
    assign outputs[5688] = layer0_outputs[5457];
    assign outputs[5689] = (layer0_outputs[5327]) | (layer0_outputs[3942]);
    assign outputs[5690] = ~(layer0_outputs[10218]);
    assign outputs[5691] = (layer0_outputs[4190]) ^ (layer0_outputs[598]);
    assign outputs[5692] = ~((layer0_outputs[6249]) ^ (layer0_outputs[2143]));
    assign outputs[5693] = (layer0_outputs[4412]) ^ (layer0_outputs[4097]);
    assign outputs[5694] = ~((layer0_outputs[934]) | (layer0_outputs[6110]));
    assign outputs[5695] = (layer0_outputs[2414]) ^ (layer0_outputs[736]);
    assign outputs[5696] = ~(layer0_outputs[1725]);
    assign outputs[5697] = layer0_outputs[2724];
    assign outputs[5698] = ~((layer0_outputs[6029]) ^ (layer0_outputs[5370]));
    assign outputs[5699] = (layer0_outputs[9698]) & (layer0_outputs[4757]);
    assign outputs[5700] = (layer0_outputs[5362]) & (layer0_outputs[8411]);
    assign outputs[5701] = ~(layer0_outputs[4631]) | (layer0_outputs[10042]);
    assign outputs[5702] = (layer0_outputs[924]) ^ (layer0_outputs[2159]);
    assign outputs[5703] = ~((layer0_outputs[6858]) | (layer0_outputs[2429]));
    assign outputs[5704] = ~((layer0_outputs[4419]) | (layer0_outputs[988]));
    assign outputs[5705] = ~((layer0_outputs[9365]) ^ (layer0_outputs[3741]));
    assign outputs[5706] = ~(layer0_outputs[3164]);
    assign outputs[5707] = ~((layer0_outputs[9248]) ^ (layer0_outputs[3264]));
    assign outputs[5708] = (layer0_outputs[4498]) ^ (layer0_outputs[7619]);
    assign outputs[5709] = layer0_outputs[3554];
    assign outputs[5710] = (layer0_outputs[1845]) & (layer0_outputs[8910]);
    assign outputs[5711] = (layer0_outputs[7563]) ^ (layer0_outputs[4700]);
    assign outputs[5712] = ~((layer0_outputs[6318]) ^ (layer0_outputs[5611]));
    assign outputs[5713] = ~((layer0_outputs[8664]) ^ (layer0_outputs[2993]));
    assign outputs[5714] = ~(layer0_outputs[9651]);
    assign outputs[5715] = layer0_outputs[4350];
    assign outputs[5716] = ~((layer0_outputs[126]) & (layer0_outputs[950]));
    assign outputs[5717] = ~((layer0_outputs[9422]) ^ (layer0_outputs[839]));
    assign outputs[5718] = ~(layer0_outputs[6208]);
    assign outputs[5719] = (layer0_outputs[2030]) ^ (layer0_outputs[6641]);
    assign outputs[5720] = layer0_outputs[2426];
    assign outputs[5721] = layer0_outputs[2862];
    assign outputs[5722] = (layer0_outputs[943]) & (layer0_outputs[7749]);
    assign outputs[5723] = ~(layer0_outputs[6501]);
    assign outputs[5724] = ~((layer0_outputs[9299]) ^ (layer0_outputs[1442]));
    assign outputs[5725] = ~(layer0_outputs[2876]);
    assign outputs[5726] = layer0_outputs[424];
    assign outputs[5727] = (layer0_outputs[3448]) ^ (layer0_outputs[6423]);
    assign outputs[5728] = (layer0_outputs[2092]) ^ (layer0_outputs[2502]);
    assign outputs[5729] = (layer0_outputs[1754]) | (layer0_outputs[9645]);
    assign outputs[5730] = ~((layer0_outputs[4711]) ^ (layer0_outputs[2887]));
    assign outputs[5731] = (layer0_outputs[8244]) ^ (layer0_outputs[903]);
    assign outputs[5732] = layer0_outputs[5212];
    assign outputs[5733] = ~((layer0_outputs[8178]) | (layer0_outputs[3438]));
    assign outputs[5734] = (layer0_outputs[4554]) & ~(layer0_outputs[5491]);
    assign outputs[5735] = ~((layer0_outputs[1721]) ^ (layer0_outputs[6555]));
    assign outputs[5736] = (layer0_outputs[9527]) & ~(layer0_outputs[4933]);
    assign outputs[5737] = ~(layer0_outputs[7059]) | (layer0_outputs[4807]);
    assign outputs[5738] = 1'b0;
    assign outputs[5739] = layer0_outputs[2372];
    assign outputs[5740] = ~((layer0_outputs[7234]) ^ (layer0_outputs[4950]));
    assign outputs[5741] = ~(layer0_outputs[4207]);
    assign outputs[5742] = ~(layer0_outputs[3687]) | (layer0_outputs[4910]);
    assign outputs[5743] = ~(layer0_outputs[6382]);
    assign outputs[5744] = layer0_outputs[5564];
    assign outputs[5745] = ~(layer0_outputs[10175]);
    assign outputs[5746] = ~(layer0_outputs[5891]) | (layer0_outputs[4018]);
    assign outputs[5747] = (layer0_outputs[9886]) & (layer0_outputs[5861]);
    assign outputs[5748] = layer0_outputs[4515];
    assign outputs[5749] = (layer0_outputs[913]) ^ (layer0_outputs[3054]);
    assign outputs[5750] = layer0_outputs[3103];
    assign outputs[5751] = (layer0_outputs[10139]) ^ (layer0_outputs[9991]);
    assign outputs[5752] = ~(layer0_outputs[8761]);
    assign outputs[5753] = ~((layer0_outputs[7720]) ^ (layer0_outputs[5751]));
    assign outputs[5754] = layer0_outputs[9080];
    assign outputs[5755] = ~((layer0_outputs[9806]) | (layer0_outputs[9783]));
    assign outputs[5756] = layer0_outputs[86];
    assign outputs[5757] = layer0_outputs[1451];
    assign outputs[5758] = ~(layer0_outputs[1050]);
    assign outputs[5759] = ~((layer0_outputs[1504]) ^ (layer0_outputs[962]));
    assign outputs[5760] = layer0_outputs[1507];
    assign outputs[5761] = ~((layer0_outputs[7019]) | (layer0_outputs[8750]));
    assign outputs[5762] = layer0_outputs[1520];
    assign outputs[5763] = (layer0_outputs[10234]) | (layer0_outputs[5578]);
    assign outputs[5764] = ~((layer0_outputs[7844]) ^ (layer0_outputs[1346]));
    assign outputs[5765] = ~((layer0_outputs[2102]) ^ (layer0_outputs[4568]));
    assign outputs[5766] = ~((layer0_outputs[4804]) ^ (layer0_outputs[8820]));
    assign outputs[5767] = ~(layer0_outputs[6437]);
    assign outputs[5768] = layer0_outputs[5591];
    assign outputs[5769] = ~((layer0_outputs[9955]) & (layer0_outputs[4651]));
    assign outputs[5770] = (layer0_outputs[7272]) ^ (layer0_outputs[1585]);
    assign outputs[5771] = layer0_outputs[5215];
    assign outputs[5772] = (layer0_outputs[1270]) ^ (layer0_outputs[7675]);
    assign outputs[5773] = (layer0_outputs[5500]) ^ (layer0_outputs[1440]);
    assign outputs[5774] = (layer0_outputs[1116]) ^ (layer0_outputs[6069]);
    assign outputs[5775] = layer0_outputs[6737];
    assign outputs[5776] = ~(layer0_outputs[6305]);
    assign outputs[5777] = (layer0_outputs[1776]) ^ (layer0_outputs[6800]);
    assign outputs[5778] = ~((layer0_outputs[5381]) ^ (layer0_outputs[653]));
    assign outputs[5779] = layer0_outputs[5448];
    assign outputs[5780] = ~(layer0_outputs[8919]);
    assign outputs[5781] = (layer0_outputs[1978]) ^ (layer0_outputs[8019]);
    assign outputs[5782] = ~((layer0_outputs[6355]) ^ (layer0_outputs[8237]));
    assign outputs[5783] = ~(layer0_outputs[3988]);
    assign outputs[5784] = ~(layer0_outputs[6307]);
    assign outputs[5785] = (layer0_outputs[9460]) | (layer0_outputs[487]);
    assign outputs[5786] = layer0_outputs[5601];
    assign outputs[5787] = layer0_outputs[7392];
    assign outputs[5788] = ~((layer0_outputs[6875]) | (layer0_outputs[546]));
    assign outputs[5789] = layer0_outputs[5215];
    assign outputs[5790] = (layer0_outputs[9012]) ^ (layer0_outputs[1015]);
    assign outputs[5791] = layer0_outputs[2139];
    assign outputs[5792] = (layer0_outputs[8586]) ^ (layer0_outputs[6113]);
    assign outputs[5793] = layer0_outputs[4542];
    assign outputs[5794] = layer0_outputs[1019];
    assign outputs[5795] = ~(layer0_outputs[7203]);
    assign outputs[5796] = (layer0_outputs[9957]) | (layer0_outputs[8094]);
    assign outputs[5797] = layer0_outputs[5657];
    assign outputs[5798] = ~(layer0_outputs[10196]) | (layer0_outputs[9873]);
    assign outputs[5799] = layer0_outputs[2869];
    assign outputs[5800] = ~((layer0_outputs[1534]) & (layer0_outputs[3919]));
    assign outputs[5801] = ~(layer0_outputs[3428]);
    assign outputs[5802] = ~((layer0_outputs[1702]) | (layer0_outputs[2658]));
    assign outputs[5803] = layer0_outputs[4839];
    assign outputs[5804] = (layer0_outputs[7471]) ^ (layer0_outputs[6939]);
    assign outputs[5805] = ~((layer0_outputs[1414]) ^ (layer0_outputs[9751]));
    assign outputs[5806] = ~(layer0_outputs[6786]) | (layer0_outputs[2725]);
    assign outputs[5807] = 1'b1;
    assign outputs[5808] = ~(layer0_outputs[8486]);
    assign outputs[5809] = (layer0_outputs[1571]) ^ (layer0_outputs[3220]);
    assign outputs[5810] = ~(layer0_outputs[7968]);
    assign outputs[5811] = ~((layer0_outputs[1362]) & (layer0_outputs[6862]));
    assign outputs[5812] = ~(layer0_outputs[2566]);
    assign outputs[5813] = layer0_outputs[6193];
    assign outputs[5814] = layer0_outputs[9768];
    assign outputs[5815] = ~((layer0_outputs[1934]) ^ (layer0_outputs[4157]));
    assign outputs[5816] = ~(layer0_outputs[8510]);
    assign outputs[5817] = ~((layer0_outputs[5490]) ^ (layer0_outputs[7028]));
    assign outputs[5818] = layer0_outputs[7067];
    assign outputs[5819] = (layer0_outputs[2034]) & ~(layer0_outputs[2835]);
    assign outputs[5820] = ~(layer0_outputs[8384]);
    assign outputs[5821] = layer0_outputs[9910];
    assign outputs[5822] = (layer0_outputs[8093]) & ~(layer0_outputs[6338]);
    assign outputs[5823] = ~(layer0_outputs[5962]) | (layer0_outputs[7526]);
    assign outputs[5824] = (layer0_outputs[6415]) ^ (layer0_outputs[9043]);
    assign outputs[5825] = layer0_outputs[527];
    assign outputs[5826] = (layer0_outputs[2238]) ^ (layer0_outputs[8072]);
    assign outputs[5827] = (layer0_outputs[8107]) ^ (layer0_outputs[919]);
    assign outputs[5828] = ~((layer0_outputs[4225]) | (layer0_outputs[4126]));
    assign outputs[5829] = ~((layer0_outputs[2389]) & (layer0_outputs[5417]));
    assign outputs[5830] = ~(layer0_outputs[2531]);
    assign outputs[5831] = ~(layer0_outputs[3253]);
    assign outputs[5832] = ~(layer0_outputs[1654]) | (layer0_outputs[7587]);
    assign outputs[5833] = ~((layer0_outputs[7215]) ^ (layer0_outputs[10193]));
    assign outputs[5834] = ~(layer0_outputs[3742]);
    assign outputs[5835] = ~(layer0_outputs[6204]);
    assign outputs[5836] = layer0_outputs[2116];
    assign outputs[5837] = ~((layer0_outputs[6473]) ^ (layer0_outputs[3706]));
    assign outputs[5838] = ~((layer0_outputs[9794]) ^ (layer0_outputs[4974]));
    assign outputs[5839] = ~((layer0_outputs[6120]) ^ (layer0_outputs[2105]));
    assign outputs[5840] = ~((layer0_outputs[8629]) & (layer0_outputs[8211]));
    assign outputs[5841] = ~(layer0_outputs[6441]);
    assign outputs[5842] = (layer0_outputs[3218]) ^ (layer0_outputs[5178]);
    assign outputs[5843] = layer0_outputs[508];
    assign outputs[5844] = (layer0_outputs[5875]) ^ (layer0_outputs[1008]);
    assign outputs[5845] = layer0_outputs[9333];
    assign outputs[5846] = layer0_outputs[6757];
    assign outputs[5847] = layer0_outputs[10200];
    assign outputs[5848] = ~(layer0_outputs[7633]);
    assign outputs[5849] = ~((layer0_outputs[2962]) ^ (layer0_outputs[3475]));
    assign outputs[5850] = (layer0_outputs[4216]) ^ (layer0_outputs[9138]);
    assign outputs[5851] = layer0_outputs[3115];
    assign outputs[5852] = layer0_outputs[2595];
    assign outputs[5853] = ~(layer0_outputs[4082]);
    assign outputs[5854] = ~((layer0_outputs[7861]) ^ (layer0_outputs[5256]));
    assign outputs[5855] = ~((layer0_outputs[7950]) & (layer0_outputs[7014]));
    assign outputs[5856] = layer0_outputs[10082];
    assign outputs[5857] = ~(layer0_outputs[9759]);
    assign outputs[5858] = ~(layer0_outputs[3769]) | (layer0_outputs[8295]);
    assign outputs[5859] = layer0_outputs[7076];
    assign outputs[5860] = layer0_outputs[7335];
    assign outputs[5861] = layer0_outputs[7478];
    assign outputs[5862] = (layer0_outputs[3599]) & (layer0_outputs[6434]);
    assign outputs[5863] = layer0_outputs[6433];
    assign outputs[5864] = (layer0_outputs[7079]) ^ (layer0_outputs[8918]);
    assign outputs[5865] = (layer0_outputs[7103]) ^ (layer0_outputs[4080]);
    assign outputs[5866] = (layer0_outputs[465]) | (layer0_outputs[4582]);
    assign outputs[5867] = (layer0_outputs[9643]) & (layer0_outputs[482]);
    assign outputs[5868] = ~((layer0_outputs[6404]) ^ (layer0_outputs[7197]));
    assign outputs[5869] = (layer0_outputs[4044]) ^ (layer0_outputs[1570]);
    assign outputs[5870] = ~(layer0_outputs[2453]);
    assign outputs[5871] = layer0_outputs[2673];
    assign outputs[5872] = layer0_outputs[838];
    assign outputs[5873] = layer0_outputs[8220];
    assign outputs[5874] = (layer0_outputs[1275]) & (layer0_outputs[3009]);
    assign outputs[5875] = ~(layer0_outputs[1331]);
    assign outputs[5876] = ~(layer0_outputs[9933]);
    assign outputs[5877] = ~((layer0_outputs[3664]) ^ (layer0_outputs[8575]));
    assign outputs[5878] = ~(layer0_outputs[9112]);
    assign outputs[5879] = ~((layer0_outputs[3013]) ^ (layer0_outputs[9242]));
    assign outputs[5880] = ~((layer0_outputs[4921]) ^ (layer0_outputs[9376]));
    assign outputs[5881] = ~((layer0_outputs[4788]) & (layer0_outputs[3316]));
    assign outputs[5882] = layer0_outputs[2509];
    assign outputs[5883] = ~((layer0_outputs[2705]) ^ (layer0_outputs[1765]));
    assign outputs[5884] = ~((layer0_outputs[6241]) ^ (layer0_outputs[5650]));
    assign outputs[5885] = layer0_outputs[6144];
    assign outputs[5886] = ~(layer0_outputs[10140]);
    assign outputs[5887] = ~(layer0_outputs[4896]);
    assign outputs[5888] = ~(layer0_outputs[6582]);
    assign outputs[5889] = ~(layer0_outputs[9316]);
    assign outputs[5890] = layer0_outputs[866];
    assign outputs[5891] = (layer0_outputs[6299]) ^ (layer0_outputs[5974]);
    assign outputs[5892] = layer0_outputs[5053];
    assign outputs[5893] = ~((layer0_outputs[891]) ^ (layer0_outputs[3448]));
    assign outputs[5894] = layer0_outputs[1101];
    assign outputs[5895] = layer0_outputs[8348];
    assign outputs[5896] = ~((layer0_outputs[6847]) ^ (layer0_outputs[8168]));
    assign outputs[5897] = ~(layer0_outputs[8906]);
    assign outputs[5898] = (layer0_outputs[3383]) ^ (layer0_outputs[7110]);
    assign outputs[5899] = ~((layer0_outputs[8144]) ^ (layer0_outputs[7232]));
    assign outputs[5900] = ~(layer0_outputs[5151]) | (layer0_outputs[734]);
    assign outputs[5901] = ~(layer0_outputs[4281]);
    assign outputs[5902] = ~((layer0_outputs[10178]) & (layer0_outputs[6425]));
    assign outputs[5903] = ~(layer0_outputs[4030]);
    assign outputs[5904] = ~(layer0_outputs[4409]);
    assign outputs[5905] = (layer0_outputs[397]) ^ (layer0_outputs[4818]);
    assign outputs[5906] = ~(layer0_outputs[6715]);
    assign outputs[5907] = ~(layer0_outputs[2901]);
    assign outputs[5908] = (layer0_outputs[2518]) ^ (layer0_outputs[686]);
    assign outputs[5909] = (layer0_outputs[4925]) ^ (layer0_outputs[352]);
    assign outputs[5910] = ~(layer0_outputs[3845]);
    assign outputs[5911] = layer0_outputs[6131];
    assign outputs[5912] = ~((layer0_outputs[4345]) ^ (layer0_outputs[3739]));
    assign outputs[5913] = ~((layer0_outputs[4547]) ^ (layer0_outputs[2648]));
    assign outputs[5914] = ~((layer0_outputs[353]) ^ (layer0_outputs[5999]));
    assign outputs[5915] = layer0_outputs[506];
    assign outputs[5916] = (layer0_outputs[5953]) ^ (layer0_outputs[6811]);
    assign outputs[5917] = (layer0_outputs[10228]) & (layer0_outputs[3051]);
    assign outputs[5918] = (layer0_outputs[3625]) | (layer0_outputs[6077]);
    assign outputs[5919] = layer0_outputs[9166];
    assign outputs[5920] = layer0_outputs[1498];
    assign outputs[5921] = ~(layer0_outputs[9944]) | (layer0_outputs[1017]);
    assign outputs[5922] = ~(layer0_outputs[3690]);
    assign outputs[5923] = ~(layer0_outputs[2667]);
    assign outputs[5924] = (layer0_outputs[9667]) & ~(layer0_outputs[869]);
    assign outputs[5925] = ~(layer0_outputs[8695]) | (layer0_outputs[9348]);
    assign outputs[5926] = ~(layer0_outputs[3026]);
    assign outputs[5927] = layer0_outputs[6077];
    assign outputs[5928] = ~(layer0_outputs[7878]);
    assign outputs[5929] = ~((layer0_outputs[7155]) & (layer0_outputs[4214]));
    assign outputs[5930] = ~((layer0_outputs[3415]) ^ (layer0_outputs[3219]));
    assign outputs[5931] = ~(layer0_outputs[3760]);
    assign outputs[5932] = ~(layer0_outputs[6700]);
    assign outputs[5933] = ~(layer0_outputs[1057]);
    assign outputs[5934] = (layer0_outputs[7426]) & ~(layer0_outputs[7489]);
    assign outputs[5935] = layer0_outputs[1564];
    assign outputs[5936] = ~(layer0_outputs[1135]);
    assign outputs[5937] = layer0_outputs[7505];
    assign outputs[5938] = ~((layer0_outputs[9266]) & (layer0_outputs[9674]));
    assign outputs[5939] = layer0_outputs[9216];
    assign outputs[5940] = layer0_outputs[2868];
    assign outputs[5941] = layer0_outputs[9607];
    assign outputs[5942] = layer0_outputs[7790];
    assign outputs[5943] = (layer0_outputs[1105]) | (layer0_outputs[8262]);
    assign outputs[5944] = (layer0_outputs[7769]) ^ (layer0_outputs[7997]);
    assign outputs[5945] = (layer0_outputs[4911]) & (layer0_outputs[937]);
    assign outputs[5946] = (layer0_outputs[4146]) | (layer0_outputs[7773]);
    assign outputs[5947] = layer0_outputs[7063];
    assign outputs[5948] = ~(layer0_outputs[1016]);
    assign outputs[5949] = ~(layer0_outputs[1051]);
    assign outputs[5950] = layer0_outputs[1001];
    assign outputs[5951] = ~(layer0_outputs[262]);
    assign outputs[5952] = layer0_outputs[2971];
    assign outputs[5953] = (layer0_outputs[3134]) ^ (layer0_outputs[7210]);
    assign outputs[5954] = ~((layer0_outputs[157]) ^ (layer0_outputs[3406]));
    assign outputs[5955] = ~(layer0_outputs[7503]);
    assign outputs[5956] = (layer0_outputs[3628]) ^ (layer0_outputs[1036]);
    assign outputs[5957] = ~((layer0_outputs[280]) | (layer0_outputs[3300]));
    assign outputs[5958] = ~((layer0_outputs[8737]) ^ (layer0_outputs[5355]));
    assign outputs[5959] = (layer0_outputs[1892]) & ~(layer0_outputs[9327]);
    assign outputs[5960] = layer0_outputs[1885];
    assign outputs[5961] = ~(layer0_outputs[5413]);
    assign outputs[5962] = ~(layer0_outputs[137]);
    assign outputs[5963] = layer0_outputs[1494];
    assign outputs[5964] = ~(layer0_outputs[8302]) | (layer0_outputs[7660]);
    assign outputs[5965] = ~(layer0_outputs[7050]);
    assign outputs[5966] = ~(layer0_outputs[4538]);
    assign outputs[5967] = ~((layer0_outputs[9018]) ^ (layer0_outputs[8727]));
    assign outputs[5968] = ~((layer0_outputs[6344]) | (layer0_outputs[7241]));
    assign outputs[5969] = layer0_outputs[2793];
    assign outputs[5970] = (layer0_outputs[8136]) ^ (layer0_outputs[4235]);
    assign outputs[5971] = layer0_outputs[2997];
    assign outputs[5972] = layer0_outputs[2820];
    assign outputs[5973] = layer0_outputs[7721];
    assign outputs[5974] = layer0_outputs[5420];
    assign outputs[5975] = (layer0_outputs[7686]) ^ (layer0_outputs[7184]);
    assign outputs[5976] = ~(layer0_outputs[261]);
    assign outputs[5977] = ~(layer0_outputs[1441]) | (layer0_outputs[1423]);
    assign outputs[5978] = (layer0_outputs[454]) ^ (layer0_outputs[145]);
    assign outputs[5979] = ~(layer0_outputs[1350]);
    assign outputs[5980] = ~(layer0_outputs[5551]);
    assign outputs[5981] = (layer0_outputs[6827]) ^ (layer0_outputs[1666]);
    assign outputs[5982] = (layer0_outputs[5876]) ^ (layer0_outputs[464]);
    assign outputs[5983] = ~((layer0_outputs[3468]) & (layer0_outputs[4778]));
    assign outputs[5984] = (layer0_outputs[4017]) ^ (layer0_outputs[8977]);
    assign outputs[5985] = (layer0_outputs[16]) ^ (layer0_outputs[1356]);
    assign outputs[5986] = (layer0_outputs[8650]) ^ (layer0_outputs[3522]);
    assign outputs[5987] = ~(layer0_outputs[1293]);
    assign outputs[5988] = layer0_outputs[4418];
    assign outputs[5989] = ~(layer0_outputs[4545]);
    assign outputs[5990] = ~(layer0_outputs[5489]) | (layer0_outputs[9825]);
    assign outputs[5991] = layer0_outputs[2233];
    assign outputs[5992] = (layer0_outputs[8244]) | (layer0_outputs[9421]);
    assign outputs[5993] = ~(layer0_outputs[8587]) | (layer0_outputs[5923]);
    assign outputs[5994] = ~(layer0_outputs[7271]) | (layer0_outputs[9785]);
    assign outputs[5995] = ~((layer0_outputs[8422]) ^ (layer0_outputs[6105]));
    assign outputs[5996] = (layer0_outputs[4161]) | (layer0_outputs[5272]);
    assign outputs[5997] = ~(layer0_outputs[9593]) | (layer0_outputs[663]);
    assign outputs[5998] = layer0_outputs[7462];
    assign outputs[5999] = (layer0_outputs[6340]) ^ (layer0_outputs[8054]);
    assign outputs[6000] = layer0_outputs[4640];
    assign outputs[6001] = ~(layer0_outputs[6196]);
    assign outputs[6002] = (layer0_outputs[6246]) & (layer0_outputs[7398]);
    assign outputs[6003] = ~(layer0_outputs[8521]);
    assign outputs[6004] = ~(layer0_outputs[5335]);
    assign outputs[6005] = layer0_outputs[7074];
    assign outputs[6006] = (layer0_outputs[8133]) & (layer0_outputs[3022]);
    assign outputs[6007] = ~(layer0_outputs[453]) | (layer0_outputs[3133]);
    assign outputs[6008] = layer0_outputs[6278];
    assign outputs[6009] = ~((layer0_outputs[5048]) ^ (layer0_outputs[8102]));
    assign outputs[6010] = ~(layer0_outputs[3863]);
    assign outputs[6011] = (layer0_outputs[1646]) | (layer0_outputs[3916]);
    assign outputs[6012] = ~(layer0_outputs[8594]);
    assign outputs[6013] = ~(layer0_outputs[77]) | (layer0_outputs[6578]);
    assign outputs[6014] = ~((layer0_outputs[5298]) ^ (layer0_outputs[2691]));
    assign outputs[6015] = ~((layer0_outputs[5368]) ^ (layer0_outputs[9909]));
    assign outputs[6016] = layer0_outputs[679];
    assign outputs[6017] = ~(layer0_outputs[5781]);
    assign outputs[6018] = layer0_outputs[1494];
    assign outputs[6019] = ~(layer0_outputs[5466]) | (layer0_outputs[9403]);
    assign outputs[6020] = (layer0_outputs[494]) | (layer0_outputs[5025]);
    assign outputs[6021] = (layer0_outputs[7278]) & ~(layer0_outputs[2866]);
    assign outputs[6022] = (layer0_outputs[8158]) | (layer0_outputs[1313]);
    assign outputs[6023] = (layer0_outputs[2169]) ^ (layer0_outputs[4473]);
    assign outputs[6024] = (layer0_outputs[2463]) ^ (layer0_outputs[1398]);
    assign outputs[6025] = ~(layer0_outputs[1693]);
    assign outputs[6026] = layer0_outputs[7636];
    assign outputs[6027] = (layer0_outputs[10126]) & (layer0_outputs[588]);
    assign outputs[6028] = ~((layer0_outputs[6810]) ^ (layer0_outputs[3188]));
    assign outputs[6029] = layer0_outputs[3083];
    assign outputs[6030] = (layer0_outputs[4852]) ^ (layer0_outputs[10171]);
    assign outputs[6031] = layer0_outputs[6054];
    assign outputs[6032] = ~(layer0_outputs[4293]) | (layer0_outputs[2653]);
    assign outputs[6033] = (layer0_outputs[2885]) & ~(layer0_outputs[5697]);
    assign outputs[6034] = ~((layer0_outputs[9034]) ^ (layer0_outputs[4265]));
    assign outputs[6035] = (layer0_outputs[1027]) ^ (layer0_outputs[1979]);
    assign outputs[6036] = (layer0_outputs[1034]) | (layer0_outputs[2980]);
    assign outputs[6037] = (layer0_outputs[5035]) ^ (layer0_outputs[8131]);
    assign outputs[6038] = ~(layer0_outputs[9770]);
    assign outputs[6039] = ~(layer0_outputs[5335]);
    assign outputs[6040] = ~((layer0_outputs[693]) | (layer0_outputs[7718]));
    assign outputs[6041] = layer0_outputs[1261];
    assign outputs[6042] = (layer0_outputs[7326]) & ~(layer0_outputs[1733]);
    assign outputs[6043] = ~((layer0_outputs[5247]) ^ (layer0_outputs[9796]));
    assign outputs[6044] = (layer0_outputs[8585]) ^ (layer0_outputs[2356]);
    assign outputs[6045] = layer0_outputs[5327];
    assign outputs[6046] = (layer0_outputs[9708]) ^ (layer0_outputs[9070]);
    assign outputs[6047] = layer0_outputs[9687];
    assign outputs[6048] = ~((layer0_outputs[3954]) ^ (layer0_outputs[4765]));
    assign outputs[6049] = (layer0_outputs[5507]) | (layer0_outputs[7774]);
    assign outputs[6050] = layer0_outputs[8259];
    assign outputs[6051] = ~((layer0_outputs[3723]) ^ (layer0_outputs[3636]));
    assign outputs[6052] = (layer0_outputs[10064]) ^ (layer0_outputs[6422]);
    assign outputs[6053] = ~(layer0_outputs[6375]);
    assign outputs[6054] = ~(layer0_outputs[7404]) | (layer0_outputs[5317]);
    assign outputs[6055] = 1'b1;
    assign outputs[6056] = layer0_outputs[2726];
    assign outputs[6057] = ~(layer0_outputs[1035]);
    assign outputs[6058] = (layer0_outputs[9072]) ^ (layer0_outputs[7128]);
    assign outputs[6059] = (layer0_outputs[5559]) & (layer0_outputs[9797]);
    assign outputs[6060] = ~(layer0_outputs[4247]);
    assign outputs[6061] = ~(layer0_outputs[2928]) | (layer0_outputs[7042]);
    assign outputs[6062] = ~((layer0_outputs[2188]) ^ (layer0_outputs[6215]));
    assign outputs[6063] = ~((layer0_outputs[9388]) | (layer0_outputs[2565]));
    assign outputs[6064] = (layer0_outputs[4899]) & ~(layer0_outputs[7653]);
    assign outputs[6065] = layer0_outputs[3301];
    assign outputs[6066] = layer0_outputs[3123];
    assign outputs[6067] = ~((layer0_outputs[4227]) ^ (layer0_outputs[9986]));
    assign outputs[6068] = layer0_outputs[2662];
    assign outputs[6069] = ~(layer0_outputs[1167]) | (layer0_outputs[6549]);
    assign outputs[6070] = (layer0_outputs[2388]) & (layer0_outputs[9562]);
    assign outputs[6071] = (layer0_outputs[1272]) | (layer0_outputs[4322]);
    assign outputs[6072] = ~((layer0_outputs[4105]) & (layer0_outputs[5555]));
    assign outputs[6073] = layer0_outputs[7467];
    assign outputs[6074] = ~((layer0_outputs[4521]) | (layer0_outputs[6044]));
    assign outputs[6075] = ~(layer0_outputs[4566]);
    assign outputs[6076] = (layer0_outputs[7159]) ^ (layer0_outputs[6718]);
    assign outputs[6077] = layer0_outputs[7631];
    assign outputs[6078] = ~((layer0_outputs[5490]) ^ (layer0_outputs[248]));
    assign outputs[6079] = ~((layer0_outputs[9716]) & (layer0_outputs[8046]));
    assign outputs[6080] = ~(layer0_outputs[4403]);
    assign outputs[6081] = ~((layer0_outputs[9416]) ^ (layer0_outputs[6211]));
    assign outputs[6082] = ~(layer0_outputs[7932]);
    assign outputs[6083] = layer0_outputs[8377];
    assign outputs[6084] = layer0_outputs[8296];
    assign outputs[6085] = (layer0_outputs[8023]) ^ (layer0_outputs[3158]);
    assign outputs[6086] = ~(layer0_outputs[10208]);
    assign outputs[6087] = (layer0_outputs[344]) ^ (layer0_outputs[3161]);
    assign outputs[6088] = (layer0_outputs[5115]) ^ (layer0_outputs[8482]);
    assign outputs[6089] = layer0_outputs[6157];
    assign outputs[6090] = ~(layer0_outputs[9641]);
    assign outputs[6091] = ~(layer0_outputs[7906]);
    assign outputs[6092] = layer0_outputs[2347];
    assign outputs[6093] = ~(layer0_outputs[9353]);
    assign outputs[6094] = ~(layer0_outputs[3659]);
    assign outputs[6095] = ~((layer0_outputs[6041]) ^ (layer0_outputs[8809]));
    assign outputs[6096] = ~((layer0_outputs[375]) ^ (layer0_outputs[494]));
    assign outputs[6097] = ~(layer0_outputs[4746]);
    assign outputs[6098] = layer0_outputs[7608];
    assign outputs[6099] = (layer0_outputs[7413]) ^ (layer0_outputs[8711]);
    assign outputs[6100] = (layer0_outputs[6825]) ^ (layer0_outputs[1060]);
    assign outputs[6101] = layer0_outputs[1277];
    assign outputs[6102] = ~(layer0_outputs[709]);
    assign outputs[6103] = layer0_outputs[5329];
    assign outputs[6104] = ~((layer0_outputs[7120]) ^ (layer0_outputs[3516]));
    assign outputs[6105] = ~((layer0_outputs[3016]) ^ (layer0_outputs[2840]));
    assign outputs[6106] = layer0_outputs[6999];
    assign outputs[6107] = ~(layer0_outputs[5998]);
    assign outputs[6108] = (layer0_outputs[898]) & ~(layer0_outputs[9498]);
    assign outputs[6109] = layer0_outputs[1014];
    assign outputs[6110] = layer0_outputs[8671];
    assign outputs[6111] = ~(layer0_outputs[3773]) | (layer0_outputs[7770]);
    assign outputs[6112] = ~((layer0_outputs[2785]) ^ (layer0_outputs[5745]));
    assign outputs[6113] = ~((layer0_outputs[6338]) ^ (layer0_outputs[1382]));
    assign outputs[6114] = ~(layer0_outputs[5775]) | (layer0_outputs[8669]);
    assign outputs[6115] = ~(layer0_outputs[2803]) | (layer0_outputs[8879]);
    assign outputs[6116] = ~(layer0_outputs[10109]);
    assign outputs[6117] = ~(layer0_outputs[5592]);
    assign outputs[6118] = (layer0_outputs[711]) ^ (layer0_outputs[6188]);
    assign outputs[6119] = ~(layer0_outputs[5383]);
    assign outputs[6120] = layer0_outputs[3461];
    assign outputs[6121] = layer0_outputs[7488];
    assign outputs[6122] = (layer0_outputs[7621]) & (layer0_outputs[5450]);
    assign outputs[6123] = (layer0_outputs[532]) & (layer0_outputs[8130]);
    assign outputs[6124] = ~(layer0_outputs[8361]);
    assign outputs[6125] = layer0_outputs[519];
    assign outputs[6126] = (layer0_outputs[2396]) ^ (layer0_outputs[8219]);
    assign outputs[6127] = ~(layer0_outputs[5894]) | (layer0_outputs[5649]);
    assign outputs[6128] = ~((layer0_outputs[2044]) | (layer0_outputs[9289]));
    assign outputs[6129] = layer0_outputs[9915];
    assign outputs[6130] = ~((layer0_outputs[371]) | (layer0_outputs[9619]));
    assign outputs[6131] = ~(layer0_outputs[502]);
    assign outputs[6132] = ~(layer0_outputs[5600]);
    assign outputs[6133] = (layer0_outputs[8820]) & ~(layer0_outputs[412]);
    assign outputs[6134] = (layer0_outputs[1842]) ^ (layer0_outputs[536]);
    assign outputs[6135] = ~(layer0_outputs[8026]);
    assign outputs[6136] = layer0_outputs[6429];
    assign outputs[6137] = ~(layer0_outputs[128]);
    assign outputs[6138] = (layer0_outputs[7761]) ^ (layer0_outputs[3621]);
    assign outputs[6139] = layer0_outputs[1717];
    assign outputs[6140] = ~(layer0_outputs[9735]);
    assign outputs[6141] = ~((layer0_outputs[322]) ^ (layer0_outputs[368]));
    assign outputs[6142] = ~((layer0_outputs[6548]) ^ (layer0_outputs[4639]));
    assign outputs[6143] = ~(layer0_outputs[4666]);
    assign outputs[6144] = ~(layer0_outputs[3752]);
    assign outputs[6145] = ~(layer0_outputs[3934]);
    assign outputs[6146] = layer0_outputs[2745];
    assign outputs[6147] = ~((layer0_outputs[72]) & (layer0_outputs[4958]));
    assign outputs[6148] = layer0_outputs[504];
    assign outputs[6149] = ~((layer0_outputs[1063]) ^ (layer0_outputs[3090]));
    assign outputs[6150] = ~(layer0_outputs[9349]);
    assign outputs[6151] = ~(layer0_outputs[6956]);
    assign outputs[6152] = ~((layer0_outputs[10090]) ^ (layer0_outputs[7647]));
    assign outputs[6153] = ~(layer0_outputs[2683]);
    assign outputs[6154] = layer0_outputs[3543];
    assign outputs[6155] = ~(layer0_outputs[269]);
    assign outputs[6156] = layer0_outputs[2216];
    assign outputs[6157] = ~((layer0_outputs[7231]) ^ (layer0_outputs[9733]));
    assign outputs[6158] = ~(layer0_outputs[4353]);
    assign outputs[6159] = layer0_outputs[7694];
    assign outputs[6160] = ~(layer0_outputs[5077]);
    assign outputs[6161] = ~(layer0_outputs[161]);
    assign outputs[6162] = ~((layer0_outputs[7417]) & (layer0_outputs[8170]));
    assign outputs[6163] = ~(layer0_outputs[3313]);
    assign outputs[6164] = (layer0_outputs[3340]) & ~(layer0_outputs[6473]);
    assign outputs[6165] = ~(layer0_outputs[4705]) | (layer0_outputs[3813]);
    assign outputs[6166] = layer0_outputs[5854];
    assign outputs[6167] = ~(layer0_outputs[8287]);
    assign outputs[6168] = ~(layer0_outputs[7090]);
    assign outputs[6169] = layer0_outputs[7425];
    assign outputs[6170] = (layer0_outputs[8596]) ^ (layer0_outputs[6843]);
    assign outputs[6171] = ~((layer0_outputs[8800]) | (layer0_outputs[2056]));
    assign outputs[6172] = ~((layer0_outputs[85]) ^ (layer0_outputs[7387]));
    assign outputs[6173] = layer0_outputs[4127];
    assign outputs[6174] = ~(layer0_outputs[6349]);
    assign outputs[6175] = layer0_outputs[555];
    assign outputs[6176] = ~((layer0_outputs[5325]) ^ (layer0_outputs[2027]));
    assign outputs[6177] = layer0_outputs[1386];
    assign outputs[6178] = ~((layer0_outputs[9545]) | (layer0_outputs[1214]));
    assign outputs[6179] = ~((layer0_outputs[5336]) ^ (layer0_outputs[7311]));
    assign outputs[6180] = layer0_outputs[7265];
    assign outputs[6181] = ~(layer0_outputs[5431]);
    assign outputs[6182] = ~(layer0_outputs[3146]);
    assign outputs[6183] = (layer0_outputs[3344]) & ~(layer0_outputs[15]);
    assign outputs[6184] = layer0_outputs[815];
    assign outputs[6185] = ~(layer0_outputs[8269]);
    assign outputs[6186] = layer0_outputs[3975];
    assign outputs[6187] = layer0_outputs[7798];
    assign outputs[6188] = ~(layer0_outputs[9278]);
    assign outputs[6189] = ~((layer0_outputs[866]) & (layer0_outputs[9521]));
    assign outputs[6190] = (layer0_outputs[4750]) & ~(layer0_outputs[9666]);
    assign outputs[6191] = layer0_outputs[4934];
    assign outputs[6192] = ~((layer0_outputs[8216]) ^ (layer0_outputs[2204]));
    assign outputs[6193] = ~((layer0_outputs[2217]) | (layer0_outputs[7503]));
    assign outputs[6194] = (layer0_outputs[4897]) & ~(layer0_outputs[6662]);
    assign outputs[6195] = (layer0_outputs[9345]) ^ (layer0_outputs[7754]);
    assign outputs[6196] = ~(layer0_outputs[3815]);
    assign outputs[6197] = layer0_outputs[9655];
    assign outputs[6198] = ~(layer0_outputs[8203]);
    assign outputs[6199] = layer0_outputs[6656];
    assign outputs[6200] = ~(layer0_outputs[9666]);
    assign outputs[6201] = ~((layer0_outputs[7784]) ^ (layer0_outputs[6235]));
    assign outputs[6202] = (layer0_outputs[3725]) & ~(layer0_outputs[4064]);
    assign outputs[6203] = ~(layer0_outputs[2090]);
    assign outputs[6204] = layer0_outputs[6585];
    assign outputs[6205] = (layer0_outputs[5730]) & ~(layer0_outputs[313]);
    assign outputs[6206] = ~(layer0_outputs[953]);
    assign outputs[6207] = layer0_outputs[3755];
    assign outputs[6208] = (layer0_outputs[6173]) & ~(layer0_outputs[1561]);
    assign outputs[6209] = layer0_outputs[167];
    assign outputs[6210] = (layer0_outputs[4362]) & ~(layer0_outputs[5177]);
    assign outputs[6211] = ~(layer0_outputs[10185]);
    assign outputs[6212] = ~(layer0_outputs[5580]);
    assign outputs[6213] = ~(layer0_outputs[7676]);
    assign outputs[6214] = layer0_outputs[3228];
    assign outputs[6215] = layer0_outputs[4481];
    assign outputs[6216] = ~(layer0_outputs[2951]);
    assign outputs[6217] = layer0_outputs[6219];
    assign outputs[6218] = ~(layer0_outputs[8967]);
    assign outputs[6219] = ~(layer0_outputs[3719]);
    assign outputs[6220] = ~(layer0_outputs[9489]);
    assign outputs[6221] = (layer0_outputs[8814]) ^ (layer0_outputs[6785]);
    assign outputs[6222] = ~(layer0_outputs[2481]) | (layer0_outputs[8402]);
    assign outputs[6223] = (layer0_outputs[5275]) & ~(layer0_outputs[5771]);
    assign outputs[6224] = layer0_outputs[8964];
    assign outputs[6225] = ~(layer0_outputs[9763]);
    assign outputs[6226] = (layer0_outputs[5]) ^ (layer0_outputs[2214]);
    assign outputs[6227] = ~(layer0_outputs[9463]);
    assign outputs[6228] = (layer0_outputs[1821]) & ~(layer0_outputs[567]);
    assign outputs[6229] = ~((layer0_outputs[10138]) | (layer0_outputs[303]));
    assign outputs[6230] = ~(layer0_outputs[6365]);
    assign outputs[6231] = layer0_outputs[5562];
    assign outputs[6232] = ~(layer0_outputs[4193]) | (layer0_outputs[3068]);
    assign outputs[6233] = ~(layer0_outputs[5762]);
    assign outputs[6234] = (layer0_outputs[7994]) & (layer0_outputs[7354]);
    assign outputs[6235] = layer0_outputs[4517];
    assign outputs[6236] = (layer0_outputs[2572]) ^ (layer0_outputs[98]);
    assign outputs[6237] = layer0_outputs[2948];
    assign outputs[6238] = ~((layer0_outputs[5873]) | (layer0_outputs[3484]));
    assign outputs[6239] = (layer0_outputs[6871]) & (layer0_outputs[5754]);
    assign outputs[6240] = layer0_outputs[4974];
    assign outputs[6241] = layer0_outputs[1642];
    assign outputs[6242] = layer0_outputs[7523];
    assign outputs[6243] = ~((layer0_outputs[2721]) | (layer0_outputs[2794]));
    assign outputs[6244] = layer0_outputs[7287];
    assign outputs[6245] = (layer0_outputs[2521]) & ~(layer0_outputs[9332]);
    assign outputs[6246] = ~(layer0_outputs[6456]);
    assign outputs[6247] = ~((layer0_outputs[2217]) & (layer0_outputs[2859]));
    assign outputs[6248] = (layer0_outputs[2343]) & ~(layer0_outputs[6781]);
    assign outputs[6249] = ~(layer0_outputs[7038]);
    assign outputs[6250] = ~((layer0_outputs[9572]) | (layer0_outputs[4622]));
    assign outputs[6251] = ~((layer0_outputs[5988]) ^ (layer0_outputs[713]));
    assign outputs[6252] = ~(layer0_outputs[3893]);
    assign outputs[6253] = layer0_outputs[6739];
    assign outputs[6254] = layer0_outputs[818];
    assign outputs[6255] = layer0_outputs[428];
    assign outputs[6256] = layer0_outputs[6679];
    assign outputs[6257] = ~(layer0_outputs[6897]);
    assign outputs[6258] = ~(layer0_outputs[3012]);
    assign outputs[6259] = (layer0_outputs[253]) ^ (layer0_outputs[5978]);
    assign outputs[6260] = ~(layer0_outputs[3360]);
    assign outputs[6261] = layer0_outputs[6732];
    assign outputs[6262] = ~(layer0_outputs[8404]);
    assign outputs[6263] = ~(layer0_outputs[5726]);
    assign outputs[6264] = (layer0_outputs[7068]) ^ (layer0_outputs[1225]);
    assign outputs[6265] = ~(layer0_outputs[1230]);
    assign outputs[6266] = (layer0_outputs[3455]) ^ (layer0_outputs[1449]);
    assign outputs[6267] = (layer0_outputs[8209]) & ~(layer0_outputs[3510]);
    assign outputs[6268] = layer0_outputs[7742];
    assign outputs[6269] = (layer0_outputs[10144]) & ~(layer0_outputs[2464]);
    assign outputs[6270] = layer0_outputs[5861];
    assign outputs[6271] = ~((layer0_outputs[2843]) ^ (layer0_outputs[9476]));
    assign outputs[6272] = layer0_outputs[7034];
    assign outputs[6273] = (layer0_outputs[4905]) ^ (layer0_outputs[2972]);
    assign outputs[6274] = layer0_outputs[7233];
    assign outputs[6275] = ~(layer0_outputs[7922]);
    assign outputs[6276] = (layer0_outputs[3347]) & ~(layer0_outputs[321]);
    assign outputs[6277] = ~(layer0_outputs[5638]);
    assign outputs[6278] = layer0_outputs[907];
    assign outputs[6279] = ~((layer0_outputs[4628]) | (layer0_outputs[116]));
    assign outputs[6280] = ~(layer0_outputs[6153]);
    assign outputs[6281] = layer0_outputs[9591];
    assign outputs[6282] = 1'b1;
    assign outputs[6283] = (layer0_outputs[3266]) & ~(layer0_outputs[9720]);
    assign outputs[6284] = layer0_outputs[7734];
    assign outputs[6285] = ~(layer0_outputs[3944]) | (layer0_outputs[5298]);
    assign outputs[6286] = ~((layer0_outputs[2213]) ^ (layer0_outputs[9871]));
    assign outputs[6287] = (layer0_outputs[6331]) ^ (layer0_outputs[9920]);
    assign outputs[6288] = ~(layer0_outputs[1626]);
    assign outputs[6289] = (layer0_outputs[4567]) | (layer0_outputs[4691]);
    assign outputs[6290] = layer0_outputs[5386];
    assign outputs[6291] = (layer0_outputs[2538]) & ~(layer0_outputs[6742]);
    assign outputs[6292] = layer0_outputs[6974];
    assign outputs[6293] = ~(layer0_outputs[4906]);
    assign outputs[6294] = ~(layer0_outputs[1439]) | (layer0_outputs[8960]);
    assign outputs[6295] = layer0_outputs[3607];
    assign outputs[6296] = layer0_outputs[4526];
    assign outputs[6297] = (layer0_outputs[8270]) & ~(layer0_outputs[8420]);
    assign outputs[6298] = ~((layer0_outputs[10127]) ^ (layer0_outputs[2382]));
    assign outputs[6299] = ~(layer0_outputs[9933]);
    assign outputs[6300] = layer0_outputs[5786];
    assign outputs[6301] = ~(layer0_outputs[6686]);
    assign outputs[6302] = (layer0_outputs[10101]) & ~(layer0_outputs[3807]);
    assign outputs[6303] = (layer0_outputs[3979]) & ~(layer0_outputs[2024]);
    assign outputs[6304] = ~(layer0_outputs[2790]);
    assign outputs[6305] = (layer0_outputs[9424]) ^ (layer0_outputs[6889]);
    assign outputs[6306] = ~(layer0_outputs[10102]);
    assign outputs[6307] = (layer0_outputs[5379]) & (layer0_outputs[4335]);
    assign outputs[6308] = ~((layer0_outputs[5290]) ^ (layer0_outputs[9862]));
    assign outputs[6309] = layer0_outputs[7005];
    assign outputs[6310] = (layer0_outputs[4532]) & ~(layer0_outputs[10091]);
    assign outputs[6311] = layer0_outputs[8008];
    assign outputs[6312] = ~((layer0_outputs[6564]) ^ (layer0_outputs[5603]));
    assign outputs[6313] = ~(layer0_outputs[4307]);
    assign outputs[6314] = ~((layer0_outputs[7227]) | (layer0_outputs[2973]));
    assign outputs[6315] = layer0_outputs[7259];
    assign outputs[6316] = (layer0_outputs[9005]) ^ (layer0_outputs[2272]);
    assign outputs[6317] = layer0_outputs[1291];
    assign outputs[6318] = (layer0_outputs[803]) & (layer0_outputs[9385]);
    assign outputs[6319] = (layer0_outputs[1913]) | (layer0_outputs[2687]);
    assign outputs[6320] = (layer0_outputs[9300]) | (layer0_outputs[6511]);
    assign outputs[6321] = layer0_outputs[9132];
    assign outputs[6322] = (layer0_outputs[2946]) & ~(layer0_outputs[4546]);
    assign outputs[6323] = (layer0_outputs[3880]) & (layer0_outputs[5806]);
    assign outputs[6324] = ~(layer0_outputs[8238]) | (layer0_outputs[1922]);
    assign outputs[6325] = ~(layer0_outputs[6431]);
    assign outputs[6326] = (layer0_outputs[4795]) & ~(layer0_outputs[3102]);
    assign outputs[6327] = layer0_outputs[6856];
    assign outputs[6328] = ~((layer0_outputs[2284]) | (layer0_outputs[7417]));
    assign outputs[6329] = (layer0_outputs[9623]) | (layer0_outputs[2802]);
    assign outputs[6330] = ~(layer0_outputs[4968]);
    assign outputs[6331] = layer0_outputs[9457];
    assign outputs[6332] = ~(layer0_outputs[3863]);
    assign outputs[6333] = (layer0_outputs[8332]) & ~(layer0_outputs[1147]);
    assign outputs[6334] = ~((layer0_outputs[4798]) | (layer0_outputs[2696]));
    assign outputs[6335] = (layer0_outputs[4989]) ^ (layer0_outputs[4374]);
    assign outputs[6336] = ~(layer0_outputs[9969]);
    assign outputs[6337] = layer0_outputs[2764];
    assign outputs[6338] = ~(layer0_outputs[9411]);
    assign outputs[6339] = layer0_outputs[10209];
    assign outputs[6340] = ~(layer0_outputs[3446]);
    assign outputs[6341] = (layer0_outputs[10237]) | (layer0_outputs[212]);
    assign outputs[6342] = (layer0_outputs[5137]) & (layer0_outputs[9475]);
    assign outputs[6343] = ~(layer0_outputs[967]);
    assign outputs[6344] = layer0_outputs[597];
    assign outputs[6345] = ~(layer0_outputs[8374]);
    assign outputs[6346] = layer0_outputs[7039];
    assign outputs[6347] = layer0_outputs[8553];
    assign outputs[6348] = (layer0_outputs[723]) ^ (layer0_outputs[3608]);
    assign outputs[6349] = ~(layer0_outputs[1212]);
    assign outputs[6350] = layer0_outputs[7998];
    assign outputs[6351] = ~((layer0_outputs[1077]) | (layer0_outputs[8821]));
    assign outputs[6352] = layer0_outputs[204];
    assign outputs[6353] = (layer0_outputs[8699]) ^ (layer0_outputs[2593]);
    assign outputs[6354] = ~(layer0_outputs[1463]) | (layer0_outputs[9918]);
    assign outputs[6355] = layer0_outputs[4647];
    assign outputs[6356] = ~(layer0_outputs[3852]);
    assign outputs[6357] = (layer0_outputs[4812]) ^ (layer0_outputs[2032]);
    assign outputs[6358] = ~(layer0_outputs[2317]);
    assign outputs[6359] = (layer0_outputs[4249]) & ~(layer0_outputs[4960]);
    assign outputs[6360] = layer0_outputs[8947];
    assign outputs[6361] = layer0_outputs[5147];
    assign outputs[6362] = layer0_outputs[7626];
    assign outputs[6363] = layer0_outputs[619];
    assign outputs[6364] = ~(layer0_outputs[10077]);
    assign outputs[6365] = ~(layer0_outputs[3422]);
    assign outputs[6366] = ~(layer0_outputs[5619]) | (layer0_outputs[555]);
    assign outputs[6367] = ~((layer0_outputs[7903]) & (layer0_outputs[8869]));
    assign outputs[6368] = layer0_outputs[2751];
    assign outputs[6369] = ~(layer0_outputs[4927]);
    assign outputs[6370] = ~((layer0_outputs[118]) ^ (layer0_outputs[7341]));
    assign outputs[6371] = (layer0_outputs[7547]) & ~(layer0_outputs[1379]);
    assign outputs[6372] = layer0_outputs[2385];
    assign outputs[6373] = layer0_outputs[3414];
    assign outputs[6374] = ~(layer0_outputs[7258]);
    assign outputs[6375] = (layer0_outputs[6546]) & ~(layer0_outputs[6402]);
    assign outputs[6376] = (layer0_outputs[8309]) ^ (layer0_outputs[6042]);
    assign outputs[6377] = ~((layer0_outputs[5555]) & (layer0_outputs[6709]));
    assign outputs[6378] = layer0_outputs[2863];
    assign outputs[6379] = ~(layer0_outputs[9681]);
    assign outputs[6380] = layer0_outputs[5932];
    assign outputs[6381] = (layer0_outputs[2124]) & ~(layer0_outputs[1756]);
    assign outputs[6382] = layer0_outputs[8063];
    assign outputs[6383] = ~(layer0_outputs[9860]) | (layer0_outputs[4438]);
    assign outputs[6384] = ~(layer0_outputs[492]);
    assign outputs[6385] = ~(layer0_outputs[832]);
    assign outputs[6386] = ~(layer0_outputs[1052]);
    assign outputs[6387] = ~(layer0_outputs[8087]);
    assign outputs[6388] = ~((layer0_outputs[9136]) | (layer0_outputs[5032]));
    assign outputs[6389] = (layer0_outputs[2046]) ^ (layer0_outputs[6780]);
    assign outputs[6390] = ~(layer0_outputs[9649]);
    assign outputs[6391] = (layer0_outputs[1068]) & (layer0_outputs[9798]);
    assign outputs[6392] = ~((layer0_outputs[1409]) ^ (layer0_outputs[8195]));
    assign outputs[6393] = ~(layer0_outputs[492]);
    assign outputs[6394] = layer0_outputs[183];
    assign outputs[6395] = ~(layer0_outputs[3247]) | (layer0_outputs[622]);
    assign outputs[6396] = (layer0_outputs[9]) & ~(layer0_outputs[5048]);
    assign outputs[6397] = layer0_outputs[2498];
    assign outputs[6398] = layer0_outputs[2373];
    assign outputs[6399] = layer0_outputs[652];
    assign outputs[6400] = (layer0_outputs[5944]) & ~(layer0_outputs[1947]);
    assign outputs[6401] = ~((layer0_outputs[3507]) & (layer0_outputs[2247]));
    assign outputs[6402] = ~(layer0_outputs[5965]);
    assign outputs[6403] = layer0_outputs[8161];
    assign outputs[6404] = ~((layer0_outputs[6293]) | (layer0_outputs[8354]));
    assign outputs[6405] = (layer0_outputs[3821]) ^ (layer0_outputs[3036]);
    assign outputs[6406] = ~(layer0_outputs[7045]);
    assign outputs[6407] = layer0_outputs[909];
    assign outputs[6408] = ~(layer0_outputs[5388]) | (layer0_outputs[2791]);
    assign outputs[6409] = ~((layer0_outputs[3278]) ^ (layer0_outputs[4129]));
    assign outputs[6410] = ~(layer0_outputs[7448]);
    assign outputs[6411] = ~(layer0_outputs[5581]);
    assign outputs[6412] = (layer0_outputs[8334]) & ~(layer0_outputs[10162]);
    assign outputs[6413] = ~(layer0_outputs[2140]);
    assign outputs[6414] = (layer0_outputs[8044]) & ~(layer0_outputs[8095]);
    assign outputs[6415] = ~((layer0_outputs[4643]) ^ (layer0_outputs[8114]));
    assign outputs[6416] = (layer0_outputs[6284]) & ~(layer0_outputs[5478]);
    assign outputs[6417] = ~(layer0_outputs[9398]) | (layer0_outputs[4702]);
    assign outputs[6418] = layer0_outputs[2183];
    assign outputs[6419] = ~((layer0_outputs[1318]) ^ (layer0_outputs[5828]));
    assign outputs[6420] = ~(layer0_outputs[6260]);
    assign outputs[6421] = ~(layer0_outputs[7841]);
    assign outputs[6422] = ~(layer0_outputs[4878]);
    assign outputs[6423] = ~(layer0_outputs[2922]);
    assign outputs[6424] = ~(layer0_outputs[4299]);
    assign outputs[6425] = ~((layer0_outputs[3252]) ^ (layer0_outputs[1138]));
    assign outputs[6426] = (layer0_outputs[4516]) & ~(layer0_outputs[6488]);
    assign outputs[6427] = layer0_outputs[648];
    assign outputs[6428] = ~((layer0_outputs[2720]) ^ (layer0_outputs[3711]));
    assign outputs[6429] = ~(layer0_outputs[1288]);
    assign outputs[6430] = layer0_outputs[2186];
    assign outputs[6431] = (layer0_outputs[351]) ^ (layer0_outputs[5640]);
    assign outputs[6432] = layer0_outputs[7842];
    assign outputs[6433] = ~(layer0_outputs[4531]) | (layer0_outputs[813]);
    assign outputs[6434] = ~(layer0_outputs[5283]);
    assign outputs[6435] = layer0_outputs[6616];
    assign outputs[6436] = ~(layer0_outputs[10007]);
    assign outputs[6437] = ~(layer0_outputs[541]);
    assign outputs[6438] = layer0_outputs[1659];
    assign outputs[6439] = ~(layer0_outputs[5143]);
    assign outputs[6440] = ~(layer0_outputs[2856]) | (layer0_outputs[6254]);
    assign outputs[6441] = ~(layer0_outputs[3802]) | (layer0_outputs[1638]);
    assign outputs[6442] = ~(layer0_outputs[9566]);
    assign outputs[6443] = ~(layer0_outputs[287]) | (layer0_outputs[1291]);
    assign outputs[6444] = ~(layer0_outputs[6394]);
    assign outputs[6445] = ~(layer0_outputs[5701]);
    assign outputs[6446] = (layer0_outputs[5210]) & ~(layer0_outputs[9844]);
    assign outputs[6447] = ~(layer0_outputs[2810]);
    assign outputs[6448] = layer0_outputs[325];
    assign outputs[6449] = (layer0_outputs[1560]) ^ (layer0_outputs[2302]);
    assign outputs[6450] = ~(layer0_outputs[4762]) | (layer0_outputs[1054]);
    assign outputs[6451] = ~(layer0_outputs[8488]) | (layer0_outputs[2813]);
    assign outputs[6452] = layer0_outputs[7194];
    assign outputs[6453] = ~((layer0_outputs[1530]) ^ (layer0_outputs[2183]));
    assign outputs[6454] = ~(layer0_outputs[7375]);
    assign outputs[6455] = (layer0_outputs[8676]) | (layer0_outputs[2875]);
    assign outputs[6456] = ~(layer0_outputs[11]);
    assign outputs[6457] = (layer0_outputs[4096]) & (layer0_outputs[3316]);
    assign outputs[6458] = (layer0_outputs[6872]) & ~(layer0_outputs[10118]);
    assign outputs[6459] = ~(layer0_outputs[2569]);
    assign outputs[6460] = (layer0_outputs[7772]) & ~(layer0_outputs[4283]);
    assign outputs[6461] = (layer0_outputs[6085]) ^ (layer0_outputs[3886]);
    assign outputs[6462] = ~(layer0_outputs[224]);
    assign outputs[6463] = (layer0_outputs[6256]) & ~(layer0_outputs[1676]);
    assign outputs[6464] = layer0_outputs[9230];
    assign outputs[6465] = ~(layer0_outputs[8324]);
    assign outputs[6466] = ~((layer0_outputs[5514]) ^ (layer0_outputs[5128]));
    assign outputs[6467] = layer0_outputs[7054];
    assign outputs[6468] = ~(layer0_outputs[1762]) | (layer0_outputs[7864]);
    assign outputs[6469] = (layer0_outputs[2744]) & ~(layer0_outputs[2424]);
    assign outputs[6470] = ~((layer0_outputs[3411]) ^ (layer0_outputs[1038]));
    assign outputs[6471] = (layer0_outputs[6778]) | (layer0_outputs[6747]);
    assign outputs[6472] = ~((layer0_outputs[9692]) | (layer0_outputs[3104]));
    assign outputs[6473] = ~(layer0_outputs[4342]);
    assign outputs[6474] = (layer0_outputs[7767]) | (layer0_outputs[2525]);
    assign outputs[6475] = (layer0_outputs[6536]) & ~(layer0_outputs[10088]);
    assign outputs[6476] = layer0_outputs[6810];
    assign outputs[6477] = layer0_outputs[9760];
    assign outputs[6478] = ~(layer0_outputs[161]);
    assign outputs[6479] = ~(layer0_outputs[1129]);
    assign outputs[6480] = ~((layer0_outputs[3949]) ^ (layer0_outputs[5074]));
    assign outputs[6481] = layer0_outputs[7054];
    assign outputs[6482] = layer0_outputs[1980];
    assign outputs[6483] = (layer0_outputs[7626]) ^ (layer0_outputs[7628]);
    assign outputs[6484] = ~((layer0_outputs[8631]) & (layer0_outputs[4815]));
    assign outputs[6485] = ~(layer0_outputs[9286]) | (layer0_outputs[3839]);
    assign outputs[6486] = layer0_outputs[49];
    assign outputs[6487] = layer0_outputs[3998];
    assign outputs[6488] = layer0_outputs[4028];
    assign outputs[6489] = ~((layer0_outputs[2941]) | (layer0_outputs[1743]));
    assign outputs[6490] = layer0_outputs[5830];
    assign outputs[6491] = (layer0_outputs[4359]) & ~(layer0_outputs[5706]);
    assign outputs[6492] = (layer0_outputs[259]) ^ (layer0_outputs[3936]);
    assign outputs[6493] = ~(layer0_outputs[7606]);
    assign outputs[6494] = (layer0_outputs[3737]) & ~(layer0_outputs[3213]);
    assign outputs[6495] = ~(layer0_outputs[6318]);
    assign outputs[6496] = ~(layer0_outputs[3509]) | (layer0_outputs[10026]);
    assign outputs[6497] = ~((layer0_outputs[8367]) ^ (layer0_outputs[7896]));
    assign outputs[6498] = ~(layer0_outputs[4525]);
    assign outputs[6499] = layer0_outputs[665];
    assign outputs[6500] = layer0_outputs[7764];
    assign outputs[6501] = layer0_outputs[6129];
    assign outputs[6502] = layer0_outputs[53];
    assign outputs[6503] = (layer0_outputs[6011]) & ~(layer0_outputs[8834]);
    assign outputs[6504] = ~(layer0_outputs[7324]);
    assign outputs[6505] = ~(layer0_outputs[6131]);
    assign outputs[6506] = ~((layer0_outputs[5232]) | (layer0_outputs[5408]));
    assign outputs[6507] = ~(layer0_outputs[3215]);
    assign outputs[6508] = ~(layer0_outputs[8899]);
    assign outputs[6509] = (layer0_outputs[6985]) & ~(layer0_outputs[9370]);
    assign outputs[6510] = (layer0_outputs[7367]) ^ (layer0_outputs[8075]);
    assign outputs[6511] = (layer0_outputs[2110]) & (layer0_outputs[4069]);
    assign outputs[6512] = (layer0_outputs[3256]) & ~(layer0_outputs[1959]);
    assign outputs[6513] = ~(layer0_outputs[5464]);
    assign outputs[6514] = (layer0_outputs[1000]) & ~(layer0_outputs[8772]);
    assign outputs[6515] = layer0_outputs[4354];
    assign outputs[6516] = ~(layer0_outputs[7979]);
    assign outputs[6517] = layer0_outputs[8721];
    assign outputs[6518] = ~(layer0_outputs[10063]);
    assign outputs[6519] = layer0_outputs[4670];
    assign outputs[6520] = ~(layer0_outputs[4464]);
    assign outputs[6521] = ~(layer0_outputs[2338]);
    assign outputs[6522] = ~(layer0_outputs[662]);
    assign outputs[6523] = layer0_outputs[2967];
    assign outputs[6524] = ~(layer0_outputs[5512]) | (layer0_outputs[1579]);
    assign outputs[6525] = ~(layer0_outputs[5293]);
    assign outputs[6526] = ~(layer0_outputs[117]);
    assign outputs[6527] = (layer0_outputs[9699]) & ~(layer0_outputs[2075]);
    assign outputs[6528] = (layer0_outputs[8322]) | (layer0_outputs[5429]);
    assign outputs[6529] = (layer0_outputs[3914]) ^ (layer0_outputs[6801]);
    assign outputs[6530] = ~((layer0_outputs[7194]) ^ (layer0_outputs[3772]));
    assign outputs[6531] = layer0_outputs[6413];
    assign outputs[6532] = ~((layer0_outputs[8777]) & (layer0_outputs[2254]));
    assign outputs[6533] = ~(layer0_outputs[4067]);
    assign outputs[6534] = layer0_outputs[8769];
    assign outputs[6535] = layer0_outputs[5090];
    assign outputs[6536] = ~(layer0_outputs[6653]);
    assign outputs[6537] = ~(layer0_outputs[5154]);
    assign outputs[6538] = layer0_outputs[464];
    assign outputs[6539] = ~(layer0_outputs[861]);
    assign outputs[6540] = (layer0_outputs[8069]) & ~(layer0_outputs[2954]);
    assign outputs[6541] = (layer0_outputs[5255]) & (layer0_outputs[406]);
    assign outputs[6542] = ~(layer0_outputs[4656]);
    assign outputs[6543] = layer0_outputs[6846];
    assign outputs[6544] = ~(layer0_outputs[9698]) | (layer0_outputs[7061]);
    assign outputs[6545] = ~(layer0_outputs[7031]);
    assign outputs[6546] = ~(layer0_outputs[8609]);
    assign outputs[6547] = (layer0_outputs[1475]) ^ (layer0_outputs[558]);
    assign outputs[6548] = ~(layer0_outputs[6134]);
    assign outputs[6549] = ~(layer0_outputs[2337]);
    assign outputs[6550] = layer0_outputs[3309];
    assign outputs[6551] = ~(layer0_outputs[6159]);
    assign outputs[6552] = ~((layer0_outputs[7448]) & (layer0_outputs[1310]));
    assign outputs[6553] = ~((layer0_outputs[2479]) & (layer0_outputs[8439]));
    assign outputs[6554] = ~(layer0_outputs[745]);
    assign outputs[6555] = ~(layer0_outputs[2833]);
    assign outputs[6556] = ~(layer0_outputs[9488]);
    assign outputs[6557] = (layer0_outputs[9606]) & (layer0_outputs[8175]);
    assign outputs[6558] = (layer0_outputs[7695]) ^ (layer0_outputs[78]);
    assign outputs[6559] = ~((layer0_outputs[6693]) | (layer0_outputs[4783]));
    assign outputs[6560] = ~(layer0_outputs[5822]) | (layer0_outputs[5221]);
    assign outputs[6561] = (layer0_outputs[2239]) ^ (layer0_outputs[359]);
    assign outputs[6562] = ~(layer0_outputs[7536]);
    assign outputs[6563] = ~(layer0_outputs[9985]);
    assign outputs[6564] = ~(layer0_outputs[3285]);
    assign outputs[6565] = ~(layer0_outputs[6014]);
    assign outputs[6566] = ~(layer0_outputs[7140]);
    assign outputs[6567] = layer0_outputs[3741];
    assign outputs[6568] = ~(layer0_outputs[9972]);
    assign outputs[6569] = (layer0_outputs[10154]) & ~(layer0_outputs[362]);
    assign outputs[6570] = (layer0_outputs[1892]) ^ (layer0_outputs[5625]);
    assign outputs[6571] = ~((layer0_outputs[208]) ^ (layer0_outputs[83]));
    assign outputs[6572] = (layer0_outputs[783]) & ~(layer0_outputs[1136]);
    assign outputs[6573] = ~(layer0_outputs[9899]) | (layer0_outputs[1473]);
    assign outputs[6574] = layer0_outputs[1742];
    assign outputs[6575] = ~(layer0_outputs[10110]);
    assign outputs[6576] = (layer0_outputs[2181]) & ~(layer0_outputs[9436]);
    assign outputs[6577] = layer0_outputs[7199];
    assign outputs[6578] = layer0_outputs[5725];
    assign outputs[6579] = (layer0_outputs[7093]) & ~(layer0_outputs[2194]);
    assign outputs[6580] = (layer0_outputs[6965]) & (layer0_outputs[4771]);
    assign outputs[6581] = ~(layer0_outputs[9943]) | (layer0_outputs[6479]);
    assign outputs[6582] = (layer0_outputs[2478]) ^ (layer0_outputs[512]);
    assign outputs[6583] = ~(layer0_outputs[6674]);
    assign outputs[6584] = ~((layer0_outputs[6501]) ^ (layer0_outputs[107]));
    assign outputs[6585] = ~(layer0_outputs[10102]);
    assign outputs[6586] = ~(layer0_outputs[8486]);
    assign outputs[6587] = layer0_outputs[4301];
    assign outputs[6588] = ~(layer0_outputs[6252]);
    assign outputs[6589] = layer0_outputs[4225];
    assign outputs[6590] = ~(layer0_outputs[1099]);
    assign outputs[6591] = layer0_outputs[7402];
    assign outputs[6592] = layer0_outputs[10111];
    assign outputs[6593] = (layer0_outputs[3359]) & (layer0_outputs[4595]);
    assign outputs[6594] = layer0_outputs[2161];
    assign outputs[6595] = ~((layer0_outputs[3973]) & (layer0_outputs[7186]));
    assign outputs[6596] = layer0_outputs[3045];
    assign outputs[6597] = ~(layer0_outputs[5450]) | (layer0_outputs[7538]);
    assign outputs[6598] = layer0_outputs[5454];
    assign outputs[6599] = layer0_outputs[1773];
    assign outputs[6600] = ~((layer0_outputs[3996]) | (layer0_outputs[8098]));
    assign outputs[6601] = ~(layer0_outputs[192]);
    assign outputs[6602] = ~(layer0_outputs[9290]) | (layer0_outputs[8065]);
    assign outputs[6603] = (layer0_outputs[1854]) & (layer0_outputs[6959]);
    assign outputs[6604] = (layer0_outputs[3295]) & (layer0_outputs[360]);
    assign outputs[6605] = layer0_outputs[8673];
    assign outputs[6606] = layer0_outputs[7319];
    assign outputs[6607] = ~((layer0_outputs[2699]) | (layer0_outputs[7156]));
    assign outputs[6608] = ~((layer0_outputs[5839]) | (layer0_outputs[5687]));
    assign outputs[6609] = (layer0_outputs[5420]) & (layer0_outputs[2415]);
    assign outputs[6610] = (layer0_outputs[1128]) ^ (layer0_outputs[5083]);
    assign outputs[6611] = layer0_outputs[1573];
    assign outputs[6612] = (layer0_outputs[5371]) & (layer0_outputs[124]);
    assign outputs[6613] = layer0_outputs[9915];
    assign outputs[6614] = ~(layer0_outputs[7625]);
    assign outputs[6615] = layer0_outputs[7094];
    assign outputs[6616] = (layer0_outputs[2480]) & (layer0_outputs[3003]);
    assign outputs[6617] = ~(layer0_outputs[9830]);
    assign outputs[6618] = ~((layer0_outputs[722]) | (layer0_outputs[2098]));
    assign outputs[6619] = ~(layer0_outputs[9863]) | (layer0_outputs[6036]);
    assign outputs[6620] = layer0_outputs[8397];
    assign outputs[6621] = layer0_outputs[5231];
    assign outputs[6622] = ~((layer0_outputs[4891]) | (layer0_outputs[6775]));
    assign outputs[6623] = ~(layer0_outputs[7209]);
    assign outputs[6624] = ~((layer0_outputs[5195]) | (layer0_outputs[7639]));
    assign outputs[6625] = layer0_outputs[1736];
    assign outputs[6626] = layer0_outputs[9414];
    assign outputs[6627] = ~(layer0_outputs[2702]);
    assign outputs[6628] = ~(layer0_outputs[2391]);
    assign outputs[6629] = layer0_outputs[8247];
    assign outputs[6630] = ~(layer0_outputs[2250]);
    assign outputs[6631] = (layer0_outputs[1037]) ^ (layer0_outputs[4309]);
    assign outputs[6632] = layer0_outputs[1218];
    assign outputs[6633] = ~(layer0_outputs[3959]);
    assign outputs[6634] = layer0_outputs[9142];
    assign outputs[6635] = ~(layer0_outputs[8382]) | (layer0_outputs[17]);
    assign outputs[6636] = (layer0_outputs[7064]) & (layer0_outputs[4652]);
    assign outputs[6637] = (layer0_outputs[2444]) ^ (layer0_outputs[1614]);
    assign outputs[6638] = ~(layer0_outputs[5009]) | (layer0_outputs[5656]);
    assign outputs[6639] = layer0_outputs[6467];
    assign outputs[6640] = ~(layer0_outputs[390]) | (layer0_outputs[3311]);
    assign outputs[6641] = ~((layer0_outputs[10122]) ^ (layer0_outputs[3070]));
    assign outputs[6642] = ~((layer0_outputs[2339]) | (layer0_outputs[968]));
    assign outputs[6643] = ~(layer0_outputs[5111]) | (layer0_outputs[9418]);
    assign outputs[6644] = (layer0_outputs[2777]) ^ (layer0_outputs[5515]);
    assign outputs[6645] = ~((layer0_outputs[6454]) ^ (layer0_outputs[8636]));
    assign outputs[6646] = layer0_outputs[9765];
    assign outputs[6647] = (layer0_outputs[5086]) ^ (layer0_outputs[557]);
    assign outputs[6648] = layer0_outputs[5161];
    assign outputs[6649] = ~(layer0_outputs[6169]);
    assign outputs[6650] = ~((layer0_outputs[9264]) ^ (layer0_outputs[10186]));
    assign outputs[6651] = ~((layer0_outputs[3600]) | (layer0_outputs[5905]));
    assign outputs[6652] = ~((layer0_outputs[5208]) | (layer0_outputs[7408]));
    assign outputs[6653] = (layer0_outputs[723]) ^ (layer0_outputs[6959]);
    assign outputs[6654] = ~(layer0_outputs[3431]) | (layer0_outputs[765]);
    assign outputs[6655] = layer0_outputs[2059];
    assign outputs[6656] = layer0_outputs[7183];
    assign outputs[6657] = ~(layer0_outputs[7379]);
    assign outputs[6658] = ~(layer0_outputs[1789]);
    assign outputs[6659] = ~((layer0_outputs[9908]) & (layer0_outputs[7691]));
    assign outputs[6660] = layer0_outputs[7491];
    assign outputs[6661] = (layer0_outputs[6898]) & (layer0_outputs[3275]);
    assign outputs[6662] = ~(layer0_outputs[2458]);
    assign outputs[6663] = ~((layer0_outputs[3194]) ^ (layer0_outputs[7509]));
    assign outputs[6664] = layer0_outputs[6973];
    assign outputs[6665] = layer0_outputs[430];
    assign outputs[6666] = ~(layer0_outputs[2856]);
    assign outputs[6667] = ~(layer0_outputs[8191]);
    assign outputs[6668] = layer0_outputs[5013];
    assign outputs[6669] = layer0_outputs[8775];
    assign outputs[6670] = (layer0_outputs[8911]) & ~(layer0_outputs[3667]);
    assign outputs[6671] = (layer0_outputs[1223]) ^ (layer0_outputs[5121]);
    assign outputs[6672] = (layer0_outputs[3617]) & ~(layer0_outputs[4653]);
    assign outputs[6673] = ~(layer0_outputs[4655]);
    assign outputs[6674] = ~((layer0_outputs[4753]) ^ (layer0_outputs[6671]));
    assign outputs[6675] = ~(layer0_outputs[8533]);
    assign outputs[6676] = layer0_outputs[5134];
    assign outputs[6677] = layer0_outputs[4544];
    assign outputs[6678] = ~((layer0_outputs[8509]) | (layer0_outputs[6759]));
    assign outputs[6679] = ~(layer0_outputs[7018]);
    assign outputs[6680] = ~((layer0_outputs[949]) | (layer0_outputs[6032]));
    assign outputs[6681] = ~((layer0_outputs[6571]) | (layer0_outputs[2422]));
    assign outputs[6682] = ~(layer0_outputs[9860]) | (layer0_outputs[6008]);
    assign outputs[6683] = ~((layer0_outputs[7978]) ^ (layer0_outputs[6692]));
    assign outputs[6684] = ~((layer0_outputs[6282]) & (layer0_outputs[9763]));
    assign outputs[6685] = ~(layer0_outputs[5246]) | (layer0_outputs[5848]);
    assign outputs[6686] = ~(layer0_outputs[2820]) | (layer0_outputs[10048]);
    assign outputs[6687] = ~((layer0_outputs[7235]) | (layer0_outputs[8450]));
    assign outputs[6688] = ~(layer0_outputs[5937]);
    assign outputs[6689] = ~(layer0_outputs[5171]);
    assign outputs[6690] = ~(layer0_outputs[7777]);
    assign outputs[6691] = layer0_outputs[629];
    assign outputs[6692] = (layer0_outputs[3592]) & (layer0_outputs[2509]);
    assign outputs[6693] = layer0_outputs[6792];
    assign outputs[6694] = ~(layer0_outputs[8908]);
    assign outputs[6695] = ~((layer0_outputs[4645]) | (layer0_outputs[3890]));
    assign outputs[6696] = (layer0_outputs[5318]) ^ (layer0_outputs[8978]);
    assign outputs[6697] = ~(layer0_outputs[4630]);
    assign outputs[6698] = ~(layer0_outputs[7895]);
    assign outputs[6699] = (layer0_outputs[8706]) | (layer0_outputs[4549]);
    assign outputs[6700] = (layer0_outputs[19]) ^ (layer0_outputs[3228]);
    assign outputs[6701] = layer0_outputs[4451];
    assign outputs[6702] = ~((layer0_outputs[9232]) ^ (layer0_outputs[1052]));
    assign outputs[6703] = ~(layer0_outputs[8205]) | (layer0_outputs[4794]);
    assign outputs[6704] = layer0_outputs[8249];
    assign outputs[6705] = (layer0_outputs[3647]) & ~(layer0_outputs[5121]);
    assign outputs[6706] = layer0_outputs[7221];
    assign outputs[6707] = ~(layer0_outputs[589]);
    assign outputs[6708] = ~((layer0_outputs[6561]) | (layer0_outputs[1548]));
    assign outputs[6709] = layer0_outputs[2225];
    assign outputs[6710] = ~(layer0_outputs[9810]);
    assign outputs[6711] = ~((layer0_outputs[889]) ^ (layer0_outputs[6829]));
    assign outputs[6712] = ~(layer0_outputs[7184]);
    assign outputs[6713] = ~(layer0_outputs[684]);
    assign outputs[6714] = ~(layer0_outputs[4262]);
    assign outputs[6715] = layer0_outputs[4285];
    assign outputs[6716] = layer0_outputs[4928];
    assign outputs[6717] = ~((layer0_outputs[8758]) | (layer0_outputs[6580]));
    assign outputs[6718] = ~(layer0_outputs[5866]) | (layer0_outputs[314]);
    assign outputs[6719] = ~(layer0_outputs[3180]);
    assign outputs[6720] = (layer0_outputs[283]) & ~(layer0_outputs[7556]);
    assign outputs[6721] = layer0_outputs[9786];
    assign outputs[6722] = ~(layer0_outputs[227]);
    assign outputs[6723] = (layer0_outputs[2117]) & ~(layer0_outputs[5724]);
    assign outputs[6724] = layer0_outputs[929];
    assign outputs[6725] = ~(layer0_outputs[5984]);
    assign outputs[6726] = (layer0_outputs[3897]) & ~(layer0_outputs[8708]);
    assign outputs[6727] = layer0_outputs[804];
    assign outputs[6728] = ~(layer0_outputs[9365]);
    assign outputs[6729] = ~((layer0_outputs[8773]) ^ (layer0_outputs[8914]));
    assign outputs[6730] = layer0_outputs[384];
    assign outputs[6731] = ~(layer0_outputs[6633]);
    assign outputs[6732] = (layer0_outputs[2188]) & ~(layer0_outputs[4884]);
    assign outputs[6733] = (layer0_outputs[5647]) | (layer0_outputs[940]);
    assign outputs[6734] = (layer0_outputs[2741]) ^ (layer0_outputs[6]);
    assign outputs[6735] = ~((layer0_outputs[7794]) ^ (layer0_outputs[5737]));
    assign outputs[6736] = ~((layer0_outputs[6824]) ^ (layer0_outputs[8401]));
    assign outputs[6737] = (layer0_outputs[7437]) & ~(layer0_outputs[9603]);
    assign outputs[6738] = ~(layer0_outputs[4649]);
    assign outputs[6739] = ~((layer0_outputs[5012]) | (layer0_outputs[10057]));
    assign outputs[6740] = (layer0_outputs[4110]) & ~(layer0_outputs[6695]);
    assign outputs[6741] = ~(layer0_outputs[3297]);
    assign outputs[6742] = ~(layer0_outputs[1077]);
    assign outputs[6743] = ~(layer0_outputs[7208]);
    assign outputs[6744] = ~(layer0_outputs[74]) | (layer0_outputs[6299]);
    assign outputs[6745] = ~(layer0_outputs[9073]);
    assign outputs[6746] = ~((layer0_outputs[8257]) ^ (layer0_outputs[8278]));
    assign outputs[6747] = (layer0_outputs[7276]) ^ (layer0_outputs[7617]);
    assign outputs[6748] = ~(layer0_outputs[8655]);
    assign outputs[6749] = ~((layer0_outputs[7230]) ^ (layer0_outputs[6332]));
    assign outputs[6750] = ~((layer0_outputs[714]) | (layer0_outputs[10050]));
    assign outputs[6751] = (layer0_outputs[10081]) & (layer0_outputs[1090]);
    assign outputs[6752] = ~((layer0_outputs[4401]) & (layer0_outputs[9256]));
    assign outputs[6753] = layer0_outputs[450];
    assign outputs[6754] = ~((layer0_outputs[4188]) ^ (layer0_outputs[5301]));
    assign outputs[6755] = ~((layer0_outputs[3826]) & (layer0_outputs[4058]));
    assign outputs[6756] = (layer0_outputs[6191]) & ~(layer0_outputs[9914]);
    assign outputs[6757] = ~(layer0_outputs[115]) | (layer0_outputs[9769]);
    assign outputs[6758] = (layer0_outputs[4829]) ^ (layer0_outputs[4229]);
    assign outputs[6759] = layer0_outputs[8884];
    assign outputs[6760] = (layer0_outputs[8388]) & ~(layer0_outputs[1645]);
    assign outputs[6761] = (layer0_outputs[3148]) & ~(layer0_outputs[3336]);
    assign outputs[6762] = ~((layer0_outputs[2236]) | (layer0_outputs[6896]));
    assign outputs[6763] = layer0_outputs[482];
    assign outputs[6764] = ~((layer0_outputs[9015]) & (layer0_outputs[661]));
    assign outputs[6765] = ~(layer0_outputs[6507]);
    assign outputs[6766] = ~((layer0_outputs[3613]) | (layer0_outputs[9276]));
    assign outputs[6767] = ~((layer0_outputs[6692]) ^ (layer0_outputs[4873]));
    assign outputs[6768] = ~(layer0_outputs[3689]);
    assign outputs[6769] = ~(layer0_outputs[7258]);
    assign outputs[6770] = ~((layer0_outputs[2817]) | (layer0_outputs[2853]));
    assign outputs[6771] = ~(layer0_outputs[2020]);
    assign outputs[6772] = ~((layer0_outputs[8542]) ^ (layer0_outputs[5167]));
    assign outputs[6773] = ~(layer0_outputs[5831]);
    assign outputs[6774] = ~(layer0_outputs[6456]);
    assign outputs[6775] = ~((layer0_outputs[8652]) | (layer0_outputs[5569]));
    assign outputs[6776] = (layer0_outputs[5392]) & (layer0_outputs[6251]);
    assign outputs[6777] = (layer0_outputs[4713]) ^ (layer0_outputs[7591]);
    assign outputs[6778] = ~(layer0_outputs[3757]) | (layer0_outputs[2310]);
    assign outputs[6779] = ~(layer0_outputs[4063]) | (layer0_outputs[6556]);
    assign outputs[6780] = ~(layer0_outputs[7159]);
    assign outputs[6781] = layer0_outputs[9760];
    assign outputs[6782] = layer0_outputs[2751];
    assign outputs[6783] = layer0_outputs[6231];
    assign outputs[6784] = (layer0_outputs[7309]) & ~(layer0_outputs[824]);
    assign outputs[6785] = (layer0_outputs[3635]) | (layer0_outputs[4561]);
    assign outputs[6786] = ~(layer0_outputs[5390]);
    assign outputs[6787] = ~((layer0_outputs[1111]) ^ (layer0_outputs[8005]));
    assign outputs[6788] = ~((layer0_outputs[1156]) & (layer0_outputs[6619]));
    assign outputs[6789] = layer0_outputs[3172];
    assign outputs[6790] = (layer0_outputs[9108]) & (layer0_outputs[4110]);
    assign outputs[6791] = ~(layer0_outputs[7020]);
    assign outputs[6792] = layer0_outputs[3072];
    assign outputs[6793] = layer0_outputs[9600];
    assign outputs[6794] = ~((layer0_outputs[7322]) & (layer0_outputs[1372]));
    assign outputs[6795] = ~(layer0_outputs[2438]);
    assign outputs[6796] = ~(layer0_outputs[3457]);
    assign outputs[6797] = ~(layer0_outputs[4011]) | (layer0_outputs[1961]);
    assign outputs[6798] = ~(layer0_outputs[8615]);
    assign outputs[6799] = layer0_outputs[10160];
    assign outputs[6800] = (layer0_outputs[7938]) ^ (layer0_outputs[4985]);
    assign outputs[6801] = (layer0_outputs[566]) & (layer0_outputs[6298]);
    assign outputs[6802] = layer0_outputs[6717];
    assign outputs[6803] = ~((layer0_outputs[6844]) & (layer0_outputs[5802]));
    assign outputs[6804] = ~(layer0_outputs[5823]);
    assign outputs[6805] = layer0_outputs[8830];
    assign outputs[6806] = ~((layer0_outputs[5863]) ^ (layer0_outputs[4636]));
    assign outputs[6807] = layer0_outputs[554];
    assign outputs[6808] = ~((layer0_outputs[9487]) | (layer0_outputs[5328]));
    assign outputs[6809] = (layer0_outputs[8864]) ^ (layer0_outputs[4985]);
    assign outputs[6810] = layer0_outputs[8088];
    assign outputs[6811] = ~((layer0_outputs[8141]) | (layer0_outputs[3044]));
    assign outputs[6812] = layer0_outputs[8672];
    assign outputs[6813] = ~((layer0_outputs[567]) | (layer0_outputs[8237]));
    assign outputs[6814] = (layer0_outputs[4959]) & ~(layer0_outputs[7257]);
    assign outputs[6815] = (layer0_outputs[365]) ^ (layer0_outputs[9227]);
    assign outputs[6816] = (layer0_outputs[1352]) ^ (layer0_outputs[7978]);
    assign outputs[6817] = (layer0_outputs[7548]) ^ (layer0_outputs[938]);
    assign outputs[6818] = layer0_outputs[7689];
    assign outputs[6819] = ~(layer0_outputs[1407]);
    assign outputs[6820] = (layer0_outputs[627]) ^ (layer0_outputs[4492]);
    assign outputs[6821] = ~((layer0_outputs[6688]) & (layer0_outputs[6112]));
    assign outputs[6822] = ~((layer0_outputs[2050]) & (layer0_outputs[4305]));
    assign outputs[6823] = ~(layer0_outputs[2710]);
    assign outputs[6824] = ~((layer0_outputs[3832]) | (layer0_outputs[1233]));
    assign outputs[6825] = ~(layer0_outputs[5686]);
    assign outputs[6826] = layer0_outputs[3480];
    assign outputs[6827] = ~((layer0_outputs[9375]) ^ (layer0_outputs[2518]));
    assign outputs[6828] = (layer0_outputs[461]) ^ (layer0_outputs[5676]);
    assign outputs[6829] = ~((layer0_outputs[7980]) ^ (layer0_outputs[3325]));
    assign outputs[6830] = (layer0_outputs[32]) ^ (layer0_outputs[2457]);
    assign outputs[6831] = layer0_outputs[9675];
    assign outputs[6832] = ~(layer0_outputs[5509]);
    assign outputs[6833] = layer0_outputs[9815];
    assign outputs[6834] = ~(layer0_outputs[6795]);
    assign outputs[6835] = ~(layer0_outputs[8329]);
    assign outputs[6836] = ~((layer0_outputs[489]) ^ (layer0_outputs[6947]));
    assign outputs[6837] = (layer0_outputs[9135]) & ~(layer0_outputs[1016]);
    assign outputs[6838] = ~((layer0_outputs[1725]) | (layer0_outputs[2516]));
    assign outputs[6839] = ~(layer0_outputs[8991]);
    assign outputs[6840] = ~((layer0_outputs[4936]) ^ (layer0_outputs[4039]));
    assign outputs[6841] = (layer0_outputs[7887]) & ~(layer0_outputs[6565]);
    assign outputs[6842] = ~((layer0_outputs[9991]) & (layer0_outputs[9914]));
    assign outputs[6843] = ~(layer0_outputs[1652]);
    assign outputs[6844] = ~(layer0_outputs[7854]) | (layer0_outputs[2343]);
    assign outputs[6845] = ~((layer0_outputs[8472]) ^ (layer0_outputs[7336]));
    assign outputs[6846] = ~((layer0_outputs[8375]) ^ (layer0_outputs[4990]));
    assign outputs[6847] = layer0_outputs[7446];
    assign outputs[6848] = (layer0_outputs[2279]) & ~(layer0_outputs[347]);
    assign outputs[6849] = layer0_outputs[3986];
    assign outputs[6850] = (layer0_outputs[8253]) | (layer0_outputs[6593]);
    assign outputs[6851] = ~(layer0_outputs[9269]);
    assign outputs[6852] = layer0_outputs[4470];
    assign outputs[6853] = (layer0_outputs[943]) ^ (layer0_outputs[2284]);
    assign outputs[6854] = (layer0_outputs[6507]) ^ (layer0_outputs[9350]);
    assign outputs[6855] = ~(layer0_outputs[2205]);
    assign outputs[6856] = ~((layer0_outputs[4536]) | (layer0_outputs[305]));
    assign outputs[6857] = ~(layer0_outputs[9800]);
    assign outputs[6858] = layer0_outputs[2697];
    assign outputs[6859] = layer0_outputs[8219];
    assign outputs[6860] = (layer0_outputs[9253]) & (layer0_outputs[5528]);
    assign outputs[6861] = layer0_outputs[5279];
    assign outputs[6862] = layer0_outputs[9932];
    assign outputs[6863] = ~(layer0_outputs[489]) | (layer0_outputs[4606]);
    assign outputs[6864] = (layer0_outputs[5867]) & ~(layer0_outputs[6568]);
    assign outputs[6865] = ~(layer0_outputs[9140]);
    assign outputs[6866] = (layer0_outputs[9869]) & (layer0_outputs[2782]);
    assign outputs[6867] = layer0_outputs[2996];
    assign outputs[6868] = layer0_outputs[2295];
    assign outputs[6869] = layer0_outputs[5186];
    assign outputs[6870] = layer0_outputs[10180];
    assign outputs[6871] = layer0_outputs[1024];
    assign outputs[6872] = ~(layer0_outputs[7828]);
    assign outputs[6873] = layer0_outputs[6168];
    assign outputs[6874] = layer0_outputs[3521];
    assign outputs[6875] = ~(layer0_outputs[2853]);
    assign outputs[6876] = layer0_outputs[2586];
    assign outputs[6877] = (layer0_outputs[6384]) & ~(layer0_outputs[4218]);
    assign outputs[6878] = layer0_outputs[7776];
    assign outputs[6879] = (layer0_outputs[1518]) & ~(layer0_outputs[3191]);
    assign outputs[6880] = layer0_outputs[363];
    assign outputs[6881] = ~(layer0_outputs[3049]);
    assign outputs[6882] = layer0_outputs[2462];
    assign outputs[6883] = ~(layer0_outputs[6471]);
    assign outputs[6884] = ~(layer0_outputs[712]);
    assign outputs[6885] = layer0_outputs[3972];
    assign outputs[6886] = layer0_outputs[10018];
    assign outputs[6887] = (layer0_outputs[6334]) & (layer0_outputs[4441]);
    assign outputs[6888] = layer0_outputs[5924];
    assign outputs[6889] = (layer0_outputs[995]) ^ (layer0_outputs[8736]);
    assign outputs[6890] = layer0_outputs[5694];
    assign outputs[6891] = (layer0_outputs[2695]) & ~(layer0_outputs[7223]);
    assign outputs[6892] = layer0_outputs[9758];
    assign outputs[6893] = ~((layer0_outputs[1995]) & (layer0_outputs[2836]));
    assign outputs[6894] = ~(layer0_outputs[9784]);
    assign outputs[6895] = (layer0_outputs[1825]) & ~(layer0_outputs[3342]);
    assign outputs[6896] = ~((layer0_outputs[7399]) ^ (layer0_outputs[2834]));
    assign outputs[6897] = ~(layer0_outputs[1974]);
    assign outputs[6898] = layer0_outputs[9588];
    assign outputs[6899] = ~(layer0_outputs[4803]);
    assign outputs[6900] = ~(layer0_outputs[1675]);
    assign outputs[6901] = (layer0_outputs[8680]) & ~(layer0_outputs[6849]);
    assign outputs[6902] = ~(layer0_outputs[5188]);
    assign outputs[6903] = ~((layer0_outputs[5347]) | (layer0_outputs[8652]));
    assign outputs[6904] = ~(layer0_outputs[6714]);
    assign outputs[6905] = layer0_outputs[2934];
    assign outputs[6906] = (layer0_outputs[8363]) ^ (layer0_outputs[802]);
    assign outputs[6907] = layer0_outputs[8273];
    assign outputs[6908] = ~((layer0_outputs[9615]) | (layer0_outputs[4269]));
    assign outputs[6909] = layer0_outputs[8076];
    assign outputs[6910] = (layer0_outputs[8855]) & (layer0_outputs[35]);
    assign outputs[6911] = ~(layer0_outputs[1689]);
    assign outputs[6912] = (layer0_outputs[6256]) & ~(layer0_outputs[787]);
    assign outputs[6913] = ~(layer0_outputs[3962]);
    assign outputs[6914] = layer0_outputs[9088];
    assign outputs[6915] = ~((layer0_outputs[3190]) | (layer0_outputs[1469]));
    assign outputs[6916] = layer0_outputs[3529];
    assign outputs[6917] = ~(layer0_outputs[5978]);
    assign outputs[6918] = ~(layer0_outputs[8572]);
    assign outputs[6919] = ~((layer0_outputs[9522]) | (layer0_outputs[4457]));
    assign outputs[6920] = ~(layer0_outputs[8722]);
    assign outputs[6921] = ~(layer0_outputs[5393]);
    assign outputs[6922] = layer0_outputs[601];
    assign outputs[6923] = ~(layer0_outputs[2804]);
    assign outputs[6924] = (layer0_outputs[5127]) ^ (layer0_outputs[6051]);
    assign outputs[6925] = (layer0_outputs[2340]) & ~(layer0_outputs[6694]);
    assign outputs[6926] = ~(layer0_outputs[9819]);
    assign outputs[6927] = ~(layer0_outputs[7914]) | (layer0_outputs[7697]);
    assign outputs[6928] = layer0_outputs[10061];
    assign outputs[6929] = layer0_outputs[8515];
    assign outputs[6930] = (layer0_outputs[500]) & ~(layer0_outputs[7276]);
    assign outputs[6931] = ~((layer0_outputs[1042]) | (layer0_outputs[6994]));
    assign outputs[6932] = (layer0_outputs[3557]) & ~(layer0_outputs[10203]);
    assign outputs[6933] = (layer0_outputs[3734]) & ~(layer0_outputs[10168]);
    assign outputs[6934] = ~((layer0_outputs[4514]) ^ (layer0_outputs[753]));
    assign outputs[6935] = ~(layer0_outputs[8130]) | (layer0_outputs[1918]);
    assign outputs[6936] = layer0_outputs[891];
    assign outputs[6937] = layer0_outputs[5844];
    assign outputs[6938] = layer0_outputs[8199];
    assign outputs[6939] = layer0_outputs[8360];
    assign outputs[6940] = layer0_outputs[9921];
    assign outputs[6941] = ~((layer0_outputs[7586]) | (layer0_outputs[3258]));
    assign outputs[6942] = ~((layer0_outputs[6444]) & (layer0_outputs[7362]));
    assign outputs[6943] = layer0_outputs[7091];
    assign outputs[6944] = ~(layer0_outputs[593]);
    assign outputs[6945] = layer0_outputs[9532];
    assign outputs[6946] = (layer0_outputs[1735]) & ~(layer0_outputs[4778]);
    assign outputs[6947] = ~(layer0_outputs[8842]);
    assign outputs[6948] = ~(layer0_outputs[1893]);
    assign outputs[6949] = (layer0_outputs[2542]) & (layer0_outputs[3727]);
    assign outputs[6950] = layer0_outputs[6728];
    assign outputs[6951] = (layer0_outputs[9964]) & ~(layer0_outputs[2707]);
    assign outputs[6952] = layer0_outputs[5738];
    assign outputs[6953] = ~(layer0_outputs[2350]);
    assign outputs[6954] = layer0_outputs[4112];
    assign outputs[6955] = ~(layer0_outputs[4224]);
    assign outputs[6956] = ~(layer0_outputs[1377]);
    assign outputs[6957] = layer0_outputs[10129];
    assign outputs[6958] = ~(layer0_outputs[564]);
    assign outputs[6959] = layer0_outputs[3380];
    assign outputs[6960] = ~(layer0_outputs[9460]);
    assign outputs[6961] = (layer0_outputs[4575]) & ~(layer0_outputs[7845]);
    assign outputs[6962] = ~(layer0_outputs[1491]);
    assign outputs[6963] = layer0_outputs[5764];
    assign outputs[6964] = (layer0_outputs[5693]) & (layer0_outputs[360]);
    assign outputs[6965] = ~((layer0_outputs[6772]) ^ (layer0_outputs[5191]));
    assign outputs[6966] = ~((layer0_outputs[3390]) | (layer0_outputs[238]));
    assign outputs[6967] = layer0_outputs[4717];
    assign outputs[6968] = ~((layer0_outputs[878]) | (layer0_outputs[1715]));
    assign outputs[6969] = (layer0_outputs[6232]) ^ (layer0_outputs[3960]);
    assign outputs[6970] = (layer0_outputs[3177]) & (layer0_outputs[9869]);
    assign outputs[6971] = layer0_outputs[6792];
    assign outputs[6972] = ~((layer0_outputs[4808]) ^ (layer0_outputs[1254]));
    assign outputs[6973] = layer0_outputs[6746];
    assign outputs[6974] = ~(layer0_outputs[9670]);
    assign outputs[6975] = ~(layer0_outputs[2622]);
    assign outputs[6976] = ~(layer0_outputs[7355]);
    assign outputs[6977] = layer0_outputs[3140];
    assign outputs[6978] = layer0_outputs[7709];
    assign outputs[6979] = (layer0_outputs[9357]) & (layer0_outputs[5397]);
    assign outputs[6980] = (layer0_outputs[2944]) & (layer0_outputs[7878]);
    assign outputs[6981] = ~(layer0_outputs[5534]);
    assign outputs[6982] = ~(layer0_outputs[8353]);
    assign outputs[6983] = layer0_outputs[7034];
    assign outputs[6984] = ~(layer0_outputs[2701]);
    assign outputs[6985] = layer0_outputs[3379];
    assign outputs[6986] = ~(layer0_outputs[833]);
    assign outputs[6987] = ~(layer0_outputs[1066]);
    assign outputs[6988] = (layer0_outputs[2588]) ^ (layer0_outputs[2098]);
    assign outputs[6989] = ~((layer0_outputs[1879]) | (layer0_outputs[2477]));
    assign outputs[6990] = layer0_outputs[6646];
    assign outputs[6991] = (layer0_outputs[2881]) & ~(layer0_outputs[5724]);
    assign outputs[6992] = ~(layer0_outputs[5345]);
    assign outputs[6993] = layer0_outputs[9098];
    assign outputs[6994] = (layer0_outputs[7307]) & ~(layer0_outputs[9660]);
    assign outputs[6995] = ~(layer0_outputs[9547]);
    assign outputs[6996] = layer0_outputs[1807];
    assign outputs[6997] = ~(layer0_outputs[3544]);
    assign outputs[6998] = layer0_outputs[6012];
    assign outputs[6999] = ~((layer0_outputs[6770]) & (layer0_outputs[3156]));
    assign outputs[7000] = layer0_outputs[13];
    assign outputs[7001] = ~(layer0_outputs[3843]);
    assign outputs[7002] = layer0_outputs[10081];
    assign outputs[7003] = ~(layer0_outputs[2254]);
    assign outputs[7004] = (layer0_outputs[6962]) & ~(layer0_outputs[447]);
    assign outputs[7005] = ~(layer0_outputs[4877]);
    assign outputs[7006] = ~((layer0_outputs[5394]) ^ (layer0_outputs[432]));
    assign outputs[7007] = layer0_outputs[7524];
    assign outputs[7008] = ~(layer0_outputs[2921]);
    assign outputs[7009] = layer0_outputs[7027];
    assign outputs[7010] = ~(layer0_outputs[1476]) | (layer0_outputs[3798]);
    assign outputs[7011] = ~(layer0_outputs[7154]);
    assign outputs[7012] = ~(layer0_outputs[1709]);
    assign outputs[7013] = layer0_outputs[9875];
    assign outputs[7014] = layer0_outputs[4075];
    assign outputs[7015] = (layer0_outputs[3149]) & ~(layer0_outputs[9587]);
    assign outputs[7016] = ~((layer0_outputs[9968]) | (layer0_outputs[3249]));
    assign outputs[7017] = ~(layer0_outputs[10172]);
    assign outputs[7018] = ~(layer0_outputs[7904]);
    assign outputs[7019] = layer0_outputs[2573];
    assign outputs[7020] = ~(layer0_outputs[3536]);
    assign outputs[7021] = ~((layer0_outputs[6048]) ^ (layer0_outputs[9093]));
    assign outputs[7022] = ~(layer0_outputs[10179]);
    assign outputs[7023] = ~(layer0_outputs[1727]);
    assign outputs[7024] = ~(layer0_outputs[809]);
    assign outputs[7025] = ~(layer0_outputs[5246]);
    assign outputs[7026] = ~(layer0_outputs[498]) | (layer0_outputs[9038]);
    assign outputs[7027] = ~((layer0_outputs[2012]) ^ (layer0_outputs[538]));
    assign outputs[7028] = layer0_outputs[234];
    assign outputs[7029] = ~(layer0_outputs[3227]);
    assign outputs[7030] = ~(layer0_outputs[9315]);
    assign outputs[7031] = ~((layer0_outputs[4613]) | (layer0_outputs[6657]));
    assign outputs[7032] = ~(layer0_outputs[5245]);
    assign outputs[7033] = (layer0_outputs[5755]) ^ (layer0_outputs[4478]);
    assign outputs[7034] = (layer0_outputs[9459]) & ~(layer0_outputs[8577]);
    assign outputs[7035] = (layer0_outputs[4562]) & (layer0_outputs[970]);
    assign outputs[7036] = ~(layer0_outputs[4926]);
    assign outputs[7037] = ~(layer0_outputs[3886]);
    assign outputs[7038] = ~(layer0_outputs[4857]);
    assign outputs[7039] = ~(layer0_outputs[6804]);
    assign outputs[7040] = layer0_outputs[7780];
    assign outputs[7041] = ~(layer0_outputs[9107]);
    assign outputs[7042] = (layer0_outputs[7501]) & ~(layer0_outputs[7526]);
    assign outputs[7043] = layer0_outputs[7570];
    assign outputs[7044] = (layer0_outputs[1778]) & ~(layer0_outputs[5697]);
    assign outputs[7045] = (layer0_outputs[6933]) ^ (layer0_outputs[10198]);
    assign outputs[7046] = layer0_outputs[1648];
    assign outputs[7047] = ~(layer0_outputs[8975]);
    assign outputs[7048] = ~(layer0_outputs[9578]);
    assign outputs[7049] = ~((layer0_outputs[9384]) | (layer0_outputs[1263]));
    assign outputs[7050] = ~(layer0_outputs[6628]);
    assign outputs[7051] = ~(layer0_outputs[2438]);
    assign outputs[7052] = layer0_outputs[2132];
    assign outputs[7053] = ~(layer0_outputs[5330]);
    assign outputs[7054] = layer0_outputs[2037];
    assign outputs[7055] = ~(layer0_outputs[5493]);
    assign outputs[7056] = layer0_outputs[4970];
    assign outputs[7057] = layer0_outputs[5725];
    assign outputs[7058] = ~(layer0_outputs[3856]);
    assign outputs[7059] = (layer0_outputs[4530]) & ~(layer0_outputs[3403]);
    assign outputs[7060] = layer0_outputs[3144];
    assign outputs[7061] = ~(layer0_outputs[2933]);
    assign outputs[7062] = ~(layer0_outputs[3198]) | (layer0_outputs[5741]);
    assign outputs[7063] = (layer0_outputs[654]) & (layer0_outputs[8283]);
    assign outputs[7064] = ~(layer0_outputs[7935]);
    assign outputs[7065] = layer0_outputs[3840];
    assign outputs[7066] = layer0_outputs[3485];
    assign outputs[7067] = layer0_outputs[7584];
    assign outputs[7068] = layer0_outputs[5040];
    assign outputs[7069] = layer0_outputs[3163];
    assign outputs[7070] = ~((layer0_outputs[5478]) | (layer0_outputs[1608]));
    assign outputs[7071] = ~(layer0_outputs[1826]);
    assign outputs[7072] = layer0_outputs[1259];
    assign outputs[7073] = layer0_outputs[5927];
    assign outputs[7074] = layer0_outputs[3687];
    assign outputs[7075] = layer0_outputs[1480];
    assign outputs[7076] = ~(layer0_outputs[4195]);
    assign outputs[7077] = layer0_outputs[6654];
    assign outputs[7078] = ~((layer0_outputs[6076]) ^ (layer0_outputs[6748]));
    assign outputs[7079] = ~(layer0_outputs[9127]);
    assign outputs[7080] = (layer0_outputs[10162]) ^ (layer0_outputs[769]);
    assign outputs[7081] = ~(layer0_outputs[7266]);
    assign outputs[7082] = (layer0_outputs[5263]) & ~(layer0_outputs[9229]);
    assign outputs[7083] = ~(layer0_outputs[6658]);
    assign outputs[7084] = ~(layer0_outputs[9865]);
    assign outputs[7085] = ~((layer0_outputs[3387]) ^ (layer0_outputs[5702]));
    assign outputs[7086] = layer0_outputs[6250];
    assign outputs[7087] = ~(layer0_outputs[455]) | (layer0_outputs[1474]);
    assign outputs[7088] = (layer0_outputs[8712]) & ~(layer0_outputs[8688]);
    assign outputs[7089] = ~(layer0_outputs[190]);
    assign outputs[7090] = layer0_outputs[7282];
    assign outputs[7091] = (layer0_outputs[7172]) & ~(layer0_outputs[3774]);
    assign outputs[7092] = ~(layer0_outputs[1687]);
    assign outputs[7093] = layer0_outputs[5747];
    assign outputs[7094] = layer0_outputs[428];
    assign outputs[7095] = ~((layer0_outputs[3671]) ^ (layer0_outputs[1720]));
    assign outputs[7096] = ~(layer0_outputs[5572]);
    assign outputs[7097] = ~((layer0_outputs[1064]) | (layer0_outputs[3377]));
    assign outputs[7098] = ~(layer0_outputs[9774]);
    assign outputs[7099] = layer0_outputs[4764];
    assign outputs[7100] = layer0_outputs[8279];
    assign outputs[7101] = layer0_outputs[1162];
    assign outputs[7102] = layer0_outputs[689];
    assign outputs[7103] = ~(layer0_outputs[10006]);
    assign outputs[7104] = ~(layer0_outputs[9924]);
    assign outputs[7105] = ~((layer0_outputs[287]) ^ (layer0_outputs[3064]));
    assign outputs[7106] = layer0_outputs[141];
    assign outputs[7107] = layer0_outputs[5830];
    assign outputs[7108] = ~(layer0_outputs[10051]);
    assign outputs[7109] = (layer0_outputs[10119]) ^ (layer0_outputs[3478]);
    assign outputs[7110] = (layer0_outputs[450]) & ~(layer0_outputs[7238]);
    assign outputs[7111] = (layer0_outputs[9518]) & ~(layer0_outputs[9386]);
    assign outputs[7112] = layer0_outputs[9251];
    assign outputs[7113] = (layer0_outputs[4756]) & ~(layer0_outputs[717]);
    assign outputs[7114] = layer0_outputs[1980];
    assign outputs[7115] = layer0_outputs[1952];
    assign outputs[7116] = (layer0_outputs[3409]) & (layer0_outputs[5254]);
    assign outputs[7117] = ~(layer0_outputs[7376]);
    assign outputs[7118] = ~((layer0_outputs[9316]) & (layer0_outputs[6485]));
    assign outputs[7119] = (layer0_outputs[6890]) & (layer0_outputs[3681]);
    assign outputs[7120] = ~(layer0_outputs[6602]) | (layer0_outputs[2488]);
    assign outputs[7121] = layer0_outputs[3130];
    assign outputs[7122] = ~(layer0_outputs[5302]) | (layer0_outputs[5213]);
    assign outputs[7123] = ~(layer0_outputs[4490]);
    assign outputs[7124] = ~(layer0_outputs[997]);
    assign outputs[7125] = ~(layer0_outputs[2806]) | (layer0_outputs[7666]);
    assign outputs[7126] = ~(layer0_outputs[5081]);
    assign outputs[7127] = ~(layer0_outputs[1326]) | (layer0_outputs[1140]);
    assign outputs[7128] = layer0_outputs[4437];
    assign outputs[7129] = layer0_outputs[8694];
    assign outputs[7130] = ~(layer0_outputs[7313]);
    assign outputs[7131] = layer0_outputs[8173];
    assign outputs[7132] = (layer0_outputs[361]) ^ (layer0_outputs[7482]);
    assign outputs[7133] = (layer0_outputs[5148]) | (layer0_outputs[6807]);
    assign outputs[7134] = (layer0_outputs[8065]) & (layer0_outputs[8]);
    assign outputs[7135] = layer0_outputs[3754];
    assign outputs[7136] = ~((layer0_outputs[825]) | (layer0_outputs[1971]));
    assign outputs[7137] = layer0_outputs[2816];
    assign outputs[7138] = ~((layer0_outputs[6459]) | (layer0_outputs[981]));
    assign outputs[7139] = (layer0_outputs[7553]) | (layer0_outputs[9585]);
    assign outputs[7140] = (layer0_outputs[1210]) & ~(layer0_outputs[1587]);
    assign outputs[7141] = (layer0_outputs[9707]) & ~(layer0_outputs[946]);
    assign outputs[7142] = ~(layer0_outputs[4085]);
    assign outputs[7143] = ~((layer0_outputs[5970]) ^ (layer0_outputs[1617]));
    assign outputs[7144] = layer0_outputs[3983];
    assign outputs[7145] = (layer0_outputs[1966]) & ~(layer0_outputs[2790]);
    assign outputs[7146] = layer0_outputs[6010];
    assign outputs[7147] = (layer0_outputs[852]) & (layer0_outputs[8844]);
    assign outputs[7148] = ~(layer0_outputs[1387]);
    assign outputs[7149] = ~(layer0_outputs[708]);
    assign outputs[7150] = ~(layer0_outputs[2459]);
    assign outputs[7151] = ~((layer0_outputs[3984]) & (layer0_outputs[2437]));
    assign outputs[7152] = (layer0_outputs[1330]) & (layer0_outputs[8886]);
    assign outputs[7153] = layer0_outputs[9310];
    assign outputs[7154] = layer0_outputs[9679];
    assign outputs[7155] = layer0_outputs[8773];
    assign outputs[7156] = ~(layer0_outputs[5961]);
    assign outputs[7157] = layer0_outputs[4590];
    assign outputs[7158] = (layer0_outputs[1925]) ^ (layer0_outputs[2489]);
    assign outputs[7159] = layer0_outputs[3986];
    assign outputs[7160] = layer0_outputs[1332];
    assign outputs[7161] = (layer0_outputs[6728]) ^ (layer0_outputs[2846]);
    assign outputs[7162] = ~(layer0_outputs[7041]);
    assign outputs[7163] = (layer0_outputs[3693]) ^ (layer0_outputs[9957]);
    assign outputs[7164] = ~((layer0_outputs[3275]) ^ (layer0_outputs[9861]));
    assign outputs[7165] = ~((layer0_outputs[2408]) & (layer0_outputs[4906]));
    assign outputs[7166] = (layer0_outputs[3574]) ^ (layer0_outputs[1843]);
    assign outputs[7167] = (layer0_outputs[3280]) & ~(layer0_outputs[6150]);
    assign outputs[7168] = ~(layer0_outputs[3034]);
    assign outputs[7169] = layer0_outputs[666];
    assign outputs[7170] = layer0_outputs[7574];
    assign outputs[7171] = ~(layer0_outputs[2590]) | (layer0_outputs[303]);
    assign outputs[7172] = ~(layer0_outputs[8204]);
    assign outputs[7173] = layer0_outputs[7763];
    assign outputs[7174] = ~(layer0_outputs[2372]);
    assign outputs[7175] = (layer0_outputs[2383]) & ~(layer0_outputs[7286]);
    assign outputs[7176] = layer0_outputs[1602];
    assign outputs[7177] = ~(layer0_outputs[9977]);
    assign outputs[7178] = ~((layer0_outputs[9720]) ^ (layer0_outputs[8358]));
    assign outputs[7179] = (layer0_outputs[9506]) & ~(layer0_outputs[9754]);
    assign outputs[7180] = ~(layer0_outputs[7523]);
    assign outputs[7181] = layer0_outputs[10133];
    assign outputs[7182] = (layer0_outputs[2337]) & (layer0_outputs[477]);
    assign outputs[7183] = layer0_outputs[4103];
    assign outputs[7184] = layer0_outputs[4443];
    assign outputs[7185] = layer0_outputs[3537];
    assign outputs[7186] = ~((layer0_outputs[9014]) | (layer0_outputs[6957]));
    assign outputs[7187] = ~((layer0_outputs[7299]) ^ (layer0_outputs[856]));
    assign outputs[7188] = ~(layer0_outputs[3732]);
    assign outputs[7189] = ~(layer0_outputs[4187]);
    assign outputs[7190] = (layer0_outputs[3556]) & ~(layer0_outputs[2447]);
    assign outputs[7191] = ~(layer0_outputs[8873]);
    assign outputs[7192] = (layer0_outputs[9362]) & ~(layer0_outputs[2540]);
    assign outputs[7193] = (layer0_outputs[5630]) & ~(layer0_outputs[5573]);
    assign outputs[7194] = (layer0_outputs[3216]) & ~(layer0_outputs[6519]);
    assign outputs[7195] = layer0_outputs[4541];
    assign outputs[7196] = layer0_outputs[3883];
    assign outputs[7197] = (layer0_outputs[6789]) & ~(layer0_outputs[6676]);
    assign outputs[7198] = layer0_outputs[7601];
    assign outputs[7199] = layer0_outputs[9212];
    assign outputs[7200] = ~((layer0_outputs[2391]) ^ (layer0_outputs[4106]));
    assign outputs[7201] = layer0_outputs[5171];
    assign outputs[7202] = ~(layer0_outputs[1874]);
    assign outputs[7203] = layer0_outputs[462];
    assign outputs[7204] = layer0_outputs[244];
    assign outputs[7205] = (layer0_outputs[5073]) | (layer0_outputs[8583]);
    assign outputs[7206] = (layer0_outputs[8213]) ^ (layer0_outputs[4754]);
    assign outputs[7207] = ~((layer0_outputs[3598]) ^ (layer0_outputs[382]));
    assign outputs[7208] = (layer0_outputs[9688]) ^ (layer0_outputs[2743]);
    assign outputs[7209] = ~((layer0_outputs[2160]) ^ (layer0_outputs[7497]));
    assign outputs[7210] = ~(layer0_outputs[3681]);
    assign outputs[7211] = layer0_outputs[6797];
    assign outputs[7212] = ~(layer0_outputs[10115]);
    assign outputs[7213] = layer0_outputs[6034];
    assign outputs[7214] = layer0_outputs[4723];
    assign outputs[7215] = ~(layer0_outputs[9621]) | (layer0_outputs[1701]);
    assign outputs[7216] = (layer0_outputs[651]) ^ (layer0_outputs[5076]);
    assign outputs[7217] = ~(layer0_outputs[6249]) | (layer0_outputs[975]);
    assign outputs[7218] = layer0_outputs[1147];
    assign outputs[7219] = (layer0_outputs[7851]) | (layer0_outputs[2497]);
    assign outputs[7220] = ~((layer0_outputs[7866]) ^ (layer0_outputs[4159]));
    assign outputs[7221] = layer0_outputs[9427];
    assign outputs[7222] = (layer0_outputs[4385]) ^ (layer0_outputs[3703]);
    assign outputs[7223] = layer0_outputs[4947];
    assign outputs[7224] = (layer0_outputs[6990]) & ~(layer0_outputs[1345]);
    assign outputs[7225] = (layer0_outputs[6663]) ^ (layer0_outputs[4792]);
    assign outputs[7226] = (layer0_outputs[4335]) & ~(layer0_outputs[9490]);
    assign outputs[7227] = ~(layer0_outputs[3654]);
    assign outputs[7228] = (layer0_outputs[1575]) & ~(layer0_outputs[1408]);
    assign outputs[7229] = ~(layer0_outputs[9762]);
    assign outputs[7230] = (layer0_outputs[6333]) | (layer0_outputs[6515]);
    assign outputs[7231] = (layer0_outputs[4912]) ^ (layer0_outputs[3878]);
    assign outputs[7232] = ~(layer0_outputs[7196]) | (layer0_outputs[6201]);
    assign outputs[7233] = ~(layer0_outputs[9341]);
    assign outputs[7234] = ~((layer0_outputs[885]) ^ (layer0_outputs[3846]));
    assign outputs[7235] = (layer0_outputs[7025]) | (layer0_outputs[4905]);
    assign outputs[7236] = ~((layer0_outputs[3859]) | (layer0_outputs[5371]));
    assign outputs[7237] = (layer0_outputs[4419]) & (layer0_outputs[637]);
    assign outputs[7238] = layer0_outputs[5783];
    assign outputs[7239] = layer0_outputs[9928];
    assign outputs[7240] = ~(layer0_outputs[1239]);
    assign outputs[7241] = (layer0_outputs[6002]) & ~(layer0_outputs[3219]);
    assign outputs[7242] = (layer0_outputs[1309]) & (layer0_outputs[10074]);
    assign outputs[7243] = (layer0_outputs[6542]) ^ (layer0_outputs[3098]);
    assign outputs[7244] = ~((layer0_outputs[2633]) | (layer0_outputs[1211]));
    assign outputs[7245] = (layer0_outputs[8996]) & ~(layer0_outputs[7151]);
    assign outputs[7246] = ~((layer0_outputs[3907]) | (layer0_outputs[4768]));
    assign outputs[7247] = ~(layer0_outputs[10190]) | (layer0_outputs[6802]);
    assign outputs[7248] = (layer0_outputs[4399]) | (layer0_outputs[4609]);
    assign outputs[7249] = ~((layer0_outputs[9142]) ^ (layer0_outputs[2889]));
    assign outputs[7250] = layer0_outputs[8004];
    assign outputs[7251] = ~((layer0_outputs[9685]) ^ (layer0_outputs[5084]));
    assign outputs[7252] = ~(layer0_outputs[6852]);
    assign outputs[7253] = ~(layer0_outputs[4010]) | (layer0_outputs[9087]);
    assign outputs[7254] = ~(layer0_outputs[8531]) | (layer0_outputs[5804]);
    assign outputs[7255] = ~(layer0_outputs[2362]);
    assign outputs[7256] = ~(layer0_outputs[8402]);
    assign outputs[7257] = ~(layer0_outputs[6793]);
    assign outputs[7258] = ~(layer0_outputs[6263]);
    assign outputs[7259] = (layer0_outputs[4162]) & (layer0_outputs[1091]);
    assign outputs[7260] = (layer0_outputs[2375]) & (layer0_outputs[3853]);
    assign outputs[7261] = (layer0_outputs[1568]) & ~(layer0_outputs[2500]);
    assign outputs[7262] = (layer0_outputs[4264]) ^ (layer0_outputs[456]);
    assign outputs[7263] = (layer0_outputs[8363]) & ~(layer0_outputs[6418]);
    assign outputs[7264] = (layer0_outputs[4222]) ^ (layer0_outputs[6961]);
    assign outputs[7265] = (layer0_outputs[3829]) & ~(layer0_outputs[9154]);
    assign outputs[7266] = layer0_outputs[5869];
    assign outputs[7267] = (layer0_outputs[1237]) & ~(layer0_outputs[4967]);
    assign outputs[7268] = layer0_outputs[7715];
    assign outputs[7269] = (layer0_outputs[1860]) & (layer0_outputs[5745]);
    assign outputs[7270] = ~((layer0_outputs[1023]) ^ (layer0_outputs[27]));
    assign outputs[7271] = layer0_outputs[7101];
    assign outputs[7272] = (layer0_outputs[7520]) ^ (layer0_outputs[10125]);
    assign outputs[7273] = layer0_outputs[5111];
    assign outputs[7274] = ~(layer0_outputs[4488]);
    assign outputs[7275] = (layer0_outputs[5821]) ^ (layer0_outputs[8827]);
    assign outputs[7276] = layer0_outputs[254];
    assign outputs[7277] = layer0_outputs[571];
    assign outputs[7278] = ~((layer0_outputs[8413]) & (layer0_outputs[8280]));
    assign outputs[7279] = ~((layer0_outputs[6308]) ^ (layer0_outputs[9224]));
    assign outputs[7280] = (layer0_outputs[1189]) | (layer0_outputs[5465]);
    assign outputs[7281] = (layer0_outputs[8738]) & (layer0_outputs[3898]);
    assign outputs[7282] = (layer0_outputs[2383]) & ~(layer0_outputs[4470]);
    assign outputs[7283] = (layer0_outputs[7226]) & ~(layer0_outputs[9596]);
    assign outputs[7284] = (layer0_outputs[3403]) & ~(layer0_outputs[8913]);
    assign outputs[7285] = ~((layer0_outputs[5028]) & (layer0_outputs[7006]));
    assign outputs[7286] = layer0_outputs[6341];
    assign outputs[7287] = ~((layer0_outputs[4071]) ^ (layer0_outputs[8439]));
    assign outputs[7288] = ~(layer0_outputs[4163]);
    assign outputs[7289] = layer0_outputs[9306];
    assign outputs[7290] = ~(layer0_outputs[5916]);
    assign outputs[7291] = ~(layer0_outputs[4682]);
    assign outputs[7292] = ~(layer0_outputs[6255]);
    assign outputs[7293] = ~(layer0_outputs[9882]);
    assign outputs[7294] = ~((layer0_outputs[8123]) & (layer0_outputs[9513]));
    assign outputs[7295] = layer0_outputs[7320];
    assign outputs[7296] = (layer0_outputs[5905]) ^ (layer0_outputs[3751]);
    assign outputs[7297] = ~(layer0_outputs[6396]);
    assign outputs[7298] = (layer0_outputs[936]) & ~(layer0_outputs[9243]);
    assign outputs[7299] = layer0_outputs[9925];
    assign outputs[7300] = ~((layer0_outputs[10024]) & (layer0_outputs[2544]));
    assign outputs[7301] = ~(layer0_outputs[978]);
    assign outputs[7302] = ~((layer0_outputs[2508]) | (layer0_outputs[3649]));
    assign outputs[7303] = (layer0_outputs[5645]) ^ (layer0_outputs[5333]);
    assign outputs[7304] = ~(layer0_outputs[1437]);
    assign outputs[7305] = layer0_outputs[3245];
    assign outputs[7306] = (layer0_outputs[9386]) | (layer0_outputs[4566]);
    assign outputs[7307] = layer0_outputs[6513];
    assign outputs[7308] = ~((layer0_outputs[5075]) | (layer0_outputs[583]));
    assign outputs[7309] = ~(layer0_outputs[5057]) | (layer0_outputs[1274]);
    assign outputs[7310] = (layer0_outputs[4638]) & ~(layer0_outputs[3491]);
    assign outputs[7311] = ~((layer0_outputs[1504]) | (layer0_outputs[9875]));
    assign outputs[7312] = ~(layer0_outputs[1786]);
    assign outputs[7313] = ~(layer0_outputs[8788]);
    assign outputs[7314] = ~(layer0_outputs[5779]);
    assign outputs[7315] = layer0_outputs[5449];
    assign outputs[7316] = (layer0_outputs[3783]) & ~(layer0_outputs[5203]);
    assign outputs[7317] = ~(layer0_outputs[401]);
    assign outputs[7318] = (layer0_outputs[6065]) ^ (layer0_outputs[1144]);
    assign outputs[7319] = ~(layer0_outputs[3657]);
    assign outputs[7320] = layer0_outputs[9894];
    assign outputs[7321] = ~(layer0_outputs[2712]);
    assign outputs[7322] = ~(layer0_outputs[2916]);
    assign outputs[7323] = layer0_outputs[6466];
    assign outputs[7324] = (layer0_outputs[4762]) & ~(layer0_outputs[4922]);
    assign outputs[7325] = layer0_outputs[3119];
    assign outputs[7326] = ~(layer0_outputs[6339]);
    assign outputs[7327] = ~(layer0_outputs[7782]);
    assign outputs[7328] = layer0_outputs[6092];
    assign outputs[7329] = layer0_outputs[3642];
    assign outputs[7330] = (layer0_outputs[7405]) & ~(layer0_outputs[5649]);
    assign outputs[7331] = ~(layer0_outputs[1631]);
    assign outputs[7332] = layer0_outputs[10012];
    assign outputs[7333] = layer0_outputs[8850];
    assign outputs[7334] = (layer0_outputs[1965]) | (layer0_outputs[8740]);
    assign outputs[7335] = ~(layer0_outputs[6058]);
    assign outputs[7336] = layer0_outputs[1125];
    assign outputs[7337] = (layer0_outputs[6387]) ^ (layer0_outputs[3858]);
    assign outputs[7338] = ~(layer0_outputs[5666]);
    assign outputs[7339] = layer0_outputs[1741];
    assign outputs[7340] = layer0_outputs[6817];
    assign outputs[7341] = ~((layer0_outputs[2178]) | (layer0_outputs[1477]));
    assign outputs[7342] = (layer0_outputs[7321]) & ~(layer0_outputs[5488]);
    assign outputs[7343] = ~((layer0_outputs[449]) ^ (layer0_outputs[5960]));
    assign outputs[7344] = ~((layer0_outputs[6742]) | (layer0_outputs[9534]));
    assign outputs[7345] = layer0_outputs[3780];
    assign outputs[7346] = ~((layer0_outputs[6451]) ^ (layer0_outputs[6245]));
    assign outputs[7347] = ~((layer0_outputs[8428]) ^ (layer0_outputs[9979]));
    assign outputs[7348] = (layer0_outputs[8067]) ^ (layer0_outputs[3227]);
    assign outputs[7349] = layer0_outputs[7937];
    assign outputs[7350] = ~(layer0_outputs[2223]) | (layer0_outputs[5925]);
    assign outputs[7351] = (layer0_outputs[4881]) & ~(layer0_outputs[9200]);
    assign outputs[7352] = (layer0_outputs[6741]) ^ (layer0_outputs[7651]);
    assign outputs[7353] = (layer0_outputs[514]) | (layer0_outputs[3938]);
    assign outputs[7354] = ~(layer0_outputs[2121]);
    assign outputs[7355] = ~(layer0_outputs[7817]);
    assign outputs[7356] = (layer0_outputs[8874]) | (layer0_outputs[3001]);
    assign outputs[7357] = (layer0_outputs[7378]) & (layer0_outputs[2670]);
    assign outputs[7358] = ~(layer0_outputs[6803]);
    assign outputs[7359] = (layer0_outputs[550]) & (layer0_outputs[7830]);
    assign outputs[7360] = (layer0_outputs[5306]) & (layer0_outputs[7182]);
    assign outputs[7361] = ~((layer0_outputs[105]) & (layer0_outputs[30]));
    assign outputs[7362] = (layer0_outputs[3935]) & ~(layer0_outputs[6213]);
    assign outputs[7363] = (layer0_outputs[106]) & ~(layer0_outputs[9682]);
    assign outputs[7364] = (layer0_outputs[6009]) & ~(layer0_outputs[2449]);
    assign outputs[7365] = ~((layer0_outputs[8915]) ^ (layer0_outputs[2783]));
    assign outputs[7366] = layer0_outputs[7891];
    assign outputs[7367] = ~((layer0_outputs[7583]) ^ (layer0_outputs[8492]));
    assign outputs[7368] = ~(layer0_outputs[3867]);
    assign outputs[7369] = (layer0_outputs[9319]) & ~(layer0_outputs[6987]);
    assign outputs[7370] = ~((layer0_outputs[5760]) ^ (layer0_outputs[964]));
    assign outputs[7371] = layer0_outputs[9684];
    assign outputs[7372] = (layer0_outputs[6661]) & (layer0_outputs[1191]);
    assign outputs[7373] = (layer0_outputs[526]) & ~(layer0_outputs[540]);
    assign outputs[7374] = (layer0_outputs[8166]) ^ (layer0_outputs[7092]);
    assign outputs[7375] = (layer0_outputs[2246]) ^ (layer0_outputs[6461]);
    assign outputs[7376] = layer0_outputs[4361];
    assign outputs[7377] = layer0_outputs[1663];
    assign outputs[7378] = (layer0_outputs[463]) ^ (layer0_outputs[9718]);
    assign outputs[7379] = ~(layer0_outputs[8491]);
    assign outputs[7380] = ~((layer0_outputs[4577]) | (layer0_outputs[2958]));
    assign outputs[7381] = (layer0_outputs[4961]) & ~(layer0_outputs[2623]);
    assign outputs[7382] = 1'b0;
    assign outputs[7383] = ~(layer0_outputs[8208]);
    assign outputs[7384] = (layer0_outputs[5665]) & ~(layer0_outputs[1588]);
    assign outputs[7385] = ~(layer0_outputs[5057]);
    assign outputs[7386] = (layer0_outputs[2475]) & ~(layer0_outputs[3869]);
    assign outputs[7387] = ~(layer0_outputs[6437]);
    assign outputs[7388] = layer0_outputs[8338];
    assign outputs[7389] = (layer0_outputs[1607]) & (layer0_outputs[472]);
    assign outputs[7390] = (layer0_outputs[5466]) & ~(layer0_outputs[5367]);
    assign outputs[7391] = ~(layer0_outputs[9989]);
    assign outputs[7392] = ~(layer0_outputs[193]);
    assign outputs[7393] = ~((layer0_outputs[2586]) & (layer0_outputs[8109]));
    assign outputs[7394] = ~(layer0_outputs[6961]);
    assign outputs[7395] = ~(layer0_outputs[4069]) | (layer0_outputs[3781]);
    assign outputs[7396] = (layer0_outputs[7832]) & (layer0_outputs[7533]);
    assign outputs[7397] = (layer0_outputs[8999]) & ~(layer0_outputs[9470]);
    assign outputs[7398] = ~(layer0_outputs[7936]);
    assign outputs[7399] = (layer0_outputs[7502]) & ~(layer0_outputs[751]);
    assign outputs[7400] = (layer0_outputs[10040]) ^ (layer0_outputs[1876]);
    assign outputs[7401] = ~(layer0_outputs[63]);
    assign outputs[7402] = layer0_outputs[1663];
    assign outputs[7403] = (layer0_outputs[2123]) | (layer0_outputs[8403]);
    assign outputs[7404] = layer0_outputs[6063];
    assign outputs[7405] = layer0_outputs[4074];
    assign outputs[7406] = (layer0_outputs[7100]) ^ (layer0_outputs[5293]);
    assign outputs[7407] = ~((layer0_outputs[9446]) & (layer0_outputs[9711]));
    assign outputs[7408] = ~(layer0_outputs[4158]);
    assign outputs[7409] = ~((layer0_outputs[8485]) ^ (layer0_outputs[1015]));
    assign outputs[7410] = layer0_outputs[8471];
    assign outputs[7411] = ~(layer0_outputs[7345]) | (layer0_outputs[8840]);
    assign outputs[7412] = ~(layer0_outputs[8994]);
    assign outputs[7413] = ~(layer0_outputs[10019]);
    assign outputs[7414] = ~(layer0_outputs[753]);
    assign outputs[7415] = ~(layer0_outputs[255]);
    assign outputs[7416] = ~((layer0_outputs[2605]) ^ (layer0_outputs[8291]));
    assign outputs[7417] = ~(layer0_outputs[8400]);
    assign outputs[7418] = (layer0_outputs[5526]) & ~(layer0_outputs[1919]);
    assign outputs[7419] = ~(layer0_outputs[5013]);
    assign outputs[7420] = ~((layer0_outputs[702]) ^ (layer0_outputs[2932]));
    assign outputs[7421] = (layer0_outputs[1485]) ^ (layer0_outputs[10035]);
    assign outputs[7422] = (layer0_outputs[1383]) ^ (layer0_outputs[3561]);
    assign outputs[7423] = ~(layer0_outputs[3235]);
    assign outputs[7424] = ~(layer0_outputs[193]);
    assign outputs[7425] = (layer0_outputs[2401]) & (layer0_outputs[4216]);
    assign outputs[7426] = ~((layer0_outputs[1827]) | (layer0_outputs[9304]));
    assign outputs[7427] = ~(layer0_outputs[9658]);
    assign outputs[7428] = layer0_outputs[3476];
    assign outputs[7429] = ~(layer0_outputs[9959]);
    assign outputs[7430] = layer0_outputs[6516];
    assign outputs[7431] = (layer0_outputs[742]) & ~(layer0_outputs[2455]);
    assign outputs[7432] = ~(layer0_outputs[2348]);
    assign outputs[7433] = ~(layer0_outputs[2380]) | (layer0_outputs[8789]);
    assign outputs[7434] = layer0_outputs[4576];
    assign outputs[7435] = ~(layer0_outputs[4687]);
    assign outputs[7436] = layer0_outputs[6900];
    assign outputs[7437] = ~(layer0_outputs[575]);
    assign outputs[7438] = ~(layer0_outputs[9842]);
    assign outputs[7439] = (layer0_outputs[5554]) & ~(layer0_outputs[4127]);
    assign outputs[7440] = layer0_outputs[2359];
    assign outputs[7441] = layer0_outputs[4742];
    assign outputs[7442] = layer0_outputs[9032];
    assign outputs[7443] = ~(layer0_outputs[2259]);
    assign outputs[7444] = layer0_outputs[10225];
    assign outputs[7445] = layer0_outputs[4149];
    assign outputs[7446] = ~(layer0_outputs[9050]);
    assign outputs[7447] = (layer0_outputs[1131]) ^ (layer0_outputs[4277]);
    assign outputs[7448] = ~((layer0_outputs[6076]) | (layer0_outputs[9962]));
    assign outputs[7449] = ~(layer0_outputs[6766]);
    assign outputs[7450] = (layer0_outputs[1184]) & (layer0_outputs[2071]);
    assign outputs[7451] = ~(layer0_outputs[8280]);
    assign outputs[7452] = ~(layer0_outputs[1075]);
    assign outputs[7453] = layer0_outputs[7179];
    assign outputs[7454] = ~(layer0_outputs[9291]);
    assign outputs[7455] = (layer0_outputs[61]) & (layer0_outputs[302]);
    assign outputs[7456] = (layer0_outputs[8763]) & (layer0_outputs[9892]);
    assign outputs[7457] = (layer0_outputs[3554]) & ~(layer0_outputs[6043]);
    assign outputs[7458] = layer0_outputs[490];
    assign outputs[7459] = (layer0_outputs[1018]) | (layer0_outputs[3176]);
    assign outputs[7460] = ~(layer0_outputs[4121]) | (layer0_outputs[4395]);
    assign outputs[7461] = layer0_outputs[7987];
    assign outputs[7462] = (layer0_outputs[3276]) & ~(layer0_outputs[1127]);
    assign outputs[7463] = (layer0_outputs[5235]) ^ (layer0_outputs[1440]);
    assign outputs[7464] = (layer0_outputs[4895]) & ~(layer0_outputs[4991]);
    assign outputs[7465] = ~(layer0_outputs[3114]);
    assign outputs[7466] = ~((layer0_outputs[6189]) | (layer0_outputs[9105]));
    assign outputs[7467] = layer0_outputs[8504];
    assign outputs[7468] = ~((layer0_outputs[1744]) ^ (layer0_outputs[8904]));
    assign outputs[7469] = (layer0_outputs[7678]) & (layer0_outputs[8182]);
    assign outputs[7470] = ~(layer0_outputs[4412]);
    assign outputs[7471] = (layer0_outputs[9832]) & ~(layer0_outputs[9419]);
    assign outputs[7472] = (layer0_outputs[4692]) & (layer0_outputs[5843]);
    assign outputs[7473] = (layer0_outputs[5567]) & ~(layer0_outputs[1867]);
    assign outputs[7474] = ~(layer0_outputs[2985]);
    assign outputs[7475] = layer0_outputs[7805];
    assign outputs[7476] = ~((layer0_outputs[6625]) | (layer0_outputs[7011]));
    assign outputs[7477] = ~((layer0_outputs[6858]) | (layer0_outputs[6411]));
    assign outputs[7478] = (layer0_outputs[1167]) ^ (layer0_outputs[1487]);
    assign outputs[7479] = (layer0_outputs[7850]) | (layer0_outputs[1501]);
    assign outputs[7480] = (layer0_outputs[4021]) | (layer0_outputs[2172]);
    assign outputs[7481] = (layer0_outputs[10110]) ^ (layer0_outputs[4003]);
    assign outputs[7482] = layer0_outputs[7958];
    assign outputs[7483] = (layer0_outputs[7649]) & (layer0_outputs[9846]);
    assign outputs[7484] = layer0_outputs[10210];
    assign outputs[7485] = (layer0_outputs[4929]) & ~(layer0_outputs[3465]);
    assign outputs[7486] = (layer0_outputs[4497]) ^ (layer0_outputs[9283]);
    assign outputs[7487] = ~(layer0_outputs[7948]) | (layer0_outputs[595]);
    assign outputs[7488] = (layer0_outputs[3624]) & ~(layer0_outputs[4083]);
    assign outputs[7489] = layer0_outputs[2585];
    assign outputs[7490] = layer0_outputs[8991];
    assign outputs[7491] = ~(layer0_outputs[6656]);
    assign outputs[7492] = ~(layer0_outputs[8561]);
    assign outputs[7493] = (layer0_outputs[2166]) & ~(layer0_outputs[7515]);
    assign outputs[7494] = ~(layer0_outputs[3718]);
    assign outputs[7495] = ~(layer0_outputs[3662]);
    assign outputs[7496] = ~((layer0_outputs[8286]) & (layer0_outputs[8818]));
    assign outputs[7497] = ~(layer0_outputs[7998]);
    assign outputs[7498] = ~(layer0_outputs[5189]);
    assign outputs[7499] = (layer0_outputs[7714]) ^ (layer0_outputs[10184]);
    assign outputs[7500] = ~(layer0_outputs[1495]);
    assign outputs[7501] = layer0_outputs[423];
    assign outputs[7502] = ~((layer0_outputs[6526]) ^ (layer0_outputs[8598]));
    assign outputs[7503] = (layer0_outputs[3601]) ^ (layer0_outputs[7188]);
    assign outputs[7504] = (layer0_outputs[4166]) & ~(layer0_outputs[819]);
    assign outputs[7505] = ~(layer0_outputs[9632]);
    assign outputs[7506] = layer0_outputs[3138];
    assign outputs[7507] = (layer0_outputs[9041]) & ~(layer0_outputs[1636]);
    assign outputs[7508] = ~(layer0_outputs[525]);
    assign outputs[7509] = layer0_outputs[783];
    assign outputs[7510] = (layer0_outputs[9452]) & (layer0_outputs[5613]);
    assign outputs[7511] = (layer0_outputs[2610]) ^ (layer0_outputs[7546]);
    assign outputs[7512] = layer0_outputs[1903];
    assign outputs[7513] = (layer0_outputs[1951]) ^ (layer0_outputs[7035]);
    assign outputs[7514] = (layer0_outputs[5265]) & (layer0_outputs[7995]);
    assign outputs[7515] = layer0_outputs[9601];
    assign outputs[7516] = ~(layer0_outputs[591]);
    assign outputs[7517] = ~((layer0_outputs[4199]) ^ (layer0_outputs[2249]));
    assign outputs[7518] = ~((layer0_outputs[2206]) | (layer0_outputs[1516]));
    assign outputs[7519] = (layer0_outputs[5020]) | (layer0_outputs[9045]);
    assign outputs[7520] = ~(layer0_outputs[4139]);
    assign outputs[7521] = layer0_outputs[3753];
    assign outputs[7522] = layer0_outputs[7376];
    assign outputs[7523] = (layer0_outputs[1546]) & ~(layer0_outputs[194]);
    assign outputs[7524] = layer0_outputs[2149];
    assign outputs[7525] = layer0_outputs[2855];
    assign outputs[7526] = ~((layer0_outputs[2344]) ^ (layer0_outputs[24]));
    assign outputs[7527] = (layer0_outputs[7416]) & ~(layer0_outputs[4861]);
    assign outputs[7528] = ~(layer0_outputs[963]);
    assign outputs[7529] = ~((layer0_outputs[2358]) | (layer0_outputs[3595]));
    assign outputs[7530] = layer0_outputs[8000];
    assign outputs[7531] = (layer0_outputs[917]) & ~(layer0_outputs[10113]);
    assign outputs[7532] = layer0_outputs[7855];
    assign outputs[7533] = (layer0_outputs[5018]) & ~(layer0_outputs[5401]);
    assign outputs[7534] = ~(layer0_outputs[6654]) | (layer0_outputs[7359]);
    assign outputs[7535] = (layer0_outputs[3823]) & ~(layer0_outputs[5179]);
    assign outputs[7536] = ~(layer0_outputs[1556]);
    assign outputs[7537] = ~((layer0_outputs[7732]) | (layer0_outputs[5024]));
    assign outputs[7538] = ~((layer0_outputs[2226]) | (layer0_outputs[1298]));
    assign outputs[7539] = ~(layer0_outputs[8229]);
    assign outputs[7540] = ~((layer0_outputs[1153]) | (layer0_outputs[6004]));
    assign outputs[7541] = ~((layer0_outputs[3565]) ^ (layer0_outputs[3640]));
    assign outputs[7542] = layer0_outputs[4665];
    assign outputs[7543] = (layer0_outputs[5626]) & ~(layer0_outputs[10134]);
    assign outputs[7544] = ~(layer0_outputs[1540]);
    assign outputs[7545] = (layer0_outputs[2180]) & ~(layer0_outputs[603]);
    assign outputs[7546] = layer0_outputs[8039];
    assign outputs[7547] = (layer0_outputs[8853]) & (layer0_outputs[6313]);
    assign outputs[7548] = (layer0_outputs[10104]) & (layer0_outputs[4152]);
    assign outputs[7549] = ~((layer0_outputs[1335]) ^ (layer0_outputs[9479]));
    assign outputs[7550] = layer0_outputs[89];
    assign outputs[7551] = (layer0_outputs[7410]) & (layer0_outputs[9608]);
    assign outputs[7552] = ~(layer0_outputs[8823]);
    assign outputs[7553] = ~(layer0_outputs[6733]);
    assign outputs[7554] = (layer0_outputs[264]) & ~(layer0_outputs[9956]);
    assign outputs[7555] = layer0_outputs[4496];
    assign outputs[7556] = ~((layer0_outputs[2565]) ^ (layer0_outputs[4326]));
    assign outputs[7557] = (layer0_outputs[7414]) & ~(layer0_outputs[2435]);
    assign outputs[7558] = (layer0_outputs[6153]) | (layer0_outputs[9294]);
    assign outputs[7559] = layer0_outputs[6866];
    assign outputs[7560] = ~(layer0_outputs[8684]);
    assign outputs[7561] = (layer0_outputs[1215]) & ~(layer0_outputs[9671]);
    assign outputs[7562] = (layer0_outputs[5037]) & ~(layer0_outputs[9252]);
    assign outputs[7563] = ~(layer0_outputs[4670]);
    assign outputs[7564] = ~(layer0_outputs[8252]);
    assign outputs[7565] = layer0_outputs[4677];
    assign outputs[7566] = ~(layer0_outputs[2538]);
    assign outputs[7567] = layer0_outputs[6878];
    assign outputs[7568] = ~(layer0_outputs[4989]);
    assign outputs[7569] = ~((layer0_outputs[2922]) ^ (layer0_outputs[2154]));
    assign outputs[7570] = (layer0_outputs[7148]) & ~(layer0_outputs[7058]);
    assign outputs[7571] = layer0_outputs[4954];
    assign outputs[7572] = layer0_outputs[4196];
    assign outputs[7573] = ~(layer0_outputs[3155]);
    assign outputs[7574] = (layer0_outputs[789]) & (layer0_outputs[2397]);
    assign outputs[7575] = (layer0_outputs[4920]) ^ (layer0_outputs[3203]);
    assign outputs[7576] = (layer0_outputs[8889]) & (layer0_outputs[7872]);
    assign outputs[7577] = (layer0_outputs[2149]) ^ (layer0_outputs[4410]);
    assign outputs[7578] = layer0_outputs[5010];
    assign outputs[7579] = ~((layer0_outputs[9981]) ^ (layer0_outputs[1904]));
    assign outputs[7580] = layer0_outputs[5462];
    assign outputs[7581] = layer0_outputs[1923];
    assign outputs[7582] = layer0_outputs[8042];
    assign outputs[7583] = (layer0_outputs[6466]) & ~(layer0_outputs[9267]);
    assign outputs[7584] = (layer0_outputs[5834]) ^ (layer0_outputs[7672]);
    assign outputs[7585] = ~(layer0_outputs[2747]);
    assign outputs[7586] = ~(layer0_outputs[8934]);
    assign outputs[7587] = (layer0_outputs[3672]) & (layer0_outputs[1309]);
    assign outputs[7588] = layer0_outputs[5193];
    assign outputs[7589] = layer0_outputs[8731];
    assign outputs[7590] = layer0_outputs[6053];
    assign outputs[7591] = ~(layer0_outputs[4967]);
    assign outputs[7592] = (layer0_outputs[8632]) ^ (layer0_outputs[7916]);
    assign outputs[7593] = ~(layer0_outputs[3477]);
    assign outputs[7594] = layer0_outputs[4793];
    assign outputs[7595] = ~(layer0_outputs[6758]) | (layer0_outputs[5341]);
    assign outputs[7596] = layer0_outputs[8619];
    assign outputs[7597] = ~((layer0_outputs[6559]) | (layer0_outputs[5343]));
    assign outputs[7598] = layer0_outputs[3041];
    assign outputs[7599] = ~(layer0_outputs[5772]);
    assign outputs[7600] = ~(layer0_outputs[7360]);
    assign outputs[7601] = layer0_outputs[2365];
    assign outputs[7602] = (layer0_outputs[1668]) ^ (layer0_outputs[7487]);
    assign outputs[7603] = ~(layer0_outputs[6815]);
    assign outputs[7604] = ~((layer0_outputs[7792]) | (layer0_outputs[5428]));
    assign outputs[7605] = (layer0_outputs[6771]) ^ (layer0_outputs[9300]);
    assign outputs[7606] = ~(layer0_outputs[6047]);
    assign outputs[7607] = ~(layer0_outputs[2967]);
    assign outputs[7608] = layer0_outputs[6475];
    assign outputs[7609] = (layer0_outputs[9145]) & ~(layer0_outputs[5430]);
    assign outputs[7610] = (layer0_outputs[5642]) & ~(layer0_outputs[10008]);
    assign outputs[7611] = ~(layer0_outputs[9466]);
    assign outputs[7612] = layer0_outputs[1118];
    assign outputs[7613] = (layer0_outputs[3819]) & ~(layer0_outputs[3972]);
    assign outputs[7614] = ~(layer0_outputs[3818]);
    assign outputs[7615] = ~(layer0_outputs[2491]);
    assign outputs[7616] = ~(layer0_outputs[3942]);
    assign outputs[7617] = layer0_outputs[4485];
    assign outputs[7618] = (layer0_outputs[4543]) ^ (layer0_outputs[6964]);
    assign outputs[7619] = ~(layer0_outputs[4774]) | (layer0_outputs[9825]);
    assign outputs[7620] = ~((layer0_outputs[1740]) ^ (layer0_outputs[9037]));
    assign outputs[7621] = (layer0_outputs[4191]) & ~(layer0_outputs[2974]);
    assign outputs[7622] = layer0_outputs[9384];
    assign outputs[7623] = layer0_outputs[7477];
    assign outputs[7624] = layer0_outputs[7729];
    assign outputs[7625] = ~(layer0_outputs[6963]);
    assign outputs[7626] = layer0_outputs[2365];
    assign outputs[7627] = ~(layer0_outputs[1437]);
    assign outputs[7628] = ~(layer0_outputs[8088]);
    assign outputs[7629] = ~(layer0_outputs[4716]);
    assign outputs[7630] = (layer0_outputs[5726]) & (layer0_outputs[9023]);
    assign outputs[7631] = (layer0_outputs[6913]) & ~(layer0_outputs[6233]);
    assign outputs[7632] = ~(layer0_outputs[7403]);
    assign outputs[7633] = (layer0_outputs[4601]) & (layer0_outputs[5922]);
    assign outputs[7634] = (layer0_outputs[4404]) & ~(layer0_outputs[40]);
    assign outputs[7635] = layer0_outputs[5399];
    assign outputs[7636] = (layer0_outputs[4484]) & ~(layer0_outputs[704]);
    assign outputs[7637] = layer0_outputs[7460];
    assign outputs[7638] = (layer0_outputs[3702]) & (layer0_outputs[8540]);
    assign outputs[7639] = ~(layer0_outputs[8643]) | (layer0_outputs[608]);
    assign outputs[7640] = (layer0_outputs[3556]) ^ (layer0_outputs[10032]);
    assign outputs[7641] = ~(layer0_outputs[4841]);
    assign outputs[7642] = ~((layer0_outputs[5032]) ^ (layer0_outputs[7119]));
    assign outputs[7643] = (layer0_outputs[3944]) & ~(layer0_outputs[1329]);
    assign outputs[7644] = (layer0_outputs[8762]) & ~(layer0_outputs[2860]);
    assign outputs[7645] = (layer0_outputs[8048]) & ~(layer0_outputs[9833]);
    assign outputs[7646] = ~(layer0_outputs[10194]);
    assign outputs[7647] = (layer0_outputs[2004]) & (layer0_outputs[1728]);
    assign outputs[7648] = layer0_outputs[9324];
    assign outputs[7649] = ~(layer0_outputs[5294]);
    assign outputs[7650] = ~(layer0_outputs[9974]);
    assign outputs[7651] = layer0_outputs[537];
    assign outputs[7652] = layer0_outputs[3968];
    assign outputs[7653] = (layer0_outputs[2646]) & ~(layer0_outputs[6897]);
    assign outputs[7654] = (layer0_outputs[4527]) & (layer0_outputs[10014]);
    assign outputs[7655] = (layer0_outputs[1378]) ^ (layer0_outputs[8428]);
    assign outputs[7656] = ~(layer0_outputs[3823]);
    assign outputs[7657] = (layer0_outputs[2184]) & (layer0_outputs[6751]);
    assign outputs[7658] = (layer0_outputs[7874]) & ~(layer0_outputs[7176]);
    assign outputs[7659] = layer0_outputs[7681];
    assign outputs[7660] = ~((layer0_outputs[2825]) ^ (layer0_outputs[6712]));
    assign outputs[7661] = ~(layer0_outputs[8716]);
    assign outputs[7662] = (layer0_outputs[4415]) & ~(layer0_outputs[1071]);
    assign outputs[7663] = layer0_outputs[2472];
    assign outputs[7664] = ~(layer0_outputs[7956]);
    assign outputs[7665] = layer0_outputs[4038];
    assign outputs[7666] = ~((layer0_outputs[7836]) ^ (layer0_outputs[5361]));
    assign outputs[7667] = (layer0_outputs[733]) & ~(layer0_outputs[8997]);
    assign outputs[7668] = ~((layer0_outputs[5963]) ^ (layer0_outputs[4834]));
    assign outputs[7669] = layer0_outputs[5957];
    assign outputs[7670] = (layer0_outputs[2050]) & (layer0_outputs[4009]);
    assign outputs[7671] = ~((layer0_outputs[6806]) | (layer0_outputs[6690]));
    assign outputs[7672] = (layer0_outputs[3193]) & ~(layer0_outputs[1951]);
    assign outputs[7673] = (layer0_outputs[8271]) ^ (layer0_outputs[3189]);
    assign outputs[7674] = (layer0_outputs[7796]) ^ (layer0_outputs[7810]);
    assign outputs[7675] = ~((layer0_outputs[6971]) | (layer0_outputs[8849]));
    assign outputs[7676] = (layer0_outputs[9272]) ^ (layer0_outputs[1206]);
    assign outputs[7677] = layer0_outputs[7009];
    assign outputs[7678] = layer0_outputs[7852];
    assign outputs[7679] = (layer0_outputs[854]) ^ (layer0_outputs[7455]);
    assign outputs[7680] = ~(layer0_outputs[9502]);
    assign outputs[7681] = (layer0_outputs[2445]) & ~(layer0_outputs[7206]);
    assign outputs[7682] = layer0_outputs[9984];
    assign outputs[7683] = (layer0_outputs[1056]) & (layer0_outputs[3819]);
    assign outputs[7684] = ~((layer0_outputs[4689]) | (layer0_outputs[962]));
    assign outputs[7685] = (layer0_outputs[4583]) & ~(layer0_outputs[6735]);
    assign outputs[7686] = ~(layer0_outputs[2886]) | (layer0_outputs[8956]);
    assign outputs[7687] = layer0_outputs[6038];
    assign outputs[7688] = layer0_outputs[8509];
    assign outputs[7689] = ~(layer0_outputs[6383]);
    assign outputs[7690] = ~(layer0_outputs[8014]);
    assign outputs[7691] = ~(layer0_outputs[8470]);
    assign outputs[7692] = layer0_outputs[3170];
    assign outputs[7693] = layer0_outputs[4724];
    assign outputs[7694] = (layer0_outputs[5295]) ^ (layer0_outputs[8416]);
    assign outputs[7695] = ~(layer0_outputs[9890]);
    assign outputs[7696] = ~(layer0_outputs[3551]);
    assign outputs[7697] = ~(layer0_outputs[8266]);
    assign outputs[7698] = layer0_outputs[1847];
    assign outputs[7699] = layer0_outputs[9827];
    assign outputs[7700] = ~(layer0_outputs[5403]);
    assign outputs[7701] = ~((layer0_outputs[4597]) | (layer0_outputs[6335]));
    assign outputs[7702] = ~(layer0_outputs[2710]);
    assign outputs[7703] = (layer0_outputs[6120]) & ~(layer0_outputs[2924]);
    assign outputs[7704] = layer0_outputs[9297];
    assign outputs[7705] = ~(layer0_outputs[4169]);
    assign outputs[7706] = (layer0_outputs[3193]) & ~(layer0_outputs[2773]);
    assign outputs[7707] = ~(layer0_outputs[953]);
    assign outputs[7708] = layer0_outputs[7683];
    assign outputs[7709] = ~(layer0_outputs[6679]);
    assign outputs[7710] = (layer0_outputs[4835]) & ~(layer0_outputs[4917]);
    assign outputs[7711] = (layer0_outputs[6214]) ^ (layer0_outputs[3889]);
    assign outputs[7712] = ~(layer0_outputs[10143]);
    assign outputs[7713] = layer0_outputs[3545];
    assign outputs[7714] = layer0_outputs[6615];
    assign outputs[7715] = layer0_outputs[6266];
    assign outputs[7716] = ~((layer0_outputs[2890]) | (layer0_outputs[6864]));
    assign outputs[7717] = ~(layer0_outputs[5684]);
    assign outputs[7718] = ~(layer0_outputs[2208]);
    assign outputs[7719] = ~(layer0_outputs[9449]);
    assign outputs[7720] = layer0_outputs[497];
    assign outputs[7721] = (layer0_outputs[3261]) & ~(layer0_outputs[4580]);
    assign outputs[7722] = layer0_outputs[10235];
    assign outputs[7723] = (layer0_outputs[5928]) & ~(layer0_outputs[7139]);
    assign outputs[7724] = ~((layer0_outputs[7429]) | (layer0_outputs[2155]));
    assign outputs[7725] = layer0_outputs[9276];
    assign outputs[7726] = layer0_outputs[7531];
    assign outputs[7727] = ~(layer0_outputs[1158]);
    assign outputs[7728] = ~((layer0_outputs[8121]) | (layer0_outputs[2828]));
    assign outputs[7729] = ~((layer0_outputs[1992]) ^ (layer0_outputs[2862]));
    assign outputs[7730] = ~(layer0_outputs[8140]);
    assign outputs[7731] = layer0_outputs[5345];
    assign outputs[7732] = ~(layer0_outputs[8720]);
    assign outputs[7733] = ~(layer0_outputs[2001]);
    assign outputs[7734] = (layer0_outputs[1979]) & (layer0_outputs[9858]);
    assign outputs[7735] = layer0_outputs[5872];
    assign outputs[7736] = (layer0_outputs[3808]) ^ (layer0_outputs[7621]);
    assign outputs[7737] = ~((layer0_outputs[4341]) ^ (layer0_outputs[5007]));
    assign outputs[7738] = layer0_outputs[6968];
    assign outputs[7739] = (layer0_outputs[9613]) & ~(layer0_outputs[1403]);
    assign outputs[7740] = (layer0_outputs[6977]) & ~(layer0_outputs[8979]);
    assign outputs[7741] = (layer0_outputs[4383]) ^ (layer0_outputs[5930]);
    assign outputs[7742] = ~(layer0_outputs[4223]);
    assign outputs[7743] = (layer0_outputs[470]) | (layer0_outputs[371]);
    assign outputs[7744] = ~(layer0_outputs[8120]);
    assign outputs[7745] = (layer0_outputs[3535]) | (layer0_outputs[2419]);
    assign outputs[7746] = layer0_outputs[8785];
    assign outputs[7747] = (layer0_outputs[999]) & ~(layer0_outputs[6704]);
    assign outputs[7748] = layer0_outputs[5673];
    assign outputs[7749] = (layer0_outputs[7202]) ^ (layer0_outputs[1204]);
    assign outputs[7750] = (layer0_outputs[7765]) & ~(layer0_outputs[8322]);
    assign outputs[7751] = (layer0_outputs[3878]) & (layer0_outputs[8383]);
    assign outputs[7752] = ~((layer0_outputs[8207]) | (layer0_outputs[7092]));
    assign outputs[7753] = (layer0_outputs[9030]) ^ (layer0_outputs[972]);
    assign outputs[7754] = (layer0_outputs[8180]) & ~(layer0_outputs[6681]);
    assign outputs[7755] = ~((layer0_outputs[5667]) | (layer0_outputs[10037]));
    assign outputs[7756] = layer0_outputs[10125];
    assign outputs[7757] = layer0_outputs[667];
    assign outputs[7758] = layer0_outputs[2507];
    assign outputs[7759] = ~((layer0_outputs[1365]) & (layer0_outputs[7875]));
    assign outputs[7760] = ~(layer0_outputs[5041]);
    assign outputs[7761] = layer0_outputs[2941];
    assign outputs[7762] = ~((layer0_outputs[4610]) | (layer0_outputs[2506]));
    assign outputs[7763] = layer0_outputs[88];
    assign outputs[7764] = ~((layer0_outputs[7711]) ^ (layer0_outputs[5577]));
    assign outputs[7765] = ~(layer0_outputs[132]);
    assign outputs[7766] = (layer0_outputs[6201]) | (layer0_outputs[7718]);
    assign outputs[7767] = (layer0_outputs[530]) ^ (layer0_outputs[839]);
    assign outputs[7768] = ~((layer0_outputs[9739]) ^ (layer0_outputs[8859]));
    assign outputs[7769] = layer0_outputs[10152];
    assign outputs[7770] = layer0_outputs[9670];
    assign outputs[7771] = layer0_outputs[8852];
    assign outputs[7772] = ~(layer0_outputs[1072]);
    assign outputs[7773] = ~((layer0_outputs[3338]) ^ (layer0_outputs[8638]));
    assign outputs[7774] = ~(layer0_outputs[104]);
    assign outputs[7775] = ~(layer0_outputs[290]) | (layer0_outputs[3289]);
    assign outputs[7776] = layer0_outputs[9290];
    assign outputs[7777] = ~(layer0_outputs[5350]);
    assign outputs[7778] = layer0_outputs[788];
    assign outputs[7779] = (layer0_outputs[3436]) & ~(layer0_outputs[8423]);
    assign outputs[7780] = (layer0_outputs[4918]) ^ (layer0_outputs[2617]);
    assign outputs[7781] = (layer0_outputs[1249]) ^ (layer0_outputs[6212]);
    assign outputs[7782] = (layer0_outputs[6374]) & ~(layer0_outputs[8877]);
    assign outputs[7783] = (layer0_outputs[4641]) & ~(layer0_outputs[6673]);
    assign outputs[7784] = (layer0_outputs[3248]) ^ (layer0_outputs[5416]);
    assign outputs[7785] = ~((layer0_outputs[9430]) ^ (layer0_outputs[7701]));
    assign outputs[7786] = ~(layer0_outputs[1784]);
    assign outputs[7787] = layer0_outputs[5355];
    assign outputs[7788] = ~(layer0_outputs[79]);
    assign outputs[7789] = ~((layer0_outputs[4094]) | (layer0_outputs[1484]));
    assign outputs[7790] = (layer0_outputs[1721]) & ~(layer0_outputs[6139]);
    assign outputs[7791] = (layer0_outputs[1321]) & ~(layer0_outputs[8472]);
    assign outputs[7792] = ~((layer0_outputs[3218]) | (layer0_outputs[1950]));
    assign outputs[7793] = ~(layer0_outputs[2992]);
    assign outputs[7794] = (layer0_outputs[291]) ^ (layer0_outputs[5934]);
    assign outputs[7795] = (layer0_outputs[6608]) & ~(layer0_outputs[3881]);
    assign outputs[7796] = ~(layer0_outputs[3020]) | (layer0_outputs[7965]);
    assign outputs[7797] = ~(layer0_outputs[9958]);
    assign outputs[7798] = (layer0_outputs[7226]) ^ (layer0_outputs[7696]);
    assign outputs[7799] = (layer0_outputs[7795]) ^ (layer0_outputs[7256]);
    assign outputs[7800] = ~((layer0_outputs[4893]) | (layer0_outputs[797]));
    assign outputs[7801] = ~(layer0_outputs[7839]);
    assign outputs[7802] = layer0_outputs[5949];
    assign outputs[7803] = ~(layer0_outputs[6157]);
    assign outputs[7804] = ~(layer0_outputs[9287]);
    assign outputs[7805] = ~((layer0_outputs[2937]) | (layer0_outputs[9469]));
    assign outputs[7806] = ~((layer0_outputs[7959]) ^ (layer0_outputs[8815]));
    assign outputs[7807] = ~(layer0_outputs[3263]);
    assign outputs[7808] = ~((layer0_outputs[6243]) ^ (layer0_outputs[7351]));
    assign outputs[7809] = ~((layer0_outputs[9811]) ^ (layer0_outputs[1341]));
    assign outputs[7810] = layer0_outputs[1098];
    assign outputs[7811] = layer0_outputs[2268];
    assign outputs[7812] = ~(layer0_outputs[3629]);
    assign outputs[7813] = layer0_outputs[4868];
    assign outputs[7814] = layer0_outputs[8620];
    assign outputs[7815] = ~(layer0_outputs[8813]);
    assign outputs[7816] = (layer0_outputs[9983]) & ~(layer0_outputs[8040]);
    assign outputs[7817] = ~((layer0_outputs[1468]) ^ (layer0_outputs[8814]));
    assign outputs[7818] = ~(layer0_outputs[183]);
    assign outputs[7819] = (layer0_outputs[4289]) & ~(layer0_outputs[9751]);
    assign outputs[7820] = layer0_outputs[9271];
    assign outputs[7821] = (layer0_outputs[9778]) & ~(layer0_outputs[5286]);
    assign outputs[7822] = layer0_outputs[5708];
    assign outputs[7823] = layer0_outputs[4581];
    assign outputs[7824] = ~(layer0_outputs[7960]);
    assign outputs[7825] = ~(layer0_outputs[7432]);
    assign outputs[7826] = layer0_outputs[4879];
    assign outputs[7827] = (layer0_outputs[8157]) & ~(layer0_outputs[6646]);
    assign outputs[7828] = ~((layer0_outputs[3905]) ^ (layer0_outputs[4159]));
    assign outputs[7829] = (layer0_outputs[2293]) & ~(layer0_outputs[4374]);
    assign outputs[7830] = (layer0_outputs[2930]) & ~(layer0_outputs[3582]);
    assign outputs[7831] = layer0_outputs[3450];
    assign outputs[7832] = layer0_outputs[5278];
    assign outputs[7833] = ~(layer0_outputs[6400]) | (layer0_outputs[4389]);
    assign outputs[7834] = layer0_outputs[9086];
    assign outputs[7835] = layer0_outputs[137];
    assign outputs[7836] = (layer0_outputs[6217]) & ~(layer0_outputs[4220]);
    assign outputs[7837] = (layer0_outputs[6928]) & (layer0_outputs[7268]);
    assign outputs[7838] = layer0_outputs[3804];
    assign outputs[7839] = (layer0_outputs[144]) & ~(layer0_outputs[8672]);
    assign outputs[7840] = ~((layer0_outputs[7118]) ^ (layer0_outputs[2669]));
    assign outputs[7841] = layer0_outputs[1677];
    assign outputs[7842] = ~(layer0_outputs[6288]);
    assign outputs[7843] = layer0_outputs[10152];
    assign outputs[7844] = ~(layer0_outputs[7868]);
    assign outputs[7845] = ~((layer0_outputs[8880]) | (layer0_outputs[4981]));
    assign outputs[7846] = ~(layer0_outputs[1835]);
    assign outputs[7847] = (layer0_outputs[8654]) | (layer0_outputs[3759]);
    assign outputs[7848] = (layer0_outputs[7806]) & (layer0_outputs[5691]);
    assign outputs[7849] = (layer0_outputs[9678]) & ~(layer0_outputs[8554]);
    assign outputs[7850] = (layer0_outputs[9624]) & (layer0_outputs[196]);
    assign outputs[7851] = (layer0_outputs[7840]) & ~(layer0_outputs[10036]);
    assign outputs[7852] = ~(layer0_outputs[6137]);
    assign outputs[7853] = ~(layer0_outputs[7848]);
    assign outputs[7854] = ~(layer0_outputs[6569]) | (layer0_outputs[4418]);
    assign outputs[7855] = ~((layer0_outputs[1806]) ^ (layer0_outputs[7730]));
    assign outputs[7856] = layer0_outputs[7357];
    assign outputs[7857] = layer0_outputs[7807];
    assign outputs[7858] = layer0_outputs[2596];
    assign outputs[7859] = layer0_outputs[3758];
    assign outputs[7860] = ~(layer0_outputs[5809]);
    assign outputs[7861] = ~(layer0_outputs[8871]);
    assign outputs[7862] = layer0_outputs[3119];
    assign outputs[7863] = ~(layer0_outputs[6597]);
    assign outputs[7864] = ~((layer0_outputs[5868]) ^ (layer0_outputs[4299]));
    assign outputs[7865] = (layer0_outputs[3465]) & ~(layer0_outputs[603]);
    assign outputs[7866] = ~(layer0_outputs[1787]);
    assign outputs[7867] = ~(layer0_outputs[6428]);
    assign outputs[7868] = (layer0_outputs[5124]) & (layer0_outputs[922]);
    assign outputs[7869] = layer0_outputs[6771];
    assign outputs[7870] = (layer0_outputs[9757]) ^ (layer0_outputs[5539]);
    assign outputs[7871] = ~((layer0_outputs[9782]) | (layer0_outputs[3239]));
    assign outputs[7872] = (layer0_outputs[2280]) & ~(layer0_outputs[5982]);
    assign outputs[7873] = layer0_outputs[394];
    assign outputs[7874] = ~(layer0_outputs[7849]);
    assign outputs[7875] = (layer0_outputs[1188]) ^ (layer0_outputs[7530]);
    assign outputs[7876] = ~(layer0_outputs[5657]) | (layer0_outputs[7587]);
    assign outputs[7877] = ~(layer0_outputs[1327]);
    assign outputs[7878] = layer0_outputs[5251];
    assign outputs[7879] = ~(layer0_outputs[1846]) | (layer0_outputs[8149]);
    assign outputs[7880] = (layer0_outputs[1788]) & ~(layer0_outputs[6395]);
    assign outputs[7881] = (layer0_outputs[8283]) & ~(layer0_outputs[2142]);
    assign outputs[7882] = ~(layer0_outputs[7642]);
    assign outputs[7883] = ~((layer0_outputs[8969]) | (layer0_outputs[3833]));
    assign outputs[7884] = layer0_outputs[9870];
    assign outputs[7885] = layer0_outputs[9701];
    assign outputs[7886] = ~(layer0_outputs[6684]);
    assign outputs[7887] = layer0_outputs[7081];
    assign outputs[7888] = layer0_outputs[1626];
    assign outputs[7889] = layer0_outputs[3770];
    assign outputs[7890] = layer0_outputs[9580];
    assign outputs[7891] = (layer0_outputs[6972]) & (layer0_outputs[7893]);
    assign outputs[7892] = ~(layer0_outputs[3742]);
    assign outputs[7893] = ~((layer0_outputs[4855]) ^ (layer0_outputs[8235]));
    assign outputs[7894] = ~(layer0_outputs[1324]);
    assign outputs[7895] = ~((layer0_outputs[4854]) ^ (layer0_outputs[6091]));
    assign outputs[7896] = (layer0_outputs[5257]) & ~(layer0_outputs[8193]);
    assign outputs[7897] = layer0_outputs[2464];
    assign outputs[7898] = ~(layer0_outputs[6562]);
    assign outputs[7899] = ~(layer0_outputs[1276]);
    assign outputs[7900] = ~(layer0_outputs[4499]);
    assign outputs[7901] = (layer0_outputs[9756]) & ~(layer0_outputs[2229]);
    assign outputs[7902] = ~((layer0_outputs[2083]) ^ (layer0_outputs[2144]));
    assign outputs[7903] = layer0_outputs[8230];
    assign outputs[7904] = ~(layer0_outputs[243]);
    assign outputs[7905] = ~(layer0_outputs[6888]);
    assign outputs[7906] = (layer0_outputs[9210]) ^ (layer0_outputs[2662]);
    assign outputs[7907] = (layer0_outputs[4573]) ^ (layer0_outputs[10187]);
    assign outputs[7908] = (layer0_outputs[8961]) ^ (layer0_outputs[4850]);
    assign outputs[7909] = layer0_outputs[9192];
    assign outputs[7910] = (layer0_outputs[8081]) & ~(layer0_outputs[3740]);
    assign outputs[7911] = ~(layer0_outputs[234]);
    assign outputs[7912] = ~(layer0_outputs[1375]);
    assign outputs[7913] = ~(layer0_outputs[6992]);
    assign outputs[7914] = layer0_outputs[1587];
    assign outputs[7915] = ~(layer0_outputs[889]);
    assign outputs[7916] = (layer0_outputs[2861]) & ~(layer0_outputs[7781]);
    assign outputs[7917] = (layer0_outputs[701]) & ~(layer0_outputs[10027]);
    assign outputs[7918] = (layer0_outputs[9631]) & (layer0_outputs[9812]);
    assign outputs[7919] = layer0_outputs[1525];
    assign outputs[7920] = ~((layer0_outputs[8565]) | (layer0_outputs[8430]));
    assign outputs[7921] = ~(layer0_outputs[867]);
    assign outputs[7922] = (layer0_outputs[6098]) & ~(layer0_outputs[7547]);
    assign outputs[7923] = ~((layer0_outputs[6520]) ^ (layer0_outputs[3624]));
    assign outputs[7924] = ~(layer0_outputs[8607]);
    assign outputs[7925] = (layer0_outputs[3153]) ^ (layer0_outputs[1128]);
    assign outputs[7926] = (layer0_outputs[6799]) & ~(layer0_outputs[6734]);
    assign outputs[7927] = ~(layer0_outputs[6108]) | (layer0_outputs[3585]);
    assign outputs[7928] = ~((layer0_outputs[8364]) ^ (layer0_outputs[6244]));
    assign outputs[7929] = layer0_outputs[3827];
    assign outputs[7930] = layer0_outputs[8412];
    assign outputs[7931] = ~(layer0_outputs[6672]) | (layer0_outputs[1993]);
    assign outputs[7932] = ~(layer0_outputs[1406]);
    assign outputs[7933] = (layer0_outputs[3871]) ^ (layer0_outputs[3380]);
    assign outputs[7934] = layer0_outputs[3574];
    assign outputs[7935] = (layer0_outputs[9217]) & (layer0_outputs[13]);
    assign outputs[7936] = layer0_outputs[5977];
    assign outputs[7937] = layer0_outputs[640];
    assign outputs[7938] = ~((layer0_outputs[8705]) | (layer0_outputs[4013]));
    assign outputs[7939] = layer0_outputs[9333];
    assign outputs[7940] = ~(layer0_outputs[3047]);
    assign outputs[7941] = layer0_outputs[9979];
    assign outputs[7942] = layer0_outputs[4290];
    assign outputs[7943] = ~(layer0_outputs[6758]);
    assign outputs[7944] = ~(layer0_outputs[5659]);
    assign outputs[7945] = ~((layer0_outputs[1844]) ^ (layer0_outputs[5865]));
    assign outputs[7946] = ~(layer0_outputs[7191]);
    assign outputs[7947] = layer0_outputs[2345];
    assign outputs[7948] = (layer0_outputs[8786]) & ~(layer0_outputs[1131]);
    assign outputs[7949] = layer0_outputs[6460];
    assign outputs[7950] = ~(layer0_outputs[3562]);
    assign outputs[7951] = layer0_outputs[3826];
    assign outputs[7952] = (layer0_outputs[89]) & (layer0_outputs[7234]);
    assign outputs[7953] = ~(layer0_outputs[8488]) | (layer0_outputs[6297]);
    assign outputs[7954] = ~((layer0_outputs[2632]) | (layer0_outputs[5948]));
    assign outputs[7955] = layer0_outputs[8597];
    assign outputs[7956] = layer0_outputs[9953];
    assign outputs[7957] = ~((layer0_outputs[3993]) ^ (layer0_outputs[7755]));
    assign outputs[7958] = layer0_outputs[2305];
    assign outputs[7959] = ~(layer0_outputs[865]);
    assign outputs[7960] = (layer0_outputs[5386]) ^ (layer0_outputs[9356]);
    assign outputs[7961] = (layer0_outputs[5563]) & ~(layer0_outputs[9742]);
    assign outputs[7962] = (layer0_outputs[4422]) & ~(layer0_outputs[4477]);
    assign outputs[7963] = (layer0_outputs[5014]) ^ (layer0_outputs[1254]);
    assign outputs[7964] = (layer0_outputs[4828]) & (layer0_outputs[5629]);
    assign outputs[7965] = ~(layer0_outputs[3286]);
    assign outputs[7966] = ~(layer0_outputs[6305]);
    assign outputs[7967] = (layer0_outputs[7591]) ^ (layer0_outputs[5874]);
    assign outputs[7968] = ~(layer0_outputs[4510]);
    assign outputs[7969] = layer0_outputs[7895];
    assign outputs[7970] = ~((layer0_outputs[7464]) | (layer0_outputs[7172]));
    assign outputs[7971] = (layer0_outputs[6062]) & (layer0_outputs[7380]);
    assign outputs[7972] = (layer0_outputs[8703]) ^ (layer0_outputs[1259]);
    assign outputs[7973] = ~(layer0_outputs[9317]);
    assign outputs[7974] = (layer0_outputs[7238]) & ~(layer0_outputs[1837]);
    assign outputs[7975] = ~((layer0_outputs[7871]) ^ (layer0_outputs[5224]));
    assign outputs[7976] = (layer0_outputs[8288]) | (layer0_outputs[8819]);
    assign outputs[7977] = ~(layer0_outputs[2934]);
    assign outputs[7978] = layer0_outputs[7320];
    assign outputs[7979] = layer0_outputs[8555];
    assign outputs[7980] = (layer0_outputs[2936]) & ~(layer0_outputs[172]);
    assign outputs[7981] = ~((layer0_outputs[9570]) | (layer0_outputs[4344]));
    assign outputs[7982] = ~(layer0_outputs[3047]);
    assign outputs[7983] = layer0_outputs[5680];
    assign outputs[7984] = layer0_outputs[1263];
    assign outputs[7985] = (layer0_outputs[8096]) ^ (layer0_outputs[6785]);
    assign outputs[7986] = ~(layer0_outputs[5879]) | (layer0_outputs[8111]);
    assign outputs[7987] = ~(layer0_outputs[2802]);
    assign outputs[7988] = ~(layer0_outputs[5276]);
    assign outputs[7989] = layer0_outputs[5722];
    assign outputs[7990] = ~((layer0_outputs[4085]) | (layer0_outputs[3058]));
    assign outputs[7991] = (layer0_outputs[1469]) ^ (layer0_outputs[4875]);
    assign outputs[7992] = ~(layer0_outputs[122]);
    assign outputs[7993] = layer0_outputs[1032];
    assign outputs[7994] = ~(layer0_outputs[2766]);
    assign outputs[7995] = ~(layer0_outputs[3224]);
    assign outputs[7996] = layer0_outputs[8475];
    assign outputs[7997] = (layer0_outputs[2630]) ^ (layer0_outputs[9388]);
    assign outputs[7998] = ~((layer0_outputs[6123]) ^ (layer0_outputs[7099]));
    assign outputs[7999] = layer0_outputs[6900];
    assign outputs[8000] = layer0_outputs[4078];
    assign outputs[8001] = layer0_outputs[1747];
    assign outputs[8002] = ~(layer0_outputs[3447]);
    assign outputs[8003] = ~(layer0_outputs[3250]);
    assign outputs[8004] = ~((layer0_outputs[9806]) | (layer0_outputs[2432]));
    assign outputs[8005] = ~((layer0_outputs[5064]) | (layer0_outputs[3714]));
    assign outputs[8006] = ~(layer0_outputs[5857]) | (layer0_outputs[6896]);
    assign outputs[8007] = ~(layer0_outputs[1730]);
    assign outputs[8008] = ~((layer0_outputs[1000]) & (layer0_outputs[2826]));
    assign outputs[8009] = ~(layer0_outputs[7622]);
    assign outputs[8010] = layer0_outputs[1207];
    assign outputs[8011] = ~(layer0_outputs[2301]);
    assign outputs[8012] = layer0_outputs[4605];
    assign outputs[8013] = layer0_outputs[3267];
    assign outputs[8014] = ~(layer0_outputs[6178]);
    assign outputs[8015] = layer0_outputs[4708];
    assign outputs[8016] = ~((layer0_outputs[3629]) | (layer0_outputs[2390]));
    assign outputs[8017] = layer0_outputs[10118];
    assign outputs[8018] = (layer0_outputs[6864]) ^ (layer0_outputs[3422]);
    assign outputs[8019] = (layer0_outputs[3895]) & ~(layer0_outputs[422]);
    assign outputs[8020] = (layer0_outputs[9847]) & ~(layer0_outputs[7834]);
    assign outputs[8021] = (layer0_outputs[7315]) & (layer0_outputs[7992]);
    assign outputs[8022] = (layer0_outputs[8111]) & ~(layer0_outputs[6787]);
    assign outputs[8023] = ~((layer0_outputs[2760]) ^ (layer0_outputs[2646]));
    assign outputs[8024] = ~((layer0_outputs[4302]) | (layer0_outputs[3862]));
    assign outputs[8025] = ~(layer0_outputs[9845]);
    assign outputs[8026] = layer0_outputs[434];
    assign outputs[8027] = (layer0_outputs[158]) ^ (layer0_outputs[8034]);
    assign outputs[8028] = ~(layer0_outputs[10105]);
    assign outputs[8029] = ~(layer0_outputs[6495]);
    assign outputs[8030] = (layer0_outputs[8127]) & ~(layer0_outputs[7967]);
    assign outputs[8031] = ~(layer0_outputs[3106]);
    assign outputs[8032] = (layer0_outputs[9118]) ^ (layer0_outputs[6584]);
    assign outputs[8033] = layer0_outputs[5748];
    assign outputs[8034] = (layer0_outputs[7888]) & ~(layer0_outputs[3239]);
    assign outputs[8035] = (layer0_outputs[8314]) & (layer0_outputs[7821]);
    assign outputs[8036] = layer0_outputs[1501];
    assign outputs[8037] = (layer0_outputs[1662]) & (layer0_outputs[6774]);
    assign outputs[8038] = ~((layer0_outputs[1068]) ^ (layer0_outputs[6716]));
    assign outputs[8039] = (layer0_outputs[5116]) & ~(layer0_outputs[6743]);
    assign outputs[8040] = layer0_outputs[6163];
    assign outputs[8041] = (layer0_outputs[8408]) ^ (layer0_outputs[5365]);
    assign outputs[8042] = layer0_outputs[2839];
    assign outputs[8043] = ~((layer0_outputs[3079]) | (layer0_outputs[7065]));
    assign outputs[8044] = ~(layer0_outputs[8240]) | (layer0_outputs[8365]);
    assign outputs[8045] = layer0_outputs[10056];
    assign outputs[8046] = layer0_outputs[5768];
    assign outputs[8047] = (layer0_outputs[8868]) & ~(layer0_outputs[3797]);
    assign outputs[8048] = ~(layer0_outputs[4820]);
    assign outputs[8049] = layer0_outputs[9980];
    assign outputs[8050] = ~(layer0_outputs[4860]);
    assign outputs[8051] = ~(layer0_outputs[5280]);
    assign outputs[8052] = layer0_outputs[3613];
    assign outputs[8053] = layer0_outputs[8443];
    assign outputs[8054] = ~(layer0_outputs[7158]);
    assign outputs[8055] = (layer0_outputs[3398]) & ~(layer0_outputs[9358]);
    assign outputs[8056] = ~((layer0_outputs[7329]) ^ (layer0_outputs[1849]));
    assign outputs[8057] = (layer0_outputs[5613]) & (layer0_outputs[6832]);
    assign outputs[8058] = layer0_outputs[2767];
    assign outputs[8059] = ~((layer0_outputs[3157]) ^ (layer0_outputs[7700]));
    assign outputs[8060] = layer0_outputs[5901];
    assign outputs[8061] = layer0_outputs[8700];
    assign outputs[8062] = ~((layer0_outputs[1497]) | (layer0_outputs[1597]));
    assign outputs[8063] = layer0_outputs[7219];
    assign outputs[8064] = ~(layer0_outputs[5137]);
    assign outputs[8065] = ~(layer0_outputs[980]);
    assign outputs[8066] = ~(layer0_outputs[8019]);
    assign outputs[8067] = ~(layer0_outputs[9000]);
    assign outputs[8068] = ~(layer0_outputs[7077]) | (layer0_outputs[9337]);
    assign outputs[8069] = ~(layer0_outputs[8110]);
    assign outputs[8070] = (layer0_outputs[8753]) & (layer0_outputs[28]);
    assign outputs[8071] = (layer0_outputs[1428]) ^ (layer0_outputs[5168]);
    assign outputs[8072] = (layer0_outputs[6326]) & ~(layer0_outputs[4836]);
    assign outputs[8073] = ~(layer0_outputs[1467]);
    assign outputs[8074] = ~((layer0_outputs[9094]) & (layer0_outputs[1852]));
    assign outputs[8075] = ~((layer0_outputs[6360]) & (layer0_outputs[3743]));
    assign outputs[8076] = ~((layer0_outputs[3937]) ^ (layer0_outputs[1843]));
    assign outputs[8077] = ~((layer0_outputs[802]) & (layer0_outputs[4411]));
    assign outputs[8078] = layer0_outputs[2427];
    assign outputs[8079] = layer0_outputs[6462];
    assign outputs[8080] = (layer0_outputs[9709]) ^ (layer0_outputs[7432]);
    assign outputs[8081] = ~((layer0_outputs[4816]) & (layer0_outputs[2600]));
    assign outputs[8082] = (layer0_outputs[537]) & ~(layer0_outputs[4814]);
    assign outputs[8083] = ~(layer0_outputs[6202]);
    assign outputs[8084] = ~(layer0_outputs[4135]);
    assign outputs[8085] = ~((layer0_outputs[2214]) ^ (layer0_outputs[6532]));
    assign outputs[8086] = (layer0_outputs[2028]) ^ (layer0_outputs[777]);
    assign outputs[8087] = ~((layer0_outputs[5919]) | (layer0_outputs[1075]));
    assign outputs[8088] = ~(layer0_outputs[5501]) | (layer0_outputs[2534]);
    assign outputs[8089] = layer0_outputs[4867];
    assign outputs[8090] = ~(layer0_outputs[9154]);
    assign outputs[8091] = ~(layer0_outputs[1569]);
    assign outputs[8092] = (layer0_outputs[4752]) & ~(layer0_outputs[2218]);
    assign outputs[8093] = (layer0_outputs[9571]) ^ (layer0_outputs[8489]);
    assign outputs[8094] = (layer0_outputs[5596]) ^ (layer0_outputs[9537]);
    assign outputs[8095] = ~(layer0_outputs[679]);
    assign outputs[8096] = ~((layer0_outputs[9064]) | (layer0_outputs[4363]));
    assign outputs[8097] = layer0_outputs[6489];
    assign outputs[8098] = layer0_outputs[8136];
    assign outputs[8099] = ~(layer0_outputs[311]);
    assign outputs[8100] = ~((layer0_outputs[5898]) ^ (layer0_outputs[1889]));
    assign outputs[8101] = (layer0_outputs[5590]) & (layer0_outputs[5984]);
    assign outputs[8102] = layer0_outputs[9868];
    assign outputs[8103] = layer0_outputs[707];
    assign outputs[8104] = layer0_outputs[9233];
    assign outputs[8105] = ~((layer0_outputs[7399]) ^ (layer0_outputs[6608]));
    assign outputs[8106] = (layer0_outputs[9036]) ^ (layer0_outputs[4848]);
    assign outputs[8107] = (layer0_outputs[6931]) & (layer0_outputs[2611]);
    assign outputs[8108] = (layer0_outputs[7306]) & ~(layer0_outputs[9155]);
    assign outputs[8109] = (layer0_outputs[6926]) & ~(layer0_outputs[3891]);
    assign outputs[8110] = layer0_outputs[1145];
    assign outputs[8111] = ~(layer0_outputs[2150]);
    assign outputs[8112] = ~((layer0_outputs[4611]) ^ (layer0_outputs[9151]));
    assign outputs[8113] = ~((layer0_outputs[6668]) ^ (layer0_outputs[6006]));
    assign outputs[8114] = (layer0_outputs[1315]) & (layer0_outputs[390]);
    assign outputs[8115] = layer0_outputs[2763];
    assign outputs[8116] = (layer0_outputs[2806]) & (layer0_outputs[6390]);
    assign outputs[8117] = (layer0_outputs[8867]) ^ (layer0_outputs[9746]);
    assign outputs[8118] = ~(layer0_outputs[5668]);
    assign outputs[8119] = (layer0_outputs[6292]) & ~(layer0_outputs[938]);
    assign outputs[8120] = (layer0_outputs[6989]) ^ (layer0_outputs[2074]);
    assign outputs[8121] = ~(layer0_outputs[5227]);
    assign outputs[8122] = (layer0_outputs[3269]) & (layer0_outputs[4460]);
    assign outputs[8123] = layer0_outputs[7197];
    assign outputs[8124] = layer0_outputs[5198];
    assign outputs[8125] = ~(layer0_outputs[8145]);
    assign outputs[8126] = (layer0_outputs[9219]) ^ (layer0_outputs[3466]);
    assign outputs[8127] = (layer0_outputs[4658]) & ~(layer0_outputs[5008]);
    assign outputs[8128] = layer0_outputs[4348];
    assign outputs[8129] = ~((layer0_outputs[7345]) ^ (layer0_outputs[558]));
    assign outputs[8130] = ~((layer0_outputs[8765]) ^ (layer0_outputs[6397]));
    assign outputs[8131] = layer0_outputs[1070];
    assign outputs[8132] = (layer0_outputs[7963]) & ~(layer0_outputs[2178]);
    assign outputs[8133] = (layer0_outputs[7031]) & ~(layer0_outputs[1194]);
    assign outputs[8134] = ~(layer0_outputs[4520]);
    assign outputs[8135] = (layer0_outputs[4712]) | (layer0_outputs[310]);
    assign outputs[8136] = (layer0_outputs[265]) | (layer0_outputs[3229]);
    assign outputs[8137] = (layer0_outputs[8447]) & (layer0_outputs[1818]);
    assign outputs[8138] = ~((layer0_outputs[2019]) ^ (layer0_outputs[3530]));
    assign outputs[8139] = ~((layer0_outputs[10027]) ^ (layer0_outputs[3242]));
    assign outputs[8140] = (layer0_outputs[5578]) & ~(layer0_outputs[285]);
    assign outputs[8141] = (layer0_outputs[7794]) & ~(layer0_outputs[2130]);
    assign outputs[8142] = ~(layer0_outputs[67]);
    assign outputs[8143] = ~((layer0_outputs[4266]) | (layer0_outputs[5346]));
    assign outputs[8144] = ~(layer0_outputs[9959]);
    assign outputs[8145] = (layer0_outputs[560]) & ~(layer0_outputs[6901]);
    assign outputs[8146] = ~(layer0_outputs[4563]);
    assign outputs[8147] = (layer0_outputs[6718]) & (layer0_outputs[2475]);
    assign outputs[8148] = ~((layer0_outputs[5549]) ^ (layer0_outputs[6084]));
    assign outputs[8149] = (layer0_outputs[7130]) ^ (layer0_outputs[9100]);
    assign outputs[8150] = (layer0_outputs[6948]) & ~(layer0_outputs[8066]);
    assign outputs[8151] = layer0_outputs[1377];
    assign outputs[8152] = (layer0_outputs[9049]) ^ (layer0_outputs[6537]);
    assign outputs[8153] = (layer0_outputs[4691]) ^ (layer0_outputs[7147]);
    assign outputs[8154] = layer0_outputs[321];
    assign outputs[8155] = ~(layer0_outputs[9223]);
    assign outputs[8156] = layer0_outputs[1273];
    assign outputs[8157] = ~((layer0_outputs[1798]) | (layer0_outputs[9779]));
    assign outputs[8158] = layer0_outputs[6357];
    assign outputs[8159] = ~(layer0_outputs[4508]);
    assign outputs[8160] = ~((layer0_outputs[3310]) | (layer0_outputs[9138]));
    assign outputs[8161] = ~((layer0_outputs[2404]) ^ (layer0_outputs[9888]));
    assign outputs[8162] = layer0_outputs[453];
    assign outputs[8163] = (layer0_outputs[7833]) ^ (layer0_outputs[2511]);
    assign outputs[8164] = (layer0_outputs[5607]) & (layer0_outputs[6867]);
    assign outputs[8165] = ~(layer0_outputs[4420]);
    assign outputs[8166] = ~((layer0_outputs[1143]) ^ (layer0_outputs[4772]));
    assign outputs[8167] = (layer0_outputs[1578]) | (layer0_outputs[8797]);
    assign outputs[8168] = ~(layer0_outputs[4087]);
    assign outputs[8169] = layer0_outputs[5145];
    assign outputs[8170] = ~(layer0_outputs[361]);
    assign outputs[8171] = ~(layer0_outputs[7461]);
    assign outputs[8172] = layer0_outputs[6552];
    assign outputs[8173] = ~(layer0_outputs[8011]);
    assign outputs[8174] = layer0_outputs[4724];
    assign outputs[8175] = ~(layer0_outputs[2744]);
    assign outputs[8176] = layer0_outputs[2375];
    assign outputs[8177] = ~(layer0_outputs[255]);
    assign outputs[8178] = layer0_outputs[1657];
    assign outputs[8179] = ~(layer0_outputs[2776]);
    assign outputs[8180] = ~((layer0_outputs[352]) | (layer0_outputs[2168]));
    assign outputs[8181] = (layer0_outputs[1255]) & ~(layer0_outputs[6881]);
    assign outputs[8182] = layer0_outputs[4450];
    assign outputs[8183] = ~(layer0_outputs[2368]) | (layer0_outputs[7046]);
    assign outputs[8184] = (layer0_outputs[7804]) ^ (layer0_outputs[186]);
    assign outputs[8185] = ~(layer0_outputs[1144]);
    assign outputs[8186] = layer0_outputs[1963];
    assign outputs[8187] = (layer0_outputs[2141]) & ~(layer0_outputs[8009]);
    assign outputs[8188] = layer0_outputs[7894];
    assign outputs[8189] = layer0_outputs[9973];
    assign outputs[8190] = (layer0_outputs[4671]) & ~(layer0_outputs[7722]);
    assign outputs[8191] = ~(layer0_outputs[251]);
    assign outputs[8192] = ~(layer0_outputs[3946]) | (layer0_outputs[6927]);
    assign outputs[8193] = (layer0_outputs[4394]) | (layer0_outputs[6886]);
    assign outputs[8194] = (layer0_outputs[3810]) ^ (layer0_outputs[7913]);
    assign outputs[8195] = ~(layer0_outputs[9017]) | (layer0_outputs[4585]);
    assign outputs[8196] = ~((layer0_outputs[9237]) ^ (layer0_outputs[8167]));
    assign outputs[8197] = layer0_outputs[2651];
    assign outputs[8198] = layer0_outputs[10041];
    assign outputs[8199] = (layer0_outputs[3167]) ^ (layer0_outputs[3859]);
    assign outputs[8200] = (layer0_outputs[8931]) ^ (layer0_outputs[8045]);
    assign outputs[8201] = (layer0_outputs[3325]) ^ (layer0_outputs[6001]);
    assign outputs[8202] = layer0_outputs[8721];
    assign outputs[8203] = (layer0_outputs[1689]) & (layer0_outputs[8876]);
    assign outputs[8204] = layer0_outputs[7490];
    assign outputs[8205] = (layer0_outputs[348]) | (layer0_outputs[7304]);
    assign outputs[8206] = (layer0_outputs[5014]) ^ (layer0_outputs[6610]);
    assign outputs[8207] = ~(layer0_outputs[2680]);
    assign outputs[8208] = ~((layer0_outputs[486]) & (layer0_outputs[6497]));
    assign outputs[8209] = ~((layer0_outputs[10204]) & (layer0_outputs[8916]));
    assign outputs[8210] = ~(layer0_outputs[2731]);
    assign outputs[8211] = ~(layer0_outputs[4024]);
    assign outputs[8212] = layer0_outputs[5169];
    assign outputs[8213] = layer0_outputs[3533];
    assign outputs[8214] = (layer0_outputs[8207]) & ~(layer0_outputs[3555]);
    assign outputs[8215] = ~((layer0_outputs[8409]) ^ (layer0_outputs[8082]));
    assign outputs[8216] = (layer0_outputs[7669]) & (layer0_outputs[3427]);
    assign outputs[8217] = ~(layer0_outputs[6136]) | (layer0_outputs[2884]);
    assign outputs[8218] = layer0_outputs[2132];
    assign outputs[8219] = ~(layer0_outputs[2687]);
    assign outputs[8220] = layer0_outputs[3969];
    assign outputs[8221] = ~((layer0_outputs[7710]) | (layer0_outputs[4084]));
    assign outputs[8222] = ~(layer0_outputs[5272]);
    assign outputs[8223] = ~((layer0_outputs[2414]) | (layer0_outputs[8511]));
    assign outputs[8224] = ~(layer0_outputs[251]) | (layer0_outputs[900]);
    assign outputs[8225] = (layer0_outputs[222]) | (layer0_outputs[9623]);
    assign outputs[8226] = ~(layer0_outputs[1841]) | (layer0_outputs[1559]);
    assign outputs[8227] = ~((layer0_outputs[5847]) ^ (layer0_outputs[1992]));
    assign outputs[8228] = ~((layer0_outputs[10063]) & (layer0_outputs[9911]));
    assign outputs[8229] = layer0_outputs[1787];
    assign outputs[8230] = layer0_outputs[4552];
    assign outputs[8231] = ~(layer0_outputs[5154]);
    assign outputs[8232] = layer0_outputs[8677];
    assign outputs[8233] = (layer0_outputs[3793]) ^ (layer0_outputs[3870]);
    assign outputs[8234] = ~((layer0_outputs[8327]) ^ (layer0_outputs[4943]));
    assign outputs[8235] = ~(layer0_outputs[3835]);
    assign outputs[8236] = layer0_outputs[6979];
    assign outputs[8237] = ~(layer0_outputs[7418]) | (layer0_outputs[4045]);
    assign outputs[8238] = ~(layer0_outputs[9433]);
    assign outputs[8239] = (layer0_outputs[6306]) & (layer0_outputs[2553]);
    assign outputs[8240] = (layer0_outputs[3626]) & ~(layer0_outputs[9919]);
    assign outputs[8241] = ~((layer0_outputs[3929]) ^ (layer0_outputs[2825]));
    assign outputs[8242] = ~(layer0_outputs[727]);
    assign outputs[8243] = ~(layer0_outputs[5159]);
    assign outputs[8244] = (layer0_outputs[124]) & ~(layer0_outputs[912]);
    assign outputs[8245] = ~(layer0_outputs[1247]);
    assign outputs[8246] = layer0_outputs[7438];
    assign outputs[8247] = ~(layer0_outputs[5942]);
    assign outputs[8248] = ~((layer0_outputs[8003]) ^ (layer0_outputs[5913]));
    assign outputs[8249] = ~((layer0_outputs[7686]) & (layer0_outputs[7463]));
    assign outputs[8250] = layer0_outputs[8354];
    assign outputs[8251] = ~(layer0_outputs[4367]) | (layer0_outputs[7420]);
    assign outputs[8252] = ~(layer0_outputs[5842]);
    assign outputs[8253] = ~(layer0_outputs[4784]);
    assign outputs[8254] = ~(layer0_outputs[4183]) | (layer0_outputs[905]);
    assign outputs[8255] = ~((layer0_outputs[4825]) ^ (layer0_outputs[4340]));
    assign outputs[8256] = ~(layer0_outputs[2929]);
    assign outputs[8257] = ~(layer0_outputs[3379]) | (layer0_outputs[6009]);
    assign outputs[8258] = ~(layer0_outputs[3438]);
    assign outputs[8259] = ~(layer0_outputs[9867]);
    assign outputs[8260] = (layer0_outputs[5891]) ^ (layer0_outputs[8038]);
    assign outputs[8261] = ~((layer0_outputs[6677]) ^ (layer0_outputs[8101]));
    assign outputs[8262] = ~((layer0_outputs[8743]) ^ (layer0_outputs[8719]));
    assign outputs[8263] = layer0_outputs[3333];
    assign outputs[8264] = layer0_outputs[5062];
    assign outputs[8265] = layer0_outputs[299];
    assign outputs[8266] = ~(layer0_outputs[6275]);
    assign outputs[8267] = ~(layer0_outputs[7039]);
    assign outputs[8268] = ~((layer0_outputs[4878]) ^ (layer0_outputs[6352]));
    assign outputs[8269] = (layer0_outputs[4551]) ^ (layer0_outputs[3352]);
    assign outputs[8270] = ~(layer0_outputs[9669]) | (layer0_outputs[4252]);
    assign outputs[8271] = layer0_outputs[8602];
    assign outputs[8272] = (layer0_outputs[8594]) | (layer0_outputs[10031]);
    assign outputs[8273] = layer0_outputs[7229];
    assign outputs[8274] = (layer0_outputs[9794]) ^ (layer0_outputs[10091]);
    assign outputs[8275] = ~((layer0_outputs[8055]) ^ (layer0_outputs[1991]));
    assign outputs[8276] = (layer0_outputs[8052]) ^ (layer0_outputs[4787]);
    assign outputs[8277] = (layer0_outputs[5350]) ^ (layer0_outputs[1861]);
    assign outputs[8278] = layer0_outputs[4143];
    assign outputs[8279] = layer0_outputs[5879];
    assign outputs[8280] = (layer0_outputs[5133]) ^ (layer0_outputs[5504]);
    assign outputs[8281] = ~(layer0_outputs[6373]);
    assign outputs[8282] = layer0_outputs[496];
    assign outputs[8283] = ~((layer0_outputs[9294]) ^ (layer0_outputs[3095]));
    assign outputs[8284] = (layer0_outputs[7077]) ^ (layer0_outputs[7962]);
    assign outputs[8285] = ~(layer0_outputs[7179]);
    assign outputs[8286] = (layer0_outputs[5542]) ^ (layer0_outputs[3548]);
    assign outputs[8287] = (layer0_outputs[1871]) ^ (layer0_outputs[3017]);
    assign outputs[8288] = ~(layer0_outputs[5999]) | (layer0_outputs[7695]);
    assign outputs[8289] = layer0_outputs[5733];
    assign outputs[8290] = (layer0_outputs[3200]) | (layer0_outputs[5468]);
    assign outputs[8291] = ~(layer0_outputs[3925]);
    assign outputs[8292] = ~(layer0_outputs[412]);
    assign outputs[8293] = (layer0_outputs[7118]) ^ (layer0_outputs[8774]);
    assign outputs[8294] = ~((layer0_outputs[9761]) | (layer0_outputs[8198]));
    assign outputs[8295] = ~(layer0_outputs[3905]);
    assign outputs[8296] = ~(layer0_outputs[8238]);
    assign outputs[8297] = ~(layer0_outputs[6114]);
    assign outputs[8298] = ~((layer0_outputs[9744]) & (layer0_outputs[2973]));
    assign outputs[8299] = layer0_outputs[1243];
    assign outputs[8300] = layer0_outputs[2191];
    assign outputs[8301] = layer0_outputs[1202];
    assign outputs[8302] = ~(layer0_outputs[7989]) | (layer0_outputs[36]);
    assign outputs[8303] = layer0_outputs[6500];
    assign outputs[8304] = ~(layer0_outputs[8180]);
    assign outputs[8305] = ~(layer0_outputs[2894]);
    assign outputs[8306] = (layer0_outputs[4084]) ^ (layer0_outputs[8383]);
    assign outputs[8307] = ~((layer0_outputs[2100]) | (layer0_outputs[528]));
    assign outputs[8308] = ~((layer0_outputs[631]) | (layer0_outputs[983]));
    assign outputs[8309] = ~(layer0_outputs[4336]);
    assign outputs[8310] = (layer0_outputs[9690]) ^ (layer0_outputs[3747]);
    assign outputs[8311] = ~(layer0_outputs[5303]) | (layer0_outputs[4811]);
    assign outputs[8312] = (layer0_outputs[1823]) ^ (layer0_outputs[10030]);
    assign outputs[8313] = ~((layer0_outputs[5893]) & (layer0_outputs[6579]));
    assign outputs[8314] = layer0_outputs[6829];
    assign outputs[8315] = (layer0_outputs[8279]) & ~(layer0_outputs[6722]);
    assign outputs[8316] = ~(layer0_outputs[6645]) | (layer0_outputs[7341]);
    assign outputs[8317] = ~((layer0_outputs[1599]) & (layer0_outputs[2688]));
    assign outputs[8318] = (layer0_outputs[7135]) ^ (layer0_outputs[7541]);
    assign outputs[8319] = layer0_outputs[1654];
    assign outputs[8320] = layer0_outputs[2309];
    assign outputs[8321] = ~((layer0_outputs[10193]) ^ (layer0_outputs[3466]));
    assign outputs[8322] = ~(layer0_outputs[9221]);
    assign outputs[8323] = layer0_outputs[3701];
    assign outputs[8324] = layer0_outputs[7766];
    assign outputs[8325] = layer0_outputs[7593];
    assign outputs[8326] = ~(layer0_outputs[7433]) | (layer0_outputs[3240]);
    assign outputs[8327] = ~(layer0_outputs[2935]);
    assign outputs[8328] = ~(layer0_outputs[6924]);
    assign outputs[8329] = layer0_outputs[4991];
    assign outputs[8330] = ~((layer0_outputs[2224]) & (layer0_outputs[9657]));
    assign outputs[8331] = (layer0_outputs[2376]) & (layer0_outputs[1257]);
    assign outputs[8332] = ~(layer0_outputs[7301]) | (layer0_outputs[9693]);
    assign outputs[8333] = ~(layer0_outputs[7871]);
    assign outputs[8334] = ~((layer0_outputs[7338]) ^ (layer0_outputs[2556]));
    assign outputs[8335] = (layer0_outputs[8648]) & ~(layer0_outputs[659]);
    assign outputs[8336] = layer0_outputs[4674];
    assign outputs[8337] = ~((layer0_outputs[4116]) ^ (layer0_outputs[3405]));
    assign outputs[8338] = (layer0_outputs[6449]) ^ (layer0_outputs[4672]);
    assign outputs[8339] = (layer0_outputs[9455]) ^ (layer0_outputs[9456]);
    assign outputs[8340] = ~(layer0_outputs[1208]) | (layer0_outputs[4964]);
    assign outputs[8341] = layer0_outputs[4048];
    assign outputs[8342] = ~(layer0_outputs[8109]) | (layer0_outputs[8990]);
    assign outputs[8343] = ~(layer0_outputs[2045]);
    assign outputs[8344] = layer0_outputs[2198];
    assign outputs[8345] = ~((layer0_outputs[5770]) ^ (layer0_outputs[296]));
    assign outputs[8346] = ~(layer0_outputs[5051]);
    assign outputs[8347] = ~(layer0_outputs[4574]) | (layer0_outputs[792]);
    assign outputs[8348] = ~(layer0_outputs[2211]);
    assign outputs[8349] = ~((layer0_outputs[7867]) ^ (layer0_outputs[763]));
    assign outputs[8350] = ~((layer0_outputs[6781]) ^ (layer0_outputs[327]));
    assign outputs[8351] = layer0_outputs[6071];
    assign outputs[8352] = (layer0_outputs[2925]) | (layer0_outputs[654]);
    assign outputs[8353] = layer0_outputs[3512];
    assign outputs[8354] = (layer0_outputs[10127]) | (layer0_outputs[7620]);
    assign outputs[8355] = layer0_outputs[525];
    assign outputs[8356] = ~((layer0_outputs[749]) ^ (layer0_outputs[4973]));
    assign outputs[8357] = ~(layer0_outputs[6302]);
    assign outputs[8358] = ~(layer0_outputs[1002]);
    assign outputs[8359] = (layer0_outputs[5915]) ^ (layer0_outputs[1260]);
    assign outputs[8360] = layer0_outputs[8796];
    assign outputs[8361] = ~(layer0_outputs[10135]);
    assign outputs[8362] = ~((layer0_outputs[9699]) & (layer0_outputs[8983]));
    assign outputs[8363] = ~(layer0_outputs[298]) | (layer0_outputs[9826]);
    assign outputs[8364] = ~(layer0_outputs[643]);
    assign outputs[8365] = ~(layer0_outputs[1915]);
    assign outputs[8366] = (layer0_outputs[9444]) ^ (layer0_outputs[9452]);
    assign outputs[8367] = (layer0_outputs[1049]) | (layer0_outputs[2988]);
    assign outputs[8368] = ~((layer0_outputs[7297]) & (layer0_outputs[2147]));
    assign outputs[8369] = ~((layer0_outputs[1982]) ^ (layer0_outputs[3066]));
    assign outputs[8370] = ~(layer0_outputs[5877]) | (layer0_outputs[334]);
    assign outputs[8371] = layer0_outputs[8099];
    assign outputs[8372] = ~(layer0_outputs[5105]);
    assign outputs[8373] = layer0_outputs[4640];
    assign outputs[8374] = ~((layer0_outputs[2641]) ^ (layer0_outputs[1946]));
    assign outputs[8375] = (layer0_outputs[4621]) ^ (layer0_outputs[6774]);
    assign outputs[8376] = ~(layer0_outputs[4651]) | (layer0_outputs[10025]);
    assign outputs[8377] = layer0_outputs[9659];
    assign outputs[8378] = ~(layer0_outputs[4100]);
    assign outputs[8379] = ~(layer0_outputs[8841]) | (layer0_outputs[4008]);
    assign outputs[8380] = ~(layer0_outputs[4091]);
    assign outputs[8381] = ~((layer0_outputs[6523]) ^ (layer0_outputs[9938]));
    assign outputs[8382] = layer0_outputs[6177];
    assign outputs[8383] = ~((layer0_outputs[4471]) ^ (layer0_outputs[1284]));
    assign outputs[8384] = ~(layer0_outputs[2815]);
    assign outputs[8385] = (layer0_outputs[2712]) ^ (layer0_outputs[7137]);
    assign outputs[8386] = (layer0_outputs[9343]) ^ (layer0_outputs[2472]);
    assign outputs[8387] = 1'b1;
    assign outputs[8388] = (layer0_outputs[1024]) ^ (layer0_outputs[7013]);
    assign outputs[8389] = (layer0_outputs[10114]) | (layer0_outputs[2433]);
    assign outputs[8390] = (layer0_outputs[2095]) ^ (layer0_outputs[2528]);
    assign outputs[8391] = ~(layer0_outputs[9457]) | (layer0_outputs[7310]);
    assign outputs[8392] = ~(layer0_outputs[645]);
    assign outputs[8393] = ~(layer0_outputs[1949]) | (layer0_outputs[8590]);
    assign outputs[8394] = ~((layer0_outputs[6494]) ^ (layer0_outputs[7692]));
    assign outputs[8395] = 1'b1;
    assign outputs[8396] = ~(layer0_outputs[9372]);
    assign outputs[8397] = ~((layer0_outputs[1630]) ^ (layer0_outputs[849]));
    assign outputs[8398] = ~((layer0_outputs[8817]) ^ (layer0_outputs[6813]));
    assign outputs[8399] = ~(layer0_outputs[4284]);
    assign outputs[8400] = ~((layer0_outputs[3868]) | (layer0_outputs[8282]));
    assign outputs[8401] = ~(layer0_outputs[9583]);
    assign outputs[8402] = ~((layer0_outputs[2320]) ^ (layer0_outputs[927]));
    assign outputs[8403] = ~((layer0_outputs[3021]) ^ (layer0_outputs[7910]));
    assign outputs[8404] = layer0_outputs[4230];
    assign outputs[8405] = ~(layer0_outputs[5498]);
    assign outputs[8406] = ~(layer0_outputs[955]);
    assign outputs[8407] = ~((layer0_outputs[9769]) ^ (layer0_outputs[3675]));
    assign outputs[8408] = layer0_outputs[5422];
    assign outputs[8409] = (layer0_outputs[8083]) & ~(layer0_outputs[6459]);
    assign outputs[8410] = ~(layer0_outputs[7535]) | (layer0_outputs[1624]);
    assign outputs[8411] = ~((layer0_outputs[6171]) ^ (layer0_outputs[4042]));
    assign outputs[8412] = ~(layer0_outputs[5906]) | (layer0_outputs[4153]);
    assign outputs[8413] = (layer0_outputs[9454]) & ~(layer0_outputs[5445]);
    assign outputs[8414] = ~(layer0_outputs[8359]);
    assign outputs[8415] = ~(layer0_outputs[4849]) | (layer0_outputs[2490]);
    assign outputs[8416] = ~(layer0_outputs[148]);
    assign outputs[8417] = ~(layer0_outputs[2286]) | (layer0_outputs[1314]);
    assign outputs[8418] = ~(layer0_outputs[1900]);
    assign outputs[8419] = ~(layer0_outputs[7613]);
    assign outputs[8420] = (layer0_outputs[6630]) ^ (layer0_outputs[7685]);
    assign outputs[8421] = layer0_outputs[3614];
    assign outputs[8422] = layer0_outputs[4528];
    assign outputs[8423] = ~(layer0_outputs[7403]) | (layer0_outputs[6206]);
    assign outputs[8424] = ~((layer0_outputs[3591]) ^ (layer0_outputs[5824]));
    assign outputs[8425] = ~((layer0_outputs[2969]) | (layer0_outputs[6705]));
    assign outputs[8426] = (layer0_outputs[4862]) & ~(layer0_outputs[10227]);
    assign outputs[8427] = ~(layer0_outputs[945]) | (layer0_outputs[1172]);
    assign outputs[8428] = ~(layer0_outputs[5260]) | (layer0_outputs[9941]);
    assign outputs[8429] = layer0_outputs[5348];
    assign outputs[8430] = layer0_outputs[6118];
    assign outputs[8431] = layer0_outputs[5788];
    assign outputs[8432] = (layer0_outputs[404]) & ~(layer0_outputs[9417]);
    assign outputs[8433] = (layer0_outputs[7123]) | (layer0_outputs[9873]);
    assign outputs[8434] = (layer0_outputs[2110]) | (layer0_outputs[6255]);
    assign outputs[8435] = ~((layer0_outputs[9003]) ^ (layer0_outputs[2735]));
    assign outputs[8436] = (layer0_outputs[31]) ^ (layer0_outputs[2128]);
    assign outputs[8437] = ~((layer0_outputs[6035]) ^ (layer0_outputs[2482]));
    assign outputs[8438] = ~(layer0_outputs[166]);
    assign outputs[8439] = ~((layer0_outputs[9382]) & (layer0_outputs[9394]));
    assign outputs[8440] = ~((layer0_outputs[4323]) ^ (layer0_outputs[2031]));
    assign outputs[8441] = (layer0_outputs[9030]) & ~(layer0_outputs[7040]);
    assign outputs[8442] = (layer0_outputs[9651]) & ~(layer0_outputs[4934]);
    assign outputs[8443] = ~(layer0_outputs[4227]);
    assign outputs[8444] = layer0_outputs[10161];
    assign outputs[8445] = ~(layer0_outputs[7528]);
    assign outputs[8446] = ~((layer0_outputs[7911]) ^ (layer0_outputs[6822]));
    assign outputs[8447] = layer0_outputs[3273];
    assign outputs[8448] = ~((layer0_outputs[2576]) & (layer0_outputs[8433]));
    assign outputs[8449] = ~((layer0_outputs[4220]) ^ (layer0_outputs[9265]));
    assign outputs[8450] = ~(layer0_outputs[8342]);
    assign outputs[8451] = layer0_outputs[8064];
    assign outputs[8452] = (layer0_outputs[6132]) & ~(layer0_outputs[7796]);
    assign outputs[8453] = (layer0_outputs[7244]) & (layer0_outputs[8571]);
    assign outputs[8454] = (layer0_outputs[3188]) ^ (layer0_outputs[599]);
    assign outputs[8455] = ~(layer0_outputs[3106]) | (layer0_outputs[9179]);
    assign outputs[8456] = ~((layer0_outputs[4863]) ^ (layer0_outputs[7252]));
    assign outputs[8457] = ~((layer0_outputs[1282]) ^ (layer0_outputs[6276]));
    assign outputs[8458] = (layer0_outputs[5185]) & ~(layer0_outputs[5175]);
    assign outputs[8459] = ~(layer0_outputs[10175]) | (layer0_outputs[9565]);
    assign outputs[8460] = ~((layer0_outputs[5187]) ^ (layer0_outputs[8744]));
    assign outputs[8461] = (layer0_outputs[8209]) ^ (layer0_outputs[8183]);
    assign outputs[8462] = ~(layer0_outputs[6192]) | (layer0_outputs[2926]);
    assign outputs[8463] = (layer0_outputs[7218]) | (layer0_outputs[3827]);
    assign outputs[8464] = ~(layer0_outputs[5338]);
    assign outputs[8465] = ~((layer0_outputs[271]) ^ (layer0_outputs[8076]));
    assign outputs[8466] = layer0_outputs[8583];
    assign outputs[8467] = ~((layer0_outputs[1731]) ^ (layer0_outputs[3337]));
    assign outputs[8468] = (layer0_outputs[10239]) ^ (layer0_outputs[8013]);
    assign outputs[8469] = layer0_outputs[245];
    assign outputs[8470] = (layer0_outputs[1929]) & ~(layer0_outputs[2145]);
    assign outputs[8471] = ~(layer0_outputs[1161]);
    assign outputs[8472] = ~(layer0_outputs[7573]);
    assign outputs[8473] = ~(layer0_outputs[5705]);
    assign outputs[8474] = ~(layer0_outputs[9924]) | (layer0_outputs[867]);
    assign outputs[8475] = ~(layer0_outputs[4000]);
    assign outputs[8476] = (layer0_outputs[7801]) ^ (layer0_outputs[8966]);
    assign outputs[8477] = ~(layer0_outputs[767]);
    assign outputs[8478] = layer0_outputs[6325];
    assign outputs[8479] = ~(layer0_outputs[9060]);
    assign outputs[8480] = (layer0_outputs[3763]) ^ (layer0_outputs[5774]);
    assign outputs[8481] = layer0_outputs[9814];
    assign outputs[8482] = ~(layer0_outputs[2079]);
    assign outputs[8483] = ~(layer0_outputs[1021]) | (layer0_outputs[3343]);
    assign outputs[8484] = (layer0_outputs[2237]) & ~(layer0_outputs[8513]);
    assign outputs[8485] = ~(layer0_outputs[1232]);
    assign outputs[8486] = (layer0_outputs[6207]) | (layer0_outputs[2746]);
    assign outputs[8487] = layer0_outputs[3328];
    assign outputs[8488] = ~(layer0_outputs[518]);
    assign outputs[8489] = (layer0_outputs[6600]) | (layer0_outputs[9891]);
    assign outputs[8490] = layer0_outputs[9203];
    assign outputs[8491] = ~((layer0_outputs[4537]) & (layer0_outputs[7018]));
    assign outputs[8492] = ~((layer0_outputs[10233]) ^ (layer0_outputs[4910]));
    assign outputs[8493] = (layer0_outputs[561]) ^ (layer0_outputs[8893]);
    assign outputs[8494] = (layer0_outputs[2689]) & ~(layer0_outputs[5216]);
    assign outputs[8495] = layer0_outputs[1628];
    assign outputs[8496] = ~(layer0_outputs[3351]) | (layer0_outputs[9252]);
    assign outputs[8497] = ~(layer0_outputs[1499]);
    assign outputs[8498] = (layer0_outputs[258]) ^ (layer0_outputs[6346]);
    assign outputs[8499] = layer0_outputs[5975];
    assign outputs[8500] = ~(layer0_outputs[1726]);
    assign outputs[8501] = ~(layer0_outputs[4489]);
    assign outputs[8502] = layer0_outputs[2455];
    assign outputs[8503] = ~((layer0_outputs[1971]) ^ (layer0_outputs[1644]));
    assign outputs[8504] = (layer0_outputs[8010]) ^ (layer0_outputs[2526]);
    assign outputs[8505] = ~(layer0_outputs[8194]);
    assign outputs[8506] = layer0_outputs[2932];
    assign outputs[8507] = layer0_outputs[6364];
    assign outputs[8508] = ~(layer0_outputs[9599]);
    assign outputs[8509] = ~((layer0_outputs[3794]) ^ (layer0_outputs[9668]));
    assign outputs[8510] = ~(layer0_outputs[9626]);
    assign outputs[8511] = ~(layer0_outputs[8331]) | (layer0_outputs[4451]);
    assign outputs[8512] = (layer0_outputs[7823]) & ~(layer0_outputs[1346]);
    assign outputs[8513] = layer0_outputs[2593];
    assign outputs[8514] = (layer0_outputs[410]) ^ (layer0_outputs[660]);
    assign outputs[8515] = (layer0_outputs[5168]) | (layer0_outputs[4452]);
    assign outputs[8516] = ~(layer0_outputs[8405]);
    assign outputs[8517] = (layer0_outputs[7143]) & ~(layer0_outputs[8982]);
    assign outputs[8518] = ~(layer0_outputs[7322]) | (layer0_outputs[4233]);
    assign outputs[8519] = ~((layer0_outputs[8715]) ^ (layer0_outputs[577]));
    assign outputs[8520] = (layer0_outputs[4035]) ^ (layer0_outputs[3703]);
    assign outputs[8521] = ~((layer0_outputs[7562]) & (layer0_outputs[4515]));
    assign outputs[8522] = layer0_outputs[4984];
    assign outputs[8523] = (layer0_outputs[9951]) ^ (layer0_outputs[9268]);
    assign outputs[8524] = ~(layer0_outputs[2170]);
    assign outputs[8525] = ~((layer0_outputs[4792]) ^ (layer0_outputs[5108]));
    assign outputs[8526] = layer0_outputs[9683];
    assign outputs[8527] = layer0_outputs[7369];
    assign outputs[8528] = (layer0_outputs[9573]) ^ (layer0_outputs[1555]);
    assign outputs[8529] = (layer0_outputs[1111]) ^ (layer0_outputs[5502]);
    assign outputs[8530] = (layer0_outputs[9594]) & ~(layer0_outputs[135]);
    assign outputs[8531] = (layer0_outputs[20]) & (layer0_outputs[8013]);
    assign outputs[8532] = ~(layer0_outputs[4253]);
    assign outputs[8533] = (layer0_outputs[3633]) & ~(layer0_outputs[770]);
    assign outputs[8534] = ~(layer0_outputs[2784]) | (layer0_outputs[5950]);
    assign outputs[8535] = layer0_outputs[849];
    assign outputs[8536] = ~(layer0_outputs[1002]);
    assign outputs[8537] = (layer0_outputs[8454]) ^ (layer0_outputs[9063]);
    assign outputs[8538] = ~(layer0_outputs[6033]);
    assign outputs[8539] = layer0_outputs[1228];
    assign outputs[8540] = ~(layer0_outputs[7047]);
    assign outputs[8541] = (layer0_outputs[5756]) & ~(layer0_outputs[1593]);
    assign outputs[8542] = ~((layer0_outputs[5806]) & (layer0_outputs[9011]));
    assign outputs[8543] = layer0_outputs[4324];
    assign outputs[8544] = (layer0_outputs[7785]) ^ (layer0_outputs[5126]);
    assign outputs[8545] = (layer0_outputs[3967]) | (layer0_outputs[2651]);
    assign outputs[8546] = layer0_outputs[6966];
    assign outputs[8547] = ~(layer0_outputs[2009]);
    assign outputs[8548] = ~((layer0_outputs[6367]) ^ (layer0_outputs[1745]));
    assign outputs[8549] = ~((layer0_outputs[1510]) ^ (layer0_outputs[376]));
    assign outputs[8550] = ~(layer0_outputs[7088]);
    assign outputs[8551] = ~((layer0_outputs[876]) & (layer0_outputs[9102]));
    assign outputs[8552] = (layer0_outputs[4266]) | (layer0_outputs[3032]);
    assign outputs[8553] = ~((layer0_outputs[2062]) & (layer0_outputs[6348]));
    assign outputs[8554] = ~(layer0_outputs[3591]);
    assign outputs[8555] = (layer0_outputs[1893]) ^ (layer0_outputs[1697]);
    assign outputs[8556] = layer0_outputs[4682];
    assign outputs[8557] = ~(layer0_outputs[1150]);
    assign outputs[8558] = ~(layer0_outputs[1124]);
    assign outputs[8559] = ~(layer0_outputs[706]) | (layer0_outputs[3533]);
    assign outputs[8560] = layer0_outputs[5282];
    assign outputs[8561] = layer0_outputs[9281];
    assign outputs[8562] = ~((layer0_outputs[3112]) ^ (layer0_outputs[4403]));
    assign outputs[8563] = (layer0_outputs[5565]) & ~(layer0_outputs[3292]);
    assign outputs[8564] = ~((layer0_outputs[8349]) | (layer0_outputs[7954]));
    assign outputs[8565] = (layer0_outputs[2602]) | (layer0_outputs[9077]);
    assign outputs[8566] = (layer0_outputs[3945]) ^ (layer0_outputs[3460]);
    assign outputs[8567] = layer0_outputs[2354];
    assign outputs[8568] = (layer0_outputs[5727]) | (layer0_outputs[9807]);
    assign outputs[8569] = (layer0_outputs[9009]) ^ (layer0_outputs[7785]);
    assign outputs[8570] = layer0_outputs[10099];
    assign outputs[8571] = layer0_outputs[8520];
    assign outputs[8572] = (layer0_outputs[3381]) | (layer0_outputs[948]);
    assign outputs[8573] = ~(layer0_outputs[955]);
    assign outputs[8574] = ~((layer0_outputs[2253]) ^ (layer0_outputs[5742]));
    assign outputs[8575] = layer0_outputs[8459];
    assign outputs[8576] = (layer0_outputs[6709]) ^ (layer0_outputs[7274]);
    assign outputs[8577] = ~((layer0_outputs[9167]) & (layer0_outputs[2569]));
    assign outputs[8578] = (layer0_outputs[4701]) ^ (layer0_outputs[916]);
    assign outputs[8579] = layer0_outputs[2227];
    assign outputs[8580] = (layer0_outputs[3071]) | (layer0_outputs[2665]);
    assign outputs[8581] = (layer0_outputs[3152]) ^ (layer0_outputs[7281]);
    assign outputs[8582] = layer0_outputs[7000];
    assign outputs[8583] = ~(layer0_outputs[4191]);
    assign outputs[8584] = ~((layer0_outputs[10227]) ^ (layer0_outputs[8585]));
    assign outputs[8585] = (layer0_outputs[1652]) ^ (layer0_outputs[4620]);
    assign outputs[8586] = layer0_outputs[1856];
    assign outputs[8587] = ~(layer0_outputs[7583]);
    assign outputs[8588] = layer0_outputs[3357];
    assign outputs[8589] = ~((layer0_outputs[1551]) ^ (layer0_outputs[2764]));
    assign outputs[8590] = ~(layer0_outputs[8790]) | (layer0_outputs[4913]);
    assign outputs[8591] = (layer0_outputs[6825]) ^ (layer0_outputs[2554]);
    assign outputs[8592] = ~((layer0_outputs[2668]) & (layer0_outputs[6183]));
    assign outputs[8593] = ~(layer0_outputs[416]) | (layer0_outputs[8746]);
    assign outputs[8594] = ~(layer0_outputs[8907]);
    assign outputs[8595] = layer0_outputs[562];
    assign outputs[8596] = ~(layer0_outputs[5965]) | (layer0_outputs[8420]);
    assign outputs[8597] = ~(layer0_outputs[6265]);
    assign outputs[8598] = ~((layer0_outputs[8595]) & (layer0_outputs[3726]));
    assign outputs[8599] = ~(layer0_outputs[1079]) | (layer0_outputs[6920]);
    assign outputs[8600] = ~((layer0_outputs[4486]) & (layer0_outputs[9887]));
    assign outputs[8601] = (layer0_outputs[772]) ^ (layer0_outputs[578]);
    assign outputs[8602] = (layer0_outputs[5799]) | (layer0_outputs[5789]);
    assign outputs[8603] = ~(layer0_outputs[5248]) | (layer0_outputs[1945]);
    assign outputs[8604] = ~((layer0_outputs[6828]) ^ (layer0_outputs[5286]));
    assign outputs[8605] = (layer0_outputs[4647]) & ~(layer0_outputs[3162]);
    assign outputs[8606] = ~((layer0_outputs[8719]) ^ (layer0_outputs[2830]));
    assign outputs[8607] = ~(layer0_outputs[5576]);
    assign outputs[8608] = ~(layer0_outputs[6615]) | (layer0_outputs[4932]);
    assign outputs[8609] = (layer0_outputs[1785]) ^ (layer0_outputs[6631]);
    assign outputs[8610] = ~((layer0_outputs[2769]) | (layer0_outputs[5845]));
    assign outputs[8611] = ~(layer0_outputs[4132]) | (layer0_outputs[3395]);
    assign outputs[8612] = (layer0_outputs[7986]) | (layer0_outputs[4268]);
    assign outputs[8613] = ~(layer0_outputs[4851]) | (layer0_outputs[5917]);
    assign outputs[8614] = ~((layer0_outputs[8397]) ^ (layer0_outputs[1026]));
    assign outputs[8615] = ~(layer0_outputs[2771]);
    assign outputs[8616] = ~(layer0_outputs[4740]);
    assign outputs[8617] = (layer0_outputs[6999]) ^ (layer0_outputs[2883]);
    assign outputs[8618] = ~(layer0_outputs[5390]) | (layer0_outputs[3531]);
    assign outputs[8619] = (layer0_outputs[7012]) ^ (layer0_outputs[5655]);
    assign outputs[8620] = ~(layer0_outputs[6873]);
    assign outputs[8621] = layer0_outputs[9972];
    assign outputs[8622] = (layer0_outputs[2384]) ^ (layer0_outputs[8523]);
    assign outputs[8623] = (layer0_outputs[8319]) ^ (layer0_outputs[9060]);
    assign outputs[8624] = layer0_outputs[4756];
    assign outputs[8625] = ~(layer0_outputs[827]);
    assign outputs[8626] = ~((layer0_outputs[9874]) ^ (layer0_outputs[7542]));
    assign outputs[8627] = ~(layer0_outputs[8371]) | (layer0_outputs[6511]);
    assign outputs[8628] = layer0_outputs[4727];
    assign outputs[8629] = ~(layer0_outputs[6869]) | (layer0_outputs[2961]);
    assign outputs[8630] = (layer0_outputs[10209]) ^ (layer0_outputs[9391]);
    assign outputs[8631] = ~(layer0_outputs[2018]) | (layer0_outputs[9678]);
    assign outputs[8632] = (layer0_outputs[4982]) ^ (layer0_outputs[5940]);
    assign outputs[8633] = ~((layer0_outputs[1472]) ^ (layer0_outputs[6484]));
    assign outputs[8634] = ~((layer0_outputs[1885]) & (layer0_outputs[4346]));
    assign outputs[8635] = ~(layer0_outputs[4331]);
    assign outputs[8636] = ~(layer0_outputs[9687]) | (layer0_outputs[7002]);
    assign outputs[8637] = ~((layer0_outputs[8614]) ^ (layer0_outputs[3]));
    assign outputs[8638] = layer0_outputs[399];
    assign outputs[8639] = (layer0_outputs[1524]) & (layer0_outputs[9512]);
    assign outputs[8640] = ~(layer0_outputs[341]);
    assign outputs[8641] = ~((layer0_outputs[4550]) ^ (layer0_outputs[4273]));
    assign outputs[8642] = layer0_outputs[3951];
    assign outputs[8643] = (layer0_outputs[7236]) ^ (layer0_outputs[8480]);
    assign outputs[8644] = ~((layer0_outputs[9231]) ^ (layer0_outputs[5739]));
    assign outputs[8645] = ~((layer0_outputs[10017]) | (layer0_outputs[7502]));
    assign outputs[8646] = (layer0_outputs[3700]) & ~(layer0_outputs[9772]);
    assign outputs[8647] = ~(layer0_outputs[3618]);
    assign outputs[8648] = ~(layer0_outputs[454]) | (layer0_outputs[6183]);
    assign outputs[8649] = layer0_outputs[1849];
    assign outputs[8650] = ~(layer0_outputs[7665]);
    assign outputs[8651] = ~(layer0_outputs[4286]);
    assign outputs[8652] = ~(layer0_outputs[3564]);
    assign outputs[8653] = ~(layer0_outputs[173]);
    assign outputs[8654] = ~(layer0_outputs[5995]) | (layer0_outputs[4693]);
    assign outputs[8655] = ~(layer0_outputs[3005]);
    assign outputs[8656] = ~(layer0_outputs[6873]);
    assign outputs[8657] = (layer0_outputs[4435]) ^ (layer0_outputs[5106]);
    assign outputs[8658] = (layer0_outputs[8298]) ^ (layer0_outputs[2556]);
    assign outputs[8659] = layer0_outputs[4827];
    assign outputs[8660] = ~(layer0_outputs[6240]);
    assign outputs[8661] = (layer0_outputs[680]) ^ (layer0_outputs[3865]);
    assign outputs[8662] = ~((layer0_outputs[9234]) & (layer0_outputs[7831]));
    assign outputs[8663] = layer0_outputs[9834];
    assign outputs[8664] = ~(layer0_outputs[10070]);
    assign outputs[8665] = ~(layer0_outputs[2158]);
    assign outputs[8666] = ~((layer0_outputs[6294]) & (layer0_outputs[6336]));
    assign outputs[8667] = (layer0_outputs[4750]) ^ (layer0_outputs[1911]);
    assign outputs[8668] = ~((layer0_outputs[8342]) ^ (layer0_outputs[5084]));
    assign outputs[8669] = layer0_outputs[2269];
    assign outputs[8670] = ~(layer0_outputs[8424]);
    assign outputs[8671] = ~((layer0_outputs[1526]) ^ (layer0_outputs[2304]));
    assign outputs[8672] = layer0_outputs[9738];
    assign outputs[8673] = ~((layer0_outputs[4136]) & (layer0_outputs[8222]));
    assign outputs[8674] = ~(layer0_outputs[3432]) | (layer0_outputs[4523]);
    assign outputs[8675] = ~(layer0_outputs[1678]) | (layer0_outputs[5141]);
    assign outputs[8676] = (layer0_outputs[3627]) & ~(layer0_outputs[9902]);
    assign outputs[8677] = (layer0_outputs[10112]) & (layer0_outputs[6487]);
    assign outputs[8678] = ~(layer0_outputs[5112]);
    assign outputs[8679] = ~((layer0_outputs[1519]) ^ (layer0_outputs[3202]));
    assign outputs[8680] = ~(layer0_outputs[7724]) | (layer0_outputs[1686]);
    assign outputs[8681] = layer0_outputs[1465];
    assign outputs[8682] = ~(layer0_outputs[8666]);
    assign outputs[8683] = ~((layer0_outputs[3439]) | (layer0_outputs[9406]));
    assign outputs[8684] = ~((layer0_outputs[1080]) ^ (layer0_outputs[2473]));
    assign outputs[8685] = layer0_outputs[7051];
    assign outputs[8686] = layer0_outputs[5132];
    assign outputs[8687] = ~(layer0_outputs[2064]);
    assign outputs[8688] = ~(layer0_outputs[2315]);
    assign outputs[8689] = ~(layer0_outputs[3237]);
    assign outputs[8690] = ~((layer0_outputs[3621]) ^ (layer0_outputs[7957]));
    assign outputs[8691] = ~((layer0_outputs[9145]) & (layer0_outputs[4426]));
    assign outputs[8692] = ~((layer0_outputs[2676]) ^ (layer0_outputs[6500]));
    assign outputs[8693] = ~(layer0_outputs[7557]) | (layer0_outputs[9479]);
    assign outputs[8694] = ~((layer0_outputs[8988]) & (layer0_outputs[3232]));
    assign outputs[8695] = ~((layer0_outputs[10003]) ^ (layer0_outputs[1817]));
    assign outputs[8696] = ~(layer0_outputs[749]);
    assign outputs[8697] = (layer0_outputs[10005]) ^ (layer0_outputs[10107]);
    assign outputs[8698] = layer0_outputs[1640];
    assign outputs[8699] = (layer0_outputs[8231]) ^ (layer0_outputs[2201]);
    assign outputs[8700] = ~(layer0_outputs[4425]);
    assign outputs[8701] = ~((layer0_outputs[93]) ^ (layer0_outputs[2809]));
    assign outputs[8702] = ~((layer0_outputs[9048]) ^ (layer0_outputs[2609]));
    assign outputs[8703] = layer0_outputs[7919];
    assign outputs[8704] = ~(layer0_outputs[3801]) | (layer0_outputs[8459]);
    assign outputs[8705] = ~(layer0_outputs[798]) | (layer0_outputs[324]);
    assign outputs[8706] = ~(layer0_outputs[1457]);
    assign outputs[8707] = layer0_outputs[8079];
    assign outputs[8708] = layer0_outputs[8780];
    assign outputs[8709] = layer0_outputs[6225];
    assign outputs[8710] = layer0_outputs[4664];
    assign outputs[8711] = (layer0_outputs[4209]) & (layer0_outputs[8380]);
    assign outputs[8712] = (layer0_outputs[4686]) | (layer0_outputs[3425]);
    assign outputs[8713] = ~((layer0_outputs[7865]) ^ (layer0_outputs[2431]));
    assign outputs[8714] = ~(layer0_outputs[2176]);
    assign outputs[8715] = ~(layer0_outputs[7659]) | (layer0_outputs[9846]);
    assign outputs[8716] = ~(layer0_outputs[5689]);
    assign outputs[8717] = ~(layer0_outputs[1478]);
    assign outputs[8718] = ~((layer0_outputs[3385]) ^ (layer0_outputs[6642]));
    assign outputs[8719] = (layer0_outputs[10166]) ^ (layer0_outputs[3223]);
    assign outputs[8720] = layer0_outputs[8296];
    assign outputs[8721] = (layer0_outputs[8368]) ^ (layer0_outputs[2713]);
    assign outputs[8722] = (layer0_outputs[2043]) | (layer0_outputs[4766]);
    assign outputs[8723] = (layer0_outputs[1517]) | (layer0_outputs[8970]);
    assign outputs[8724] = layer0_outputs[6640];
    assign outputs[8725] = ~(layer0_outputs[8359]);
    assign outputs[8726] = ~((layer0_outputs[9743]) ^ (layer0_outputs[10046]));
    assign outputs[8727] = (layer0_outputs[3349]) ^ (layer0_outputs[527]);
    assign outputs[8728] = layer0_outputs[1527];
    assign outputs[8729] = ~(layer0_outputs[851]);
    assign outputs[8730] = ~((layer0_outputs[7173]) ^ (layer0_outputs[2039]));
    assign outputs[8731] = (layer0_outputs[8519]) & ~(layer0_outputs[8346]);
    assign outputs[8732] = (layer0_outputs[9314]) ^ (layer0_outputs[7674]);
    assign outputs[8733] = layer0_outputs[1364];
    assign outputs[8734] = ~(layer0_outputs[3509]);
    assign outputs[8735] = (layer0_outputs[8487]) | (layer0_outputs[4400]);
    assign outputs[8736] = (layer0_outputs[9161]) & ~(layer0_outputs[6053]);
    assign outputs[8737] = ~(layer0_outputs[2986]) | (layer0_outputs[9982]);
    assign outputs[8738] = ~(layer0_outputs[4309]);
    assign outputs[8739] = (layer0_outputs[1496]) ^ (layer0_outputs[5880]);
    assign outputs[8740] = ~((layer0_outputs[5644]) ^ (layer0_outputs[398]));
    assign outputs[8741] = ~((layer0_outputs[9984]) & (layer0_outputs[3190]));
    assign outputs[8742] = ~(layer0_outputs[2496]);
    assign outputs[8743] = (layer0_outputs[1048]) ^ (layer0_outputs[1987]);
    assign outputs[8744] = ~(layer0_outputs[4175]) | (layer0_outputs[9306]);
    assign outputs[8745] = (layer0_outputs[1431]) ^ (layer0_outputs[6887]);
    assign outputs[8746] = layer0_outputs[4143];
    assign outputs[8747] = layer0_outputs[2839];
    assign outputs[8748] = ~(layer0_outputs[1289]);
    assign outputs[8749] = ~(layer0_outputs[8156]);
    assign outputs[8750] = (layer0_outputs[1883]) | (layer0_outputs[972]);
    assign outputs[8751] = ~(layer0_outputs[870]);
    assign outputs[8752] = layer0_outputs[1859];
    assign outputs[8753] = (layer0_outputs[2888]) ^ (layer0_outputs[7370]);
    assign outputs[8754] = layer0_outputs[8691];
    assign outputs[8755] = ~(layer0_outputs[6372]) | (layer0_outputs[2752]);
    assign outputs[8756] = (layer0_outputs[9101]) ^ (layer0_outputs[281]);
    assign outputs[8757] = ~((layer0_outputs[2463]) ^ (layer0_outputs[10174]));
    assign outputs[8758] = layer0_outputs[4759];
    assign outputs[8759] = ~((layer0_outputs[3154]) ^ (layer0_outputs[543]));
    assign outputs[8760] = ~((layer0_outputs[5113]) ^ (layer0_outputs[5542]));
    assign outputs[8761] = ~(layer0_outputs[5618]);
    assign outputs[8762] = ~(layer0_outputs[3983]);
    assign outputs[8763] = ~(layer0_outputs[8092]);
    assign outputs[8764] = ~(layer0_outputs[7183]);
    assign outputs[8765] = ~(layer0_outputs[9046]) | (layer0_outputs[6986]);
    assign outputs[8766] = ~(layer0_outputs[5584]);
    assign outputs[8767] = ~(layer0_outputs[8768]) | (layer0_outputs[5797]);
    assign outputs[8768] = ~(layer0_outputs[1248]);
    assign outputs[8769] = ~((layer0_outputs[8606]) ^ (layer0_outputs[9329]));
    assign outputs[8770] = layer0_outputs[1869];
    assign outputs[8771] = ~((layer0_outputs[2819]) ^ (layer0_outputs[6566]));
    assign outputs[8772] = ~(layer0_outputs[393]);
    assign outputs[8773] = ~((layer0_outputs[1710]) ^ (layer0_outputs[7832]));
    assign outputs[8774] = ~((layer0_outputs[8077]) ^ (layer0_outputs[2388]));
    assign outputs[8775] = ~(layer0_outputs[6328]);
    assign outputs[8776] = ~(layer0_outputs[9378]) | (layer0_outputs[647]);
    assign outputs[8777] = (layer0_outputs[4034]) ^ (layer0_outputs[4933]);
    assign outputs[8778] = (layer0_outputs[6591]) & ~(layer0_outputs[3135]);
    assign outputs[8779] = ~((layer0_outputs[2968]) | (layer0_outputs[8564]));
    assign outputs[8780] = layer0_outputs[9273];
    assign outputs[8781] = layer0_outputs[9439];
    assign outputs[8782] = ~(layer0_outputs[7355]);
    assign outputs[8783] = (layer0_outputs[7108]) & ~(layer0_outputs[2342]);
    assign outputs[8784] = (layer0_outputs[4137]) ^ (layer0_outputs[216]);
    assign outputs[8785] = ~(layer0_outputs[7949]) | (layer0_outputs[7219]);
    assign outputs[8786] = ~(layer0_outputs[4012]) | (layer0_outputs[7207]);
    assign outputs[8787] = layer0_outputs[2400];
    assign outputs[8788] = ~((layer0_outputs[1866]) ^ (layer0_outputs[4882]));
    assign outputs[8789] = (layer0_outputs[3784]) & (layer0_outputs[5283]);
    assign outputs[8790] = (layer0_outputs[9302]) ^ (layer0_outputs[2756]);
    assign outputs[8791] = ~((layer0_outputs[1909]) ^ (layer0_outputs[3032]));
    assign outputs[8792] = (layer0_outputs[8646]) & ~(layer0_outputs[1323]);
    assign outputs[8793] = (layer0_outputs[6435]) | (layer0_outputs[9002]);
    assign outputs[8794] = ~(layer0_outputs[5750]);
    assign outputs[8795] = layer0_outputs[8286];
    assign outputs[8796] = ~((layer0_outputs[6273]) ^ (layer0_outputs[4823]));
    assign outputs[8797] = ~((layer0_outputs[8201]) ^ (layer0_outputs[1520]));
    assign outputs[8798] = (layer0_outputs[3606]) ^ (layer0_outputs[6830]);
    assign outputs[8799] = (layer0_outputs[4314]) ^ (layer0_outputs[3018]);
    assign outputs[8800] = ~((layer0_outputs[1286]) ^ (layer0_outputs[85]));
    assign outputs[8801] = layer0_outputs[5650];
    assign outputs[8802] = layer0_outputs[5241];
    assign outputs[8803] = (layer0_outputs[5094]) | (layer0_outputs[618]);
    assign outputs[8804] = ~(layer0_outputs[7213]);
    assign outputs[8805] = layer0_outputs[5732];
    assign outputs[8806] = ~(layer0_outputs[2533]) | (layer0_outputs[10019]);
    assign outputs[8807] = ~((layer0_outputs[1676]) ^ (layer0_outputs[1222]));
    assign outputs[8808] = (layer0_outputs[7138]) ^ (layer0_outputs[3094]);
    assign outputs[8809] = ~(layer0_outputs[6019]);
    assign outputs[8810] = ~(layer0_outputs[393]) | (layer0_outputs[9807]);
    assign outputs[8811] = ~(layer0_outputs[1166]);
    assign outputs[8812] = ~(layer0_outputs[3143]);
    assign outputs[8813] = ~((layer0_outputs[3768]) & (layer0_outputs[2865]));
    assign outputs[8814] = (layer0_outputs[8776]) & (layer0_outputs[4962]);
    assign outputs[8815] = (layer0_outputs[8281]) | (layer0_outputs[5914]);
    assign outputs[8816] = (layer0_outputs[3906]) & ~(layer0_outputs[2755]);
    assign outputs[8817] = layer0_outputs[1886];
    assign outputs[8818] = ~((layer0_outputs[9491]) ^ (layer0_outputs[2685]));
    assign outputs[8819] = ~(layer0_outputs[1209]);
    assign outputs[8820] = (layer0_outputs[515]) ^ (layer0_outputs[5642]);
    assign outputs[8821] = ~(layer0_outputs[5791]) | (layer0_outputs[7140]);
    assign outputs[8822] = (layer0_outputs[6912]) ^ (layer0_outputs[7038]);
    assign outputs[8823] = (layer0_outputs[7111]) ^ (layer0_outputs[7374]);
    assign outputs[8824] = layer0_outputs[3263];
    assign outputs[8825] = (layer0_outputs[2574]) ^ (layer0_outputs[8974]);
    assign outputs[8826] = layer0_outputs[4570];
    assign outputs[8827] = (layer0_outputs[4168]) ^ (layer0_outputs[5716]);
    assign outputs[8828] = ~((layer0_outputs[5818]) ^ (layer0_outputs[9926]));
    assign outputs[8829] = layer0_outputs[2955];
    assign outputs[8830] = ~(layer0_outputs[7126]) | (layer0_outputs[6577]);
    assign outputs[8831] = ~(layer0_outputs[8210]);
    assign outputs[8832] = layer0_outputs[9683];
    assign outputs[8833] = ~(layer0_outputs[2640]) | (layer0_outputs[1964]);
    assign outputs[8834] = ~(layer0_outputs[3792]) | (layer0_outputs[2487]);
    assign outputs[8835] = (layer0_outputs[6571]) ^ (layer0_outputs[8386]);
    assign outputs[8836] = (layer0_outputs[3919]) ^ (layer0_outputs[7]);
    assign outputs[8837] = (layer0_outputs[8794]) | (layer0_outputs[8812]);
    assign outputs[8838] = ~((layer0_outputs[823]) ^ (layer0_outputs[4392]));
    assign outputs[8839] = ~(layer0_outputs[6946]);
    assign outputs[8840] = layer0_outputs[3471];
    assign outputs[8841] = (layer0_outputs[957]) ^ (layer0_outputs[3709]);
    assign outputs[8842] = (layer0_outputs[5617]) ^ (layer0_outputs[6060]);
    assign outputs[8843] = ~(layer0_outputs[3777]);
    assign outputs[8844] = ~(layer0_outputs[6353]);
    assign outputs[8845] = ~(layer0_outputs[6393]) | (layer0_outputs[3540]);
    assign outputs[8846] = ~(layer0_outputs[1614]);
    assign outputs[8847] = ~((layer0_outputs[1271]) ^ (layer0_outputs[9359]));
    assign outputs[8848] = layer0_outputs[1628];
    assign outputs[8849] = (layer0_outputs[7052]) & ~(layer0_outputs[3584]);
    assign outputs[8850] = layer0_outputs[7480];
    assign outputs[8851] = layer0_outputs[9552];
    assign outputs[8852] = (layer0_outputs[9347]) & (layer0_outputs[8604]);
    assign outputs[8853] = (layer0_outputs[4715]) ^ (layer0_outputs[4155]);
    assign outputs[8854] = ~(layer0_outputs[458]);
    assign outputs[8855] = layer0_outputs[5364];
    assign outputs[8856] = layer0_outputs[7684];
    assign outputs[8857] = ~(layer0_outputs[1965]);
    assign outputs[8858] = ~((layer0_outputs[114]) ^ (layer0_outputs[7221]));
    assign outputs[8859] = ~(layer0_outputs[3961]) | (layer0_outputs[332]);
    assign outputs[8860] = ~(layer0_outputs[2993]);
    assign outputs[8861] = ~(layer0_outputs[2115]);
    assign outputs[8862] = ~((layer0_outputs[3484]) & (layer0_outputs[2912]));
    assign outputs[8863] = ~(layer0_outputs[4761]);
    assign outputs[8864] = layer0_outputs[1222];
    assign outputs[8865] = (layer0_outputs[7527]) | (layer0_outputs[7540]);
    assign outputs[8866] = layer0_outputs[3691];
    assign outputs[8867] = (layer0_outputs[7462]) ^ (layer0_outputs[2305]);
    assign outputs[8868] = ~(layer0_outputs[1308]) | (layer0_outputs[5006]);
    assign outputs[8869] = (layer0_outputs[2471]) ^ (layer0_outputs[7982]);
    assign outputs[8870] = (layer0_outputs[8517]) ^ (layer0_outputs[1621]);
    assign outputs[8871] = ~(layer0_outputs[480]);
    assign outputs[8872] = ~(layer0_outputs[2837]);
    assign outputs[8873] = (layer0_outputs[7255]) & (layer0_outputs[6855]);
    assign outputs[8874] = (layer0_outputs[1533]) ^ (layer0_outputs[1474]);
    assign outputs[8875] = ~(layer0_outputs[5102]);
    assign outputs[8876] = ~((layer0_outputs[388]) ^ (layer0_outputs[1708]));
    assign outputs[8877] = (layer0_outputs[3727]) ^ (layer0_outputs[2443]);
    assign outputs[8878] = ~(layer0_outputs[8347]);
    assign outputs[8879] = layer0_outputs[6653];
    assign outputs[8880] = ~((layer0_outputs[3933]) ^ (layer0_outputs[3126]));
    assign outputs[8881] = ~((layer0_outputs[9841]) & (layer0_outputs[7634]));
    assign outputs[8882] = ~(layer0_outputs[4108]);
    assign outputs[8883] = ~((layer0_outputs[3594]) ^ (layer0_outputs[3222]));
    assign outputs[8884] = ~(layer0_outputs[164]);
    assign outputs[8885] = ~((layer0_outputs[3409]) ^ (layer0_outputs[5238]));
    assign outputs[8886] = ~((layer0_outputs[5113]) ^ (layer0_outputs[8981]));
    assign outputs[8887] = ~((layer0_outputs[3329]) ^ (layer0_outputs[1545]));
    assign outputs[8888] = ~(layer0_outputs[6604]);
    assign outputs[8889] = ~((layer0_outputs[6561]) | (layer0_outputs[890]));
    assign outputs[8890] = layer0_outputs[8187];
    assign outputs[8891] = (layer0_outputs[8268]) ^ (layer0_outputs[4158]);
    assign outputs[8892] = (layer0_outputs[7454]) & ~(layer0_outputs[4062]);
    assign outputs[8893] = ~(layer0_outputs[511]) | (layer0_outputs[5899]);
    assign outputs[8894] = ~((layer0_outputs[7112]) & (layer0_outputs[5360]));
    assign outputs[8895] = layer0_outputs[1921];
    assign outputs[8896] = ~(layer0_outputs[4509]);
    assign outputs[8897] = ~(layer0_outputs[9549]);
    assign outputs[8898] = layer0_outputs[4944];
    assign outputs[8899] = ~((layer0_outputs[9332]) & (layer0_outputs[1690]));
    assign outputs[8900] = ~(layer0_outputs[9109]);
    assign outputs[8901] = (layer0_outputs[4137]) ^ (layer0_outputs[1853]);
    assign outputs[8902] = ~(layer0_outputs[9942]) | (layer0_outputs[2768]);
    assign outputs[8903] = (layer0_outputs[6179]) | (layer0_outputs[4898]);
    assign outputs[8904] = ~(layer0_outputs[8757]);
    assign outputs[8905] = ~(layer0_outputs[8100]) | (layer0_outputs[7900]);
    assign outputs[8906] = ~(layer0_outputs[7132]);
    assign outputs[8907] = ~((layer0_outputs[3257]) ^ (layer0_outputs[6641]));
    assign outputs[8908] = ~((layer0_outputs[3080]) | (layer0_outputs[9854]));
    assign outputs[8909] = ~(layer0_outputs[248]) | (layer0_outputs[392]);
    assign outputs[8910] = layer0_outputs[6972];
    assign outputs[8911] = (layer0_outputs[6590]) ^ (layer0_outputs[3668]);
    assign outputs[8912] = ~((layer0_outputs[1405]) ^ (layer0_outputs[2769]));
    assign outputs[8913] = ~(layer0_outputs[8904]) | (layer0_outputs[3620]);
    assign outputs[8914] = layer0_outputs[1030];
    assign outputs[8915] = ~(layer0_outputs[2493]);
    assign outputs[8916] = ~(layer0_outputs[4990]);
    assign outputs[8917] = ~((layer0_outputs[6963]) ^ (layer0_outputs[5446]));
    assign outputs[8918] = ~(layer0_outputs[6040]) | (layer0_outputs[3165]);
    assign outputs[8919] = ~(layer0_outputs[6538]);
    assign outputs[8920] = ~(layer0_outputs[3137]) | (layer0_outputs[2663]);
    assign outputs[8921] = ~((layer0_outputs[836]) ^ (layer0_outputs[9123]));
    assign outputs[8922] = layer0_outputs[8677];
    assign outputs[8923] = layer0_outputs[236];
    assign outputs[8924] = ~(layer0_outputs[2995]);
    assign outputs[8925] = (layer0_outputs[9711]) & ~(layer0_outputs[7003]);
    assign outputs[8926] = ~((layer0_outputs[8092]) ^ (layer0_outputs[8310]));
    assign outputs[8927] = (layer0_outputs[9219]) | (layer0_outputs[8370]);
    assign outputs[8928] = ~(layer0_outputs[828]);
    assign outputs[8929] = ~(layer0_outputs[610]) | (layer0_outputs[5793]);
    assign outputs[8930] = (layer0_outputs[3997]) ^ (layer0_outputs[6319]);
    assign outputs[8931] = ~(layer0_outputs[7423]) | (layer0_outputs[8924]);
    assign outputs[8932] = ~((layer0_outputs[8267]) ^ (layer0_outputs[9853]));
    assign outputs[8933] = (layer0_outputs[6455]) & ~(layer0_outputs[3971]);
    assign outputs[8934] = ~(layer0_outputs[5964]);
    assign outputs[8935] = layer0_outputs[8621];
    assign outputs[8936] = (layer0_outputs[9631]) ^ (layer0_outputs[5659]);
    assign outputs[8937] = layer0_outputs[6403];
    assign outputs[8938] = ~(layer0_outputs[95]);
    assign outputs[8939] = ~(layer0_outputs[2889]);
    assign outputs[8940] = (layer0_outputs[385]) | (layer0_outputs[881]);
    assign outputs[8941] = (layer0_outputs[5594]) ^ (layer0_outputs[2849]);
    assign outputs[8942] = (layer0_outputs[8546]) | (layer0_outputs[7604]);
    assign outputs[8943] = 1'b1;
    assign outputs[8944] = (layer0_outputs[944]) & (layer0_outputs[1697]);
    assign outputs[8945] = layer0_outputs[4041];
    assign outputs[8946] = (layer0_outputs[4612]) ^ (layer0_outputs[8517]);
    assign outputs[8947] = ~((layer0_outputs[1960]) ^ (layer0_outputs[2891]));
    assign outputs[8948] = (layer0_outputs[9057]) ^ (layer0_outputs[2877]);
    assign outputs[8949] = layer0_outputs[6958];
    assign outputs[8950] = ~((layer0_outputs[1803]) ^ (layer0_outputs[4471]));
    assign outputs[8951] = (layer0_outputs[5331]) & ~(layer0_outputs[5992]);
    assign outputs[8952] = (layer0_outputs[3948]) & (layer0_outputs[2318]);
    assign outputs[8953] = layer0_outputs[668];
    assign outputs[8954] = ~(layer0_outputs[6891]);
    assign outputs[8955] = ~(layer0_outputs[10062]) | (layer0_outputs[2015]);
    assign outputs[8956] = (layer0_outputs[3656]) ^ (layer0_outputs[1159]);
    assign outputs[8957] = ~((layer0_outputs[5933]) ^ (layer0_outputs[7638]));
    assign outputs[8958] = ~(layer0_outputs[807]);
    assign outputs[8959] = (layer0_outputs[168]) & ~(layer0_outputs[6841]);
    assign outputs[8960] = (layer0_outputs[10009]) & ~(layer0_outputs[2319]);
    assign outputs[8961] = ~(layer0_outputs[3488]);
    assign outputs[8962] = ~((layer0_outputs[2363]) | (layer0_outputs[8662]));
    assign outputs[8963] = ~(layer0_outputs[1303]);
    assign outputs[8964] = (layer0_outputs[5945]) ^ (layer0_outputs[1933]);
    assign outputs[8965] = layer0_outputs[3600];
    assign outputs[8966] = (layer0_outputs[3486]) ^ (layer0_outputs[581]);
    assign outputs[8967] = ~(layer0_outputs[6983]);
    assign outputs[8968] = ~(layer0_outputs[9064]) | (layer0_outputs[8456]);
    assign outputs[8969] = (layer0_outputs[166]) ^ (layer0_outputs[1204]);
    assign outputs[8970] = ~(layer0_outputs[6452]);
    assign outputs[8971] = ~((layer0_outputs[976]) ^ (layer0_outputs[4339]));
    assign outputs[8972] = ~((layer0_outputs[4015]) & (layer0_outputs[5447]));
    assign outputs[8973] = ~((layer0_outputs[4424]) & (layer0_outputs[6816]));
    assign outputs[8974] = ~(layer0_outputs[5498]);
    assign outputs[8975] = layer0_outputs[4748];
    assign outputs[8976] = ~((layer0_outputs[7393]) ^ (layer0_outputs[2137]));
    assign outputs[8977] = layer0_outputs[6172];
    assign outputs[8978] = ~((layer0_outputs[617]) ^ (layer0_outputs[7867]));
    assign outputs[8979] = ~(layer0_outputs[6386]) | (layer0_outputs[10067]);
    assign outputs[8980] = (layer0_outputs[3310]) ^ (layer0_outputs[1557]);
    assign outputs[8981] = ~(layer0_outputs[2745]) | (layer0_outputs[5267]);
    assign outputs[8982] = layer0_outputs[5766];
    assign outputs[8983] = ~(layer0_outputs[9746]) | (layer0_outputs[3872]);
    assign outputs[8984] = (layer0_outputs[6734]) & (layer0_outputs[2250]);
    assign outputs[8985] = ~(layer0_outputs[2849]);
    assign outputs[8986] = ~(layer0_outputs[2604]) | (layer0_outputs[278]);
    assign outputs[8987] = ~(layer0_outputs[4453]);
    assign outputs[8988] = ~(layer0_outputs[9259]);
    assign outputs[8989] = ~(layer0_outputs[6093]);
    assign outputs[8990] = ~(layer0_outputs[4289]);
    assign outputs[8991] = layer0_outputs[8060];
    assign outputs[8992] = (layer0_outputs[7820]) | (layer0_outputs[5645]);
    assign outputs[8993] = (layer0_outputs[6893]) ^ (layer0_outputs[4781]);
    assign outputs[8994] = ~(layer0_outputs[9448]);
    assign outputs[8995] = ~((layer0_outputs[5251]) | (layer0_outputs[5544]));
    assign outputs[8996] = layer0_outputs[1359];
    assign outputs[8997] = (layer0_outputs[2760]) ^ (layer0_outputs[8848]);
    assign outputs[8998] = layer0_outputs[7930];
    assign outputs[8999] = layer0_outputs[1290];
    assign outputs[9000] = (layer0_outputs[4827]) | (layer0_outputs[2014]);
    assign outputs[9001] = ~((layer0_outputs[5735]) ^ (layer0_outputs[7525]));
    assign outputs[9002] = layer0_outputs[819];
    assign outputs[9003] = (layer0_outputs[718]) & (layer0_outputs[7549]);
    assign outputs[9004] = ~((layer0_outputs[5985]) & (layer0_outputs[373]));
    assign outputs[9005] = ~((layer0_outputs[1621]) & (layer0_outputs[912]));
    assign outputs[9006] = 1'b0;
    assign outputs[9007] = layer0_outputs[418];
    assign outputs[9008] = ~(layer0_outputs[3463]) | (layer0_outputs[6316]);
    assign outputs[9009] = ~(layer0_outputs[5787]);
    assign outputs[9010] = (layer0_outputs[2881]) & (layer0_outputs[4048]);
    assign outputs[9011] = ~(layer0_outputs[3345]);
    assign outputs[9012] = ~((layer0_outputs[2215]) ^ (layer0_outputs[1882]));
    assign outputs[9013] = ~(layer0_outputs[8356]);
    assign outputs[9014] = ~((layer0_outputs[8391]) ^ (layer0_outputs[20]));
    assign outputs[9015] = ~((layer0_outputs[6418]) ^ (layer0_outputs[7513]));
    assign outputs[9016] = (layer0_outputs[6291]) ^ (layer0_outputs[2018]);
    assign outputs[9017] = ~(layer0_outputs[8151]) | (layer0_outputs[7175]);
    assign outputs[9018] = ~(layer0_outputs[6623]) | (layer0_outputs[7457]);
    assign outputs[9019] = ~((layer0_outputs[9652]) & (layer0_outputs[7367]));
    assign outputs[9020] = ~(layer0_outputs[5470]) | (layer0_outputs[4123]);
    assign outputs[9021] = ~(layer0_outputs[6716]) | (layer0_outputs[190]);
    assign outputs[9022] = (layer0_outputs[7104]) ^ (layer0_outputs[8961]);
    assign outputs[9023] = layer0_outputs[181];
    assign outputs[9024] = layer0_outputs[3778];
    assign outputs[9025] = ~((layer0_outputs[4478]) & (layer0_outputs[1256]));
    assign outputs[9026] = ~(layer0_outputs[10084]) | (layer0_outputs[6245]);
    assign outputs[9027] = ~(layer0_outputs[2160]) | (layer0_outputs[2055]);
    assign outputs[9028] = ~(layer0_outputs[59]) | (layer0_outputs[5767]);
    assign outputs[9029] = ~((layer0_outputs[5135]) ^ (layer0_outputs[6901]));
    assign outputs[9030] = ~((layer0_outputs[6103]) ^ (layer0_outputs[650]));
    assign outputs[9031] = ~((layer0_outputs[1791]) ^ (layer0_outputs[3968]));
    assign outputs[9032] = ~(layer0_outputs[7049]);
    assign outputs[9033] = ~((layer0_outputs[5776]) ^ (layer0_outputs[523]));
    assign outputs[9034] = ~(layer0_outputs[7627]);
    assign outputs[9035] = layer0_outputs[7735];
    assign outputs[9036] = ~(layer0_outputs[4525]);
    assign outputs[9037] = (layer0_outputs[4406]) & (layer0_outputs[918]);
    assign outputs[9038] = (layer0_outputs[5070]) & (layer0_outputs[7283]);
    assign outputs[9039] = layer0_outputs[7162];
    assign outputs[9040] = layer0_outputs[2200];
    assign outputs[9041] = 1'b0;
    assign outputs[9042] = ~(layer0_outputs[3012]);
    assign outputs[9043] = 1'b0;
    assign outputs[9044] = (layer0_outputs[3157]) ^ (layer0_outputs[5357]);
    assign outputs[9045] = ~((layer0_outputs[6209]) ^ (layer0_outputs[5017]));
    assign outputs[9046] = ~((layer0_outputs[879]) & (layer0_outputs[493]));
    assign outputs[9047] = layer0_outputs[357];
    assign outputs[9048] = (layer0_outputs[2412]) ^ (layer0_outputs[5759]);
    assign outputs[9049] = ~(layer0_outputs[3283]);
    assign outputs[9050] = ~((layer0_outputs[5126]) ^ (layer0_outputs[9940]));
    assign outputs[9051] = layer0_outputs[4098];
    assign outputs[9052] = ~(layer0_outputs[9867]);
    assign outputs[9053] = ~(layer0_outputs[2095]);
    assign outputs[9054] = (layer0_outputs[5299]) ^ (layer0_outputs[6994]);
    assign outputs[9055] = layer0_outputs[9137];
    assign outputs[9056] = (layer0_outputs[5761]) & ~(layer0_outputs[2271]);
    assign outputs[9057] = ~(layer0_outputs[6779]);
    assign outputs[9058] = ~((layer0_outputs[7268]) ^ (layer0_outputs[10128]));
    assign outputs[9059] = (layer0_outputs[4838]) ^ (layer0_outputs[5507]);
    assign outputs[9060] = ~(layer0_outputs[3125]);
    assign outputs[9061] = layer0_outputs[1462];
    assign outputs[9062] = ~(layer0_outputs[1831]);
    assign outputs[9063] = layer0_outputs[5005];
    assign outputs[9064] = ~(layer0_outputs[4743]);
    assign outputs[9065] = (layer0_outputs[5514]) & ~(layer0_outputs[4260]);
    assign outputs[9066] = ~(layer0_outputs[9676]) | (layer0_outputs[4907]);
    assign outputs[9067] = ~((layer0_outputs[1203]) ^ (layer0_outputs[9734]));
    assign outputs[9068] = 1'b1;
    assign outputs[9069] = ~(layer0_outputs[9409]);
    assign outputs[9070] = 1'b1;
    assign outputs[9071] = layer0_outputs[6796];
    assign outputs[9072] = layer0_outputs[591];
    assign outputs[9073] = layer0_outputs[7726];
    assign outputs[9074] = ~((layer0_outputs[4141]) ^ (layer0_outputs[2151]));
    assign outputs[9075] = ~((layer0_outputs[1760]) ^ (layer0_outputs[4915]));
    assign outputs[9076] = layer0_outputs[757];
    assign outputs[9077] = ~(layer0_outputs[7666]) | (layer0_outputs[8394]);
    assign outputs[9078] = ~((layer0_outputs[6666]) ^ (layer0_outputs[3917]));
    assign outputs[9079] = (layer0_outputs[5552]) ^ (layer0_outputs[298]);
    assign outputs[9080] = (layer0_outputs[1231]) & ~(layer0_outputs[3102]);
    assign outputs[9081] = ~((layer0_outputs[5735]) & (layer0_outputs[4099]));
    assign outputs[9082] = ~(layer0_outputs[3715]);
    assign outputs[9083] = (layer0_outputs[2024]) ^ (layer0_outputs[937]);
    assign outputs[9084] = ~(layer0_outputs[7173]) | (layer0_outputs[4431]);
    assign outputs[9085] = ~(layer0_outputs[6802]);
    assign outputs[9086] = (layer0_outputs[1342]) | (layer0_outputs[8884]);
    assign outputs[9087] = ~(layer0_outputs[1482]);
    assign outputs[9088] = ~(layer0_outputs[7612]) | (layer0_outputs[950]);
    assign outputs[9089] = (layer0_outputs[4769]) ^ (layer0_outputs[9215]);
    assign outputs[9090] = ~((layer0_outputs[2255]) ^ (layer0_outputs[6850]));
    assign outputs[9091] = ~((layer0_outputs[5079]) ^ (layer0_outputs[2850]));
    assign outputs[9092] = ~((layer0_outputs[7307]) ^ (layer0_outputs[2908]));
    assign outputs[9093] = layer0_outputs[5062];
    assign outputs[9094] = ~(layer0_outputs[6637]) | (layer0_outputs[10059]);
    assign outputs[9095] = (layer0_outputs[84]) ^ (layer0_outputs[5237]);
    assign outputs[9096] = ~(layer0_outputs[7049]);
    assign outputs[9097] = ~(layer0_outputs[7622]);
    assign outputs[9098] = (layer0_outputs[5817]) & ~(layer0_outputs[4217]);
    assign outputs[9099] = ~((layer0_outputs[3701]) ^ (layer0_outputs[2697]));
    assign outputs[9100] = layer0_outputs[5698];
    assign outputs[9101] = ~((layer0_outputs[9281]) ^ (layer0_outputs[4221]));
    assign outputs[9102] = (layer0_outputs[9727]) ^ (layer0_outputs[4780]);
    assign outputs[9103] = ~((layer0_outputs[9103]) ^ (layer0_outputs[4592]));
    assign outputs[9104] = (layer0_outputs[350]) & ~(layer0_outputs[8487]);
    assign outputs[9105] = (layer0_outputs[1040]) ^ (layer0_outputs[5647]);
    assign outputs[9106] = ~(layer0_outputs[4398]);
    assign outputs[9107] = ~(layer0_outputs[1594]) | (layer0_outputs[4531]);
    assign outputs[9108] = layer0_outputs[3734];
    assign outputs[9109] = (layer0_outputs[3992]) & ~(layer0_outputs[185]);
    assign outputs[9110] = (layer0_outputs[697]) & (layer0_outputs[7246]);
    assign outputs[9111] = ~(layer0_outputs[715]);
    assign outputs[9112] = layer0_outputs[5763];
    assign outputs[9113] = ~((layer0_outputs[3850]) & (layer0_outputs[9126]));
    assign outputs[9114] = (layer0_outputs[1063]) ^ (layer0_outputs[38]);
    assign outputs[9115] = 1'b1;
    assign outputs[9116] = layer0_outputs[5909];
    assign outputs[9117] = (layer0_outputs[6990]) ^ (layer0_outputs[9872]);
    assign outputs[9118] = ~((layer0_outputs[9204]) ^ (layer0_outputs[7333]));
    assign outputs[9119] = (layer0_outputs[4006]) ^ (layer0_outputs[3761]);
    assign outputs[9120] = layer0_outputs[7055];
    assign outputs[9121] = (layer0_outputs[5200]) ^ (layer0_outputs[7535]);
    assign outputs[9122] = layer0_outputs[5503];
    assign outputs[9123] = ~((layer0_outputs[5779]) ^ (layer0_outputs[6760]));
    assign outputs[9124] = ~(layer0_outputs[8647]);
    assign outputs[9125] = ~(layer0_outputs[6894]);
    assign outputs[9126] = ~(layer0_outputs[6101]);
    assign outputs[9127] = ~(layer0_outputs[9412]);
    assign outputs[9128] = ~(layer0_outputs[1935]);
    assign outputs[9129] = (layer0_outputs[1486]) | (layer0_outputs[6532]);
    assign outputs[9130] = layer0_outputs[7300];
    assign outputs[9131] = (layer0_outputs[3417]) ^ (layer0_outputs[2635]);
    assign outputs[9132] = layer0_outputs[9567];
    assign outputs[9133] = ~((layer0_outputs[9607]) | (layer0_outputs[3928]));
    assign outputs[9134] = ~(layer0_outputs[1511]);
    assign outputs[9135] = ~((layer0_outputs[4066]) & (layer0_outputs[2386]));
    assign outputs[9136] = layer0_outputs[5004];
    assign outputs[9137] = layer0_outputs[7991];
    assign outputs[9138] = ~(layer0_outputs[9086]);
    assign outputs[9139] = ~((layer0_outputs[1783]) ^ (layer0_outputs[9158]));
    assign outputs[9140] = ~(layer0_outputs[840]) | (layer0_outputs[5838]);
    assign outputs[9141] = ~(layer0_outputs[2334]);
    assign outputs[9142] = ~((layer0_outputs[6923]) ^ (layer0_outputs[4504]));
    assign outputs[9143] = layer0_outputs[5347];
    assign outputs[9144] = (layer0_outputs[5903]) | (layer0_outputs[5414]);
    assign outputs[9145] = ~((layer0_outputs[8496]) | (layer0_outputs[1113]));
    assign outputs[9146] = (layer0_outputs[5968]) | (layer0_outputs[9674]);
    assign outputs[9147] = layer0_outputs[5793];
    assign outputs[9148] = ~((layer0_outputs[9081]) ^ (layer0_outputs[2397]));
    assign outputs[9149] = ~(layer0_outputs[9311]);
    assign outputs[9150] = ~((layer0_outputs[8498]) ^ (layer0_outputs[4468]));
    assign outputs[9151] = ~((layer0_outputs[8535]) ^ (layer0_outputs[769]));
    assign outputs[9152] = (layer0_outputs[2997]) | (layer0_outputs[4304]);
    assign outputs[9153] = ~(layer0_outputs[830]);
    assign outputs[9154] = ~(layer0_outputs[7545]);
    assign outputs[9155] = layer0_outputs[6298];
    assign outputs[9156] = (layer0_outputs[8799]) & ~(layer0_outputs[4849]);
    assign outputs[9157] = ~(layer0_outputs[5166]);
    assign outputs[9158] = ~((layer0_outputs[5627]) ^ (layer0_outputs[1561]));
    assign outputs[9159] = ~(layer0_outputs[3746]);
    assign outputs[9160] = ~((layer0_outputs[8333]) ^ (layer0_outputs[2717]));
    assign outputs[9161] = ~(layer0_outputs[8249]);
    assign outputs[9162] = ~((layer0_outputs[3019]) ^ (layer0_outputs[8031]));
    assign outputs[9163] = (layer0_outputs[4602]) ^ (layer0_outputs[8458]);
    assign outputs[9164] = ~((layer0_outputs[5091]) | (layer0_outputs[3987]));
    assign outputs[9165] = layer0_outputs[5483];
    assign outputs[9166] = ~((layer0_outputs[1447]) & (layer0_outputs[9485]));
    assign outputs[9167] = ~(layer0_outputs[4503]);
    assign outputs[9168] = (layer0_outputs[6156]) ^ (layer0_outputs[7566]);
    assign outputs[9169] = ~((layer0_outputs[5107]) ^ (layer0_outputs[9313]));
    assign outputs[9170] = ~(layer0_outputs[2572]);
    assign outputs[9171] = ~((layer0_outputs[151]) ^ (layer0_outputs[5292]));
    assign outputs[9172] = ~(layer0_outputs[703]);
    assign outputs[9173] = ~(layer0_outputs[5738]) | (layer0_outputs[9257]);
    assign outputs[9174] = ~(layer0_outputs[4584]);
    assign outputs[9175] = ~(layer0_outputs[8388]);
    assign outputs[9176] = ~(layer0_outputs[2478]);
    assign outputs[9177] = layer0_outputs[4074];
    assign outputs[9178] = layer0_outputs[9508];
    assign outputs[9179] = layer0_outputs[2706];
    assign outputs[9180] = ~((layer0_outputs[6711]) ^ (layer0_outputs[3519]));
    assign outputs[9181] = ~(layer0_outputs[1761]);
    assign outputs[9182] = ~((layer0_outputs[162]) ^ (layer0_outputs[4706]));
    assign outputs[9183] = (layer0_outputs[1514]) & (layer0_outputs[9553]);
    assign outputs[9184] = (layer0_outputs[7863]) ^ (layer0_outputs[9522]);
    assign outputs[9185] = (layer0_outputs[5369]) & (layer0_outputs[1333]);
    assign outputs[9186] = (layer0_outputs[3198]) & (layer0_outputs[9113]);
    assign outputs[9187] = ~((layer0_outputs[7934]) ^ (layer0_outputs[10222]));
    assign outputs[9188] = (layer0_outputs[607]) ^ (layer0_outputs[2404]);
    assign outputs[9189] = (layer0_outputs[80]) ^ (layer0_outputs[2640]);
    assign outputs[9190] = ~(layer0_outputs[9392]);
    assign outputs[9191] = layer0_outputs[1401];
    assign outputs[9192] = ~((layer0_outputs[2529]) ^ (layer0_outputs[9107]));
    assign outputs[9193] = ~(layer0_outputs[4808]);
    assign outputs[9194] = ~(layer0_outputs[6224]);
    assign outputs[9195] = ~(layer0_outputs[7513]) | (layer0_outputs[993]);
    assign outputs[9196] = ~((layer0_outputs[5716]) ^ (layer0_outputs[8739]));
    assign outputs[9197] = ~(layer0_outputs[5730]);
    assign outputs[9198] = layer0_outputs[4946];
    assign outputs[9199] = layer0_outputs[7946];
    assign outputs[9200] = (layer0_outputs[5002]) ^ (layer0_outputs[1883]);
    assign outputs[9201] = layer0_outputs[7059];
    assign outputs[9202] = ~(layer0_outputs[9702]) | (layer0_outputs[8040]);
    assign outputs[9203] = layer0_outputs[2976];
    assign outputs[9204] = ~((layer0_outputs[7500]) & (layer0_outputs[9996]));
    assign outputs[9205] = layer0_outputs[8990];
    assign outputs[9206] = ~(layer0_outputs[3724]);
    assign outputs[9207] = layer0_outputs[1444];
    assign outputs[9208] = ~(layer0_outputs[10111]);
    assign outputs[9209] = (layer0_outputs[3454]) ^ (layer0_outputs[7876]);
    assign outputs[9210] = ~(layer0_outputs[7959]);
    assign outputs[9211] = ~(layer0_outputs[515]) | (layer0_outputs[7332]);
    assign outputs[9212] = ~(layer0_outputs[4345]);
    assign outputs[9213] = layer0_outputs[10236];
    assign outputs[9214] = (layer0_outputs[9108]) ^ (layer0_outputs[9574]);
    assign outputs[9215] = ~((layer0_outputs[9508]) ^ (layer0_outputs[8886]));
    assign outputs[9216] = ~(layer0_outputs[3943]) | (layer0_outputs[5211]);
    assign outputs[9217] = (layer0_outputs[9222]) & ~(layer0_outputs[6287]);
    assign outputs[9218] = (layer0_outputs[7544]) & ~(layer0_outputs[5693]);
    assign outputs[9219] = ~(layer0_outputs[1913]);
    assign outputs[9220] = (layer0_outputs[1604]) & ~(layer0_outputs[2210]);
    assign outputs[9221] = layer0_outputs[6218];
    assign outputs[9222] = layer0_outputs[8797];
    assign outputs[9223] = ~(layer0_outputs[6569]);
    assign outputs[9224] = (layer0_outputs[9855]) & ~(layer0_outputs[3418]);
    assign outputs[9225] = (layer0_outputs[3678]) | (layer0_outputs[8911]);
    assign outputs[9226] = ~((layer0_outputs[5531]) & (layer0_outputs[505]));
    assign outputs[9227] = ~(layer0_outputs[6542]);
    assign outputs[9228] = layer0_outputs[9128];
    assign outputs[9229] = layer0_outputs[9968];
    assign outputs[9230] = ~((layer0_outputs[3503]) ^ (layer0_outputs[7850]));
    assign outputs[9231] = (layer0_outputs[2738]) ^ (layer0_outputs[807]);
    assign outputs[9232] = (layer0_outputs[4016]) & ~(layer0_outputs[2417]);
    assign outputs[9233] = layer0_outputs[4938];
    assign outputs[9234] = ~(layer0_outputs[6029]);
    assign outputs[9235] = layer0_outputs[477];
    assign outputs[9236] = ~((layer0_outputs[8840]) ^ (layer0_outputs[5458]));
    assign outputs[9237] = ~((layer0_outputs[9309]) ^ (layer0_outputs[4730]));
    assign outputs[9238] = ~(layer0_outputs[4408]);
    assign outputs[9239] = layer0_outputs[9141];
    assign outputs[9240] = ~(layer0_outputs[3141]);
    assign outputs[9241] = ~((layer0_outputs[3775]) | (layer0_outputs[8756]));
    assign outputs[9242] = ~(layer0_outputs[7716]);
    assign outputs[9243] = (layer0_outputs[1619]) ^ (layer0_outputs[8321]);
    assign outputs[9244] = ~((layer0_outputs[2134]) & (layer0_outputs[1146]));
    assign outputs[9245] = (layer0_outputs[877]) ^ (layer0_outputs[6301]);
    assign outputs[9246] = ~(layer0_outputs[9390]);
    assign outputs[9247] = layer0_outputs[5825];
    assign outputs[9248] = ~(layer0_outputs[7782]);
    assign outputs[9249] = layer0_outputs[9072];
    assign outputs[9250] = layer0_outputs[6039];
    assign outputs[9251] = ~(layer0_outputs[9789]);
    assign outputs[9252] = ~((layer0_outputs[2039]) ^ (layer0_outputs[4089]));
    assign outputs[9253] = (layer0_outputs[3251]) & ~(layer0_outputs[9254]);
    assign outputs[9254] = ~((layer0_outputs[5976]) ^ (layer0_outputs[3300]));
    assign outputs[9255] = ~((layer0_outputs[4821]) ^ (layer0_outputs[6381]));
    assign outputs[9256] = (layer0_outputs[8717]) & ~(layer0_outputs[1554]);
    assign outputs[9257] = ~((layer0_outputs[8035]) ^ (layer0_outputs[4832]));
    assign outputs[9258] = (layer0_outputs[604]) & (layer0_outputs[3765]);
    assign outputs[9259] = layer0_outputs[2858];
    assign outputs[9260] = ~(layer0_outputs[6872]);
    assign outputs[9261] = ~(layer0_outputs[9837]);
    assign outputs[9262] = ~(layer0_outputs[3132]);
    assign outputs[9263] = layer0_outputs[222];
    assign outputs[9264] = (layer0_outputs[4057]) & ~(layer0_outputs[4818]);
    assign outputs[9265] = (layer0_outputs[424]) & ~(layer0_outputs[3822]);
    assign outputs[9266] = (layer0_outputs[2953]) & ~(layer0_outputs[4587]);
    assign outputs[9267] = layer0_outputs[3225];
    assign outputs[9268] = (layer0_outputs[3001]) ^ (layer0_outputs[7519]);
    assign outputs[9269] = layer0_outputs[2747];
    assign outputs[9270] = (layer0_outputs[2045]) & (layer0_outputs[2838]);
    assign outputs[9271] = layer0_outputs[9831];
    assign outputs[9272] = ~((layer0_outputs[801]) ^ (layer0_outputs[2601]));
    assign outputs[9273] = ~((layer0_outputs[4467]) ^ (layer0_outputs[7754]));
    assign outputs[9274] = ~(layer0_outputs[1480]);
    assign outputs[9275] = ~(layer0_outputs[3482]);
    assign outputs[9276] = ~(layer0_outputs[3118]);
    assign outputs[9277] = (layer0_outputs[3521]) ^ (layer0_outputs[1761]);
    assign outputs[9278] = (layer0_outputs[6859]) ^ (layer0_outputs[5854]);
    assign outputs[9279] = ~(layer0_outputs[7635]);
    assign outputs[9280] = ~(layer0_outputs[843]);
    assign outputs[9281] = ~(layer0_outputs[9949]);
    assign outputs[9282] = (layer0_outputs[8203]) & (layer0_outputs[5903]);
    assign outputs[9283] = (layer0_outputs[7398]) & ~(layer0_outputs[8343]);
    assign outputs[9284] = ~(layer0_outputs[2330]);
    assign outputs[9285] = (layer0_outputs[8623]) & ~(layer0_outputs[7116]);
    assign outputs[9286] = ~(layer0_outputs[4083]);
    assign outputs[9287] = ~(layer0_outputs[10170]) | (layer0_outputs[1148]);
    assign outputs[9288] = ~((layer0_outputs[3646]) ^ (layer0_outputs[3363]));
    assign outputs[9289] = layer0_outputs[5981];
    assign outputs[9290] = (layer0_outputs[9082]) & ~(layer0_outputs[7042]);
    assign outputs[9291] = ~(layer0_outputs[3643]);
    assign outputs[9292] = (layer0_outputs[4281]) ^ (layer0_outputs[2163]);
    assign outputs[9293] = ~((layer0_outputs[4874]) | (layer0_outputs[6618]));
    assign outputs[9294] = (layer0_outputs[55]) & (layer0_outputs[2193]);
    assign outputs[9295] = (layer0_outputs[5966]) & (layer0_outputs[3291]);
    assign outputs[9296] = ~(layer0_outputs[8369]);
    assign outputs[9297] = layer0_outputs[7131];
    assign outputs[9298] = layer0_outputs[8450];
    assign outputs[9299] = ~(layer0_outputs[534]);
    assign outputs[9300] = (layer0_outputs[4231]) | (layer0_outputs[383]);
    assign outputs[9301] = layer0_outputs[5865];
    assign outputs[9302] = ~(layer0_outputs[1550]);
    assign outputs[9303] = (layer0_outputs[3924]) ^ (layer0_outputs[8717]);
    assign outputs[9304] = ~(layer0_outputs[7848]);
    assign outputs[9305] = ~(layer0_outputs[1642]);
    assign outputs[9306] = (layer0_outputs[3280]) ^ (layer0_outputs[6022]);
    assign outputs[9307] = (layer0_outputs[10210]) ^ (layer0_outputs[2126]);
    assign outputs[9308] = layer0_outputs[4149];
    assign outputs[9309] = layer0_outputs[8043];
    assign outputs[9310] = ~(layer0_outputs[9526]);
    assign outputs[9311] = ~(layer0_outputs[6477]);
    assign outputs[9312] = (layer0_outputs[1319]) & (layer0_outputs[10122]);
    assign outputs[9313] = (layer0_outputs[9055]) & ~(layer0_outputs[9600]);
    assign outputs[9314] = ~(layer0_outputs[6109]);
    assign outputs[9315] = layer0_outputs[2131];
    assign outputs[9316] = layer0_outputs[1102];
    assign outputs[9317] = ~((layer0_outputs[1361]) | (layer0_outputs[1636]));
    assign outputs[9318] = (layer0_outputs[7931]) ^ (layer0_outputs[1358]);
    assign outputs[9319] = layer0_outputs[5663];
    assign outputs[9320] = (layer0_outputs[5994]) ^ (layer0_outputs[6969]);
    assign outputs[9321] = layer0_outputs[6681];
    assign outputs[9322] = ~(layer0_outputs[9927]);
    assign outputs[9323] = (layer0_outputs[7961]) & ~(layer0_outputs[2703]);
    assign outputs[9324] = layer0_outputs[5584];
    assign outputs[9325] = ~(layer0_outputs[7036]);
    assign outputs[9326] = layer0_outputs[1623];
    assign outputs[9327] = ~((layer0_outputs[9866]) | (layer0_outputs[1268]));
    assign outputs[9328] = layer0_outputs[1673];
    assign outputs[9329] = ~((layer0_outputs[9857]) | (layer0_outputs[1283]));
    assign outputs[9330] = ~(layer0_outputs[8952]);
    assign outputs[9331] = layer0_outputs[7779];
    assign outputs[9332] = ~((layer0_outputs[2507]) ^ (layer0_outputs[4306]));
    assign outputs[9333] = ~((layer0_outputs[1977]) & (layer0_outputs[1280]));
    assign outputs[9334] = (layer0_outputs[3708]) & ~(layer0_outputs[2274]);
    assign outputs[9335] = ~(layer0_outputs[1584]);
    assign outputs[9336] = ~((layer0_outputs[9161]) ^ (layer0_outputs[4811]));
    assign outputs[9337] = ~(layer0_outputs[7001]) | (layer0_outputs[7030]);
    assign outputs[9338] = (layer0_outputs[5396]) & ~(layer0_outputs[4530]);
    assign outputs[9339] = ~((layer0_outputs[3097]) | (layer0_outputs[8973]));
    assign outputs[9340] = ~(layer0_outputs[1281]);
    assign outputs[9341] = ~(layer0_outputs[1800]);
    assign outputs[9342] = (layer0_outputs[7613]) & ~(layer0_outputs[6010]);
    assign outputs[9343] = ~(layer0_outputs[6579]);
    assign outputs[9344] = (layer0_outputs[1212]) & ~(layer0_outputs[5695]);
    assign outputs[9345] = ~(layer0_outputs[9639]);
    assign outputs[9346] = ~(layer0_outputs[8556]);
    assign outputs[9347] = ~(layer0_outputs[6853]);
    assign outputs[9348] = (layer0_outputs[3077]) ^ (layer0_outputs[8568]);
    assign outputs[9349] = (layer0_outputs[3361]) & ~(layer0_outputs[8427]);
    assign outputs[9350] = layer0_outputs[8989];
    assign outputs[9351] = (layer0_outputs[9690]) & ~(layer0_outputs[4027]);
    assign outputs[9352] = ~((layer0_outputs[6890]) | (layer0_outputs[1750]));
    assign outputs[9353] = layer0_outputs[4736];
    assign outputs[9354] = layer0_outputs[4801];
    assign outputs[9355] = (layer0_outputs[1762]) & ~(layer0_outputs[6515]);
    assign outputs[9356] = (layer0_outputs[4771]) & (layer0_outputs[115]);
    assign outputs[9357] = (layer0_outputs[3304]) & ~(layer0_outputs[2279]);
    assign outputs[9358] = ~(layer0_outputs[8958]);
    assign outputs[9359] = (layer0_outputs[6444]) & ~(layer0_outputs[1367]);
    assign outputs[9360] = layer0_outputs[5717];
    assign outputs[9361] = ~(layer0_outputs[4761]);
    assign outputs[9362] = layer0_outputs[5009];
    assign outputs[9363] = ~(layer0_outputs[7310]);
    assign outputs[9364] = ~(layer0_outputs[4246]);
    assign outputs[9365] = ~(layer0_outputs[1295]);
    assign outputs[9366] = ~((layer0_outputs[8993]) ^ (layer0_outputs[9634]));
    assign outputs[9367] = ~((layer0_outputs[2016]) | (layer0_outputs[3539]));
    assign outputs[9368] = (layer0_outputs[6583]) ^ (layer0_outputs[7037]);
    assign outputs[9369] = ~((layer0_outputs[4949]) ^ (layer0_outputs[2275]));
    assign outputs[9370] = ~(layer0_outputs[689]);
    assign outputs[9371] = (layer0_outputs[2251]) & ~(layer0_outputs[7333]);
    assign outputs[9372] = ~((layer0_outputs[5600]) | (layer0_outputs[8239]));
    assign outputs[9373] = (layer0_outputs[8826]) & ~(layer0_outputs[9163]);
    assign outputs[9374] = layer0_outputs[5441];
    assign outputs[9375] = layer0_outputs[8177];
    assign outputs[9376] = layer0_outputs[6111];
    assign outputs[9377] = (layer0_outputs[1682]) & (layer0_outputs[46]);
    assign outputs[9378] = ~(layer0_outputs[9789]);
    assign outputs[9379] = layer0_outputs[6218];
    assign outputs[9380] = ~((layer0_outputs[3175]) | (layer0_outputs[2875]));
    assign outputs[9381] = layer0_outputs[1445];
    assign outputs[9382] = (layer0_outputs[513]) & ~(layer0_outputs[5192]);
    assign outputs[9383] = (layer0_outputs[9934]) & ~(layer0_outputs[7153]);
    assign outputs[9384] = (layer0_outputs[6028]) & (layer0_outputs[7870]);
    assign outputs[9385] = ~(layer0_outputs[5477]);
    assign outputs[9386] = (layer0_outputs[8196]) & (layer0_outputs[4507]);
    assign outputs[9387] = ~((layer0_outputs[1073]) & (layer0_outputs[6964]));
    assign outputs[9388] = ~(layer0_outputs[9122]);
    assign outputs[9389] = (layer0_outputs[678]) ^ (layer0_outputs[9568]);
    assign outputs[9390] = (layer0_outputs[9175]) ^ (layer0_outputs[733]);
    assign outputs[9391] = ~((layer0_outputs[467]) ^ (layer0_outputs[1325]));
    assign outputs[9392] = (layer0_outputs[4513]) & ~(layer0_outputs[3952]);
    assign outputs[9393] = (layer0_outputs[2205]) & ~(layer0_outputs[6942]);
    assign outputs[9394] = (layer0_outputs[2047]) ^ (layer0_outputs[1318]);
    assign outputs[9395] = ~((layer0_outputs[301]) ^ (layer0_outputs[576]));
    assign outputs[9396] = ~((layer0_outputs[5538]) ^ (layer0_outputs[1619]));
    assign outputs[9397] = ~((layer0_outputs[6095]) ^ (layer0_outputs[6416]));
    assign outputs[9398] = layer0_outputs[7147];
    assign outputs[9399] = ~((layer0_outputs[1685]) | (layer0_outputs[5132]));
    assign outputs[9400] = layer0_outputs[8442];
    assign outputs[9401] = (layer0_outputs[5497]) ^ (layer0_outputs[958]);
    assign outputs[9402] = layer0_outputs[2349];
    assign outputs[9403] = (layer0_outputs[2736]) & ~(layer0_outputs[4710]);
    assign outputs[9404] = layer0_outputs[4439];
    assign outputs[9405] = ~(layer0_outputs[9379]);
    assign outputs[9406] = layer0_outputs[8251];
    assign outputs[9407] = ~(layer0_outputs[862]);
    assign outputs[9408] = ~((layer0_outputs[3307]) ^ (layer0_outputs[4830]));
    assign outputs[9409] = ~(layer0_outputs[2312]);
    assign outputs[9410] = ~((layer0_outputs[9664]) ^ (layer0_outputs[2080]));
    assign outputs[9411] = layer0_outputs[6535];
    assign outputs[9412] = ~(layer0_outputs[1742]);
    assign outputs[9413] = layer0_outputs[2209];
    assign outputs[9414] = ~(layer0_outputs[9020]);
    assign outputs[9415] = layer0_outputs[705];
    assign outputs[9416] = ~(layer0_outputs[2929]);
    assign outputs[9417] = layer0_outputs[9965];
    assign outputs[9418] = layer0_outputs[513];
    assign outputs[9419] = (layer0_outputs[2719]) ^ (layer0_outputs[9752]);
    assign outputs[9420] = (layer0_outputs[5172]) & (layer0_outputs[3673]);
    assign outputs[9421] = layer0_outputs[2153];
    assign outputs[9422] = layer0_outputs[7762];
    assign outputs[9423] = ~(layer0_outputs[82]) | (layer0_outputs[7338]);
    assign outputs[9424] = ~(layer0_outputs[4913]);
    assign outputs[9425] = (layer0_outputs[1943]) & ~(layer0_outputs[1059]);
    assign outputs[9426] = ~(layer0_outputs[1753]);
    assign outputs[9427] = ~(layer0_outputs[1831]);
    assign outputs[9428] = ~(layer0_outputs[3479]);
    assign outputs[9429] = layer0_outputs[2492];
    assign outputs[9430] = (layer0_outputs[7074]) & ~(layer0_outputs[720]);
    assign outputs[9431] = layer0_outputs[996];
    assign outputs[9432] = ~((layer0_outputs[968]) | (layer0_outputs[2301]));
    assign outputs[9433] = (layer0_outputs[10086]) & (layer0_outputs[7725]);
    assign outputs[9434] = layer0_outputs[991];
    assign outputs[9435] = layer0_outputs[7813];
    assign outputs[9436] = layer0_outputs[9663];
    assign outputs[9437] = ~((layer0_outputs[6628]) | (layer0_outputs[3144]));
    assign outputs[9438] = ~(layer0_outputs[780]);
    assign outputs[9439] = ~((layer0_outputs[7595]) | (layer0_outputs[2143]));
    assign outputs[9440] = ~(layer0_outputs[6787]);
    assign outputs[9441] = (layer0_outputs[9056]) & (layer0_outputs[8083]);
    assign outputs[9442] = ~(layer0_outputs[7425]) | (layer0_outputs[1457]);
    assign outputs[9443] = ~(layer0_outputs[8506]);
    assign outputs[9444] = layer0_outputs[2921];
    assign outputs[9445] = (layer0_outputs[7100]) | (layer0_outputs[2557]);
    assign outputs[9446] = (layer0_outputs[7152]) & (layer0_outputs[4461]);
    assign outputs[9447] = (layer0_outputs[8457]) ^ (layer0_outputs[7656]);
    assign outputs[9448] = layer0_outputs[3587];
    assign outputs[9449] = ~(layer0_outputs[4701]);
    assign outputs[9450] = (layer0_outputs[5987]) & (layer0_outputs[3074]);
    assign outputs[9451] = ~(layer0_outputs[1420]);
    assign outputs[9452] = 1'b0;
    assign outputs[9453] = (layer0_outputs[5058]) ^ (layer0_outputs[4203]);
    assign outputs[9454] = layer0_outputs[372];
    assign outputs[9455] = (layer0_outputs[649]) & (layer0_outputs[5316]);
    assign outputs[9456] = layer0_outputs[6581];
    assign outputs[9457] = ~(layer0_outputs[8225]);
    assign outputs[9458] = (layer0_outputs[7120]) & ~(layer0_outputs[8669]);
    assign outputs[9459] = ~(layer0_outputs[7620]);
    assign outputs[9460] = ~(layer0_outputs[2252]);
    assign outputs[9461] = ~((layer0_outputs[4274]) | (layer0_outputs[8808]));
    assign outputs[9462] = layer0_outputs[1316];
    assign outputs[9463] = (layer0_outputs[2441]) | (layer0_outputs[8545]);
    assign outputs[9464] = layer0_outputs[1923];
    assign outputs[9465] = ~(layer0_outputs[4248]);
    assign outputs[9466] = ~(layer0_outputs[610]);
    assign outputs[9467] = ~(layer0_outputs[18]) | (layer0_outputs[6668]);
    assign outputs[9468] = layer0_outputs[5146];
    assign outputs[9469] = layer0_outputs[9792];
    assign outputs[9470] = ~((layer0_outputs[6101]) ^ (layer0_outputs[10194]));
    assign outputs[9471] = layer0_outputs[6056];
    assign outputs[9472] = ~((layer0_outputs[7303]) ^ (layer0_outputs[8150]));
    assign outputs[9473] = ~(layer0_outputs[931]);
    assign outputs[9474] = layer0_outputs[2976];
    assign outputs[9475] = ~((layer0_outputs[4066]) | (layer0_outputs[2536]));
    assign outputs[9476] = ~(layer0_outputs[4625]);
    assign outputs[9477] = ~(layer0_outputs[766]);
    assign outputs[9478] = ~(layer0_outputs[9249]);
    assign outputs[9479] = ~(layer0_outputs[2742]) | (layer0_outputs[5142]);
    assign outputs[9480] = (layer0_outputs[3158]) & ~(layer0_outputs[7592]);
    assign outputs[9481] = ~((layer0_outputs[2729]) | (layer0_outputs[4637]));
    assign outputs[9482] = ~(layer0_outputs[2740]);
    assign outputs[9483] = (layer0_outputs[5083]) & ~(layer0_outputs[110]);
    assign outputs[9484] = ~((layer0_outputs[3437]) ^ (layer0_outputs[6083]));
    assign outputs[9485] = ~(layer0_outputs[6914]);
    assign outputs[9486] = ~((layer0_outputs[8416]) ^ (layer0_outputs[10149]));
    assign outputs[9487] = ~(layer0_outputs[7661]);
    assign outputs[9488] = (layer0_outputs[8713]) & (layer0_outputs[4120]);
    assign outputs[9489] = ~((layer0_outputs[8598]) ^ (layer0_outputs[1660]));
    assign outputs[9490] = layer0_outputs[3495];
    assign outputs[9491] = layer0_outputs[4410];
    assign outputs[9492] = ~(layer0_outputs[7058]);
    assign outputs[9493] = (layer0_outputs[9021]) ^ (layer0_outputs[2513]);
    assign outputs[9494] = (layer0_outputs[9027]) & ~(layer0_outputs[7339]);
    assign outputs[9495] = layer0_outputs[2025];
    assign outputs[9496] = ~(layer0_outputs[8845]);
    assign outputs[9497] = (layer0_outputs[6678]) & (layer0_outputs[6438]);
    assign outputs[9498] = layer0_outputs[8976];
    assign outputs[9499] = (layer0_outputs[2896]) ^ (layer0_outputs[6905]);
    assign outputs[9500] = ~(layer0_outputs[640]);
    assign outputs[9501] = (layer0_outputs[8366]) & ~(layer0_outputs[1084]);
    assign outputs[9502] = (layer0_outputs[4870]) & ~(layer0_outputs[1117]);
    assign outputs[9503] = ~((layer0_outputs[8548]) ^ (layer0_outputs[8457]));
    assign outputs[9504] = ~((layer0_outputs[9075]) | (layer0_outputs[9733]));
    assign outputs[9505] = (layer0_outputs[6493]) & ~(layer0_outputs[4550]);
    assign outputs[9506] = ~((layer0_outputs[9777]) & (layer0_outputs[9913]));
    assign outputs[9507] = ~(layer0_outputs[8023]);
    assign outputs[9508] = ~((layer0_outputs[2514]) | (layer0_outputs[7037]));
    assign outputs[9509] = layer0_outputs[873];
    assign outputs[9510] = ~(layer0_outputs[3417]);
    assign outputs[9511] = layer0_outputs[9214];
    assign outputs[9512] = layer0_outputs[8313];
    assign outputs[9513] = ~((layer0_outputs[9320]) | (layer0_outputs[10047]));
    assign outputs[9514] = (layer0_outputs[5050]) & ~(layer0_outputs[9696]);
    assign outputs[9515] = layer0_outputs[1125];
    assign outputs[9516] = ~(layer0_outputs[6194]);
    assign outputs[9517] = ~((layer0_outputs[8467]) ^ (layer0_outputs[763]));
    assign outputs[9518] = layer0_outputs[121];
    assign outputs[9519] = layer0_outputs[8950];
    assign outputs[9520] = (layer0_outputs[4257]) ^ (layer0_outputs[7920]);
    assign outputs[9521] = (layer0_outputs[6114]) ^ (layer0_outputs[5448]);
    assign outputs[9522] = layer0_outputs[7707];
    assign outputs[9523] = ~(layer0_outputs[5304]) | (layer0_outputs[9184]);
    assign outputs[9524] = ~((layer0_outputs[7599]) ^ (layer0_outputs[2366]));
    assign outputs[9525] = ~(layer0_outputs[411]) | (layer0_outputs[7499]);
    assign outputs[9526] = ~(layer0_outputs[1327]);
    assign outputs[9527] = ~(layer0_outputs[2373]);
    assign outputs[9528] = ~((layer0_outputs[5568]) ^ (layer0_outputs[9058]));
    assign outputs[9529] = (layer0_outputs[8568]) & ~(layer0_outputs[8066]);
    assign outputs[9530] = ~((layer0_outputs[3086]) ^ (layer0_outputs[1647]));
    assign outputs[9531] = ~((layer0_outputs[3658]) ^ (layer0_outputs[5356]));
    assign outputs[9532] = layer0_outputs[4758];
    assign outputs[9533] = (layer0_outputs[8529]) ^ (layer0_outputs[4788]);
    assign outputs[9534] = layer0_outputs[3388];
    assign outputs[9535] = layer0_outputs[9784];
    assign outputs[9536] = ~((layer0_outputs[3531]) | (layer0_outputs[2798]));
    assign outputs[9537] = layer0_outputs[7081];
    assign outputs[9538] = ~(layer0_outputs[6225]);
    assign outputs[9539] = ~((layer0_outputs[10101]) | (layer0_outputs[5880]));
    assign outputs[9540] = ~((layer0_outputs[9533]) ^ (layer0_outputs[9174]));
    assign outputs[9541] = (layer0_outputs[3160]) | (layer0_outputs[5789]);
    assign outputs[9542] = layer0_outputs[1195];
    assign outputs[9543] = ~((layer0_outputs[3093]) ^ (layer0_outputs[1458]));
    assign outputs[9544] = layer0_outputs[7601];
    assign outputs[9545] = layer0_outputs[2222];
    assign outputs[9546] = layer0_outputs[9353];
    assign outputs[9547] = ~(layer0_outputs[5586]);
    assign outputs[9548] = ~(layer0_outputs[6567]);
    assign outputs[9549] = (layer0_outputs[5070]) & ~(layer0_outputs[671]);
    assign outputs[9550] = layer0_outputs[824];
    assign outputs[9551] = ~(layer0_outputs[6185]);
    assign outputs[9552] = layer0_outputs[2622];
    assign outputs[9553] = ~((layer0_outputs[5656]) ^ (layer0_outputs[10048]));
    assign outputs[9554] = (layer0_outputs[4421]) | (layer0_outputs[5890]);
    assign outputs[9555] = (layer0_outputs[3371]) ^ (layer0_outputs[8112]);
    assign outputs[9556] = ~((layer0_outputs[5957]) ^ (layer0_outputs[3525]));
    assign outputs[9557] = (layer0_outputs[9732]) | (layer0_outputs[5393]);
    assign outputs[9558] = (layer0_outputs[2584]) | (layer0_outputs[7818]);
    assign outputs[9559] = ~(layer0_outputs[4696]);
    assign outputs[9560] = (layer0_outputs[10180]) ^ (layer0_outputs[6868]);
    assign outputs[9561] = layer0_outputs[4315];
    assign outputs[9562] = layer0_outputs[3874];
    assign outputs[9563] = ~(layer0_outputs[6417]);
    assign outputs[9564] = (layer0_outputs[216]) & (layer0_outputs[8942]);
    assign outputs[9565] = (layer0_outputs[8608]) ^ (layer0_outputs[6135]);
    assign outputs[9566] = (layer0_outputs[1168]) & ~(layer0_outputs[7881]);
    assign outputs[9567] = ~((layer0_outputs[4167]) ^ (layer0_outputs[5908]));
    assign outputs[9568] = ~((layer0_outputs[2530]) ^ (layer0_outputs[10142]));
    assign outputs[9569] = ~(layer0_outputs[3933]);
    assign outputs[9570] = layer0_outputs[1542];
    assign outputs[9571] = ~(layer0_outputs[3652]) | (layer0_outputs[2824]);
    assign outputs[9572] = layer0_outputs[4347];
    assign outputs[9573] = (layer0_outputs[6541]) & (layer0_outputs[9269]);
    assign outputs[9574] = (layer0_outputs[2197]) ^ (layer0_outputs[5993]);
    assign outputs[9575] = (layer0_outputs[6176]) ^ (layer0_outputs[9319]);
    assign outputs[9576] = (layer0_outputs[2704]) & ~(layer0_outputs[4121]);
    assign outputs[9577] = (layer0_outputs[3547]) & ~(layer0_outputs[3638]);
    assign outputs[9578] = (layer0_outputs[9564]) & (layer0_outputs[520]);
    assign outputs[9579] = ~((layer0_outputs[5453]) ^ (layer0_outputs[8311]));
    assign outputs[9580] = (layer0_outputs[2434]) | (layer0_outputs[8384]);
    assign outputs[9581] = layer0_outputs[1744];
    assign outputs[9582] = ~(layer0_outputs[5683]);
    assign outputs[9583] = ~((layer0_outputs[1162]) | (layer0_outputs[3683]));
    assign outputs[9584] = (layer0_outputs[3828]) | (layer0_outputs[3970]);
    assign outputs[9585] = (layer0_outputs[5535]) & (layer0_outputs[958]);
    assign outputs[9586] = ~(layer0_outputs[5851]) | (layer0_outputs[5612]);
    assign outputs[9587] = (layer0_outputs[5816]) & (layer0_outputs[7231]);
    assign outputs[9588] = ~(layer0_outputs[808]);
    assign outputs[9589] = layer0_outputs[1390];
    assign outputs[9590] = ~(layer0_outputs[9247]);
    assign outputs[9591] = ~(layer0_outputs[10163]);
    assign outputs[9592] = layer0_outputs[8174];
    assign outputs[9593] = ~(layer0_outputs[4142]) | (layer0_outputs[6632]);
    assign outputs[9594] = ~(layer0_outputs[6142]);
    assign outputs[9595] = ~(layer0_outputs[3825]) | (layer0_outputs[678]);
    assign outputs[9596] = ~((layer0_outputs[6564]) ^ (layer0_outputs[5576]));
    assign outputs[9597] = (layer0_outputs[6577]) ^ (layer0_outputs[2283]);
    assign outputs[9598] = ~(layer0_outputs[3199]) | (layer0_outputs[6062]);
    assign outputs[9599] = ~((layer0_outputs[2637]) | (layer0_outputs[1586]));
    assign outputs[9600] = ~(layer0_outputs[5477]);
    assign outputs[9601] = (layer0_outputs[3576]) & ~(layer0_outputs[673]);
    assign outputs[9602] = ~((layer0_outputs[750]) | (layer0_outputs[9764]));
    assign outputs[9603] = layer0_outputs[7512];
    assign outputs[9604] = ~(layer0_outputs[3020]);
    assign outputs[9605] = ~((layer0_outputs[5069]) & (layer0_outputs[8751]));
    assign outputs[9606] = (layer0_outputs[6683]) & ~(layer0_outputs[7539]);
    assign outputs[9607] = ~((layer0_outputs[6333]) ^ (layer0_outputs[3551]));
    assign outputs[9608] = (layer0_outputs[831]) & (layer0_outputs[1481]);
    assign outputs[9609] = (layer0_outputs[5339]) & ~(layer0_outputs[1944]);
    assign outputs[9610] = ~(layer0_outputs[3062]);
    assign outputs[9611] = (layer0_outputs[8276]) & (layer0_outputs[1405]);
    assign outputs[9612] = layer0_outputs[3500];
    assign outputs[9613] = (layer0_outputs[8297]) & (layer0_outputs[1483]);
    assign outputs[9614] = layer0_outputs[2579];
    assign outputs[9615] = ~(layer0_outputs[7973]) | (layer0_outputs[2511]);
    assign outputs[9616] = ~((layer0_outputs[7089]) ^ (layer0_outputs[2942]));
    assign outputs[9617] = ~(layer0_outputs[2614]) | (layer0_outputs[2353]);
    assign outputs[9618] = layer0_outputs[7915];
    assign outputs[9619] = ~(layer0_outputs[634]);
    assign outputs[9620] = (layer0_outputs[2876]) & (layer0_outputs[3982]);
    assign outputs[9621] = (layer0_outputs[9080]) & (layer0_outputs[5680]);
    assign outputs[9622] = ~(layer0_outputs[6736]);
    assign outputs[9623] = (layer0_outputs[5290]) | (layer0_outputs[4341]);
    assign outputs[9624] = (layer0_outputs[8119]) & ~(layer0_outputs[7402]);
    assign outputs[9625] = (layer0_outputs[281]) ^ (layer0_outputs[590]);
    assign outputs[9626] = layer0_outputs[9116];
    assign outputs[9627] = ~(layer0_outputs[1175]);
    assign outputs[9628] = ~((layer0_outputs[5459]) | (layer0_outputs[6691]));
    assign outputs[9629] = layer0_outputs[9437];
    assign outputs[9630] = (layer0_outputs[4029]) & ~(layer0_outputs[5071]);
    assign outputs[9631] = ~(layer0_outputs[7204]);
    assign outputs[9632] = (layer0_outputs[8560]) & ~(layer0_outputs[7940]);
    assign outputs[9633] = ~((layer0_outputs[7647]) | (layer0_outputs[6145]));
    assign outputs[9634] = ~((layer0_outputs[6014]) ^ (layer0_outputs[2594]));
    assign outputs[9635] = (layer0_outputs[1297]) ^ (layer0_outputs[9975]);
    assign outputs[9636] = (layer0_outputs[8955]) & (layer0_outputs[5548]);
    assign outputs[9637] = (layer0_outputs[4484]) & (layer0_outputs[9126]);
    assign outputs[9638] = ~(layer0_outputs[6517]);
    assign outputs[9639] = (layer0_outputs[5996]) & (layer0_outputs[8559]);
    assign outputs[9640] = ~((layer0_outputs[315]) ^ (layer0_outputs[6908]));
    assign outputs[9641] = ~((layer0_outputs[4102]) & (layer0_outputs[2165]));
    assign outputs[9642] = layer0_outputs[1734];
    assign outputs[9643] = ~((layer0_outputs[5815]) | (layer0_outputs[8772]));
    assign outputs[9644] = ~(layer0_outputs[574]) | (layer0_outputs[5082]);
    assign outputs[9645] = layer0_outputs[3205];
    assign outputs[9646] = ~((layer0_outputs[9232]) ^ (layer0_outputs[4089]));
    assign outputs[9647] = ~((layer0_outputs[3478]) ^ (layer0_outputs[1368]));
    assign outputs[9648] = (layer0_outputs[2199]) & ~(layer0_outputs[2292]);
    assign outputs[9649] = (layer0_outputs[5641]) & ~(layer0_outputs[4952]);
    assign outputs[9650] = (layer0_outputs[2119]) ^ (layer0_outputs[7884]);
    assign outputs[9651] = ~(layer0_outputs[1348]);
    assign outputs[9652] = (layer0_outputs[982]) & ~(layer0_outputs[3470]);
    assign outputs[9653] = layer0_outputs[8446];
    assign outputs[9654] = (layer0_outputs[147]) & ~(layer0_outputs[9755]);
    assign outputs[9655] = (layer0_outputs[1163]) & ~(layer0_outputs[5263]);
    assign outputs[9656] = ~(layer0_outputs[4481]);
    assign outputs[9657] = ~((layer0_outputs[8304]) | (layer0_outputs[6997]));
    assign outputs[9658] = (layer0_outputs[9115]) & ~(layer0_outputs[7967]);
    assign outputs[9659] = ~(layer0_outputs[9646]) | (layer0_outputs[6461]);
    assign outputs[9660] = ~(layer0_outputs[230]);
    assign outputs[9661] = (layer0_outputs[2182]) & ~(layer0_outputs[966]);
    assign outputs[9662] = ~(layer0_outputs[169]);
    assign outputs[9663] = layer0_outputs[1350];
    assign outputs[9664] = (layer0_outputs[9260]) ^ (layer0_outputs[5123]);
    assign outputs[9665] = ~((layer0_outputs[1848]) ^ (layer0_outputs[3369]));
    assign outputs[9666] = ~(layer0_outputs[7728]);
    assign outputs[9667] = layer0_outputs[1610];
    assign outputs[9668] = layer0_outputs[3713];
    assign outputs[9669] = ~((layer0_outputs[644]) ^ (layer0_outputs[1611]));
    assign outputs[9670] = ~((layer0_outputs[7287]) & (layer0_outputs[1465]));
    assign outputs[9671] = ~((layer0_outputs[8270]) & (layer0_outputs[4020]));
    assign outputs[9672] = ~(layer0_outputs[10231]);
    assign outputs[9673] = (layer0_outputs[2519]) | (layer0_outputs[8530]);
    assign outputs[9674] = ~(layer0_outputs[4189]);
    assign outputs[9675] = (layer0_outputs[7610]) & (layer0_outputs[5149]);
    assign outputs[9676] = ~(layer0_outputs[2331]);
    assign outputs[9677] = (layer0_outputs[7454]) & ~(layer0_outputs[3579]);
    assign outputs[9678] = layer0_outputs[8389];
    assign outputs[9679] = layer0_outputs[1239];
    assign outputs[9680] = ~((layer0_outputs[8469]) | (layer0_outputs[8639]));
    assign outputs[9681] = ~((layer0_outputs[10232]) ^ (layer0_outputs[4813]));
    assign outputs[9682] = (layer0_outputs[374]) ^ (layer0_outputs[7858]);
    assign outputs[9683] = layer0_outputs[2878];
    assign outputs[9684] = layer0_outputs[2954];
    assign outputs[9685] = ~(layer0_outputs[5249]);
    assign outputs[9686] = layer0_outputs[6976];
    assign outputs[9687] = (layer0_outputs[5392]) ^ (layer0_outputs[2011]);
    assign outputs[9688] = (layer0_outputs[3597]) & ~(layer0_outputs[7461]);
    assign outputs[9689] = (layer0_outputs[4357]) ^ (layer0_outputs[5313]);
    assign outputs[9690] = ~((layer0_outputs[7789]) ^ (layer0_outputs[7013]));
    assign outputs[9691] = layer0_outputs[7099];
    assign outputs[9692] = ~(layer0_outputs[8561]);
    assign outputs[9693] = ~(layer0_outputs[7537]);
    assign outputs[9694] = ~((layer0_outputs[10191]) ^ (layer0_outputs[2984]));
    assign outputs[9695] = (layer0_outputs[7196]) & ~(layer0_outputs[5025]);
    assign outputs[9696] = (layer0_outputs[5796]) ^ (layer0_outputs[9880]);
    assign outputs[9697] = ~((layer0_outputs[2781]) | (layer0_outputs[8224]));
    assign outputs[9698] = ~((layer0_outputs[8152]) ^ (layer0_outputs[633]));
    assign outputs[9699] = (layer0_outputs[929]) ^ (layer0_outputs[4308]);
    assign outputs[9700] = ~(layer0_outputs[5451]);
    assign outputs[9701] = (layer0_outputs[2349]) | (layer0_outputs[1359]);
    assign outputs[9702] = ~(layer0_outputs[9017]);
    assign outputs[9703] = ~(layer0_outputs[9996]);
    assign outputs[9704] = layer0_outputs[2190];
    assign outputs[9705] = ~((layer0_outputs[7592]) ^ (layer0_outputs[4475]));
    assign outputs[9706] = layer0_outputs[1657];
    assign outputs[9707] = ~((layer0_outputs[7102]) ^ (layer0_outputs[1264]));
    assign outputs[9708] = layer0_outputs[10029];
    assign outputs[9709] = layer0_outputs[2290];
    assign outputs[9710] = ~(layer0_outputs[4405]);
    assign outputs[9711] = (layer0_outputs[2221]) & ~(layer0_outputs[10097]);
    assign outputs[9712] = (layer0_outputs[1208]) ^ (layer0_outputs[7171]);
    assign outputs[9713] = ~((layer0_outputs[2484]) ^ (layer0_outputs[7769]));
    assign outputs[9714] = ~((layer0_outputs[3359]) ^ (layer0_outputs[9661]));
    assign outputs[9715] = (layer0_outputs[5819]) & ~(layer0_outputs[3002]);
    assign outputs[9716] = (layer0_outputs[5823]) | (layer0_outputs[5750]);
    assign outputs[9717] = ~(layer0_outputs[3725]);
    assign outputs[9718] = ~((layer0_outputs[2895]) | (layer0_outputs[1580]));
    assign outputs[9719] = layer0_outputs[5275];
    assign outputs[9720] = (layer0_outputs[4182]) ^ (layer0_outputs[1122]);
    assign outputs[9721] = (layer0_outputs[1183]) & (layer0_outputs[7937]);
    assign outputs[9722] = (layer0_outputs[6134]) & ~(layer0_outputs[9440]);
    assign outputs[9723] = layer0_outputs[8762];
    assign outputs[9724] = ~(layer0_outputs[2026]);
    assign outputs[9725] = (layer0_outputs[8382]) & (layer0_outputs[4692]);
    assign outputs[9726] = ~(layer0_outputs[1157]) | (layer0_outputs[830]);
    assign outputs[9727] = layer0_outputs[6842];
    assign outputs[9728] = (layer0_outputs[3270]) & (layer0_outputs[8875]);
    assign outputs[9729] = ~((layer0_outputs[10039]) | (layer0_outputs[9715]));
    assign outputs[9730] = (layer0_outputs[7436]) | (layer0_outputs[5046]);
    assign outputs[9731] = ~(layer0_outputs[3630]);
    assign outputs[9732] = ~(layer0_outputs[9358]);
    assign outputs[9733] = (layer0_outputs[1982]) & (layer0_outputs[6683]);
    assign outputs[9734] = (layer0_outputs[8414]) ^ (layer0_outputs[2957]);
    assign outputs[9735] = layer0_outputs[7933];
    assign outputs[9736] = (layer0_outputs[7494]) & (layer0_outputs[2659]);
    assign outputs[9737] = ~(layer0_outputs[270]);
    assign outputs[9738] = layer0_outputs[5139];
    assign outputs[9739] = ~((layer0_outputs[9999]) ^ (layer0_outputs[4519]));
    assign outputs[9740] = layer0_outputs[8597];
    assign outputs[9741] = ~(layer0_outputs[7883]);
    assign outputs[9742] = (layer0_outputs[7976]) | (layer0_outputs[8085]);
    assign outputs[9743] = layer0_outputs[1317];
    assign outputs[9744] = layer0_outputs[1301];
    assign outputs[9745] = (layer0_outputs[8401]) ^ (layer0_outputs[8026]);
    assign outputs[9746] = ~((layer0_outputs[7602]) ^ (layer0_outputs[2273]));
    assign outputs[9747] = layer0_outputs[9928];
    assign outputs[9748] = (layer0_outputs[1623]) & ~(layer0_outputs[7740]);
    assign outputs[9749] = layer0_outputs[7214];
    assign outputs[9750] = ~(layer0_outputs[3442]);
    assign outputs[9751] = ~((layer0_outputs[1084]) ^ (layer0_outputs[6729]));
    assign outputs[9752] = layer0_outputs[10020];
    assign outputs[9753] = layer0_outputs[1694];
    assign outputs[9754] = ~((layer0_outputs[4130]) | (layer0_outputs[3880]));
    assign outputs[9755] = layer0_outputs[2673];
    assign outputs[9756] = layer0_outputs[905];
    assign outputs[9757] = layer0_outputs[10078];
    assign outputs[9758] = layer0_outputs[5353];
    assign outputs[9759] = layer0_outputs[6697];
    assign outputs[9760] = ~(layer0_outputs[9551]);
    assign outputs[9761] = (layer0_outputs[5543]) ^ (layer0_outputs[887]);
    assign outputs[9762] = ~((layer0_outputs[8963]) ^ (layer0_outputs[5703]));
    assign outputs[9763] = (layer0_outputs[848]) ^ (layer0_outputs[5344]);
    assign outputs[9764] = ~((layer0_outputs[6710]) & (layer0_outputs[4810]));
    assign outputs[9765] = ~((layer0_outputs[3023]) ^ (layer0_outputs[8395]));
    assign outputs[9766] = ~(layer0_outputs[7325]);
    assign outputs[9767] = (layer0_outputs[1394]) ^ (layer0_outputs[7928]);
    assign outputs[9768] = ~(layer0_outputs[9856]);
    assign outputs[9769] = ~(layer0_outputs[7945]);
    assign outputs[9770] = (layer0_outputs[9516]) & (layer0_outputs[3400]);
    assign outputs[9771] = ~(layer0_outputs[9550]) | (layer0_outputs[3966]);
    assign outputs[9772] = ~((layer0_outputs[8037]) & (layer0_outputs[4997]));
    assign outputs[9773] = ~((layer0_outputs[6175]) ^ (layer0_outputs[1655]));
    assign outputs[9774] = (layer0_outputs[256]) ^ (layer0_outputs[3317]);
    assign outputs[9775] = ~(layer0_outputs[1523]);
    assign outputs[9776] = ~(layer0_outputs[1367]);
    assign outputs[9777] = layer0_outputs[1886];
    assign outputs[9778] = (layer0_outputs[7889]) & ~(layer0_outputs[4825]);
    assign outputs[9779] = (layer0_outputs[7411]) | (layer0_outputs[4179]);
    assign outputs[9780] = layer0_outputs[5587];
    assign outputs[9781] = ~(layer0_outputs[9220]);
    assign outputs[9782] = (layer0_outputs[1083]) ^ (layer0_outputs[8912]);
    assign outputs[9783] = (layer0_outputs[4173]) ^ (layer0_outputs[3105]);
    assign outputs[9784] = (layer0_outputs[1414]) & ~(layer0_outputs[2076]);
    assign outputs[9785] = layer0_outputs[9577];
    assign outputs[9786] = layer0_outputs[1126];
    assign outputs[9787] = layer0_outputs[7380];
    assign outputs[9788] = (layer0_outputs[1470]) & ~(layer0_outputs[9961]);
    assign outputs[9789] = layer0_outputs[6989];
    assign outputs[9790] = (layer0_outputs[2265]) ^ (layer0_outputs[9320]);
    assign outputs[9791] = ~((layer0_outputs[3141]) | (layer0_outputs[14]));
    assign outputs[9792] = (layer0_outputs[7148]) & ~(layer0_outputs[5409]);
    assign outputs[9793] = layer0_outputs[6516];
    assign outputs[9794] = layer0_outputs[1062];
    assign outputs[9795] = ~((layer0_outputs[4535]) | (layer0_outputs[7990]));
    assign outputs[9796] = layer0_outputs[9703];
    assign outputs[9797] = ~(layer0_outputs[5090]);
    assign outputs[9798] = ~((layer0_outputs[6159]) ^ (layer0_outputs[7674]));
    assign outputs[9799] = ~(layer0_outputs[1435]);
    assign outputs[9800] = layer0_outputs[7008];
    assign outputs[9801] = layer0_outputs[8968];
    assign outputs[9802] = layer0_outputs[7363];
    assign outputs[9803] = ~(layer0_outputs[2003]);
    assign outputs[9804] = (layer0_outputs[6831]) & ~(layer0_outputs[544]);
    assign outputs[9805] = (layer0_outputs[6642]) & ~(layer0_outputs[1978]);
    assign outputs[9806] = ~((layer0_outputs[653]) | (layer0_outputs[6865]));
    assign outputs[9807] = layer0_outputs[8033];
    assign outputs[9808] = layer0_outputs[6266];
    assign outputs[9809] = ~(layer0_outputs[9523]) | (layer0_outputs[3453]);
    assign outputs[9810] = ~(layer0_outputs[469]);
    assign outputs[9811] = ~(layer0_outputs[1092]);
    assign outputs[9812] = (layer0_outputs[7458]) & ~(layer0_outputs[2129]);
    assign outputs[9813] = (layer0_outputs[5081]) ^ (layer0_outputs[1858]);
    assign outputs[9814] = (layer0_outputs[9004]) ^ (layer0_outputs[8236]);
    assign outputs[9815] = layer0_outputs[5762];
    assign outputs[9816] = layer0_outputs[7343];
    assign outputs[9817] = (layer0_outputs[8202]) ^ (layer0_outputs[8429]);
    assign outputs[9818] = (layer0_outputs[9648]) & ~(layer0_outputs[5815]);
    assign outputs[9819] = layer0_outputs[5482];
    assign outputs[9820] = layer0_outputs[4210];
    assign outputs[9821] = (layer0_outputs[5284]) ^ (layer0_outputs[7136]);
    assign outputs[9822] = (layer0_outputs[332]) & ~(layer0_outputs[4097]);
    assign outputs[9823] = (layer0_outputs[7980]) & ~(layer0_outputs[10204]);
    assign outputs[9824] = (layer0_outputs[2546]) & ~(layer0_outputs[4964]);
    assign outputs[9825] = ~(layer0_outputs[6573]);
    assign outputs[9826] = layer0_outputs[8362];
    assign outputs[9827] = (layer0_outputs[1963]) & ~(layer0_outputs[5669]);
    assign outputs[9828] = ~((layer0_outputs[8686]) ^ (layer0_outputs[8933]));
    assign outputs[9829] = (layer0_outputs[539]) & ~(layer0_outputs[267]);
    assign outputs[9830] = ~(layer0_outputs[1295]);
    assign outputs[9831] = ~(layer0_outputs[2946]);
    assign outputs[9832] = (layer0_outputs[7123]) & ~(layer0_outputs[5975]);
    assign outputs[9833] = layer0_outputs[7995];
    assign outputs[9834] = ~((layer0_outputs[1986]) ^ (layer0_outputs[7281]));
    assign outputs[9835] = ~(layer0_outputs[4751]);
    assign outputs[9836] = layer0_outputs[7888];
    assign outputs[9837] = layer0_outputs[4310];
    assign outputs[9838] = ~(layer0_outputs[3790]);
    assign outputs[9839] = ~(layer0_outputs[2064]);
    assign outputs[9840] = (layer0_outputs[9824]) & ~(layer0_outputs[7713]);
    assign outputs[9841] = ~(layer0_outputs[5456]);
    assign outputs[9842] = ~(layer0_outputs[8920]);
    assign outputs[9843] = ~(layer0_outputs[625]);
    assign outputs[9844] = (layer0_outputs[1856]) & ~(layer0_outputs[4138]);
    assign outputs[9845] = layer0_outputs[5768];
    assign outputs[9846] = (layer0_outputs[9351]) ^ (layer0_outputs[5158]);
    assign outputs[9847] = ~((layer0_outputs[7080]) ^ (layer0_outputs[2682]));
    assign outputs[9848] = (layer0_outputs[132]) | (layer0_outputs[8900]);
    assign outputs[9849] = (layer0_outputs[419]) ^ (layer0_outputs[8482]);
    assign outputs[9850] = (layer0_outputs[860]) & (layer0_outputs[817]);
    assign outputs[9851] = ~(layer0_outputs[6651]);
    assign outputs[9852] = (layer0_outputs[7656]) | (layer0_outputs[899]);
    assign outputs[9853] = ~((layer0_outputs[6141]) ^ (layer0_outputs[3694]));
    assign outputs[9854] = layer0_outputs[2499];
    assign outputs[9855] = (layer0_outputs[7569]) & ~(layer0_outputs[5751]);
    assign outputs[9856] = ~(layer0_outputs[4571]);
    assign outputs[9857] = (layer0_outputs[338]) & ~(layer0_outputs[2014]);
    assign outputs[9858] = ~(layer0_outputs[153]);
    assign outputs[9859] = layer0_outputs[4552];
    assign outputs[9860] = (layer0_outputs[8647]) & (layer0_outputs[8334]);
    assign outputs[9861] = ~((layer0_outputs[5183]) | (layer0_outputs[1433]));
    assign outputs[9862] = ~(layer0_outputs[5921]);
    assign outputs[9863] = ~(layer0_outputs[7263]) | (layer0_outputs[1471]);
    assign outputs[9864] = (layer0_outputs[6003]) & ~(layer0_outputs[5956]);
    assign outputs[9865] = (layer0_outputs[8122]) ^ (layer0_outputs[6446]);
    assign outputs[9866] = ~(layer0_outputs[3134]);
    assign outputs[9867] = ~(layer0_outputs[9610]) | (layer0_outputs[5970]);
    assign outputs[9868] = ~(layer0_outputs[9669]);
    assign outputs[9869] = ~((layer0_outputs[8998]) & (layer0_outputs[1948]));
    assign outputs[9870] = ~((layer0_outputs[3187]) ^ (layer0_outputs[4019]));
    assign outputs[9871] = layer0_outputs[2809];
    assign outputs[9872] = ~(layer0_outputs[8460]);
    assign outputs[9873] = ~(layer0_outputs[858]);
    assign outputs[9874] = ~(layer0_outputs[793]);
    assign outputs[9875] = layer0_outputs[8125];
    assign outputs[9876] = layer0_outputs[4055];
    assign outputs[9877] = ~(layer0_outputs[10163]) | (layer0_outputs[8922]);
    assign outputs[9878] = ~((layer0_outputs[8346]) | (layer0_outputs[3563]));
    assign outputs[9879] = (layer0_outputs[7698]) ^ (layer0_outputs[1531]);
    assign outputs[9880] = ~(layer0_outputs[6237]);
    assign outputs[9881] = ~((layer0_outputs[7277]) & (layer0_outputs[636]));
    assign outputs[9882] = ~(layer0_outputs[4782]);
    assign outputs[9883] = ~((layer0_outputs[8657]) ^ (layer0_outputs[5376]));
    assign outputs[9884] = ~(layer0_outputs[729]);
    assign outputs[9885] = (layer0_outputs[5095]) & ~(layer0_outputs[7262]);
    assign outputs[9886] = ~(layer0_outputs[8512]);
    assign outputs[9887] = (layer0_outputs[2175]) & (layer0_outputs[4815]);
    assign outputs[9888] = ~(layer0_outputs[4386]);
    assign outputs[9889] = ~((layer0_outputs[1641]) ^ (layer0_outputs[5429]));
    assign outputs[9890] = layer0_outputs[9939];
    assign outputs[9891] = ~(layer0_outputs[8576]);
    assign outputs[9892] = ~((layer0_outputs[5207]) ^ (layer0_outputs[2135]));
    assign outputs[9893] = ~((layer0_outputs[10181]) ^ (layer0_outputs[3483]));
    assign outputs[9894] = (layer0_outputs[10103]) ^ (layer0_outputs[981]);
    assign outputs[9895] = 1'b0;
    assign outputs[9896] = ~((layer0_outputs[2850]) | (layer0_outputs[952]));
    assign outputs[9897] = ~((layer0_outputs[9001]) ^ (layer0_outputs[3721]));
    assign outputs[9898] = ~((layer0_outputs[1954]) ^ (layer0_outputs[9472]));
    assign outputs[9899] = (layer0_outputs[2377]) & ~(layer0_outputs[7905]);
    assign outputs[9900] = ~((layer0_outputs[358]) | (layer0_outputs[1990]));
    assign outputs[9901] = (layer0_outputs[3828]) & ~(layer0_outputs[4047]);
    assign outputs[9902] = ~(layer0_outputs[7925]);
    assign outputs[9903] = layer0_outputs[5309];
    assign outputs[9904] = layer0_outputs[5552];
    assign outputs[9905] = ~(layer0_outputs[2628]);
    assign outputs[9906] = ~(layer0_outputs[3969]);
    assign outputs[9907] = ~(layer0_outputs[7887]);
    assign outputs[9908] = layer0_outputs[2052];
    assign outputs[9909] = ~(layer0_outputs[4354]);
    assign outputs[9910] = ~((layer0_outputs[9866]) | (layer0_outputs[5411]));
    assign outputs[9911] = layer0_outputs[4565];
    assign outputs[9912] = layer0_outputs[10197];
    assign outputs[9913] = (layer0_outputs[9822]) & (layer0_outputs[3195]);
    assign outputs[9914] = (layer0_outputs[1541]) & ~(layer0_outputs[201]);
    assign outputs[9915] = (layer0_outputs[6884]) ^ (layer0_outputs[623]);
    assign outputs[9916] = ~((layer0_outputs[1389]) | (layer0_outputs[6417]));
    assign outputs[9917] = ~((layer0_outputs[7609]) ^ (layer0_outputs[3553]));
    assign outputs[9918] = (layer0_outputs[9561]) & ~(layer0_outputs[1304]);
    assign outputs[9919] = ~((layer0_outputs[9538]) | (layer0_outputs[7659]));
    assign outputs[9920] = layer0_outputs[6524];
    assign outputs[9921] = layer0_outputs[7663];
    assign outputs[9922] = ~((layer0_outputs[3343]) & (layer0_outputs[9657]));
    assign outputs[9923] = (layer0_outputs[257]) ^ (layer0_outputs[10147]);
    assign outputs[9924] = ~(layer0_outputs[5979]);
    assign outputs[9925] = ~((layer0_outputs[2006]) ^ (layer0_outputs[5545]));
    assign outputs[9926] = ~(layer0_outputs[7260]);
    assign outputs[9927] = ~(layer0_outputs[2615]);
    assign outputs[9928] = ~(layer0_outputs[767]);
    assign outputs[9929] = layer0_outputs[1916];
    assign outputs[9930] = ~((layer0_outputs[26]) ^ (layer0_outputs[384]));
    assign outputs[9931] = ~(layer0_outputs[2624]);
    assign outputs[9932] = ~((layer0_outputs[9969]) & (layer0_outputs[2655]));
    assign outputs[9933] = layer0_outputs[9162];
    assign outputs[9934] = (layer0_outputs[10165]) & ~(layer0_outputs[754]);
    assign outputs[9935] = ~(layer0_outputs[8978]);
    assign outputs[9936] = (layer0_outputs[9613]) & (layer0_outputs[1145]);
    assign outputs[9937] = ~(layer0_outputs[4204]);
    assign outputs[9938] = (layer0_outputs[2818]) & ~(layer0_outputs[2113]);
    assign outputs[9939] = ~((layer0_outputs[8918]) ^ (layer0_outputs[8325]));
    assign outputs[9940] = ~(layer0_outputs[40]);
    assign outputs[9941] = (layer0_outputs[2677]) ^ (layer0_outputs[1960]);
    assign outputs[9942] = (layer0_outputs[8945]) ^ (layer0_outputs[9338]);
    assign outputs[9943] = layer0_outputs[1644];
    assign outputs[9944] = ~((layer0_outputs[4588]) ^ (layer0_outputs[6339]));
    assign outputs[9945] = ~(layer0_outputs[2352]);
    assign outputs[9946] = layer0_outputs[9647];
    assign outputs[9947] = ~(layer0_outputs[8845]);
    assign outputs[9948] = (layer0_outputs[9987]) & ~(layer0_outputs[7630]);
    assign outputs[9949] = (layer0_outputs[4774]) & ~(layer0_outputs[66]);
    assign outputs[9950] = ~((layer0_outputs[7053]) | (layer0_outputs[9247]));
    assign outputs[9951] = ~((layer0_outputs[3795]) ^ (layer0_outputs[3004]));
    assign outputs[9952] = ~((layer0_outputs[2461]) ^ (layer0_outputs[6685]));
    assign outputs[9953] = layer0_outputs[4837];
    assign outputs[9954] = ~((layer0_outputs[5148]) ^ (layer0_outputs[9321]));
    assign outputs[9955] = layer0_outputs[1307];
    assign outputs[9956] = ~(layer0_outputs[3903]);
    assign outputs[9957] = ~(layer0_outputs[7243]);
    assign outputs[9958] = (layer0_outputs[2259]) ^ (layer0_outputs[5210]);
    assign outputs[9959] = (layer0_outputs[3597]) & ~(layer0_outputs[6973]);
    assign outputs[9960] = ~((layer0_outputs[9524]) ^ (layer0_outputs[3083]));
    assign outputs[9961] = (layer0_outputs[2055]) | (layer0_outputs[3429]);
    assign outputs[9962] = (layer0_outputs[4100]) & ~(layer0_outputs[7860]);
    assign outputs[9963] = (layer0_outputs[9811]) | (layer0_outputs[5940]);
    assign outputs[9964] = (layer0_outputs[7245]) ^ (layer0_outputs[6609]);
    assign outputs[9965] = ~(layer0_outputs[3217]);
    assign outputs[9966] = ~(layer0_outputs[2330]);
    assign outputs[9967] = ~((layer0_outputs[9637]) ^ (layer0_outputs[4940]));
    assign outputs[9968] = (layer0_outputs[6563]) & ~(layer0_outputs[7800]);
    assign outputs[9969] = ~(layer0_outputs[3875]);
    assign outputs[9970] = layer0_outputs[7101];
    assign outputs[9971] = layer0_outputs[9701];
    assign outputs[9972] = ~(layer0_outputs[7451]);
    assign outputs[9973] = (layer0_outputs[2410]) & ~(layer0_outputs[9293]);
    assign outputs[9974] = (layer0_outputs[1812]) & (layer0_outputs[6887]);
    assign outputs[9975] = ~(layer0_outputs[9346]);
    assign outputs[9976] = layer0_outputs[2890];
    assign outputs[9977] = layer0_outputs[1251];
    assign outputs[9978] = ~((layer0_outputs[1443]) ^ (layer0_outputs[1043]));
    assign outputs[9979] = ~(layer0_outputs[8662]);
    assign outputs[9980] = ~(layer0_outputs[7084]);
    assign outputs[9981] = (layer0_outputs[4979]) ^ (layer0_outputs[1332]);
    assign outputs[9982] = ~(layer0_outputs[2891]) | (layer0_outputs[6751]);
    assign outputs[9983] = (layer0_outputs[8560]) & ~(layer0_outputs[6777]);
    assign outputs[9984] = ~(layer0_outputs[9993]);
    assign outputs[9985] = ~((layer0_outputs[4842]) ^ (layer0_outputs[3007]));
    assign outputs[9986] = (layer0_outputs[2867]) ^ (layer0_outputs[5567]);
    assign outputs[9987] = (layer0_outputs[3678]) & ~(layer0_outputs[1339]);
    assign outputs[9988] = ~((layer0_outputs[5072]) | (layer0_outputs[2038]));
    assign outputs[9989] = layer0_outputs[9855];
    assign outputs[9990] = ~(layer0_outputs[5529]);
    assign outputs[9991] = ~(layer0_outputs[8358]);
    assign outputs[9992] = (layer0_outputs[7933]) & ~(layer0_outputs[4980]);
    assign outputs[9993] = layer0_outputs[3412];
    assign outputs[9994] = ~(layer0_outputs[4591]);
    assign outputs[9995] = layer0_outputs[10195];
    assign outputs[9996] = layer0_outputs[998];
    assign outputs[9997] = ~((layer0_outputs[8138]) ^ (layer0_outputs[3261]));
    assign outputs[9998] = (layer0_outputs[9404]) ^ (layer0_outputs[1236]);
    assign outputs[9999] = layer0_outputs[7654];
    assign outputs[10000] = ~(layer0_outputs[1497]) | (layer0_outputs[416]);
    assign outputs[10001] = ~(layer0_outputs[2913]);
    assign outputs[10002] = ~(layer0_outputs[7981]);
    assign outputs[10003] = (layer0_outputs[4195]) & ~(layer0_outputs[5896]);
    assign outputs[10004] = ~(layer0_outputs[8929]);
    assign outputs[10005] = ~(layer0_outputs[9529]) | (layer0_outputs[5006]);
    assign outputs[10006] = (layer0_outputs[661]) & ~(layer0_outputs[6854]);
    assign outputs[10007] = ~(layer0_outputs[2674]) | (layer0_outputs[1833]);
    assign outputs[10008] = ~((layer0_outputs[9931]) ^ (layer0_outputs[8689]));
    assign outputs[10009] = ~(layer0_outputs[2364]);
    assign outputs[10010] = ~(layer0_outputs[5212]);
    assign outputs[10011] = (layer0_outputs[196]) & ~(layer0_outputs[5633]);
    assign outputs[10012] = layer0_outputs[3593];
    assign outputs[10013] = layer0_outputs[6976];
    assign outputs[10014] = ~(layer0_outputs[4237]);
    assign outputs[10015] = layer0_outputs[3967];
    assign outputs[10016] = ~((layer0_outputs[6945]) & (layer0_outputs[1894]));
    assign outputs[10017] = ~(layer0_outputs[1086]);
    assign outputs[10018] = layer0_outputs[9926];
    assign outputs[10019] = ~(layer0_outputs[4694]);
    assign outputs[10020] = (layer0_outputs[4436]) & ~(layer0_outputs[3419]);
    assign outputs[10021] = (layer0_outputs[8098]) ^ (layer0_outputs[9359]);
    assign outputs[10022] = (layer0_outputs[9202]) & ~(layer0_outputs[6878]);
    assign outputs[10023] = ~((layer0_outputs[2066]) ^ (layer0_outputs[6833]));
    assign outputs[10024] = ~(layer0_outputs[7496]);
    assign outputs[10025] = ~(layer0_outputs[2158]);
    assign outputs[10026] = layer0_outputs[6671];
    assign outputs[10027] = layer0_outputs[1456];
    assign outputs[10028] = (layer0_outputs[6007]) | (layer0_outputs[2803]);
    assign outputs[10029] = (layer0_outputs[2393]) & ~(layer0_outputs[2392]);
    assign outputs[10030] = ~(layer0_outputs[3062]);
    assign outputs[10031] = (layer0_outputs[2918]) ^ (layer0_outputs[130]);
    assign outputs[10032] = layer0_outputs[9339];
    assign outputs[10033] = layer0_outputs[5501];
    assign outputs[10034] = (layer0_outputs[744]) ^ (layer0_outputs[9994]);
    assign outputs[10035] = ~((layer0_outputs[6538]) ^ (layer0_outputs[5633]));
    assign outputs[10036] = (layer0_outputs[6095]) ^ (layer0_outputs[7820]);
    assign outputs[10037] = (layer0_outputs[5900]) & ~(layer0_outputs[4095]);
    assign outputs[10038] = (layer0_outputs[3294]) & (layer0_outputs[5892]);
    assign outputs[10039] = (layer0_outputs[868]) ^ (layer0_outputs[9034]);
    assign outputs[10040] = ~((layer0_outputs[8912]) ^ (layer0_outputs[1664]));
    assign outputs[10041] = (layer0_outputs[3555]) & ~(layer0_outputs[5219]);
    assign outputs[10042] = ~((layer0_outputs[1421]) | (layer0_outputs[8000]));
    assign outputs[10043] = layer0_outputs[4856];
    assign outputs[10044] = ~(layer0_outputs[1872]);
    assign outputs[10045] = (layer0_outputs[6381]) ^ (layer0_outputs[4603]);
    assign outputs[10046] = layer0_outputs[3024];
    assign outputs[10047] = layer0_outputs[9822];
    assign outputs[10048] = ~(layer0_outputs[5078]);
    assign outputs[10049] = (layer0_outputs[3431]) & ~(layer0_outputs[7187]);
    assign outputs[10050] = layer0_outputs[8627];
    assign outputs[10051] = (layer0_outputs[7157]) | (layer0_outputs[9965]);
    assign outputs[10052] = ~(layer0_outputs[8520]);
    assign outputs[10053] = (layer0_outputs[2072]) & ~(layer0_outputs[10222]);
    assign outputs[10054] = ~(layer0_outputs[7406]);
    assign outputs[10055] = (layer0_outputs[1300]) & ~(layer0_outputs[3643]);
    assign outputs[10056] = ~(layer0_outputs[3097]);
    assign outputs[10057] = layer0_outputs[6988];
    assign outputs[10058] = ~((layer0_outputs[8466]) ^ (layer0_outputs[7060]));
    assign outputs[10059] = (layer0_outputs[2152]) ^ (layer0_outputs[5575]);
    assign outputs[10060] = (layer0_outputs[6089]) ^ (layer0_outputs[1648]);
    assign outputs[10061] = (layer0_outputs[5195]) & ~(layer0_outputs[3737]);
    assign outputs[10062] = ~(layer0_outputs[9903]);
    assign outputs[10063] = ~(layer0_outputs[4654]);
    assign outputs[10064] = (layer0_outputs[5620]) | (layer0_outputs[6035]);
    assign outputs[10065] = (layer0_outputs[6981]) & ~(layer0_outputs[1142]);
    assign outputs[10066] = ~(layer0_outputs[2156]) | (layer0_outputs[4146]);
    assign outputs[10067] = (layer0_outputs[4178]) & ~(layer0_outputs[8469]);
    assign outputs[10068] = ~(layer0_outputs[10068]);
    assign outputs[10069] = (layer0_outputs[3381]) ^ (layer0_outputs[7044]);
    assign outputs[10070] = layer0_outputs[102];
    assign outputs[10071] = layer0_outputs[731];
    assign outputs[10072] = ~(layer0_outputs[8215]);
    assign outputs[10073] = ~((layer0_outputs[784]) ^ (layer0_outputs[7145]));
    assign outputs[10074] = ~((layer0_outputs[2127]) ^ (layer0_outputs[1007]));
    assign outputs[10075] = (layer0_outputs[8571]) & (layer0_outputs[4054]);
    assign outputs[10076] = ~((layer0_outputs[5838]) | (layer0_outputs[4923]));
    assign outputs[10077] = ~(layer0_outputs[5887]);
    assign outputs[10078] = layer0_outputs[5374];
    assign outputs[10079] = ~(layer0_outputs[8673]);
    assign outputs[10080] = ~(layer0_outputs[4175]) | (layer0_outputs[1273]);
    assign outputs[10081] = ~(layer0_outputs[9589]);
    assign outputs[10082] = ~((layer0_outputs[2909]) ^ (layer0_outputs[6226]));
    assign outputs[10083] = ~(layer0_outputs[3768]);
    assign outputs[10084] = layer0_outputs[8516];
    assign outputs[10085] = ~(layer0_outputs[1193]);
    assign outputs[10086] = (layer0_outputs[8633]) & ~(layer0_outputs[1595]);
    assign outputs[10087] = (layer0_outputs[7177]) & ~(layer0_outputs[5469]);
    assign outputs[10088] = ~(layer0_outputs[1280]) | (layer0_outputs[2469]);
    assign outputs[10089] = layer0_outputs[4681];
    assign outputs[10090] = layer0_outputs[1250];
    assign outputs[10091] = (layer0_outputs[446]) & (layer0_outputs[5172]);
    assign outputs[10092] = ~(layer0_outputs[7783]);
    assign outputs[10093] = (layer0_outputs[8061]) ^ (layer0_outputs[6606]);
    assign outputs[10094] = ~(layer0_outputs[8192]);
    assign outputs[10095] = layer0_outputs[5244];
    assign outputs[10096] = ~((layer0_outputs[7344]) | (layer0_outputs[614]));
    assign outputs[10097] = (layer0_outputs[2424]) & ~(layer0_outputs[6172]);
    assign outputs[10098] = layer0_outputs[9137];
    assign outputs[10099] = ~((layer0_outputs[9381]) ^ (layer0_outputs[637]));
    assign outputs[10100] = layer0_outputs[6600];
    assign outputs[10101] = ~(layer0_outputs[4726]);
    assign outputs[10102] = ~(layer0_outputs[1231]);
    assign outputs[10103] = ~((layer0_outputs[5983]) | (layer0_outputs[8639]));
    assign outputs[10104] = layer0_outputs[7193];
    assign outputs[10105] = ~(layer0_outputs[2730]) | (layer0_outputs[7331]);
    assign outputs[10106] = layer0_outputs[1748];
    assign outputs[10107] = ~(layer0_outputs[7646]);
    assign outputs[10108] = layer0_outputs[2277];
    assign outputs[10109] = (layer0_outputs[7453]) & ~(layer0_outputs[8432]);
    assign outputs[10110] = (layer0_outputs[1234]) & ~(layer0_outputs[8105]);
    assign outputs[10111] = layer0_outputs[1141];
    assign outputs[10112] = (layer0_outputs[857]) & ~(layer0_outputs[10147]);
    assign outputs[10113] = layer0_outputs[2873];
    assign outputs[10114] = layer0_outputs[8514];
    assign outputs[10115] = layer0_outputs[1924];
    assign outputs[10116] = ~(layer0_outputs[4770]);
    assign outputs[10117] = layer0_outputs[3454];
    assign outputs[10118] = ~(layer0_outputs[8952]);
    assign outputs[10119] = ~((layer0_outputs[5184]) | (layer0_outputs[3291]));
    assign outputs[10120] = (layer0_outputs[2605]) ^ (layer0_outputs[6761]);
    assign outputs[10121] = layer0_outputs[28];
    assign outputs[10122] = ~((layer0_outputs[5767]) ^ (layer0_outputs[1546]));
    assign outputs[10123] = layer0_outputs[7297];
    assign outputs[10124] = ~(layer0_outputs[1855]) | (layer0_outputs[254]);
    assign outputs[10125] = (layer0_outputs[4830]) & (layer0_outputs[8085]);
    assign outputs[10126] = ~((layer0_outputs[7597]) | (layer0_outputs[4213]));
    assign outputs[10127] = ~(layer0_outputs[386]);
    assign outputs[10128] = ~((layer0_outputs[3159]) ^ (layer0_outputs[8470]));
    assign outputs[10129] = ~((layer0_outputs[3805]) ^ (layer0_outputs[8843]));
    assign outputs[10130] = layer0_outputs[8944];
    assign outputs[10131] = layer0_outputs[9054];
    assign outputs[10132] = (layer0_outputs[4871]) & ~(layer0_outputs[5556]);
    assign outputs[10133] = ~(layer0_outputs[501]);
    assign outputs[10134] = (layer0_outputs[5748]) ^ (layer0_outputs[9757]);
    assign outputs[10135] = layer0_outputs[6621];
    assign outputs[10136] = (layer0_outputs[10238]) ^ (layer0_outputs[8791]);
    assign outputs[10137] = layer0_outputs[4240];
    assign outputs[10138] = layer0_outputs[8864];
    assign outputs[10139] = layer0_outputs[8649];
    assign outputs[10140] = ~(layer0_outputs[2138]);
    assign outputs[10141] = ~(layer0_outputs[3781]);
    assign outputs[10142] = ~(layer0_outputs[5367]);
    assign outputs[10143] = ~(layer0_outputs[2387]);
    assign outputs[10144] = ~(layer0_outputs[7178]);
    assign outputs[10145] = layer0_outputs[1470];
    assign outputs[10146] = ~(layer0_outputs[5218]) | (layer0_outputs[1683]);
    assign outputs[10147] = ~(layer0_outputs[4128]) | (layer0_outputs[3113]);
    assign outputs[10148] = (layer0_outputs[3268]) & ~(layer0_outputs[1397]);
    assign outputs[10149] = ~((layer0_outputs[8811]) | (layer0_outputs[9254]));
    assign outputs[10150] = ~(layer0_outputs[4193]);
    assign outputs[10151] = layer0_outputs[2706];
    assign outputs[10152] = (layer0_outputs[5852]) | (layer0_outputs[6754]);
    assign outputs[10153] = layer0_outputs[7558];
    assign outputs[10154] = ~(layer0_outputs[8684]);
    assign outputs[10155] = ~((layer0_outputs[9777]) ^ (layer0_outputs[10093]));
    assign outputs[10156] = ~(layer0_outputs[99]) | (layer0_outputs[1857]);
    assign outputs[10157] = layer0_outputs[5907];
    assign outputs[10158] = ~(layer0_outputs[2505]);
    assign outputs[10159] = ~(layer0_outputs[9998]);
    assign outputs[10160] = ~(layer0_outputs[2521]) | (layer0_outputs[5019]);
    assign outputs[10161] = ~((layer0_outputs[1605]) & (layer0_outputs[597]));
    assign outputs[10162] = layer0_outputs[8366];
    assign outputs[10163] = ~((layer0_outputs[5285]) | (layer0_outputs[7764]));
    assign outputs[10164] = (layer0_outputs[7475]) & (layer0_outputs[3423]);
    assign outputs[10165] = (layer0_outputs[684]) & ~(layer0_outputs[1373]);
    assign outputs[10166] = ~(layer0_outputs[6022]);
    assign outputs[10167] = layer0_outputs[850];
    assign outputs[10168] = layer0_outputs[5846];
    assign outputs[10169] = ~((layer0_outputs[4361]) ^ (layer0_outputs[9318]));
    assign outputs[10170] = layer0_outputs[5150];
    assign outputs[10171] = ~((layer0_outputs[563]) ^ (layer0_outputs[7825]));
    assign outputs[10172] = (layer0_outputs[9790]) ^ (layer0_outputs[765]);
    assign outputs[10173] = (layer0_outputs[3669]) ^ (layer0_outputs[175]);
    assign outputs[10174] = ~(layer0_outputs[22]);
    assign outputs[10175] = (layer0_outputs[8862]) ^ (layer0_outputs[4648]);
    assign outputs[10176] = ~(layer0_outputs[7138]);
    assign outputs[10177] = ~((layer0_outputs[1320]) | (layer0_outputs[8022]));
    assign outputs[10178] = ~(layer0_outputs[9236]) | (layer0_outputs[1792]);
    assign outputs[10179] = (layer0_outputs[1574]) ^ (layer0_outputs[7481]);
    assign outputs[10180] = (layer0_outputs[3641]) & (layer0_outputs[2322]);
    assign outputs[10181] = ~(layer0_outputs[9766]) | (layer0_outputs[4715]);
    assign outputs[10182] = (layer0_outputs[5990]) & ~(layer0_outputs[8701]);
    assign outputs[10183] = (layer0_outputs[4677]) ^ (layer0_outputs[1975]);
    assign outputs[10184] = (layer0_outputs[4459]) ^ (layer0_outputs[8391]);
    assign outputs[10185] = layer0_outputs[4931];
    assign outputs[10186] = layer0_outputs[7894];
    assign outputs[10187] = ~(layer0_outputs[7700]);
    assign outputs[10188] = (layer0_outputs[2765]) & (layer0_outputs[8438]);
    assign outputs[10189] = (layer0_outputs[8837]) & ~(layer0_outputs[4916]);
    assign outputs[10190] = ~((layer0_outputs[9788]) ^ (layer0_outputs[7308]));
    assign outputs[10191] = ~((layer0_outputs[2283]) & (layer0_outputs[3030]));
    assign outputs[10192] = (layer0_outputs[2154]) ^ (layer0_outputs[2470]);
    assign outputs[10193] = ~(layer0_outputs[6216]) | (layer0_outputs[3354]);
    assign outputs[10194] = ~((layer0_outputs[4292]) ^ (layer0_outputs[4704]));
    assign outputs[10195] = layer0_outputs[3932];
    assign outputs[10196] = layer0_outputs[62];
    assign outputs[10197] = ~((layer0_outputs[3105]) ^ (layer0_outputs[2195]));
    assign outputs[10198] = (layer0_outputs[9169]) & ~(layer0_outputs[1177]);
    assign outputs[10199] = ~((layer0_outputs[8405]) & (layer0_outputs[6246]));
    assign outputs[10200] = (layer0_outputs[2715]) ^ (layer0_outputs[8557]);
    assign outputs[10201] = (layer0_outputs[10106]) & ~(layer0_outputs[2915]);
    assign outputs[10202] = (layer0_outputs[8073]) & ~(layer0_outputs[2798]);
    assign outputs[10203] = ~(layer0_outputs[9843]);
    assign outputs[10204] = (layer0_outputs[2187]) & ~(layer0_outputs[574]);
    assign outputs[10205] = (layer0_outputs[5619]) & (layer0_outputs[695]);
    assign outputs[10206] = (layer0_outputs[8655]) & (layer0_outputs[4518]);
    assign outputs[10207] = layer0_outputs[2084];
    assign outputs[10208] = layer0_outputs[3408];
    assign outputs[10209] = (layer0_outputs[463]) & ~(layer0_outputs[5939]);
    assign outputs[10210] = (layer0_outputs[6862]) ^ (layer0_outputs[6448]);
    assign outputs[10211] = (layer0_outputs[5955]) ^ (layer0_outputs[3994]);
    assign outputs[10212] = ~(layer0_outputs[8852]);
    assign outputs[10213] = (layer0_outputs[5341]) & ~(layer0_outputs[1285]);
    assign outputs[10214] = ~((layer0_outputs[5228]) ^ (layer0_outputs[9339]));
    assign outputs[10215] = ~(layer0_outputs[4908]);
    assign outputs[10216] = ~((layer0_outputs[9947]) ^ (layer0_outputs[2437]));
    assign outputs[10217] = layer0_outputs[1483];
    assign outputs[10218] = ~((layer0_outputs[6170]) | (layer0_outputs[2770]));
    assign outputs[10219] = (layer0_outputs[3573]) & (layer0_outputs[1]);
    assign outputs[10220] = layer0_outputs[987];
    assign outputs[10221] = ~(layer0_outputs[10208]);
    assign outputs[10222] = ~(layer0_outputs[127]);
    assign outputs[10223] = ~((layer0_outputs[1097]) ^ (layer0_outputs[2829]));
    assign outputs[10224] = ~((layer0_outputs[1948]) ^ (layer0_outputs[4673]));
    assign outputs[10225] = ~(layer0_outputs[7362]);
    assign outputs[10226] = ~(layer0_outputs[8335]);
    assign outputs[10227] = (layer0_outputs[6425]) | (layer0_outputs[6521]);
    assign outputs[10228] = (layer0_outputs[3446]) ^ (layer0_outputs[6715]);
    assign outputs[10229] = (layer0_outputs[8123]) & ~(layer0_outputs[5709]);
    assign outputs[10230] = ~((layer0_outputs[8108]) ^ (layer0_outputs[2260]));
    assign outputs[10231] = (layer0_outputs[2086]) & (layer0_outputs[7819]);
    assign outputs[10232] = ~((layer0_outputs[8829]) ^ (layer0_outputs[2999]));
    assign outputs[10233] = layer0_outputs[2215];
    assign outputs[10234] = ~((layer0_outputs[7577]) ^ (layer0_outputs[9919]));
    assign outputs[10235] = (layer0_outputs[5641]) & ~(layer0_outputs[5404]);
    assign outputs[10236] = ~(layer0_outputs[3100]);
    assign outputs[10237] = ~((layer0_outputs[2570]) | (layer0_outputs[7257]));
    assign outputs[10238] = layer0_outputs[2288];
    assign outputs[10239] = ~(layer0_outputs[4446]);
endmodule
