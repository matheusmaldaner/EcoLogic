library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(5119 downto 0);
    signal layer1_outputs: std_logic_vector(5119 downto 0);
    signal layer2_outputs: std_logic_vector(5119 downto 0);

begin
    layer0_outputs(0) <= not (a or b);
    layer0_outputs(1) <= a or b;
    layer0_outputs(2) <= not (a or b);
    layer0_outputs(3) <= a or b;
    layer0_outputs(4) <= a and b;
    layer0_outputs(5) <= b and not a;
    layer0_outputs(6) <= b and not a;
    layer0_outputs(7) <= a and not b;
    layer0_outputs(8) <= b and not a;
    layer0_outputs(9) <= not b;
    layer0_outputs(10) <= a xor b;
    layer0_outputs(11) <= a or b;
    layer0_outputs(12) <= a or b;
    layer0_outputs(13) <= b;
    layer0_outputs(14) <= a or b;
    layer0_outputs(15) <= not (a xor b);
    layer0_outputs(16) <= 1'b0;
    layer0_outputs(17) <= not a or b;
    layer0_outputs(18) <= not (a or b);
    layer0_outputs(19) <= a;
    layer0_outputs(20) <= not (a xor b);
    layer0_outputs(21) <= a xor b;
    layer0_outputs(22) <= not a or b;
    layer0_outputs(23) <= not a;
    layer0_outputs(24) <= a xor b;
    layer0_outputs(25) <= 1'b1;
    layer0_outputs(26) <= not b or a;
    layer0_outputs(27) <= not a;
    layer0_outputs(28) <= not b;
    layer0_outputs(29) <= a and not b;
    layer0_outputs(30) <= not (a or b);
    layer0_outputs(31) <= not a;
    layer0_outputs(32) <= not (a xor b);
    layer0_outputs(33) <= a;
    layer0_outputs(34) <= a or b;
    layer0_outputs(35) <= not (a xor b);
    layer0_outputs(36) <= not (a or b);
    layer0_outputs(37) <= 1'b1;
    layer0_outputs(38) <= a and not b;
    layer0_outputs(39) <= not b;
    layer0_outputs(40) <= not b;
    layer0_outputs(41) <= a xor b;
    layer0_outputs(42) <= a;
    layer0_outputs(43) <= not (a xor b);
    layer0_outputs(44) <= not (a or b);
    layer0_outputs(45) <= a or b;
    layer0_outputs(46) <= a or b;
    layer0_outputs(47) <= a or b;
    layer0_outputs(48) <= b;
    layer0_outputs(49) <= a and not b;
    layer0_outputs(50) <= not (a xor b);
    layer0_outputs(51) <= not b or a;
    layer0_outputs(52) <= not b;
    layer0_outputs(53) <= a xor b;
    layer0_outputs(54) <= not b;
    layer0_outputs(55) <= not a or b;
    layer0_outputs(56) <= not b or a;
    layer0_outputs(57) <= not a;
    layer0_outputs(58) <= b and not a;
    layer0_outputs(59) <= b and not a;
    layer0_outputs(60) <= a and not b;
    layer0_outputs(61) <= a or b;
    layer0_outputs(62) <= b and not a;
    layer0_outputs(63) <= not (a xor b);
    layer0_outputs(64) <= not a;
    layer0_outputs(65) <= not (a and b);
    layer0_outputs(66) <= not (a or b);
    layer0_outputs(67) <= not a;
    layer0_outputs(68) <= not b;
    layer0_outputs(69) <= a;
    layer0_outputs(70) <= not b;
    layer0_outputs(71) <= not (a or b);
    layer0_outputs(72) <= not (a or b);
    layer0_outputs(73) <= a or b;
    layer0_outputs(74) <= not (a and b);
    layer0_outputs(75) <= a;
    layer0_outputs(76) <= not (a or b);
    layer0_outputs(77) <= not (a or b);
    layer0_outputs(78) <= not (a or b);
    layer0_outputs(79) <= a xor b;
    layer0_outputs(80) <= b;
    layer0_outputs(81) <= a or b;
    layer0_outputs(82) <= not (a xor b);
    layer0_outputs(83) <= b and not a;
    layer0_outputs(84) <= a or b;
    layer0_outputs(85) <= b and not a;
    layer0_outputs(86) <= 1'b1;
    layer0_outputs(87) <= b and not a;
    layer0_outputs(88) <= a and not b;
    layer0_outputs(89) <= a or b;
    layer0_outputs(90) <= a and not b;
    layer0_outputs(91) <= a or b;
    layer0_outputs(92) <= b and not a;
    layer0_outputs(93) <= b;
    layer0_outputs(94) <= not (a xor b);
    layer0_outputs(95) <= a;
    layer0_outputs(96) <= b;
    layer0_outputs(97) <= not a or b;
    layer0_outputs(98) <= not b or a;
    layer0_outputs(99) <= not (a or b);
    layer0_outputs(100) <= a;
    layer0_outputs(101) <= not (a xor b);
    layer0_outputs(102) <= b and not a;
    layer0_outputs(103) <= a xor b;
    layer0_outputs(104) <= a or b;
    layer0_outputs(105) <= not (a or b);
    layer0_outputs(106) <= not a;
    layer0_outputs(107) <= not b;
    layer0_outputs(108) <= not b or a;
    layer0_outputs(109) <= 1'b1;
    layer0_outputs(110) <= a xor b;
    layer0_outputs(111) <= a and not b;
    layer0_outputs(112) <= a;
    layer0_outputs(113) <= not b or a;
    layer0_outputs(114) <= not a;
    layer0_outputs(115) <= a or b;
    layer0_outputs(116) <= a xor b;
    layer0_outputs(117) <= a or b;
    layer0_outputs(118) <= not a or b;
    layer0_outputs(119) <= a;
    layer0_outputs(120) <= not (a or b);
    layer0_outputs(121) <= a or b;
    layer0_outputs(122) <= not (a or b);
    layer0_outputs(123) <= a and not b;
    layer0_outputs(124) <= b and not a;
    layer0_outputs(125) <= not a;
    layer0_outputs(126) <= a and not b;
    layer0_outputs(127) <= a or b;
    layer0_outputs(128) <= a;
    layer0_outputs(129) <= not (a xor b);
    layer0_outputs(130) <= 1'b1;
    layer0_outputs(131) <= not a or b;
    layer0_outputs(132) <= not b or a;
    layer0_outputs(133) <= a and b;
    layer0_outputs(134) <= not b or a;
    layer0_outputs(135) <= 1'b1;
    layer0_outputs(136) <= a;
    layer0_outputs(137) <= not (a or b);
    layer0_outputs(138) <= a;
    layer0_outputs(139) <= not a;
    layer0_outputs(140) <= not b;
    layer0_outputs(141) <= a;
    layer0_outputs(142) <= not b or a;
    layer0_outputs(143) <= not (a or b);
    layer0_outputs(144) <= not (a xor b);
    layer0_outputs(145) <= a;
    layer0_outputs(146) <= a xor b;
    layer0_outputs(147) <= a and not b;
    layer0_outputs(148) <= a;
    layer0_outputs(149) <= 1'b0;
    layer0_outputs(150) <= a or b;
    layer0_outputs(151) <= not (a or b);
    layer0_outputs(152) <= not a;
    layer0_outputs(153) <= 1'b1;
    layer0_outputs(154) <= not b;
    layer0_outputs(155) <= not a or b;
    layer0_outputs(156) <= not a;
    layer0_outputs(157) <= not (a xor b);
    layer0_outputs(158) <= a xor b;
    layer0_outputs(159) <= not b or a;
    layer0_outputs(160) <= not (a and b);
    layer0_outputs(161) <= b and not a;
    layer0_outputs(162) <= b;
    layer0_outputs(163) <= not (a or b);
    layer0_outputs(164) <= not (a or b);
    layer0_outputs(165) <= a xor b;
    layer0_outputs(166) <= not a;
    layer0_outputs(167) <= 1'b0;
    layer0_outputs(168) <= not (a xor b);
    layer0_outputs(169) <= b and not a;
    layer0_outputs(170) <= a or b;
    layer0_outputs(171) <= not (a or b);
    layer0_outputs(172) <= not b or a;
    layer0_outputs(173) <= not (a xor b);
    layer0_outputs(174) <= not b or a;
    layer0_outputs(175) <= a or b;
    layer0_outputs(176) <= not (a xor b);
    layer0_outputs(177) <= not b or a;
    layer0_outputs(178) <= not (a xor b);
    layer0_outputs(179) <= a or b;
    layer0_outputs(180) <= a and not b;
    layer0_outputs(181) <= not b;
    layer0_outputs(182) <= a and not b;
    layer0_outputs(183) <= not (a or b);
    layer0_outputs(184) <= a xor b;
    layer0_outputs(185) <= not b;
    layer0_outputs(186) <= a xor b;
    layer0_outputs(187) <= not b;
    layer0_outputs(188) <= not (a or b);
    layer0_outputs(189) <= not a;
    layer0_outputs(190) <= a or b;
    layer0_outputs(191) <= a or b;
    layer0_outputs(192) <= b and not a;
    layer0_outputs(193) <= 1'b1;
    layer0_outputs(194) <= b and not a;
    layer0_outputs(195) <= not b;
    layer0_outputs(196) <= a and not b;
    layer0_outputs(197) <= a xor b;
    layer0_outputs(198) <= a or b;
    layer0_outputs(199) <= b and not a;
    layer0_outputs(200) <= a and b;
    layer0_outputs(201) <= a;
    layer0_outputs(202) <= b and not a;
    layer0_outputs(203) <= not (a or b);
    layer0_outputs(204) <= 1'b1;
    layer0_outputs(205) <= a or b;
    layer0_outputs(206) <= not b or a;
    layer0_outputs(207) <= not a;
    layer0_outputs(208) <= a;
    layer0_outputs(209) <= a xor b;
    layer0_outputs(210) <= not (a or b);
    layer0_outputs(211) <= b and not a;
    layer0_outputs(212) <= not a or b;
    layer0_outputs(213) <= b;
    layer0_outputs(214) <= not (a or b);
    layer0_outputs(215) <= a;
    layer0_outputs(216) <= not (a or b);
    layer0_outputs(217) <= 1'b1;
    layer0_outputs(218) <= a and not b;
    layer0_outputs(219) <= a or b;
    layer0_outputs(220) <= a xor b;
    layer0_outputs(221) <= a;
    layer0_outputs(222) <= not b;
    layer0_outputs(223) <= a and not b;
    layer0_outputs(224) <= a or b;
    layer0_outputs(225) <= b and not a;
    layer0_outputs(226) <= not b or a;
    layer0_outputs(227) <= not (a or b);
    layer0_outputs(228) <= not b;
    layer0_outputs(229) <= not (a or b);
    layer0_outputs(230) <= a or b;
    layer0_outputs(231) <= 1'b0;
    layer0_outputs(232) <= not (a or b);
    layer0_outputs(233) <= not (a or b);
    layer0_outputs(234) <= not a or b;
    layer0_outputs(235) <= not a or b;
    layer0_outputs(236) <= not a;
    layer0_outputs(237) <= not a;
    layer0_outputs(238) <= not (a xor b);
    layer0_outputs(239) <= not a or b;
    layer0_outputs(240) <= not b or a;
    layer0_outputs(241) <= a or b;
    layer0_outputs(242) <= not b or a;
    layer0_outputs(243) <= a xor b;
    layer0_outputs(244) <= not (a and b);
    layer0_outputs(245) <= a or b;
    layer0_outputs(246) <= not (a or b);
    layer0_outputs(247) <= a or b;
    layer0_outputs(248) <= not (a and b);
    layer0_outputs(249) <= a xor b;
    layer0_outputs(250) <= not (a or b);
    layer0_outputs(251) <= a;
    layer0_outputs(252) <= not a or b;
    layer0_outputs(253) <= 1'b0;
    layer0_outputs(254) <= not (a or b);
    layer0_outputs(255) <= b;
    layer0_outputs(256) <= a or b;
    layer0_outputs(257) <= a or b;
    layer0_outputs(258) <= 1'b1;
    layer0_outputs(259) <= not b or a;
    layer0_outputs(260) <= not (a xor b);
    layer0_outputs(261) <= a;
    layer0_outputs(262) <= not b;
    layer0_outputs(263) <= not (a or b);
    layer0_outputs(264) <= 1'b1;
    layer0_outputs(265) <= not (a xor b);
    layer0_outputs(266) <= not b;
    layer0_outputs(267) <= not (a or b);
    layer0_outputs(268) <= not b or a;
    layer0_outputs(269) <= not b or a;
    layer0_outputs(270) <= not (a or b);
    layer0_outputs(271) <= a and not b;
    layer0_outputs(272) <= not a;
    layer0_outputs(273) <= not a or b;
    layer0_outputs(274) <= b;
    layer0_outputs(275) <= a or b;
    layer0_outputs(276) <= b;
    layer0_outputs(277) <= 1'b1;
    layer0_outputs(278) <= a and not b;
    layer0_outputs(279) <= a xor b;
    layer0_outputs(280) <= a xor b;
    layer0_outputs(281) <= a or b;
    layer0_outputs(282) <= a and not b;
    layer0_outputs(283) <= not (a and b);
    layer0_outputs(284) <= not (a xor b);
    layer0_outputs(285) <= a;
    layer0_outputs(286) <= b;
    layer0_outputs(287) <= a;
    layer0_outputs(288) <= not (a xor b);
    layer0_outputs(289) <= not (a or b);
    layer0_outputs(290) <= a;
    layer0_outputs(291) <= 1'b0;
    layer0_outputs(292) <= b;
    layer0_outputs(293) <= a or b;
    layer0_outputs(294) <= a or b;
    layer0_outputs(295) <= a;
    layer0_outputs(296) <= a or b;
    layer0_outputs(297) <= not b;
    layer0_outputs(298) <= b;
    layer0_outputs(299) <= a or b;
    layer0_outputs(300) <= not b;
    layer0_outputs(301) <= a;
    layer0_outputs(302) <= a xor b;
    layer0_outputs(303) <= not (a or b);
    layer0_outputs(304) <= 1'b0;
    layer0_outputs(305) <= not b;
    layer0_outputs(306) <= b and not a;
    layer0_outputs(307) <= b;
    layer0_outputs(308) <= not a;
    layer0_outputs(309) <= b;
    layer0_outputs(310) <= a;
    layer0_outputs(311) <= a xor b;
    layer0_outputs(312) <= a or b;
    layer0_outputs(313) <= not (a or b);
    layer0_outputs(314) <= 1'b0;
    layer0_outputs(315) <= b;
    layer0_outputs(316) <= a or b;
    layer0_outputs(317) <= a or b;
    layer0_outputs(318) <= not (a xor b);
    layer0_outputs(319) <= not b;
    layer0_outputs(320) <= not (a xor b);
    layer0_outputs(321) <= a or b;
    layer0_outputs(322) <= 1'b0;
    layer0_outputs(323) <= a and b;
    layer0_outputs(324) <= a or b;
    layer0_outputs(325) <= a;
    layer0_outputs(326) <= a xor b;
    layer0_outputs(327) <= a or b;
    layer0_outputs(328) <= b;
    layer0_outputs(329) <= not (a xor b);
    layer0_outputs(330) <= not b;
    layer0_outputs(331) <= a and not b;
    layer0_outputs(332) <= a xor b;
    layer0_outputs(333) <= not b or a;
    layer0_outputs(334) <= a;
    layer0_outputs(335) <= not a;
    layer0_outputs(336) <= not b or a;
    layer0_outputs(337) <= not (a xor b);
    layer0_outputs(338) <= not a or b;
    layer0_outputs(339) <= b;
    layer0_outputs(340) <= b;
    layer0_outputs(341) <= a and not b;
    layer0_outputs(342) <= not b or a;
    layer0_outputs(343) <= a xor b;
    layer0_outputs(344) <= not a;
    layer0_outputs(345) <= a;
    layer0_outputs(346) <= a or b;
    layer0_outputs(347) <= not (a or b);
    layer0_outputs(348) <= not b;
    layer0_outputs(349) <= not a or b;
    layer0_outputs(350) <= a and b;
    layer0_outputs(351) <= a and not b;
    layer0_outputs(352) <= a or b;
    layer0_outputs(353) <= a or b;
    layer0_outputs(354) <= 1'b0;
    layer0_outputs(355) <= a;
    layer0_outputs(356) <= not b or a;
    layer0_outputs(357) <= not (a and b);
    layer0_outputs(358) <= a and not b;
    layer0_outputs(359) <= a xor b;
    layer0_outputs(360) <= b;
    layer0_outputs(361) <= not a;
    layer0_outputs(362) <= a and not b;
    layer0_outputs(363) <= not a or b;
    layer0_outputs(364) <= 1'b0;
    layer0_outputs(365) <= a;
    layer0_outputs(366) <= not a or b;
    layer0_outputs(367) <= not (a or b);
    layer0_outputs(368) <= not b;
    layer0_outputs(369) <= b;
    layer0_outputs(370) <= b and not a;
    layer0_outputs(371) <= b;
    layer0_outputs(372) <= not (a xor b);
    layer0_outputs(373) <= b and not a;
    layer0_outputs(374) <= a xor b;
    layer0_outputs(375) <= not b;
    layer0_outputs(376) <= b and not a;
    layer0_outputs(377) <= not (a and b);
    layer0_outputs(378) <= not (a or b);
    layer0_outputs(379) <= not b;
    layer0_outputs(380) <= b;
    layer0_outputs(381) <= a or b;
    layer0_outputs(382) <= a;
    layer0_outputs(383) <= b and not a;
    layer0_outputs(384) <= not a;
    layer0_outputs(385) <= a xor b;
    layer0_outputs(386) <= not (a or b);
    layer0_outputs(387) <= not (a or b);
    layer0_outputs(388) <= not (a or b);
    layer0_outputs(389) <= not a or b;
    layer0_outputs(390) <= a and not b;
    layer0_outputs(391) <= not a;
    layer0_outputs(392) <= not b or a;
    layer0_outputs(393) <= 1'b0;
    layer0_outputs(394) <= b and not a;
    layer0_outputs(395) <= not (a and b);
    layer0_outputs(396) <= a or b;
    layer0_outputs(397) <= a or b;
    layer0_outputs(398) <= b and not a;
    layer0_outputs(399) <= b;
    layer0_outputs(400) <= not a or b;
    layer0_outputs(401) <= a or b;
    layer0_outputs(402) <= a and not b;
    layer0_outputs(403) <= b and not a;
    layer0_outputs(404) <= 1'b1;
    layer0_outputs(405) <= not (a or b);
    layer0_outputs(406) <= a or b;
    layer0_outputs(407) <= b and not a;
    layer0_outputs(408) <= not a or b;
    layer0_outputs(409) <= not a;
    layer0_outputs(410) <= not b or a;
    layer0_outputs(411) <= a and b;
    layer0_outputs(412) <= a and not b;
    layer0_outputs(413) <= not a or b;
    layer0_outputs(414) <= not (a xor b);
    layer0_outputs(415) <= not a;
    layer0_outputs(416) <= not (a or b);
    layer0_outputs(417) <= not a or b;
    layer0_outputs(418) <= b and not a;
    layer0_outputs(419) <= not (a or b);
    layer0_outputs(420) <= a or b;
    layer0_outputs(421) <= 1'b1;
    layer0_outputs(422) <= a and not b;
    layer0_outputs(423) <= not b;
    layer0_outputs(424) <= not b or a;
    layer0_outputs(425) <= a and not b;
    layer0_outputs(426) <= b;
    layer0_outputs(427) <= not a or b;
    layer0_outputs(428) <= not a;
    layer0_outputs(429) <= not (a or b);
    layer0_outputs(430) <= not b or a;
    layer0_outputs(431) <= a and not b;
    layer0_outputs(432) <= a;
    layer0_outputs(433) <= not b or a;
    layer0_outputs(434) <= not b;
    layer0_outputs(435) <= not (a or b);
    layer0_outputs(436) <= a or b;
    layer0_outputs(437) <= not b or a;
    layer0_outputs(438) <= a;
    layer0_outputs(439) <= a xor b;
    layer0_outputs(440) <= not (a and b);
    layer0_outputs(441) <= not a;
    layer0_outputs(442) <= b and not a;
    layer0_outputs(443) <= a xor b;
    layer0_outputs(444) <= 1'b0;
    layer0_outputs(445) <= not b;
    layer0_outputs(446) <= not a;
    layer0_outputs(447) <= not b;
    layer0_outputs(448) <= not (a and b);
    layer0_outputs(449) <= not (a or b);
    layer0_outputs(450) <= a or b;
    layer0_outputs(451) <= not b;
    layer0_outputs(452) <= not (a or b);
    layer0_outputs(453) <= not (a or b);
    layer0_outputs(454) <= b and not a;
    layer0_outputs(455) <= not b;
    layer0_outputs(456) <= not b or a;
    layer0_outputs(457) <= a xor b;
    layer0_outputs(458) <= a or b;
    layer0_outputs(459) <= a xor b;
    layer0_outputs(460) <= 1'b1;
    layer0_outputs(461) <= b;
    layer0_outputs(462) <= not (a or b);
    layer0_outputs(463) <= b;
    layer0_outputs(464) <= a or b;
    layer0_outputs(465) <= not (a or b);
    layer0_outputs(466) <= a and not b;
    layer0_outputs(467) <= not (a and b);
    layer0_outputs(468) <= 1'b1;
    layer0_outputs(469) <= b;
    layer0_outputs(470) <= a xor b;
    layer0_outputs(471) <= 1'b1;
    layer0_outputs(472) <= a or b;
    layer0_outputs(473) <= not (a or b);
    layer0_outputs(474) <= not (a or b);
    layer0_outputs(475) <= a;
    layer0_outputs(476) <= a and not b;
    layer0_outputs(477) <= b and not a;
    layer0_outputs(478) <= 1'b1;
    layer0_outputs(479) <= a;
    layer0_outputs(480) <= a or b;
    layer0_outputs(481) <= not a;
    layer0_outputs(482) <= a;
    layer0_outputs(483) <= a xor b;
    layer0_outputs(484) <= not b or a;
    layer0_outputs(485) <= a xor b;
    layer0_outputs(486) <= a xor b;
    layer0_outputs(487) <= not a;
    layer0_outputs(488) <= not b or a;
    layer0_outputs(489) <= b and not a;
    layer0_outputs(490) <= not a;
    layer0_outputs(491) <= b;
    layer0_outputs(492) <= not a;
    layer0_outputs(493) <= a and not b;
    layer0_outputs(494) <= not (a or b);
    layer0_outputs(495) <= not (a and b);
    layer0_outputs(496) <= a or b;
    layer0_outputs(497) <= a;
    layer0_outputs(498) <= a and not b;
    layer0_outputs(499) <= 1'b0;
    layer0_outputs(500) <= not b;
    layer0_outputs(501) <= not (a or b);
    layer0_outputs(502) <= a;
    layer0_outputs(503) <= not a;
    layer0_outputs(504) <= a;
    layer0_outputs(505) <= not (a or b);
    layer0_outputs(506) <= not (a xor b);
    layer0_outputs(507) <= a or b;
    layer0_outputs(508) <= not (a and b);
    layer0_outputs(509) <= a xor b;
    layer0_outputs(510) <= a or b;
    layer0_outputs(511) <= not b;
    layer0_outputs(512) <= not (a xor b);
    layer0_outputs(513) <= a xor b;
    layer0_outputs(514) <= a xor b;
    layer0_outputs(515) <= a xor b;
    layer0_outputs(516) <= not (a or b);
    layer0_outputs(517) <= b;
    layer0_outputs(518) <= not (a or b);
    layer0_outputs(519) <= not a;
    layer0_outputs(520) <= a;
    layer0_outputs(521) <= a;
    layer0_outputs(522) <= a or b;
    layer0_outputs(523) <= a xor b;
    layer0_outputs(524) <= 1'b1;
    layer0_outputs(525) <= not (a or b);
    layer0_outputs(526) <= not a or b;
    layer0_outputs(527) <= not a;
    layer0_outputs(528) <= a and not b;
    layer0_outputs(529) <= not (a and b);
    layer0_outputs(530) <= b;
    layer0_outputs(531) <= a;
    layer0_outputs(532) <= not (a or b);
    layer0_outputs(533) <= not a;
    layer0_outputs(534) <= not (a xor b);
    layer0_outputs(535) <= a;
    layer0_outputs(536) <= not (a and b);
    layer0_outputs(537) <= a and b;
    layer0_outputs(538) <= not b or a;
    layer0_outputs(539) <= not a;
    layer0_outputs(540) <= not b;
    layer0_outputs(541) <= not (a or b);
    layer0_outputs(542) <= not b or a;
    layer0_outputs(543) <= not (a xor b);
    layer0_outputs(544) <= not b;
    layer0_outputs(545) <= a xor b;
    layer0_outputs(546) <= a xor b;
    layer0_outputs(547) <= a or b;
    layer0_outputs(548) <= a;
    layer0_outputs(549) <= not a;
    layer0_outputs(550) <= not (a xor b);
    layer0_outputs(551) <= b and not a;
    layer0_outputs(552) <= not (a xor b);
    layer0_outputs(553) <= not b;
    layer0_outputs(554) <= a and not b;
    layer0_outputs(555) <= not b;
    layer0_outputs(556) <= not a;
    layer0_outputs(557) <= a;
    layer0_outputs(558) <= not (a or b);
    layer0_outputs(559) <= not (a or b);
    layer0_outputs(560) <= not a;
    layer0_outputs(561) <= a or b;
    layer0_outputs(562) <= not a;
    layer0_outputs(563) <= not b or a;
    layer0_outputs(564) <= 1'b1;
    layer0_outputs(565) <= a or b;
    layer0_outputs(566) <= not a or b;
    layer0_outputs(567) <= a;
    layer0_outputs(568) <= a or b;
    layer0_outputs(569) <= not (a xor b);
    layer0_outputs(570) <= not b;
    layer0_outputs(571) <= b;
    layer0_outputs(572) <= not (a or b);
    layer0_outputs(573) <= not a or b;
    layer0_outputs(574) <= a;
    layer0_outputs(575) <= not (a or b);
    layer0_outputs(576) <= not a or b;
    layer0_outputs(577) <= not a or b;
    layer0_outputs(578) <= not (a xor b);
    layer0_outputs(579) <= not b;
    layer0_outputs(580) <= a and not b;
    layer0_outputs(581) <= b and not a;
    layer0_outputs(582) <= a or b;
    layer0_outputs(583) <= a;
    layer0_outputs(584) <= not (a and b);
    layer0_outputs(585) <= not a;
    layer0_outputs(586) <= a;
    layer0_outputs(587) <= b;
    layer0_outputs(588) <= not b;
    layer0_outputs(589) <= not (a and b);
    layer0_outputs(590) <= not a;
    layer0_outputs(591) <= not (a or b);
    layer0_outputs(592) <= b and not a;
    layer0_outputs(593) <= not (a xor b);
    layer0_outputs(594) <= not b or a;
    layer0_outputs(595) <= a xor b;
    layer0_outputs(596) <= b and not a;
    layer0_outputs(597) <= not (a xor b);
    layer0_outputs(598) <= not (a or b);
    layer0_outputs(599) <= not b or a;
    layer0_outputs(600) <= a xor b;
    layer0_outputs(601) <= a or b;
    layer0_outputs(602) <= b and not a;
    layer0_outputs(603) <= a and b;
    layer0_outputs(604) <= not b or a;
    layer0_outputs(605) <= not a or b;
    layer0_outputs(606) <= not (a or b);
    layer0_outputs(607) <= a and not b;
    layer0_outputs(608) <= b and not a;
    layer0_outputs(609) <= not a or b;
    layer0_outputs(610) <= not a;
    layer0_outputs(611) <= b;
    layer0_outputs(612) <= a xor b;
    layer0_outputs(613) <= b and not a;
    layer0_outputs(614) <= not b;
    layer0_outputs(615) <= not (a or b);
    layer0_outputs(616) <= a and b;
    layer0_outputs(617) <= a or b;
    layer0_outputs(618) <= not a;
    layer0_outputs(619) <= not a;
    layer0_outputs(620) <= b and not a;
    layer0_outputs(621) <= not (a or b);
    layer0_outputs(622) <= b and not a;
    layer0_outputs(623) <= not (a or b);
    layer0_outputs(624) <= not b or a;
    layer0_outputs(625) <= not (a or b);
    layer0_outputs(626) <= a;
    layer0_outputs(627) <= a or b;
    layer0_outputs(628) <= not b or a;
    layer0_outputs(629) <= a and not b;
    layer0_outputs(630) <= 1'b1;
    layer0_outputs(631) <= b;
    layer0_outputs(632) <= not (a or b);
    layer0_outputs(633) <= b and not a;
    layer0_outputs(634) <= not a or b;
    layer0_outputs(635) <= not (a xor b);
    layer0_outputs(636) <= not b;
    layer0_outputs(637) <= not a;
    layer0_outputs(638) <= not b or a;
    layer0_outputs(639) <= not a;
    layer0_outputs(640) <= not (a xor b);
    layer0_outputs(641) <= a xor b;
    layer0_outputs(642) <= a;
    layer0_outputs(643) <= b and not a;
    layer0_outputs(644) <= not b or a;
    layer0_outputs(645) <= not b;
    layer0_outputs(646) <= not (a xor b);
    layer0_outputs(647) <= not (a and b);
    layer0_outputs(648) <= a or b;
    layer0_outputs(649) <= not (a or b);
    layer0_outputs(650) <= a and b;
    layer0_outputs(651) <= a;
    layer0_outputs(652) <= a and not b;
    layer0_outputs(653) <= not b;
    layer0_outputs(654) <= a and b;
    layer0_outputs(655) <= not b or a;
    layer0_outputs(656) <= a or b;
    layer0_outputs(657) <= a;
    layer0_outputs(658) <= a xor b;
    layer0_outputs(659) <= a and not b;
    layer0_outputs(660) <= not (a xor b);
    layer0_outputs(661) <= a and b;
    layer0_outputs(662) <= b and not a;
    layer0_outputs(663) <= not (a and b);
    layer0_outputs(664) <= not a;
    layer0_outputs(665) <= a xor b;
    layer0_outputs(666) <= not (a xor b);
    layer0_outputs(667) <= not (a xor b);
    layer0_outputs(668) <= a or b;
    layer0_outputs(669) <= a;
    layer0_outputs(670) <= a;
    layer0_outputs(671) <= not a or b;
    layer0_outputs(672) <= b and not a;
    layer0_outputs(673) <= not b or a;
    layer0_outputs(674) <= a xor b;
    layer0_outputs(675) <= b and not a;
    layer0_outputs(676) <= b;
    layer0_outputs(677) <= b;
    layer0_outputs(678) <= not (a or b);
    layer0_outputs(679) <= a and not b;
    layer0_outputs(680) <= b;
    layer0_outputs(681) <= not a;
    layer0_outputs(682) <= not (a or b);
    layer0_outputs(683) <= a;
    layer0_outputs(684) <= not a;
    layer0_outputs(685) <= not b;
    layer0_outputs(686) <= not b;
    layer0_outputs(687) <= a or b;
    layer0_outputs(688) <= not b or a;
    layer0_outputs(689) <= a and b;
    layer0_outputs(690) <= not (a or b);
    layer0_outputs(691) <= a or b;
    layer0_outputs(692) <= a;
    layer0_outputs(693) <= not b or a;
    layer0_outputs(694) <= 1'b1;
    layer0_outputs(695) <= b and not a;
    layer0_outputs(696) <= not a;
    layer0_outputs(697) <= a xor b;
    layer0_outputs(698) <= not a;
    layer0_outputs(699) <= a or b;
    layer0_outputs(700) <= not (a or b);
    layer0_outputs(701) <= not a or b;
    layer0_outputs(702) <= b;
    layer0_outputs(703) <= b and not a;
    layer0_outputs(704) <= a;
    layer0_outputs(705) <= b;
    layer0_outputs(706) <= not (a or b);
    layer0_outputs(707) <= not a;
    layer0_outputs(708) <= not (a or b);
    layer0_outputs(709) <= b;
    layer0_outputs(710) <= 1'b1;
    layer0_outputs(711) <= not b;
    layer0_outputs(712) <= not a;
    layer0_outputs(713) <= a and not b;
    layer0_outputs(714) <= a and not b;
    layer0_outputs(715) <= not b or a;
    layer0_outputs(716) <= a xor b;
    layer0_outputs(717) <= a or b;
    layer0_outputs(718) <= not a or b;
    layer0_outputs(719) <= not (a or b);
    layer0_outputs(720) <= not (a and b);
    layer0_outputs(721) <= a and not b;
    layer0_outputs(722) <= not (a or b);
    layer0_outputs(723) <= not b or a;
    layer0_outputs(724) <= not (a and b);
    layer0_outputs(725) <= a;
    layer0_outputs(726) <= a or b;
    layer0_outputs(727) <= a or b;
    layer0_outputs(728) <= a;
    layer0_outputs(729) <= not (a or b);
    layer0_outputs(730) <= a or b;
    layer0_outputs(731) <= a and not b;
    layer0_outputs(732) <= a or b;
    layer0_outputs(733) <= a;
    layer0_outputs(734) <= a or b;
    layer0_outputs(735) <= not (a and b);
    layer0_outputs(736) <= b and not a;
    layer0_outputs(737) <= not (a or b);
    layer0_outputs(738) <= a or b;
    layer0_outputs(739) <= not (a and b);
    layer0_outputs(740) <= a or b;
    layer0_outputs(741) <= not a;
    layer0_outputs(742) <= not (a xor b);
    layer0_outputs(743) <= b;
    layer0_outputs(744) <= a or b;
    layer0_outputs(745) <= a xor b;
    layer0_outputs(746) <= not (a xor b);
    layer0_outputs(747) <= a xor b;
    layer0_outputs(748) <= 1'b0;
    layer0_outputs(749) <= not a or b;
    layer0_outputs(750) <= not a;
    layer0_outputs(751) <= not (a xor b);
    layer0_outputs(752) <= b and not a;
    layer0_outputs(753) <= a or b;
    layer0_outputs(754) <= b;
    layer0_outputs(755) <= not b or a;
    layer0_outputs(756) <= a xor b;
    layer0_outputs(757) <= not a;
    layer0_outputs(758) <= not b or a;
    layer0_outputs(759) <= b;
    layer0_outputs(760) <= not b;
    layer0_outputs(761) <= b and not a;
    layer0_outputs(762) <= b;
    layer0_outputs(763) <= not b or a;
    layer0_outputs(764) <= b;
    layer0_outputs(765) <= 1'b1;
    layer0_outputs(766) <= not b;
    layer0_outputs(767) <= b;
    layer0_outputs(768) <= a xor b;
    layer0_outputs(769) <= b;
    layer0_outputs(770) <= not b or a;
    layer0_outputs(771) <= not (a xor b);
    layer0_outputs(772) <= a xor b;
    layer0_outputs(773) <= not (a or b);
    layer0_outputs(774) <= not b or a;
    layer0_outputs(775) <= a or b;
    layer0_outputs(776) <= a and b;
    layer0_outputs(777) <= not (a or b);
    layer0_outputs(778) <= a and not b;
    layer0_outputs(779) <= b;
    layer0_outputs(780) <= b and not a;
    layer0_outputs(781) <= a or b;
    layer0_outputs(782) <= not (a or b);
    layer0_outputs(783) <= not (a xor b);
    layer0_outputs(784) <= not (a xor b);
    layer0_outputs(785) <= not b;
    layer0_outputs(786) <= b;
    layer0_outputs(787) <= not (a and b);
    layer0_outputs(788) <= a;
    layer0_outputs(789) <= not (a and b);
    layer0_outputs(790) <= 1'b1;
    layer0_outputs(791) <= a xor b;
    layer0_outputs(792) <= b and not a;
    layer0_outputs(793) <= not (a or b);
    layer0_outputs(794) <= b and not a;
    layer0_outputs(795) <= not (a xor b);
    layer0_outputs(796) <= a and not b;
    layer0_outputs(797) <= not b;
    layer0_outputs(798) <= a xor b;
    layer0_outputs(799) <= not a or b;
    layer0_outputs(800) <= not b or a;
    layer0_outputs(801) <= not (a xor b);
    layer0_outputs(802) <= a;
    layer0_outputs(803) <= not b or a;
    layer0_outputs(804) <= 1'b0;
    layer0_outputs(805) <= a or b;
    layer0_outputs(806) <= not (a or b);
    layer0_outputs(807) <= a or b;
    layer0_outputs(808) <= not (a or b);
    layer0_outputs(809) <= not a or b;
    layer0_outputs(810) <= 1'b0;
    layer0_outputs(811) <= 1'b1;
    layer0_outputs(812) <= a;
    layer0_outputs(813) <= a and b;
    layer0_outputs(814) <= not (a or b);
    layer0_outputs(815) <= not (a xor b);
    layer0_outputs(816) <= not (a or b);
    layer0_outputs(817) <= a xor b;
    layer0_outputs(818) <= not b or a;
    layer0_outputs(819) <= b;
    layer0_outputs(820) <= a or b;
    layer0_outputs(821) <= a and not b;
    layer0_outputs(822) <= a or b;
    layer0_outputs(823) <= b and not a;
    layer0_outputs(824) <= not (a or b);
    layer0_outputs(825) <= a xor b;
    layer0_outputs(826) <= not b or a;
    layer0_outputs(827) <= a or b;
    layer0_outputs(828) <= b;
    layer0_outputs(829) <= not (a xor b);
    layer0_outputs(830) <= 1'b0;
    layer0_outputs(831) <= a or b;
    layer0_outputs(832) <= not (a or b);
    layer0_outputs(833) <= not (a xor b);
    layer0_outputs(834) <= not a;
    layer0_outputs(835) <= a and not b;
    layer0_outputs(836) <= not (a or b);
    layer0_outputs(837) <= not (a or b);
    layer0_outputs(838) <= a and not b;
    layer0_outputs(839) <= not a or b;
    layer0_outputs(840) <= a or b;
    layer0_outputs(841) <= a;
    layer0_outputs(842) <= not (a or b);
    layer0_outputs(843) <= a and b;
    layer0_outputs(844) <= a;
    layer0_outputs(845) <= a or b;
    layer0_outputs(846) <= not a;
    layer0_outputs(847) <= b;
    layer0_outputs(848) <= not (a or b);
    layer0_outputs(849) <= a xor b;
    layer0_outputs(850) <= not a;
    layer0_outputs(851) <= a;
    layer0_outputs(852) <= a;
    layer0_outputs(853) <= 1'b1;
    layer0_outputs(854) <= not (a or b);
    layer0_outputs(855) <= not (a xor b);
    layer0_outputs(856) <= not b;
    layer0_outputs(857) <= not (a xor b);
    layer0_outputs(858) <= not (a xor b);
    layer0_outputs(859) <= a xor b;
    layer0_outputs(860) <= a;
    layer0_outputs(861) <= b and not a;
    layer0_outputs(862) <= not (a or b);
    layer0_outputs(863) <= not (a xor b);
    layer0_outputs(864) <= 1'b1;
    layer0_outputs(865) <= a and b;
    layer0_outputs(866) <= not b;
    layer0_outputs(867) <= a or b;
    layer0_outputs(868) <= not (a xor b);
    layer0_outputs(869) <= 1'b0;
    layer0_outputs(870) <= a;
    layer0_outputs(871) <= a xor b;
    layer0_outputs(872) <= a or b;
    layer0_outputs(873) <= not (a xor b);
    layer0_outputs(874) <= not a or b;
    layer0_outputs(875) <= not a or b;
    layer0_outputs(876) <= not a or b;
    layer0_outputs(877) <= not a or b;
    layer0_outputs(878) <= 1'b1;
    layer0_outputs(879) <= not b;
    layer0_outputs(880) <= not a or b;
    layer0_outputs(881) <= b and not a;
    layer0_outputs(882) <= a or b;
    layer0_outputs(883) <= not b;
    layer0_outputs(884) <= not (a or b);
    layer0_outputs(885) <= a xor b;
    layer0_outputs(886) <= not a or b;
    layer0_outputs(887) <= not b;
    layer0_outputs(888) <= not (a xor b);
    layer0_outputs(889) <= not (a or b);
    layer0_outputs(890) <= b and not a;
    layer0_outputs(891) <= 1'b0;
    layer0_outputs(892) <= a xor b;
    layer0_outputs(893) <= a;
    layer0_outputs(894) <= not (a or b);
    layer0_outputs(895) <= not a or b;
    layer0_outputs(896) <= not (a or b);
    layer0_outputs(897) <= a or b;
    layer0_outputs(898) <= not b;
    layer0_outputs(899) <= b;
    layer0_outputs(900) <= 1'b0;
    layer0_outputs(901) <= b and not a;
    layer0_outputs(902) <= a or b;
    layer0_outputs(903) <= a xor b;
    layer0_outputs(904) <= not a;
    layer0_outputs(905) <= not (a or b);
    layer0_outputs(906) <= not a;
    layer0_outputs(907) <= a and not b;
    layer0_outputs(908) <= not b or a;
    layer0_outputs(909) <= a xor b;
    layer0_outputs(910) <= a or b;
    layer0_outputs(911) <= a;
    layer0_outputs(912) <= a;
    layer0_outputs(913) <= not (a or b);
    layer0_outputs(914) <= not b or a;
    layer0_outputs(915) <= a and not b;
    layer0_outputs(916) <= a xor b;
    layer0_outputs(917) <= a xor b;
    layer0_outputs(918) <= a;
    layer0_outputs(919) <= b and not a;
    layer0_outputs(920) <= a;
    layer0_outputs(921) <= b;
    layer0_outputs(922) <= not (a and b);
    layer0_outputs(923) <= a;
    layer0_outputs(924) <= a or b;
    layer0_outputs(925) <= a and not b;
    layer0_outputs(926) <= not (a or b);
    layer0_outputs(927) <= a and not b;
    layer0_outputs(928) <= not (a and b);
    layer0_outputs(929) <= a and not b;
    layer0_outputs(930) <= not a;
    layer0_outputs(931) <= not b;
    layer0_outputs(932) <= not (a and b);
    layer0_outputs(933) <= a and not b;
    layer0_outputs(934) <= b and not a;
    layer0_outputs(935) <= a;
    layer0_outputs(936) <= b;
    layer0_outputs(937) <= not a;
    layer0_outputs(938) <= not (a or b);
    layer0_outputs(939) <= not (a or b);
    layer0_outputs(940) <= not (a or b);
    layer0_outputs(941) <= a;
    layer0_outputs(942) <= a xor b;
    layer0_outputs(943) <= a or b;
    layer0_outputs(944) <= not (a and b);
    layer0_outputs(945) <= a;
    layer0_outputs(946) <= a xor b;
    layer0_outputs(947) <= a;
    layer0_outputs(948) <= a or b;
    layer0_outputs(949) <= not a;
    layer0_outputs(950) <= not (a xor b);
    layer0_outputs(951) <= not b or a;
    layer0_outputs(952) <= not (a xor b);
    layer0_outputs(953) <= a;
    layer0_outputs(954) <= a xor b;
    layer0_outputs(955) <= not a or b;
    layer0_outputs(956) <= not (a and b);
    layer0_outputs(957) <= b and not a;
    layer0_outputs(958) <= not (a or b);
    layer0_outputs(959) <= 1'b0;
    layer0_outputs(960) <= not b or a;
    layer0_outputs(961) <= b and not a;
    layer0_outputs(962) <= a and b;
    layer0_outputs(963) <= a or b;
    layer0_outputs(964) <= not b or a;
    layer0_outputs(965) <= a xor b;
    layer0_outputs(966) <= a;
    layer0_outputs(967) <= not (a or b);
    layer0_outputs(968) <= b;
    layer0_outputs(969) <= not (a xor b);
    layer0_outputs(970) <= not a;
    layer0_outputs(971) <= not b or a;
    layer0_outputs(972) <= not a;
    layer0_outputs(973) <= a or b;
    layer0_outputs(974) <= not (a and b);
    layer0_outputs(975) <= a and not b;
    layer0_outputs(976) <= not (a or b);
    layer0_outputs(977) <= a;
    layer0_outputs(978) <= not (a or b);
    layer0_outputs(979) <= not (a xor b);
    layer0_outputs(980) <= not b;
    layer0_outputs(981) <= 1'b0;
    layer0_outputs(982) <= 1'b1;
    layer0_outputs(983) <= b and not a;
    layer0_outputs(984) <= not (a xor b);
    layer0_outputs(985) <= b;
    layer0_outputs(986) <= not b;
    layer0_outputs(987) <= a and not b;
    layer0_outputs(988) <= not (a xor b);
    layer0_outputs(989) <= b and not a;
    layer0_outputs(990) <= a;
    layer0_outputs(991) <= not (a or b);
    layer0_outputs(992) <= not a or b;
    layer0_outputs(993) <= a and not b;
    layer0_outputs(994) <= not (a and b);
    layer0_outputs(995) <= not (a or b);
    layer0_outputs(996) <= not b;
    layer0_outputs(997) <= a or b;
    layer0_outputs(998) <= a and not b;
    layer0_outputs(999) <= not (a or b);
    layer0_outputs(1000) <= a and b;
    layer0_outputs(1001) <= a and not b;
    layer0_outputs(1002) <= a or b;
    layer0_outputs(1003) <= not a;
    layer0_outputs(1004) <= b;
    layer0_outputs(1005) <= a;
    layer0_outputs(1006) <= b;
    layer0_outputs(1007) <= a or b;
    layer0_outputs(1008) <= 1'b1;
    layer0_outputs(1009) <= not a;
    layer0_outputs(1010) <= a or b;
    layer0_outputs(1011) <= not (a or b);
    layer0_outputs(1012) <= not (a xor b);
    layer0_outputs(1013) <= not (a or b);
    layer0_outputs(1014) <= not (a xor b);
    layer0_outputs(1015) <= not b or a;
    layer0_outputs(1016) <= b and not a;
    layer0_outputs(1017) <= not a or b;
    layer0_outputs(1018) <= a and b;
    layer0_outputs(1019) <= not (a xor b);
    layer0_outputs(1020) <= not a;
    layer0_outputs(1021) <= not b;
    layer0_outputs(1022) <= a or b;
    layer0_outputs(1023) <= b;
    layer0_outputs(1024) <= b;
    layer0_outputs(1025) <= 1'b0;
    layer0_outputs(1026) <= b;
    layer0_outputs(1027) <= a or b;
    layer0_outputs(1028) <= b and not a;
    layer0_outputs(1029) <= not (a or b);
    layer0_outputs(1030) <= not (a xor b);
    layer0_outputs(1031) <= b;
    layer0_outputs(1032) <= b and not a;
    layer0_outputs(1033) <= not (a or b);
    layer0_outputs(1034) <= a and not b;
    layer0_outputs(1035) <= a or b;
    layer0_outputs(1036) <= a or b;
    layer0_outputs(1037) <= a xor b;
    layer0_outputs(1038) <= not a;
    layer0_outputs(1039) <= a and not b;
    layer0_outputs(1040) <= 1'b1;
    layer0_outputs(1041) <= not b or a;
    layer0_outputs(1042) <= a and not b;
    layer0_outputs(1043) <= a xor b;
    layer0_outputs(1044) <= not (a or b);
    layer0_outputs(1045) <= not (a xor b);
    layer0_outputs(1046) <= not (a xor b);
    layer0_outputs(1047) <= not (a xor b);
    layer0_outputs(1048) <= a and b;
    layer0_outputs(1049) <= not a;
    layer0_outputs(1050) <= not a or b;
    layer0_outputs(1051) <= not a or b;
    layer0_outputs(1052) <= a xor b;
    layer0_outputs(1053) <= not b or a;
    layer0_outputs(1054) <= not a or b;
    layer0_outputs(1055) <= 1'b0;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= a and b;
    layer0_outputs(1058) <= not b;
    layer0_outputs(1059) <= not (a and b);
    layer0_outputs(1060) <= not a;
    layer0_outputs(1061) <= not b or a;
    layer0_outputs(1062) <= a or b;
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= not (a or b);
    layer0_outputs(1065) <= 1'b0;
    layer0_outputs(1066) <= not b;
    layer0_outputs(1067) <= not b or a;
    layer0_outputs(1068) <= a xor b;
    layer0_outputs(1069) <= not (a xor b);
    layer0_outputs(1070) <= not (a xor b);
    layer0_outputs(1071) <= a or b;
    layer0_outputs(1072) <= not (a xor b);
    layer0_outputs(1073) <= not b or a;
    layer0_outputs(1074) <= a;
    layer0_outputs(1075) <= not b;
    layer0_outputs(1076) <= a and not b;
    layer0_outputs(1077) <= not (a or b);
    layer0_outputs(1078) <= a and not b;
    layer0_outputs(1079) <= b and not a;
    layer0_outputs(1080) <= a or b;
    layer0_outputs(1081) <= b;
    layer0_outputs(1082) <= a;
    layer0_outputs(1083) <= a xor b;
    layer0_outputs(1084) <= b;
    layer0_outputs(1085) <= a or b;
    layer0_outputs(1086) <= a and b;
    layer0_outputs(1087) <= not (a xor b);
    layer0_outputs(1088) <= a;
    layer0_outputs(1089) <= a;
    layer0_outputs(1090) <= not b;
    layer0_outputs(1091) <= not (a xor b);
    layer0_outputs(1092) <= 1'b0;
    layer0_outputs(1093) <= not a;
    layer0_outputs(1094) <= not b;
    layer0_outputs(1095) <= a;
    layer0_outputs(1096) <= not b or a;
    layer0_outputs(1097) <= a;
    layer0_outputs(1098) <= not (a or b);
    layer0_outputs(1099) <= not a;
    layer0_outputs(1100) <= b;
    layer0_outputs(1101) <= not (a or b);
    layer0_outputs(1102) <= a xor b;
    layer0_outputs(1103) <= not (a xor b);
    layer0_outputs(1104) <= b and not a;
    layer0_outputs(1105) <= a;
    layer0_outputs(1106) <= b;
    layer0_outputs(1107) <= a xor b;
    layer0_outputs(1108) <= a or b;
    layer0_outputs(1109) <= not (a or b);
    layer0_outputs(1110) <= not a;
    layer0_outputs(1111) <= not a;
    layer0_outputs(1112) <= 1'b0;
    layer0_outputs(1113) <= not b or a;
    layer0_outputs(1114) <= a xor b;
    layer0_outputs(1115) <= b and not a;
    layer0_outputs(1116) <= not a;
    layer0_outputs(1117) <= not (a or b);
    layer0_outputs(1118) <= a or b;
    layer0_outputs(1119) <= not (a or b);
    layer0_outputs(1120) <= not a;
    layer0_outputs(1121) <= a and not b;
    layer0_outputs(1122) <= a and b;
    layer0_outputs(1123) <= a and b;
    layer0_outputs(1124) <= not b or a;
    layer0_outputs(1125) <= not (a or b);
    layer0_outputs(1126) <= a xor b;
    layer0_outputs(1127) <= 1'b1;
    layer0_outputs(1128) <= not (a xor b);
    layer0_outputs(1129) <= not (a or b);
    layer0_outputs(1130) <= not a;
    layer0_outputs(1131) <= not (a or b);
    layer0_outputs(1132) <= not (a or b);
    layer0_outputs(1133) <= not (a or b);
    layer0_outputs(1134) <= b;
    layer0_outputs(1135) <= a or b;
    layer0_outputs(1136) <= not b;
    layer0_outputs(1137) <= not (a or b);
    layer0_outputs(1138) <= a or b;
    layer0_outputs(1139) <= not a or b;
    layer0_outputs(1140) <= 1'b0;
    layer0_outputs(1141) <= a or b;
    layer0_outputs(1142) <= not a;
    layer0_outputs(1143) <= 1'b1;
    layer0_outputs(1144) <= not (a or b);
    layer0_outputs(1145) <= not (a or b);
    layer0_outputs(1146) <= a or b;
    layer0_outputs(1147) <= a or b;
    layer0_outputs(1148) <= not b;
    layer0_outputs(1149) <= not (a xor b);
    layer0_outputs(1150) <= not (a or b);
    layer0_outputs(1151) <= a xor b;
    layer0_outputs(1152) <= b;
    layer0_outputs(1153) <= not (a and b);
    layer0_outputs(1154) <= a or b;
    layer0_outputs(1155) <= not a;
    layer0_outputs(1156) <= 1'b1;
    layer0_outputs(1157) <= not b or a;
    layer0_outputs(1158) <= a;
    layer0_outputs(1159) <= b;
    layer0_outputs(1160) <= a or b;
    layer0_outputs(1161) <= not (a and b);
    layer0_outputs(1162) <= b;
    layer0_outputs(1163) <= a and not b;
    layer0_outputs(1164) <= not a or b;
    layer0_outputs(1165) <= not (a and b);
    layer0_outputs(1166) <= a and not b;
    layer0_outputs(1167) <= not (a and b);
    layer0_outputs(1168) <= a or b;
    layer0_outputs(1169) <= b;
    layer0_outputs(1170) <= not (a and b);
    layer0_outputs(1171) <= not a;
    layer0_outputs(1172) <= 1'b0;
    layer0_outputs(1173) <= not a;
    layer0_outputs(1174) <= not b or a;
    layer0_outputs(1175) <= a;
    layer0_outputs(1176) <= a and not b;
    layer0_outputs(1177) <= not (a xor b);
    layer0_outputs(1178) <= a;
    layer0_outputs(1179) <= not b;
    layer0_outputs(1180) <= a xor b;
    layer0_outputs(1181) <= a or b;
    layer0_outputs(1182) <= a;
    layer0_outputs(1183) <= 1'b1;
    layer0_outputs(1184) <= a;
    layer0_outputs(1185) <= not a;
    layer0_outputs(1186) <= a;
    layer0_outputs(1187) <= a or b;
    layer0_outputs(1188) <= not b or a;
    layer0_outputs(1189) <= a xor b;
    layer0_outputs(1190) <= not a;
    layer0_outputs(1191) <= a or b;
    layer0_outputs(1192) <= not a or b;
    layer0_outputs(1193) <= a and not b;
    layer0_outputs(1194) <= not b;
    layer0_outputs(1195) <= not b or a;
    layer0_outputs(1196) <= not (a or b);
    layer0_outputs(1197) <= not a or b;
    layer0_outputs(1198) <= not (a xor b);
    layer0_outputs(1199) <= 1'b1;
    layer0_outputs(1200) <= not b;
    layer0_outputs(1201) <= not a;
    layer0_outputs(1202) <= not (a xor b);
    layer0_outputs(1203) <= not (a or b);
    layer0_outputs(1204) <= a or b;
    layer0_outputs(1205) <= a and not b;
    layer0_outputs(1206) <= not (a or b);
    layer0_outputs(1207) <= b;
    layer0_outputs(1208) <= not (a xor b);
    layer0_outputs(1209) <= not a;
    layer0_outputs(1210) <= not (a or b);
    layer0_outputs(1211) <= not (a xor b);
    layer0_outputs(1212) <= a or b;
    layer0_outputs(1213) <= a;
    layer0_outputs(1214) <= not a or b;
    layer0_outputs(1215) <= a and b;
    layer0_outputs(1216) <= not b or a;
    layer0_outputs(1217) <= not a;
    layer0_outputs(1218) <= not a or b;
    layer0_outputs(1219) <= b and not a;
    layer0_outputs(1220) <= not b;
    layer0_outputs(1221) <= not (a or b);
    layer0_outputs(1222) <= not (a or b);
    layer0_outputs(1223) <= a;
    layer0_outputs(1224) <= a xor b;
    layer0_outputs(1225) <= not (a xor b);
    layer0_outputs(1226) <= not b or a;
    layer0_outputs(1227) <= not a;
    layer0_outputs(1228) <= a;
    layer0_outputs(1229) <= not (a or b);
    layer0_outputs(1230) <= not b or a;
    layer0_outputs(1231) <= not b or a;
    layer0_outputs(1232) <= a and not b;
    layer0_outputs(1233) <= not (a or b);
    layer0_outputs(1234) <= not (a or b);
    layer0_outputs(1235) <= a or b;
    layer0_outputs(1236) <= 1'b1;
    layer0_outputs(1237) <= not b;
    layer0_outputs(1238) <= b;
    layer0_outputs(1239) <= not a;
    layer0_outputs(1240) <= not a;
    layer0_outputs(1241) <= a;
    layer0_outputs(1242) <= not (a or b);
    layer0_outputs(1243) <= a and b;
    layer0_outputs(1244) <= not b or a;
    layer0_outputs(1245) <= a xor b;
    layer0_outputs(1246) <= a and not b;
    layer0_outputs(1247) <= a and b;
    layer0_outputs(1248) <= a or b;
    layer0_outputs(1249) <= a xor b;
    layer0_outputs(1250) <= a or b;
    layer0_outputs(1251) <= not a;
    layer0_outputs(1252) <= 1'b1;
    layer0_outputs(1253) <= a or b;
    layer0_outputs(1254) <= not (a or b);
    layer0_outputs(1255) <= a or b;
    layer0_outputs(1256) <= b and not a;
    layer0_outputs(1257) <= not (a xor b);
    layer0_outputs(1258) <= not b or a;
    layer0_outputs(1259) <= a;
    layer0_outputs(1260) <= a or b;
    layer0_outputs(1261) <= not a;
    layer0_outputs(1262) <= a or b;
    layer0_outputs(1263) <= a and b;
    layer0_outputs(1264) <= not (a or b);
    layer0_outputs(1265) <= a xor b;
    layer0_outputs(1266) <= a and not b;
    layer0_outputs(1267) <= not (a and b);
    layer0_outputs(1268) <= not (a or b);
    layer0_outputs(1269) <= a;
    layer0_outputs(1270) <= not (a and b);
    layer0_outputs(1271) <= a;
    layer0_outputs(1272) <= not (a xor b);
    layer0_outputs(1273) <= b and not a;
    layer0_outputs(1274) <= b and not a;
    layer0_outputs(1275) <= 1'b1;
    layer0_outputs(1276) <= not (a xor b);
    layer0_outputs(1277) <= not b;
    layer0_outputs(1278) <= not a;
    layer0_outputs(1279) <= a;
    layer0_outputs(1280) <= a and not b;
    layer0_outputs(1281) <= b;
    layer0_outputs(1282) <= b;
    layer0_outputs(1283) <= not b or a;
    layer0_outputs(1284) <= b;
    layer0_outputs(1285) <= b and not a;
    layer0_outputs(1286) <= not a or b;
    layer0_outputs(1287) <= a xor b;
    layer0_outputs(1288) <= not a or b;
    layer0_outputs(1289) <= not (a xor b);
    layer0_outputs(1290) <= not (a xor b);
    layer0_outputs(1291) <= not b or a;
    layer0_outputs(1292) <= not (a xor b);
    layer0_outputs(1293) <= not b;
    layer0_outputs(1294) <= a and b;
    layer0_outputs(1295) <= not (a xor b);
    layer0_outputs(1296) <= not (a xor b);
    layer0_outputs(1297) <= a;
    layer0_outputs(1298) <= 1'b0;
    layer0_outputs(1299) <= not b or a;
    layer0_outputs(1300) <= 1'b1;
    layer0_outputs(1301) <= b;
    layer0_outputs(1302) <= b;
    layer0_outputs(1303) <= b and not a;
    layer0_outputs(1304) <= not (a or b);
    layer0_outputs(1305) <= a;
    layer0_outputs(1306) <= a xor b;
    layer0_outputs(1307) <= not b or a;
    layer0_outputs(1308) <= not (a or b);
    layer0_outputs(1309) <= a or b;
    layer0_outputs(1310) <= not b;
    layer0_outputs(1311) <= a and not b;
    layer0_outputs(1312) <= b and not a;
    layer0_outputs(1313) <= not b;
    layer0_outputs(1314) <= b;
    layer0_outputs(1315) <= not (a xor b);
    layer0_outputs(1316) <= b and not a;
    layer0_outputs(1317) <= not (a xor b);
    layer0_outputs(1318) <= b;
    layer0_outputs(1319) <= not b;
    layer0_outputs(1320) <= a or b;
    layer0_outputs(1321) <= a or b;
    layer0_outputs(1322) <= a or b;
    layer0_outputs(1323) <= b and not a;
    layer0_outputs(1324) <= b;
    layer0_outputs(1325) <= a and b;
    layer0_outputs(1326) <= a or b;
    layer0_outputs(1327) <= b;
    layer0_outputs(1328) <= not a;
    layer0_outputs(1329) <= not b or a;
    layer0_outputs(1330) <= b;
    layer0_outputs(1331) <= not (a or b);
    layer0_outputs(1332) <= not b;
    layer0_outputs(1333) <= a or b;
    layer0_outputs(1334) <= b;
    layer0_outputs(1335) <= b and not a;
    layer0_outputs(1336) <= a xor b;
    layer0_outputs(1337) <= not b or a;
    layer0_outputs(1338) <= a xor b;
    layer0_outputs(1339) <= not a or b;
    layer0_outputs(1340) <= not a;
    layer0_outputs(1341) <= not (a xor b);
    layer0_outputs(1342) <= a and not b;
    layer0_outputs(1343) <= not (a xor b);
    layer0_outputs(1344) <= a and not b;
    layer0_outputs(1345) <= not (a or b);
    layer0_outputs(1346) <= not (a and b);
    layer0_outputs(1347) <= not b or a;
    layer0_outputs(1348) <= a or b;
    layer0_outputs(1349) <= a or b;
    layer0_outputs(1350) <= 1'b1;
    layer0_outputs(1351) <= a or b;
    layer0_outputs(1352) <= a;
    layer0_outputs(1353) <= a and not b;
    layer0_outputs(1354) <= not (a xor b);
    layer0_outputs(1355) <= not b;
    layer0_outputs(1356) <= b and not a;
    layer0_outputs(1357) <= b;
    layer0_outputs(1358) <= b;
    layer0_outputs(1359) <= b;
    layer0_outputs(1360) <= not (a xor b);
    layer0_outputs(1361) <= not (a or b);
    layer0_outputs(1362) <= not (a xor b);
    layer0_outputs(1363) <= a;
    layer0_outputs(1364) <= not (a or b);
    layer0_outputs(1365) <= a or b;
    layer0_outputs(1366) <= not a or b;
    layer0_outputs(1367) <= b and not a;
    layer0_outputs(1368) <= not b or a;
    layer0_outputs(1369) <= not a or b;
    layer0_outputs(1370) <= a or b;
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= 1'b1;
    layer0_outputs(1373) <= not (a and b);
    layer0_outputs(1374) <= not a;
    layer0_outputs(1375) <= a;
    layer0_outputs(1376) <= not a;
    layer0_outputs(1377) <= a and not b;
    layer0_outputs(1378) <= b and not a;
    layer0_outputs(1379) <= not (a xor b);
    layer0_outputs(1380) <= not b or a;
    layer0_outputs(1381) <= a and not b;
    layer0_outputs(1382) <= b;
    layer0_outputs(1383) <= not a;
    layer0_outputs(1384) <= not (a or b);
    layer0_outputs(1385) <= a or b;
    layer0_outputs(1386) <= a and not b;
    layer0_outputs(1387) <= 1'b1;
    layer0_outputs(1388) <= a xor b;
    layer0_outputs(1389) <= not (a or b);
    layer0_outputs(1390) <= a;
    layer0_outputs(1391) <= b;
    layer0_outputs(1392) <= a and not b;
    layer0_outputs(1393) <= a;
    layer0_outputs(1394) <= not (a or b);
    layer0_outputs(1395) <= not (a or b);
    layer0_outputs(1396) <= not a or b;
    layer0_outputs(1397) <= b and not a;
    layer0_outputs(1398) <= b;
    layer0_outputs(1399) <= a;
    layer0_outputs(1400) <= b and not a;
    layer0_outputs(1401) <= not (a xor b);
    layer0_outputs(1402) <= not (a or b);
    layer0_outputs(1403) <= b and not a;
    layer0_outputs(1404) <= a or b;
    layer0_outputs(1405) <= not a or b;
    layer0_outputs(1406) <= not (a or b);
    layer0_outputs(1407) <= not (a xor b);
    layer0_outputs(1408) <= b and not a;
    layer0_outputs(1409) <= 1'b0;
    layer0_outputs(1410) <= not (a xor b);
    layer0_outputs(1411) <= not (a or b);
    layer0_outputs(1412) <= a and b;
    layer0_outputs(1413) <= a;
    layer0_outputs(1414) <= not a;
    layer0_outputs(1415) <= b;
    layer0_outputs(1416) <= a;
    layer0_outputs(1417) <= a;
    layer0_outputs(1418) <= not (a xor b);
    layer0_outputs(1419) <= not a;
    layer0_outputs(1420) <= a or b;
    layer0_outputs(1421) <= not (a or b);
    layer0_outputs(1422) <= not (a or b);
    layer0_outputs(1423) <= not b;
    layer0_outputs(1424) <= a;
    layer0_outputs(1425) <= not b;
    layer0_outputs(1426) <= not (a xor b);
    layer0_outputs(1427) <= a;
    layer0_outputs(1428) <= b and not a;
    layer0_outputs(1429) <= not b or a;
    layer0_outputs(1430) <= b;
    layer0_outputs(1431) <= not (a or b);
    layer0_outputs(1432) <= not (a or b);
    layer0_outputs(1433) <= b;
    layer0_outputs(1434) <= a;
    layer0_outputs(1435) <= 1'b0;
    layer0_outputs(1436) <= a and not b;
    layer0_outputs(1437) <= a;
    layer0_outputs(1438) <= a or b;
    layer0_outputs(1439) <= a xor b;
    layer0_outputs(1440) <= not b or a;
    layer0_outputs(1441) <= not a;
    layer0_outputs(1442) <= b and not a;
    layer0_outputs(1443) <= a or b;
    layer0_outputs(1444) <= a and not b;
    layer0_outputs(1445) <= a or b;
    layer0_outputs(1446) <= a and not b;
    layer0_outputs(1447) <= not b;
    layer0_outputs(1448) <= not b or a;
    layer0_outputs(1449) <= not a or b;
    layer0_outputs(1450) <= not (a and b);
    layer0_outputs(1451) <= b;
    layer0_outputs(1452) <= not b or a;
    layer0_outputs(1453) <= a and b;
    layer0_outputs(1454) <= a or b;
    layer0_outputs(1455) <= not b;
    layer0_outputs(1456) <= a xor b;
    layer0_outputs(1457) <= a;
    layer0_outputs(1458) <= a xor b;
    layer0_outputs(1459) <= not (a and b);
    layer0_outputs(1460) <= b and not a;
    layer0_outputs(1461) <= b;
    layer0_outputs(1462) <= b;
    layer0_outputs(1463) <= not (a or b);
    layer0_outputs(1464) <= not (a or b);
    layer0_outputs(1465) <= a and b;
    layer0_outputs(1466) <= a xor b;
    layer0_outputs(1467) <= a or b;
    layer0_outputs(1468) <= 1'b0;
    layer0_outputs(1469) <= not a;
    layer0_outputs(1470) <= not (a or b);
    layer0_outputs(1471) <= not a or b;
    layer0_outputs(1472) <= not a;
    layer0_outputs(1473) <= not a;
    layer0_outputs(1474) <= a and not b;
    layer0_outputs(1475) <= not (a and b);
    layer0_outputs(1476) <= a and b;
    layer0_outputs(1477) <= not (a xor b);
    layer0_outputs(1478) <= a;
    layer0_outputs(1479) <= not (a or b);
    layer0_outputs(1480) <= not a;
    layer0_outputs(1481) <= a;
    layer0_outputs(1482) <= not (a xor b);
    layer0_outputs(1483) <= b;
    layer0_outputs(1484) <= b;
    layer0_outputs(1485) <= not b;
    layer0_outputs(1486) <= not (a and b);
    layer0_outputs(1487) <= 1'b0;
    layer0_outputs(1488) <= a and not b;
    layer0_outputs(1489) <= not (a or b);
    layer0_outputs(1490) <= not (a and b);
    layer0_outputs(1491) <= not (a and b);
    layer0_outputs(1492) <= not (a xor b);
    layer0_outputs(1493) <= 1'b1;
    layer0_outputs(1494) <= a and not b;
    layer0_outputs(1495) <= not (a and b);
    layer0_outputs(1496) <= not a;
    layer0_outputs(1497) <= not a;
    layer0_outputs(1498) <= not (a or b);
    layer0_outputs(1499) <= not (a or b);
    layer0_outputs(1500) <= not (a xor b);
    layer0_outputs(1501) <= not b;
    layer0_outputs(1502) <= not b;
    layer0_outputs(1503) <= 1'b1;
    layer0_outputs(1504) <= a xor b;
    layer0_outputs(1505) <= a or b;
    layer0_outputs(1506) <= not (a and b);
    layer0_outputs(1507) <= not (a or b);
    layer0_outputs(1508) <= b and not a;
    layer0_outputs(1509) <= not a;
    layer0_outputs(1510) <= not (a or b);
    layer0_outputs(1511) <= not (a xor b);
    layer0_outputs(1512) <= not a or b;
    layer0_outputs(1513) <= a xor b;
    layer0_outputs(1514) <= a or b;
    layer0_outputs(1515) <= a and b;
    layer0_outputs(1516) <= not a;
    layer0_outputs(1517) <= b and not a;
    layer0_outputs(1518) <= a and not b;
    layer0_outputs(1519) <= not b or a;
    layer0_outputs(1520) <= not (a or b);
    layer0_outputs(1521) <= not (a or b);
    layer0_outputs(1522) <= a xor b;
    layer0_outputs(1523) <= a xor b;
    layer0_outputs(1524) <= not b;
    layer0_outputs(1525) <= not (a xor b);
    layer0_outputs(1526) <= not a;
    layer0_outputs(1527) <= a;
    layer0_outputs(1528) <= a and not b;
    layer0_outputs(1529) <= not b or a;
    layer0_outputs(1530) <= not b or a;
    layer0_outputs(1531) <= not (a or b);
    layer0_outputs(1532) <= not (a or b);
    layer0_outputs(1533) <= not (a xor b);
    layer0_outputs(1534) <= not b or a;
    layer0_outputs(1535) <= a;
    layer0_outputs(1536) <= not a;
    layer0_outputs(1537) <= a or b;
    layer0_outputs(1538) <= 1'b0;
    layer0_outputs(1539) <= not (a or b);
    layer0_outputs(1540) <= a or b;
    layer0_outputs(1541) <= b;
    layer0_outputs(1542) <= not (a or b);
    layer0_outputs(1543) <= b and not a;
    layer0_outputs(1544) <= a or b;
    layer0_outputs(1545) <= b;
    layer0_outputs(1546) <= b;
    layer0_outputs(1547) <= not a;
    layer0_outputs(1548) <= a and b;
    layer0_outputs(1549) <= not b;
    layer0_outputs(1550) <= a or b;
    layer0_outputs(1551) <= not (a or b);
    layer0_outputs(1552) <= not b;
    layer0_outputs(1553) <= a xor b;
    layer0_outputs(1554) <= a and not b;
    layer0_outputs(1555) <= not a or b;
    layer0_outputs(1556) <= b;
    layer0_outputs(1557) <= a;
    layer0_outputs(1558) <= a and not b;
    layer0_outputs(1559) <= not (a xor b);
    layer0_outputs(1560) <= b;
    layer0_outputs(1561) <= not a;
    layer0_outputs(1562) <= not (a or b);
    layer0_outputs(1563) <= b;
    layer0_outputs(1564) <= a or b;
    layer0_outputs(1565) <= not (a or b);
    layer0_outputs(1566) <= not b or a;
    layer0_outputs(1567) <= a and not b;
    layer0_outputs(1568) <= a and not b;
    layer0_outputs(1569) <= b and not a;
    layer0_outputs(1570) <= not b;
    layer0_outputs(1571) <= not (a and b);
    layer0_outputs(1572) <= not a;
    layer0_outputs(1573) <= a xor b;
    layer0_outputs(1574) <= b and not a;
    layer0_outputs(1575) <= a;
    layer0_outputs(1576) <= not a or b;
    layer0_outputs(1577) <= a xor b;
    layer0_outputs(1578) <= b and not a;
    layer0_outputs(1579) <= not (a or b);
    layer0_outputs(1580) <= not b or a;
    layer0_outputs(1581) <= b;
    layer0_outputs(1582) <= b;
    layer0_outputs(1583) <= b;
    layer0_outputs(1584) <= not a;
    layer0_outputs(1585) <= not (a xor b);
    layer0_outputs(1586) <= not (a or b);
    layer0_outputs(1587) <= not b;
    layer0_outputs(1588) <= not b or a;
    layer0_outputs(1589) <= not (a xor b);
    layer0_outputs(1590) <= a or b;
    layer0_outputs(1591) <= a;
    layer0_outputs(1592) <= not (a or b);
    layer0_outputs(1593) <= b and not a;
    layer0_outputs(1594) <= a or b;
    layer0_outputs(1595) <= not (a or b);
    layer0_outputs(1596) <= not b or a;
    layer0_outputs(1597) <= a or b;
    layer0_outputs(1598) <= a or b;
    layer0_outputs(1599) <= not (a or b);
    layer0_outputs(1600) <= not (a or b);
    layer0_outputs(1601) <= not a or b;
    layer0_outputs(1602) <= 1'b0;
    layer0_outputs(1603) <= not a or b;
    layer0_outputs(1604) <= a xor b;
    layer0_outputs(1605) <= not b or a;
    layer0_outputs(1606) <= not a or b;
    layer0_outputs(1607) <= not (a or b);
    layer0_outputs(1608) <= 1'b0;
    layer0_outputs(1609) <= 1'b0;
    layer0_outputs(1610) <= not b or a;
    layer0_outputs(1611) <= not a or b;
    layer0_outputs(1612) <= a;
    layer0_outputs(1613) <= not b or a;
    layer0_outputs(1614) <= 1'b0;
    layer0_outputs(1615) <= a;
    layer0_outputs(1616) <= a;
    layer0_outputs(1617) <= not b or a;
    layer0_outputs(1618) <= a or b;
    layer0_outputs(1619) <= not (a or b);
    layer0_outputs(1620) <= a xor b;
    layer0_outputs(1621) <= not b or a;
    layer0_outputs(1622) <= not a;
    layer0_outputs(1623) <= a or b;
    layer0_outputs(1624) <= not (a or b);
    layer0_outputs(1625) <= a and b;
    layer0_outputs(1626) <= not b or a;
    layer0_outputs(1627) <= not a;
    layer0_outputs(1628) <= not (a or b);
    layer0_outputs(1629) <= a xor b;
    layer0_outputs(1630) <= a and not b;
    layer0_outputs(1631) <= not a;
    layer0_outputs(1632) <= b and not a;
    layer0_outputs(1633) <= not a;
    layer0_outputs(1634) <= not b or a;
    layer0_outputs(1635) <= not b or a;
    layer0_outputs(1636) <= a;
    layer0_outputs(1637) <= not a;
    layer0_outputs(1638) <= not a or b;
    layer0_outputs(1639) <= 1'b0;
    layer0_outputs(1640) <= not b or a;
    layer0_outputs(1641) <= not (a or b);
    layer0_outputs(1642) <= a xor b;
    layer0_outputs(1643) <= a;
    layer0_outputs(1644) <= a xor b;
    layer0_outputs(1645) <= not (a or b);
    layer0_outputs(1646) <= a and not b;
    layer0_outputs(1647) <= a or b;
    layer0_outputs(1648) <= not a;
    layer0_outputs(1649) <= not b;
    layer0_outputs(1650) <= a xor b;
    layer0_outputs(1651) <= a or b;
    layer0_outputs(1652) <= a xor b;
    layer0_outputs(1653) <= a;
    layer0_outputs(1654) <= not b or a;
    layer0_outputs(1655) <= not a or b;
    layer0_outputs(1656) <= a xor b;
    layer0_outputs(1657) <= not (a or b);
    layer0_outputs(1658) <= b;
    layer0_outputs(1659) <= a and not b;
    layer0_outputs(1660) <= a;
    layer0_outputs(1661) <= b and not a;
    layer0_outputs(1662) <= a and b;
    layer0_outputs(1663) <= not b or a;
    layer0_outputs(1664) <= b;
    layer0_outputs(1665) <= a;
    layer0_outputs(1666) <= b;
    layer0_outputs(1667) <= not b;
    layer0_outputs(1668) <= not b;
    layer0_outputs(1669) <= not a;
    layer0_outputs(1670) <= b;
    layer0_outputs(1671) <= not (a and b);
    layer0_outputs(1672) <= not b or a;
    layer0_outputs(1673) <= b;
    layer0_outputs(1674) <= not (a xor b);
    layer0_outputs(1675) <= a or b;
    layer0_outputs(1676) <= b;
    layer0_outputs(1677) <= not (a or b);
    layer0_outputs(1678) <= a or b;
    layer0_outputs(1679) <= b and not a;
    layer0_outputs(1680) <= not b or a;
    layer0_outputs(1681) <= not a;
    layer0_outputs(1682) <= not a or b;
    layer0_outputs(1683) <= a or b;
    layer0_outputs(1684) <= 1'b1;
    layer0_outputs(1685) <= not (a or b);
    layer0_outputs(1686) <= not b;
    layer0_outputs(1687) <= not (a xor b);
    layer0_outputs(1688) <= a and b;
    layer0_outputs(1689) <= b;
    layer0_outputs(1690) <= not (a xor b);
    layer0_outputs(1691) <= a and not b;
    layer0_outputs(1692) <= a;
    layer0_outputs(1693) <= not (a xor b);
    layer0_outputs(1694) <= a xor b;
    layer0_outputs(1695) <= not a or b;
    layer0_outputs(1696) <= a or b;
    layer0_outputs(1697) <= not a or b;
    layer0_outputs(1698) <= a and not b;
    layer0_outputs(1699) <= not a;
    layer0_outputs(1700) <= not b;
    layer0_outputs(1701) <= b;
    layer0_outputs(1702) <= b;
    layer0_outputs(1703) <= 1'b0;
    layer0_outputs(1704) <= a;
    layer0_outputs(1705) <= a;
    layer0_outputs(1706) <= not (a xor b);
    layer0_outputs(1707) <= a;
    layer0_outputs(1708) <= not (a or b);
    layer0_outputs(1709) <= b;
    layer0_outputs(1710) <= a xor b;
    layer0_outputs(1711) <= a and b;
    layer0_outputs(1712) <= not a or b;
    layer0_outputs(1713) <= not b;
    layer0_outputs(1714) <= not (a and b);
    layer0_outputs(1715) <= 1'b1;
    layer0_outputs(1716) <= not (a xor b);
    layer0_outputs(1717) <= not a;
    layer0_outputs(1718) <= not a;
    layer0_outputs(1719) <= a xor b;
    layer0_outputs(1720) <= not (a or b);
    layer0_outputs(1721) <= b;
    layer0_outputs(1722) <= a and not b;
    layer0_outputs(1723) <= b;
    layer0_outputs(1724) <= b;
    layer0_outputs(1725) <= not a or b;
    layer0_outputs(1726) <= not (a and b);
    layer0_outputs(1727) <= not b or a;
    layer0_outputs(1728) <= b and not a;
    layer0_outputs(1729) <= a xor b;
    layer0_outputs(1730) <= a;
    layer0_outputs(1731) <= not a or b;
    layer0_outputs(1732) <= not (a xor b);
    layer0_outputs(1733) <= not b or a;
    layer0_outputs(1734) <= not b or a;
    layer0_outputs(1735) <= not (a or b);
    layer0_outputs(1736) <= b and not a;
    layer0_outputs(1737) <= not b;
    layer0_outputs(1738) <= a xor b;
    layer0_outputs(1739) <= not (a or b);
    layer0_outputs(1740) <= b;
    layer0_outputs(1741) <= b and not a;
    layer0_outputs(1742) <= a and b;
    layer0_outputs(1743) <= a or b;
    layer0_outputs(1744) <= a or b;
    layer0_outputs(1745) <= not a;
    layer0_outputs(1746) <= not (a or b);
    layer0_outputs(1747) <= not b or a;
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= b and not a;
    layer0_outputs(1750) <= b;
    layer0_outputs(1751) <= a or b;
    layer0_outputs(1752) <= not (a or b);
    layer0_outputs(1753) <= not b;
    layer0_outputs(1754) <= not a;
    layer0_outputs(1755) <= not a;
    layer0_outputs(1756) <= a and not b;
    layer0_outputs(1757) <= not a or b;
    layer0_outputs(1758) <= not a;
    layer0_outputs(1759) <= b;
    layer0_outputs(1760) <= not (a and b);
    layer0_outputs(1761) <= not (a or b);
    layer0_outputs(1762) <= not b;
    layer0_outputs(1763) <= a;
    layer0_outputs(1764) <= a or b;
    layer0_outputs(1765) <= a and not b;
    layer0_outputs(1766) <= not (a or b);
    layer0_outputs(1767) <= a or b;
    layer0_outputs(1768) <= a or b;
    layer0_outputs(1769) <= not b;
    layer0_outputs(1770) <= a;
    layer0_outputs(1771) <= b;
    layer0_outputs(1772) <= not b or a;
    layer0_outputs(1773) <= not b;
    layer0_outputs(1774) <= b and not a;
    layer0_outputs(1775) <= not a or b;
    layer0_outputs(1776) <= 1'b0;
    layer0_outputs(1777) <= not b or a;
    layer0_outputs(1778) <= a xor b;
    layer0_outputs(1779) <= a and b;
    layer0_outputs(1780) <= a or b;
    layer0_outputs(1781) <= a or b;
    layer0_outputs(1782) <= a or b;
    layer0_outputs(1783) <= not (a or b);
    layer0_outputs(1784) <= b;
    layer0_outputs(1785) <= not a;
    layer0_outputs(1786) <= not (a xor b);
    layer0_outputs(1787) <= b and not a;
    layer0_outputs(1788) <= b;
    layer0_outputs(1789) <= not (a xor b);
    layer0_outputs(1790) <= not b;
    layer0_outputs(1791) <= not (a or b);
    layer0_outputs(1792) <= a xor b;
    layer0_outputs(1793) <= not b or a;
    layer0_outputs(1794) <= a and not b;
    layer0_outputs(1795) <= not (a and b);
    layer0_outputs(1796) <= not a or b;
    layer0_outputs(1797) <= not b;
    layer0_outputs(1798) <= not (a or b);
    layer0_outputs(1799) <= a or b;
    layer0_outputs(1800) <= b and not a;
    layer0_outputs(1801) <= not (a xor b);
    layer0_outputs(1802) <= 1'b0;
    layer0_outputs(1803) <= not b;
    layer0_outputs(1804) <= a or b;
    layer0_outputs(1805) <= a or b;
    layer0_outputs(1806) <= a and not b;
    layer0_outputs(1807) <= a or b;
    layer0_outputs(1808) <= not b or a;
    layer0_outputs(1809) <= a and not b;
    layer0_outputs(1810) <= a;
    layer0_outputs(1811) <= a or b;
    layer0_outputs(1812) <= not (a or b);
    layer0_outputs(1813) <= not (a or b);
    layer0_outputs(1814) <= not (a or b);
    layer0_outputs(1815) <= a and not b;
    layer0_outputs(1816) <= not (a or b);
    layer0_outputs(1817) <= a and not b;
    layer0_outputs(1818) <= not (a or b);
    layer0_outputs(1819) <= not (a xor b);
    layer0_outputs(1820) <= a xor b;
    layer0_outputs(1821) <= a or b;
    layer0_outputs(1822) <= not a or b;
    layer0_outputs(1823) <= a or b;
    layer0_outputs(1824) <= not b or a;
    layer0_outputs(1825) <= not (a xor b);
    layer0_outputs(1826) <= b;
    layer0_outputs(1827) <= a or b;
    layer0_outputs(1828) <= b;
    layer0_outputs(1829) <= not (a xor b);
    layer0_outputs(1830) <= not (a or b);
    layer0_outputs(1831) <= not (a xor b);
    layer0_outputs(1832) <= not (a or b);
    layer0_outputs(1833) <= a or b;
    layer0_outputs(1834) <= a xor b;
    layer0_outputs(1835) <= b and not a;
    layer0_outputs(1836) <= a;
    layer0_outputs(1837) <= not a;
    layer0_outputs(1838) <= a and b;
    layer0_outputs(1839) <= a and not b;
    layer0_outputs(1840) <= a;
    layer0_outputs(1841) <= not b;
    layer0_outputs(1842) <= a;
    layer0_outputs(1843) <= b;
    layer0_outputs(1844) <= not (a or b);
    layer0_outputs(1845) <= not (a or b);
    layer0_outputs(1846) <= a;
    layer0_outputs(1847) <= not b;
    layer0_outputs(1848) <= not b or a;
    layer0_outputs(1849) <= not b;
    layer0_outputs(1850) <= b;
    layer0_outputs(1851) <= not a;
    layer0_outputs(1852) <= not a or b;
    layer0_outputs(1853) <= a or b;
    layer0_outputs(1854) <= not b;
    layer0_outputs(1855) <= not (a or b);
    layer0_outputs(1856) <= a;
    layer0_outputs(1857) <= not b;
    layer0_outputs(1858) <= a or b;
    layer0_outputs(1859) <= b and not a;
    layer0_outputs(1860) <= not (a xor b);
    layer0_outputs(1861) <= b;
    layer0_outputs(1862) <= not a;
    layer0_outputs(1863) <= not b;
    layer0_outputs(1864) <= a and not b;
    layer0_outputs(1865) <= not (a and b);
    layer0_outputs(1866) <= b and not a;
    layer0_outputs(1867) <= not a or b;
    layer0_outputs(1868) <= a or b;
    layer0_outputs(1869) <= not (a or b);
    layer0_outputs(1870) <= not a;
    layer0_outputs(1871) <= b and not a;
    layer0_outputs(1872) <= not a or b;
    layer0_outputs(1873) <= not (a or b);
    layer0_outputs(1874) <= not a;
    layer0_outputs(1875) <= not (a xor b);
    layer0_outputs(1876) <= not b;
    layer0_outputs(1877) <= b;
    layer0_outputs(1878) <= 1'b0;
    layer0_outputs(1879) <= not a;
    layer0_outputs(1880) <= 1'b1;
    layer0_outputs(1881) <= not (a or b);
    layer0_outputs(1882) <= not b;
    layer0_outputs(1883) <= b;
    layer0_outputs(1884) <= not (a or b);
    layer0_outputs(1885) <= a;
    layer0_outputs(1886) <= not a;
    layer0_outputs(1887) <= a or b;
    layer0_outputs(1888) <= not (a and b);
    layer0_outputs(1889) <= a;
    layer0_outputs(1890) <= b;
    layer0_outputs(1891) <= not (a or b);
    layer0_outputs(1892) <= a or b;
    layer0_outputs(1893) <= not (a or b);
    layer0_outputs(1894) <= not b;
    layer0_outputs(1895) <= not (a or b);
    layer0_outputs(1896) <= b and not a;
    layer0_outputs(1897) <= b and not a;
    layer0_outputs(1898) <= not a;
    layer0_outputs(1899) <= b and not a;
    layer0_outputs(1900) <= not (a and b);
    layer0_outputs(1901) <= not a;
    layer0_outputs(1902) <= not (a xor b);
    layer0_outputs(1903) <= not a or b;
    layer0_outputs(1904) <= a xor b;
    layer0_outputs(1905) <= a;
    layer0_outputs(1906) <= a xor b;
    layer0_outputs(1907) <= not a;
    layer0_outputs(1908) <= not (a xor b);
    layer0_outputs(1909) <= a and not b;
    layer0_outputs(1910) <= a and not b;
    layer0_outputs(1911) <= not a;
    layer0_outputs(1912) <= not (a xor b);
    layer0_outputs(1913) <= not (a xor b);
    layer0_outputs(1914) <= not b;
    layer0_outputs(1915) <= a xor b;
    layer0_outputs(1916) <= a;
    layer0_outputs(1917) <= not (a xor b);
    layer0_outputs(1918) <= b and not a;
    layer0_outputs(1919) <= b;
    layer0_outputs(1920) <= not b;
    layer0_outputs(1921) <= not (a or b);
    layer0_outputs(1922) <= a and b;
    layer0_outputs(1923) <= not (a and b);
    layer0_outputs(1924) <= a or b;
    layer0_outputs(1925) <= not (a or b);
    layer0_outputs(1926) <= b and not a;
    layer0_outputs(1927) <= not a;
    layer0_outputs(1928) <= not b or a;
    layer0_outputs(1929) <= a xor b;
    layer0_outputs(1930) <= b and not a;
    layer0_outputs(1931) <= a or b;
    layer0_outputs(1932) <= a or b;
    layer0_outputs(1933) <= a xor b;
    layer0_outputs(1934) <= not b or a;
    layer0_outputs(1935) <= a or b;
    layer0_outputs(1936) <= not a;
    layer0_outputs(1937) <= b;
    layer0_outputs(1938) <= not b;
    layer0_outputs(1939) <= a xor b;
    layer0_outputs(1940) <= a xor b;
    layer0_outputs(1941) <= a and b;
    layer0_outputs(1942) <= not a;
    layer0_outputs(1943) <= a and not b;
    layer0_outputs(1944) <= not a;
    layer0_outputs(1945) <= not b;
    layer0_outputs(1946) <= not a;
    layer0_outputs(1947) <= b;
    layer0_outputs(1948) <= not (a xor b);
    layer0_outputs(1949) <= not a;
    layer0_outputs(1950) <= not (a xor b);
    layer0_outputs(1951) <= not b or a;
    layer0_outputs(1952) <= a or b;
    layer0_outputs(1953) <= b and not a;
    layer0_outputs(1954) <= a or b;
    layer0_outputs(1955) <= not (a xor b);
    layer0_outputs(1956) <= b;
    layer0_outputs(1957) <= b;
    layer0_outputs(1958) <= not b;
    layer0_outputs(1959) <= a and not b;
    layer0_outputs(1960) <= b and not a;
    layer0_outputs(1961) <= not (a xor b);
    layer0_outputs(1962) <= a or b;
    layer0_outputs(1963) <= a or b;
    layer0_outputs(1964) <= not a or b;
    layer0_outputs(1965) <= not a;
    layer0_outputs(1966) <= not (a or b);
    layer0_outputs(1967) <= not a or b;
    layer0_outputs(1968) <= a;
    layer0_outputs(1969) <= not a;
    layer0_outputs(1970) <= not (a xor b);
    layer0_outputs(1971) <= not (a or b);
    layer0_outputs(1972) <= not (a or b);
    layer0_outputs(1973) <= b and not a;
    layer0_outputs(1974) <= not a;
    layer0_outputs(1975) <= a or b;
    layer0_outputs(1976) <= not b;
    layer0_outputs(1977) <= not (a or b);
    layer0_outputs(1978) <= not (a or b);
    layer0_outputs(1979) <= not (a or b);
    layer0_outputs(1980) <= a;
    layer0_outputs(1981) <= a and not b;
    layer0_outputs(1982) <= not (a xor b);
    layer0_outputs(1983) <= not (a or b);
    layer0_outputs(1984) <= a;
    layer0_outputs(1985) <= not a or b;
    layer0_outputs(1986) <= a and not b;
    layer0_outputs(1987) <= a;
    layer0_outputs(1988) <= not (a or b);
    layer0_outputs(1989) <= a or b;
    layer0_outputs(1990) <= not a or b;
    layer0_outputs(1991) <= not (a and b);
    layer0_outputs(1992) <= not b;
    layer0_outputs(1993) <= a and not b;
    layer0_outputs(1994) <= a or b;
    layer0_outputs(1995) <= a or b;
    layer0_outputs(1996) <= not b;
    layer0_outputs(1997) <= not (a xor b);
    layer0_outputs(1998) <= a and not b;
    layer0_outputs(1999) <= not (a or b);
    layer0_outputs(2000) <= b;
    layer0_outputs(2001) <= a or b;
    layer0_outputs(2002) <= a and not b;
    layer0_outputs(2003) <= not b or a;
    layer0_outputs(2004) <= not a or b;
    layer0_outputs(2005) <= not a;
    layer0_outputs(2006) <= not b;
    layer0_outputs(2007) <= 1'b0;
    layer0_outputs(2008) <= a and not b;
    layer0_outputs(2009) <= a and not b;
    layer0_outputs(2010) <= not (a and b);
    layer0_outputs(2011) <= b and not a;
    layer0_outputs(2012) <= 1'b0;
    layer0_outputs(2013) <= a or b;
    layer0_outputs(2014) <= b and not a;
    layer0_outputs(2015) <= a;
    layer0_outputs(2016) <= a or b;
    layer0_outputs(2017) <= a and b;
    layer0_outputs(2018) <= a or b;
    layer0_outputs(2019) <= b;
    layer0_outputs(2020) <= not (a or b);
    layer0_outputs(2021) <= not b;
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= a;
    layer0_outputs(2024) <= not (a or b);
    layer0_outputs(2025) <= a or b;
    layer0_outputs(2026) <= a and not b;
    layer0_outputs(2027) <= not b;
    layer0_outputs(2028) <= a and not b;
    layer0_outputs(2029) <= a or b;
    layer0_outputs(2030) <= not b or a;
    layer0_outputs(2031) <= not a;
    layer0_outputs(2032) <= not a or b;
    layer0_outputs(2033) <= b;
    layer0_outputs(2034) <= not a or b;
    layer0_outputs(2035) <= a;
    layer0_outputs(2036) <= not (a or b);
    layer0_outputs(2037) <= not b;
    layer0_outputs(2038) <= a;
    layer0_outputs(2039) <= not (a or b);
    layer0_outputs(2040) <= not a;
    layer0_outputs(2041) <= not (a xor b);
    layer0_outputs(2042) <= not b;
    layer0_outputs(2043) <= a or b;
    layer0_outputs(2044) <= a;
    layer0_outputs(2045) <= not a;
    layer0_outputs(2046) <= not (a or b);
    layer0_outputs(2047) <= not a or b;
    layer0_outputs(2048) <= a;
    layer0_outputs(2049) <= not (a or b);
    layer0_outputs(2050) <= not a;
    layer0_outputs(2051) <= not a;
    layer0_outputs(2052) <= b and not a;
    layer0_outputs(2053) <= a or b;
    layer0_outputs(2054) <= 1'b1;
    layer0_outputs(2055) <= not (a xor b);
    layer0_outputs(2056) <= not b;
    layer0_outputs(2057) <= a or b;
    layer0_outputs(2058) <= a xor b;
    layer0_outputs(2059) <= not b or a;
    layer0_outputs(2060) <= a xor b;
    layer0_outputs(2061) <= not a;
    layer0_outputs(2062) <= not a or b;
    layer0_outputs(2063) <= b;
    layer0_outputs(2064) <= a;
    layer0_outputs(2065) <= not b or a;
    layer0_outputs(2066) <= a and not b;
    layer0_outputs(2067) <= a and not b;
    layer0_outputs(2068) <= 1'b0;
    layer0_outputs(2069) <= b and not a;
    layer0_outputs(2070) <= not b or a;
    layer0_outputs(2071) <= not (a xor b);
    layer0_outputs(2072) <= not (a xor b);
    layer0_outputs(2073) <= not b;
    layer0_outputs(2074) <= b;
    layer0_outputs(2075) <= not (a or b);
    layer0_outputs(2076) <= a or b;
    layer0_outputs(2077) <= a xor b;
    layer0_outputs(2078) <= b;
    layer0_outputs(2079) <= a;
    layer0_outputs(2080) <= 1'b1;
    layer0_outputs(2081) <= not b or a;
    layer0_outputs(2082) <= b and not a;
    layer0_outputs(2083) <= a and b;
    layer0_outputs(2084) <= a xor b;
    layer0_outputs(2085) <= not (a or b);
    layer0_outputs(2086) <= a or b;
    layer0_outputs(2087) <= not (a or b);
    layer0_outputs(2088) <= a xor b;
    layer0_outputs(2089) <= a xor b;
    layer0_outputs(2090) <= b and not a;
    layer0_outputs(2091) <= not (a xor b);
    layer0_outputs(2092) <= not (a or b);
    layer0_outputs(2093) <= b;
    layer0_outputs(2094) <= not b or a;
    layer0_outputs(2095) <= not b or a;
    layer0_outputs(2096) <= not (a xor b);
    layer0_outputs(2097) <= not a;
    layer0_outputs(2098) <= a;
    layer0_outputs(2099) <= a and not b;
    layer0_outputs(2100) <= b;
    layer0_outputs(2101) <= not (a or b);
    layer0_outputs(2102) <= not a;
    layer0_outputs(2103) <= a or b;
    layer0_outputs(2104) <= a and b;
    layer0_outputs(2105) <= 1'b0;
    layer0_outputs(2106) <= a or b;
    layer0_outputs(2107) <= a and not b;
    layer0_outputs(2108) <= a;
    layer0_outputs(2109) <= a or b;
    layer0_outputs(2110) <= not a;
    layer0_outputs(2111) <= not a;
    layer0_outputs(2112) <= 1'b1;
    layer0_outputs(2113) <= not (a xor b);
    layer0_outputs(2114) <= b and not a;
    layer0_outputs(2115) <= not b;
    layer0_outputs(2116) <= b and not a;
    layer0_outputs(2117) <= not a or b;
    layer0_outputs(2118) <= not a or b;
    layer0_outputs(2119) <= b and not a;
    layer0_outputs(2120) <= not a or b;
    layer0_outputs(2121) <= a or b;
    layer0_outputs(2122) <= a or b;
    layer0_outputs(2123) <= a;
    layer0_outputs(2124) <= 1'b1;
    layer0_outputs(2125) <= not b or a;
    layer0_outputs(2126) <= not (a and b);
    layer0_outputs(2127) <= not b;
    layer0_outputs(2128) <= not a;
    layer0_outputs(2129) <= a xor b;
    layer0_outputs(2130) <= not (a xor b);
    layer0_outputs(2131) <= a or b;
    layer0_outputs(2132) <= not (a or b);
    layer0_outputs(2133) <= 1'b1;
    layer0_outputs(2134) <= b and not a;
    layer0_outputs(2135) <= not (a xor b);
    layer0_outputs(2136) <= not b;
    layer0_outputs(2137) <= b and not a;
    layer0_outputs(2138) <= not b;
    layer0_outputs(2139) <= 1'b1;
    layer0_outputs(2140) <= a or b;
    layer0_outputs(2141) <= a xor b;
    layer0_outputs(2142) <= a;
    layer0_outputs(2143) <= a;
    layer0_outputs(2144) <= not (a or b);
    layer0_outputs(2145) <= not (a or b);
    layer0_outputs(2146) <= not (a or b);
    layer0_outputs(2147) <= a and not b;
    layer0_outputs(2148) <= not a;
    layer0_outputs(2149) <= a;
    layer0_outputs(2150) <= a or b;
    layer0_outputs(2151) <= b;
    layer0_outputs(2152) <= not (a xor b);
    layer0_outputs(2153) <= a xor b;
    layer0_outputs(2154) <= not a or b;
    layer0_outputs(2155) <= a or b;
    layer0_outputs(2156) <= not (a xor b);
    layer0_outputs(2157) <= not b;
    layer0_outputs(2158) <= b;
    layer0_outputs(2159) <= not (a or b);
    layer0_outputs(2160) <= a;
    layer0_outputs(2161) <= a and not b;
    layer0_outputs(2162) <= not a or b;
    layer0_outputs(2163) <= not (a or b);
    layer0_outputs(2164) <= a;
    layer0_outputs(2165) <= not (a or b);
    layer0_outputs(2166) <= a xor b;
    layer0_outputs(2167) <= a or b;
    layer0_outputs(2168) <= not a or b;
    layer0_outputs(2169) <= not (a or b);
    layer0_outputs(2170) <= not a or b;
    layer0_outputs(2171) <= not b;
    layer0_outputs(2172) <= 1'b0;
    layer0_outputs(2173) <= a or b;
    layer0_outputs(2174) <= not a or b;
    layer0_outputs(2175) <= 1'b1;
    layer0_outputs(2176) <= a xor b;
    layer0_outputs(2177) <= not b;
    layer0_outputs(2178) <= not a;
    layer0_outputs(2179) <= b;
    layer0_outputs(2180) <= not (a xor b);
    layer0_outputs(2181) <= not b or a;
    layer0_outputs(2182) <= b;
    layer0_outputs(2183) <= a or b;
    layer0_outputs(2184) <= a and not b;
    layer0_outputs(2185) <= a;
    layer0_outputs(2186) <= not b or a;
    layer0_outputs(2187) <= a or b;
    layer0_outputs(2188) <= a or b;
    layer0_outputs(2189) <= not (a xor b);
    layer0_outputs(2190) <= not (a xor b);
    layer0_outputs(2191) <= 1'b1;
    layer0_outputs(2192) <= not a;
    layer0_outputs(2193) <= not (a or b);
    layer0_outputs(2194) <= a or b;
    layer0_outputs(2195) <= a xor b;
    layer0_outputs(2196) <= b;
    layer0_outputs(2197) <= not (a or b);
    layer0_outputs(2198) <= not (a and b);
    layer0_outputs(2199) <= not (a or b);
    layer0_outputs(2200) <= a;
    layer0_outputs(2201) <= not (a xor b);
    layer0_outputs(2202) <= a and not b;
    layer0_outputs(2203) <= not (a and b);
    layer0_outputs(2204) <= not a;
    layer0_outputs(2205) <= a and not b;
    layer0_outputs(2206) <= not (a xor b);
    layer0_outputs(2207) <= not (a and b);
    layer0_outputs(2208) <= a;
    layer0_outputs(2209) <= a xor b;
    layer0_outputs(2210) <= not (a xor b);
    layer0_outputs(2211) <= not b or a;
    layer0_outputs(2212) <= a xor b;
    layer0_outputs(2213) <= b and not a;
    layer0_outputs(2214) <= b;
    layer0_outputs(2215) <= a xor b;
    layer0_outputs(2216) <= b;
    layer0_outputs(2217) <= b;
    layer0_outputs(2218) <= not b;
    layer0_outputs(2219) <= not (a or b);
    layer0_outputs(2220) <= not a or b;
    layer0_outputs(2221) <= a or b;
    layer0_outputs(2222) <= not (a or b);
    layer0_outputs(2223) <= not b;
    layer0_outputs(2224) <= a or b;
    layer0_outputs(2225) <= 1'b1;
    layer0_outputs(2226) <= not (a or b);
    layer0_outputs(2227) <= 1'b1;
    layer0_outputs(2228) <= b and not a;
    layer0_outputs(2229) <= 1'b1;
    layer0_outputs(2230) <= not (a or b);
    layer0_outputs(2231) <= a xor b;
    layer0_outputs(2232) <= a or b;
    layer0_outputs(2233) <= not a or b;
    layer0_outputs(2234) <= not (a or b);
    layer0_outputs(2235) <= 1'b0;
    layer0_outputs(2236) <= not b or a;
    layer0_outputs(2237) <= a;
    layer0_outputs(2238) <= a xor b;
    layer0_outputs(2239) <= a and b;
    layer0_outputs(2240) <= b and not a;
    layer0_outputs(2241) <= a or b;
    layer0_outputs(2242) <= not a;
    layer0_outputs(2243) <= not b or a;
    layer0_outputs(2244) <= b and not a;
    layer0_outputs(2245) <= 1'b0;
    layer0_outputs(2246) <= not a;
    layer0_outputs(2247) <= a and not b;
    layer0_outputs(2248) <= b and not a;
    layer0_outputs(2249) <= a or b;
    layer0_outputs(2250) <= not a or b;
    layer0_outputs(2251) <= b;
    layer0_outputs(2252) <= not (a xor b);
    layer0_outputs(2253) <= not a;
    layer0_outputs(2254) <= not a or b;
    layer0_outputs(2255) <= a or b;
    layer0_outputs(2256) <= not (a xor b);
    layer0_outputs(2257) <= not b;
    layer0_outputs(2258) <= not (a or b);
    layer0_outputs(2259) <= b;
    layer0_outputs(2260) <= b;
    layer0_outputs(2261) <= not (a xor b);
    layer0_outputs(2262) <= a or b;
    layer0_outputs(2263) <= not (a or b);
    layer0_outputs(2264) <= a and not b;
    layer0_outputs(2265) <= a xor b;
    layer0_outputs(2266) <= not (a or b);
    layer0_outputs(2267) <= not (a or b);
    layer0_outputs(2268) <= not (a or b);
    layer0_outputs(2269) <= b and not a;
    layer0_outputs(2270) <= not b;
    layer0_outputs(2271) <= not b;
    layer0_outputs(2272) <= a;
    layer0_outputs(2273) <= not (a xor b);
    layer0_outputs(2274) <= a and b;
    layer0_outputs(2275) <= 1'b0;
    layer0_outputs(2276) <= a or b;
    layer0_outputs(2277) <= not b;
    layer0_outputs(2278) <= not a;
    layer0_outputs(2279) <= not (a or b);
    layer0_outputs(2280) <= not (a or b);
    layer0_outputs(2281) <= not (a and b);
    layer0_outputs(2282) <= a xor b;
    layer0_outputs(2283) <= b and not a;
    layer0_outputs(2284) <= a and b;
    layer0_outputs(2285) <= b;
    layer0_outputs(2286) <= not (a xor b);
    layer0_outputs(2287) <= a or b;
    layer0_outputs(2288) <= b;
    layer0_outputs(2289) <= a;
    layer0_outputs(2290) <= not (a and b);
    layer0_outputs(2291) <= not b or a;
    layer0_outputs(2292) <= not (a or b);
    layer0_outputs(2293) <= not b;
    layer0_outputs(2294) <= a xor b;
    layer0_outputs(2295) <= a or b;
    layer0_outputs(2296) <= a or b;
    layer0_outputs(2297) <= a or b;
    layer0_outputs(2298) <= not (a or b);
    layer0_outputs(2299) <= not b;
    layer0_outputs(2300) <= not (a or b);
    layer0_outputs(2301) <= b and not a;
    layer0_outputs(2302) <= not a or b;
    layer0_outputs(2303) <= a;
    layer0_outputs(2304) <= not (a or b);
    layer0_outputs(2305) <= not a;
    layer0_outputs(2306) <= b and not a;
    layer0_outputs(2307) <= not b;
    layer0_outputs(2308) <= not b or a;
    layer0_outputs(2309) <= a xor b;
    layer0_outputs(2310) <= a and b;
    layer0_outputs(2311) <= not b;
    layer0_outputs(2312) <= a and not b;
    layer0_outputs(2313) <= not (a or b);
    layer0_outputs(2314) <= a and not b;
    layer0_outputs(2315) <= not (a or b);
    layer0_outputs(2316) <= not a;
    layer0_outputs(2317) <= a;
    layer0_outputs(2318) <= 1'b1;
    layer0_outputs(2319) <= not b;
    layer0_outputs(2320) <= b and not a;
    layer0_outputs(2321) <= not a;
    layer0_outputs(2322) <= b and not a;
    layer0_outputs(2323) <= a or b;
    layer0_outputs(2324) <= b and not a;
    layer0_outputs(2325) <= not (a xor b);
    layer0_outputs(2326) <= a xor b;
    layer0_outputs(2327) <= a or b;
    layer0_outputs(2328) <= not a;
    layer0_outputs(2329) <= not (a or b);
    layer0_outputs(2330) <= not b or a;
    layer0_outputs(2331) <= a or b;
    layer0_outputs(2332) <= a xor b;
    layer0_outputs(2333) <= not b;
    layer0_outputs(2334) <= not (a and b);
    layer0_outputs(2335) <= a xor b;
    layer0_outputs(2336) <= a;
    layer0_outputs(2337) <= a and not b;
    layer0_outputs(2338) <= a and not b;
    layer0_outputs(2339) <= b and not a;
    layer0_outputs(2340) <= a;
    layer0_outputs(2341) <= b and not a;
    layer0_outputs(2342) <= not b;
    layer0_outputs(2343) <= a or b;
    layer0_outputs(2344) <= not b or a;
    layer0_outputs(2345) <= a xor b;
    layer0_outputs(2346) <= 1'b0;
    layer0_outputs(2347) <= not b;
    layer0_outputs(2348) <= not (a or b);
    layer0_outputs(2349) <= a or b;
    layer0_outputs(2350) <= not (a and b);
    layer0_outputs(2351) <= a or b;
    layer0_outputs(2352) <= 1'b0;
    layer0_outputs(2353) <= not b;
    layer0_outputs(2354) <= a and not b;
    layer0_outputs(2355) <= b;
    layer0_outputs(2356) <= a or b;
    layer0_outputs(2357) <= a and not b;
    layer0_outputs(2358) <= not (a and b);
    layer0_outputs(2359) <= not (a xor b);
    layer0_outputs(2360) <= not a or b;
    layer0_outputs(2361) <= not a;
    layer0_outputs(2362) <= not (a and b);
    layer0_outputs(2363) <= not (a or b);
    layer0_outputs(2364) <= a and b;
    layer0_outputs(2365) <= not a or b;
    layer0_outputs(2366) <= a xor b;
    layer0_outputs(2367) <= not a or b;
    layer0_outputs(2368) <= a;
    layer0_outputs(2369) <= not (a or b);
    layer0_outputs(2370) <= a xor b;
    layer0_outputs(2371) <= b;
    layer0_outputs(2372) <= not b or a;
    layer0_outputs(2373) <= not (a and b);
    layer0_outputs(2374) <= a or b;
    layer0_outputs(2375) <= a and not b;
    layer0_outputs(2376) <= not b or a;
    layer0_outputs(2377) <= not (a xor b);
    layer0_outputs(2378) <= a or b;
    layer0_outputs(2379) <= a or b;
    layer0_outputs(2380) <= b and not a;
    layer0_outputs(2381) <= b and not a;
    layer0_outputs(2382) <= not b;
    layer0_outputs(2383) <= not a;
    layer0_outputs(2384) <= not a;
    layer0_outputs(2385) <= not (a and b);
    layer0_outputs(2386) <= a xor b;
    layer0_outputs(2387) <= b and not a;
    layer0_outputs(2388) <= not b;
    layer0_outputs(2389) <= not b or a;
    layer0_outputs(2390) <= a xor b;
    layer0_outputs(2391) <= not a or b;
    layer0_outputs(2392) <= a xor b;
    layer0_outputs(2393) <= 1'b1;
    layer0_outputs(2394) <= b;
    layer0_outputs(2395) <= not (a or b);
    layer0_outputs(2396) <= not (a or b);
    layer0_outputs(2397) <= a or b;
    layer0_outputs(2398) <= a;
    layer0_outputs(2399) <= a or b;
    layer0_outputs(2400) <= a xor b;
    layer0_outputs(2401) <= not (a or b);
    layer0_outputs(2402) <= not a or b;
    layer0_outputs(2403) <= a and b;
    layer0_outputs(2404) <= not (a or b);
    layer0_outputs(2405) <= b and not a;
    layer0_outputs(2406) <= not a;
    layer0_outputs(2407) <= not a or b;
    layer0_outputs(2408) <= a;
    layer0_outputs(2409) <= not b or a;
    layer0_outputs(2410) <= 1'b1;
    layer0_outputs(2411) <= not (a or b);
    layer0_outputs(2412) <= not b;
    layer0_outputs(2413) <= a xor b;
    layer0_outputs(2414) <= a or b;
    layer0_outputs(2415) <= b and not a;
    layer0_outputs(2416) <= a xor b;
    layer0_outputs(2417) <= not (a or b);
    layer0_outputs(2418) <= a;
    layer0_outputs(2419) <= a or b;
    layer0_outputs(2420) <= 1'b0;
    layer0_outputs(2421) <= a;
    layer0_outputs(2422) <= a or b;
    layer0_outputs(2423) <= 1'b1;
    layer0_outputs(2424) <= not b;
    layer0_outputs(2425) <= not a;
    layer0_outputs(2426) <= not b or a;
    layer0_outputs(2427) <= not (a or b);
    layer0_outputs(2428) <= a and not b;
    layer0_outputs(2429) <= not (a or b);
    layer0_outputs(2430) <= not (a and b);
    layer0_outputs(2431) <= 1'b0;
    layer0_outputs(2432) <= a;
    layer0_outputs(2433) <= not (a or b);
    layer0_outputs(2434) <= not a or b;
    layer0_outputs(2435) <= b;
    layer0_outputs(2436) <= a xor b;
    layer0_outputs(2437) <= a;
    layer0_outputs(2438) <= a and not b;
    layer0_outputs(2439) <= not b;
    layer0_outputs(2440) <= a xor b;
    layer0_outputs(2441) <= not a or b;
    layer0_outputs(2442) <= not b or a;
    layer0_outputs(2443) <= b;
    layer0_outputs(2444) <= a and not b;
    layer0_outputs(2445) <= b;
    layer0_outputs(2446) <= b and not a;
    layer0_outputs(2447) <= not (a or b);
    layer0_outputs(2448) <= not (a xor b);
    layer0_outputs(2449) <= 1'b0;
    layer0_outputs(2450) <= not (a or b);
    layer0_outputs(2451) <= a;
    layer0_outputs(2452) <= 1'b1;
    layer0_outputs(2453) <= b;
    layer0_outputs(2454) <= not (a xor b);
    layer0_outputs(2455) <= not (a and b);
    layer0_outputs(2456) <= a or b;
    layer0_outputs(2457) <= b and not a;
    layer0_outputs(2458) <= not b or a;
    layer0_outputs(2459) <= not a;
    layer0_outputs(2460) <= a or b;
    layer0_outputs(2461) <= a and not b;
    layer0_outputs(2462) <= not b;
    layer0_outputs(2463) <= a;
    layer0_outputs(2464) <= b and not a;
    layer0_outputs(2465) <= 1'b1;
    layer0_outputs(2466) <= a or b;
    layer0_outputs(2467) <= b and not a;
    layer0_outputs(2468) <= a;
    layer0_outputs(2469) <= not a or b;
    layer0_outputs(2470) <= not (a or b);
    layer0_outputs(2471) <= not a or b;
    layer0_outputs(2472) <= not (a or b);
    layer0_outputs(2473) <= a or b;
    layer0_outputs(2474) <= b;
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= 1'b1;
    layer0_outputs(2477) <= b and not a;
    layer0_outputs(2478) <= not (a and b);
    layer0_outputs(2479) <= not (a or b);
    layer0_outputs(2480) <= a;
    layer0_outputs(2481) <= not a or b;
    layer0_outputs(2482) <= a or b;
    layer0_outputs(2483) <= not (a xor b);
    layer0_outputs(2484) <= a or b;
    layer0_outputs(2485) <= b and not a;
    layer0_outputs(2486) <= not (a xor b);
    layer0_outputs(2487) <= not a or b;
    layer0_outputs(2488) <= b and not a;
    layer0_outputs(2489) <= not (a or b);
    layer0_outputs(2490) <= not a;
    layer0_outputs(2491) <= not (a or b);
    layer0_outputs(2492) <= not b;
    layer0_outputs(2493) <= not b or a;
    layer0_outputs(2494) <= a or b;
    layer0_outputs(2495) <= not (a or b);
    layer0_outputs(2496) <= b;
    layer0_outputs(2497) <= 1'b1;
    layer0_outputs(2498) <= 1'b1;
    layer0_outputs(2499) <= not (a or b);
    layer0_outputs(2500) <= a or b;
    layer0_outputs(2501) <= not a;
    layer0_outputs(2502) <= not (a or b);
    layer0_outputs(2503) <= a;
    layer0_outputs(2504) <= a xor b;
    layer0_outputs(2505) <= not (a xor b);
    layer0_outputs(2506) <= 1'b1;
    layer0_outputs(2507) <= not a;
    layer0_outputs(2508) <= a or b;
    layer0_outputs(2509) <= a and not b;
    layer0_outputs(2510) <= not a;
    layer0_outputs(2511) <= not a;
    layer0_outputs(2512) <= not a or b;
    layer0_outputs(2513) <= 1'b0;
    layer0_outputs(2514) <= not (a or b);
    layer0_outputs(2515) <= b;
    layer0_outputs(2516) <= not (a or b);
    layer0_outputs(2517) <= b;
    layer0_outputs(2518) <= not b;
    layer0_outputs(2519) <= a and not b;
    layer0_outputs(2520) <= not a or b;
    layer0_outputs(2521) <= not a;
    layer0_outputs(2522) <= not a;
    layer0_outputs(2523) <= not b or a;
    layer0_outputs(2524) <= not a;
    layer0_outputs(2525) <= a xor b;
    layer0_outputs(2526) <= a;
    layer0_outputs(2527) <= a or b;
    layer0_outputs(2528) <= a or b;
    layer0_outputs(2529) <= not (a and b);
    layer0_outputs(2530) <= not a;
    layer0_outputs(2531) <= a xor b;
    layer0_outputs(2532) <= not b;
    layer0_outputs(2533) <= not b or a;
    layer0_outputs(2534) <= not (a xor b);
    layer0_outputs(2535) <= not b;
    layer0_outputs(2536) <= not b or a;
    layer0_outputs(2537) <= 1'b1;
    layer0_outputs(2538) <= b;
    layer0_outputs(2539) <= a;
    layer0_outputs(2540) <= not (a xor b);
    layer0_outputs(2541) <= a;
    layer0_outputs(2542) <= not a;
    layer0_outputs(2543) <= 1'b0;
    layer0_outputs(2544) <= not a;
    layer0_outputs(2545) <= a or b;
    layer0_outputs(2546) <= b;
    layer0_outputs(2547) <= not a or b;
    layer0_outputs(2548) <= not a;
    layer0_outputs(2549) <= not (a xor b);
    layer0_outputs(2550) <= not a;
    layer0_outputs(2551) <= not (a or b);
    layer0_outputs(2552) <= b and not a;
    layer0_outputs(2553) <= not (a or b);
    layer0_outputs(2554) <= a;
    layer0_outputs(2555) <= not b or a;
    layer0_outputs(2556) <= a xor b;
    layer0_outputs(2557) <= b;
    layer0_outputs(2558) <= b;
    layer0_outputs(2559) <= b;
    layer0_outputs(2560) <= b and not a;
    layer0_outputs(2561) <= not (a and b);
    layer0_outputs(2562) <= not a or b;
    layer0_outputs(2563) <= not (a xor b);
    layer0_outputs(2564) <= b;
    layer0_outputs(2565) <= not a or b;
    layer0_outputs(2566) <= not (a xor b);
    layer0_outputs(2567) <= a xor b;
    layer0_outputs(2568) <= a or b;
    layer0_outputs(2569) <= not b;
    layer0_outputs(2570) <= 1'b1;
    layer0_outputs(2571) <= not b;
    layer0_outputs(2572) <= a and not b;
    layer0_outputs(2573) <= not a;
    layer0_outputs(2574) <= a or b;
    layer0_outputs(2575) <= a or b;
    layer0_outputs(2576) <= not b or a;
    layer0_outputs(2577) <= not (a xor b);
    layer0_outputs(2578) <= b;
    layer0_outputs(2579) <= a and not b;
    layer0_outputs(2580) <= not (a or b);
    layer0_outputs(2581) <= a;
    layer0_outputs(2582) <= b and not a;
    layer0_outputs(2583) <= b;
    layer0_outputs(2584) <= a and not b;
    layer0_outputs(2585) <= not (a xor b);
    layer0_outputs(2586) <= a and not b;
    layer0_outputs(2587) <= not (a or b);
    layer0_outputs(2588) <= not (a or b);
    layer0_outputs(2589) <= not (a xor b);
    layer0_outputs(2590) <= not (a or b);
    layer0_outputs(2591) <= not a;
    layer0_outputs(2592) <= a or b;
    layer0_outputs(2593) <= not a or b;
    layer0_outputs(2594) <= not a;
    layer0_outputs(2595) <= not a or b;
    layer0_outputs(2596) <= a or b;
    layer0_outputs(2597) <= not b;
    layer0_outputs(2598) <= a or b;
    layer0_outputs(2599) <= 1'b1;
    layer0_outputs(2600) <= not b;
    layer0_outputs(2601) <= a;
    layer0_outputs(2602) <= not b or a;
    layer0_outputs(2603) <= not (a or b);
    layer0_outputs(2604) <= not b;
    layer0_outputs(2605) <= a and not b;
    layer0_outputs(2606) <= b and not a;
    layer0_outputs(2607) <= a and not b;
    layer0_outputs(2608) <= not b or a;
    layer0_outputs(2609) <= a xor b;
    layer0_outputs(2610) <= not a or b;
    layer0_outputs(2611) <= not a;
    layer0_outputs(2612) <= not b;
    layer0_outputs(2613) <= a xor b;
    layer0_outputs(2614) <= a or b;
    layer0_outputs(2615) <= a or b;
    layer0_outputs(2616) <= a or b;
    layer0_outputs(2617) <= not (a or b);
    layer0_outputs(2618) <= not (a xor b);
    layer0_outputs(2619) <= a;
    layer0_outputs(2620) <= a or b;
    layer0_outputs(2621) <= not a;
    layer0_outputs(2622) <= not b;
    layer0_outputs(2623) <= a and not b;
    layer0_outputs(2624) <= not a or b;
    layer0_outputs(2625) <= not a;
    layer0_outputs(2626) <= a xor b;
    layer0_outputs(2627) <= not b;
    layer0_outputs(2628) <= a xor b;
    layer0_outputs(2629) <= not b;
    layer0_outputs(2630) <= not (a and b);
    layer0_outputs(2631) <= not (a xor b);
    layer0_outputs(2632) <= not (a and b);
    layer0_outputs(2633) <= a;
    layer0_outputs(2634) <= not a or b;
    layer0_outputs(2635) <= a or b;
    layer0_outputs(2636) <= not (a or b);
    layer0_outputs(2637) <= not a;
    layer0_outputs(2638) <= a;
    layer0_outputs(2639) <= not a or b;
    layer0_outputs(2640) <= not a;
    layer0_outputs(2641) <= a;
    layer0_outputs(2642) <= a and not b;
    layer0_outputs(2643) <= not (a or b);
    layer0_outputs(2644) <= 1'b1;
    layer0_outputs(2645) <= 1'b1;
    layer0_outputs(2646) <= not b;
    layer0_outputs(2647) <= b and not a;
    layer0_outputs(2648) <= not a or b;
    layer0_outputs(2649) <= 1'b1;
    layer0_outputs(2650) <= b;
    layer0_outputs(2651) <= a and not b;
    layer0_outputs(2652) <= b;
    layer0_outputs(2653) <= 1'b0;
    layer0_outputs(2654) <= a;
    layer0_outputs(2655) <= 1'b1;
    layer0_outputs(2656) <= not b;
    layer0_outputs(2657) <= not (a xor b);
    layer0_outputs(2658) <= b and not a;
    layer0_outputs(2659) <= not b or a;
    layer0_outputs(2660) <= a xor b;
    layer0_outputs(2661) <= 1'b0;
    layer0_outputs(2662) <= 1'b0;
    layer0_outputs(2663) <= a xor b;
    layer0_outputs(2664) <= not (a or b);
    layer0_outputs(2665) <= a xor b;
    layer0_outputs(2666) <= 1'b0;
    layer0_outputs(2667) <= 1'b0;
    layer0_outputs(2668) <= not b or a;
    layer0_outputs(2669) <= a;
    layer0_outputs(2670) <= b;
    layer0_outputs(2671) <= not (a or b);
    layer0_outputs(2672) <= not b or a;
    layer0_outputs(2673) <= a;
    layer0_outputs(2674) <= b and not a;
    layer0_outputs(2675) <= a and not b;
    layer0_outputs(2676) <= not b;
    layer0_outputs(2677) <= a;
    layer0_outputs(2678) <= a and not b;
    layer0_outputs(2679) <= b;
    layer0_outputs(2680) <= b and not a;
    layer0_outputs(2681) <= not a or b;
    layer0_outputs(2682) <= not (a and b);
    layer0_outputs(2683) <= a and not b;
    layer0_outputs(2684) <= not b;
    layer0_outputs(2685) <= not b;
    layer0_outputs(2686) <= not a or b;
    layer0_outputs(2687) <= a or b;
    layer0_outputs(2688) <= a;
    layer0_outputs(2689) <= a or b;
    layer0_outputs(2690) <= b;
    layer0_outputs(2691) <= not a;
    layer0_outputs(2692) <= a and not b;
    layer0_outputs(2693) <= a;
    layer0_outputs(2694) <= not a;
    layer0_outputs(2695) <= not a;
    layer0_outputs(2696) <= not a or b;
    layer0_outputs(2697) <= not a;
    layer0_outputs(2698) <= not b;
    layer0_outputs(2699) <= not (a or b);
    layer0_outputs(2700) <= a and not b;
    layer0_outputs(2701) <= not (a xor b);
    layer0_outputs(2702) <= not b or a;
    layer0_outputs(2703) <= b and not a;
    layer0_outputs(2704) <= not a;
    layer0_outputs(2705) <= a xor b;
    layer0_outputs(2706) <= not a;
    layer0_outputs(2707) <= not (a and b);
    layer0_outputs(2708) <= a xor b;
    layer0_outputs(2709) <= not a or b;
    layer0_outputs(2710) <= not a;
    layer0_outputs(2711) <= 1'b1;
    layer0_outputs(2712) <= not (a xor b);
    layer0_outputs(2713) <= a and not b;
    layer0_outputs(2714) <= b and not a;
    layer0_outputs(2715) <= not a or b;
    layer0_outputs(2716) <= a and not b;
    layer0_outputs(2717) <= not (a xor b);
    layer0_outputs(2718) <= not a;
    layer0_outputs(2719) <= not (a and b);
    layer0_outputs(2720) <= a and b;
    layer0_outputs(2721) <= not a or b;
    layer0_outputs(2722) <= 1'b0;
    layer0_outputs(2723) <= not (a or b);
    layer0_outputs(2724) <= not a;
    layer0_outputs(2725) <= b and not a;
    layer0_outputs(2726) <= a or b;
    layer0_outputs(2727) <= not (a xor b);
    layer0_outputs(2728) <= a xor b;
    layer0_outputs(2729) <= not (a or b);
    layer0_outputs(2730) <= a and not b;
    layer0_outputs(2731) <= not (a and b);
    layer0_outputs(2732) <= a or b;
    layer0_outputs(2733) <= not (a or b);
    layer0_outputs(2734) <= not (a or b);
    layer0_outputs(2735) <= b and not a;
    layer0_outputs(2736) <= b;
    layer0_outputs(2737) <= 1'b1;
    layer0_outputs(2738) <= not b;
    layer0_outputs(2739) <= not (a or b);
    layer0_outputs(2740) <= not b or a;
    layer0_outputs(2741) <= 1'b1;
    layer0_outputs(2742) <= a and b;
    layer0_outputs(2743) <= b and not a;
    layer0_outputs(2744) <= not b;
    layer0_outputs(2745) <= not a or b;
    layer0_outputs(2746) <= a xor b;
    layer0_outputs(2747) <= not a;
    layer0_outputs(2748) <= 1'b0;
    layer0_outputs(2749) <= b and not a;
    layer0_outputs(2750) <= not a;
    layer0_outputs(2751) <= not b;
    layer0_outputs(2752) <= not a or b;
    layer0_outputs(2753) <= not (a or b);
    layer0_outputs(2754) <= a or b;
    layer0_outputs(2755) <= b and not a;
    layer0_outputs(2756) <= not a;
    layer0_outputs(2757) <= b and not a;
    layer0_outputs(2758) <= a;
    layer0_outputs(2759) <= not a;
    layer0_outputs(2760) <= b and not a;
    layer0_outputs(2761) <= b and not a;
    layer0_outputs(2762) <= not b or a;
    layer0_outputs(2763) <= b;
    layer0_outputs(2764) <= a xor b;
    layer0_outputs(2765) <= b;
    layer0_outputs(2766) <= a and not b;
    layer0_outputs(2767) <= not a;
    layer0_outputs(2768) <= a or b;
    layer0_outputs(2769) <= b;
    layer0_outputs(2770) <= b;
    layer0_outputs(2771) <= not a or b;
    layer0_outputs(2772) <= a or b;
    layer0_outputs(2773) <= b and not a;
    layer0_outputs(2774) <= not (a or b);
    layer0_outputs(2775) <= not a or b;
    layer0_outputs(2776) <= not b;
    layer0_outputs(2777) <= a and b;
    layer0_outputs(2778) <= not a;
    layer0_outputs(2779) <= not (a and b);
    layer0_outputs(2780) <= 1'b0;
    layer0_outputs(2781) <= a and b;
    layer0_outputs(2782) <= 1'b1;
    layer0_outputs(2783) <= not a;
    layer0_outputs(2784) <= 1'b0;
    layer0_outputs(2785) <= not b or a;
    layer0_outputs(2786) <= b;
    layer0_outputs(2787) <= 1'b1;
    layer0_outputs(2788) <= a;
    layer0_outputs(2789) <= not (a and b);
    layer0_outputs(2790) <= a and not b;
    layer0_outputs(2791) <= a and b;
    layer0_outputs(2792) <= a or b;
    layer0_outputs(2793) <= not a;
    layer0_outputs(2794) <= 1'b1;
    layer0_outputs(2795) <= not (a or b);
    layer0_outputs(2796) <= b;
    layer0_outputs(2797) <= not b;
    layer0_outputs(2798) <= not a;
    layer0_outputs(2799) <= a or b;
    layer0_outputs(2800) <= not b;
    layer0_outputs(2801) <= not a or b;
    layer0_outputs(2802) <= not a or b;
    layer0_outputs(2803) <= a or b;
    layer0_outputs(2804) <= not b;
    layer0_outputs(2805) <= b;
    layer0_outputs(2806) <= a;
    layer0_outputs(2807) <= a;
    layer0_outputs(2808) <= not a;
    layer0_outputs(2809) <= not a;
    layer0_outputs(2810) <= not a or b;
    layer0_outputs(2811) <= a and b;
    layer0_outputs(2812) <= not (a or b);
    layer0_outputs(2813) <= a and not b;
    layer0_outputs(2814) <= a and not b;
    layer0_outputs(2815) <= not (a or b);
    layer0_outputs(2816) <= b;
    layer0_outputs(2817) <= not b;
    layer0_outputs(2818) <= not (a xor b);
    layer0_outputs(2819) <= not a;
    layer0_outputs(2820) <= 1'b0;
    layer0_outputs(2821) <= a and not b;
    layer0_outputs(2822) <= a and not b;
    layer0_outputs(2823) <= not (a or b);
    layer0_outputs(2824) <= a;
    layer0_outputs(2825) <= not (a or b);
    layer0_outputs(2826) <= not (a xor b);
    layer0_outputs(2827) <= not a or b;
    layer0_outputs(2828) <= not b;
    layer0_outputs(2829) <= a and not b;
    layer0_outputs(2830) <= 1'b0;
    layer0_outputs(2831) <= not b or a;
    layer0_outputs(2832) <= b and not a;
    layer0_outputs(2833) <= a or b;
    layer0_outputs(2834) <= 1'b0;
    layer0_outputs(2835) <= not a;
    layer0_outputs(2836) <= not (a or b);
    layer0_outputs(2837) <= b and not a;
    layer0_outputs(2838) <= a xor b;
    layer0_outputs(2839) <= 1'b0;
    layer0_outputs(2840) <= b and not a;
    layer0_outputs(2841) <= a;
    layer0_outputs(2842) <= a or b;
    layer0_outputs(2843) <= not b;
    layer0_outputs(2844) <= a or b;
    layer0_outputs(2845) <= not b or a;
    layer0_outputs(2846) <= not (a xor b);
    layer0_outputs(2847) <= not a or b;
    layer0_outputs(2848) <= not (a or b);
    layer0_outputs(2849) <= a and b;
    layer0_outputs(2850) <= not (a xor b);
    layer0_outputs(2851) <= 1'b1;
    layer0_outputs(2852) <= not (a or b);
    layer0_outputs(2853) <= not (a xor b);
    layer0_outputs(2854) <= not a or b;
    layer0_outputs(2855) <= not b;
    layer0_outputs(2856) <= b and not a;
    layer0_outputs(2857) <= not (a or b);
    layer0_outputs(2858) <= not (a or b);
    layer0_outputs(2859) <= a and b;
    layer0_outputs(2860) <= not a;
    layer0_outputs(2861) <= 1'b1;
    layer0_outputs(2862) <= not b;
    layer0_outputs(2863) <= not a;
    layer0_outputs(2864) <= a;
    layer0_outputs(2865) <= a or b;
    layer0_outputs(2866) <= not b or a;
    layer0_outputs(2867) <= a or b;
    layer0_outputs(2868) <= not (a or b);
    layer0_outputs(2869) <= b and not a;
    layer0_outputs(2870) <= not b;
    layer0_outputs(2871) <= a and b;
    layer0_outputs(2872) <= not b or a;
    layer0_outputs(2873) <= a xor b;
    layer0_outputs(2874) <= not b or a;
    layer0_outputs(2875) <= a;
    layer0_outputs(2876) <= b;
    layer0_outputs(2877) <= a or b;
    layer0_outputs(2878) <= not (a xor b);
    layer0_outputs(2879) <= b;
    layer0_outputs(2880) <= not (a and b);
    layer0_outputs(2881) <= a;
    layer0_outputs(2882) <= not b or a;
    layer0_outputs(2883) <= not a or b;
    layer0_outputs(2884) <= not a;
    layer0_outputs(2885) <= b and not a;
    layer0_outputs(2886) <= a or b;
    layer0_outputs(2887) <= a xor b;
    layer0_outputs(2888) <= a and b;
    layer0_outputs(2889) <= not (a or b);
    layer0_outputs(2890) <= not (a or b);
    layer0_outputs(2891) <= b and not a;
    layer0_outputs(2892) <= a or b;
    layer0_outputs(2893) <= b and not a;
    layer0_outputs(2894) <= a or b;
    layer0_outputs(2895) <= not a or b;
    layer0_outputs(2896) <= 1'b1;
    layer0_outputs(2897) <= a and b;
    layer0_outputs(2898) <= not (a or b);
    layer0_outputs(2899) <= not a or b;
    layer0_outputs(2900) <= not b or a;
    layer0_outputs(2901) <= a xor b;
    layer0_outputs(2902) <= a or b;
    layer0_outputs(2903) <= a xor b;
    layer0_outputs(2904) <= 1'b0;
    layer0_outputs(2905) <= a or b;
    layer0_outputs(2906) <= 1'b0;
    layer0_outputs(2907) <= not a or b;
    layer0_outputs(2908) <= not a;
    layer0_outputs(2909) <= b;
    layer0_outputs(2910) <= not a;
    layer0_outputs(2911) <= a and b;
    layer0_outputs(2912) <= b and not a;
    layer0_outputs(2913) <= a xor b;
    layer0_outputs(2914) <= b;
    layer0_outputs(2915) <= not (a or b);
    layer0_outputs(2916) <= a and not b;
    layer0_outputs(2917) <= a or b;
    layer0_outputs(2918) <= not (a or b);
    layer0_outputs(2919) <= a or b;
    layer0_outputs(2920) <= 1'b1;
    layer0_outputs(2921) <= not (a or b);
    layer0_outputs(2922) <= not (a or b);
    layer0_outputs(2923) <= 1'b0;
    layer0_outputs(2924) <= not (a or b);
    layer0_outputs(2925) <= b;
    layer0_outputs(2926) <= b;
    layer0_outputs(2927) <= not (a or b);
    layer0_outputs(2928) <= b;
    layer0_outputs(2929) <= not a;
    layer0_outputs(2930) <= not (a or b);
    layer0_outputs(2931) <= not (a or b);
    layer0_outputs(2932) <= not b;
    layer0_outputs(2933) <= not (a and b);
    layer0_outputs(2934) <= not a or b;
    layer0_outputs(2935) <= b;
    layer0_outputs(2936) <= a and not b;
    layer0_outputs(2937) <= a;
    layer0_outputs(2938) <= not a;
    layer0_outputs(2939) <= a xor b;
    layer0_outputs(2940) <= b and not a;
    layer0_outputs(2941) <= not a;
    layer0_outputs(2942) <= b and not a;
    layer0_outputs(2943) <= not a;
    layer0_outputs(2944) <= not a or b;
    layer0_outputs(2945) <= not b;
    layer0_outputs(2946) <= a and not b;
    layer0_outputs(2947) <= not a or b;
    layer0_outputs(2948) <= b;
    layer0_outputs(2949) <= not (a xor b);
    layer0_outputs(2950) <= a or b;
    layer0_outputs(2951) <= a and not b;
    layer0_outputs(2952) <= not (a or b);
    layer0_outputs(2953) <= not (a xor b);
    layer0_outputs(2954) <= not (a or b);
    layer0_outputs(2955) <= 1'b0;
    layer0_outputs(2956) <= b and not a;
    layer0_outputs(2957) <= a;
    layer0_outputs(2958) <= not b;
    layer0_outputs(2959) <= b and not a;
    layer0_outputs(2960) <= not b or a;
    layer0_outputs(2961) <= a or b;
    layer0_outputs(2962) <= not (a or b);
    layer0_outputs(2963) <= a and not b;
    layer0_outputs(2964) <= not (a or b);
    layer0_outputs(2965) <= 1'b0;
    layer0_outputs(2966) <= 1'b0;
    layer0_outputs(2967) <= not b or a;
    layer0_outputs(2968) <= not a or b;
    layer0_outputs(2969) <= a or b;
    layer0_outputs(2970) <= not (a xor b);
    layer0_outputs(2971) <= not b;
    layer0_outputs(2972) <= not b;
    layer0_outputs(2973) <= not (a xor b);
    layer0_outputs(2974) <= a and not b;
    layer0_outputs(2975) <= a or b;
    layer0_outputs(2976) <= a or b;
    layer0_outputs(2977) <= not (a or b);
    layer0_outputs(2978) <= a or b;
    layer0_outputs(2979) <= a;
    layer0_outputs(2980) <= not (a or b);
    layer0_outputs(2981) <= a;
    layer0_outputs(2982) <= a xor b;
    layer0_outputs(2983) <= b and not a;
    layer0_outputs(2984) <= a or b;
    layer0_outputs(2985) <= a xor b;
    layer0_outputs(2986) <= not a;
    layer0_outputs(2987) <= a;
    layer0_outputs(2988) <= not (a xor b);
    layer0_outputs(2989) <= not b;
    layer0_outputs(2990) <= not a;
    layer0_outputs(2991) <= not (a or b);
    layer0_outputs(2992) <= not (a or b);
    layer0_outputs(2993) <= 1'b0;
    layer0_outputs(2994) <= b;
    layer0_outputs(2995) <= a;
    layer0_outputs(2996) <= a or b;
    layer0_outputs(2997) <= a and not b;
    layer0_outputs(2998) <= a;
    layer0_outputs(2999) <= a and not b;
    layer0_outputs(3000) <= not b or a;
    layer0_outputs(3001) <= not (a xor b);
    layer0_outputs(3002) <= a or b;
    layer0_outputs(3003) <= b;
    layer0_outputs(3004) <= not b;
    layer0_outputs(3005) <= not (a or b);
    layer0_outputs(3006) <= a xor b;
    layer0_outputs(3007) <= a;
    layer0_outputs(3008) <= a xor b;
    layer0_outputs(3009) <= a and not b;
    layer0_outputs(3010) <= not b or a;
    layer0_outputs(3011) <= a or b;
    layer0_outputs(3012) <= b and not a;
    layer0_outputs(3013) <= not (a xor b);
    layer0_outputs(3014) <= not a;
    layer0_outputs(3015) <= not (a or b);
    layer0_outputs(3016) <= not (a xor b);
    layer0_outputs(3017) <= a or b;
    layer0_outputs(3018) <= 1'b1;
    layer0_outputs(3019) <= b and not a;
    layer0_outputs(3020) <= not (a or b);
    layer0_outputs(3021) <= a;
    layer0_outputs(3022) <= not b or a;
    layer0_outputs(3023) <= b and not a;
    layer0_outputs(3024) <= a and not b;
    layer0_outputs(3025) <= a xor b;
    layer0_outputs(3026) <= a or b;
    layer0_outputs(3027) <= a or b;
    layer0_outputs(3028) <= not (a or b);
    layer0_outputs(3029) <= not a or b;
    layer0_outputs(3030) <= a and b;
    layer0_outputs(3031) <= not a;
    layer0_outputs(3032) <= not b or a;
    layer0_outputs(3033) <= not b or a;
    layer0_outputs(3034) <= 1'b1;
    layer0_outputs(3035) <= 1'b1;
    layer0_outputs(3036) <= not b;
    layer0_outputs(3037) <= not (a xor b);
    layer0_outputs(3038) <= 1'b1;
    layer0_outputs(3039) <= not a or b;
    layer0_outputs(3040) <= not (a and b);
    layer0_outputs(3041) <= a;
    layer0_outputs(3042) <= a;
    layer0_outputs(3043) <= a or b;
    layer0_outputs(3044) <= not b;
    layer0_outputs(3045) <= a and b;
    layer0_outputs(3046) <= not (a or b);
    layer0_outputs(3047) <= b;
    layer0_outputs(3048) <= not a;
    layer0_outputs(3049) <= not (a xor b);
    layer0_outputs(3050) <= a and b;
    layer0_outputs(3051) <= not a or b;
    layer0_outputs(3052) <= b;
    layer0_outputs(3053) <= a xor b;
    layer0_outputs(3054) <= not (a and b);
    layer0_outputs(3055) <= a xor b;
    layer0_outputs(3056) <= not (a or b);
    layer0_outputs(3057) <= not (a or b);
    layer0_outputs(3058) <= not a or b;
    layer0_outputs(3059) <= not a;
    layer0_outputs(3060) <= not b or a;
    layer0_outputs(3061) <= not a or b;
    layer0_outputs(3062) <= a or b;
    layer0_outputs(3063) <= not b or a;
    layer0_outputs(3064) <= not (a xor b);
    layer0_outputs(3065) <= 1'b0;
    layer0_outputs(3066) <= b;
    layer0_outputs(3067) <= a;
    layer0_outputs(3068) <= a or b;
    layer0_outputs(3069) <= not b or a;
    layer0_outputs(3070) <= b;
    layer0_outputs(3071) <= b;
    layer0_outputs(3072) <= a;
    layer0_outputs(3073) <= b;
    layer0_outputs(3074) <= a xor b;
    layer0_outputs(3075) <= a or b;
    layer0_outputs(3076) <= not b or a;
    layer0_outputs(3077) <= not b;
    layer0_outputs(3078) <= a and not b;
    layer0_outputs(3079) <= not b or a;
    layer0_outputs(3080) <= not a;
    layer0_outputs(3081) <= b;
    layer0_outputs(3082) <= a xor b;
    layer0_outputs(3083) <= not (a or b);
    layer0_outputs(3084) <= not b;
    layer0_outputs(3085) <= not (a or b);
    layer0_outputs(3086) <= not a;
    layer0_outputs(3087) <= not b or a;
    layer0_outputs(3088) <= not b;
    layer0_outputs(3089) <= a or b;
    layer0_outputs(3090) <= not b;
    layer0_outputs(3091) <= not a;
    layer0_outputs(3092) <= not (a or b);
    layer0_outputs(3093) <= not (a xor b);
    layer0_outputs(3094) <= not b or a;
    layer0_outputs(3095) <= 1'b1;
    layer0_outputs(3096) <= not a or b;
    layer0_outputs(3097) <= not b or a;
    layer0_outputs(3098) <= not b or a;
    layer0_outputs(3099) <= not a or b;
    layer0_outputs(3100) <= not b or a;
    layer0_outputs(3101) <= a or b;
    layer0_outputs(3102) <= not (a or b);
    layer0_outputs(3103) <= 1'b0;
    layer0_outputs(3104) <= not a;
    layer0_outputs(3105) <= not (a xor b);
    layer0_outputs(3106) <= not a or b;
    layer0_outputs(3107) <= a or b;
    layer0_outputs(3108) <= not (a or b);
    layer0_outputs(3109) <= not (a and b);
    layer0_outputs(3110) <= a xor b;
    layer0_outputs(3111) <= not (a or b);
    layer0_outputs(3112) <= a or b;
    layer0_outputs(3113) <= not b;
    layer0_outputs(3114) <= b;
    layer0_outputs(3115) <= not a;
    layer0_outputs(3116) <= not a;
    layer0_outputs(3117) <= b;
    layer0_outputs(3118) <= a or b;
    layer0_outputs(3119) <= not a;
    layer0_outputs(3120) <= a and b;
    layer0_outputs(3121) <= a or b;
    layer0_outputs(3122) <= not (a or b);
    layer0_outputs(3123) <= a and not b;
    layer0_outputs(3124) <= b;
    layer0_outputs(3125) <= not a or b;
    layer0_outputs(3126) <= b;
    layer0_outputs(3127) <= not a;
    layer0_outputs(3128) <= b;
    layer0_outputs(3129) <= a;
    layer0_outputs(3130) <= a;
    layer0_outputs(3131) <= not b or a;
    layer0_outputs(3132) <= a;
    layer0_outputs(3133) <= a;
    layer0_outputs(3134) <= a and b;
    layer0_outputs(3135) <= not (a or b);
    layer0_outputs(3136) <= not b or a;
    layer0_outputs(3137) <= not (a or b);
    layer0_outputs(3138) <= 1'b1;
    layer0_outputs(3139) <= a or b;
    layer0_outputs(3140) <= not (a or b);
    layer0_outputs(3141) <= a xor b;
    layer0_outputs(3142) <= not (a or b);
    layer0_outputs(3143) <= b;
    layer0_outputs(3144) <= not a;
    layer0_outputs(3145) <= not (a or b);
    layer0_outputs(3146) <= not b;
    layer0_outputs(3147) <= 1'b0;
    layer0_outputs(3148) <= b and not a;
    layer0_outputs(3149) <= a;
    layer0_outputs(3150) <= not (a or b);
    layer0_outputs(3151) <= a xor b;
    layer0_outputs(3152) <= 1'b0;
    layer0_outputs(3153) <= not (a xor b);
    layer0_outputs(3154) <= not (a xor b);
    layer0_outputs(3155) <= 1'b1;
    layer0_outputs(3156) <= a;
    layer0_outputs(3157) <= not a;
    layer0_outputs(3158) <= not b or a;
    layer0_outputs(3159) <= b;
    layer0_outputs(3160) <= not b or a;
    layer0_outputs(3161) <= a and not b;
    layer0_outputs(3162) <= a and not b;
    layer0_outputs(3163) <= a or b;
    layer0_outputs(3164) <= b;
    layer0_outputs(3165) <= b and not a;
    layer0_outputs(3166) <= a and not b;
    layer0_outputs(3167) <= not a or b;
    layer0_outputs(3168) <= a;
    layer0_outputs(3169) <= a or b;
    layer0_outputs(3170) <= not (a or b);
    layer0_outputs(3171) <= not a or b;
    layer0_outputs(3172) <= 1'b0;
    layer0_outputs(3173) <= not (a and b);
    layer0_outputs(3174) <= a or b;
    layer0_outputs(3175) <= a or b;
    layer0_outputs(3176) <= a;
    layer0_outputs(3177) <= a;
    layer0_outputs(3178) <= not a or b;
    layer0_outputs(3179) <= not b or a;
    layer0_outputs(3180) <= not a or b;
    layer0_outputs(3181) <= a or b;
    layer0_outputs(3182) <= not (a or b);
    layer0_outputs(3183) <= not (a or b);
    layer0_outputs(3184) <= not b or a;
    layer0_outputs(3185) <= a;
    layer0_outputs(3186) <= not b or a;
    layer0_outputs(3187) <= not a or b;
    layer0_outputs(3188) <= a or b;
    layer0_outputs(3189) <= a;
    layer0_outputs(3190) <= b;
    layer0_outputs(3191) <= not b;
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= not a;
    layer0_outputs(3194) <= not a or b;
    layer0_outputs(3195) <= not b;
    layer0_outputs(3196) <= not (a or b);
    layer0_outputs(3197) <= not (a or b);
    layer0_outputs(3198) <= a and not b;
    layer0_outputs(3199) <= a xor b;
    layer0_outputs(3200) <= a or b;
    layer0_outputs(3201) <= 1'b0;
    layer0_outputs(3202) <= a or b;
    layer0_outputs(3203) <= a xor b;
    layer0_outputs(3204) <= not a;
    layer0_outputs(3205) <= not (a or b);
    layer0_outputs(3206) <= a xor b;
    layer0_outputs(3207) <= not a or b;
    layer0_outputs(3208) <= not (a or b);
    layer0_outputs(3209) <= a;
    layer0_outputs(3210) <= a or b;
    layer0_outputs(3211) <= not b or a;
    layer0_outputs(3212) <= b and not a;
    layer0_outputs(3213) <= not (a or b);
    layer0_outputs(3214) <= 1'b1;
    layer0_outputs(3215) <= a xor b;
    layer0_outputs(3216) <= not (a or b);
    layer0_outputs(3217) <= not (a or b);
    layer0_outputs(3218) <= not (a xor b);
    layer0_outputs(3219) <= not b or a;
    layer0_outputs(3220) <= not (a xor b);
    layer0_outputs(3221) <= not a;
    layer0_outputs(3222) <= a or b;
    layer0_outputs(3223) <= not a;
    layer0_outputs(3224) <= a or b;
    layer0_outputs(3225) <= a or b;
    layer0_outputs(3226) <= not (a or b);
    layer0_outputs(3227) <= b;
    layer0_outputs(3228) <= b and not a;
    layer0_outputs(3229) <= not a or b;
    layer0_outputs(3230) <= not (a or b);
    layer0_outputs(3231) <= not b;
    layer0_outputs(3232) <= b;
    layer0_outputs(3233) <= not (a or b);
    layer0_outputs(3234) <= a or b;
    layer0_outputs(3235) <= not a or b;
    layer0_outputs(3236) <= not b;
    layer0_outputs(3237) <= not (a xor b);
    layer0_outputs(3238) <= not (a or b);
    layer0_outputs(3239) <= not a or b;
    layer0_outputs(3240) <= not b;
    layer0_outputs(3241) <= b;
    layer0_outputs(3242) <= a and b;
    layer0_outputs(3243) <= a;
    layer0_outputs(3244) <= 1'b1;
    layer0_outputs(3245) <= not a;
    layer0_outputs(3246) <= not b or a;
    layer0_outputs(3247) <= not a;
    layer0_outputs(3248) <= a or b;
    layer0_outputs(3249) <= a and b;
    layer0_outputs(3250) <= not (a xor b);
    layer0_outputs(3251) <= not (a or b);
    layer0_outputs(3252) <= not a;
    layer0_outputs(3253) <= a or b;
    layer0_outputs(3254) <= not a;
    layer0_outputs(3255) <= a or b;
    layer0_outputs(3256) <= a or b;
    layer0_outputs(3257) <= b;
    layer0_outputs(3258) <= a and not b;
    layer0_outputs(3259) <= a and b;
    layer0_outputs(3260) <= not b;
    layer0_outputs(3261) <= a xor b;
    layer0_outputs(3262) <= a or b;
    layer0_outputs(3263) <= a;
    layer0_outputs(3264) <= a xor b;
    layer0_outputs(3265) <= not a or b;
    layer0_outputs(3266) <= not a or b;
    layer0_outputs(3267) <= not b;
    layer0_outputs(3268) <= a or b;
    layer0_outputs(3269) <= b and not a;
    layer0_outputs(3270) <= not (a or b);
    layer0_outputs(3271) <= a and not b;
    layer0_outputs(3272) <= not (a or b);
    layer0_outputs(3273) <= a and not b;
    layer0_outputs(3274) <= not b or a;
    layer0_outputs(3275) <= not b;
    layer0_outputs(3276) <= not a or b;
    layer0_outputs(3277) <= not (a and b);
    layer0_outputs(3278) <= a and not b;
    layer0_outputs(3279) <= 1'b0;
    layer0_outputs(3280) <= not a;
    layer0_outputs(3281) <= a xor b;
    layer0_outputs(3282) <= a xor b;
    layer0_outputs(3283) <= not a or b;
    layer0_outputs(3284) <= not (a or b);
    layer0_outputs(3285) <= a and not b;
    layer0_outputs(3286) <= a;
    layer0_outputs(3287) <= a or b;
    layer0_outputs(3288) <= a or b;
    layer0_outputs(3289) <= a and not b;
    layer0_outputs(3290) <= not (a or b);
    layer0_outputs(3291) <= not a;
    layer0_outputs(3292) <= b and not a;
    layer0_outputs(3293) <= not b;
    layer0_outputs(3294) <= b and not a;
    layer0_outputs(3295) <= not b or a;
    layer0_outputs(3296) <= not (a xor b);
    layer0_outputs(3297) <= b and not a;
    layer0_outputs(3298) <= b and not a;
    layer0_outputs(3299) <= a and not b;
    layer0_outputs(3300) <= b;
    layer0_outputs(3301) <= a or b;
    layer0_outputs(3302) <= b and not a;
    layer0_outputs(3303) <= not b or a;
    layer0_outputs(3304) <= not (a or b);
    layer0_outputs(3305) <= b;
    layer0_outputs(3306) <= not (a xor b);
    layer0_outputs(3307) <= b and not a;
    layer0_outputs(3308) <= a or b;
    layer0_outputs(3309) <= a;
    layer0_outputs(3310) <= a or b;
    layer0_outputs(3311) <= not a;
    layer0_outputs(3312) <= a or b;
    layer0_outputs(3313) <= a or b;
    layer0_outputs(3314) <= not b or a;
    layer0_outputs(3315) <= not (a xor b);
    layer0_outputs(3316) <= a or b;
    layer0_outputs(3317) <= b;
    layer0_outputs(3318) <= a and not b;
    layer0_outputs(3319) <= a or b;
    layer0_outputs(3320) <= not a;
    layer0_outputs(3321) <= not b or a;
    layer0_outputs(3322) <= not b;
    layer0_outputs(3323) <= not a;
    layer0_outputs(3324) <= a or b;
    layer0_outputs(3325) <= b;
    layer0_outputs(3326) <= not a;
    layer0_outputs(3327) <= b;
    layer0_outputs(3328) <= a;
    layer0_outputs(3329) <= a or b;
    layer0_outputs(3330) <= not b or a;
    layer0_outputs(3331) <= a or b;
    layer0_outputs(3332) <= a;
    layer0_outputs(3333) <= not (a or b);
    layer0_outputs(3334) <= b;
    layer0_outputs(3335) <= a or b;
    layer0_outputs(3336) <= b;
    layer0_outputs(3337) <= a or b;
    layer0_outputs(3338) <= not (a or b);
    layer0_outputs(3339) <= a or b;
    layer0_outputs(3340) <= a xor b;
    layer0_outputs(3341) <= not a;
    layer0_outputs(3342) <= a or b;
    layer0_outputs(3343) <= not b;
    layer0_outputs(3344) <= not a;
    layer0_outputs(3345) <= not (a xor b);
    layer0_outputs(3346) <= not b or a;
    layer0_outputs(3347) <= a or b;
    layer0_outputs(3348) <= not (a and b);
    layer0_outputs(3349) <= not (a xor b);
    layer0_outputs(3350) <= a or b;
    layer0_outputs(3351) <= not (a xor b);
    layer0_outputs(3352) <= not (a xor b);
    layer0_outputs(3353) <= not (a or b);
    layer0_outputs(3354) <= b;
    layer0_outputs(3355) <= not (a or b);
    layer0_outputs(3356) <= not (a or b);
    layer0_outputs(3357) <= 1'b0;
    layer0_outputs(3358) <= not (a and b);
    layer0_outputs(3359) <= a;
    layer0_outputs(3360) <= b and not a;
    layer0_outputs(3361) <= not (a xor b);
    layer0_outputs(3362) <= b;
    layer0_outputs(3363) <= a;
    layer0_outputs(3364) <= a;
    layer0_outputs(3365) <= not (a or b);
    layer0_outputs(3366) <= a and b;
    layer0_outputs(3367) <= not b;
    layer0_outputs(3368) <= 1'b0;
    layer0_outputs(3369) <= a and b;
    layer0_outputs(3370) <= not (a xor b);
    layer0_outputs(3371) <= not a or b;
    layer0_outputs(3372) <= not (a xor b);
    layer0_outputs(3373) <= b;
    layer0_outputs(3374) <= not (a xor b);
    layer0_outputs(3375) <= not b;
    layer0_outputs(3376) <= not b;
    layer0_outputs(3377) <= not b or a;
    layer0_outputs(3378) <= not b;
    layer0_outputs(3379) <= a and not b;
    layer0_outputs(3380) <= b and not a;
    layer0_outputs(3381) <= not a;
    layer0_outputs(3382) <= a or b;
    layer0_outputs(3383) <= a;
    layer0_outputs(3384) <= not b or a;
    layer0_outputs(3385) <= a or b;
    layer0_outputs(3386) <= a or b;
    layer0_outputs(3387) <= not (a or b);
    layer0_outputs(3388) <= a or b;
    layer0_outputs(3389) <= not (a and b);
    layer0_outputs(3390) <= not (a or b);
    layer0_outputs(3391) <= not b;
    layer0_outputs(3392) <= a and not b;
    layer0_outputs(3393) <= a or b;
    layer0_outputs(3394) <= b;
    layer0_outputs(3395) <= b;
    layer0_outputs(3396) <= 1'b1;
    layer0_outputs(3397) <= a xor b;
    layer0_outputs(3398) <= a or b;
    layer0_outputs(3399) <= not b;
    layer0_outputs(3400) <= not a;
    layer0_outputs(3401) <= not b or a;
    layer0_outputs(3402) <= a or b;
    layer0_outputs(3403) <= not a or b;
    layer0_outputs(3404) <= not b or a;
    layer0_outputs(3405) <= a and not b;
    layer0_outputs(3406) <= not b;
    layer0_outputs(3407) <= not (a or b);
    layer0_outputs(3408) <= not b or a;
    layer0_outputs(3409) <= a xor b;
    layer0_outputs(3410) <= not b or a;
    layer0_outputs(3411) <= a;
    layer0_outputs(3412) <= not b;
    layer0_outputs(3413) <= not b;
    layer0_outputs(3414) <= not (a xor b);
    layer0_outputs(3415) <= a or b;
    layer0_outputs(3416) <= not b or a;
    layer0_outputs(3417) <= not b or a;
    layer0_outputs(3418) <= not (a and b);
    layer0_outputs(3419) <= not a;
    layer0_outputs(3420) <= b;
    layer0_outputs(3421) <= not a or b;
    layer0_outputs(3422) <= not (a and b);
    layer0_outputs(3423) <= not b or a;
    layer0_outputs(3424) <= 1'b0;
    layer0_outputs(3425) <= not a;
    layer0_outputs(3426) <= a xor b;
    layer0_outputs(3427) <= not (a xor b);
    layer0_outputs(3428) <= not a;
    layer0_outputs(3429) <= not a or b;
    layer0_outputs(3430) <= a and b;
    layer0_outputs(3431) <= not (a or b);
    layer0_outputs(3432) <= a and not b;
    layer0_outputs(3433) <= not b or a;
    layer0_outputs(3434) <= 1'b0;
    layer0_outputs(3435) <= 1'b0;
    layer0_outputs(3436) <= not b or a;
    layer0_outputs(3437) <= not (a xor b);
    layer0_outputs(3438) <= not (a or b);
    layer0_outputs(3439) <= a or b;
    layer0_outputs(3440) <= not (a xor b);
    layer0_outputs(3441) <= a;
    layer0_outputs(3442) <= a or b;
    layer0_outputs(3443) <= not a or b;
    layer0_outputs(3444) <= a xor b;
    layer0_outputs(3445) <= not (a or b);
    layer0_outputs(3446) <= not (a xor b);
    layer0_outputs(3447) <= a;
    layer0_outputs(3448) <= a;
    layer0_outputs(3449) <= not (a and b);
    layer0_outputs(3450) <= a and not b;
    layer0_outputs(3451) <= not a or b;
    layer0_outputs(3452) <= 1'b1;
    layer0_outputs(3453) <= not a or b;
    layer0_outputs(3454) <= not b or a;
    layer0_outputs(3455) <= not a;
    layer0_outputs(3456) <= a;
    layer0_outputs(3457) <= a and not b;
    layer0_outputs(3458) <= a;
    layer0_outputs(3459) <= a xor b;
    layer0_outputs(3460) <= a and not b;
    layer0_outputs(3461) <= not (a or b);
    layer0_outputs(3462) <= a or b;
    layer0_outputs(3463) <= not a;
    layer0_outputs(3464) <= not (a xor b);
    layer0_outputs(3465) <= a or b;
    layer0_outputs(3466) <= a or b;
    layer0_outputs(3467) <= a or b;
    layer0_outputs(3468) <= b;
    layer0_outputs(3469) <= not a;
    layer0_outputs(3470) <= a or b;
    layer0_outputs(3471) <= not a;
    layer0_outputs(3472) <= not a or b;
    layer0_outputs(3473) <= a and not b;
    layer0_outputs(3474) <= a and b;
    layer0_outputs(3475) <= b and not a;
    layer0_outputs(3476) <= not a or b;
    layer0_outputs(3477) <= a and not b;
    layer0_outputs(3478) <= not a or b;
    layer0_outputs(3479) <= not a or b;
    layer0_outputs(3480) <= a and b;
    layer0_outputs(3481) <= not b;
    layer0_outputs(3482) <= not b or a;
    layer0_outputs(3483) <= not b or a;
    layer0_outputs(3484) <= a xor b;
    layer0_outputs(3485) <= a and not b;
    layer0_outputs(3486) <= b and not a;
    layer0_outputs(3487) <= not (a or b);
    layer0_outputs(3488) <= not b or a;
    layer0_outputs(3489) <= not (a or b);
    layer0_outputs(3490) <= a or b;
    layer0_outputs(3491) <= a or b;
    layer0_outputs(3492) <= not (a or b);
    layer0_outputs(3493) <= a xor b;
    layer0_outputs(3494) <= a xor b;
    layer0_outputs(3495) <= b;
    layer0_outputs(3496) <= a;
    layer0_outputs(3497) <= not (a or b);
    layer0_outputs(3498) <= not (a or b);
    layer0_outputs(3499) <= a xor b;
    layer0_outputs(3500) <= not b or a;
    layer0_outputs(3501) <= not a;
    layer0_outputs(3502) <= not (a or b);
    layer0_outputs(3503) <= not b;
    layer0_outputs(3504) <= a;
    layer0_outputs(3505) <= b and not a;
    layer0_outputs(3506) <= b;
    layer0_outputs(3507) <= not (a or b);
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= b;
    layer0_outputs(3510) <= not (a and b);
    layer0_outputs(3511) <= not (a xor b);
    layer0_outputs(3512) <= not (a xor b);
    layer0_outputs(3513) <= a or b;
    layer0_outputs(3514) <= not a;
    layer0_outputs(3515) <= a and b;
    layer0_outputs(3516) <= not b;
    layer0_outputs(3517) <= not (a or b);
    layer0_outputs(3518) <= not b or a;
    layer0_outputs(3519) <= a xor b;
    layer0_outputs(3520) <= not a or b;
    layer0_outputs(3521) <= b and not a;
    layer0_outputs(3522) <= b and not a;
    layer0_outputs(3523) <= a and not b;
    layer0_outputs(3524) <= not a or b;
    layer0_outputs(3525) <= a and not b;
    layer0_outputs(3526) <= not (a xor b);
    layer0_outputs(3527) <= not b;
    layer0_outputs(3528) <= not (a or b);
    layer0_outputs(3529) <= a or b;
    layer0_outputs(3530) <= a or b;
    layer0_outputs(3531) <= not b;
    layer0_outputs(3532) <= not a or b;
    layer0_outputs(3533) <= b and not a;
    layer0_outputs(3534) <= not a;
    layer0_outputs(3535) <= a xor b;
    layer0_outputs(3536) <= a or b;
    layer0_outputs(3537) <= not b;
    layer0_outputs(3538) <= a and b;
    layer0_outputs(3539) <= not (a or b);
    layer0_outputs(3540) <= a or b;
    layer0_outputs(3541) <= not a;
    layer0_outputs(3542) <= not (a or b);
    layer0_outputs(3543) <= a and not b;
    layer0_outputs(3544) <= a;
    layer0_outputs(3545) <= 1'b1;
    layer0_outputs(3546) <= not (a or b);
    layer0_outputs(3547) <= not (a xor b);
    layer0_outputs(3548) <= b;
    layer0_outputs(3549) <= not b;
    layer0_outputs(3550) <= not (a xor b);
    layer0_outputs(3551) <= a and not b;
    layer0_outputs(3552) <= a;
    layer0_outputs(3553) <= a xor b;
    layer0_outputs(3554) <= b and not a;
    layer0_outputs(3555) <= not (a or b);
    layer0_outputs(3556) <= not (a or b);
    layer0_outputs(3557) <= not a;
    layer0_outputs(3558) <= not (a or b);
    layer0_outputs(3559) <= a or b;
    layer0_outputs(3560) <= not (a or b);
    layer0_outputs(3561) <= not (a xor b);
    layer0_outputs(3562) <= b;
    layer0_outputs(3563) <= not a;
    layer0_outputs(3564) <= a or b;
    layer0_outputs(3565) <= not b;
    layer0_outputs(3566) <= b;
    layer0_outputs(3567) <= not b or a;
    layer0_outputs(3568) <= b and not a;
    layer0_outputs(3569) <= a and not b;
    layer0_outputs(3570) <= a or b;
    layer0_outputs(3571) <= not a or b;
    layer0_outputs(3572) <= not b;
    layer0_outputs(3573) <= a xor b;
    layer0_outputs(3574) <= not a;
    layer0_outputs(3575) <= not b or a;
    layer0_outputs(3576) <= b and not a;
    layer0_outputs(3577) <= not (a xor b);
    layer0_outputs(3578) <= not b or a;
    layer0_outputs(3579) <= 1'b0;
    layer0_outputs(3580) <= a xor b;
    layer0_outputs(3581) <= not (a or b);
    layer0_outputs(3582) <= not (a or b);
    layer0_outputs(3583) <= not a;
    layer0_outputs(3584) <= a and b;
    layer0_outputs(3585) <= not (a or b);
    layer0_outputs(3586) <= 1'b1;
    layer0_outputs(3587) <= b;
    layer0_outputs(3588) <= b;
    layer0_outputs(3589) <= not (a or b);
    layer0_outputs(3590) <= not (a or b);
    layer0_outputs(3591) <= a and not b;
    layer0_outputs(3592) <= not a;
    layer0_outputs(3593) <= a xor b;
    layer0_outputs(3594) <= not b;
    layer0_outputs(3595) <= not a or b;
    layer0_outputs(3596) <= not b;
    layer0_outputs(3597) <= b;
    layer0_outputs(3598) <= a or b;
    layer0_outputs(3599) <= not (a xor b);
    layer0_outputs(3600) <= a or b;
    layer0_outputs(3601) <= a;
    layer0_outputs(3602) <= a or b;
    layer0_outputs(3603) <= not a or b;
    layer0_outputs(3604) <= a;
    layer0_outputs(3605) <= not (a or b);
    layer0_outputs(3606) <= not (a xor b);
    layer0_outputs(3607) <= a;
    layer0_outputs(3608) <= b;
    layer0_outputs(3609) <= not (a xor b);
    layer0_outputs(3610) <= a or b;
    layer0_outputs(3611) <= a or b;
    layer0_outputs(3612) <= not a;
    layer0_outputs(3613) <= a or b;
    layer0_outputs(3614) <= not a or b;
    layer0_outputs(3615) <= a;
    layer0_outputs(3616) <= a and not b;
    layer0_outputs(3617) <= not (a or b);
    layer0_outputs(3618) <= a or b;
    layer0_outputs(3619) <= a or b;
    layer0_outputs(3620) <= b;
    layer0_outputs(3621) <= a or b;
    layer0_outputs(3622) <= a xor b;
    layer0_outputs(3623) <= not (a or b);
    layer0_outputs(3624) <= not a;
    layer0_outputs(3625) <= not b;
    layer0_outputs(3626) <= a;
    layer0_outputs(3627) <= a or b;
    layer0_outputs(3628) <= not (a or b);
    layer0_outputs(3629) <= b and not a;
    layer0_outputs(3630) <= not b or a;
    layer0_outputs(3631) <= not (a or b);
    layer0_outputs(3632) <= a and not b;
    layer0_outputs(3633) <= not b or a;
    layer0_outputs(3634) <= b and not a;
    layer0_outputs(3635) <= not a;
    layer0_outputs(3636) <= a;
    layer0_outputs(3637) <= 1'b0;
    layer0_outputs(3638) <= not (a or b);
    layer0_outputs(3639) <= not b or a;
    layer0_outputs(3640) <= not a or b;
    layer0_outputs(3641) <= a and b;
    layer0_outputs(3642) <= a or b;
    layer0_outputs(3643) <= not (a or b);
    layer0_outputs(3644) <= not (a or b);
    layer0_outputs(3645) <= not (a xor b);
    layer0_outputs(3646) <= 1'b1;
    layer0_outputs(3647) <= a and b;
    layer0_outputs(3648) <= 1'b1;
    layer0_outputs(3649) <= a and b;
    layer0_outputs(3650) <= not (a xor b);
    layer0_outputs(3651) <= 1'b0;
    layer0_outputs(3652) <= not (a or b);
    layer0_outputs(3653) <= not b;
    layer0_outputs(3654) <= a xor b;
    layer0_outputs(3655) <= not b or a;
    layer0_outputs(3656) <= a;
    layer0_outputs(3657) <= not a;
    layer0_outputs(3658) <= a or b;
    layer0_outputs(3659) <= not b;
    layer0_outputs(3660) <= not b or a;
    layer0_outputs(3661) <= a or b;
    layer0_outputs(3662) <= not a;
    layer0_outputs(3663) <= a and not b;
    layer0_outputs(3664) <= not b or a;
    layer0_outputs(3665) <= not a;
    layer0_outputs(3666) <= a or b;
    layer0_outputs(3667) <= a or b;
    layer0_outputs(3668) <= a xor b;
    layer0_outputs(3669) <= not b;
    layer0_outputs(3670) <= a and not b;
    layer0_outputs(3671) <= b and not a;
    layer0_outputs(3672) <= a and not b;
    layer0_outputs(3673) <= a and b;
    layer0_outputs(3674) <= a or b;
    layer0_outputs(3675) <= b and not a;
    layer0_outputs(3676) <= not a or b;
    layer0_outputs(3677) <= a xor b;
    layer0_outputs(3678) <= a;
    layer0_outputs(3679) <= a;
    layer0_outputs(3680) <= not a or b;
    layer0_outputs(3681) <= not (a xor b);
    layer0_outputs(3682) <= not b;
    layer0_outputs(3683) <= not (a and b);
    layer0_outputs(3684) <= b and not a;
    layer0_outputs(3685) <= b and not a;
    layer0_outputs(3686) <= not (a and b);
    layer0_outputs(3687) <= a or b;
    layer0_outputs(3688) <= not (a xor b);
    layer0_outputs(3689) <= not (a xor b);
    layer0_outputs(3690) <= b;
    layer0_outputs(3691) <= not a or b;
    layer0_outputs(3692) <= a or b;
    layer0_outputs(3693) <= a and not b;
    layer0_outputs(3694) <= not (a or b);
    layer0_outputs(3695) <= not (a or b);
    layer0_outputs(3696) <= not a or b;
    layer0_outputs(3697) <= a or b;
    layer0_outputs(3698) <= a xor b;
    layer0_outputs(3699) <= a xor b;
    layer0_outputs(3700) <= a;
    layer0_outputs(3701) <= not (a or b);
    layer0_outputs(3702) <= a or b;
    layer0_outputs(3703) <= a or b;
    layer0_outputs(3704) <= not (a or b);
    layer0_outputs(3705) <= a and b;
    layer0_outputs(3706) <= b;
    layer0_outputs(3707) <= not a or b;
    layer0_outputs(3708) <= b and not a;
    layer0_outputs(3709) <= a;
    layer0_outputs(3710) <= not a or b;
    layer0_outputs(3711) <= b and not a;
    layer0_outputs(3712) <= 1'b0;
    layer0_outputs(3713) <= a or b;
    layer0_outputs(3714) <= a;
    layer0_outputs(3715) <= a or b;
    layer0_outputs(3716) <= b and not a;
    layer0_outputs(3717) <= not (a or b);
    layer0_outputs(3718) <= not a or b;
    layer0_outputs(3719) <= not (a or b);
    layer0_outputs(3720) <= a or b;
    layer0_outputs(3721) <= not b or a;
    layer0_outputs(3722) <= a;
    layer0_outputs(3723) <= not (a or b);
    layer0_outputs(3724) <= a xor b;
    layer0_outputs(3725) <= not a;
    layer0_outputs(3726) <= not (a and b);
    layer0_outputs(3727) <= not b or a;
    layer0_outputs(3728) <= a and not b;
    layer0_outputs(3729) <= b;
    layer0_outputs(3730) <= not b or a;
    layer0_outputs(3731) <= not a;
    layer0_outputs(3732) <= b;
    layer0_outputs(3733) <= b;
    layer0_outputs(3734) <= a xor b;
    layer0_outputs(3735) <= not b or a;
    layer0_outputs(3736) <= not (a or b);
    layer0_outputs(3737) <= 1'b0;
    layer0_outputs(3738) <= not (a or b);
    layer0_outputs(3739) <= a and not b;
    layer0_outputs(3740) <= not a;
    layer0_outputs(3741) <= not b;
    layer0_outputs(3742) <= not (a and b);
    layer0_outputs(3743) <= a;
    layer0_outputs(3744) <= a and not b;
    layer0_outputs(3745) <= not a;
    layer0_outputs(3746) <= not (a xor b);
    layer0_outputs(3747) <= not b;
    layer0_outputs(3748) <= not b or a;
    layer0_outputs(3749) <= b;
    layer0_outputs(3750) <= b;
    layer0_outputs(3751) <= not a or b;
    layer0_outputs(3752) <= not b;
    layer0_outputs(3753) <= not b;
    layer0_outputs(3754) <= b;
    layer0_outputs(3755) <= b and not a;
    layer0_outputs(3756) <= not b;
    layer0_outputs(3757) <= a or b;
    layer0_outputs(3758) <= not (a xor b);
    layer0_outputs(3759) <= a and not b;
    layer0_outputs(3760) <= not b or a;
    layer0_outputs(3761) <= b;
    layer0_outputs(3762) <= a and not b;
    layer0_outputs(3763) <= a xor b;
    layer0_outputs(3764) <= not a or b;
    layer0_outputs(3765) <= not b;
    layer0_outputs(3766) <= a;
    layer0_outputs(3767) <= not a or b;
    layer0_outputs(3768) <= a or b;
    layer0_outputs(3769) <= not b or a;
    layer0_outputs(3770) <= a or b;
    layer0_outputs(3771) <= not (a or b);
    layer0_outputs(3772) <= a xor b;
    layer0_outputs(3773) <= 1'b0;
    layer0_outputs(3774) <= not (a xor b);
    layer0_outputs(3775) <= not a;
    layer0_outputs(3776) <= not (a or b);
    layer0_outputs(3777) <= a and b;
    layer0_outputs(3778) <= not b or a;
    layer0_outputs(3779) <= a;
    layer0_outputs(3780) <= a and not b;
    layer0_outputs(3781) <= not (a or b);
    layer0_outputs(3782) <= a xor b;
    layer0_outputs(3783) <= not a;
    layer0_outputs(3784) <= not (a or b);
    layer0_outputs(3785) <= not b or a;
    layer0_outputs(3786) <= not (a or b);
    layer0_outputs(3787) <= not a;
    layer0_outputs(3788) <= not b or a;
    layer0_outputs(3789) <= not a or b;
    layer0_outputs(3790) <= a or b;
    layer0_outputs(3791) <= not b or a;
    layer0_outputs(3792) <= a;
    layer0_outputs(3793) <= b;
    layer0_outputs(3794) <= a or b;
    layer0_outputs(3795) <= not a;
    layer0_outputs(3796) <= a or b;
    layer0_outputs(3797) <= not (a or b);
    layer0_outputs(3798) <= 1'b0;
    layer0_outputs(3799) <= a xor b;
    layer0_outputs(3800) <= 1'b1;
    layer0_outputs(3801) <= b and not a;
    layer0_outputs(3802) <= not b;
    layer0_outputs(3803) <= a;
    layer0_outputs(3804) <= b;
    layer0_outputs(3805) <= a xor b;
    layer0_outputs(3806) <= not (a and b);
    layer0_outputs(3807) <= b;
    layer0_outputs(3808) <= not (a or b);
    layer0_outputs(3809) <= not b or a;
    layer0_outputs(3810) <= 1'b1;
    layer0_outputs(3811) <= not (a or b);
    layer0_outputs(3812) <= a xor b;
    layer0_outputs(3813) <= a or b;
    layer0_outputs(3814) <= not (a xor b);
    layer0_outputs(3815) <= b and not a;
    layer0_outputs(3816) <= not (a xor b);
    layer0_outputs(3817) <= not (a or b);
    layer0_outputs(3818) <= not (a or b);
    layer0_outputs(3819) <= a;
    layer0_outputs(3820) <= not b;
    layer0_outputs(3821) <= not b or a;
    layer0_outputs(3822) <= not b;
    layer0_outputs(3823) <= not (a or b);
    layer0_outputs(3824) <= a or b;
    layer0_outputs(3825) <= a xor b;
    layer0_outputs(3826) <= a and not b;
    layer0_outputs(3827) <= b;
    layer0_outputs(3828) <= a xor b;
    layer0_outputs(3829) <= not (a or b);
    layer0_outputs(3830) <= a and not b;
    layer0_outputs(3831) <= a or b;
    layer0_outputs(3832) <= not (a or b);
    layer0_outputs(3833) <= not (a and b);
    layer0_outputs(3834) <= b;
    layer0_outputs(3835) <= a or b;
    layer0_outputs(3836) <= b and not a;
    layer0_outputs(3837) <= not (a and b);
    layer0_outputs(3838) <= a or b;
    layer0_outputs(3839) <= a or b;
    layer0_outputs(3840) <= a or b;
    layer0_outputs(3841) <= not b or a;
    layer0_outputs(3842) <= not b or a;
    layer0_outputs(3843) <= a and not b;
    layer0_outputs(3844) <= a or b;
    layer0_outputs(3845) <= not b or a;
    layer0_outputs(3846) <= 1'b0;
    layer0_outputs(3847) <= a xor b;
    layer0_outputs(3848) <= a or b;
    layer0_outputs(3849) <= a;
    layer0_outputs(3850) <= a or b;
    layer0_outputs(3851) <= a or b;
    layer0_outputs(3852) <= b;
    layer0_outputs(3853) <= not b;
    layer0_outputs(3854) <= not b;
    layer0_outputs(3855) <= not a;
    layer0_outputs(3856) <= b and not a;
    layer0_outputs(3857) <= not a;
    layer0_outputs(3858) <= 1'b0;
    layer0_outputs(3859) <= b;
    layer0_outputs(3860) <= not (a xor b);
    layer0_outputs(3861) <= a;
    layer0_outputs(3862) <= a or b;
    layer0_outputs(3863) <= b;
    layer0_outputs(3864) <= 1'b1;
    layer0_outputs(3865) <= a and b;
    layer0_outputs(3866) <= a or b;
    layer0_outputs(3867) <= a;
    layer0_outputs(3868) <= not a;
    layer0_outputs(3869) <= not (a or b);
    layer0_outputs(3870) <= not (a or b);
    layer0_outputs(3871) <= a or b;
    layer0_outputs(3872) <= a;
    layer0_outputs(3873) <= not b;
    layer0_outputs(3874) <= a;
    layer0_outputs(3875) <= a or b;
    layer0_outputs(3876) <= b and not a;
    layer0_outputs(3877) <= a xor b;
    layer0_outputs(3878) <= b;
    layer0_outputs(3879) <= b and not a;
    layer0_outputs(3880) <= not b or a;
    layer0_outputs(3881) <= not b or a;
    layer0_outputs(3882) <= not (a xor b);
    layer0_outputs(3883) <= not b;
    layer0_outputs(3884) <= not b;
    layer0_outputs(3885) <= a;
    layer0_outputs(3886) <= not (a or b);
    layer0_outputs(3887) <= not (a or b);
    layer0_outputs(3888) <= not (a or b);
    layer0_outputs(3889) <= not a or b;
    layer0_outputs(3890) <= 1'b1;
    layer0_outputs(3891) <= a and not b;
    layer0_outputs(3892) <= a and not b;
    layer0_outputs(3893) <= a or b;
    layer0_outputs(3894) <= not b or a;
    layer0_outputs(3895) <= a;
    layer0_outputs(3896) <= a;
    layer0_outputs(3897) <= not (a and b);
    layer0_outputs(3898) <= b and not a;
    layer0_outputs(3899) <= a xor b;
    layer0_outputs(3900) <= b and not a;
    layer0_outputs(3901) <= not b or a;
    layer0_outputs(3902) <= not a or b;
    layer0_outputs(3903) <= not a or b;
    layer0_outputs(3904) <= a or b;
    layer0_outputs(3905) <= a or b;
    layer0_outputs(3906) <= a and not b;
    layer0_outputs(3907) <= 1'b0;
    layer0_outputs(3908) <= not (a xor b);
    layer0_outputs(3909) <= not b or a;
    layer0_outputs(3910) <= a and not b;
    layer0_outputs(3911) <= not (a xor b);
    layer0_outputs(3912) <= not (a or b);
    layer0_outputs(3913) <= not a or b;
    layer0_outputs(3914) <= not a;
    layer0_outputs(3915) <= not (a or b);
    layer0_outputs(3916) <= a and not b;
    layer0_outputs(3917) <= not b or a;
    layer0_outputs(3918) <= a xor b;
    layer0_outputs(3919) <= not b;
    layer0_outputs(3920) <= not a or b;
    layer0_outputs(3921) <= not (a or b);
    layer0_outputs(3922) <= not (a or b);
    layer0_outputs(3923) <= not (a or b);
    layer0_outputs(3924) <= not a;
    layer0_outputs(3925) <= b and not a;
    layer0_outputs(3926) <= not a or b;
    layer0_outputs(3927) <= a;
    layer0_outputs(3928) <= a or b;
    layer0_outputs(3929) <= not (a xor b);
    layer0_outputs(3930) <= not (a or b);
    layer0_outputs(3931) <= a and not b;
    layer0_outputs(3932) <= not a or b;
    layer0_outputs(3933) <= not b;
    layer0_outputs(3934) <= a or b;
    layer0_outputs(3935) <= not b or a;
    layer0_outputs(3936) <= a xor b;
    layer0_outputs(3937) <= not (a or b);
    layer0_outputs(3938) <= not a;
    layer0_outputs(3939) <= not b;
    layer0_outputs(3940) <= not a;
    layer0_outputs(3941) <= not (a and b);
    layer0_outputs(3942) <= not (a or b);
    layer0_outputs(3943) <= not b;
    layer0_outputs(3944) <= not (a xor b);
    layer0_outputs(3945) <= not (a and b);
    layer0_outputs(3946) <= not (a and b);
    layer0_outputs(3947) <= not b or a;
    layer0_outputs(3948) <= a or b;
    layer0_outputs(3949) <= b;
    layer0_outputs(3950) <= not a;
    layer0_outputs(3951) <= a xor b;
    layer0_outputs(3952) <= not (a or b);
    layer0_outputs(3953) <= a or b;
    layer0_outputs(3954) <= b;
    layer0_outputs(3955) <= not b or a;
    layer0_outputs(3956) <= not (a or b);
    layer0_outputs(3957) <= not a or b;
    layer0_outputs(3958) <= a and b;
    layer0_outputs(3959) <= 1'b0;
    layer0_outputs(3960) <= a;
    layer0_outputs(3961) <= b;
    layer0_outputs(3962) <= not a or b;
    layer0_outputs(3963) <= a xor b;
    layer0_outputs(3964) <= a or b;
    layer0_outputs(3965) <= not b;
    layer0_outputs(3966) <= not (a or b);
    layer0_outputs(3967) <= not b;
    layer0_outputs(3968) <= not (a or b);
    layer0_outputs(3969) <= 1'b1;
    layer0_outputs(3970) <= not (a or b);
    layer0_outputs(3971) <= not a or b;
    layer0_outputs(3972) <= a;
    layer0_outputs(3973) <= not b;
    layer0_outputs(3974) <= b;
    layer0_outputs(3975) <= not a;
    layer0_outputs(3976) <= not (a xor b);
    layer0_outputs(3977) <= a xor b;
    layer0_outputs(3978) <= not (a and b);
    layer0_outputs(3979) <= a;
    layer0_outputs(3980) <= b;
    layer0_outputs(3981) <= not (a or b);
    layer0_outputs(3982) <= not (a or b);
    layer0_outputs(3983) <= not (a or b);
    layer0_outputs(3984) <= not a;
    layer0_outputs(3985) <= a;
    layer0_outputs(3986) <= a or b;
    layer0_outputs(3987) <= not (a and b);
    layer0_outputs(3988) <= b;
    layer0_outputs(3989) <= a xor b;
    layer0_outputs(3990) <= a or b;
    layer0_outputs(3991) <= a or b;
    layer0_outputs(3992) <= a xor b;
    layer0_outputs(3993) <= a and not b;
    layer0_outputs(3994) <= not (a and b);
    layer0_outputs(3995) <= a and not b;
    layer0_outputs(3996) <= b and not a;
    layer0_outputs(3997) <= a or b;
    layer0_outputs(3998) <= not a or b;
    layer0_outputs(3999) <= b;
    layer0_outputs(4000) <= b;
    layer0_outputs(4001) <= a or b;
    layer0_outputs(4002) <= not (a and b);
    layer0_outputs(4003) <= not (a or b);
    layer0_outputs(4004) <= not (a or b);
    layer0_outputs(4005) <= not a or b;
    layer0_outputs(4006) <= not (a or b);
    layer0_outputs(4007) <= not (a xor b);
    layer0_outputs(4008) <= 1'b1;
    layer0_outputs(4009) <= not a or b;
    layer0_outputs(4010) <= not a;
    layer0_outputs(4011) <= a or b;
    layer0_outputs(4012) <= not a;
    layer0_outputs(4013) <= not a;
    layer0_outputs(4014) <= a and not b;
    layer0_outputs(4015) <= a and not b;
    layer0_outputs(4016) <= b;
    layer0_outputs(4017) <= not a or b;
    layer0_outputs(4018) <= a xor b;
    layer0_outputs(4019) <= a xor b;
    layer0_outputs(4020) <= not (a or b);
    layer0_outputs(4021) <= b and not a;
    layer0_outputs(4022) <= not b;
    layer0_outputs(4023) <= not b or a;
    layer0_outputs(4024) <= a or b;
    layer0_outputs(4025) <= not a or b;
    layer0_outputs(4026) <= b;
    layer0_outputs(4027) <= not a or b;
    layer0_outputs(4028) <= not (a and b);
    layer0_outputs(4029) <= a or b;
    layer0_outputs(4030) <= not (a xor b);
    layer0_outputs(4031) <= a and not b;
    layer0_outputs(4032) <= a;
    layer0_outputs(4033) <= a or b;
    layer0_outputs(4034) <= b and not a;
    layer0_outputs(4035) <= a or b;
    layer0_outputs(4036) <= a xor b;
    layer0_outputs(4037) <= not a;
    layer0_outputs(4038) <= a;
    layer0_outputs(4039) <= not a;
    layer0_outputs(4040) <= a and b;
    layer0_outputs(4041) <= not a or b;
    layer0_outputs(4042) <= not (a or b);
    layer0_outputs(4043) <= a;
    layer0_outputs(4044) <= a and not b;
    layer0_outputs(4045) <= b;
    layer0_outputs(4046) <= not (a xor b);
    layer0_outputs(4047) <= a;
    layer0_outputs(4048) <= not a;
    layer0_outputs(4049) <= b and not a;
    layer0_outputs(4050) <= a xor b;
    layer0_outputs(4051) <= a;
    layer0_outputs(4052) <= b;
    layer0_outputs(4053) <= b and not a;
    layer0_outputs(4054) <= not (a or b);
    layer0_outputs(4055) <= a;
    layer0_outputs(4056) <= not (a or b);
    layer0_outputs(4057) <= not b or a;
    layer0_outputs(4058) <= not b;
    layer0_outputs(4059) <= not (a xor b);
    layer0_outputs(4060) <= b;
    layer0_outputs(4061) <= not b;
    layer0_outputs(4062) <= b;
    layer0_outputs(4063) <= not (a xor b);
    layer0_outputs(4064) <= a and not b;
    layer0_outputs(4065) <= not (a and b);
    layer0_outputs(4066) <= not a or b;
    layer0_outputs(4067) <= not a or b;
    layer0_outputs(4068) <= not b;
    layer0_outputs(4069) <= b and not a;
    layer0_outputs(4070) <= a and not b;
    layer0_outputs(4071) <= a or b;
    layer0_outputs(4072) <= not (a or b);
    layer0_outputs(4073) <= not b;
    layer0_outputs(4074) <= not a or b;
    layer0_outputs(4075) <= not a or b;
    layer0_outputs(4076) <= a;
    layer0_outputs(4077) <= a or b;
    layer0_outputs(4078) <= a and b;
    layer0_outputs(4079) <= not (a or b);
    layer0_outputs(4080) <= not (a or b);
    layer0_outputs(4081) <= not b or a;
    layer0_outputs(4082) <= 1'b0;
    layer0_outputs(4083) <= a and b;
    layer0_outputs(4084) <= not a or b;
    layer0_outputs(4085) <= not b or a;
    layer0_outputs(4086) <= a and not b;
    layer0_outputs(4087) <= not a or b;
    layer0_outputs(4088) <= not (a xor b);
    layer0_outputs(4089) <= b and not a;
    layer0_outputs(4090) <= not a;
    layer0_outputs(4091) <= not (a or b);
    layer0_outputs(4092) <= b;
    layer0_outputs(4093) <= not b;
    layer0_outputs(4094) <= not (a and b);
    layer0_outputs(4095) <= a or b;
    layer0_outputs(4096) <= a or b;
    layer0_outputs(4097) <= b;
    layer0_outputs(4098) <= not (a xor b);
    layer0_outputs(4099) <= a;
    layer0_outputs(4100) <= a;
    layer0_outputs(4101) <= not a or b;
    layer0_outputs(4102) <= not a;
    layer0_outputs(4103) <= not a or b;
    layer0_outputs(4104) <= 1'b0;
    layer0_outputs(4105) <= a;
    layer0_outputs(4106) <= not (a xor b);
    layer0_outputs(4107) <= not b or a;
    layer0_outputs(4108) <= b;
    layer0_outputs(4109) <= not (a xor b);
    layer0_outputs(4110) <= a xor b;
    layer0_outputs(4111) <= not a;
    layer0_outputs(4112) <= a or b;
    layer0_outputs(4113) <= a and b;
    layer0_outputs(4114) <= a and not b;
    layer0_outputs(4115) <= not a or b;
    layer0_outputs(4116) <= a or b;
    layer0_outputs(4117) <= b;
    layer0_outputs(4118) <= not b;
    layer0_outputs(4119) <= a xor b;
    layer0_outputs(4120) <= a or b;
    layer0_outputs(4121) <= not a or b;
    layer0_outputs(4122) <= a xor b;
    layer0_outputs(4123) <= 1'b1;
    layer0_outputs(4124) <= a or b;
    layer0_outputs(4125) <= a and not b;
    layer0_outputs(4126) <= a or b;
    layer0_outputs(4127) <= not (a xor b);
    layer0_outputs(4128) <= a xor b;
    layer0_outputs(4129) <= b;
    layer0_outputs(4130) <= not b or a;
    layer0_outputs(4131) <= not (a and b);
    layer0_outputs(4132) <= not b or a;
    layer0_outputs(4133) <= 1'b0;
    layer0_outputs(4134) <= a xor b;
    layer0_outputs(4135) <= b;
    layer0_outputs(4136) <= not (a or b);
    layer0_outputs(4137) <= not (a xor b);
    layer0_outputs(4138) <= b and not a;
    layer0_outputs(4139) <= not b;
    layer0_outputs(4140) <= 1'b0;
    layer0_outputs(4141) <= not a or b;
    layer0_outputs(4142) <= a or b;
    layer0_outputs(4143) <= a or b;
    layer0_outputs(4144) <= a and not b;
    layer0_outputs(4145) <= not (a xor b);
    layer0_outputs(4146) <= not a or b;
    layer0_outputs(4147) <= not (a xor b);
    layer0_outputs(4148) <= not b or a;
    layer0_outputs(4149) <= b;
    layer0_outputs(4150) <= not (a and b);
    layer0_outputs(4151) <= a and not b;
    layer0_outputs(4152) <= b and not a;
    layer0_outputs(4153) <= not a or b;
    layer0_outputs(4154) <= a or b;
    layer0_outputs(4155) <= not b;
    layer0_outputs(4156) <= b;
    layer0_outputs(4157) <= a and not b;
    layer0_outputs(4158) <= not a or b;
    layer0_outputs(4159) <= b and not a;
    layer0_outputs(4160) <= b and not a;
    layer0_outputs(4161) <= not a;
    layer0_outputs(4162) <= 1'b0;
    layer0_outputs(4163) <= a xor b;
    layer0_outputs(4164) <= not b or a;
    layer0_outputs(4165) <= not (a or b);
    layer0_outputs(4166) <= a and not b;
    layer0_outputs(4167) <= not b or a;
    layer0_outputs(4168) <= not a;
    layer0_outputs(4169) <= not (a or b);
    layer0_outputs(4170) <= 1'b1;
    layer0_outputs(4171) <= not b or a;
    layer0_outputs(4172) <= not (a or b);
    layer0_outputs(4173) <= not (a xor b);
    layer0_outputs(4174) <= b;
    layer0_outputs(4175) <= a or b;
    layer0_outputs(4176) <= b;
    layer0_outputs(4177) <= a;
    layer0_outputs(4178) <= a and not b;
    layer0_outputs(4179) <= b;
    layer0_outputs(4180) <= not b;
    layer0_outputs(4181) <= a;
    layer0_outputs(4182) <= a xor b;
    layer0_outputs(4183) <= not b or a;
    layer0_outputs(4184) <= a;
    layer0_outputs(4185) <= a and not b;
    layer0_outputs(4186) <= a;
    layer0_outputs(4187) <= a xor b;
    layer0_outputs(4188) <= not (a xor b);
    layer0_outputs(4189) <= not a;
    layer0_outputs(4190) <= b and not a;
    layer0_outputs(4191) <= not (a xor b);
    layer0_outputs(4192) <= a or b;
    layer0_outputs(4193) <= a and not b;
    layer0_outputs(4194) <= a or b;
    layer0_outputs(4195) <= a and not b;
    layer0_outputs(4196) <= not (a or b);
    layer0_outputs(4197) <= not a or b;
    layer0_outputs(4198) <= not (a xor b);
    layer0_outputs(4199) <= a and b;
    layer0_outputs(4200) <= not a;
    layer0_outputs(4201) <= b and not a;
    layer0_outputs(4202) <= not (a or b);
    layer0_outputs(4203) <= a and b;
    layer0_outputs(4204) <= not (a or b);
    layer0_outputs(4205) <= not b;
    layer0_outputs(4206) <= 1'b0;
    layer0_outputs(4207) <= not (a xor b);
    layer0_outputs(4208) <= not b;
    layer0_outputs(4209) <= not b;
    layer0_outputs(4210) <= 1'b0;
    layer0_outputs(4211) <= 1'b0;
    layer0_outputs(4212) <= not b;
    layer0_outputs(4213) <= b;
    layer0_outputs(4214) <= not (a or b);
    layer0_outputs(4215) <= not a;
    layer0_outputs(4216) <= a xor b;
    layer0_outputs(4217) <= not (a xor b);
    layer0_outputs(4218) <= not (a or b);
    layer0_outputs(4219) <= not (a xor b);
    layer0_outputs(4220) <= not (a xor b);
    layer0_outputs(4221) <= not (a xor b);
    layer0_outputs(4222) <= not a or b;
    layer0_outputs(4223) <= b;
    layer0_outputs(4224) <= a xor b;
    layer0_outputs(4225) <= a xor b;
    layer0_outputs(4226) <= not b or a;
    layer0_outputs(4227) <= b and not a;
    layer0_outputs(4228) <= a;
    layer0_outputs(4229) <= not (a and b);
    layer0_outputs(4230) <= not b;
    layer0_outputs(4231) <= a and b;
    layer0_outputs(4232) <= a xor b;
    layer0_outputs(4233) <= 1'b1;
    layer0_outputs(4234) <= not (a or b);
    layer0_outputs(4235) <= not a or b;
    layer0_outputs(4236) <= not (a xor b);
    layer0_outputs(4237) <= a;
    layer0_outputs(4238) <= not b;
    layer0_outputs(4239) <= not (a or b);
    layer0_outputs(4240) <= not b;
    layer0_outputs(4241) <= a xor b;
    layer0_outputs(4242) <= not (a xor b);
    layer0_outputs(4243) <= not (a or b);
    layer0_outputs(4244) <= a xor b;
    layer0_outputs(4245) <= not a or b;
    layer0_outputs(4246) <= not a or b;
    layer0_outputs(4247) <= not (a and b);
    layer0_outputs(4248) <= not b;
    layer0_outputs(4249) <= not a or b;
    layer0_outputs(4250) <= not b;
    layer0_outputs(4251) <= not (a and b);
    layer0_outputs(4252) <= a;
    layer0_outputs(4253) <= not (a and b);
    layer0_outputs(4254) <= not a or b;
    layer0_outputs(4255) <= 1'b0;
    layer0_outputs(4256) <= a or b;
    layer0_outputs(4257) <= a and b;
    layer0_outputs(4258) <= a or b;
    layer0_outputs(4259) <= a xor b;
    layer0_outputs(4260) <= not (a or b);
    layer0_outputs(4261) <= not (a or b);
    layer0_outputs(4262) <= 1'b0;
    layer0_outputs(4263) <= not (a xor b);
    layer0_outputs(4264) <= a xor b;
    layer0_outputs(4265) <= not a or b;
    layer0_outputs(4266) <= not (a xor b);
    layer0_outputs(4267) <= a and not b;
    layer0_outputs(4268) <= b;
    layer0_outputs(4269) <= b;
    layer0_outputs(4270) <= a xor b;
    layer0_outputs(4271) <= not b;
    layer0_outputs(4272) <= b and not a;
    layer0_outputs(4273) <= b;
    layer0_outputs(4274) <= a and b;
    layer0_outputs(4275) <= 1'b1;
    layer0_outputs(4276) <= not (a and b);
    layer0_outputs(4277) <= 1'b1;
    layer0_outputs(4278) <= not a;
    layer0_outputs(4279) <= a or b;
    layer0_outputs(4280) <= not a;
    layer0_outputs(4281) <= b;
    layer0_outputs(4282) <= not b;
    layer0_outputs(4283) <= a or b;
    layer0_outputs(4284) <= not (a or b);
    layer0_outputs(4285) <= 1'b0;
    layer0_outputs(4286) <= a xor b;
    layer0_outputs(4287) <= a xor b;
    layer0_outputs(4288) <= not b or a;
    layer0_outputs(4289) <= not b or a;
    layer0_outputs(4290) <= a;
    layer0_outputs(4291) <= not (a or b);
    layer0_outputs(4292) <= a and b;
    layer0_outputs(4293) <= not (a xor b);
    layer0_outputs(4294) <= not b or a;
    layer0_outputs(4295) <= not b;
    layer0_outputs(4296) <= not (a or b);
    layer0_outputs(4297) <= a or b;
    layer0_outputs(4298) <= not (a or b);
    layer0_outputs(4299) <= not (a or b);
    layer0_outputs(4300) <= not (a xor b);
    layer0_outputs(4301) <= not (a or b);
    layer0_outputs(4302) <= not a;
    layer0_outputs(4303) <= a;
    layer0_outputs(4304) <= a or b;
    layer0_outputs(4305) <= a or b;
    layer0_outputs(4306) <= a;
    layer0_outputs(4307) <= not (a xor b);
    layer0_outputs(4308) <= 1'b0;
    layer0_outputs(4309) <= a or b;
    layer0_outputs(4310) <= a xor b;
    layer0_outputs(4311) <= a or b;
    layer0_outputs(4312) <= a and not b;
    layer0_outputs(4313) <= a;
    layer0_outputs(4314) <= not b or a;
    layer0_outputs(4315) <= not b;
    layer0_outputs(4316) <= b;
    layer0_outputs(4317) <= not (a xor b);
    layer0_outputs(4318) <= a;
    layer0_outputs(4319) <= b;
    layer0_outputs(4320) <= a;
    layer0_outputs(4321) <= a xor b;
    layer0_outputs(4322) <= not b or a;
    layer0_outputs(4323) <= a xor b;
    layer0_outputs(4324) <= a xor b;
    layer0_outputs(4325) <= not a or b;
    layer0_outputs(4326) <= a;
    layer0_outputs(4327) <= a or b;
    layer0_outputs(4328) <= not b;
    layer0_outputs(4329) <= not (a xor b);
    layer0_outputs(4330) <= a or b;
    layer0_outputs(4331) <= 1'b0;
    layer0_outputs(4332) <= not (a xor b);
    layer0_outputs(4333) <= not (a xor b);
    layer0_outputs(4334) <= a or b;
    layer0_outputs(4335) <= a and b;
    layer0_outputs(4336) <= not a;
    layer0_outputs(4337) <= b;
    layer0_outputs(4338) <= a or b;
    layer0_outputs(4339) <= not (a or b);
    layer0_outputs(4340) <= a;
    layer0_outputs(4341) <= not a or b;
    layer0_outputs(4342) <= a;
    layer0_outputs(4343) <= not a or b;
    layer0_outputs(4344) <= b;
    layer0_outputs(4345) <= 1'b0;
    layer0_outputs(4346) <= a;
    layer0_outputs(4347) <= a;
    layer0_outputs(4348) <= a;
    layer0_outputs(4349) <= b;
    layer0_outputs(4350) <= a;
    layer0_outputs(4351) <= 1'b0;
    layer0_outputs(4352) <= b;
    layer0_outputs(4353) <= a and not b;
    layer0_outputs(4354) <= not (a or b);
    layer0_outputs(4355) <= not b or a;
    layer0_outputs(4356) <= a xor b;
    layer0_outputs(4357) <= b;
    layer0_outputs(4358) <= a and not b;
    layer0_outputs(4359) <= not b;
    layer0_outputs(4360) <= b and not a;
    layer0_outputs(4361) <= not a or b;
    layer0_outputs(4362) <= not (a and b);
    layer0_outputs(4363) <= not b or a;
    layer0_outputs(4364) <= a and b;
    layer0_outputs(4365) <= not (a xor b);
    layer0_outputs(4366) <= not (a xor b);
    layer0_outputs(4367) <= a xor b;
    layer0_outputs(4368) <= a or b;
    layer0_outputs(4369) <= not (a xor b);
    layer0_outputs(4370) <= not (a or b);
    layer0_outputs(4371) <= not b or a;
    layer0_outputs(4372) <= a and b;
    layer0_outputs(4373) <= a xor b;
    layer0_outputs(4374) <= a;
    layer0_outputs(4375) <= not (a xor b);
    layer0_outputs(4376) <= 1'b0;
    layer0_outputs(4377) <= not (a and b);
    layer0_outputs(4378) <= not b or a;
    layer0_outputs(4379) <= not (a or b);
    layer0_outputs(4380) <= a xor b;
    layer0_outputs(4381) <= not a or b;
    layer0_outputs(4382) <= not (a xor b);
    layer0_outputs(4383) <= a and not b;
    layer0_outputs(4384) <= b;
    layer0_outputs(4385) <= b;
    layer0_outputs(4386) <= b;
    layer0_outputs(4387) <= a and not b;
    layer0_outputs(4388) <= a;
    layer0_outputs(4389) <= not (a or b);
    layer0_outputs(4390) <= a xor b;
    layer0_outputs(4391) <= not a;
    layer0_outputs(4392) <= b;
    layer0_outputs(4393) <= not b or a;
    layer0_outputs(4394) <= a and not b;
    layer0_outputs(4395) <= b and not a;
    layer0_outputs(4396) <= a;
    layer0_outputs(4397) <= b;
    layer0_outputs(4398) <= a and not b;
    layer0_outputs(4399) <= a and not b;
    layer0_outputs(4400) <= not (a or b);
    layer0_outputs(4401) <= b;
    layer0_outputs(4402) <= a xor b;
    layer0_outputs(4403) <= not a or b;
    layer0_outputs(4404) <= not b;
    layer0_outputs(4405) <= not (a xor b);
    layer0_outputs(4406) <= b;
    layer0_outputs(4407) <= not (a and b);
    layer0_outputs(4408) <= not (a xor b);
    layer0_outputs(4409) <= not (a or b);
    layer0_outputs(4410) <= not (a or b);
    layer0_outputs(4411) <= a or b;
    layer0_outputs(4412) <= not (a and b);
    layer0_outputs(4413) <= a xor b;
    layer0_outputs(4414) <= not (a or b);
    layer0_outputs(4415) <= not (a or b);
    layer0_outputs(4416) <= b and not a;
    layer0_outputs(4417) <= not (a xor b);
    layer0_outputs(4418) <= b;
    layer0_outputs(4419) <= not b;
    layer0_outputs(4420) <= a and not b;
    layer0_outputs(4421) <= not (a xor b);
    layer0_outputs(4422) <= a and not b;
    layer0_outputs(4423) <= not a or b;
    layer0_outputs(4424) <= b;
    layer0_outputs(4425) <= b and not a;
    layer0_outputs(4426) <= not (a or b);
    layer0_outputs(4427) <= not (a or b);
    layer0_outputs(4428) <= not b;
    layer0_outputs(4429) <= not a;
    layer0_outputs(4430) <= a xor b;
    layer0_outputs(4431) <= a;
    layer0_outputs(4432) <= not (a xor b);
    layer0_outputs(4433) <= a xor b;
    layer0_outputs(4434) <= b;
    layer0_outputs(4435) <= not (a or b);
    layer0_outputs(4436) <= not (a or b);
    layer0_outputs(4437) <= a and not b;
    layer0_outputs(4438) <= a or b;
    layer0_outputs(4439) <= not a or b;
    layer0_outputs(4440) <= not (a or b);
    layer0_outputs(4441) <= not a or b;
    layer0_outputs(4442) <= b;
    layer0_outputs(4443) <= 1'b1;
    layer0_outputs(4444) <= a xor b;
    layer0_outputs(4445) <= not (a xor b);
    layer0_outputs(4446) <= a;
    layer0_outputs(4447) <= a xor b;
    layer0_outputs(4448) <= a xor b;
    layer0_outputs(4449) <= not (a or b);
    layer0_outputs(4450) <= a;
    layer0_outputs(4451) <= not (a or b);
    layer0_outputs(4452) <= a or b;
    layer0_outputs(4453) <= a or b;
    layer0_outputs(4454) <= a xor b;
    layer0_outputs(4455) <= not a;
    layer0_outputs(4456) <= b and not a;
    layer0_outputs(4457) <= not a;
    layer0_outputs(4458) <= 1'b0;
    layer0_outputs(4459) <= not (a xor b);
    layer0_outputs(4460) <= b and not a;
    layer0_outputs(4461) <= a or b;
    layer0_outputs(4462) <= a and b;
    layer0_outputs(4463) <= not b;
    layer0_outputs(4464) <= not b or a;
    layer0_outputs(4465) <= a and b;
    layer0_outputs(4466) <= not b or a;
    layer0_outputs(4467) <= 1'b1;
    layer0_outputs(4468) <= a and not b;
    layer0_outputs(4469) <= not b;
    layer0_outputs(4470) <= a or b;
    layer0_outputs(4471) <= a and not b;
    layer0_outputs(4472) <= not (a xor b);
    layer0_outputs(4473) <= not (a or b);
    layer0_outputs(4474) <= a or b;
    layer0_outputs(4475) <= a and not b;
    layer0_outputs(4476) <= not a;
    layer0_outputs(4477) <= not a or b;
    layer0_outputs(4478) <= not a;
    layer0_outputs(4479) <= not (a xor b);
    layer0_outputs(4480) <= a and not b;
    layer0_outputs(4481) <= a;
    layer0_outputs(4482) <= a or b;
    layer0_outputs(4483) <= b;
    layer0_outputs(4484) <= a;
    layer0_outputs(4485) <= not (a or b);
    layer0_outputs(4486) <= not (a and b);
    layer0_outputs(4487) <= b and not a;
    layer0_outputs(4488) <= b and not a;
    layer0_outputs(4489) <= not (a or b);
    layer0_outputs(4490) <= not (a xor b);
    layer0_outputs(4491) <= a;
    layer0_outputs(4492) <= not b;
    layer0_outputs(4493) <= not (a and b);
    layer0_outputs(4494) <= 1'b0;
    layer0_outputs(4495) <= not b;
    layer0_outputs(4496) <= not (a xor b);
    layer0_outputs(4497) <= b;
    layer0_outputs(4498) <= not (a xor b);
    layer0_outputs(4499) <= not b or a;
    layer0_outputs(4500) <= a xor b;
    layer0_outputs(4501) <= not a;
    layer0_outputs(4502) <= 1'b0;
    layer0_outputs(4503) <= not (a or b);
    layer0_outputs(4504) <= not (a xor b);
    layer0_outputs(4505) <= b;
    layer0_outputs(4506) <= not (a xor b);
    layer0_outputs(4507) <= a or b;
    layer0_outputs(4508) <= a and not b;
    layer0_outputs(4509) <= a or b;
    layer0_outputs(4510) <= not b;
    layer0_outputs(4511) <= a;
    layer0_outputs(4512) <= 1'b1;
    layer0_outputs(4513) <= not (a or b);
    layer0_outputs(4514) <= not a or b;
    layer0_outputs(4515) <= not (a or b);
    layer0_outputs(4516) <= b and not a;
    layer0_outputs(4517) <= a and not b;
    layer0_outputs(4518) <= not b;
    layer0_outputs(4519) <= not a or b;
    layer0_outputs(4520) <= not (a xor b);
    layer0_outputs(4521) <= a or b;
    layer0_outputs(4522) <= a xor b;
    layer0_outputs(4523) <= not a or b;
    layer0_outputs(4524) <= a;
    layer0_outputs(4525) <= not (a or b);
    layer0_outputs(4526) <= not (a or b);
    layer0_outputs(4527) <= a and b;
    layer0_outputs(4528) <= 1'b1;
    layer0_outputs(4529) <= not a;
    layer0_outputs(4530) <= not (a or b);
    layer0_outputs(4531) <= b;
    layer0_outputs(4532) <= not a;
    layer0_outputs(4533) <= a xor b;
    layer0_outputs(4534) <= not a or b;
    layer0_outputs(4535) <= not (a xor b);
    layer0_outputs(4536) <= a or b;
    layer0_outputs(4537) <= a;
    layer0_outputs(4538) <= not a;
    layer0_outputs(4539) <= not (a or b);
    layer0_outputs(4540) <= a or b;
    layer0_outputs(4541) <= not b or a;
    layer0_outputs(4542) <= b;
    layer0_outputs(4543) <= not b or a;
    layer0_outputs(4544) <= not a;
    layer0_outputs(4545) <= not a or b;
    layer0_outputs(4546) <= not (a or b);
    layer0_outputs(4547) <= not b;
    layer0_outputs(4548) <= a xor b;
    layer0_outputs(4549) <= not b or a;
    layer0_outputs(4550) <= a xor b;
    layer0_outputs(4551) <= b;
    layer0_outputs(4552) <= a or b;
    layer0_outputs(4553) <= not (a or b);
    layer0_outputs(4554) <= a or b;
    layer0_outputs(4555) <= not a or b;
    layer0_outputs(4556) <= b and not a;
    layer0_outputs(4557) <= a;
    layer0_outputs(4558) <= not a or b;
    layer0_outputs(4559) <= not (a xor b);
    layer0_outputs(4560) <= a and not b;
    layer0_outputs(4561) <= a;
    layer0_outputs(4562) <= not (a or b);
    layer0_outputs(4563) <= a xor b;
    layer0_outputs(4564) <= not b or a;
    layer0_outputs(4565) <= a xor b;
    layer0_outputs(4566) <= not (a or b);
    layer0_outputs(4567) <= a or b;
    layer0_outputs(4568) <= a or b;
    layer0_outputs(4569) <= not (a or b);
    layer0_outputs(4570) <= b and not a;
    layer0_outputs(4571) <= a and not b;
    layer0_outputs(4572) <= not b or a;
    layer0_outputs(4573) <= a or b;
    layer0_outputs(4574) <= b and not a;
    layer0_outputs(4575) <= a and b;
    layer0_outputs(4576) <= not (a xor b);
    layer0_outputs(4577) <= not (a and b);
    layer0_outputs(4578) <= not (a or b);
    layer0_outputs(4579) <= not b or a;
    layer0_outputs(4580) <= a xor b;
    layer0_outputs(4581) <= 1'b0;
    layer0_outputs(4582) <= 1'b1;
    layer0_outputs(4583) <= a or b;
    layer0_outputs(4584) <= b;
    layer0_outputs(4585) <= a;
    layer0_outputs(4586) <= a;
    layer0_outputs(4587) <= 1'b1;
    layer0_outputs(4588) <= a or b;
    layer0_outputs(4589) <= not (a or b);
    layer0_outputs(4590) <= a and not b;
    layer0_outputs(4591) <= a and b;
    layer0_outputs(4592) <= a and not b;
    layer0_outputs(4593) <= b and not a;
    layer0_outputs(4594) <= not (a and b);
    layer0_outputs(4595) <= not b or a;
    layer0_outputs(4596) <= not b or a;
    layer0_outputs(4597) <= not a or b;
    layer0_outputs(4598) <= not b;
    layer0_outputs(4599) <= not b;
    layer0_outputs(4600) <= not a;
    layer0_outputs(4601) <= a or b;
    layer0_outputs(4602) <= not a or b;
    layer0_outputs(4603) <= not b;
    layer0_outputs(4604) <= not (a or b);
    layer0_outputs(4605) <= a or b;
    layer0_outputs(4606) <= not (a or b);
    layer0_outputs(4607) <= not (a and b);
    layer0_outputs(4608) <= not b;
    layer0_outputs(4609) <= a or b;
    layer0_outputs(4610) <= not a or b;
    layer0_outputs(4611) <= 1'b0;
    layer0_outputs(4612) <= not a or b;
    layer0_outputs(4613) <= not b;
    layer0_outputs(4614) <= not b or a;
    layer0_outputs(4615) <= a;
    layer0_outputs(4616) <= a or b;
    layer0_outputs(4617) <= not b;
    layer0_outputs(4618) <= not (a xor b);
    layer0_outputs(4619) <= not b;
    layer0_outputs(4620) <= not b;
    layer0_outputs(4621) <= 1'b1;
    layer0_outputs(4622) <= not (a xor b);
    layer0_outputs(4623) <= not (a xor b);
    layer0_outputs(4624) <= not (a xor b);
    layer0_outputs(4625) <= b;
    layer0_outputs(4626) <= not (a xor b);
    layer0_outputs(4627) <= a xor b;
    layer0_outputs(4628) <= not b;
    layer0_outputs(4629) <= not b;
    layer0_outputs(4630) <= not (a and b);
    layer0_outputs(4631) <= not (a or b);
    layer0_outputs(4632) <= not a or b;
    layer0_outputs(4633) <= not (a or b);
    layer0_outputs(4634) <= not b;
    layer0_outputs(4635) <= a xor b;
    layer0_outputs(4636) <= not (a or b);
    layer0_outputs(4637) <= a and not b;
    layer0_outputs(4638) <= a and b;
    layer0_outputs(4639) <= not b;
    layer0_outputs(4640) <= a;
    layer0_outputs(4641) <= not a;
    layer0_outputs(4642) <= a xor b;
    layer0_outputs(4643) <= a xor b;
    layer0_outputs(4644) <= not (a and b);
    layer0_outputs(4645) <= not (a and b);
    layer0_outputs(4646) <= a xor b;
    layer0_outputs(4647) <= b;
    layer0_outputs(4648) <= not b or a;
    layer0_outputs(4649) <= a and not b;
    layer0_outputs(4650) <= 1'b0;
    layer0_outputs(4651) <= not (a or b);
    layer0_outputs(4652) <= a and not b;
    layer0_outputs(4653) <= b and not a;
    layer0_outputs(4654) <= not b or a;
    layer0_outputs(4655) <= 1'b0;
    layer0_outputs(4656) <= a or b;
    layer0_outputs(4657) <= a or b;
    layer0_outputs(4658) <= not (a xor b);
    layer0_outputs(4659) <= b;
    layer0_outputs(4660) <= a xor b;
    layer0_outputs(4661) <= not (a or b);
    layer0_outputs(4662) <= not (a or b);
    layer0_outputs(4663) <= not (a or b);
    layer0_outputs(4664) <= b and not a;
    layer0_outputs(4665) <= not (a or b);
    layer0_outputs(4666) <= a or b;
    layer0_outputs(4667) <= not a or b;
    layer0_outputs(4668) <= not (a xor b);
    layer0_outputs(4669) <= not (a and b);
    layer0_outputs(4670) <= a or b;
    layer0_outputs(4671) <= a xor b;
    layer0_outputs(4672) <= not b or a;
    layer0_outputs(4673) <= a xor b;
    layer0_outputs(4674) <= a;
    layer0_outputs(4675) <= 1'b0;
    layer0_outputs(4676) <= 1'b0;
    layer0_outputs(4677) <= not a or b;
    layer0_outputs(4678) <= not a or b;
    layer0_outputs(4679) <= a xor b;
    layer0_outputs(4680) <= not a;
    layer0_outputs(4681) <= a and not b;
    layer0_outputs(4682) <= b;
    layer0_outputs(4683) <= not a;
    layer0_outputs(4684) <= not b;
    layer0_outputs(4685) <= a and b;
    layer0_outputs(4686) <= a or b;
    layer0_outputs(4687) <= b and not a;
    layer0_outputs(4688) <= b;
    layer0_outputs(4689) <= not (a xor b);
    layer0_outputs(4690) <= b;
    layer0_outputs(4691) <= not b;
    layer0_outputs(4692) <= not (a or b);
    layer0_outputs(4693) <= not b;
    layer0_outputs(4694) <= not (a xor b);
    layer0_outputs(4695) <= a xor b;
    layer0_outputs(4696) <= a or b;
    layer0_outputs(4697) <= not (a or b);
    layer0_outputs(4698) <= a xor b;
    layer0_outputs(4699) <= b;
    layer0_outputs(4700) <= not b;
    layer0_outputs(4701) <= not (a xor b);
    layer0_outputs(4702) <= not b;
    layer0_outputs(4703) <= b;
    layer0_outputs(4704) <= not b;
    layer0_outputs(4705) <= not (a and b);
    layer0_outputs(4706) <= not (a or b);
    layer0_outputs(4707) <= a and not b;
    layer0_outputs(4708) <= a and not b;
    layer0_outputs(4709) <= a xor b;
    layer0_outputs(4710) <= a xor b;
    layer0_outputs(4711) <= not (a or b);
    layer0_outputs(4712) <= not (a and b);
    layer0_outputs(4713) <= not (a xor b);
    layer0_outputs(4714) <= not (a xor b);
    layer0_outputs(4715) <= not (a xor b);
    layer0_outputs(4716) <= not (a or b);
    layer0_outputs(4717) <= not b or a;
    layer0_outputs(4718) <= not b;
    layer0_outputs(4719) <= a or b;
    layer0_outputs(4720) <= not (a or b);
    layer0_outputs(4721) <= a and not b;
    layer0_outputs(4722) <= not a or b;
    layer0_outputs(4723) <= not (a or b);
    layer0_outputs(4724) <= a xor b;
    layer0_outputs(4725) <= not a;
    layer0_outputs(4726) <= 1'b1;
    layer0_outputs(4727) <= not (a xor b);
    layer0_outputs(4728) <= a or b;
    layer0_outputs(4729) <= not b;
    layer0_outputs(4730) <= 1'b0;
    layer0_outputs(4731) <= b and not a;
    layer0_outputs(4732) <= b;
    layer0_outputs(4733) <= not (a xor b);
    layer0_outputs(4734) <= b and not a;
    layer0_outputs(4735) <= not a;
    layer0_outputs(4736) <= a;
    layer0_outputs(4737) <= not b or a;
    layer0_outputs(4738) <= not a or b;
    layer0_outputs(4739) <= not a;
    layer0_outputs(4740) <= not b or a;
    layer0_outputs(4741) <= not (a xor b);
    layer0_outputs(4742) <= b;
    layer0_outputs(4743) <= not (a or b);
    layer0_outputs(4744) <= a or b;
    layer0_outputs(4745) <= a or b;
    layer0_outputs(4746) <= a;
    layer0_outputs(4747) <= not (a or b);
    layer0_outputs(4748) <= not (a xor b);
    layer0_outputs(4749) <= a and not b;
    layer0_outputs(4750) <= not b;
    layer0_outputs(4751) <= a and not b;
    layer0_outputs(4752) <= a or b;
    layer0_outputs(4753) <= not (a or b);
    layer0_outputs(4754) <= not a or b;
    layer0_outputs(4755) <= b;
    layer0_outputs(4756) <= not b;
    layer0_outputs(4757) <= not (a xor b);
    layer0_outputs(4758) <= a xor b;
    layer0_outputs(4759) <= a;
    layer0_outputs(4760) <= b and not a;
    layer0_outputs(4761) <= not b or a;
    layer0_outputs(4762) <= a or b;
    layer0_outputs(4763) <= b;
    layer0_outputs(4764) <= a and b;
    layer0_outputs(4765) <= not a;
    layer0_outputs(4766) <= a or b;
    layer0_outputs(4767) <= b;
    layer0_outputs(4768) <= not (a or b);
    layer0_outputs(4769) <= a or b;
    layer0_outputs(4770) <= not (a xor b);
    layer0_outputs(4771) <= not a;
    layer0_outputs(4772) <= not a or b;
    layer0_outputs(4773) <= a or b;
    layer0_outputs(4774) <= not b;
    layer0_outputs(4775) <= a;
    layer0_outputs(4776) <= not (a or b);
    layer0_outputs(4777) <= b and not a;
    layer0_outputs(4778) <= a and not b;
    layer0_outputs(4779) <= a;
    layer0_outputs(4780) <= a and not b;
    layer0_outputs(4781) <= not b;
    layer0_outputs(4782) <= a and not b;
    layer0_outputs(4783) <= 1'b1;
    layer0_outputs(4784) <= not (a xor b);
    layer0_outputs(4785) <= a or b;
    layer0_outputs(4786) <= a or b;
    layer0_outputs(4787) <= a or b;
    layer0_outputs(4788) <= a or b;
    layer0_outputs(4789) <= a and b;
    layer0_outputs(4790) <= b and not a;
    layer0_outputs(4791) <= a and not b;
    layer0_outputs(4792) <= b;
    layer0_outputs(4793) <= not a or b;
    layer0_outputs(4794) <= a xor b;
    layer0_outputs(4795) <= not a;
    layer0_outputs(4796) <= b and not a;
    layer0_outputs(4797) <= not (a or b);
    layer0_outputs(4798) <= not b;
    layer0_outputs(4799) <= a or b;
    layer0_outputs(4800) <= 1'b0;
    layer0_outputs(4801) <= a or b;
    layer0_outputs(4802) <= a xor b;
    layer0_outputs(4803) <= a xor b;
    layer0_outputs(4804) <= not a or b;
    layer0_outputs(4805) <= a or b;
    layer0_outputs(4806) <= not (a or b);
    layer0_outputs(4807) <= not b;
    layer0_outputs(4808) <= a xor b;
    layer0_outputs(4809) <= not b;
    layer0_outputs(4810) <= not b or a;
    layer0_outputs(4811) <= not a or b;
    layer0_outputs(4812) <= not (a or b);
    layer0_outputs(4813) <= not (a and b);
    layer0_outputs(4814) <= a or b;
    layer0_outputs(4815) <= b;
    layer0_outputs(4816) <= b and not a;
    layer0_outputs(4817) <= not (a xor b);
    layer0_outputs(4818) <= 1'b0;
    layer0_outputs(4819) <= not b or a;
    layer0_outputs(4820) <= not a;
    layer0_outputs(4821) <= b and not a;
    layer0_outputs(4822) <= not a;
    layer0_outputs(4823) <= not b or a;
    layer0_outputs(4824) <= a xor b;
    layer0_outputs(4825) <= not a;
    layer0_outputs(4826) <= a and not b;
    layer0_outputs(4827) <= not (a xor b);
    layer0_outputs(4828) <= not b;
    layer0_outputs(4829) <= a xor b;
    layer0_outputs(4830) <= 1'b1;
    layer0_outputs(4831) <= a and b;
    layer0_outputs(4832) <= not a or b;
    layer0_outputs(4833) <= a and not b;
    layer0_outputs(4834) <= b;
    layer0_outputs(4835) <= not (a or b);
    layer0_outputs(4836) <= not a;
    layer0_outputs(4837) <= a or b;
    layer0_outputs(4838) <= a xor b;
    layer0_outputs(4839) <= a or b;
    layer0_outputs(4840) <= not b;
    layer0_outputs(4841) <= a xor b;
    layer0_outputs(4842) <= not a;
    layer0_outputs(4843) <= a;
    layer0_outputs(4844) <= not b or a;
    layer0_outputs(4845) <= b;
    layer0_outputs(4846) <= a and b;
    layer0_outputs(4847) <= not (a or b);
    layer0_outputs(4848) <= b;
    layer0_outputs(4849) <= a;
    layer0_outputs(4850) <= not (a xor b);
    layer0_outputs(4851) <= 1'b0;
    layer0_outputs(4852) <= b;
    layer0_outputs(4853) <= b;
    layer0_outputs(4854) <= not (a and b);
    layer0_outputs(4855) <= not (a or b);
    layer0_outputs(4856) <= a xor b;
    layer0_outputs(4857) <= not (a or b);
    layer0_outputs(4858) <= not (a xor b);
    layer0_outputs(4859) <= not (a or b);
    layer0_outputs(4860) <= not a;
    layer0_outputs(4861) <= not (a xor b);
    layer0_outputs(4862) <= a or b;
    layer0_outputs(4863) <= not (a or b);
    layer0_outputs(4864) <= b and not a;
    layer0_outputs(4865) <= not b or a;
    layer0_outputs(4866) <= not a;
    layer0_outputs(4867) <= not (a xor b);
    layer0_outputs(4868) <= not b;
    layer0_outputs(4869) <= 1'b0;
    layer0_outputs(4870) <= not (a or b);
    layer0_outputs(4871) <= not (a or b);
    layer0_outputs(4872) <= not (a or b);
    layer0_outputs(4873) <= b;
    layer0_outputs(4874) <= not b or a;
    layer0_outputs(4875) <= not (a xor b);
    layer0_outputs(4876) <= a and b;
    layer0_outputs(4877) <= not b or a;
    layer0_outputs(4878) <= b;
    layer0_outputs(4879) <= a;
    layer0_outputs(4880) <= not a;
    layer0_outputs(4881) <= b;
    layer0_outputs(4882) <= a and b;
    layer0_outputs(4883) <= not a;
    layer0_outputs(4884) <= 1'b0;
    layer0_outputs(4885) <= not a;
    layer0_outputs(4886) <= a xor b;
    layer0_outputs(4887) <= not b;
    layer0_outputs(4888) <= not a;
    layer0_outputs(4889) <= a or b;
    layer0_outputs(4890) <= a or b;
    layer0_outputs(4891) <= a;
    layer0_outputs(4892) <= a and b;
    layer0_outputs(4893) <= not a;
    layer0_outputs(4894) <= a or b;
    layer0_outputs(4895) <= a;
    layer0_outputs(4896) <= not a;
    layer0_outputs(4897) <= a or b;
    layer0_outputs(4898) <= not b;
    layer0_outputs(4899) <= a xor b;
    layer0_outputs(4900) <= not a;
    layer0_outputs(4901) <= b;
    layer0_outputs(4902) <= a and not b;
    layer0_outputs(4903) <= b;
    layer0_outputs(4904) <= a and not b;
    layer0_outputs(4905) <= not a;
    layer0_outputs(4906) <= a xor b;
    layer0_outputs(4907) <= a or b;
    layer0_outputs(4908) <= not (a or b);
    layer0_outputs(4909) <= not a;
    layer0_outputs(4910) <= a;
    layer0_outputs(4911) <= 1'b1;
    layer0_outputs(4912) <= a and not b;
    layer0_outputs(4913) <= a or b;
    layer0_outputs(4914) <= not (a and b);
    layer0_outputs(4915) <= a;
    layer0_outputs(4916) <= not b or a;
    layer0_outputs(4917) <= 1'b1;
    layer0_outputs(4918) <= b and not a;
    layer0_outputs(4919) <= a xor b;
    layer0_outputs(4920) <= not (a or b);
    layer0_outputs(4921) <= not (a or b);
    layer0_outputs(4922) <= a xor b;
    layer0_outputs(4923) <= a xor b;
    layer0_outputs(4924) <= a or b;
    layer0_outputs(4925) <= b;
    layer0_outputs(4926) <= b and not a;
    layer0_outputs(4927) <= not b or a;
    layer0_outputs(4928) <= not a;
    layer0_outputs(4929) <= a or b;
    layer0_outputs(4930) <= not (a or b);
    layer0_outputs(4931) <= b and not a;
    layer0_outputs(4932) <= not b or a;
    layer0_outputs(4933) <= a;
    layer0_outputs(4934) <= not (a xor b);
    layer0_outputs(4935) <= not b;
    layer0_outputs(4936) <= not b;
    layer0_outputs(4937) <= not b or a;
    layer0_outputs(4938) <= not b or a;
    layer0_outputs(4939) <= a and not b;
    layer0_outputs(4940) <= not (a or b);
    layer0_outputs(4941) <= not (a xor b);
    layer0_outputs(4942) <= not a;
    layer0_outputs(4943) <= a;
    layer0_outputs(4944) <= not (a xor b);
    layer0_outputs(4945) <= not (a or b);
    layer0_outputs(4946) <= a or b;
    layer0_outputs(4947) <= not a or b;
    layer0_outputs(4948) <= not (a xor b);
    layer0_outputs(4949) <= a xor b;
    layer0_outputs(4950) <= a and not b;
    layer0_outputs(4951) <= 1'b1;
    layer0_outputs(4952) <= b and not a;
    layer0_outputs(4953) <= not a;
    layer0_outputs(4954) <= not (a xor b);
    layer0_outputs(4955) <= a or b;
    layer0_outputs(4956) <= a or b;
    layer0_outputs(4957) <= not a;
    layer0_outputs(4958) <= a and b;
    layer0_outputs(4959) <= a;
    layer0_outputs(4960) <= not b;
    layer0_outputs(4961) <= not (a xor b);
    layer0_outputs(4962) <= not (a or b);
    layer0_outputs(4963) <= a or b;
    layer0_outputs(4964) <= not (a or b);
    layer0_outputs(4965) <= a and not b;
    layer0_outputs(4966) <= a or b;
    layer0_outputs(4967) <= a and not b;
    layer0_outputs(4968) <= b and not a;
    layer0_outputs(4969) <= b;
    layer0_outputs(4970) <= b;
    layer0_outputs(4971) <= b and not a;
    layer0_outputs(4972) <= b;
    layer0_outputs(4973) <= not b or a;
    layer0_outputs(4974) <= a xor b;
    layer0_outputs(4975) <= a and b;
    layer0_outputs(4976) <= a or b;
    layer0_outputs(4977) <= not b or a;
    layer0_outputs(4978) <= not b;
    layer0_outputs(4979) <= b;
    layer0_outputs(4980) <= a and b;
    layer0_outputs(4981) <= 1'b1;
    layer0_outputs(4982) <= a xor b;
    layer0_outputs(4983) <= not a;
    layer0_outputs(4984) <= not b or a;
    layer0_outputs(4985) <= a;
    layer0_outputs(4986) <= not (a or b);
    layer0_outputs(4987) <= a xor b;
    layer0_outputs(4988) <= not (a or b);
    layer0_outputs(4989) <= not (a and b);
    layer0_outputs(4990) <= a and not b;
    layer0_outputs(4991) <= not (a xor b);
    layer0_outputs(4992) <= not a;
    layer0_outputs(4993) <= not b;
    layer0_outputs(4994) <= not a;
    layer0_outputs(4995) <= not (a or b);
    layer0_outputs(4996) <= not (a xor b);
    layer0_outputs(4997) <= not b;
    layer0_outputs(4998) <= 1'b1;
    layer0_outputs(4999) <= b and not a;
    layer0_outputs(5000) <= not (a or b);
    layer0_outputs(5001) <= not (a and b);
    layer0_outputs(5002) <= not a;
    layer0_outputs(5003) <= a or b;
    layer0_outputs(5004) <= 1'b0;
    layer0_outputs(5005) <= not (a xor b);
    layer0_outputs(5006) <= b and not a;
    layer0_outputs(5007) <= not a or b;
    layer0_outputs(5008) <= 1'b1;
    layer0_outputs(5009) <= not a;
    layer0_outputs(5010) <= 1'b0;
    layer0_outputs(5011) <= a;
    layer0_outputs(5012) <= b and not a;
    layer0_outputs(5013) <= not (a or b);
    layer0_outputs(5014) <= a or b;
    layer0_outputs(5015) <= not b or a;
    layer0_outputs(5016) <= not (a xor b);
    layer0_outputs(5017) <= not a or b;
    layer0_outputs(5018) <= a xor b;
    layer0_outputs(5019) <= a or b;
    layer0_outputs(5020) <= not a or b;
    layer0_outputs(5021) <= not a;
    layer0_outputs(5022) <= not a;
    layer0_outputs(5023) <= a or b;
    layer0_outputs(5024) <= not b or a;
    layer0_outputs(5025) <= not (a or b);
    layer0_outputs(5026) <= a or b;
    layer0_outputs(5027) <= not a;
    layer0_outputs(5028) <= b and not a;
    layer0_outputs(5029) <= not (a xor b);
    layer0_outputs(5030) <= not b or a;
    layer0_outputs(5031) <= 1'b0;
    layer0_outputs(5032) <= b;
    layer0_outputs(5033) <= not (a or b);
    layer0_outputs(5034) <= b and not a;
    layer0_outputs(5035) <= not (a or b);
    layer0_outputs(5036) <= not (a xor b);
    layer0_outputs(5037) <= not b;
    layer0_outputs(5038) <= not (a or b);
    layer0_outputs(5039) <= not (a xor b);
    layer0_outputs(5040) <= a or b;
    layer0_outputs(5041) <= a;
    layer0_outputs(5042) <= a;
    layer0_outputs(5043) <= not b or a;
    layer0_outputs(5044) <= b;
    layer0_outputs(5045) <= not (a or b);
    layer0_outputs(5046) <= b and not a;
    layer0_outputs(5047) <= not (a or b);
    layer0_outputs(5048) <= a and not b;
    layer0_outputs(5049) <= a;
    layer0_outputs(5050) <= a or b;
    layer0_outputs(5051) <= b;
    layer0_outputs(5052) <= a xor b;
    layer0_outputs(5053) <= not a;
    layer0_outputs(5054) <= a or b;
    layer0_outputs(5055) <= b and not a;
    layer0_outputs(5056) <= not (a or b);
    layer0_outputs(5057) <= not (a or b);
    layer0_outputs(5058) <= 1'b1;
    layer0_outputs(5059) <= a or b;
    layer0_outputs(5060) <= a;
    layer0_outputs(5061) <= a;
    layer0_outputs(5062) <= not b;
    layer0_outputs(5063) <= a or b;
    layer0_outputs(5064) <= not a or b;
    layer0_outputs(5065) <= not (a or b);
    layer0_outputs(5066) <= not b;
    layer0_outputs(5067) <= not (a xor b);
    layer0_outputs(5068) <= not (a xor b);
    layer0_outputs(5069) <= a;
    layer0_outputs(5070) <= not (a xor b);
    layer0_outputs(5071) <= not (a and b);
    layer0_outputs(5072) <= 1'b0;
    layer0_outputs(5073) <= a or b;
    layer0_outputs(5074) <= a or b;
    layer0_outputs(5075) <= not a or b;
    layer0_outputs(5076) <= not b or a;
    layer0_outputs(5077) <= a xor b;
    layer0_outputs(5078) <= not a or b;
    layer0_outputs(5079) <= a or b;
    layer0_outputs(5080) <= not a or b;
    layer0_outputs(5081) <= b and not a;
    layer0_outputs(5082) <= not (a and b);
    layer0_outputs(5083) <= not (a or b);
    layer0_outputs(5084) <= a or b;
    layer0_outputs(5085) <= 1'b0;
    layer0_outputs(5086) <= not (a or b);
    layer0_outputs(5087) <= b;
    layer0_outputs(5088) <= a or b;
    layer0_outputs(5089) <= a or b;
    layer0_outputs(5090) <= not (a xor b);
    layer0_outputs(5091) <= a and not b;
    layer0_outputs(5092) <= b;
    layer0_outputs(5093) <= b and not a;
    layer0_outputs(5094) <= not (a or b);
    layer0_outputs(5095) <= a and not b;
    layer0_outputs(5096) <= not (a xor b);
    layer0_outputs(5097) <= not (a or b);
    layer0_outputs(5098) <= b and not a;
    layer0_outputs(5099) <= a xor b;
    layer0_outputs(5100) <= b and not a;
    layer0_outputs(5101) <= b and not a;
    layer0_outputs(5102) <= a xor b;
    layer0_outputs(5103) <= not (a or b);
    layer0_outputs(5104) <= b and not a;
    layer0_outputs(5105) <= not (a or b);
    layer0_outputs(5106) <= not a;
    layer0_outputs(5107) <= b;
    layer0_outputs(5108) <= a or b;
    layer0_outputs(5109) <= a;
    layer0_outputs(5110) <= a xor b;
    layer0_outputs(5111) <= not a or b;
    layer0_outputs(5112) <= b;
    layer0_outputs(5113) <= not b;
    layer0_outputs(5114) <= b;
    layer0_outputs(5115) <= not b or a;
    layer0_outputs(5116) <= a;
    layer0_outputs(5117) <= a;
    layer0_outputs(5118) <= a xor b;
    layer0_outputs(5119) <= 1'b1;
    layer1_outputs(0) <= a xor b;
    layer1_outputs(1) <= a;
    layer1_outputs(2) <= not b;
    layer1_outputs(3) <= not b;
    layer1_outputs(4) <= a and not b;
    layer1_outputs(5) <= b;
    layer1_outputs(6) <= a;
    layer1_outputs(7) <= not a;
    layer1_outputs(8) <= not b;
    layer1_outputs(9) <= b;
    layer1_outputs(10) <= b;
    layer1_outputs(11) <= b;
    layer1_outputs(12) <= not (a or b);
    layer1_outputs(13) <= not b;
    layer1_outputs(14) <= not (a xor b);
    layer1_outputs(15) <= b;
    layer1_outputs(16) <= not (a xor b);
    layer1_outputs(17) <= b and not a;
    layer1_outputs(18) <= b;
    layer1_outputs(19) <= a;
    layer1_outputs(20) <= not b;
    layer1_outputs(21) <= not a;
    layer1_outputs(22) <= a and not b;
    layer1_outputs(23) <= not (a xor b);
    layer1_outputs(24) <= not a;
    layer1_outputs(25) <= a and not b;
    layer1_outputs(26) <= not a;
    layer1_outputs(27) <= not b or a;
    layer1_outputs(28) <= b;
    layer1_outputs(29) <= not (a and b);
    layer1_outputs(30) <= a;
    layer1_outputs(31) <= a or b;
    layer1_outputs(32) <= a or b;
    layer1_outputs(33) <= not a;
    layer1_outputs(34) <= a xor b;
    layer1_outputs(35) <= not a or b;
    layer1_outputs(36) <= a;
    layer1_outputs(37) <= a;
    layer1_outputs(38) <= not (a and b);
    layer1_outputs(39) <= not b or a;
    layer1_outputs(40) <= not (a and b);
    layer1_outputs(41) <= not (a or b);
    layer1_outputs(42) <= not a;
    layer1_outputs(43) <= not (a and b);
    layer1_outputs(44) <= a xor b;
    layer1_outputs(45) <= b and not a;
    layer1_outputs(46) <= not (a and b);
    layer1_outputs(47) <= not a;
    layer1_outputs(48) <= not b;
    layer1_outputs(49) <= b;
    layer1_outputs(50) <= not b or a;
    layer1_outputs(51) <= a or b;
    layer1_outputs(52) <= not a or b;
    layer1_outputs(53) <= not (a or b);
    layer1_outputs(54) <= not a;
    layer1_outputs(55) <= not b or a;
    layer1_outputs(56) <= not a or b;
    layer1_outputs(57) <= not a;
    layer1_outputs(58) <= 1'b0;
    layer1_outputs(59) <= not a;
    layer1_outputs(60) <= not (a xor b);
    layer1_outputs(61) <= not (a xor b);
    layer1_outputs(62) <= not b or a;
    layer1_outputs(63) <= not a;
    layer1_outputs(64) <= not (a xor b);
    layer1_outputs(65) <= not b or a;
    layer1_outputs(66) <= not (a or b);
    layer1_outputs(67) <= not a or b;
    layer1_outputs(68) <= not a or b;
    layer1_outputs(69) <= a;
    layer1_outputs(70) <= b;
    layer1_outputs(71) <= a or b;
    layer1_outputs(72) <= a xor b;
    layer1_outputs(73) <= a and not b;
    layer1_outputs(74) <= not a or b;
    layer1_outputs(75) <= not (a xor b);
    layer1_outputs(76) <= a xor b;
    layer1_outputs(77) <= not (a or b);
    layer1_outputs(78) <= not (a xor b);
    layer1_outputs(79) <= not (a xor b);
    layer1_outputs(80) <= not (a or b);
    layer1_outputs(81) <= not b or a;
    layer1_outputs(82) <= b and not a;
    layer1_outputs(83) <= not (a and b);
    layer1_outputs(84) <= a;
    layer1_outputs(85) <= not b;
    layer1_outputs(86) <= not b;
    layer1_outputs(87) <= a or b;
    layer1_outputs(88) <= b and not a;
    layer1_outputs(89) <= not b;
    layer1_outputs(90) <= not a or b;
    layer1_outputs(91) <= a and b;
    layer1_outputs(92) <= a or b;
    layer1_outputs(93) <= not a;
    layer1_outputs(94) <= not (a or b);
    layer1_outputs(95) <= a xor b;
    layer1_outputs(96) <= a or b;
    layer1_outputs(97) <= not a;
    layer1_outputs(98) <= not a or b;
    layer1_outputs(99) <= b;
    layer1_outputs(100) <= b;
    layer1_outputs(101) <= not (a or b);
    layer1_outputs(102) <= not b;
    layer1_outputs(103) <= not b;
    layer1_outputs(104) <= not (a and b);
    layer1_outputs(105) <= not a;
    layer1_outputs(106) <= a;
    layer1_outputs(107) <= a and not b;
    layer1_outputs(108) <= a;
    layer1_outputs(109) <= a and not b;
    layer1_outputs(110) <= b and not a;
    layer1_outputs(111) <= not b;
    layer1_outputs(112) <= not (a or b);
    layer1_outputs(113) <= b and not a;
    layer1_outputs(114) <= a and b;
    layer1_outputs(115) <= a and b;
    layer1_outputs(116) <= a and not b;
    layer1_outputs(117) <= not (a xor b);
    layer1_outputs(118) <= not (a xor b);
    layer1_outputs(119) <= not a;
    layer1_outputs(120) <= a xor b;
    layer1_outputs(121) <= not (a and b);
    layer1_outputs(122) <= not a;
    layer1_outputs(123) <= b and not a;
    layer1_outputs(124) <= not (a and b);
    layer1_outputs(125) <= a and not b;
    layer1_outputs(126) <= not (a and b);
    layer1_outputs(127) <= a;
    layer1_outputs(128) <= not a or b;
    layer1_outputs(129) <= not (a xor b);
    layer1_outputs(130) <= a and not b;
    layer1_outputs(131) <= a and b;
    layer1_outputs(132) <= not b or a;
    layer1_outputs(133) <= not b or a;
    layer1_outputs(134) <= b;
    layer1_outputs(135) <= not (a and b);
    layer1_outputs(136) <= 1'b1;
    layer1_outputs(137) <= not b or a;
    layer1_outputs(138) <= a and b;
    layer1_outputs(139) <= not b;
    layer1_outputs(140) <= not b or a;
    layer1_outputs(141) <= not b or a;
    layer1_outputs(142) <= a and not b;
    layer1_outputs(143) <= b;
    layer1_outputs(144) <= 1'b0;
    layer1_outputs(145) <= b;
    layer1_outputs(146) <= not b or a;
    layer1_outputs(147) <= not b or a;
    layer1_outputs(148) <= a and b;
    layer1_outputs(149) <= a;
    layer1_outputs(150) <= not b or a;
    layer1_outputs(151) <= not b;
    layer1_outputs(152) <= not a or b;
    layer1_outputs(153) <= 1'b1;
    layer1_outputs(154) <= 1'b1;
    layer1_outputs(155) <= not a;
    layer1_outputs(156) <= b and not a;
    layer1_outputs(157) <= not b;
    layer1_outputs(158) <= not (a xor b);
    layer1_outputs(159) <= not b;
    layer1_outputs(160) <= a;
    layer1_outputs(161) <= not b;
    layer1_outputs(162) <= not a;
    layer1_outputs(163) <= not a or b;
    layer1_outputs(164) <= not (a or b);
    layer1_outputs(165) <= a and b;
    layer1_outputs(166) <= b;
    layer1_outputs(167) <= a or b;
    layer1_outputs(168) <= not (a xor b);
    layer1_outputs(169) <= not b or a;
    layer1_outputs(170) <= 1'b0;
    layer1_outputs(171) <= not b;
    layer1_outputs(172) <= a or b;
    layer1_outputs(173) <= not b;
    layer1_outputs(174) <= not b;
    layer1_outputs(175) <= not a;
    layer1_outputs(176) <= 1'b1;
    layer1_outputs(177) <= b and not a;
    layer1_outputs(178) <= b;
    layer1_outputs(179) <= a;
    layer1_outputs(180) <= b;
    layer1_outputs(181) <= a;
    layer1_outputs(182) <= b;
    layer1_outputs(183) <= not (a xor b);
    layer1_outputs(184) <= a and not b;
    layer1_outputs(185) <= not b or a;
    layer1_outputs(186) <= not a or b;
    layer1_outputs(187) <= not b or a;
    layer1_outputs(188) <= a or b;
    layer1_outputs(189) <= not (a and b);
    layer1_outputs(190) <= b and not a;
    layer1_outputs(191) <= not a;
    layer1_outputs(192) <= b;
    layer1_outputs(193) <= a xor b;
    layer1_outputs(194) <= a and b;
    layer1_outputs(195) <= b;
    layer1_outputs(196) <= a and not b;
    layer1_outputs(197) <= not a;
    layer1_outputs(198) <= not a or b;
    layer1_outputs(199) <= not (a or b);
    layer1_outputs(200) <= not (a and b);
    layer1_outputs(201) <= b;
    layer1_outputs(202) <= a and b;
    layer1_outputs(203) <= 1'b0;
    layer1_outputs(204) <= not b;
    layer1_outputs(205) <= a xor b;
    layer1_outputs(206) <= a xor b;
    layer1_outputs(207) <= a and not b;
    layer1_outputs(208) <= a xor b;
    layer1_outputs(209) <= not a or b;
    layer1_outputs(210) <= not a;
    layer1_outputs(211) <= a;
    layer1_outputs(212) <= a;
    layer1_outputs(213) <= not b;
    layer1_outputs(214) <= a;
    layer1_outputs(215) <= a xor b;
    layer1_outputs(216) <= 1'b1;
    layer1_outputs(217) <= a;
    layer1_outputs(218) <= a;
    layer1_outputs(219) <= b and not a;
    layer1_outputs(220) <= not (a and b);
    layer1_outputs(221) <= not (a and b);
    layer1_outputs(222) <= not (a and b);
    layer1_outputs(223) <= not b;
    layer1_outputs(224) <= a;
    layer1_outputs(225) <= not b or a;
    layer1_outputs(226) <= not b or a;
    layer1_outputs(227) <= not b or a;
    layer1_outputs(228) <= not (a xor b);
    layer1_outputs(229) <= not b or a;
    layer1_outputs(230) <= not a or b;
    layer1_outputs(231) <= not b;
    layer1_outputs(232) <= b and not a;
    layer1_outputs(233) <= not b or a;
    layer1_outputs(234) <= b and not a;
    layer1_outputs(235) <= not a;
    layer1_outputs(236) <= b;
    layer1_outputs(237) <= b and not a;
    layer1_outputs(238) <= b and not a;
    layer1_outputs(239) <= a and b;
    layer1_outputs(240) <= b and not a;
    layer1_outputs(241) <= a or b;
    layer1_outputs(242) <= b and not a;
    layer1_outputs(243) <= not b;
    layer1_outputs(244) <= b;
    layer1_outputs(245) <= not (a and b);
    layer1_outputs(246) <= not a or b;
    layer1_outputs(247) <= a;
    layer1_outputs(248) <= b;
    layer1_outputs(249) <= a and b;
    layer1_outputs(250) <= a;
    layer1_outputs(251) <= a xor b;
    layer1_outputs(252) <= not a;
    layer1_outputs(253) <= not b;
    layer1_outputs(254) <= b;
    layer1_outputs(255) <= b and not a;
    layer1_outputs(256) <= a;
    layer1_outputs(257) <= b;
    layer1_outputs(258) <= a or b;
    layer1_outputs(259) <= a and b;
    layer1_outputs(260) <= not b or a;
    layer1_outputs(261) <= not a;
    layer1_outputs(262) <= not a or b;
    layer1_outputs(263) <= a xor b;
    layer1_outputs(264) <= not (a and b);
    layer1_outputs(265) <= a or b;
    layer1_outputs(266) <= not (a xor b);
    layer1_outputs(267) <= not (a and b);
    layer1_outputs(268) <= not b;
    layer1_outputs(269) <= not (a and b);
    layer1_outputs(270) <= not a;
    layer1_outputs(271) <= not b;
    layer1_outputs(272) <= b;
    layer1_outputs(273) <= not (a or b);
    layer1_outputs(274) <= a;
    layer1_outputs(275) <= 1'b0;
    layer1_outputs(276) <= b;
    layer1_outputs(277) <= a and b;
    layer1_outputs(278) <= not a;
    layer1_outputs(279) <= a;
    layer1_outputs(280) <= not b;
    layer1_outputs(281) <= not b or a;
    layer1_outputs(282) <= not (a xor b);
    layer1_outputs(283) <= a;
    layer1_outputs(284) <= b and not a;
    layer1_outputs(285) <= a and not b;
    layer1_outputs(286) <= not b;
    layer1_outputs(287) <= a;
    layer1_outputs(288) <= 1'b0;
    layer1_outputs(289) <= a and not b;
    layer1_outputs(290) <= not (a and b);
    layer1_outputs(291) <= not b;
    layer1_outputs(292) <= 1'b0;
    layer1_outputs(293) <= a and not b;
    layer1_outputs(294) <= b;
    layer1_outputs(295) <= b;
    layer1_outputs(296) <= not a or b;
    layer1_outputs(297) <= a or b;
    layer1_outputs(298) <= b and not a;
    layer1_outputs(299) <= a;
    layer1_outputs(300) <= a or b;
    layer1_outputs(301) <= not a or b;
    layer1_outputs(302) <= not a;
    layer1_outputs(303) <= 1'b0;
    layer1_outputs(304) <= a xor b;
    layer1_outputs(305) <= a or b;
    layer1_outputs(306) <= not (a xor b);
    layer1_outputs(307) <= b;
    layer1_outputs(308) <= a xor b;
    layer1_outputs(309) <= a and b;
    layer1_outputs(310) <= a;
    layer1_outputs(311) <= b;
    layer1_outputs(312) <= b and not a;
    layer1_outputs(313) <= not (a xor b);
    layer1_outputs(314) <= not (a xor b);
    layer1_outputs(315) <= not a;
    layer1_outputs(316) <= b and not a;
    layer1_outputs(317) <= not (a xor b);
    layer1_outputs(318) <= a and b;
    layer1_outputs(319) <= b;
    layer1_outputs(320) <= not (a and b);
    layer1_outputs(321) <= not b;
    layer1_outputs(322) <= not b or a;
    layer1_outputs(323) <= not a or b;
    layer1_outputs(324) <= not a;
    layer1_outputs(325) <= a and b;
    layer1_outputs(326) <= not b;
    layer1_outputs(327) <= 1'b0;
    layer1_outputs(328) <= a and not b;
    layer1_outputs(329) <= a and b;
    layer1_outputs(330) <= not (a and b);
    layer1_outputs(331) <= not b;
    layer1_outputs(332) <= a or b;
    layer1_outputs(333) <= not a;
    layer1_outputs(334) <= b and not a;
    layer1_outputs(335) <= not (a or b);
    layer1_outputs(336) <= a or b;
    layer1_outputs(337) <= not b;
    layer1_outputs(338) <= a;
    layer1_outputs(339) <= not (a xor b);
    layer1_outputs(340) <= not b or a;
    layer1_outputs(341) <= not (a and b);
    layer1_outputs(342) <= b and not a;
    layer1_outputs(343) <= a and b;
    layer1_outputs(344) <= not a or b;
    layer1_outputs(345) <= not (a or b);
    layer1_outputs(346) <= not (a and b);
    layer1_outputs(347) <= a;
    layer1_outputs(348) <= not (a and b);
    layer1_outputs(349) <= not (a xor b);
    layer1_outputs(350) <= a xor b;
    layer1_outputs(351) <= b;
    layer1_outputs(352) <= b and not a;
    layer1_outputs(353) <= a xor b;
    layer1_outputs(354) <= a xor b;
    layer1_outputs(355) <= b;
    layer1_outputs(356) <= a;
    layer1_outputs(357) <= not (a or b);
    layer1_outputs(358) <= not (a or b);
    layer1_outputs(359) <= not b or a;
    layer1_outputs(360) <= not b or a;
    layer1_outputs(361) <= not a or b;
    layer1_outputs(362) <= a;
    layer1_outputs(363) <= a and b;
    layer1_outputs(364) <= a or b;
    layer1_outputs(365) <= a or b;
    layer1_outputs(366) <= a and not b;
    layer1_outputs(367) <= a and not b;
    layer1_outputs(368) <= not (a xor b);
    layer1_outputs(369) <= a;
    layer1_outputs(370) <= b;
    layer1_outputs(371) <= a and not b;
    layer1_outputs(372) <= not a;
    layer1_outputs(373) <= a and b;
    layer1_outputs(374) <= a;
    layer1_outputs(375) <= not (a xor b);
    layer1_outputs(376) <= b and not a;
    layer1_outputs(377) <= a;
    layer1_outputs(378) <= not (a and b);
    layer1_outputs(379) <= a and not b;
    layer1_outputs(380) <= b and not a;
    layer1_outputs(381) <= b and not a;
    layer1_outputs(382) <= a xor b;
    layer1_outputs(383) <= not a or b;
    layer1_outputs(384) <= b;
    layer1_outputs(385) <= a;
    layer1_outputs(386) <= not (a xor b);
    layer1_outputs(387) <= not (a or b);
    layer1_outputs(388) <= not b;
    layer1_outputs(389) <= not a;
    layer1_outputs(390) <= a and b;
    layer1_outputs(391) <= not a;
    layer1_outputs(392) <= not (a and b);
    layer1_outputs(393) <= not b or a;
    layer1_outputs(394) <= not b;
    layer1_outputs(395) <= a;
    layer1_outputs(396) <= not (a and b);
    layer1_outputs(397) <= a;
    layer1_outputs(398) <= b;
    layer1_outputs(399) <= not (a xor b);
    layer1_outputs(400) <= a or b;
    layer1_outputs(401) <= a and b;
    layer1_outputs(402) <= not b or a;
    layer1_outputs(403) <= b and not a;
    layer1_outputs(404) <= a and not b;
    layer1_outputs(405) <= b and not a;
    layer1_outputs(406) <= not (a and b);
    layer1_outputs(407) <= a;
    layer1_outputs(408) <= not (a and b);
    layer1_outputs(409) <= a and not b;
    layer1_outputs(410) <= not (a and b);
    layer1_outputs(411) <= a xor b;
    layer1_outputs(412) <= a xor b;
    layer1_outputs(413) <= not a;
    layer1_outputs(414) <= b and not a;
    layer1_outputs(415) <= not a or b;
    layer1_outputs(416) <= a;
    layer1_outputs(417) <= b;
    layer1_outputs(418) <= a;
    layer1_outputs(419) <= b and not a;
    layer1_outputs(420) <= not (a xor b);
    layer1_outputs(421) <= not b;
    layer1_outputs(422) <= not (a or b);
    layer1_outputs(423) <= not b;
    layer1_outputs(424) <= a or b;
    layer1_outputs(425) <= a and not b;
    layer1_outputs(426) <= b and not a;
    layer1_outputs(427) <= not b or a;
    layer1_outputs(428) <= a;
    layer1_outputs(429) <= a;
    layer1_outputs(430) <= a xor b;
    layer1_outputs(431) <= not a;
    layer1_outputs(432) <= b;
    layer1_outputs(433) <= not (a xor b);
    layer1_outputs(434) <= a and not b;
    layer1_outputs(435) <= not b or a;
    layer1_outputs(436) <= a and b;
    layer1_outputs(437) <= not (a and b);
    layer1_outputs(438) <= a;
    layer1_outputs(439) <= not b;
    layer1_outputs(440) <= not b;
    layer1_outputs(441) <= not (a and b);
    layer1_outputs(442) <= a or b;
    layer1_outputs(443) <= a or b;
    layer1_outputs(444) <= a;
    layer1_outputs(445) <= 1'b1;
    layer1_outputs(446) <= b and not a;
    layer1_outputs(447) <= a and b;
    layer1_outputs(448) <= not b;
    layer1_outputs(449) <= not a or b;
    layer1_outputs(450) <= not b or a;
    layer1_outputs(451) <= not (a xor b);
    layer1_outputs(452) <= a or b;
    layer1_outputs(453) <= a or b;
    layer1_outputs(454) <= not (a xor b);
    layer1_outputs(455) <= not (a and b);
    layer1_outputs(456) <= b;
    layer1_outputs(457) <= b and not a;
    layer1_outputs(458) <= b and not a;
    layer1_outputs(459) <= b and not a;
    layer1_outputs(460) <= b and not a;
    layer1_outputs(461) <= not (a or b);
    layer1_outputs(462) <= not a or b;
    layer1_outputs(463) <= not (a or b);
    layer1_outputs(464) <= not (a or b);
    layer1_outputs(465) <= not a;
    layer1_outputs(466) <= not (a and b);
    layer1_outputs(467) <= a or b;
    layer1_outputs(468) <= not (a and b);
    layer1_outputs(469) <= a and b;
    layer1_outputs(470) <= not (a and b);
    layer1_outputs(471) <= not a or b;
    layer1_outputs(472) <= a and b;
    layer1_outputs(473) <= 1'b1;
    layer1_outputs(474) <= not (a and b);
    layer1_outputs(475) <= a xor b;
    layer1_outputs(476) <= not (a xor b);
    layer1_outputs(477) <= a;
    layer1_outputs(478) <= not (a xor b);
    layer1_outputs(479) <= a and b;
    layer1_outputs(480) <= not (a and b);
    layer1_outputs(481) <= not a or b;
    layer1_outputs(482) <= b;
    layer1_outputs(483) <= not a or b;
    layer1_outputs(484) <= not b or a;
    layer1_outputs(485) <= not (a or b);
    layer1_outputs(486) <= not b or a;
    layer1_outputs(487) <= not a or b;
    layer1_outputs(488) <= 1'b1;
    layer1_outputs(489) <= a xor b;
    layer1_outputs(490) <= not (a and b);
    layer1_outputs(491) <= not a;
    layer1_outputs(492) <= b;
    layer1_outputs(493) <= not a;
    layer1_outputs(494) <= a and not b;
    layer1_outputs(495) <= not b;
    layer1_outputs(496) <= a and b;
    layer1_outputs(497) <= not a;
    layer1_outputs(498) <= a or b;
    layer1_outputs(499) <= not (a xor b);
    layer1_outputs(500) <= a and not b;
    layer1_outputs(501) <= not a;
    layer1_outputs(502) <= b;
    layer1_outputs(503) <= not b;
    layer1_outputs(504) <= not a or b;
    layer1_outputs(505) <= b and not a;
    layer1_outputs(506) <= a and not b;
    layer1_outputs(507) <= b;
    layer1_outputs(508) <= a;
    layer1_outputs(509) <= a and b;
    layer1_outputs(510) <= not b or a;
    layer1_outputs(511) <= not (a and b);
    layer1_outputs(512) <= a xor b;
    layer1_outputs(513) <= a or b;
    layer1_outputs(514) <= not (a xor b);
    layer1_outputs(515) <= not a or b;
    layer1_outputs(516) <= not b or a;
    layer1_outputs(517) <= not a;
    layer1_outputs(518) <= b;
    layer1_outputs(519) <= not b;
    layer1_outputs(520) <= not (a or b);
    layer1_outputs(521) <= a and not b;
    layer1_outputs(522) <= a and b;
    layer1_outputs(523) <= b;
    layer1_outputs(524) <= a and b;
    layer1_outputs(525) <= not a;
    layer1_outputs(526) <= a xor b;
    layer1_outputs(527) <= not (a and b);
    layer1_outputs(528) <= not (a and b);
    layer1_outputs(529) <= not b or a;
    layer1_outputs(530) <= not a;
    layer1_outputs(531) <= b and not a;
    layer1_outputs(532) <= not b;
    layer1_outputs(533) <= b and not a;
    layer1_outputs(534) <= not (a or b);
    layer1_outputs(535) <= a xor b;
    layer1_outputs(536) <= not b;
    layer1_outputs(537) <= not b;
    layer1_outputs(538) <= a;
    layer1_outputs(539) <= not (a or b);
    layer1_outputs(540) <= a xor b;
    layer1_outputs(541) <= not b;
    layer1_outputs(542) <= a and not b;
    layer1_outputs(543) <= not a or b;
    layer1_outputs(544) <= b;
    layer1_outputs(545) <= not (a or b);
    layer1_outputs(546) <= a;
    layer1_outputs(547) <= 1'b0;
    layer1_outputs(548) <= not b;
    layer1_outputs(549) <= a and b;
    layer1_outputs(550) <= not b;
    layer1_outputs(551) <= a and b;
    layer1_outputs(552) <= a and not b;
    layer1_outputs(553) <= not b;
    layer1_outputs(554) <= 1'b0;
    layer1_outputs(555) <= b and not a;
    layer1_outputs(556) <= not (a xor b);
    layer1_outputs(557) <= a xor b;
    layer1_outputs(558) <= a or b;
    layer1_outputs(559) <= a xor b;
    layer1_outputs(560) <= not (a xor b);
    layer1_outputs(561) <= not a;
    layer1_outputs(562) <= not b;
    layer1_outputs(563) <= not a or b;
    layer1_outputs(564) <= a xor b;
    layer1_outputs(565) <= a xor b;
    layer1_outputs(566) <= not b or a;
    layer1_outputs(567) <= not a;
    layer1_outputs(568) <= not a or b;
    layer1_outputs(569) <= a and not b;
    layer1_outputs(570) <= not a;
    layer1_outputs(571) <= 1'b1;
    layer1_outputs(572) <= a and b;
    layer1_outputs(573) <= not (a xor b);
    layer1_outputs(574) <= not b;
    layer1_outputs(575) <= not a;
    layer1_outputs(576) <= a;
    layer1_outputs(577) <= 1'b1;
    layer1_outputs(578) <= a and b;
    layer1_outputs(579) <= not a;
    layer1_outputs(580) <= a;
    layer1_outputs(581) <= a and b;
    layer1_outputs(582) <= a or b;
    layer1_outputs(583) <= b and not a;
    layer1_outputs(584) <= not (a or b);
    layer1_outputs(585) <= not (a xor b);
    layer1_outputs(586) <= not b;
    layer1_outputs(587) <= 1'b0;
    layer1_outputs(588) <= b and not a;
    layer1_outputs(589) <= not a or b;
    layer1_outputs(590) <= not b;
    layer1_outputs(591) <= not (a xor b);
    layer1_outputs(592) <= 1'b1;
    layer1_outputs(593) <= a and not b;
    layer1_outputs(594) <= b and not a;
    layer1_outputs(595) <= a xor b;
    layer1_outputs(596) <= not (a and b);
    layer1_outputs(597) <= not (a and b);
    layer1_outputs(598) <= not (a or b);
    layer1_outputs(599) <= not b;
    layer1_outputs(600) <= b and not a;
    layer1_outputs(601) <= a or b;
    layer1_outputs(602) <= not b;
    layer1_outputs(603) <= a and b;
    layer1_outputs(604) <= 1'b0;
    layer1_outputs(605) <= not a or b;
    layer1_outputs(606) <= not a;
    layer1_outputs(607) <= a;
    layer1_outputs(608) <= a and not b;
    layer1_outputs(609) <= a;
    layer1_outputs(610) <= not (a or b);
    layer1_outputs(611) <= b;
    layer1_outputs(612) <= not (a or b);
    layer1_outputs(613) <= not (a xor b);
    layer1_outputs(614) <= not (a or b);
    layer1_outputs(615) <= a xor b;
    layer1_outputs(616) <= a;
    layer1_outputs(617) <= a or b;
    layer1_outputs(618) <= not b or a;
    layer1_outputs(619) <= b;
    layer1_outputs(620) <= not a;
    layer1_outputs(621) <= a and b;
    layer1_outputs(622) <= a and not b;
    layer1_outputs(623) <= 1'b1;
    layer1_outputs(624) <= not b or a;
    layer1_outputs(625) <= a and b;
    layer1_outputs(626) <= not b;
    layer1_outputs(627) <= not (a xor b);
    layer1_outputs(628) <= a;
    layer1_outputs(629) <= not a or b;
    layer1_outputs(630) <= not (a and b);
    layer1_outputs(631) <= a and not b;
    layer1_outputs(632) <= not b or a;
    layer1_outputs(633) <= not b;
    layer1_outputs(634) <= not (a and b);
    layer1_outputs(635) <= b;
    layer1_outputs(636) <= not (a and b);
    layer1_outputs(637) <= a and not b;
    layer1_outputs(638) <= not b or a;
    layer1_outputs(639) <= a or b;
    layer1_outputs(640) <= not a;
    layer1_outputs(641) <= a;
    layer1_outputs(642) <= a and not b;
    layer1_outputs(643) <= a xor b;
    layer1_outputs(644) <= not (a or b);
    layer1_outputs(645) <= a and not b;
    layer1_outputs(646) <= not (a or b);
    layer1_outputs(647) <= 1'b0;
    layer1_outputs(648) <= a and b;
    layer1_outputs(649) <= not a;
    layer1_outputs(650) <= b and not a;
    layer1_outputs(651) <= not (a and b);
    layer1_outputs(652) <= not (a or b);
    layer1_outputs(653) <= a or b;
    layer1_outputs(654) <= a or b;
    layer1_outputs(655) <= a and b;
    layer1_outputs(656) <= not a;
    layer1_outputs(657) <= a xor b;
    layer1_outputs(658) <= not b or a;
    layer1_outputs(659) <= a;
    layer1_outputs(660) <= a and not b;
    layer1_outputs(661) <= a xor b;
    layer1_outputs(662) <= b;
    layer1_outputs(663) <= not (a xor b);
    layer1_outputs(664) <= not b;
    layer1_outputs(665) <= a and b;
    layer1_outputs(666) <= a xor b;
    layer1_outputs(667) <= b;
    layer1_outputs(668) <= a and not b;
    layer1_outputs(669) <= a and b;
    layer1_outputs(670) <= a and not b;
    layer1_outputs(671) <= not b or a;
    layer1_outputs(672) <= not b or a;
    layer1_outputs(673) <= not b;
    layer1_outputs(674) <= not (a and b);
    layer1_outputs(675) <= not (a and b);
    layer1_outputs(676) <= not a;
    layer1_outputs(677) <= a;
    layer1_outputs(678) <= not (a or b);
    layer1_outputs(679) <= a or b;
    layer1_outputs(680) <= not (a or b);
    layer1_outputs(681) <= a;
    layer1_outputs(682) <= not b or a;
    layer1_outputs(683) <= b and not a;
    layer1_outputs(684) <= a and b;
    layer1_outputs(685) <= not (a or b);
    layer1_outputs(686) <= not (a and b);
    layer1_outputs(687) <= not (a xor b);
    layer1_outputs(688) <= not (a or b);
    layer1_outputs(689) <= a xor b;
    layer1_outputs(690) <= a or b;
    layer1_outputs(691) <= a and not b;
    layer1_outputs(692) <= not (a xor b);
    layer1_outputs(693) <= not (a and b);
    layer1_outputs(694) <= b;
    layer1_outputs(695) <= b and not a;
    layer1_outputs(696) <= b;
    layer1_outputs(697) <= a;
    layer1_outputs(698) <= a or b;
    layer1_outputs(699) <= b;
    layer1_outputs(700) <= a and b;
    layer1_outputs(701) <= a xor b;
    layer1_outputs(702) <= not b or a;
    layer1_outputs(703) <= not (a or b);
    layer1_outputs(704) <= a xor b;
    layer1_outputs(705) <= b and not a;
    layer1_outputs(706) <= a xor b;
    layer1_outputs(707) <= not b or a;
    layer1_outputs(708) <= not a or b;
    layer1_outputs(709) <= b;
    layer1_outputs(710) <= not a or b;
    layer1_outputs(711) <= a;
    layer1_outputs(712) <= b;
    layer1_outputs(713) <= 1'b1;
    layer1_outputs(714) <= a;
    layer1_outputs(715) <= not a;
    layer1_outputs(716) <= not a;
    layer1_outputs(717) <= not b;
    layer1_outputs(718) <= not (a xor b);
    layer1_outputs(719) <= a xor b;
    layer1_outputs(720) <= not b;
    layer1_outputs(721) <= not b;
    layer1_outputs(722) <= not b;
    layer1_outputs(723) <= not a;
    layer1_outputs(724) <= not (a or b);
    layer1_outputs(725) <= not a;
    layer1_outputs(726) <= b and not a;
    layer1_outputs(727) <= not (a and b);
    layer1_outputs(728) <= not b or a;
    layer1_outputs(729) <= a and not b;
    layer1_outputs(730) <= a xor b;
    layer1_outputs(731) <= not (a xor b);
    layer1_outputs(732) <= a and not b;
    layer1_outputs(733) <= not a or b;
    layer1_outputs(734) <= a and b;
    layer1_outputs(735) <= b and not a;
    layer1_outputs(736) <= a or b;
    layer1_outputs(737) <= not (a and b);
    layer1_outputs(738) <= not a or b;
    layer1_outputs(739) <= not a or b;
    layer1_outputs(740) <= a;
    layer1_outputs(741) <= a;
    layer1_outputs(742) <= b;
    layer1_outputs(743) <= not b or a;
    layer1_outputs(744) <= a and b;
    layer1_outputs(745) <= not (a and b);
    layer1_outputs(746) <= not b;
    layer1_outputs(747) <= not b;
    layer1_outputs(748) <= 1'b0;
    layer1_outputs(749) <= a and not b;
    layer1_outputs(750) <= a;
    layer1_outputs(751) <= not (a or b);
    layer1_outputs(752) <= b and not a;
    layer1_outputs(753) <= not b;
    layer1_outputs(754) <= a or b;
    layer1_outputs(755) <= not b;
    layer1_outputs(756) <= b and not a;
    layer1_outputs(757) <= not b;
    layer1_outputs(758) <= not b;
    layer1_outputs(759) <= not b;
    layer1_outputs(760) <= a xor b;
    layer1_outputs(761) <= not (a or b);
    layer1_outputs(762) <= a or b;
    layer1_outputs(763) <= b;
    layer1_outputs(764) <= a or b;
    layer1_outputs(765) <= a and not b;
    layer1_outputs(766) <= a and b;
    layer1_outputs(767) <= not (a xor b);
    layer1_outputs(768) <= 1'b0;
    layer1_outputs(769) <= not a or b;
    layer1_outputs(770) <= b;
    layer1_outputs(771) <= a;
    layer1_outputs(772) <= a and not b;
    layer1_outputs(773) <= not (a xor b);
    layer1_outputs(774) <= not (a xor b);
    layer1_outputs(775) <= not a or b;
    layer1_outputs(776) <= b;
    layer1_outputs(777) <= a and not b;
    layer1_outputs(778) <= a;
    layer1_outputs(779) <= a xor b;
    layer1_outputs(780) <= not (a or b);
    layer1_outputs(781) <= b;
    layer1_outputs(782) <= a and not b;
    layer1_outputs(783) <= a or b;
    layer1_outputs(784) <= 1'b0;
    layer1_outputs(785) <= not (a or b);
    layer1_outputs(786) <= not b or a;
    layer1_outputs(787) <= not b;
    layer1_outputs(788) <= a or b;
    layer1_outputs(789) <= a and b;
    layer1_outputs(790) <= not a;
    layer1_outputs(791) <= not (a or b);
    layer1_outputs(792) <= not (a or b);
    layer1_outputs(793) <= not (a or b);
    layer1_outputs(794) <= a and b;
    layer1_outputs(795) <= not (a xor b);
    layer1_outputs(796) <= b;
    layer1_outputs(797) <= a xor b;
    layer1_outputs(798) <= not b;
    layer1_outputs(799) <= a;
    layer1_outputs(800) <= not b;
    layer1_outputs(801) <= a;
    layer1_outputs(802) <= not b;
    layer1_outputs(803) <= b;
    layer1_outputs(804) <= not b or a;
    layer1_outputs(805) <= a and b;
    layer1_outputs(806) <= not b or a;
    layer1_outputs(807) <= a and not b;
    layer1_outputs(808) <= a xor b;
    layer1_outputs(809) <= b and not a;
    layer1_outputs(810) <= a and b;
    layer1_outputs(811) <= a;
    layer1_outputs(812) <= not (a or b);
    layer1_outputs(813) <= a or b;
    layer1_outputs(814) <= not a;
    layer1_outputs(815) <= not (a xor b);
    layer1_outputs(816) <= not b;
    layer1_outputs(817) <= not b or a;
    layer1_outputs(818) <= not b;
    layer1_outputs(819) <= not (a and b);
    layer1_outputs(820) <= not (a or b);
    layer1_outputs(821) <= 1'b0;
    layer1_outputs(822) <= b;
    layer1_outputs(823) <= a and not b;
    layer1_outputs(824) <= a and b;
    layer1_outputs(825) <= 1'b0;
    layer1_outputs(826) <= b;
    layer1_outputs(827) <= not (a xor b);
    layer1_outputs(828) <= a;
    layer1_outputs(829) <= a or b;
    layer1_outputs(830) <= not b or a;
    layer1_outputs(831) <= not b;
    layer1_outputs(832) <= not b or a;
    layer1_outputs(833) <= not a;
    layer1_outputs(834) <= a and b;
    layer1_outputs(835) <= not (a or b);
    layer1_outputs(836) <= a and not b;
    layer1_outputs(837) <= a;
    layer1_outputs(838) <= a;
    layer1_outputs(839) <= a and b;
    layer1_outputs(840) <= not a;
    layer1_outputs(841) <= b and not a;
    layer1_outputs(842) <= not a or b;
    layer1_outputs(843) <= a;
    layer1_outputs(844) <= b;
    layer1_outputs(845) <= not a;
    layer1_outputs(846) <= b;
    layer1_outputs(847) <= not (a and b);
    layer1_outputs(848) <= a and not b;
    layer1_outputs(849) <= not a or b;
    layer1_outputs(850) <= not (a xor b);
    layer1_outputs(851) <= a and not b;
    layer1_outputs(852) <= not b or a;
    layer1_outputs(853) <= a and b;
    layer1_outputs(854) <= not (a xor b);
    layer1_outputs(855) <= a and not b;
    layer1_outputs(856) <= b and not a;
    layer1_outputs(857) <= not (a or b);
    layer1_outputs(858) <= not (a xor b);
    layer1_outputs(859) <= a;
    layer1_outputs(860) <= not b or a;
    layer1_outputs(861) <= not a;
    layer1_outputs(862) <= b and not a;
    layer1_outputs(863) <= a and b;
    layer1_outputs(864) <= a;
    layer1_outputs(865) <= b and not a;
    layer1_outputs(866) <= not a or b;
    layer1_outputs(867) <= a;
    layer1_outputs(868) <= 1'b0;
    layer1_outputs(869) <= a;
    layer1_outputs(870) <= a;
    layer1_outputs(871) <= not a;
    layer1_outputs(872) <= a;
    layer1_outputs(873) <= b;
    layer1_outputs(874) <= b;
    layer1_outputs(875) <= a xor b;
    layer1_outputs(876) <= not b or a;
    layer1_outputs(877) <= a;
    layer1_outputs(878) <= not b or a;
    layer1_outputs(879) <= not a;
    layer1_outputs(880) <= a or b;
    layer1_outputs(881) <= b;
    layer1_outputs(882) <= not a or b;
    layer1_outputs(883) <= not (a xor b);
    layer1_outputs(884) <= b and not a;
    layer1_outputs(885) <= not b or a;
    layer1_outputs(886) <= a;
    layer1_outputs(887) <= not b;
    layer1_outputs(888) <= not a or b;
    layer1_outputs(889) <= a xor b;
    layer1_outputs(890) <= not b;
    layer1_outputs(891) <= not (a xor b);
    layer1_outputs(892) <= a and not b;
    layer1_outputs(893) <= not (a or b);
    layer1_outputs(894) <= a;
    layer1_outputs(895) <= b;
    layer1_outputs(896) <= a or b;
    layer1_outputs(897) <= a and not b;
    layer1_outputs(898) <= not (a or b);
    layer1_outputs(899) <= not (a and b);
    layer1_outputs(900) <= not b;
    layer1_outputs(901) <= not a;
    layer1_outputs(902) <= not a or b;
    layer1_outputs(903) <= a and b;
    layer1_outputs(904) <= a and b;
    layer1_outputs(905) <= a;
    layer1_outputs(906) <= not b or a;
    layer1_outputs(907) <= a;
    layer1_outputs(908) <= a and not b;
    layer1_outputs(909) <= a and not b;
    layer1_outputs(910) <= a and b;
    layer1_outputs(911) <= not a;
    layer1_outputs(912) <= a and not b;
    layer1_outputs(913) <= a and not b;
    layer1_outputs(914) <= a and b;
    layer1_outputs(915) <= a and not b;
    layer1_outputs(916) <= not b;
    layer1_outputs(917) <= not (a and b);
    layer1_outputs(918) <= not (a or b);
    layer1_outputs(919) <= a;
    layer1_outputs(920) <= 1'b0;
    layer1_outputs(921) <= b and not a;
    layer1_outputs(922) <= not (a or b);
    layer1_outputs(923) <= not b or a;
    layer1_outputs(924) <= a;
    layer1_outputs(925) <= not b;
    layer1_outputs(926) <= not a or b;
    layer1_outputs(927) <= a and b;
    layer1_outputs(928) <= not (a or b);
    layer1_outputs(929) <= a;
    layer1_outputs(930) <= a xor b;
    layer1_outputs(931) <= a or b;
    layer1_outputs(932) <= a and b;
    layer1_outputs(933) <= b;
    layer1_outputs(934) <= not a or b;
    layer1_outputs(935) <= a or b;
    layer1_outputs(936) <= not a or b;
    layer1_outputs(937) <= a and b;
    layer1_outputs(938) <= not a or b;
    layer1_outputs(939) <= not (a and b);
    layer1_outputs(940) <= not (a xor b);
    layer1_outputs(941) <= not b or a;
    layer1_outputs(942) <= not a;
    layer1_outputs(943) <= not b or a;
    layer1_outputs(944) <= b and not a;
    layer1_outputs(945) <= 1'b1;
    layer1_outputs(946) <= b and not a;
    layer1_outputs(947) <= not b;
    layer1_outputs(948) <= a and b;
    layer1_outputs(949) <= a xor b;
    layer1_outputs(950) <= not a or b;
    layer1_outputs(951) <= not a;
    layer1_outputs(952) <= not a or b;
    layer1_outputs(953) <= not (a and b);
    layer1_outputs(954) <= not (a or b);
    layer1_outputs(955) <= b and not a;
    layer1_outputs(956) <= not a;
    layer1_outputs(957) <= b and not a;
    layer1_outputs(958) <= not (a and b);
    layer1_outputs(959) <= a;
    layer1_outputs(960) <= 1'b0;
    layer1_outputs(961) <= not (a xor b);
    layer1_outputs(962) <= not a;
    layer1_outputs(963) <= b;
    layer1_outputs(964) <= not a or b;
    layer1_outputs(965) <= a;
    layer1_outputs(966) <= not a;
    layer1_outputs(967) <= not b or a;
    layer1_outputs(968) <= not (a and b);
    layer1_outputs(969) <= not (a xor b);
    layer1_outputs(970) <= not b;
    layer1_outputs(971) <= a;
    layer1_outputs(972) <= not (a xor b);
    layer1_outputs(973) <= a or b;
    layer1_outputs(974) <= not b;
    layer1_outputs(975) <= a;
    layer1_outputs(976) <= b;
    layer1_outputs(977) <= not b;
    layer1_outputs(978) <= a xor b;
    layer1_outputs(979) <= not a or b;
    layer1_outputs(980) <= a xor b;
    layer1_outputs(981) <= not b;
    layer1_outputs(982) <= a;
    layer1_outputs(983) <= not (a and b);
    layer1_outputs(984) <= a;
    layer1_outputs(985) <= not (a xor b);
    layer1_outputs(986) <= a and not b;
    layer1_outputs(987) <= b and not a;
    layer1_outputs(988) <= a and not b;
    layer1_outputs(989) <= not b;
    layer1_outputs(990) <= b and not a;
    layer1_outputs(991) <= not (a or b);
    layer1_outputs(992) <= 1'b1;
    layer1_outputs(993) <= a xor b;
    layer1_outputs(994) <= b and not a;
    layer1_outputs(995) <= not a;
    layer1_outputs(996) <= a and not b;
    layer1_outputs(997) <= not a;
    layer1_outputs(998) <= not (a xor b);
    layer1_outputs(999) <= b;
    layer1_outputs(1000) <= a;
    layer1_outputs(1001) <= a and not b;
    layer1_outputs(1002) <= not (a and b);
    layer1_outputs(1003) <= not a;
    layer1_outputs(1004) <= not a or b;
    layer1_outputs(1005) <= not a or b;
    layer1_outputs(1006) <= not a or b;
    layer1_outputs(1007) <= b and not a;
    layer1_outputs(1008) <= a and not b;
    layer1_outputs(1009) <= not a or b;
    layer1_outputs(1010) <= not b or a;
    layer1_outputs(1011) <= a and not b;
    layer1_outputs(1012) <= b;
    layer1_outputs(1013) <= a;
    layer1_outputs(1014) <= a or b;
    layer1_outputs(1015) <= b and not a;
    layer1_outputs(1016) <= a or b;
    layer1_outputs(1017) <= not b or a;
    layer1_outputs(1018) <= a and b;
    layer1_outputs(1019) <= a and b;
    layer1_outputs(1020) <= a and not b;
    layer1_outputs(1021) <= a;
    layer1_outputs(1022) <= not b or a;
    layer1_outputs(1023) <= b;
    layer1_outputs(1024) <= not b or a;
    layer1_outputs(1025) <= not b;
    layer1_outputs(1026) <= not (a xor b);
    layer1_outputs(1027) <= not a;
    layer1_outputs(1028) <= a or b;
    layer1_outputs(1029) <= a and not b;
    layer1_outputs(1030) <= a;
    layer1_outputs(1031) <= a;
    layer1_outputs(1032) <= a and b;
    layer1_outputs(1033) <= not (a or b);
    layer1_outputs(1034) <= not b or a;
    layer1_outputs(1035) <= not (a or b);
    layer1_outputs(1036) <= not (a and b);
    layer1_outputs(1037) <= b and not a;
    layer1_outputs(1038) <= not b or a;
    layer1_outputs(1039) <= not (a or b);
    layer1_outputs(1040) <= a or b;
    layer1_outputs(1041) <= not (a and b);
    layer1_outputs(1042) <= not b;
    layer1_outputs(1043) <= not (a xor b);
    layer1_outputs(1044) <= b;
    layer1_outputs(1045) <= not b or a;
    layer1_outputs(1046) <= not (a or b);
    layer1_outputs(1047) <= b;
    layer1_outputs(1048) <= not a;
    layer1_outputs(1049) <= b;
    layer1_outputs(1050) <= not b or a;
    layer1_outputs(1051) <= a and b;
    layer1_outputs(1052) <= 1'b1;
    layer1_outputs(1053) <= b;
    layer1_outputs(1054) <= a;
    layer1_outputs(1055) <= not b;
    layer1_outputs(1056) <= not a or b;
    layer1_outputs(1057) <= b;
    layer1_outputs(1058) <= a and not b;
    layer1_outputs(1059) <= a;
    layer1_outputs(1060) <= not a;
    layer1_outputs(1061) <= a and not b;
    layer1_outputs(1062) <= b;
    layer1_outputs(1063) <= a;
    layer1_outputs(1064) <= not a or b;
    layer1_outputs(1065) <= not a or b;
    layer1_outputs(1066) <= not b;
    layer1_outputs(1067) <= not a;
    layer1_outputs(1068) <= not b;
    layer1_outputs(1069) <= not (a or b);
    layer1_outputs(1070) <= not a or b;
    layer1_outputs(1071) <= a;
    layer1_outputs(1072) <= a or b;
    layer1_outputs(1073) <= a and b;
    layer1_outputs(1074) <= not (a xor b);
    layer1_outputs(1075) <= not a;
    layer1_outputs(1076) <= a xor b;
    layer1_outputs(1077) <= a xor b;
    layer1_outputs(1078) <= b and not a;
    layer1_outputs(1079) <= a;
    layer1_outputs(1080) <= not a or b;
    layer1_outputs(1081) <= not b or a;
    layer1_outputs(1082) <= not b;
    layer1_outputs(1083) <= 1'b1;
    layer1_outputs(1084) <= not (a xor b);
    layer1_outputs(1085) <= not a or b;
    layer1_outputs(1086) <= a and b;
    layer1_outputs(1087) <= not (a or b);
    layer1_outputs(1088) <= not a or b;
    layer1_outputs(1089) <= b;
    layer1_outputs(1090) <= not (a or b);
    layer1_outputs(1091) <= not b or a;
    layer1_outputs(1092) <= not b or a;
    layer1_outputs(1093) <= a and b;
    layer1_outputs(1094) <= not b or a;
    layer1_outputs(1095) <= not a or b;
    layer1_outputs(1096) <= a and b;
    layer1_outputs(1097) <= not a or b;
    layer1_outputs(1098) <= a and b;
    layer1_outputs(1099) <= not a;
    layer1_outputs(1100) <= not (a and b);
    layer1_outputs(1101) <= not b or a;
    layer1_outputs(1102) <= not a or b;
    layer1_outputs(1103) <= not a or b;
    layer1_outputs(1104) <= not b or a;
    layer1_outputs(1105) <= a and not b;
    layer1_outputs(1106) <= not b;
    layer1_outputs(1107) <= b and not a;
    layer1_outputs(1108) <= b;
    layer1_outputs(1109) <= a or b;
    layer1_outputs(1110) <= 1'b1;
    layer1_outputs(1111) <= not a or b;
    layer1_outputs(1112) <= a xor b;
    layer1_outputs(1113) <= a and b;
    layer1_outputs(1114) <= a or b;
    layer1_outputs(1115) <= a;
    layer1_outputs(1116) <= not b or a;
    layer1_outputs(1117) <= not (a or b);
    layer1_outputs(1118) <= not (a xor b);
    layer1_outputs(1119) <= not (a and b);
    layer1_outputs(1120) <= not (a xor b);
    layer1_outputs(1121) <= not a;
    layer1_outputs(1122) <= a and not b;
    layer1_outputs(1123) <= a;
    layer1_outputs(1124) <= a and b;
    layer1_outputs(1125) <= a;
    layer1_outputs(1126) <= not a or b;
    layer1_outputs(1127) <= not (a xor b);
    layer1_outputs(1128) <= not (a and b);
    layer1_outputs(1129) <= 1'b0;
    layer1_outputs(1130) <= not b or a;
    layer1_outputs(1131) <= b;
    layer1_outputs(1132) <= not a;
    layer1_outputs(1133) <= a and not b;
    layer1_outputs(1134) <= a and b;
    layer1_outputs(1135) <= not a;
    layer1_outputs(1136) <= not a;
    layer1_outputs(1137) <= not a;
    layer1_outputs(1138) <= 1'b1;
    layer1_outputs(1139) <= not b or a;
    layer1_outputs(1140) <= a;
    layer1_outputs(1141) <= b;
    layer1_outputs(1142) <= a;
    layer1_outputs(1143) <= not a;
    layer1_outputs(1144) <= not (a or b);
    layer1_outputs(1145) <= a and b;
    layer1_outputs(1146) <= not (a xor b);
    layer1_outputs(1147) <= a xor b;
    layer1_outputs(1148) <= not a or b;
    layer1_outputs(1149) <= not a or b;
    layer1_outputs(1150) <= not (a and b);
    layer1_outputs(1151) <= a;
    layer1_outputs(1152) <= not (a xor b);
    layer1_outputs(1153) <= not (a or b);
    layer1_outputs(1154) <= not (a and b);
    layer1_outputs(1155) <= not a or b;
    layer1_outputs(1156) <= not (a and b);
    layer1_outputs(1157) <= a or b;
    layer1_outputs(1158) <= a;
    layer1_outputs(1159) <= a and not b;
    layer1_outputs(1160) <= not (a xor b);
    layer1_outputs(1161) <= a and not b;
    layer1_outputs(1162) <= not b;
    layer1_outputs(1163) <= not b;
    layer1_outputs(1164) <= b and not a;
    layer1_outputs(1165) <= a and b;
    layer1_outputs(1166) <= b and not a;
    layer1_outputs(1167) <= not b or a;
    layer1_outputs(1168) <= not b;
    layer1_outputs(1169) <= b;
    layer1_outputs(1170) <= a and not b;
    layer1_outputs(1171) <= b and not a;
    layer1_outputs(1172) <= a and b;
    layer1_outputs(1173) <= not (a and b);
    layer1_outputs(1174) <= not b or a;
    layer1_outputs(1175) <= not a;
    layer1_outputs(1176) <= b;
    layer1_outputs(1177) <= not b or a;
    layer1_outputs(1178) <= b and not a;
    layer1_outputs(1179) <= not a or b;
    layer1_outputs(1180) <= a and not b;
    layer1_outputs(1181) <= not (a xor b);
    layer1_outputs(1182) <= a or b;
    layer1_outputs(1183) <= not a;
    layer1_outputs(1184) <= not (a and b);
    layer1_outputs(1185) <= not a;
    layer1_outputs(1186) <= not a;
    layer1_outputs(1187) <= a and not b;
    layer1_outputs(1188) <= a xor b;
    layer1_outputs(1189) <= a or b;
    layer1_outputs(1190) <= not a or b;
    layer1_outputs(1191) <= not a or b;
    layer1_outputs(1192) <= a and b;
    layer1_outputs(1193) <= a xor b;
    layer1_outputs(1194) <= not a;
    layer1_outputs(1195) <= a or b;
    layer1_outputs(1196) <= b;
    layer1_outputs(1197) <= not (a xor b);
    layer1_outputs(1198) <= not (a or b);
    layer1_outputs(1199) <= b;
    layer1_outputs(1200) <= not b;
    layer1_outputs(1201) <= not a;
    layer1_outputs(1202) <= a;
    layer1_outputs(1203) <= not b;
    layer1_outputs(1204) <= not (a xor b);
    layer1_outputs(1205) <= a or b;
    layer1_outputs(1206) <= not a or b;
    layer1_outputs(1207) <= not b;
    layer1_outputs(1208) <= not (a or b);
    layer1_outputs(1209) <= a and not b;
    layer1_outputs(1210) <= not (a xor b);
    layer1_outputs(1211) <= not a;
    layer1_outputs(1212) <= a;
    layer1_outputs(1213) <= not b;
    layer1_outputs(1214) <= a xor b;
    layer1_outputs(1215) <= a and b;
    layer1_outputs(1216) <= b;
    layer1_outputs(1217) <= not a or b;
    layer1_outputs(1218) <= b;
    layer1_outputs(1219) <= b;
    layer1_outputs(1220) <= b and not a;
    layer1_outputs(1221) <= a and b;
    layer1_outputs(1222) <= not b;
    layer1_outputs(1223) <= not a;
    layer1_outputs(1224) <= a and b;
    layer1_outputs(1225) <= a and b;
    layer1_outputs(1226) <= not b or a;
    layer1_outputs(1227) <= b and not a;
    layer1_outputs(1228) <= not (a xor b);
    layer1_outputs(1229) <= a and not b;
    layer1_outputs(1230) <= not b or a;
    layer1_outputs(1231) <= b and not a;
    layer1_outputs(1232) <= b and not a;
    layer1_outputs(1233) <= not a or b;
    layer1_outputs(1234) <= not b or a;
    layer1_outputs(1235) <= not b or a;
    layer1_outputs(1236) <= not (a xor b);
    layer1_outputs(1237) <= not a;
    layer1_outputs(1238) <= not a;
    layer1_outputs(1239) <= a and b;
    layer1_outputs(1240) <= not (a or b);
    layer1_outputs(1241) <= not (a and b);
    layer1_outputs(1242) <= not a;
    layer1_outputs(1243) <= a or b;
    layer1_outputs(1244) <= a xor b;
    layer1_outputs(1245) <= not b or a;
    layer1_outputs(1246) <= not b or a;
    layer1_outputs(1247) <= a or b;
    layer1_outputs(1248) <= a;
    layer1_outputs(1249) <= not a;
    layer1_outputs(1250) <= not b or a;
    layer1_outputs(1251) <= b and not a;
    layer1_outputs(1252) <= a xor b;
    layer1_outputs(1253) <= a and b;
    layer1_outputs(1254) <= a and b;
    layer1_outputs(1255) <= a or b;
    layer1_outputs(1256) <= not b or a;
    layer1_outputs(1257) <= not b or a;
    layer1_outputs(1258) <= a and not b;
    layer1_outputs(1259) <= a or b;
    layer1_outputs(1260) <= 1'b1;
    layer1_outputs(1261) <= not a;
    layer1_outputs(1262) <= a;
    layer1_outputs(1263) <= a and b;
    layer1_outputs(1264) <= not (a and b);
    layer1_outputs(1265) <= not b;
    layer1_outputs(1266) <= not b;
    layer1_outputs(1267) <= b;
    layer1_outputs(1268) <= not b;
    layer1_outputs(1269) <= not b;
    layer1_outputs(1270) <= a and b;
    layer1_outputs(1271) <= not b;
    layer1_outputs(1272) <= not a;
    layer1_outputs(1273) <= 1'b1;
    layer1_outputs(1274) <= not b;
    layer1_outputs(1275) <= not (a xor b);
    layer1_outputs(1276) <= a and b;
    layer1_outputs(1277) <= not (a xor b);
    layer1_outputs(1278) <= a;
    layer1_outputs(1279) <= 1'b1;
    layer1_outputs(1280) <= a;
    layer1_outputs(1281) <= a;
    layer1_outputs(1282) <= a or b;
    layer1_outputs(1283) <= 1'b1;
    layer1_outputs(1284) <= a xor b;
    layer1_outputs(1285) <= a or b;
    layer1_outputs(1286) <= not (a xor b);
    layer1_outputs(1287) <= a or b;
    layer1_outputs(1288) <= not (a xor b);
    layer1_outputs(1289) <= a xor b;
    layer1_outputs(1290) <= b;
    layer1_outputs(1291) <= not a;
    layer1_outputs(1292) <= not a or b;
    layer1_outputs(1293) <= 1'b0;
    layer1_outputs(1294) <= not b;
    layer1_outputs(1295) <= not b;
    layer1_outputs(1296) <= b and not a;
    layer1_outputs(1297) <= not a;
    layer1_outputs(1298) <= a;
    layer1_outputs(1299) <= a;
    layer1_outputs(1300) <= not b;
    layer1_outputs(1301) <= b and not a;
    layer1_outputs(1302) <= a;
    layer1_outputs(1303) <= not a;
    layer1_outputs(1304) <= b;
    layer1_outputs(1305) <= not a;
    layer1_outputs(1306) <= not a;
    layer1_outputs(1307) <= not b or a;
    layer1_outputs(1308) <= b;
    layer1_outputs(1309) <= not (a or b);
    layer1_outputs(1310) <= not (a xor b);
    layer1_outputs(1311) <= not (a xor b);
    layer1_outputs(1312) <= a and b;
    layer1_outputs(1313) <= not (a or b);
    layer1_outputs(1314) <= a;
    layer1_outputs(1315) <= not a or b;
    layer1_outputs(1316) <= a;
    layer1_outputs(1317) <= not b or a;
    layer1_outputs(1318) <= not b or a;
    layer1_outputs(1319) <= a or b;
    layer1_outputs(1320) <= a and b;
    layer1_outputs(1321) <= a and not b;
    layer1_outputs(1322) <= not b;
    layer1_outputs(1323) <= not b or a;
    layer1_outputs(1324) <= not b or a;
    layer1_outputs(1325) <= not (a or b);
    layer1_outputs(1326) <= not (a xor b);
    layer1_outputs(1327) <= a or b;
    layer1_outputs(1328) <= a or b;
    layer1_outputs(1329) <= not (a or b);
    layer1_outputs(1330) <= not a;
    layer1_outputs(1331) <= a xor b;
    layer1_outputs(1332) <= not b;
    layer1_outputs(1333) <= b;
    layer1_outputs(1334) <= a or b;
    layer1_outputs(1335) <= b;
    layer1_outputs(1336) <= a or b;
    layer1_outputs(1337) <= b;
    layer1_outputs(1338) <= a and b;
    layer1_outputs(1339) <= not a or b;
    layer1_outputs(1340) <= b and not a;
    layer1_outputs(1341) <= a;
    layer1_outputs(1342) <= not a;
    layer1_outputs(1343) <= not a or b;
    layer1_outputs(1344) <= not b;
    layer1_outputs(1345) <= not a;
    layer1_outputs(1346) <= a;
    layer1_outputs(1347) <= a;
    layer1_outputs(1348) <= not b;
    layer1_outputs(1349) <= not (a and b);
    layer1_outputs(1350) <= b and not a;
    layer1_outputs(1351) <= 1'b0;
    layer1_outputs(1352) <= a or b;
    layer1_outputs(1353) <= not b;
    layer1_outputs(1354) <= not b;
    layer1_outputs(1355) <= b and not a;
    layer1_outputs(1356) <= a and not b;
    layer1_outputs(1357) <= not b;
    layer1_outputs(1358) <= a and b;
    layer1_outputs(1359) <= not (a or b);
    layer1_outputs(1360) <= b;
    layer1_outputs(1361) <= a;
    layer1_outputs(1362) <= not b;
    layer1_outputs(1363) <= not b;
    layer1_outputs(1364) <= not b or a;
    layer1_outputs(1365) <= b and not a;
    layer1_outputs(1366) <= a and b;
    layer1_outputs(1367) <= a;
    layer1_outputs(1368) <= a and not b;
    layer1_outputs(1369) <= a and b;
    layer1_outputs(1370) <= not b or a;
    layer1_outputs(1371) <= not b or a;
    layer1_outputs(1372) <= not (a xor b);
    layer1_outputs(1373) <= not b or a;
    layer1_outputs(1374) <= not b;
    layer1_outputs(1375) <= b and not a;
    layer1_outputs(1376) <= a xor b;
    layer1_outputs(1377) <= a;
    layer1_outputs(1378) <= a;
    layer1_outputs(1379) <= a and b;
    layer1_outputs(1380) <= b;
    layer1_outputs(1381) <= not (a and b);
    layer1_outputs(1382) <= a;
    layer1_outputs(1383) <= not b or a;
    layer1_outputs(1384) <= b;
    layer1_outputs(1385) <= a xor b;
    layer1_outputs(1386) <= not b or a;
    layer1_outputs(1387) <= not b or a;
    layer1_outputs(1388) <= not b or a;
    layer1_outputs(1389) <= not (a and b);
    layer1_outputs(1390) <= a;
    layer1_outputs(1391) <= a and not b;
    layer1_outputs(1392) <= not (a or b);
    layer1_outputs(1393) <= a;
    layer1_outputs(1394) <= a and b;
    layer1_outputs(1395) <= not (a xor b);
    layer1_outputs(1396) <= not (a or b);
    layer1_outputs(1397) <= not a;
    layer1_outputs(1398) <= not (a xor b);
    layer1_outputs(1399) <= a and b;
    layer1_outputs(1400) <= not b;
    layer1_outputs(1401) <= not b;
    layer1_outputs(1402) <= a and not b;
    layer1_outputs(1403) <= not a or b;
    layer1_outputs(1404) <= not (a xor b);
    layer1_outputs(1405) <= not a;
    layer1_outputs(1406) <= b and not a;
    layer1_outputs(1407) <= a xor b;
    layer1_outputs(1408) <= a and not b;
    layer1_outputs(1409) <= b;
    layer1_outputs(1410) <= a;
    layer1_outputs(1411) <= a or b;
    layer1_outputs(1412) <= not b or a;
    layer1_outputs(1413) <= not b;
    layer1_outputs(1414) <= not b or a;
    layer1_outputs(1415) <= not b;
    layer1_outputs(1416) <= a;
    layer1_outputs(1417) <= not a;
    layer1_outputs(1418) <= b and not a;
    layer1_outputs(1419) <= b;
    layer1_outputs(1420) <= a and b;
    layer1_outputs(1421) <= a;
    layer1_outputs(1422) <= not b or a;
    layer1_outputs(1423) <= a xor b;
    layer1_outputs(1424) <= not (a xor b);
    layer1_outputs(1425) <= not (a and b);
    layer1_outputs(1426) <= a and not b;
    layer1_outputs(1427) <= a;
    layer1_outputs(1428) <= a;
    layer1_outputs(1429) <= not a or b;
    layer1_outputs(1430) <= not a;
    layer1_outputs(1431) <= not (a xor b);
    layer1_outputs(1432) <= b and not a;
    layer1_outputs(1433) <= b and not a;
    layer1_outputs(1434) <= not (a xor b);
    layer1_outputs(1435) <= b and not a;
    layer1_outputs(1436) <= b and not a;
    layer1_outputs(1437) <= a and b;
    layer1_outputs(1438) <= a;
    layer1_outputs(1439) <= a;
    layer1_outputs(1440) <= not (a or b);
    layer1_outputs(1441) <= b;
    layer1_outputs(1442) <= a;
    layer1_outputs(1443) <= not a;
    layer1_outputs(1444) <= not a;
    layer1_outputs(1445) <= not b;
    layer1_outputs(1446) <= a or b;
    layer1_outputs(1447) <= a and not b;
    layer1_outputs(1448) <= a or b;
    layer1_outputs(1449) <= a xor b;
    layer1_outputs(1450) <= not b;
    layer1_outputs(1451) <= not a;
    layer1_outputs(1452) <= a and not b;
    layer1_outputs(1453) <= not b or a;
    layer1_outputs(1454) <= not a;
    layer1_outputs(1455) <= not a or b;
    layer1_outputs(1456) <= a or b;
    layer1_outputs(1457) <= not (a and b);
    layer1_outputs(1458) <= b;
    layer1_outputs(1459) <= a or b;
    layer1_outputs(1460) <= a and b;
    layer1_outputs(1461) <= a and b;
    layer1_outputs(1462) <= a and b;
    layer1_outputs(1463) <= 1'b1;
    layer1_outputs(1464) <= b;
    layer1_outputs(1465) <= not b;
    layer1_outputs(1466) <= b and not a;
    layer1_outputs(1467) <= not (a and b);
    layer1_outputs(1468) <= b;
    layer1_outputs(1469) <= not (a xor b);
    layer1_outputs(1470) <= a xor b;
    layer1_outputs(1471) <= not a or b;
    layer1_outputs(1472) <= not b or a;
    layer1_outputs(1473) <= not a or b;
    layer1_outputs(1474) <= not a or b;
    layer1_outputs(1475) <= a and b;
    layer1_outputs(1476) <= b;
    layer1_outputs(1477) <= b and not a;
    layer1_outputs(1478) <= a;
    layer1_outputs(1479) <= b and not a;
    layer1_outputs(1480) <= a;
    layer1_outputs(1481) <= not b;
    layer1_outputs(1482) <= a or b;
    layer1_outputs(1483) <= b and not a;
    layer1_outputs(1484) <= a;
    layer1_outputs(1485) <= not (a and b);
    layer1_outputs(1486) <= not b or a;
    layer1_outputs(1487) <= 1'b0;
    layer1_outputs(1488) <= b;
    layer1_outputs(1489) <= a;
    layer1_outputs(1490) <= not b;
    layer1_outputs(1491) <= not b or a;
    layer1_outputs(1492) <= b;
    layer1_outputs(1493) <= not b;
    layer1_outputs(1494) <= not (a and b);
    layer1_outputs(1495) <= a xor b;
    layer1_outputs(1496) <= 1'b1;
    layer1_outputs(1497) <= a or b;
    layer1_outputs(1498) <= not a;
    layer1_outputs(1499) <= a and b;
    layer1_outputs(1500) <= a or b;
    layer1_outputs(1501) <= not a;
    layer1_outputs(1502) <= a and b;
    layer1_outputs(1503) <= not (a and b);
    layer1_outputs(1504) <= b;
    layer1_outputs(1505) <= a;
    layer1_outputs(1506) <= a;
    layer1_outputs(1507) <= not b;
    layer1_outputs(1508) <= a and not b;
    layer1_outputs(1509) <= not b or a;
    layer1_outputs(1510) <= not a or b;
    layer1_outputs(1511) <= b;
    layer1_outputs(1512) <= b;
    layer1_outputs(1513) <= not b;
    layer1_outputs(1514) <= a and not b;
    layer1_outputs(1515) <= a xor b;
    layer1_outputs(1516) <= b and not a;
    layer1_outputs(1517) <= a and b;
    layer1_outputs(1518) <= a and b;
    layer1_outputs(1519) <= not b or a;
    layer1_outputs(1520) <= not (a or b);
    layer1_outputs(1521) <= not b;
    layer1_outputs(1522) <= a and b;
    layer1_outputs(1523) <= not b or a;
    layer1_outputs(1524) <= a xor b;
    layer1_outputs(1525) <= a;
    layer1_outputs(1526) <= b and not a;
    layer1_outputs(1527) <= a;
    layer1_outputs(1528) <= a and not b;
    layer1_outputs(1529) <= a;
    layer1_outputs(1530) <= not (a xor b);
    layer1_outputs(1531) <= not a;
    layer1_outputs(1532) <= a or b;
    layer1_outputs(1533) <= a or b;
    layer1_outputs(1534) <= not a;
    layer1_outputs(1535) <= b and not a;
    layer1_outputs(1536) <= not a;
    layer1_outputs(1537) <= not (a or b);
    layer1_outputs(1538) <= b;
    layer1_outputs(1539) <= a xor b;
    layer1_outputs(1540) <= a;
    layer1_outputs(1541) <= not a;
    layer1_outputs(1542) <= not b or a;
    layer1_outputs(1543) <= b;
    layer1_outputs(1544) <= not b or a;
    layer1_outputs(1545) <= b;
    layer1_outputs(1546) <= a or b;
    layer1_outputs(1547) <= not b;
    layer1_outputs(1548) <= a xor b;
    layer1_outputs(1549) <= not a or b;
    layer1_outputs(1550) <= not (a xor b);
    layer1_outputs(1551) <= not (a and b);
    layer1_outputs(1552) <= not (a or b);
    layer1_outputs(1553) <= a and b;
    layer1_outputs(1554) <= a;
    layer1_outputs(1555) <= not b;
    layer1_outputs(1556) <= a;
    layer1_outputs(1557) <= a and b;
    layer1_outputs(1558) <= not b;
    layer1_outputs(1559) <= a xor b;
    layer1_outputs(1560) <= a and not b;
    layer1_outputs(1561) <= a and not b;
    layer1_outputs(1562) <= b;
    layer1_outputs(1563) <= b and not a;
    layer1_outputs(1564) <= a xor b;
    layer1_outputs(1565) <= not b or a;
    layer1_outputs(1566) <= a or b;
    layer1_outputs(1567) <= 1'b0;
    layer1_outputs(1568) <= a xor b;
    layer1_outputs(1569) <= b;
    layer1_outputs(1570) <= b;
    layer1_outputs(1571) <= not (a xor b);
    layer1_outputs(1572) <= a;
    layer1_outputs(1573) <= 1'b1;
    layer1_outputs(1574) <= not b;
    layer1_outputs(1575) <= 1'b1;
    layer1_outputs(1576) <= a;
    layer1_outputs(1577) <= b;
    layer1_outputs(1578) <= not b;
    layer1_outputs(1579) <= b;
    layer1_outputs(1580) <= not (a xor b);
    layer1_outputs(1581) <= b and not a;
    layer1_outputs(1582) <= a and not b;
    layer1_outputs(1583) <= a and b;
    layer1_outputs(1584) <= a or b;
    layer1_outputs(1585) <= not b or a;
    layer1_outputs(1586) <= not (a and b);
    layer1_outputs(1587) <= b and not a;
    layer1_outputs(1588) <= not (a and b);
    layer1_outputs(1589) <= b;
    layer1_outputs(1590) <= a;
    layer1_outputs(1591) <= a;
    layer1_outputs(1592) <= not (a xor b);
    layer1_outputs(1593) <= a or b;
    layer1_outputs(1594) <= a;
    layer1_outputs(1595) <= not (a and b);
    layer1_outputs(1596) <= a and not b;
    layer1_outputs(1597) <= a;
    layer1_outputs(1598) <= a;
    layer1_outputs(1599) <= not (a xor b);
    layer1_outputs(1600) <= b;
    layer1_outputs(1601) <= not (a or b);
    layer1_outputs(1602) <= not a;
    layer1_outputs(1603) <= b;
    layer1_outputs(1604) <= a xor b;
    layer1_outputs(1605) <= not a;
    layer1_outputs(1606) <= not b;
    layer1_outputs(1607) <= a;
    layer1_outputs(1608) <= not a;
    layer1_outputs(1609) <= a;
    layer1_outputs(1610) <= not (a xor b);
    layer1_outputs(1611) <= a and b;
    layer1_outputs(1612) <= a or b;
    layer1_outputs(1613) <= a and not b;
    layer1_outputs(1614) <= b;
    layer1_outputs(1615) <= 1'b1;
    layer1_outputs(1616) <= a;
    layer1_outputs(1617) <= b and not a;
    layer1_outputs(1618) <= not (a and b);
    layer1_outputs(1619) <= not a;
    layer1_outputs(1620) <= 1'b1;
    layer1_outputs(1621) <= a or b;
    layer1_outputs(1622) <= not a;
    layer1_outputs(1623) <= not (a or b);
    layer1_outputs(1624) <= b and not a;
    layer1_outputs(1625) <= b;
    layer1_outputs(1626) <= a and b;
    layer1_outputs(1627) <= b;
    layer1_outputs(1628) <= not a or b;
    layer1_outputs(1629) <= a;
    layer1_outputs(1630) <= a and b;
    layer1_outputs(1631) <= not b;
    layer1_outputs(1632) <= b;
    layer1_outputs(1633) <= not (a xor b);
    layer1_outputs(1634) <= a or b;
    layer1_outputs(1635) <= a;
    layer1_outputs(1636) <= a or b;
    layer1_outputs(1637) <= not a or b;
    layer1_outputs(1638) <= not (a xor b);
    layer1_outputs(1639) <= not (a and b);
    layer1_outputs(1640) <= not (a xor b);
    layer1_outputs(1641) <= b and not a;
    layer1_outputs(1642) <= not b;
    layer1_outputs(1643) <= not b or a;
    layer1_outputs(1644) <= not b or a;
    layer1_outputs(1645) <= not b;
    layer1_outputs(1646) <= b;
    layer1_outputs(1647) <= a;
    layer1_outputs(1648) <= b and not a;
    layer1_outputs(1649) <= not a or b;
    layer1_outputs(1650) <= not (a or b);
    layer1_outputs(1651) <= not a or b;
    layer1_outputs(1652) <= 1'b0;
    layer1_outputs(1653) <= a;
    layer1_outputs(1654) <= not (a or b);
    layer1_outputs(1655) <= a and b;
    layer1_outputs(1656) <= a;
    layer1_outputs(1657) <= not (a and b);
    layer1_outputs(1658) <= not (a and b);
    layer1_outputs(1659) <= not (a and b);
    layer1_outputs(1660) <= a;
    layer1_outputs(1661) <= not b or a;
    layer1_outputs(1662) <= not (a xor b);
    layer1_outputs(1663) <= not a or b;
    layer1_outputs(1664) <= a;
    layer1_outputs(1665) <= a and b;
    layer1_outputs(1666) <= a or b;
    layer1_outputs(1667) <= a;
    layer1_outputs(1668) <= not a;
    layer1_outputs(1669) <= not (a or b);
    layer1_outputs(1670) <= not a;
    layer1_outputs(1671) <= not (a and b);
    layer1_outputs(1672) <= not a;
    layer1_outputs(1673) <= not (a and b);
    layer1_outputs(1674) <= a and b;
    layer1_outputs(1675) <= not (a xor b);
    layer1_outputs(1676) <= b and not a;
    layer1_outputs(1677) <= a and not b;
    layer1_outputs(1678) <= not b;
    layer1_outputs(1679) <= b;
    layer1_outputs(1680) <= not a or b;
    layer1_outputs(1681) <= a and not b;
    layer1_outputs(1682) <= not (a or b);
    layer1_outputs(1683) <= 1'b0;
    layer1_outputs(1684) <= b and not a;
    layer1_outputs(1685) <= not (a xor b);
    layer1_outputs(1686) <= a or b;
    layer1_outputs(1687) <= a and b;
    layer1_outputs(1688) <= a and not b;
    layer1_outputs(1689) <= a or b;
    layer1_outputs(1690) <= not b;
    layer1_outputs(1691) <= not a or b;
    layer1_outputs(1692) <= not b;
    layer1_outputs(1693) <= not b or a;
    layer1_outputs(1694) <= a and not b;
    layer1_outputs(1695) <= b;
    layer1_outputs(1696) <= a;
    layer1_outputs(1697) <= a and b;
    layer1_outputs(1698) <= a and not b;
    layer1_outputs(1699) <= not (a xor b);
    layer1_outputs(1700) <= not a or b;
    layer1_outputs(1701) <= b;
    layer1_outputs(1702) <= not a or b;
    layer1_outputs(1703) <= a and not b;
    layer1_outputs(1704) <= not (a and b);
    layer1_outputs(1705) <= not b or a;
    layer1_outputs(1706) <= b;
    layer1_outputs(1707) <= not a or b;
    layer1_outputs(1708) <= not (a and b);
    layer1_outputs(1709) <= a and not b;
    layer1_outputs(1710) <= not b;
    layer1_outputs(1711) <= a and b;
    layer1_outputs(1712) <= a and not b;
    layer1_outputs(1713) <= a and b;
    layer1_outputs(1714) <= a and not b;
    layer1_outputs(1715) <= b and not a;
    layer1_outputs(1716) <= a xor b;
    layer1_outputs(1717) <= b and not a;
    layer1_outputs(1718) <= not (a and b);
    layer1_outputs(1719) <= not (a xor b);
    layer1_outputs(1720) <= a and not b;
    layer1_outputs(1721) <= not (a and b);
    layer1_outputs(1722) <= a and b;
    layer1_outputs(1723) <= a and not b;
    layer1_outputs(1724) <= not a or b;
    layer1_outputs(1725) <= a xor b;
    layer1_outputs(1726) <= not a;
    layer1_outputs(1727) <= a or b;
    layer1_outputs(1728) <= not b or a;
    layer1_outputs(1729) <= not (a and b);
    layer1_outputs(1730) <= a and b;
    layer1_outputs(1731) <= a;
    layer1_outputs(1732) <= b and not a;
    layer1_outputs(1733) <= not b or a;
    layer1_outputs(1734) <= a;
    layer1_outputs(1735) <= a or b;
    layer1_outputs(1736) <= a;
    layer1_outputs(1737) <= b and not a;
    layer1_outputs(1738) <= a and not b;
    layer1_outputs(1739) <= b;
    layer1_outputs(1740) <= not (a xor b);
    layer1_outputs(1741) <= not b or a;
    layer1_outputs(1742) <= a;
    layer1_outputs(1743) <= a and not b;
    layer1_outputs(1744) <= b;
    layer1_outputs(1745) <= not b;
    layer1_outputs(1746) <= not (a or b);
    layer1_outputs(1747) <= a;
    layer1_outputs(1748) <= not b or a;
    layer1_outputs(1749) <= a or b;
    layer1_outputs(1750) <= not b;
    layer1_outputs(1751) <= not (a or b);
    layer1_outputs(1752) <= not b or a;
    layer1_outputs(1753) <= a and not b;
    layer1_outputs(1754) <= b;
    layer1_outputs(1755) <= 1'b0;
    layer1_outputs(1756) <= 1'b1;
    layer1_outputs(1757) <= not b;
    layer1_outputs(1758) <= a and b;
    layer1_outputs(1759) <= not a or b;
    layer1_outputs(1760) <= not b or a;
    layer1_outputs(1761) <= a or b;
    layer1_outputs(1762) <= not b or a;
    layer1_outputs(1763) <= a and not b;
    layer1_outputs(1764) <= not (a and b);
    layer1_outputs(1765) <= a and not b;
    layer1_outputs(1766) <= not a or b;
    layer1_outputs(1767) <= b;
    layer1_outputs(1768) <= not b;
    layer1_outputs(1769) <= not (a or b);
    layer1_outputs(1770) <= not b;
    layer1_outputs(1771) <= a and b;
    layer1_outputs(1772) <= not (a or b);
    layer1_outputs(1773) <= 1'b0;
    layer1_outputs(1774) <= not b or a;
    layer1_outputs(1775) <= not (a xor b);
    layer1_outputs(1776) <= not (a or b);
    layer1_outputs(1777) <= not (a xor b);
    layer1_outputs(1778) <= not (a and b);
    layer1_outputs(1779) <= 1'b1;
    layer1_outputs(1780) <= not b;
    layer1_outputs(1781) <= b and not a;
    layer1_outputs(1782) <= not b;
    layer1_outputs(1783) <= not (a xor b);
    layer1_outputs(1784) <= not (a or b);
    layer1_outputs(1785) <= not (a and b);
    layer1_outputs(1786) <= a and b;
    layer1_outputs(1787) <= b and not a;
    layer1_outputs(1788) <= not a;
    layer1_outputs(1789) <= a and not b;
    layer1_outputs(1790) <= not (a or b);
    layer1_outputs(1791) <= a or b;
    layer1_outputs(1792) <= b;
    layer1_outputs(1793) <= a;
    layer1_outputs(1794) <= not b or a;
    layer1_outputs(1795) <= a and b;
    layer1_outputs(1796) <= 1'b0;
    layer1_outputs(1797) <= 1'b0;
    layer1_outputs(1798) <= not (a xor b);
    layer1_outputs(1799) <= not b;
    layer1_outputs(1800) <= not (a and b);
    layer1_outputs(1801) <= not b;
    layer1_outputs(1802) <= not a or b;
    layer1_outputs(1803) <= a and not b;
    layer1_outputs(1804) <= not (a and b);
    layer1_outputs(1805) <= not (a or b);
    layer1_outputs(1806) <= not b or a;
    layer1_outputs(1807) <= not a;
    layer1_outputs(1808) <= not a;
    layer1_outputs(1809) <= a and not b;
    layer1_outputs(1810) <= not (a and b);
    layer1_outputs(1811) <= not a;
    layer1_outputs(1812) <= not (a or b);
    layer1_outputs(1813) <= b;
    layer1_outputs(1814) <= a or b;
    layer1_outputs(1815) <= a and b;
    layer1_outputs(1816) <= not (a or b);
    layer1_outputs(1817) <= not a;
    layer1_outputs(1818) <= a and b;
    layer1_outputs(1819) <= not (a and b);
    layer1_outputs(1820) <= not (a and b);
    layer1_outputs(1821) <= b;
    layer1_outputs(1822) <= b and not a;
    layer1_outputs(1823) <= a or b;
    layer1_outputs(1824) <= a and not b;
    layer1_outputs(1825) <= not (a or b);
    layer1_outputs(1826) <= a or b;
    layer1_outputs(1827) <= a and b;
    layer1_outputs(1828) <= a xor b;
    layer1_outputs(1829) <= not a or b;
    layer1_outputs(1830) <= a and not b;
    layer1_outputs(1831) <= a;
    layer1_outputs(1832) <= b and not a;
    layer1_outputs(1833) <= not (a xor b);
    layer1_outputs(1834) <= 1'b0;
    layer1_outputs(1835) <= not b or a;
    layer1_outputs(1836) <= not a;
    layer1_outputs(1837) <= not (a and b);
    layer1_outputs(1838) <= a and not b;
    layer1_outputs(1839) <= a;
    layer1_outputs(1840) <= a xor b;
    layer1_outputs(1841) <= a;
    layer1_outputs(1842) <= not b;
    layer1_outputs(1843) <= a;
    layer1_outputs(1844) <= a or b;
    layer1_outputs(1845) <= a;
    layer1_outputs(1846) <= a;
    layer1_outputs(1847) <= a and not b;
    layer1_outputs(1848) <= not (a or b);
    layer1_outputs(1849) <= a xor b;
    layer1_outputs(1850) <= b;
    layer1_outputs(1851) <= a and b;
    layer1_outputs(1852) <= not b or a;
    layer1_outputs(1853) <= a and b;
    layer1_outputs(1854) <= not (a xor b);
    layer1_outputs(1855) <= a xor b;
    layer1_outputs(1856) <= not b;
    layer1_outputs(1857) <= not b;
    layer1_outputs(1858) <= b and not a;
    layer1_outputs(1859) <= a;
    layer1_outputs(1860) <= a and b;
    layer1_outputs(1861) <= 1'b1;
    layer1_outputs(1862) <= a and not b;
    layer1_outputs(1863) <= not (a xor b);
    layer1_outputs(1864) <= a and not b;
    layer1_outputs(1865) <= a and b;
    layer1_outputs(1866) <= b;
    layer1_outputs(1867) <= b and not a;
    layer1_outputs(1868) <= a or b;
    layer1_outputs(1869) <= not (a or b);
    layer1_outputs(1870) <= not a or b;
    layer1_outputs(1871) <= a xor b;
    layer1_outputs(1872) <= a and b;
    layer1_outputs(1873) <= b;
    layer1_outputs(1874) <= a and not b;
    layer1_outputs(1875) <= a or b;
    layer1_outputs(1876) <= not (a xor b);
    layer1_outputs(1877) <= not (a or b);
    layer1_outputs(1878) <= a and b;
    layer1_outputs(1879) <= not a or b;
    layer1_outputs(1880) <= not a;
    layer1_outputs(1881) <= 1'b1;
    layer1_outputs(1882) <= not b or a;
    layer1_outputs(1883) <= not (a or b);
    layer1_outputs(1884) <= a or b;
    layer1_outputs(1885) <= a and b;
    layer1_outputs(1886) <= not b or a;
    layer1_outputs(1887) <= a and not b;
    layer1_outputs(1888) <= b and not a;
    layer1_outputs(1889) <= not a or b;
    layer1_outputs(1890) <= a;
    layer1_outputs(1891) <= a;
    layer1_outputs(1892) <= b and not a;
    layer1_outputs(1893) <= not b;
    layer1_outputs(1894) <= not (a or b);
    layer1_outputs(1895) <= not a or b;
    layer1_outputs(1896) <= a or b;
    layer1_outputs(1897) <= a or b;
    layer1_outputs(1898) <= a and not b;
    layer1_outputs(1899) <= a and b;
    layer1_outputs(1900) <= b and not a;
    layer1_outputs(1901) <= b;
    layer1_outputs(1902) <= a and not b;
    layer1_outputs(1903) <= not b;
    layer1_outputs(1904) <= a;
    layer1_outputs(1905) <= a or b;
    layer1_outputs(1906) <= a and not b;
    layer1_outputs(1907) <= a and b;
    layer1_outputs(1908) <= not a or b;
    layer1_outputs(1909) <= not (a and b);
    layer1_outputs(1910) <= 1'b0;
    layer1_outputs(1911) <= a and not b;
    layer1_outputs(1912) <= a or b;
    layer1_outputs(1913) <= not b or a;
    layer1_outputs(1914) <= a xor b;
    layer1_outputs(1915) <= b and not a;
    layer1_outputs(1916) <= not b;
    layer1_outputs(1917) <= not b or a;
    layer1_outputs(1918) <= b;
    layer1_outputs(1919) <= b;
    layer1_outputs(1920) <= not a or b;
    layer1_outputs(1921) <= not a;
    layer1_outputs(1922) <= not b or a;
    layer1_outputs(1923) <= not a;
    layer1_outputs(1924) <= not (a xor b);
    layer1_outputs(1925) <= a and b;
    layer1_outputs(1926) <= a or b;
    layer1_outputs(1927) <= a;
    layer1_outputs(1928) <= a and b;
    layer1_outputs(1929) <= a;
    layer1_outputs(1930) <= not b;
    layer1_outputs(1931) <= not b;
    layer1_outputs(1932) <= not b;
    layer1_outputs(1933) <= not a;
    layer1_outputs(1934) <= a xor b;
    layer1_outputs(1935) <= a and b;
    layer1_outputs(1936) <= b and not a;
    layer1_outputs(1937) <= b;
    layer1_outputs(1938) <= b and not a;
    layer1_outputs(1939) <= b and not a;
    layer1_outputs(1940) <= b;
    layer1_outputs(1941) <= not (a or b);
    layer1_outputs(1942) <= a xor b;
    layer1_outputs(1943) <= a or b;
    layer1_outputs(1944) <= b;
    layer1_outputs(1945) <= b;
    layer1_outputs(1946) <= b and not a;
    layer1_outputs(1947) <= not b;
    layer1_outputs(1948) <= a or b;
    layer1_outputs(1949) <= not (a xor b);
    layer1_outputs(1950) <= not b;
    layer1_outputs(1951) <= a or b;
    layer1_outputs(1952) <= a and b;
    layer1_outputs(1953) <= not b;
    layer1_outputs(1954) <= not a;
    layer1_outputs(1955) <= not a or b;
    layer1_outputs(1956) <= a and b;
    layer1_outputs(1957) <= not a or b;
    layer1_outputs(1958) <= not a;
    layer1_outputs(1959) <= not (a xor b);
    layer1_outputs(1960) <= not (a or b);
    layer1_outputs(1961) <= b;
    layer1_outputs(1962) <= not (a or b);
    layer1_outputs(1963) <= not b or a;
    layer1_outputs(1964) <= a and not b;
    layer1_outputs(1965) <= a xor b;
    layer1_outputs(1966) <= b and not a;
    layer1_outputs(1967) <= a and b;
    layer1_outputs(1968) <= not b or a;
    layer1_outputs(1969) <= not b or a;
    layer1_outputs(1970) <= b and not a;
    layer1_outputs(1971) <= a;
    layer1_outputs(1972) <= not (a xor b);
    layer1_outputs(1973) <= not b;
    layer1_outputs(1974) <= a;
    layer1_outputs(1975) <= a;
    layer1_outputs(1976) <= not (a or b);
    layer1_outputs(1977) <= not (a or b);
    layer1_outputs(1978) <= a and b;
    layer1_outputs(1979) <= a and b;
    layer1_outputs(1980) <= a and not b;
    layer1_outputs(1981) <= b;
    layer1_outputs(1982) <= not (a and b);
    layer1_outputs(1983) <= not b or a;
    layer1_outputs(1984) <= not a;
    layer1_outputs(1985) <= not a;
    layer1_outputs(1986) <= not a or b;
    layer1_outputs(1987) <= 1'b1;
    layer1_outputs(1988) <= b and not a;
    layer1_outputs(1989) <= not (a and b);
    layer1_outputs(1990) <= a and b;
    layer1_outputs(1991) <= not b;
    layer1_outputs(1992) <= a or b;
    layer1_outputs(1993) <= a;
    layer1_outputs(1994) <= a and b;
    layer1_outputs(1995) <= b and not a;
    layer1_outputs(1996) <= not (a and b);
    layer1_outputs(1997) <= not b or a;
    layer1_outputs(1998) <= not a;
    layer1_outputs(1999) <= not (a and b);
    layer1_outputs(2000) <= b and not a;
    layer1_outputs(2001) <= b and not a;
    layer1_outputs(2002) <= not (a xor b);
    layer1_outputs(2003) <= a;
    layer1_outputs(2004) <= 1'b1;
    layer1_outputs(2005) <= a or b;
    layer1_outputs(2006) <= b and not a;
    layer1_outputs(2007) <= b;
    layer1_outputs(2008) <= not a or b;
    layer1_outputs(2009) <= not b;
    layer1_outputs(2010) <= not a or b;
    layer1_outputs(2011) <= not a;
    layer1_outputs(2012) <= not (a and b);
    layer1_outputs(2013) <= b and not a;
    layer1_outputs(2014) <= not b or a;
    layer1_outputs(2015) <= b;
    layer1_outputs(2016) <= b;
    layer1_outputs(2017) <= not a;
    layer1_outputs(2018) <= a xor b;
    layer1_outputs(2019) <= not a;
    layer1_outputs(2020) <= b;
    layer1_outputs(2021) <= not b or a;
    layer1_outputs(2022) <= not b;
    layer1_outputs(2023) <= not (a or b);
    layer1_outputs(2024) <= not a;
    layer1_outputs(2025) <= b;
    layer1_outputs(2026) <= a or b;
    layer1_outputs(2027) <= not b;
    layer1_outputs(2028) <= a;
    layer1_outputs(2029) <= not b or a;
    layer1_outputs(2030) <= not b;
    layer1_outputs(2031) <= not a or b;
    layer1_outputs(2032) <= a or b;
    layer1_outputs(2033) <= a;
    layer1_outputs(2034) <= a;
    layer1_outputs(2035) <= b;
    layer1_outputs(2036) <= a and b;
    layer1_outputs(2037) <= not (a xor b);
    layer1_outputs(2038) <= a or b;
    layer1_outputs(2039) <= not a;
    layer1_outputs(2040) <= a and not b;
    layer1_outputs(2041) <= a;
    layer1_outputs(2042) <= not (a or b);
    layer1_outputs(2043) <= not a;
    layer1_outputs(2044) <= a and b;
    layer1_outputs(2045) <= b and not a;
    layer1_outputs(2046) <= not (a or b);
    layer1_outputs(2047) <= not (a or b);
    layer1_outputs(2048) <= not (a or b);
    layer1_outputs(2049) <= not (a and b);
    layer1_outputs(2050) <= a;
    layer1_outputs(2051) <= b and not a;
    layer1_outputs(2052) <= b;
    layer1_outputs(2053) <= not a or b;
    layer1_outputs(2054) <= not a;
    layer1_outputs(2055) <= not b;
    layer1_outputs(2056) <= a;
    layer1_outputs(2057) <= not b;
    layer1_outputs(2058) <= a or b;
    layer1_outputs(2059) <= a and b;
    layer1_outputs(2060) <= a or b;
    layer1_outputs(2061) <= not (a xor b);
    layer1_outputs(2062) <= not b or a;
    layer1_outputs(2063) <= not (a xor b);
    layer1_outputs(2064) <= a;
    layer1_outputs(2065) <= not (a and b);
    layer1_outputs(2066) <= not a or b;
    layer1_outputs(2067) <= a and not b;
    layer1_outputs(2068) <= not b;
    layer1_outputs(2069) <= not (a xor b);
    layer1_outputs(2070) <= a xor b;
    layer1_outputs(2071) <= a and not b;
    layer1_outputs(2072) <= not b or a;
    layer1_outputs(2073) <= a or b;
    layer1_outputs(2074) <= a and not b;
    layer1_outputs(2075) <= b;
    layer1_outputs(2076) <= not b;
    layer1_outputs(2077) <= a xor b;
    layer1_outputs(2078) <= not (a xor b);
    layer1_outputs(2079) <= b;
    layer1_outputs(2080) <= a and not b;
    layer1_outputs(2081) <= a or b;
    layer1_outputs(2082) <= not b or a;
    layer1_outputs(2083) <= not (a or b);
    layer1_outputs(2084) <= not b;
    layer1_outputs(2085) <= not (a xor b);
    layer1_outputs(2086) <= a and b;
    layer1_outputs(2087) <= a xor b;
    layer1_outputs(2088) <= b;
    layer1_outputs(2089) <= not a;
    layer1_outputs(2090) <= b and not a;
    layer1_outputs(2091) <= a xor b;
    layer1_outputs(2092) <= not a or b;
    layer1_outputs(2093) <= not (a or b);
    layer1_outputs(2094) <= b;
    layer1_outputs(2095) <= not (a xor b);
    layer1_outputs(2096) <= not b or a;
    layer1_outputs(2097) <= a xor b;
    layer1_outputs(2098) <= not b;
    layer1_outputs(2099) <= not a;
    layer1_outputs(2100) <= not a or b;
    layer1_outputs(2101) <= not a;
    layer1_outputs(2102) <= not b or a;
    layer1_outputs(2103) <= not a or b;
    layer1_outputs(2104) <= a or b;
    layer1_outputs(2105) <= not a;
    layer1_outputs(2106) <= a;
    layer1_outputs(2107) <= not (a or b);
    layer1_outputs(2108) <= a;
    layer1_outputs(2109) <= a or b;
    layer1_outputs(2110) <= a or b;
    layer1_outputs(2111) <= a and b;
    layer1_outputs(2112) <= not a;
    layer1_outputs(2113) <= not b or a;
    layer1_outputs(2114) <= a and b;
    layer1_outputs(2115) <= not (a xor b);
    layer1_outputs(2116) <= b and not a;
    layer1_outputs(2117) <= a xor b;
    layer1_outputs(2118) <= not a;
    layer1_outputs(2119) <= not b or a;
    layer1_outputs(2120) <= b;
    layer1_outputs(2121) <= b;
    layer1_outputs(2122) <= not b or a;
    layer1_outputs(2123) <= 1'b1;
    layer1_outputs(2124) <= not b;
    layer1_outputs(2125) <= b;
    layer1_outputs(2126) <= a xor b;
    layer1_outputs(2127) <= not a or b;
    layer1_outputs(2128) <= not a or b;
    layer1_outputs(2129) <= not b;
    layer1_outputs(2130) <= not a;
    layer1_outputs(2131) <= a and not b;
    layer1_outputs(2132) <= a and not b;
    layer1_outputs(2133) <= not a;
    layer1_outputs(2134) <= not (a xor b);
    layer1_outputs(2135) <= b and not a;
    layer1_outputs(2136) <= not (a xor b);
    layer1_outputs(2137) <= b and not a;
    layer1_outputs(2138) <= a;
    layer1_outputs(2139) <= not (a and b);
    layer1_outputs(2140) <= a and b;
    layer1_outputs(2141) <= a;
    layer1_outputs(2142) <= not b;
    layer1_outputs(2143) <= a and not b;
    layer1_outputs(2144) <= a xor b;
    layer1_outputs(2145) <= not a;
    layer1_outputs(2146) <= not (a and b);
    layer1_outputs(2147) <= not (a xor b);
    layer1_outputs(2148) <= a and not b;
    layer1_outputs(2149) <= b;
    layer1_outputs(2150) <= not b or a;
    layer1_outputs(2151) <= a;
    layer1_outputs(2152) <= not (a and b);
    layer1_outputs(2153) <= not b;
    layer1_outputs(2154) <= not b;
    layer1_outputs(2155) <= a and not b;
    layer1_outputs(2156) <= a and not b;
    layer1_outputs(2157) <= a xor b;
    layer1_outputs(2158) <= not (a xor b);
    layer1_outputs(2159) <= not a;
    layer1_outputs(2160) <= not b;
    layer1_outputs(2161) <= not (a and b);
    layer1_outputs(2162) <= b and not a;
    layer1_outputs(2163) <= not a;
    layer1_outputs(2164) <= a;
    layer1_outputs(2165) <= a;
    layer1_outputs(2166) <= not (a xor b);
    layer1_outputs(2167) <= a and not b;
    layer1_outputs(2168) <= not (a or b);
    layer1_outputs(2169) <= not a or b;
    layer1_outputs(2170) <= not (a xor b);
    layer1_outputs(2171) <= not (a xor b);
    layer1_outputs(2172) <= not a or b;
    layer1_outputs(2173) <= not b;
    layer1_outputs(2174) <= a and b;
    layer1_outputs(2175) <= a or b;
    layer1_outputs(2176) <= not a;
    layer1_outputs(2177) <= a;
    layer1_outputs(2178) <= a and b;
    layer1_outputs(2179) <= not (a and b);
    layer1_outputs(2180) <= not (a and b);
    layer1_outputs(2181) <= a and b;
    layer1_outputs(2182) <= not (a and b);
    layer1_outputs(2183) <= a and not b;
    layer1_outputs(2184) <= not a;
    layer1_outputs(2185) <= not (a and b);
    layer1_outputs(2186) <= a xor b;
    layer1_outputs(2187) <= a;
    layer1_outputs(2188) <= not b;
    layer1_outputs(2189) <= not a;
    layer1_outputs(2190) <= b and not a;
    layer1_outputs(2191) <= a xor b;
    layer1_outputs(2192) <= not b;
    layer1_outputs(2193) <= 1'b1;
    layer1_outputs(2194) <= not a;
    layer1_outputs(2195) <= a and b;
    layer1_outputs(2196) <= 1'b0;
    layer1_outputs(2197) <= a and not b;
    layer1_outputs(2198) <= not b or a;
    layer1_outputs(2199) <= b;
    layer1_outputs(2200) <= b and not a;
    layer1_outputs(2201) <= not a;
    layer1_outputs(2202) <= a;
    layer1_outputs(2203) <= not b;
    layer1_outputs(2204) <= not (a xor b);
    layer1_outputs(2205) <= not (a and b);
    layer1_outputs(2206) <= b and not a;
    layer1_outputs(2207) <= b and not a;
    layer1_outputs(2208) <= 1'b0;
    layer1_outputs(2209) <= a and not b;
    layer1_outputs(2210) <= b and not a;
    layer1_outputs(2211) <= a;
    layer1_outputs(2212) <= not b or a;
    layer1_outputs(2213) <= a or b;
    layer1_outputs(2214) <= a xor b;
    layer1_outputs(2215) <= not b or a;
    layer1_outputs(2216) <= not (a or b);
    layer1_outputs(2217) <= not b;
    layer1_outputs(2218) <= not (a or b);
    layer1_outputs(2219) <= a;
    layer1_outputs(2220) <= 1'b0;
    layer1_outputs(2221) <= not b;
    layer1_outputs(2222) <= a or b;
    layer1_outputs(2223) <= not (a xor b);
    layer1_outputs(2224) <= a xor b;
    layer1_outputs(2225) <= not b or a;
    layer1_outputs(2226) <= b and not a;
    layer1_outputs(2227) <= not (a or b);
    layer1_outputs(2228) <= not (a and b);
    layer1_outputs(2229) <= not b;
    layer1_outputs(2230) <= a and not b;
    layer1_outputs(2231) <= not a or b;
    layer1_outputs(2232) <= not (a xor b);
    layer1_outputs(2233) <= b and not a;
    layer1_outputs(2234) <= 1'b1;
    layer1_outputs(2235) <= a or b;
    layer1_outputs(2236) <= not (a and b);
    layer1_outputs(2237) <= a and not b;
    layer1_outputs(2238) <= not b;
    layer1_outputs(2239) <= a or b;
    layer1_outputs(2240) <= 1'b1;
    layer1_outputs(2241) <= not a or b;
    layer1_outputs(2242) <= not (a or b);
    layer1_outputs(2243) <= a and b;
    layer1_outputs(2244) <= a or b;
    layer1_outputs(2245) <= a;
    layer1_outputs(2246) <= not (a and b);
    layer1_outputs(2247) <= b;
    layer1_outputs(2248) <= a and not b;
    layer1_outputs(2249) <= not a;
    layer1_outputs(2250) <= not a;
    layer1_outputs(2251) <= not (a xor b);
    layer1_outputs(2252) <= not a or b;
    layer1_outputs(2253) <= not a;
    layer1_outputs(2254) <= not (a xor b);
    layer1_outputs(2255) <= not b;
    layer1_outputs(2256) <= a or b;
    layer1_outputs(2257) <= b and not a;
    layer1_outputs(2258) <= not b or a;
    layer1_outputs(2259) <= a and not b;
    layer1_outputs(2260) <= a and b;
    layer1_outputs(2261) <= b;
    layer1_outputs(2262) <= not b;
    layer1_outputs(2263) <= a xor b;
    layer1_outputs(2264) <= not a;
    layer1_outputs(2265) <= not (a xor b);
    layer1_outputs(2266) <= a;
    layer1_outputs(2267) <= not a;
    layer1_outputs(2268) <= a;
    layer1_outputs(2269) <= b and not a;
    layer1_outputs(2270) <= 1'b1;
    layer1_outputs(2271) <= a;
    layer1_outputs(2272) <= not (a xor b);
    layer1_outputs(2273) <= b and not a;
    layer1_outputs(2274) <= not a or b;
    layer1_outputs(2275) <= not a or b;
    layer1_outputs(2276) <= not (a or b);
    layer1_outputs(2277) <= a or b;
    layer1_outputs(2278) <= a and b;
    layer1_outputs(2279) <= a xor b;
    layer1_outputs(2280) <= not b;
    layer1_outputs(2281) <= a or b;
    layer1_outputs(2282) <= not a or b;
    layer1_outputs(2283) <= b;
    layer1_outputs(2284) <= a and not b;
    layer1_outputs(2285) <= a and b;
    layer1_outputs(2286) <= b and not a;
    layer1_outputs(2287) <= a and not b;
    layer1_outputs(2288) <= a or b;
    layer1_outputs(2289) <= a or b;
    layer1_outputs(2290) <= a xor b;
    layer1_outputs(2291) <= not b or a;
    layer1_outputs(2292) <= not a or b;
    layer1_outputs(2293) <= b;
    layer1_outputs(2294) <= not (a and b);
    layer1_outputs(2295) <= not (a or b);
    layer1_outputs(2296) <= b;
    layer1_outputs(2297) <= b;
    layer1_outputs(2298) <= not (a xor b);
    layer1_outputs(2299) <= not b;
    layer1_outputs(2300) <= b;
    layer1_outputs(2301) <= b and not a;
    layer1_outputs(2302) <= not (a or b);
    layer1_outputs(2303) <= a and b;
    layer1_outputs(2304) <= not (a and b);
    layer1_outputs(2305) <= a;
    layer1_outputs(2306) <= not (a and b);
    layer1_outputs(2307) <= not b or a;
    layer1_outputs(2308) <= not a or b;
    layer1_outputs(2309) <= not b or a;
    layer1_outputs(2310) <= not b or a;
    layer1_outputs(2311) <= not (a and b);
    layer1_outputs(2312) <= not (a xor b);
    layer1_outputs(2313) <= a;
    layer1_outputs(2314) <= not a;
    layer1_outputs(2315) <= a;
    layer1_outputs(2316) <= not (a or b);
    layer1_outputs(2317) <= b;
    layer1_outputs(2318) <= b;
    layer1_outputs(2319) <= a and b;
    layer1_outputs(2320) <= b;
    layer1_outputs(2321) <= b and not a;
    layer1_outputs(2322) <= a xor b;
    layer1_outputs(2323) <= not a;
    layer1_outputs(2324) <= not b;
    layer1_outputs(2325) <= not b or a;
    layer1_outputs(2326) <= b and not a;
    layer1_outputs(2327) <= not b;
    layer1_outputs(2328) <= 1'b1;
    layer1_outputs(2329) <= a and not b;
    layer1_outputs(2330) <= not a or b;
    layer1_outputs(2331) <= not b;
    layer1_outputs(2332) <= not a;
    layer1_outputs(2333) <= not a;
    layer1_outputs(2334) <= not (a or b);
    layer1_outputs(2335) <= not (a or b);
    layer1_outputs(2336) <= not a;
    layer1_outputs(2337) <= b;
    layer1_outputs(2338) <= not a or b;
    layer1_outputs(2339) <= b;
    layer1_outputs(2340) <= b;
    layer1_outputs(2341) <= a and b;
    layer1_outputs(2342) <= not a or b;
    layer1_outputs(2343) <= 1'b0;
    layer1_outputs(2344) <= a and not b;
    layer1_outputs(2345) <= a and not b;
    layer1_outputs(2346) <= not b;
    layer1_outputs(2347) <= b and not a;
    layer1_outputs(2348) <= a xor b;
    layer1_outputs(2349) <= not b or a;
    layer1_outputs(2350) <= b and not a;
    layer1_outputs(2351) <= not b;
    layer1_outputs(2352) <= not b;
    layer1_outputs(2353) <= a and not b;
    layer1_outputs(2354) <= a;
    layer1_outputs(2355) <= not b;
    layer1_outputs(2356) <= not (a and b);
    layer1_outputs(2357) <= b;
    layer1_outputs(2358) <= a;
    layer1_outputs(2359) <= not a or b;
    layer1_outputs(2360) <= a and b;
    layer1_outputs(2361) <= not b or a;
    layer1_outputs(2362) <= not b;
    layer1_outputs(2363) <= not a or b;
    layer1_outputs(2364) <= not (a or b);
    layer1_outputs(2365) <= not (a or b);
    layer1_outputs(2366) <= not b;
    layer1_outputs(2367) <= b and not a;
    layer1_outputs(2368) <= a;
    layer1_outputs(2369) <= a or b;
    layer1_outputs(2370) <= not a;
    layer1_outputs(2371) <= a and b;
    layer1_outputs(2372) <= a or b;
    layer1_outputs(2373) <= a and b;
    layer1_outputs(2374) <= b and not a;
    layer1_outputs(2375) <= not b or a;
    layer1_outputs(2376) <= a or b;
    layer1_outputs(2377) <= a and not b;
    layer1_outputs(2378) <= not b;
    layer1_outputs(2379) <= b;
    layer1_outputs(2380) <= 1'b0;
    layer1_outputs(2381) <= not a;
    layer1_outputs(2382) <= not a or b;
    layer1_outputs(2383) <= not a or b;
    layer1_outputs(2384) <= b and not a;
    layer1_outputs(2385) <= a and b;
    layer1_outputs(2386) <= a and b;
    layer1_outputs(2387) <= a and b;
    layer1_outputs(2388) <= a;
    layer1_outputs(2389) <= not b or a;
    layer1_outputs(2390) <= a and b;
    layer1_outputs(2391) <= not (a and b);
    layer1_outputs(2392) <= 1'b1;
    layer1_outputs(2393) <= not (a or b);
    layer1_outputs(2394) <= a and b;
    layer1_outputs(2395) <= not (a and b);
    layer1_outputs(2396) <= b;
    layer1_outputs(2397) <= not b or a;
    layer1_outputs(2398) <= not a or b;
    layer1_outputs(2399) <= b and not a;
    layer1_outputs(2400) <= b and not a;
    layer1_outputs(2401) <= not (a or b);
    layer1_outputs(2402) <= not b or a;
    layer1_outputs(2403) <= not a or b;
    layer1_outputs(2404) <= a or b;
    layer1_outputs(2405) <= not b;
    layer1_outputs(2406) <= not b;
    layer1_outputs(2407) <= not (a and b);
    layer1_outputs(2408) <= not (a or b);
    layer1_outputs(2409) <= not b or a;
    layer1_outputs(2410) <= a and b;
    layer1_outputs(2411) <= a or b;
    layer1_outputs(2412) <= not (a and b);
    layer1_outputs(2413) <= not b;
    layer1_outputs(2414) <= a;
    layer1_outputs(2415) <= not a or b;
    layer1_outputs(2416) <= b and not a;
    layer1_outputs(2417) <= not b;
    layer1_outputs(2418) <= a;
    layer1_outputs(2419) <= a xor b;
    layer1_outputs(2420) <= b;
    layer1_outputs(2421) <= not (a and b);
    layer1_outputs(2422) <= b;
    layer1_outputs(2423) <= not a;
    layer1_outputs(2424) <= a xor b;
    layer1_outputs(2425) <= a;
    layer1_outputs(2426) <= b;
    layer1_outputs(2427) <= not a or b;
    layer1_outputs(2428) <= a;
    layer1_outputs(2429) <= not b or a;
    layer1_outputs(2430) <= a;
    layer1_outputs(2431) <= b and not a;
    layer1_outputs(2432) <= b and not a;
    layer1_outputs(2433) <= not (a xor b);
    layer1_outputs(2434) <= a xor b;
    layer1_outputs(2435) <= not a;
    layer1_outputs(2436) <= not (a xor b);
    layer1_outputs(2437) <= not a;
    layer1_outputs(2438) <= a and not b;
    layer1_outputs(2439) <= b;
    layer1_outputs(2440) <= a and not b;
    layer1_outputs(2441) <= a;
    layer1_outputs(2442) <= b;
    layer1_outputs(2443) <= not (a xor b);
    layer1_outputs(2444) <= a and not b;
    layer1_outputs(2445) <= a xor b;
    layer1_outputs(2446) <= a;
    layer1_outputs(2447) <= not (a or b);
    layer1_outputs(2448) <= a and not b;
    layer1_outputs(2449) <= not a or b;
    layer1_outputs(2450) <= not a or b;
    layer1_outputs(2451) <= 1'b0;
    layer1_outputs(2452) <= b;
    layer1_outputs(2453) <= a;
    layer1_outputs(2454) <= not (a or b);
    layer1_outputs(2455) <= not b or a;
    layer1_outputs(2456) <= a and b;
    layer1_outputs(2457) <= not (a or b);
    layer1_outputs(2458) <= a and b;
    layer1_outputs(2459) <= not a;
    layer1_outputs(2460) <= not (a xor b);
    layer1_outputs(2461) <= not (a xor b);
    layer1_outputs(2462) <= b;
    layer1_outputs(2463) <= not (a xor b);
    layer1_outputs(2464) <= b and not a;
    layer1_outputs(2465) <= not b;
    layer1_outputs(2466) <= a or b;
    layer1_outputs(2467) <= not (a xor b);
    layer1_outputs(2468) <= not a or b;
    layer1_outputs(2469) <= not a or b;
    layer1_outputs(2470) <= a or b;
    layer1_outputs(2471) <= not b or a;
    layer1_outputs(2472) <= not b or a;
    layer1_outputs(2473) <= not b;
    layer1_outputs(2474) <= a and b;
    layer1_outputs(2475) <= not b;
    layer1_outputs(2476) <= a or b;
    layer1_outputs(2477) <= a and not b;
    layer1_outputs(2478) <= not a or b;
    layer1_outputs(2479) <= a and b;
    layer1_outputs(2480) <= not (a or b);
    layer1_outputs(2481) <= a and b;
    layer1_outputs(2482) <= b;
    layer1_outputs(2483) <= not b;
    layer1_outputs(2484) <= not a;
    layer1_outputs(2485) <= b;
    layer1_outputs(2486) <= not a or b;
    layer1_outputs(2487) <= b;
    layer1_outputs(2488) <= a and not b;
    layer1_outputs(2489) <= not b or a;
    layer1_outputs(2490) <= b;
    layer1_outputs(2491) <= not b;
    layer1_outputs(2492) <= not (a and b);
    layer1_outputs(2493) <= a and b;
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= not (a and b);
    layer1_outputs(2496) <= 1'b0;
    layer1_outputs(2497) <= not b;
    layer1_outputs(2498) <= a;
    layer1_outputs(2499) <= not (a xor b);
    layer1_outputs(2500) <= not b or a;
    layer1_outputs(2501) <= not a;
    layer1_outputs(2502) <= not (a and b);
    layer1_outputs(2503) <= b;
    layer1_outputs(2504) <= not (a xor b);
    layer1_outputs(2505) <= a or b;
    layer1_outputs(2506) <= not a or b;
    layer1_outputs(2507) <= b;
    layer1_outputs(2508) <= not a;
    layer1_outputs(2509) <= a;
    layer1_outputs(2510) <= b and not a;
    layer1_outputs(2511) <= 1'b0;
    layer1_outputs(2512) <= not (a or b);
    layer1_outputs(2513) <= not (a and b);
    layer1_outputs(2514) <= not b or a;
    layer1_outputs(2515) <= b;
    layer1_outputs(2516) <= b and not a;
    layer1_outputs(2517) <= a and b;
    layer1_outputs(2518) <= not b or a;
    layer1_outputs(2519) <= not (a xor b);
    layer1_outputs(2520) <= a and b;
    layer1_outputs(2521) <= not a or b;
    layer1_outputs(2522) <= 1'b1;
    layer1_outputs(2523) <= not (a or b);
    layer1_outputs(2524) <= a or b;
    layer1_outputs(2525) <= not b or a;
    layer1_outputs(2526) <= not b;
    layer1_outputs(2527) <= not b;
    layer1_outputs(2528) <= b;
    layer1_outputs(2529) <= not a;
    layer1_outputs(2530) <= 1'b0;
    layer1_outputs(2531) <= a or b;
    layer1_outputs(2532) <= b and not a;
    layer1_outputs(2533) <= a;
    layer1_outputs(2534) <= a and b;
    layer1_outputs(2535) <= not a;
    layer1_outputs(2536) <= a xor b;
    layer1_outputs(2537) <= b;
    layer1_outputs(2538) <= a;
    layer1_outputs(2539) <= a or b;
    layer1_outputs(2540) <= not (a xor b);
    layer1_outputs(2541) <= not a or b;
    layer1_outputs(2542) <= not b or a;
    layer1_outputs(2543) <= not b or a;
    layer1_outputs(2544) <= not b;
    layer1_outputs(2545) <= not b or a;
    layer1_outputs(2546) <= a and b;
    layer1_outputs(2547) <= not (a or b);
    layer1_outputs(2548) <= not a or b;
    layer1_outputs(2549) <= not a;
    layer1_outputs(2550) <= not (a or b);
    layer1_outputs(2551) <= b and not a;
    layer1_outputs(2552) <= not (a and b);
    layer1_outputs(2553) <= b;
    layer1_outputs(2554) <= not (a or b);
    layer1_outputs(2555) <= a and b;
    layer1_outputs(2556) <= b and not a;
    layer1_outputs(2557) <= a and b;
    layer1_outputs(2558) <= a xor b;
    layer1_outputs(2559) <= not b;
    layer1_outputs(2560) <= not b or a;
    layer1_outputs(2561) <= not b or a;
    layer1_outputs(2562) <= a or b;
    layer1_outputs(2563) <= a;
    layer1_outputs(2564) <= a and b;
    layer1_outputs(2565) <= not a or b;
    layer1_outputs(2566) <= a xor b;
    layer1_outputs(2567) <= a and b;
    layer1_outputs(2568) <= not (a and b);
    layer1_outputs(2569) <= a or b;
    layer1_outputs(2570) <= not (a or b);
    layer1_outputs(2571) <= not a or b;
    layer1_outputs(2572) <= not a;
    layer1_outputs(2573) <= a or b;
    layer1_outputs(2574) <= not a;
    layer1_outputs(2575) <= not (a xor b);
    layer1_outputs(2576) <= not a;
    layer1_outputs(2577) <= not (a or b);
    layer1_outputs(2578) <= not (a xor b);
    layer1_outputs(2579) <= not a;
    layer1_outputs(2580) <= a or b;
    layer1_outputs(2581) <= not b;
    layer1_outputs(2582) <= b and not a;
    layer1_outputs(2583) <= a and b;
    layer1_outputs(2584) <= a or b;
    layer1_outputs(2585) <= not a or b;
    layer1_outputs(2586) <= not (a or b);
    layer1_outputs(2587) <= not b;
    layer1_outputs(2588) <= b;
    layer1_outputs(2589) <= b and not a;
    layer1_outputs(2590) <= not b or a;
    layer1_outputs(2591) <= not b or a;
    layer1_outputs(2592) <= not b;
    layer1_outputs(2593) <= not b or a;
    layer1_outputs(2594) <= 1'b1;
    layer1_outputs(2595) <= a or b;
    layer1_outputs(2596) <= b and not a;
    layer1_outputs(2597) <= a and b;
    layer1_outputs(2598) <= a and not b;
    layer1_outputs(2599) <= a and b;
    layer1_outputs(2600) <= a or b;
    layer1_outputs(2601) <= not (a or b);
    layer1_outputs(2602) <= b and not a;
    layer1_outputs(2603) <= not a or b;
    layer1_outputs(2604) <= a;
    layer1_outputs(2605) <= a and b;
    layer1_outputs(2606) <= b;
    layer1_outputs(2607) <= not (a and b);
    layer1_outputs(2608) <= a;
    layer1_outputs(2609) <= b;
    layer1_outputs(2610) <= not (a xor b);
    layer1_outputs(2611) <= not b;
    layer1_outputs(2612) <= b;
    layer1_outputs(2613) <= b;
    layer1_outputs(2614) <= b;
    layer1_outputs(2615) <= 1'b0;
    layer1_outputs(2616) <= not a or b;
    layer1_outputs(2617) <= not b;
    layer1_outputs(2618) <= b and not a;
    layer1_outputs(2619) <= a;
    layer1_outputs(2620) <= a or b;
    layer1_outputs(2621) <= not b or a;
    layer1_outputs(2622) <= not (a and b);
    layer1_outputs(2623) <= not (a xor b);
    layer1_outputs(2624) <= a;
    layer1_outputs(2625) <= not (a xor b);
    layer1_outputs(2626) <= not b;
    layer1_outputs(2627) <= a or b;
    layer1_outputs(2628) <= not a or b;
    layer1_outputs(2629) <= b;
    layer1_outputs(2630) <= not b or a;
    layer1_outputs(2631) <= not b or a;
    layer1_outputs(2632) <= not b;
    layer1_outputs(2633) <= not (a and b);
    layer1_outputs(2634) <= not (a or b);
    layer1_outputs(2635) <= not b;
    layer1_outputs(2636) <= not a;
    layer1_outputs(2637) <= a or b;
    layer1_outputs(2638) <= b and not a;
    layer1_outputs(2639) <= not (a or b);
    layer1_outputs(2640) <= a and b;
    layer1_outputs(2641) <= not (a and b);
    layer1_outputs(2642) <= a;
    layer1_outputs(2643) <= 1'b0;
    layer1_outputs(2644) <= not a or b;
    layer1_outputs(2645) <= not b;
    layer1_outputs(2646) <= a and b;
    layer1_outputs(2647) <= 1'b0;
    layer1_outputs(2648) <= not (a xor b);
    layer1_outputs(2649) <= not b or a;
    layer1_outputs(2650) <= a and b;
    layer1_outputs(2651) <= not b;
    layer1_outputs(2652) <= a;
    layer1_outputs(2653) <= a and b;
    layer1_outputs(2654) <= b;
    layer1_outputs(2655) <= a or b;
    layer1_outputs(2656) <= not a or b;
    layer1_outputs(2657) <= b and not a;
    layer1_outputs(2658) <= not a;
    layer1_outputs(2659) <= a or b;
    layer1_outputs(2660) <= b;
    layer1_outputs(2661) <= b;
    layer1_outputs(2662) <= a;
    layer1_outputs(2663) <= b;
    layer1_outputs(2664) <= 1'b0;
    layer1_outputs(2665) <= not a or b;
    layer1_outputs(2666) <= a and not b;
    layer1_outputs(2667) <= a;
    layer1_outputs(2668) <= not (a or b);
    layer1_outputs(2669) <= a and not b;
    layer1_outputs(2670) <= a or b;
    layer1_outputs(2671) <= not (a xor b);
    layer1_outputs(2672) <= not (a and b);
    layer1_outputs(2673) <= 1'b0;
    layer1_outputs(2674) <= not (a xor b);
    layer1_outputs(2675) <= a and b;
    layer1_outputs(2676) <= b;
    layer1_outputs(2677) <= b and not a;
    layer1_outputs(2678) <= a xor b;
    layer1_outputs(2679) <= a xor b;
    layer1_outputs(2680) <= b and not a;
    layer1_outputs(2681) <= a and b;
    layer1_outputs(2682) <= a and b;
    layer1_outputs(2683) <= a or b;
    layer1_outputs(2684) <= not (a or b);
    layer1_outputs(2685) <= b and not a;
    layer1_outputs(2686) <= b;
    layer1_outputs(2687) <= b and not a;
    layer1_outputs(2688) <= b;
    layer1_outputs(2689) <= not a;
    layer1_outputs(2690) <= not (a or b);
    layer1_outputs(2691) <= 1'b1;
    layer1_outputs(2692) <= not a;
    layer1_outputs(2693) <= a or b;
    layer1_outputs(2694) <= a and not b;
    layer1_outputs(2695) <= not (a and b);
    layer1_outputs(2696) <= a xor b;
    layer1_outputs(2697) <= not a;
    layer1_outputs(2698) <= b;
    layer1_outputs(2699) <= not b;
    layer1_outputs(2700) <= b and not a;
    layer1_outputs(2701) <= a or b;
    layer1_outputs(2702) <= not a or b;
    layer1_outputs(2703) <= a and b;
    layer1_outputs(2704) <= a;
    layer1_outputs(2705) <= not (a xor b);
    layer1_outputs(2706) <= b and not a;
    layer1_outputs(2707) <= not b or a;
    layer1_outputs(2708) <= not b or a;
    layer1_outputs(2709) <= not b;
    layer1_outputs(2710) <= not a;
    layer1_outputs(2711) <= a;
    layer1_outputs(2712) <= b and not a;
    layer1_outputs(2713) <= not (a xor b);
    layer1_outputs(2714) <= b;
    layer1_outputs(2715) <= not b;
    layer1_outputs(2716) <= a;
    layer1_outputs(2717) <= a xor b;
    layer1_outputs(2718) <= not b;
    layer1_outputs(2719) <= a;
    layer1_outputs(2720) <= a or b;
    layer1_outputs(2721) <= not b;
    layer1_outputs(2722) <= 1'b0;
    layer1_outputs(2723) <= 1'b1;
    layer1_outputs(2724) <= not (a and b);
    layer1_outputs(2725) <= a or b;
    layer1_outputs(2726) <= not a;
    layer1_outputs(2727) <= a and not b;
    layer1_outputs(2728) <= b;
    layer1_outputs(2729) <= not a;
    layer1_outputs(2730) <= not (a and b);
    layer1_outputs(2731) <= not b;
    layer1_outputs(2732) <= a xor b;
    layer1_outputs(2733) <= not a or b;
    layer1_outputs(2734) <= not (a xor b);
    layer1_outputs(2735) <= a and not b;
    layer1_outputs(2736) <= a and not b;
    layer1_outputs(2737) <= not a or b;
    layer1_outputs(2738) <= not a;
    layer1_outputs(2739) <= not (a and b);
    layer1_outputs(2740) <= a and not b;
    layer1_outputs(2741) <= not a or b;
    layer1_outputs(2742) <= not a or b;
    layer1_outputs(2743) <= a and b;
    layer1_outputs(2744) <= not b or a;
    layer1_outputs(2745) <= b;
    layer1_outputs(2746) <= not b;
    layer1_outputs(2747) <= not (a or b);
    layer1_outputs(2748) <= a and b;
    layer1_outputs(2749) <= not a or b;
    layer1_outputs(2750) <= not b or a;
    layer1_outputs(2751) <= not (a or b);
    layer1_outputs(2752) <= a;
    layer1_outputs(2753) <= a or b;
    layer1_outputs(2754) <= a;
    layer1_outputs(2755) <= a and b;
    layer1_outputs(2756) <= a xor b;
    layer1_outputs(2757) <= not (a or b);
    layer1_outputs(2758) <= a and not b;
    layer1_outputs(2759) <= not b;
    layer1_outputs(2760) <= not b or a;
    layer1_outputs(2761) <= not a or b;
    layer1_outputs(2762) <= a or b;
    layer1_outputs(2763) <= not (a and b);
    layer1_outputs(2764) <= a xor b;
    layer1_outputs(2765) <= not a;
    layer1_outputs(2766) <= a xor b;
    layer1_outputs(2767) <= not (a or b);
    layer1_outputs(2768) <= not (a and b);
    layer1_outputs(2769) <= a xor b;
    layer1_outputs(2770) <= a or b;
    layer1_outputs(2771) <= not (a or b);
    layer1_outputs(2772) <= b and not a;
    layer1_outputs(2773) <= not b;
    layer1_outputs(2774) <= a;
    layer1_outputs(2775) <= a xor b;
    layer1_outputs(2776) <= b;
    layer1_outputs(2777) <= not (a or b);
    layer1_outputs(2778) <= not b;
    layer1_outputs(2779) <= b and not a;
    layer1_outputs(2780) <= b and not a;
    layer1_outputs(2781) <= not a;
    layer1_outputs(2782) <= b;
    layer1_outputs(2783) <= not b or a;
    layer1_outputs(2784) <= 1'b1;
    layer1_outputs(2785) <= not a or b;
    layer1_outputs(2786) <= b;
    layer1_outputs(2787) <= not a or b;
    layer1_outputs(2788) <= not (a and b);
    layer1_outputs(2789) <= a or b;
    layer1_outputs(2790) <= a;
    layer1_outputs(2791) <= not b;
    layer1_outputs(2792) <= b;
    layer1_outputs(2793) <= b;
    layer1_outputs(2794) <= not a;
    layer1_outputs(2795) <= not a;
    layer1_outputs(2796) <= a or b;
    layer1_outputs(2797) <= b and not a;
    layer1_outputs(2798) <= a;
    layer1_outputs(2799) <= a xor b;
    layer1_outputs(2800) <= b;
    layer1_outputs(2801) <= a or b;
    layer1_outputs(2802) <= not b or a;
    layer1_outputs(2803) <= not (a or b);
    layer1_outputs(2804) <= a;
    layer1_outputs(2805) <= not a;
    layer1_outputs(2806) <= b;
    layer1_outputs(2807) <= b and not a;
    layer1_outputs(2808) <= a and not b;
    layer1_outputs(2809) <= not (a xor b);
    layer1_outputs(2810) <= 1'b1;
    layer1_outputs(2811) <= not (a xor b);
    layer1_outputs(2812) <= not b or a;
    layer1_outputs(2813) <= a and b;
    layer1_outputs(2814) <= not (a xor b);
    layer1_outputs(2815) <= a;
    layer1_outputs(2816) <= a or b;
    layer1_outputs(2817) <= a or b;
    layer1_outputs(2818) <= a or b;
    layer1_outputs(2819) <= a and not b;
    layer1_outputs(2820) <= a or b;
    layer1_outputs(2821) <= a or b;
    layer1_outputs(2822) <= a;
    layer1_outputs(2823) <= b;
    layer1_outputs(2824) <= not a;
    layer1_outputs(2825) <= a and not b;
    layer1_outputs(2826) <= not b;
    layer1_outputs(2827) <= a or b;
    layer1_outputs(2828) <= b and not a;
    layer1_outputs(2829) <= not (a or b);
    layer1_outputs(2830) <= a;
    layer1_outputs(2831) <= not (a xor b);
    layer1_outputs(2832) <= a;
    layer1_outputs(2833) <= not a or b;
    layer1_outputs(2834) <= a;
    layer1_outputs(2835) <= b;
    layer1_outputs(2836) <= b;
    layer1_outputs(2837) <= a and not b;
    layer1_outputs(2838) <= not a;
    layer1_outputs(2839) <= a xor b;
    layer1_outputs(2840) <= a;
    layer1_outputs(2841) <= a;
    layer1_outputs(2842) <= a xor b;
    layer1_outputs(2843) <= b;
    layer1_outputs(2844) <= not b;
    layer1_outputs(2845) <= not b;
    layer1_outputs(2846) <= b and not a;
    layer1_outputs(2847) <= a;
    layer1_outputs(2848) <= b;
    layer1_outputs(2849) <= not a;
    layer1_outputs(2850) <= not b;
    layer1_outputs(2851) <= not (a or b);
    layer1_outputs(2852) <= not a;
    layer1_outputs(2853) <= b and not a;
    layer1_outputs(2854) <= not a or b;
    layer1_outputs(2855) <= not b;
    layer1_outputs(2856) <= a;
    layer1_outputs(2857) <= not b or a;
    layer1_outputs(2858) <= a xor b;
    layer1_outputs(2859) <= a or b;
    layer1_outputs(2860) <= b;
    layer1_outputs(2861) <= b;
    layer1_outputs(2862) <= not b or a;
    layer1_outputs(2863) <= not (a or b);
    layer1_outputs(2864) <= a xor b;
    layer1_outputs(2865) <= a and not b;
    layer1_outputs(2866) <= a;
    layer1_outputs(2867) <= a xor b;
    layer1_outputs(2868) <= not a;
    layer1_outputs(2869) <= a and b;
    layer1_outputs(2870) <= b;
    layer1_outputs(2871) <= not a;
    layer1_outputs(2872) <= b;
    layer1_outputs(2873) <= a;
    layer1_outputs(2874) <= not a or b;
    layer1_outputs(2875) <= not b or a;
    layer1_outputs(2876) <= not a or b;
    layer1_outputs(2877) <= a and not b;
    layer1_outputs(2878) <= not b;
    layer1_outputs(2879) <= not a;
    layer1_outputs(2880) <= b;
    layer1_outputs(2881) <= a;
    layer1_outputs(2882) <= not b;
    layer1_outputs(2883) <= b;
    layer1_outputs(2884) <= not a;
    layer1_outputs(2885) <= not a;
    layer1_outputs(2886) <= b and not a;
    layer1_outputs(2887) <= not b;
    layer1_outputs(2888) <= 1'b1;
    layer1_outputs(2889) <= not b or a;
    layer1_outputs(2890) <= not b;
    layer1_outputs(2891) <= not b;
    layer1_outputs(2892) <= a or b;
    layer1_outputs(2893) <= a xor b;
    layer1_outputs(2894) <= not b;
    layer1_outputs(2895) <= not a or b;
    layer1_outputs(2896) <= a and b;
    layer1_outputs(2897) <= not (a xor b);
    layer1_outputs(2898) <= not a;
    layer1_outputs(2899) <= a;
    layer1_outputs(2900) <= not b;
    layer1_outputs(2901) <= not a or b;
    layer1_outputs(2902) <= not (a or b);
    layer1_outputs(2903) <= not b;
    layer1_outputs(2904) <= not (a or b);
    layer1_outputs(2905) <= not (a xor b);
    layer1_outputs(2906) <= a and not b;
    layer1_outputs(2907) <= a and not b;
    layer1_outputs(2908) <= b and not a;
    layer1_outputs(2909) <= a;
    layer1_outputs(2910) <= not (a or b);
    layer1_outputs(2911) <= not a;
    layer1_outputs(2912) <= a;
    layer1_outputs(2913) <= a or b;
    layer1_outputs(2914) <= not b or a;
    layer1_outputs(2915) <= not a;
    layer1_outputs(2916) <= not a or b;
    layer1_outputs(2917) <= a;
    layer1_outputs(2918) <= a xor b;
    layer1_outputs(2919) <= not b;
    layer1_outputs(2920) <= not (a and b);
    layer1_outputs(2921) <= a or b;
    layer1_outputs(2922) <= a and not b;
    layer1_outputs(2923) <= a;
    layer1_outputs(2924) <= not b;
    layer1_outputs(2925) <= a or b;
    layer1_outputs(2926) <= b and not a;
    layer1_outputs(2927) <= a;
    layer1_outputs(2928) <= a xor b;
    layer1_outputs(2929) <= a;
    layer1_outputs(2930) <= b;
    layer1_outputs(2931) <= a;
    layer1_outputs(2932) <= not (a and b);
    layer1_outputs(2933) <= not b or a;
    layer1_outputs(2934) <= not (a xor b);
    layer1_outputs(2935) <= a xor b;
    layer1_outputs(2936) <= not a;
    layer1_outputs(2937) <= a and b;
    layer1_outputs(2938) <= b;
    layer1_outputs(2939) <= not a;
    layer1_outputs(2940) <= not a;
    layer1_outputs(2941) <= 1'b1;
    layer1_outputs(2942) <= a and b;
    layer1_outputs(2943) <= not (a and b);
    layer1_outputs(2944) <= a or b;
    layer1_outputs(2945) <= not a or b;
    layer1_outputs(2946) <= b;
    layer1_outputs(2947) <= not b;
    layer1_outputs(2948) <= b;
    layer1_outputs(2949) <= a or b;
    layer1_outputs(2950) <= a;
    layer1_outputs(2951) <= not b or a;
    layer1_outputs(2952) <= not b;
    layer1_outputs(2953) <= a;
    layer1_outputs(2954) <= not a;
    layer1_outputs(2955) <= a or b;
    layer1_outputs(2956) <= a;
    layer1_outputs(2957) <= a xor b;
    layer1_outputs(2958) <= a and not b;
    layer1_outputs(2959) <= a;
    layer1_outputs(2960) <= a or b;
    layer1_outputs(2961) <= not b or a;
    layer1_outputs(2962) <= not (a xor b);
    layer1_outputs(2963) <= not b;
    layer1_outputs(2964) <= b;
    layer1_outputs(2965) <= not a;
    layer1_outputs(2966) <= b;
    layer1_outputs(2967) <= a;
    layer1_outputs(2968) <= a or b;
    layer1_outputs(2969) <= b and not a;
    layer1_outputs(2970) <= a and not b;
    layer1_outputs(2971) <= not a;
    layer1_outputs(2972) <= a or b;
    layer1_outputs(2973) <= not (a xor b);
    layer1_outputs(2974) <= not b;
    layer1_outputs(2975) <= a;
    layer1_outputs(2976) <= not b or a;
    layer1_outputs(2977) <= a and not b;
    layer1_outputs(2978) <= not (a and b);
    layer1_outputs(2979) <= a;
    layer1_outputs(2980) <= 1'b1;
    layer1_outputs(2981) <= a and b;
    layer1_outputs(2982) <= b;
    layer1_outputs(2983) <= a;
    layer1_outputs(2984) <= a and b;
    layer1_outputs(2985) <= b and not a;
    layer1_outputs(2986) <= a and b;
    layer1_outputs(2987) <= not a;
    layer1_outputs(2988) <= b;
    layer1_outputs(2989) <= a and b;
    layer1_outputs(2990) <= b and not a;
    layer1_outputs(2991) <= a and not b;
    layer1_outputs(2992) <= not b;
    layer1_outputs(2993) <= a or b;
    layer1_outputs(2994) <= not (a or b);
    layer1_outputs(2995) <= a;
    layer1_outputs(2996) <= not (a or b);
    layer1_outputs(2997) <= not (a and b);
    layer1_outputs(2998) <= b;
    layer1_outputs(2999) <= not a;
    layer1_outputs(3000) <= a or b;
    layer1_outputs(3001) <= not (a xor b);
    layer1_outputs(3002) <= not (a xor b);
    layer1_outputs(3003) <= b and not a;
    layer1_outputs(3004) <= a and not b;
    layer1_outputs(3005) <= b and not a;
    layer1_outputs(3006) <= b;
    layer1_outputs(3007) <= a or b;
    layer1_outputs(3008) <= a or b;
    layer1_outputs(3009) <= a;
    layer1_outputs(3010) <= a and b;
    layer1_outputs(3011) <= a;
    layer1_outputs(3012) <= a;
    layer1_outputs(3013) <= not (a xor b);
    layer1_outputs(3014) <= not (a and b);
    layer1_outputs(3015) <= a and b;
    layer1_outputs(3016) <= a and not b;
    layer1_outputs(3017) <= b;
    layer1_outputs(3018) <= a;
    layer1_outputs(3019) <= a;
    layer1_outputs(3020) <= not (a or b);
    layer1_outputs(3021) <= a;
    layer1_outputs(3022) <= b;
    layer1_outputs(3023) <= not a;
    layer1_outputs(3024) <= not b;
    layer1_outputs(3025) <= not a;
    layer1_outputs(3026) <= b;
    layer1_outputs(3027) <= not a;
    layer1_outputs(3028) <= a and not b;
    layer1_outputs(3029) <= a;
    layer1_outputs(3030) <= not b;
    layer1_outputs(3031) <= not (a and b);
    layer1_outputs(3032) <= a xor b;
    layer1_outputs(3033) <= b and not a;
    layer1_outputs(3034) <= not (a or b);
    layer1_outputs(3035) <= not a;
    layer1_outputs(3036) <= a and not b;
    layer1_outputs(3037) <= not b or a;
    layer1_outputs(3038) <= not a;
    layer1_outputs(3039) <= a xor b;
    layer1_outputs(3040) <= not (a or b);
    layer1_outputs(3041) <= a or b;
    layer1_outputs(3042) <= 1'b0;
    layer1_outputs(3043) <= not b or a;
    layer1_outputs(3044) <= b and not a;
    layer1_outputs(3045) <= a or b;
    layer1_outputs(3046) <= 1'b1;
    layer1_outputs(3047) <= b;
    layer1_outputs(3048) <= a or b;
    layer1_outputs(3049) <= not (a and b);
    layer1_outputs(3050) <= a xor b;
    layer1_outputs(3051) <= not b or a;
    layer1_outputs(3052) <= not a or b;
    layer1_outputs(3053) <= a and b;
    layer1_outputs(3054) <= a or b;
    layer1_outputs(3055) <= a or b;
    layer1_outputs(3056) <= not (a and b);
    layer1_outputs(3057) <= a;
    layer1_outputs(3058) <= a or b;
    layer1_outputs(3059) <= not a;
    layer1_outputs(3060) <= a xor b;
    layer1_outputs(3061) <= a and not b;
    layer1_outputs(3062) <= not (a xor b);
    layer1_outputs(3063) <= not (a xor b);
    layer1_outputs(3064) <= not (a or b);
    layer1_outputs(3065) <= a and b;
    layer1_outputs(3066) <= not (a and b);
    layer1_outputs(3067) <= a or b;
    layer1_outputs(3068) <= a and b;
    layer1_outputs(3069) <= a and b;
    layer1_outputs(3070) <= not b or a;
    layer1_outputs(3071) <= not (a and b);
    layer1_outputs(3072) <= not (a or b);
    layer1_outputs(3073) <= not (a and b);
    layer1_outputs(3074) <= a and not b;
    layer1_outputs(3075) <= a and not b;
    layer1_outputs(3076) <= not b or a;
    layer1_outputs(3077) <= not (a and b);
    layer1_outputs(3078) <= not a or b;
    layer1_outputs(3079) <= a and not b;
    layer1_outputs(3080) <= b;
    layer1_outputs(3081) <= a;
    layer1_outputs(3082) <= a or b;
    layer1_outputs(3083) <= a and b;
    layer1_outputs(3084) <= not b;
    layer1_outputs(3085) <= not (a xor b);
    layer1_outputs(3086) <= b;
    layer1_outputs(3087) <= not b;
    layer1_outputs(3088) <= not (a or b);
    layer1_outputs(3089) <= a;
    layer1_outputs(3090) <= a;
    layer1_outputs(3091) <= 1'b1;
    layer1_outputs(3092) <= b and not a;
    layer1_outputs(3093) <= b;
    layer1_outputs(3094) <= a and b;
    layer1_outputs(3095) <= a;
    layer1_outputs(3096) <= not b or a;
    layer1_outputs(3097) <= not (a or b);
    layer1_outputs(3098) <= not b;
    layer1_outputs(3099) <= a xor b;
    layer1_outputs(3100) <= a or b;
    layer1_outputs(3101) <= not a;
    layer1_outputs(3102) <= a or b;
    layer1_outputs(3103) <= a and b;
    layer1_outputs(3104) <= a and b;
    layer1_outputs(3105) <= a and not b;
    layer1_outputs(3106) <= a and b;
    layer1_outputs(3107) <= not (a xor b);
    layer1_outputs(3108) <= not (a xor b);
    layer1_outputs(3109) <= not a or b;
    layer1_outputs(3110) <= a xor b;
    layer1_outputs(3111) <= a and not b;
    layer1_outputs(3112) <= a xor b;
    layer1_outputs(3113) <= not b or a;
    layer1_outputs(3114) <= b and not a;
    layer1_outputs(3115) <= a;
    layer1_outputs(3116) <= not (a and b);
    layer1_outputs(3117) <= not (a xor b);
    layer1_outputs(3118) <= b;
    layer1_outputs(3119) <= b;
    layer1_outputs(3120) <= a or b;
    layer1_outputs(3121) <= not a or b;
    layer1_outputs(3122) <= a;
    layer1_outputs(3123) <= not (a or b);
    layer1_outputs(3124) <= not (a xor b);
    layer1_outputs(3125) <= a;
    layer1_outputs(3126) <= a xor b;
    layer1_outputs(3127) <= not (a xor b);
    layer1_outputs(3128) <= not (a and b);
    layer1_outputs(3129) <= b;
    layer1_outputs(3130) <= b;
    layer1_outputs(3131) <= a;
    layer1_outputs(3132) <= not b;
    layer1_outputs(3133) <= a xor b;
    layer1_outputs(3134) <= not (a or b);
    layer1_outputs(3135) <= not (a or b);
    layer1_outputs(3136) <= b and not a;
    layer1_outputs(3137) <= b and not a;
    layer1_outputs(3138) <= not (a xor b);
    layer1_outputs(3139) <= not (a or b);
    layer1_outputs(3140) <= not (a or b);
    layer1_outputs(3141) <= a and not b;
    layer1_outputs(3142) <= b and not a;
    layer1_outputs(3143) <= a;
    layer1_outputs(3144) <= not (a xor b);
    layer1_outputs(3145) <= not (a xor b);
    layer1_outputs(3146) <= a and not b;
    layer1_outputs(3147) <= not (a or b);
    layer1_outputs(3148) <= not (a or b);
    layer1_outputs(3149) <= not (a and b);
    layer1_outputs(3150) <= not (a and b);
    layer1_outputs(3151) <= a or b;
    layer1_outputs(3152) <= a;
    layer1_outputs(3153) <= not b;
    layer1_outputs(3154) <= not (a or b);
    layer1_outputs(3155) <= not b;
    layer1_outputs(3156) <= not (a and b);
    layer1_outputs(3157) <= a and b;
    layer1_outputs(3158) <= not (a or b);
    layer1_outputs(3159) <= not a;
    layer1_outputs(3160) <= b and not a;
    layer1_outputs(3161) <= not (a and b);
    layer1_outputs(3162) <= a;
    layer1_outputs(3163) <= a or b;
    layer1_outputs(3164) <= not b;
    layer1_outputs(3165) <= a and b;
    layer1_outputs(3166) <= not (a xor b);
    layer1_outputs(3167) <= a and b;
    layer1_outputs(3168) <= 1'b0;
    layer1_outputs(3169) <= not (a and b);
    layer1_outputs(3170) <= 1'b0;
    layer1_outputs(3171) <= not a;
    layer1_outputs(3172) <= not b or a;
    layer1_outputs(3173) <= a xor b;
    layer1_outputs(3174) <= not (a xor b);
    layer1_outputs(3175) <= a;
    layer1_outputs(3176) <= b;
    layer1_outputs(3177) <= b;
    layer1_outputs(3178) <= a;
    layer1_outputs(3179) <= not b;
    layer1_outputs(3180) <= b and not a;
    layer1_outputs(3181) <= a;
    layer1_outputs(3182) <= not b or a;
    layer1_outputs(3183) <= a and b;
    layer1_outputs(3184) <= a and b;
    layer1_outputs(3185) <= not a or b;
    layer1_outputs(3186) <= not a or b;
    layer1_outputs(3187) <= a and not b;
    layer1_outputs(3188) <= a xor b;
    layer1_outputs(3189) <= a or b;
    layer1_outputs(3190) <= a and not b;
    layer1_outputs(3191) <= not (a and b);
    layer1_outputs(3192) <= not a;
    layer1_outputs(3193) <= b and not a;
    layer1_outputs(3194) <= a and not b;
    layer1_outputs(3195) <= not b or a;
    layer1_outputs(3196) <= not b;
    layer1_outputs(3197) <= not a;
    layer1_outputs(3198) <= not (a or b);
    layer1_outputs(3199) <= not a;
    layer1_outputs(3200) <= not b;
    layer1_outputs(3201) <= a;
    layer1_outputs(3202) <= a and b;
    layer1_outputs(3203) <= a xor b;
    layer1_outputs(3204) <= b;
    layer1_outputs(3205) <= a or b;
    layer1_outputs(3206) <= a and b;
    layer1_outputs(3207) <= 1'b1;
    layer1_outputs(3208) <= not (a and b);
    layer1_outputs(3209) <= not b;
    layer1_outputs(3210) <= not a or b;
    layer1_outputs(3211) <= not a;
    layer1_outputs(3212) <= not b;
    layer1_outputs(3213) <= a or b;
    layer1_outputs(3214) <= a and b;
    layer1_outputs(3215) <= not b;
    layer1_outputs(3216) <= not a or b;
    layer1_outputs(3217) <= not b;
    layer1_outputs(3218) <= not b or a;
    layer1_outputs(3219) <= 1'b1;
    layer1_outputs(3220) <= a xor b;
    layer1_outputs(3221) <= a and b;
    layer1_outputs(3222) <= not b;
    layer1_outputs(3223) <= not b or a;
    layer1_outputs(3224) <= not b or a;
    layer1_outputs(3225) <= not a;
    layer1_outputs(3226) <= a;
    layer1_outputs(3227) <= a;
    layer1_outputs(3228) <= b;
    layer1_outputs(3229) <= b;
    layer1_outputs(3230) <= not (a xor b);
    layer1_outputs(3231) <= a and not b;
    layer1_outputs(3232) <= not b;
    layer1_outputs(3233) <= b and not a;
    layer1_outputs(3234) <= not (a xor b);
    layer1_outputs(3235) <= a and b;
    layer1_outputs(3236) <= not b;
    layer1_outputs(3237) <= not a or b;
    layer1_outputs(3238) <= not a;
    layer1_outputs(3239) <= not (a or b);
    layer1_outputs(3240) <= not a;
    layer1_outputs(3241) <= not a;
    layer1_outputs(3242) <= not a or b;
    layer1_outputs(3243) <= not b or a;
    layer1_outputs(3244) <= b;
    layer1_outputs(3245) <= b;
    layer1_outputs(3246) <= not a;
    layer1_outputs(3247) <= not a;
    layer1_outputs(3248) <= b and not a;
    layer1_outputs(3249) <= a;
    layer1_outputs(3250) <= a or b;
    layer1_outputs(3251) <= not (a and b);
    layer1_outputs(3252) <= a and b;
    layer1_outputs(3253) <= a xor b;
    layer1_outputs(3254) <= a and not b;
    layer1_outputs(3255) <= a and b;
    layer1_outputs(3256) <= a or b;
    layer1_outputs(3257) <= a and b;
    layer1_outputs(3258) <= not (a and b);
    layer1_outputs(3259) <= not a;
    layer1_outputs(3260) <= not b or a;
    layer1_outputs(3261) <= b and not a;
    layer1_outputs(3262) <= a;
    layer1_outputs(3263) <= a;
    layer1_outputs(3264) <= not a or b;
    layer1_outputs(3265) <= not (a and b);
    layer1_outputs(3266) <= not b;
    layer1_outputs(3267) <= a;
    layer1_outputs(3268) <= b and not a;
    layer1_outputs(3269) <= a and not b;
    layer1_outputs(3270) <= 1'b0;
    layer1_outputs(3271) <= not b or a;
    layer1_outputs(3272) <= not a;
    layer1_outputs(3273) <= not (a and b);
    layer1_outputs(3274) <= b and not a;
    layer1_outputs(3275) <= a xor b;
    layer1_outputs(3276) <= b;
    layer1_outputs(3277) <= a and b;
    layer1_outputs(3278) <= b and not a;
    layer1_outputs(3279) <= b;
    layer1_outputs(3280) <= 1'b0;
    layer1_outputs(3281) <= not a or b;
    layer1_outputs(3282) <= 1'b0;
    layer1_outputs(3283) <= not (a and b);
    layer1_outputs(3284) <= 1'b1;
    layer1_outputs(3285) <= not (a or b);
    layer1_outputs(3286) <= not a;
    layer1_outputs(3287) <= b and not a;
    layer1_outputs(3288) <= b;
    layer1_outputs(3289) <= a or b;
    layer1_outputs(3290) <= not (a or b);
    layer1_outputs(3291) <= b;
    layer1_outputs(3292) <= not (a or b);
    layer1_outputs(3293) <= a and not b;
    layer1_outputs(3294) <= a xor b;
    layer1_outputs(3295) <= a and b;
    layer1_outputs(3296) <= not (a or b);
    layer1_outputs(3297) <= b;
    layer1_outputs(3298) <= b;
    layer1_outputs(3299) <= not (a and b);
    layer1_outputs(3300) <= b;
    layer1_outputs(3301) <= not (a and b);
    layer1_outputs(3302) <= not a or b;
    layer1_outputs(3303) <= not a or b;
    layer1_outputs(3304) <= not (a xor b);
    layer1_outputs(3305) <= a and b;
    layer1_outputs(3306) <= not a or b;
    layer1_outputs(3307) <= not (a or b);
    layer1_outputs(3308) <= a and b;
    layer1_outputs(3309) <= b and not a;
    layer1_outputs(3310) <= b and not a;
    layer1_outputs(3311) <= b;
    layer1_outputs(3312) <= not (a and b);
    layer1_outputs(3313) <= a and not b;
    layer1_outputs(3314) <= a or b;
    layer1_outputs(3315) <= not b;
    layer1_outputs(3316) <= not a or b;
    layer1_outputs(3317) <= a and b;
    layer1_outputs(3318) <= b;
    layer1_outputs(3319) <= a xor b;
    layer1_outputs(3320) <= not b;
    layer1_outputs(3321) <= not (a xor b);
    layer1_outputs(3322) <= not (a xor b);
    layer1_outputs(3323) <= not (a and b);
    layer1_outputs(3324) <= not b;
    layer1_outputs(3325) <= b and not a;
    layer1_outputs(3326) <= b;
    layer1_outputs(3327) <= a and not b;
    layer1_outputs(3328) <= not b;
    layer1_outputs(3329) <= not a or b;
    layer1_outputs(3330) <= not (a xor b);
    layer1_outputs(3331) <= a;
    layer1_outputs(3332) <= not (a or b);
    layer1_outputs(3333) <= a xor b;
    layer1_outputs(3334) <= not a or b;
    layer1_outputs(3335) <= a xor b;
    layer1_outputs(3336) <= not a;
    layer1_outputs(3337) <= not (a xor b);
    layer1_outputs(3338) <= a;
    layer1_outputs(3339) <= b;
    layer1_outputs(3340) <= b and not a;
    layer1_outputs(3341) <= 1'b1;
    layer1_outputs(3342) <= a;
    layer1_outputs(3343) <= not b or a;
    layer1_outputs(3344) <= not a or b;
    layer1_outputs(3345) <= not b or a;
    layer1_outputs(3346) <= a and not b;
    layer1_outputs(3347) <= not b;
    layer1_outputs(3348) <= not (a xor b);
    layer1_outputs(3349) <= not b;
    layer1_outputs(3350) <= b and not a;
    layer1_outputs(3351) <= not a;
    layer1_outputs(3352) <= b;
    layer1_outputs(3353) <= b;
    layer1_outputs(3354) <= b;
    layer1_outputs(3355) <= not a or b;
    layer1_outputs(3356) <= a and not b;
    layer1_outputs(3357) <= a and b;
    layer1_outputs(3358) <= 1'b1;
    layer1_outputs(3359) <= not a;
    layer1_outputs(3360) <= not a or b;
    layer1_outputs(3361) <= not (a or b);
    layer1_outputs(3362) <= a or b;
    layer1_outputs(3363) <= not b;
    layer1_outputs(3364) <= b;
    layer1_outputs(3365) <= b;
    layer1_outputs(3366) <= b;
    layer1_outputs(3367) <= not a or b;
    layer1_outputs(3368) <= a and b;
    layer1_outputs(3369) <= not b;
    layer1_outputs(3370) <= a or b;
    layer1_outputs(3371) <= not (a and b);
    layer1_outputs(3372) <= not (a and b);
    layer1_outputs(3373) <= not a or b;
    layer1_outputs(3374) <= a;
    layer1_outputs(3375) <= not (a and b);
    layer1_outputs(3376) <= not b or a;
    layer1_outputs(3377) <= a;
    layer1_outputs(3378) <= a or b;
    layer1_outputs(3379) <= a and b;
    layer1_outputs(3380) <= a and b;
    layer1_outputs(3381) <= not a or b;
    layer1_outputs(3382) <= b and not a;
    layer1_outputs(3383) <= not a or b;
    layer1_outputs(3384) <= not a or b;
    layer1_outputs(3385) <= a or b;
    layer1_outputs(3386) <= a;
    layer1_outputs(3387) <= not a;
    layer1_outputs(3388) <= a;
    layer1_outputs(3389) <= a and not b;
    layer1_outputs(3390) <= a;
    layer1_outputs(3391) <= b and not a;
    layer1_outputs(3392) <= not (a xor b);
    layer1_outputs(3393) <= a;
    layer1_outputs(3394) <= a or b;
    layer1_outputs(3395) <= a or b;
    layer1_outputs(3396) <= a and not b;
    layer1_outputs(3397) <= a;
    layer1_outputs(3398) <= a or b;
    layer1_outputs(3399) <= a and b;
    layer1_outputs(3400) <= not a or b;
    layer1_outputs(3401) <= not a;
    layer1_outputs(3402) <= a;
    layer1_outputs(3403) <= a;
    layer1_outputs(3404) <= not (a xor b);
    layer1_outputs(3405) <= b and not a;
    layer1_outputs(3406) <= a and b;
    layer1_outputs(3407) <= not a or b;
    layer1_outputs(3408) <= not (a or b);
    layer1_outputs(3409) <= b;
    layer1_outputs(3410) <= b;
    layer1_outputs(3411) <= b and not a;
    layer1_outputs(3412) <= a;
    layer1_outputs(3413) <= 1'b0;
    layer1_outputs(3414) <= not (a and b);
    layer1_outputs(3415) <= a xor b;
    layer1_outputs(3416) <= a and b;
    layer1_outputs(3417) <= a xor b;
    layer1_outputs(3418) <= not (a and b);
    layer1_outputs(3419) <= b;
    layer1_outputs(3420) <= b;
    layer1_outputs(3421) <= not (a and b);
    layer1_outputs(3422) <= not a or b;
    layer1_outputs(3423) <= 1'b1;
    layer1_outputs(3424) <= 1'b0;
    layer1_outputs(3425) <= a and not b;
    layer1_outputs(3426) <= not a or b;
    layer1_outputs(3427) <= not (a and b);
    layer1_outputs(3428) <= 1'b0;
    layer1_outputs(3429) <= 1'b0;
    layer1_outputs(3430) <= not a or b;
    layer1_outputs(3431) <= not a;
    layer1_outputs(3432) <= b;
    layer1_outputs(3433) <= not (a or b);
    layer1_outputs(3434) <= not a or b;
    layer1_outputs(3435) <= a or b;
    layer1_outputs(3436) <= a xor b;
    layer1_outputs(3437) <= not b or a;
    layer1_outputs(3438) <= not (a xor b);
    layer1_outputs(3439) <= not a;
    layer1_outputs(3440) <= a;
    layer1_outputs(3441) <= not a;
    layer1_outputs(3442) <= b;
    layer1_outputs(3443) <= b;
    layer1_outputs(3444) <= not a or b;
    layer1_outputs(3445) <= not a;
    layer1_outputs(3446) <= not b;
    layer1_outputs(3447) <= b;
    layer1_outputs(3448) <= not (a xor b);
    layer1_outputs(3449) <= not (a or b);
    layer1_outputs(3450) <= b and not a;
    layer1_outputs(3451) <= a xor b;
    layer1_outputs(3452) <= a xor b;
    layer1_outputs(3453) <= not (a or b);
    layer1_outputs(3454) <= a and not b;
    layer1_outputs(3455) <= not a or b;
    layer1_outputs(3456) <= a and b;
    layer1_outputs(3457) <= a xor b;
    layer1_outputs(3458) <= a and b;
    layer1_outputs(3459) <= a;
    layer1_outputs(3460) <= not a or b;
    layer1_outputs(3461) <= not b;
    layer1_outputs(3462) <= a and b;
    layer1_outputs(3463) <= 1'b0;
    layer1_outputs(3464) <= not b or a;
    layer1_outputs(3465) <= not (a or b);
    layer1_outputs(3466) <= b and not a;
    layer1_outputs(3467) <= a;
    layer1_outputs(3468) <= b;
    layer1_outputs(3469) <= 1'b0;
    layer1_outputs(3470) <= not b;
    layer1_outputs(3471) <= not (a or b);
    layer1_outputs(3472) <= not a;
    layer1_outputs(3473) <= not (a xor b);
    layer1_outputs(3474) <= 1'b0;
    layer1_outputs(3475) <= a and b;
    layer1_outputs(3476) <= not (a and b);
    layer1_outputs(3477) <= not a;
    layer1_outputs(3478) <= not b or a;
    layer1_outputs(3479) <= not (a xor b);
    layer1_outputs(3480) <= a;
    layer1_outputs(3481) <= b;
    layer1_outputs(3482) <= not b;
    layer1_outputs(3483) <= not a or b;
    layer1_outputs(3484) <= not b or a;
    layer1_outputs(3485) <= a and not b;
    layer1_outputs(3486) <= a or b;
    layer1_outputs(3487) <= a xor b;
    layer1_outputs(3488) <= not (a and b);
    layer1_outputs(3489) <= not a;
    layer1_outputs(3490) <= not (a xor b);
    layer1_outputs(3491) <= b and not a;
    layer1_outputs(3492) <= a and b;
    layer1_outputs(3493) <= not b;
    layer1_outputs(3494) <= not (a or b);
    layer1_outputs(3495) <= not b;
    layer1_outputs(3496) <= a;
    layer1_outputs(3497) <= not a;
    layer1_outputs(3498) <= not a;
    layer1_outputs(3499) <= 1'b1;
    layer1_outputs(3500) <= a xor b;
    layer1_outputs(3501) <= a or b;
    layer1_outputs(3502) <= a;
    layer1_outputs(3503) <= a and b;
    layer1_outputs(3504) <= a and b;
    layer1_outputs(3505) <= b and not a;
    layer1_outputs(3506) <= not (a and b);
    layer1_outputs(3507) <= a or b;
    layer1_outputs(3508) <= not b;
    layer1_outputs(3509) <= not (a or b);
    layer1_outputs(3510) <= not (a xor b);
    layer1_outputs(3511) <= a and b;
    layer1_outputs(3512) <= a and not b;
    layer1_outputs(3513) <= b and not a;
    layer1_outputs(3514) <= a and b;
    layer1_outputs(3515) <= a and not b;
    layer1_outputs(3516) <= not (a and b);
    layer1_outputs(3517) <= b;
    layer1_outputs(3518) <= not (a xor b);
    layer1_outputs(3519) <= b;
    layer1_outputs(3520) <= not a;
    layer1_outputs(3521) <= b and not a;
    layer1_outputs(3522) <= a;
    layer1_outputs(3523) <= not b;
    layer1_outputs(3524) <= not a;
    layer1_outputs(3525) <= not b;
    layer1_outputs(3526) <= b;
    layer1_outputs(3527) <= a xor b;
    layer1_outputs(3528) <= a or b;
    layer1_outputs(3529) <= not b;
    layer1_outputs(3530) <= not b;
    layer1_outputs(3531) <= a and not b;
    layer1_outputs(3532) <= a;
    layer1_outputs(3533) <= not b or a;
    layer1_outputs(3534) <= not b;
    layer1_outputs(3535) <= a or b;
    layer1_outputs(3536) <= not a or b;
    layer1_outputs(3537) <= a;
    layer1_outputs(3538) <= not b;
    layer1_outputs(3539) <= not (a xor b);
    layer1_outputs(3540) <= not (a xor b);
    layer1_outputs(3541) <= not (a or b);
    layer1_outputs(3542) <= not (a or b);
    layer1_outputs(3543) <= not b or a;
    layer1_outputs(3544) <= not a;
    layer1_outputs(3545) <= not b;
    layer1_outputs(3546) <= a xor b;
    layer1_outputs(3547) <= a xor b;
    layer1_outputs(3548) <= not a or b;
    layer1_outputs(3549) <= a and not b;
    layer1_outputs(3550) <= a or b;
    layer1_outputs(3551) <= not a;
    layer1_outputs(3552) <= not (a and b);
    layer1_outputs(3553) <= not b or a;
    layer1_outputs(3554) <= b;
    layer1_outputs(3555) <= b;
    layer1_outputs(3556) <= a;
    layer1_outputs(3557) <= a;
    layer1_outputs(3558) <= not (a or b);
    layer1_outputs(3559) <= a and not b;
    layer1_outputs(3560) <= a xor b;
    layer1_outputs(3561) <= not b or a;
    layer1_outputs(3562) <= not (a xor b);
    layer1_outputs(3563) <= a and not b;
    layer1_outputs(3564) <= a or b;
    layer1_outputs(3565) <= a and not b;
    layer1_outputs(3566) <= 1'b0;
    layer1_outputs(3567) <= not (a or b);
    layer1_outputs(3568) <= a;
    layer1_outputs(3569) <= a;
    layer1_outputs(3570) <= a and b;
    layer1_outputs(3571) <= not b;
    layer1_outputs(3572) <= not (a or b);
    layer1_outputs(3573) <= a and b;
    layer1_outputs(3574) <= not (a and b);
    layer1_outputs(3575) <= not (a or b);
    layer1_outputs(3576) <= b;
    layer1_outputs(3577) <= not (a and b);
    layer1_outputs(3578) <= not (a xor b);
    layer1_outputs(3579) <= a;
    layer1_outputs(3580) <= a and not b;
    layer1_outputs(3581) <= b and not a;
    layer1_outputs(3582) <= a;
    layer1_outputs(3583) <= not b or a;
    layer1_outputs(3584) <= not (a and b);
    layer1_outputs(3585) <= a and b;
    layer1_outputs(3586) <= b;
    layer1_outputs(3587) <= not a or b;
    layer1_outputs(3588) <= a xor b;
    layer1_outputs(3589) <= 1'b0;
    layer1_outputs(3590) <= b and not a;
    layer1_outputs(3591) <= a or b;
    layer1_outputs(3592) <= not (a or b);
    layer1_outputs(3593) <= not b or a;
    layer1_outputs(3594) <= not a or b;
    layer1_outputs(3595) <= a and b;
    layer1_outputs(3596) <= b;
    layer1_outputs(3597) <= 1'b0;
    layer1_outputs(3598) <= a;
    layer1_outputs(3599) <= b;
    layer1_outputs(3600) <= not (a and b);
    layer1_outputs(3601) <= a;
    layer1_outputs(3602) <= not a or b;
    layer1_outputs(3603) <= a;
    layer1_outputs(3604) <= a and b;
    layer1_outputs(3605) <= a and not b;
    layer1_outputs(3606) <= a or b;
    layer1_outputs(3607) <= a or b;
    layer1_outputs(3608) <= not a;
    layer1_outputs(3609) <= not (a xor b);
    layer1_outputs(3610) <= a;
    layer1_outputs(3611) <= not a or b;
    layer1_outputs(3612) <= not b or a;
    layer1_outputs(3613) <= a;
    layer1_outputs(3614) <= 1'b0;
    layer1_outputs(3615) <= a and b;
    layer1_outputs(3616) <= 1'b1;
    layer1_outputs(3617) <= a or b;
    layer1_outputs(3618) <= a;
    layer1_outputs(3619) <= not (a xor b);
    layer1_outputs(3620) <= not a;
    layer1_outputs(3621) <= not (a or b);
    layer1_outputs(3622) <= a;
    layer1_outputs(3623) <= a and not b;
    layer1_outputs(3624) <= a;
    layer1_outputs(3625) <= a and b;
    layer1_outputs(3626) <= not b;
    layer1_outputs(3627) <= a and not b;
    layer1_outputs(3628) <= not (a xor b);
    layer1_outputs(3629) <= not b or a;
    layer1_outputs(3630) <= b and not a;
    layer1_outputs(3631) <= not a or b;
    layer1_outputs(3632) <= not b;
    layer1_outputs(3633) <= a and not b;
    layer1_outputs(3634) <= not (a and b);
    layer1_outputs(3635) <= not a or b;
    layer1_outputs(3636) <= a and b;
    layer1_outputs(3637) <= not a;
    layer1_outputs(3638) <= a and not b;
    layer1_outputs(3639) <= not b;
    layer1_outputs(3640) <= b;
    layer1_outputs(3641) <= b and not a;
    layer1_outputs(3642) <= a;
    layer1_outputs(3643) <= not (a and b);
    layer1_outputs(3644) <= b;
    layer1_outputs(3645) <= not a;
    layer1_outputs(3646) <= not b;
    layer1_outputs(3647) <= a or b;
    layer1_outputs(3648) <= b and not a;
    layer1_outputs(3649) <= b and not a;
    layer1_outputs(3650) <= b;
    layer1_outputs(3651) <= a and not b;
    layer1_outputs(3652) <= 1'b1;
    layer1_outputs(3653) <= not a;
    layer1_outputs(3654) <= not (a or b);
    layer1_outputs(3655) <= not (a and b);
    layer1_outputs(3656) <= not a or b;
    layer1_outputs(3657) <= not a;
    layer1_outputs(3658) <= not a or b;
    layer1_outputs(3659) <= 1'b0;
    layer1_outputs(3660) <= not (a and b);
    layer1_outputs(3661) <= a and not b;
    layer1_outputs(3662) <= 1'b0;
    layer1_outputs(3663) <= b;
    layer1_outputs(3664) <= a and not b;
    layer1_outputs(3665) <= a or b;
    layer1_outputs(3666) <= a xor b;
    layer1_outputs(3667) <= not b;
    layer1_outputs(3668) <= a or b;
    layer1_outputs(3669) <= a xor b;
    layer1_outputs(3670) <= not a;
    layer1_outputs(3671) <= a or b;
    layer1_outputs(3672) <= a and not b;
    layer1_outputs(3673) <= a and not b;
    layer1_outputs(3674) <= not (a or b);
    layer1_outputs(3675) <= a;
    layer1_outputs(3676) <= not a;
    layer1_outputs(3677) <= 1'b1;
    layer1_outputs(3678) <= a or b;
    layer1_outputs(3679) <= a and b;
    layer1_outputs(3680) <= a and b;
    layer1_outputs(3681) <= not (a xor b);
    layer1_outputs(3682) <= a;
    layer1_outputs(3683) <= a or b;
    layer1_outputs(3684) <= a and b;
    layer1_outputs(3685) <= a;
    layer1_outputs(3686) <= not b or a;
    layer1_outputs(3687) <= not (a and b);
    layer1_outputs(3688) <= a;
    layer1_outputs(3689) <= not a;
    layer1_outputs(3690) <= a;
    layer1_outputs(3691) <= a xor b;
    layer1_outputs(3692) <= not (a and b);
    layer1_outputs(3693) <= not a;
    layer1_outputs(3694) <= not a;
    layer1_outputs(3695) <= b;
    layer1_outputs(3696) <= a or b;
    layer1_outputs(3697) <= b and not a;
    layer1_outputs(3698) <= a xor b;
    layer1_outputs(3699) <= not b;
    layer1_outputs(3700) <= not (a or b);
    layer1_outputs(3701) <= a and not b;
    layer1_outputs(3702) <= not b or a;
    layer1_outputs(3703) <= not a;
    layer1_outputs(3704) <= a xor b;
    layer1_outputs(3705) <= not b;
    layer1_outputs(3706) <= b and not a;
    layer1_outputs(3707) <= a and b;
    layer1_outputs(3708) <= b;
    layer1_outputs(3709) <= a;
    layer1_outputs(3710) <= a and b;
    layer1_outputs(3711) <= not (a and b);
    layer1_outputs(3712) <= not (a and b);
    layer1_outputs(3713) <= 1'b0;
    layer1_outputs(3714) <= not (a or b);
    layer1_outputs(3715) <= a and not b;
    layer1_outputs(3716) <= not (a and b);
    layer1_outputs(3717) <= not a;
    layer1_outputs(3718) <= a and not b;
    layer1_outputs(3719) <= b and not a;
    layer1_outputs(3720) <= a and b;
    layer1_outputs(3721) <= not (a or b);
    layer1_outputs(3722) <= a or b;
    layer1_outputs(3723) <= not (a and b);
    layer1_outputs(3724) <= not b or a;
    layer1_outputs(3725) <= b and not a;
    layer1_outputs(3726) <= not b or a;
    layer1_outputs(3727) <= a and not b;
    layer1_outputs(3728) <= not a or b;
    layer1_outputs(3729) <= not (a xor b);
    layer1_outputs(3730) <= a xor b;
    layer1_outputs(3731) <= not a or b;
    layer1_outputs(3732) <= not (a or b);
    layer1_outputs(3733) <= a xor b;
    layer1_outputs(3734) <= b and not a;
    layer1_outputs(3735) <= not a or b;
    layer1_outputs(3736) <= b;
    layer1_outputs(3737) <= 1'b1;
    layer1_outputs(3738) <= not a;
    layer1_outputs(3739) <= not (a xor b);
    layer1_outputs(3740) <= not a;
    layer1_outputs(3741) <= a and b;
    layer1_outputs(3742) <= a;
    layer1_outputs(3743) <= not b or a;
    layer1_outputs(3744) <= b;
    layer1_outputs(3745) <= a and not b;
    layer1_outputs(3746) <= not a or b;
    layer1_outputs(3747) <= not a or b;
    layer1_outputs(3748) <= a and b;
    layer1_outputs(3749) <= b;
    layer1_outputs(3750) <= not a;
    layer1_outputs(3751) <= not a;
    layer1_outputs(3752) <= not (a xor b);
    layer1_outputs(3753) <= a or b;
    layer1_outputs(3754) <= a or b;
    layer1_outputs(3755) <= not b or a;
    layer1_outputs(3756) <= not b;
    layer1_outputs(3757) <= not b;
    layer1_outputs(3758) <= 1'b1;
    layer1_outputs(3759) <= a;
    layer1_outputs(3760) <= not (a xor b);
    layer1_outputs(3761) <= a or b;
    layer1_outputs(3762) <= not b;
    layer1_outputs(3763) <= not a;
    layer1_outputs(3764) <= not a;
    layer1_outputs(3765) <= not a;
    layer1_outputs(3766) <= not (a xor b);
    layer1_outputs(3767) <= not a;
    layer1_outputs(3768) <= a or b;
    layer1_outputs(3769) <= b and not a;
    layer1_outputs(3770) <= a;
    layer1_outputs(3771) <= not b;
    layer1_outputs(3772) <= b and not a;
    layer1_outputs(3773) <= a;
    layer1_outputs(3774) <= not (a or b);
    layer1_outputs(3775) <= a xor b;
    layer1_outputs(3776) <= a and not b;
    layer1_outputs(3777) <= 1'b0;
    layer1_outputs(3778) <= not (a and b);
    layer1_outputs(3779) <= b;
    layer1_outputs(3780) <= not b;
    layer1_outputs(3781) <= not (a or b);
    layer1_outputs(3782) <= a;
    layer1_outputs(3783) <= not a;
    layer1_outputs(3784) <= not (a xor b);
    layer1_outputs(3785) <= a or b;
    layer1_outputs(3786) <= a;
    layer1_outputs(3787) <= not a;
    layer1_outputs(3788) <= a or b;
    layer1_outputs(3789) <= not a or b;
    layer1_outputs(3790) <= a xor b;
    layer1_outputs(3791) <= not a or b;
    layer1_outputs(3792) <= a xor b;
    layer1_outputs(3793) <= a and not b;
    layer1_outputs(3794) <= not a or b;
    layer1_outputs(3795) <= a and not b;
    layer1_outputs(3796) <= a and b;
    layer1_outputs(3797) <= not a or b;
    layer1_outputs(3798) <= a;
    layer1_outputs(3799) <= not (a or b);
    layer1_outputs(3800) <= not (a xor b);
    layer1_outputs(3801) <= a and b;
    layer1_outputs(3802) <= not a;
    layer1_outputs(3803) <= b;
    layer1_outputs(3804) <= not a or b;
    layer1_outputs(3805) <= 1'b1;
    layer1_outputs(3806) <= not a or b;
    layer1_outputs(3807) <= b and not a;
    layer1_outputs(3808) <= 1'b1;
    layer1_outputs(3809) <= a;
    layer1_outputs(3810) <= not (a and b);
    layer1_outputs(3811) <= not (a or b);
    layer1_outputs(3812) <= a or b;
    layer1_outputs(3813) <= a or b;
    layer1_outputs(3814) <= b and not a;
    layer1_outputs(3815) <= a;
    layer1_outputs(3816) <= b;
    layer1_outputs(3817) <= a and not b;
    layer1_outputs(3818) <= b;
    layer1_outputs(3819) <= not a or b;
    layer1_outputs(3820) <= not (a xor b);
    layer1_outputs(3821) <= not (a and b);
    layer1_outputs(3822) <= not (a or b);
    layer1_outputs(3823) <= 1'b0;
    layer1_outputs(3824) <= a;
    layer1_outputs(3825) <= a xor b;
    layer1_outputs(3826) <= not a or b;
    layer1_outputs(3827) <= b and not a;
    layer1_outputs(3828) <= not (a or b);
    layer1_outputs(3829) <= not (a or b);
    layer1_outputs(3830) <= a and b;
    layer1_outputs(3831) <= b and not a;
    layer1_outputs(3832) <= not a;
    layer1_outputs(3833) <= b;
    layer1_outputs(3834) <= a and not b;
    layer1_outputs(3835) <= a and b;
    layer1_outputs(3836) <= b;
    layer1_outputs(3837) <= b and not a;
    layer1_outputs(3838) <= a or b;
    layer1_outputs(3839) <= not (a and b);
    layer1_outputs(3840) <= not a or b;
    layer1_outputs(3841) <= not a;
    layer1_outputs(3842) <= not a;
    layer1_outputs(3843) <= not b or a;
    layer1_outputs(3844) <= b and not a;
    layer1_outputs(3845) <= not b or a;
    layer1_outputs(3846) <= not a;
    layer1_outputs(3847) <= not a or b;
    layer1_outputs(3848) <= a or b;
    layer1_outputs(3849) <= b;
    layer1_outputs(3850) <= not a or b;
    layer1_outputs(3851) <= not b or a;
    layer1_outputs(3852) <= a and not b;
    layer1_outputs(3853) <= a or b;
    layer1_outputs(3854) <= b;
    layer1_outputs(3855) <= not a or b;
    layer1_outputs(3856) <= not b or a;
    layer1_outputs(3857) <= not (a and b);
    layer1_outputs(3858) <= not b;
    layer1_outputs(3859) <= 1'b1;
    layer1_outputs(3860) <= a xor b;
    layer1_outputs(3861) <= not a;
    layer1_outputs(3862) <= not a;
    layer1_outputs(3863) <= b;
    layer1_outputs(3864) <= not (a or b);
    layer1_outputs(3865) <= not (a and b);
    layer1_outputs(3866) <= a xor b;
    layer1_outputs(3867) <= not b or a;
    layer1_outputs(3868) <= not b;
    layer1_outputs(3869) <= a;
    layer1_outputs(3870) <= a and not b;
    layer1_outputs(3871) <= not (a or b);
    layer1_outputs(3872) <= 1'b1;
    layer1_outputs(3873) <= a;
    layer1_outputs(3874) <= not a;
    layer1_outputs(3875) <= a;
    layer1_outputs(3876) <= a and b;
    layer1_outputs(3877) <= a;
    layer1_outputs(3878) <= not b;
    layer1_outputs(3879) <= a and b;
    layer1_outputs(3880) <= not b;
    layer1_outputs(3881) <= not a;
    layer1_outputs(3882) <= not (a or b);
    layer1_outputs(3883) <= not b;
    layer1_outputs(3884) <= not b;
    layer1_outputs(3885) <= b and not a;
    layer1_outputs(3886) <= a xor b;
    layer1_outputs(3887) <= a and b;
    layer1_outputs(3888) <= not b;
    layer1_outputs(3889) <= not a or b;
    layer1_outputs(3890) <= not b or a;
    layer1_outputs(3891) <= a and not b;
    layer1_outputs(3892) <= not (a xor b);
    layer1_outputs(3893) <= a and b;
    layer1_outputs(3894) <= not a;
    layer1_outputs(3895) <= not a or b;
    layer1_outputs(3896) <= not b or a;
    layer1_outputs(3897) <= a or b;
    layer1_outputs(3898) <= a;
    layer1_outputs(3899) <= a and not b;
    layer1_outputs(3900) <= not (a and b);
    layer1_outputs(3901) <= not b;
    layer1_outputs(3902) <= not (a or b);
    layer1_outputs(3903) <= not (a or b);
    layer1_outputs(3904) <= a and b;
    layer1_outputs(3905) <= b and not a;
    layer1_outputs(3906) <= not b;
    layer1_outputs(3907) <= a;
    layer1_outputs(3908) <= a xor b;
    layer1_outputs(3909) <= not a;
    layer1_outputs(3910) <= a and not b;
    layer1_outputs(3911) <= a or b;
    layer1_outputs(3912) <= not b;
    layer1_outputs(3913) <= not a;
    layer1_outputs(3914) <= not (a xor b);
    layer1_outputs(3915) <= b;
    layer1_outputs(3916) <= 1'b0;
    layer1_outputs(3917) <= not a;
    layer1_outputs(3918) <= not (a and b);
    layer1_outputs(3919) <= not (a or b);
    layer1_outputs(3920) <= a;
    layer1_outputs(3921) <= a and not b;
    layer1_outputs(3922) <= b;
    layer1_outputs(3923) <= b;
    layer1_outputs(3924) <= 1'b0;
    layer1_outputs(3925) <= b and not a;
    layer1_outputs(3926) <= not b or a;
    layer1_outputs(3927) <= not a or b;
    layer1_outputs(3928) <= not (a or b);
    layer1_outputs(3929) <= a xor b;
    layer1_outputs(3930) <= not (a and b);
    layer1_outputs(3931) <= not (a or b);
    layer1_outputs(3932) <= a and b;
    layer1_outputs(3933) <= not (a and b);
    layer1_outputs(3934) <= a and b;
    layer1_outputs(3935) <= 1'b1;
    layer1_outputs(3936) <= not b;
    layer1_outputs(3937) <= b and not a;
    layer1_outputs(3938) <= not b or a;
    layer1_outputs(3939) <= a or b;
    layer1_outputs(3940) <= a;
    layer1_outputs(3941) <= a;
    layer1_outputs(3942) <= not b;
    layer1_outputs(3943) <= b;
    layer1_outputs(3944) <= b and not a;
    layer1_outputs(3945) <= b;
    layer1_outputs(3946) <= not (a and b);
    layer1_outputs(3947) <= not b or a;
    layer1_outputs(3948) <= a xor b;
    layer1_outputs(3949) <= not a;
    layer1_outputs(3950) <= b;
    layer1_outputs(3951) <= not (a xor b);
    layer1_outputs(3952) <= not (a or b);
    layer1_outputs(3953) <= a and b;
    layer1_outputs(3954) <= b;
    layer1_outputs(3955) <= b;
    layer1_outputs(3956) <= a and not b;
    layer1_outputs(3957) <= a or b;
    layer1_outputs(3958) <= a;
    layer1_outputs(3959) <= a xor b;
    layer1_outputs(3960) <= a or b;
    layer1_outputs(3961) <= a and not b;
    layer1_outputs(3962) <= not (a or b);
    layer1_outputs(3963) <= not a or b;
    layer1_outputs(3964) <= b and not a;
    layer1_outputs(3965) <= not (a xor b);
    layer1_outputs(3966) <= not (a or b);
    layer1_outputs(3967) <= not b;
    layer1_outputs(3968) <= a xor b;
    layer1_outputs(3969) <= not a;
    layer1_outputs(3970) <= b and not a;
    layer1_outputs(3971) <= not a or b;
    layer1_outputs(3972) <= b and not a;
    layer1_outputs(3973) <= b;
    layer1_outputs(3974) <= a;
    layer1_outputs(3975) <= a xor b;
    layer1_outputs(3976) <= not (a xor b);
    layer1_outputs(3977) <= a and b;
    layer1_outputs(3978) <= a;
    layer1_outputs(3979) <= b and not a;
    layer1_outputs(3980) <= not (a and b);
    layer1_outputs(3981) <= b and not a;
    layer1_outputs(3982) <= b and not a;
    layer1_outputs(3983) <= not (a or b);
    layer1_outputs(3984) <= a;
    layer1_outputs(3985) <= a xor b;
    layer1_outputs(3986) <= not a or b;
    layer1_outputs(3987) <= a and not b;
    layer1_outputs(3988) <= not (a or b);
    layer1_outputs(3989) <= a and not b;
    layer1_outputs(3990) <= a;
    layer1_outputs(3991) <= not (a or b);
    layer1_outputs(3992) <= a or b;
    layer1_outputs(3993) <= not b;
    layer1_outputs(3994) <= not a;
    layer1_outputs(3995) <= not (a and b);
    layer1_outputs(3996) <= not (a xor b);
    layer1_outputs(3997) <= not (a or b);
    layer1_outputs(3998) <= a;
    layer1_outputs(3999) <= not b or a;
    layer1_outputs(4000) <= not a;
    layer1_outputs(4001) <= not (a or b);
    layer1_outputs(4002) <= not a;
    layer1_outputs(4003) <= not a;
    layer1_outputs(4004) <= a or b;
    layer1_outputs(4005) <= a and b;
    layer1_outputs(4006) <= a or b;
    layer1_outputs(4007) <= not a;
    layer1_outputs(4008) <= a or b;
    layer1_outputs(4009) <= a or b;
    layer1_outputs(4010) <= not (a and b);
    layer1_outputs(4011) <= 1'b0;
    layer1_outputs(4012) <= not (a and b);
    layer1_outputs(4013) <= not b or a;
    layer1_outputs(4014) <= b and not a;
    layer1_outputs(4015) <= a xor b;
    layer1_outputs(4016) <= a;
    layer1_outputs(4017) <= a xor b;
    layer1_outputs(4018) <= not (a or b);
    layer1_outputs(4019) <= b;
    layer1_outputs(4020) <= not a;
    layer1_outputs(4021) <= b;
    layer1_outputs(4022) <= a and b;
    layer1_outputs(4023) <= a and not b;
    layer1_outputs(4024) <= not a;
    layer1_outputs(4025) <= a;
    layer1_outputs(4026) <= a and b;
    layer1_outputs(4027) <= not a or b;
    layer1_outputs(4028) <= not a or b;
    layer1_outputs(4029) <= a and not b;
    layer1_outputs(4030) <= a;
    layer1_outputs(4031) <= a and not b;
    layer1_outputs(4032) <= not b or a;
    layer1_outputs(4033) <= b and not a;
    layer1_outputs(4034) <= not (a and b);
    layer1_outputs(4035) <= not b;
    layer1_outputs(4036) <= a xor b;
    layer1_outputs(4037) <= a and b;
    layer1_outputs(4038) <= not b;
    layer1_outputs(4039) <= not b or a;
    layer1_outputs(4040) <= not b;
    layer1_outputs(4041) <= a;
    layer1_outputs(4042) <= not (a and b);
    layer1_outputs(4043) <= not b or a;
    layer1_outputs(4044) <= not (a and b);
    layer1_outputs(4045) <= a xor b;
    layer1_outputs(4046) <= a and not b;
    layer1_outputs(4047) <= not (a xor b);
    layer1_outputs(4048) <= a and b;
    layer1_outputs(4049) <= 1'b0;
    layer1_outputs(4050) <= not b;
    layer1_outputs(4051) <= a or b;
    layer1_outputs(4052) <= a xor b;
    layer1_outputs(4053) <= not b or a;
    layer1_outputs(4054) <= not a or b;
    layer1_outputs(4055) <= not (a or b);
    layer1_outputs(4056) <= a;
    layer1_outputs(4057) <= a xor b;
    layer1_outputs(4058) <= a and b;
    layer1_outputs(4059) <= not (a and b);
    layer1_outputs(4060) <= a or b;
    layer1_outputs(4061) <= not b;
    layer1_outputs(4062) <= a and b;
    layer1_outputs(4063) <= b and not a;
    layer1_outputs(4064) <= a or b;
    layer1_outputs(4065) <= not b;
    layer1_outputs(4066) <= not (a or b);
    layer1_outputs(4067) <= not a or b;
    layer1_outputs(4068) <= b;
    layer1_outputs(4069) <= a;
    layer1_outputs(4070) <= b;
    layer1_outputs(4071) <= not b or a;
    layer1_outputs(4072) <= not a or b;
    layer1_outputs(4073) <= not a or b;
    layer1_outputs(4074) <= b and not a;
    layer1_outputs(4075) <= a and not b;
    layer1_outputs(4076) <= b;
    layer1_outputs(4077) <= not a;
    layer1_outputs(4078) <= not b or a;
    layer1_outputs(4079) <= b and not a;
    layer1_outputs(4080) <= not a;
    layer1_outputs(4081) <= not b;
    layer1_outputs(4082) <= a and not b;
    layer1_outputs(4083) <= not a;
    layer1_outputs(4084) <= b;
    layer1_outputs(4085) <= 1'b0;
    layer1_outputs(4086) <= not (a xor b);
    layer1_outputs(4087) <= a and b;
    layer1_outputs(4088) <= b;
    layer1_outputs(4089) <= b and not a;
    layer1_outputs(4090) <= b;
    layer1_outputs(4091) <= not (a or b);
    layer1_outputs(4092) <= not a;
    layer1_outputs(4093) <= not a or b;
    layer1_outputs(4094) <= not a;
    layer1_outputs(4095) <= not b or a;
    layer1_outputs(4096) <= a xor b;
    layer1_outputs(4097) <= a;
    layer1_outputs(4098) <= not b or a;
    layer1_outputs(4099) <= b;
    layer1_outputs(4100) <= not a;
    layer1_outputs(4101) <= not (a and b);
    layer1_outputs(4102) <= not (a xor b);
    layer1_outputs(4103) <= a xor b;
    layer1_outputs(4104) <= not (a or b);
    layer1_outputs(4105) <= a xor b;
    layer1_outputs(4106) <= b and not a;
    layer1_outputs(4107) <= b and not a;
    layer1_outputs(4108) <= not b;
    layer1_outputs(4109) <= not a or b;
    layer1_outputs(4110) <= a and not b;
    layer1_outputs(4111) <= not (a and b);
    layer1_outputs(4112) <= a;
    layer1_outputs(4113) <= a xor b;
    layer1_outputs(4114) <= not a or b;
    layer1_outputs(4115) <= b and not a;
    layer1_outputs(4116) <= b and not a;
    layer1_outputs(4117) <= a and not b;
    layer1_outputs(4118) <= a;
    layer1_outputs(4119) <= b;
    layer1_outputs(4120) <= a or b;
    layer1_outputs(4121) <= a or b;
    layer1_outputs(4122) <= not a;
    layer1_outputs(4123) <= b and not a;
    layer1_outputs(4124) <= b and not a;
    layer1_outputs(4125) <= not a;
    layer1_outputs(4126) <= b;
    layer1_outputs(4127) <= not b or a;
    layer1_outputs(4128) <= not b;
    layer1_outputs(4129) <= a and not b;
    layer1_outputs(4130) <= not (a or b);
    layer1_outputs(4131) <= a and not b;
    layer1_outputs(4132) <= not (a or b);
    layer1_outputs(4133) <= a and b;
    layer1_outputs(4134) <= b and not a;
    layer1_outputs(4135) <= not a;
    layer1_outputs(4136) <= not (a and b);
    layer1_outputs(4137) <= not (a xor b);
    layer1_outputs(4138) <= b and not a;
    layer1_outputs(4139) <= not a;
    layer1_outputs(4140) <= not (a xor b);
    layer1_outputs(4141) <= not b;
    layer1_outputs(4142) <= not (a xor b);
    layer1_outputs(4143) <= b and not a;
    layer1_outputs(4144) <= not a or b;
    layer1_outputs(4145) <= a;
    layer1_outputs(4146) <= a or b;
    layer1_outputs(4147) <= not (a and b);
    layer1_outputs(4148) <= not b;
    layer1_outputs(4149) <= not b;
    layer1_outputs(4150) <= not b or a;
    layer1_outputs(4151) <= not a or b;
    layer1_outputs(4152) <= a;
    layer1_outputs(4153) <= a or b;
    layer1_outputs(4154) <= not (a and b);
    layer1_outputs(4155) <= not (a and b);
    layer1_outputs(4156) <= a;
    layer1_outputs(4157) <= 1'b1;
    layer1_outputs(4158) <= not (a and b);
    layer1_outputs(4159) <= not (a xor b);
    layer1_outputs(4160) <= not (a or b);
    layer1_outputs(4161) <= not (a or b);
    layer1_outputs(4162) <= b and not a;
    layer1_outputs(4163) <= a;
    layer1_outputs(4164) <= a or b;
    layer1_outputs(4165) <= a or b;
    layer1_outputs(4166) <= a or b;
    layer1_outputs(4167) <= a or b;
    layer1_outputs(4168) <= a and b;
    layer1_outputs(4169) <= a or b;
    layer1_outputs(4170) <= a xor b;
    layer1_outputs(4171) <= not (a and b);
    layer1_outputs(4172) <= a xor b;
    layer1_outputs(4173) <= not (a or b);
    layer1_outputs(4174) <= a xor b;
    layer1_outputs(4175) <= a and b;
    layer1_outputs(4176) <= b and not a;
    layer1_outputs(4177) <= a;
    layer1_outputs(4178) <= not a or b;
    layer1_outputs(4179) <= not b;
    layer1_outputs(4180) <= not (a and b);
    layer1_outputs(4181) <= a;
    layer1_outputs(4182) <= not (a xor b);
    layer1_outputs(4183) <= not b or a;
    layer1_outputs(4184) <= a or b;
    layer1_outputs(4185) <= not a or b;
    layer1_outputs(4186) <= not b;
    layer1_outputs(4187) <= b;
    layer1_outputs(4188) <= not b or a;
    layer1_outputs(4189) <= b and not a;
    layer1_outputs(4190) <= not (a or b);
    layer1_outputs(4191) <= not (a or b);
    layer1_outputs(4192) <= not b or a;
    layer1_outputs(4193) <= not b or a;
    layer1_outputs(4194) <= a and not b;
    layer1_outputs(4195) <= not a;
    layer1_outputs(4196) <= not b;
    layer1_outputs(4197) <= b;
    layer1_outputs(4198) <= not a or b;
    layer1_outputs(4199) <= not a or b;
    layer1_outputs(4200) <= a and not b;
    layer1_outputs(4201) <= b and not a;
    layer1_outputs(4202) <= a and not b;
    layer1_outputs(4203) <= not b;
    layer1_outputs(4204) <= a;
    layer1_outputs(4205) <= not (a and b);
    layer1_outputs(4206) <= b and not a;
    layer1_outputs(4207) <= 1'b1;
    layer1_outputs(4208) <= a and not b;
    layer1_outputs(4209) <= not a or b;
    layer1_outputs(4210) <= not b;
    layer1_outputs(4211) <= not b or a;
    layer1_outputs(4212) <= not b or a;
    layer1_outputs(4213) <= not (a or b);
    layer1_outputs(4214) <= b;
    layer1_outputs(4215) <= a and b;
    layer1_outputs(4216) <= not b;
    layer1_outputs(4217) <= not a;
    layer1_outputs(4218) <= not b or a;
    layer1_outputs(4219) <= a and b;
    layer1_outputs(4220) <= b and not a;
    layer1_outputs(4221) <= b and not a;
    layer1_outputs(4222) <= not b;
    layer1_outputs(4223) <= not a;
    layer1_outputs(4224) <= not b or a;
    layer1_outputs(4225) <= a or b;
    layer1_outputs(4226) <= not a or b;
    layer1_outputs(4227) <= not (a or b);
    layer1_outputs(4228) <= a xor b;
    layer1_outputs(4229) <= not (a and b);
    layer1_outputs(4230) <= 1'b1;
    layer1_outputs(4231) <= not b;
    layer1_outputs(4232) <= a xor b;
    layer1_outputs(4233) <= a;
    layer1_outputs(4234) <= a and not b;
    layer1_outputs(4235) <= not b;
    layer1_outputs(4236) <= a xor b;
    layer1_outputs(4237) <= not a;
    layer1_outputs(4238) <= a or b;
    layer1_outputs(4239) <= not b or a;
    layer1_outputs(4240) <= a;
    layer1_outputs(4241) <= a;
    layer1_outputs(4242) <= b and not a;
    layer1_outputs(4243) <= not b;
    layer1_outputs(4244) <= not (a or b);
    layer1_outputs(4245) <= not a;
    layer1_outputs(4246) <= a and b;
    layer1_outputs(4247) <= a or b;
    layer1_outputs(4248) <= a;
    layer1_outputs(4249) <= not b or a;
    layer1_outputs(4250) <= not (a and b);
    layer1_outputs(4251) <= 1'b0;
    layer1_outputs(4252) <= a and b;
    layer1_outputs(4253) <= a or b;
    layer1_outputs(4254) <= a;
    layer1_outputs(4255) <= not b;
    layer1_outputs(4256) <= a and b;
    layer1_outputs(4257) <= not (a xor b);
    layer1_outputs(4258) <= not (a and b);
    layer1_outputs(4259) <= not a or b;
    layer1_outputs(4260) <= not (a and b);
    layer1_outputs(4261) <= a xor b;
    layer1_outputs(4262) <= a xor b;
    layer1_outputs(4263) <= b;
    layer1_outputs(4264) <= a;
    layer1_outputs(4265) <= a or b;
    layer1_outputs(4266) <= not b;
    layer1_outputs(4267) <= not b or a;
    layer1_outputs(4268) <= not a;
    layer1_outputs(4269) <= a and not b;
    layer1_outputs(4270) <= b;
    layer1_outputs(4271) <= not a;
    layer1_outputs(4272) <= a;
    layer1_outputs(4273) <= a and b;
    layer1_outputs(4274) <= a and not b;
    layer1_outputs(4275) <= a and b;
    layer1_outputs(4276) <= a or b;
    layer1_outputs(4277) <= a and b;
    layer1_outputs(4278) <= not b or a;
    layer1_outputs(4279) <= a or b;
    layer1_outputs(4280) <= not a;
    layer1_outputs(4281) <= a and not b;
    layer1_outputs(4282) <= not (a xor b);
    layer1_outputs(4283) <= not b or a;
    layer1_outputs(4284) <= not b or a;
    layer1_outputs(4285) <= not a or b;
    layer1_outputs(4286) <= a and not b;
    layer1_outputs(4287) <= not a;
    layer1_outputs(4288) <= b;
    layer1_outputs(4289) <= b and not a;
    layer1_outputs(4290) <= not a or b;
    layer1_outputs(4291) <= b;
    layer1_outputs(4292) <= not b;
    layer1_outputs(4293) <= not (a and b);
    layer1_outputs(4294) <= a and not b;
    layer1_outputs(4295) <= a and not b;
    layer1_outputs(4296) <= not b or a;
    layer1_outputs(4297) <= b;
    layer1_outputs(4298) <= not (a or b);
    layer1_outputs(4299) <= a and not b;
    layer1_outputs(4300) <= not a or b;
    layer1_outputs(4301) <= a and not b;
    layer1_outputs(4302) <= b;
    layer1_outputs(4303) <= not a or b;
    layer1_outputs(4304) <= not b or a;
    layer1_outputs(4305) <= a and b;
    layer1_outputs(4306) <= not a;
    layer1_outputs(4307) <= b;
    layer1_outputs(4308) <= not b;
    layer1_outputs(4309) <= not (a or b);
    layer1_outputs(4310) <= not (a and b);
    layer1_outputs(4311) <= b;
    layer1_outputs(4312) <= not (a and b);
    layer1_outputs(4313) <= a;
    layer1_outputs(4314) <= not b;
    layer1_outputs(4315) <= not (a and b);
    layer1_outputs(4316) <= b;
    layer1_outputs(4317) <= not (a or b);
    layer1_outputs(4318) <= not b or a;
    layer1_outputs(4319) <= b;
    layer1_outputs(4320) <= a;
    layer1_outputs(4321) <= not (a and b);
    layer1_outputs(4322) <= a or b;
    layer1_outputs(4323) <= b;
    layer1_outputs(4324) <= not a or b;
    layer1_outputs(4325) <= not a or b;
    layer1_outputs(4326) <= not (a or b);
    layer1_outputs(4327) <= b and not a;
    layer1_outputs(4328) <= b and not a;
    layer1_outputs(4329) <= b and not a;
    layer1_outputs(4330) <= not b or a;
    layer1_outputs(4331) <= not a;
    layer1_outputs(4332) <= not (a and b);
    layer1_outputs(4333) <= not (a or b);
    layer1_outputs(4334) <= b and not a;
    layer1_outputs(4335) <= a or b;
    layer1_outputs(4336) <= not b or a;
    layer1_outputs(4337) <= not a or b;
    layer1_outputs(4338) <= not b;
    layer1_outputs(4339) <= b;
    layer1_outputs(4340) <= a and not b;
    layer1_outputs(4341) <= not b;
    layer1_outputs(4342) <= not (a xor b);
    layer1_outputs(4343) <= not (a and b);
    layer1_outputs(4344) <= b and not a;
    layer1_outputs(4345) <= not b or a;
    layer1_outputs(4346) <= a xor b;
    layer1_outputs(4347) <= a xor b;
    layer1_outputs(4348) <= a and b;
    layer1_outputs(4349) <= b and not a;
    layer1_outputs(4350) <= a xor b;
    layer1_outputs(4351) <= a xor b;
    layer1_outputs(4352) <= b;
    layer1_outputs(4353) <= a and not b;
    layer1_outputs(4354) <= not b;
    layer1_outputs(4355) <= not (a and b);
    layer1_outputs(4356) <= b;
    layer1_outputs(4357) <= not (a xor b);
    layer1_outputs(4358) <= not b;
    layer1_outputs(4359) <= 1'b1;
    layer1_outputs(4360) <= not (a or b);
    layer1_outputs(4361) <= not a;
    layer1_outputs(4362) <= not (a or b);
    layer1_outputs(4363) <= a;
    layer1_outputs(4364) <= not a;
    layer1_outputs(4365) <= a xor b;
    layer1_outputs(4366) <= not a;
    layer1_outputs(4367) <= not (a or b);
    layer1_outputs(4368) <= a xor b;
    layer1_outputs(4369) <= a;
    layer1_outputs(4370) <= not (a and b);
    layer1_outputs(4371) <= a;
    layer1_outputs(4372) <= not a or b;
    layer1_outputs(4373) <= a xor b;
    layer1_outputs(4374) <= not (a and b);
    layer1_outputs(4375) <= not a;
    layer1_outputs(4376) <= a and b;
    layer1_outputs(4377) <= not a or b;
    layer1_outputs(4378) <= not (a or b);
    layer1_outputs(4379) <= not (a and b);
    layer1_outputs(4380) <= a;
    layer1_outputs(4381) <= b;
    layer1_outputs(4382) <= not (a xor b);
    layer1_outputs(4383) <= not b;
    layer1_outputs(4384) <= b and not a;
    layer1_outputs(4385) <= a and b;
    layer1_outputs(4386) <= a or b;
    layer1_outputs(4387) <= not (a xor b);
    layer1_outputs(4388) <= 1'b1;
    layer1_outputs(4389) <= a and not b;
    layer1_outputs(4390) <= a xor b;
    layer1_outputs(4391) <= b;
    layer1_outputs(4392) <= b;
    layer1_outputs(4393) <= a or b;
    layer1_outputs(4394) <= not (a or b);
    layer1_outputs(4395) <= not b or a;
    layer1_outputs(4396) <= a and not b;
    layer1_outputs(4397) <= not (a or b);
    layer1_outputs(4398) <= not (a or b);
    layer1_outputs(4399) <= not (a xor b);
    layer1_outputs(4400) <= a and not b;
    layer1_outputs(4401) <= not (a or b);
    layer1_outputs(4402) <= a;
    layer1_outputs(4403) <= not b or a;
    layer1_outputs(4404) <= a and not b;
    layer1_outputs(4405) <= not b;
    layer1_outputs(4406) <= a and b;
    layer1_outputs(4407) <= a xor b;
    layer1_outputs(4408) <= not (a and b);
    layer1_outputs(4409) <= a and b;
    layer1_outputs(4410) <= 1'b1;
    layer1_outputs(4411) <= not (a or b);
    layer1_outputs(4412) <= a xor b;
    layer1_outputs(4413) <= a or b;
    layer1_outputs(4414) <= b;
    layer1_outputs(4415) <= not a or b;
    layer1_outputs(4416) <= a and not b;
    layer1_outputs(4417) <= not (a or b);
    layer1_outputs(4418) <= b;
    layer1_outputs(4419) <= not b or a;
    layer1_outputs(4420) <= b;
    layer1_outputs(4421) <= not b or a;
    layer1_outputs(4422) <= not a or b;
    layer1_outputs(4423) <= not a;
    layer1_outputs(4424) <= not a or b;
    layer1_outputs(4425) <= not a or b;
    layer1_outputs(4426) <= not b or a;
    layer1_outputs(4427) <= not a;
    layer1_outputs(4428) <= b;
    layer1_outputs(4429) <= not (a or b);
    layer1_outputs(4430) <= a or b;
    layer1_outputs(4431) <= a or b;
    layer1_outputs(4432) <= a and not b;
    layer1_outputs(4433) <= a and b;
    layer1_outputs(4434) <= not a;
    layer1_outputs(4435) <= b;
    layer1_outputs(4436) <= a or b;
    layer1_outputs(4437) <= not a or b;
    layer1_outputs(4438) <= not (a xor b);
    layer1_outputs(4439) <= 1'b0;
    layer1_outputs(4440) <= b and not a;
    layer1_outputs(4441) <= not b or a;
    layer1_outputs(4442) <= not (a xor b);
    layer1_outputs(4443) <= a or b;
    layer1_outputs(4444) <= a or b;
    layer1_outputs(4445) <= b and not a;
    layer1_outputs(4446) <= not a;
    layer1_outputs(4447) <= not (a or b);
    layer1_outputs(4448) <= b and not a;
    layer1_outputs(4449) <= not a;
    layer1_outputs(4450) <= b;
    layer1_outputs(4451) <= not a;
    layer1_outputs(4452) <= a and b;
    layer1_outputs(4453) <= not a or b;
    layer1_outputs(4454) <= not (a and b);
    layer1_outputs(4455) <= b;
    layer1_outputs(4456) <= not b or a;
    layer1_outputs(4457) <= a;
    layer1_outputs(4458) <= b and not a;
    layer1_outputs(4459) <= a and b;
    layer1_outputs(4460) <= not a;
    layer1_outputs(4461) <= a and not b;
    layer1_outputs(4462) <= not a or b;
    layer1_outputs(4463) <= a and b;
    layer1_outputs(4464) <= a xor b;
    layer1_outputs(4465) <= a;
    layer1_outputs(4466) <= not a;
    layer1_outputs(4467) <= not (a and b);
    layer1_outputs(4468) <= not (a and b);
    layer1_outputs(4469) <= b;
    layer1_outputs(4470) <= not (a or b);
    layer1_outputs(4471) <= not (a and b);
    layer1_outputs(4472) <= not a;
    layer1_outputs(4473) <= a;
    layer1_outputs(4474) <= a and b;
    layer1_outputs(4475) <= b and not a;
    layer1_outputs(4476) <= a xor b;
    layer1_outputs(4477) <= a and b;
    layer1_outputs(4478) <= not a or b;
    layer1_outputs(4479) <= b and not a;
    layer1_outputs(4480) <= not (a xor b);
    layer1_outputs(4481) <= not b or a;
    layer1_outputs(4482) <= a;
    layer1_outputs(4483) <= not b;
    layer1_outputs(4484) <= a and not b;
    layer1_outputs(4485) <= b;
    layer1_outputs(4486) <= a and not b;
    layer1_outputs(4487) <= a and not b;
    layer1_outputs(4488) <= not a or b;
    layer1_outputs(4489) <= not (a xor b);
    layer1_outputs(4490) <= not a;
    layer1_outputs(4491) <= not b or a;
    layer1_outputs(4492) <= a;
    layer1_outputs(4493) <= a and b;
    layer1_outputs(4494) <= a;
    layer1_outputs(4495) <= not b;
    layer1_outputs(4496) <= not b or a;
    layer1_outputs(4497) <= a and not b;
    layer1_outputs(4498) <= a xor b;
    layer1_outputs(4499) <= b;
    layer1_outputs(4500) <= not b or a;
    layer1_outputs(4501) <= a and not b;
    layer1_outputs(4502) <= a xor b;
    layer1_outputs(4503) <= a and not b;
    layer1_outputs(4504) <= a and b;
    layer1_outputs(4505) <= a and b;
    layer1_outputs(4506) <= b;
    layer1_outputs(4507) <= not a;
    layer1_outputs(4508) <= not (a xor b);
    layer1_outputs(4509) <= not b or a;
    layer1_outputs(4510) <= a xor b;
    layer1_outputs(4511) <= a and b;
    layer1_outputs(4512) <= a or b;
    layer1_outputs(4513) <= not (a or b);
    layer1_outputs(4514) <= not (a xor b);
    layer1_outputs(4515) <= 1'b1;
    layer1_outputs(4516) <= a xor b;
    layer1_outputs(4517) <= a and not b;
    layer1_outputs(4518) <= not (a xor b);
    layer1_outputs(4519) <= b and not a;
    layer1_outputs(4520) <= not (a or b);
    layer1_outputs(4521) <= a xor b;
    layer1_outputs(4522) <= a xor b;
    layer1_outputs(4523) <= a or b;
    layer1_outputs(4524) <= b;
    layer1_outputs(4525) <= a xor b;
    layer1_outputs(4526) <= b;
    layer1_outputs(4527) <= a or b;
    layer1_outputs(4528) <= a and b;
    layer1_outputs(4529) <= a xor b;
    layer1_outputs(4530) <= a and not b;
    layer1_outputs(4531) <= 1'b1;
    layer1_outputs(4532) <= not (a and b);
    layer1_outputs(4533) <= b;
    layer1_outputs(4534) <= not a or b;
    layer1_outputs(4535) <= b;
    layer1_outputs(4536) <= not a;
    layer1_outputs(4537) <= not a or b;
    layer1_outputs(4538) <= a xor b;
    layer1_outputs(4539) <= not (a xor b);
    layer1_outputs(4540) <= 1'b1;
    layer1_outputs(4541) <= not (a or b);
    layer1_outputs(4542) <= not a;
    layer1_outputs(4543) <= not (a xor b);
    layer1_outputs(4544) <= a and b;
    layer1_outputs(4545) <= not a;
    layer1_outputs(4546) <= not a;
    layer1_outputs(4547) <= not a;
    layer1_outputs(4548) <= a;
    layer1_outputs(4549) <= not a or b;
    layer1_outputs(4550) <= a;
    layer1_outputs(4551) <= 1'b0;
    layer1_outputs(4552) <= b;
    layer1_outputs(4553) <= not (a or b);
    layer1_outputs(4554) <= a;
    layer1_outputs(4555) <= not (a xor b);
    layer1_outputs(4556) <= not b or a;
    layer1_outputs(4557) <= not (a and b);
    layer1_outputs(4558) <= not (a or b);
    layer1_outputs(4559) <= not b or a;
    layer1_outputs(4560) <= a xor b;
    layer1_outputs(4561) <= a;
    layer1_outputs(4562) <= not a;
    layer1_outputs(4563) <= not a or b;
    layer1_outputs(4564) <= b and not a;
    layer1_outputs(4565) <= a or b;
    layer1_outputs(4566) <= 1'b1;
    layer1_outputs(4567) <= not a or b;
    layer1_outputs(4568) <= a and not b;
    layer1_outputs(4569) <= a xor b;
    layer1_outputs(4570) <= a and b;
    layer1_outputs(4571) <= a and b;
    layer1_outputs(4572) <= not b or a;
    layer1_outputs(4573) <= a xor b;
    layer1_outputs(4574) <= a xor b;
    layer1_outputs(4575) <= b;
    layer1_outputs(4576) <= b;
    layer1_outputs(4577) <= not a;
    layer1_outputs(4578) <= b;
    layer1_outputs(4579) <= not a;
    layer1_outputs(4580) <= b;
    layer1_outputs(4581) <= not a or b;
    layer1_outputs(4582) <= b;
    layer1_outputs(4583) <= not (a or b);
    layer1_outputs(4584) <= not (a and b);
    layer1_outputs(4585) <= a and not b;
    layer1_outputs(4586) <= a;
    layer1_outputs(4587) <= a and not b;
    layer1_outputs(4588) <= not (a xor b);
    layer1_outputs(4589) <= a;
    layer1_outputs(4590) <= not a or b;
    layer1_outputs(4591) <= a xor b;
    layer1_outputs(4592) <= a and not b;
    layer1_outputs(4593) <= a and b;
    layer1_outputs(4594) <= not (a or b);
    layer1_outputs(4595) <= b;
    layer1_outputs(4596) <= a and not b;
    layer1_outputs(4597) <= b and not a;
    layer1_outputs(4598) <= b and not a;
    layer1_outputs(4599) <= a or b;
    layer1_outputs(4600) <= a and not b;
    layer1_outputs(4601) <= b;
    layer1_outputs(4602) <= a or b;
    layer1_outputs(4603) <= b;
    layer1_outputs(4604) <= not (a or b);
    layer1_outputs(4605) <= a xor b;
    layer1_outputs(4606) <= a or b;
    layer1_outputs(4607) <= not a;
    layer1_outputs(4608) <= a xor b;
    layer1_outputs(4609) <= not b or a;
    layer1_outputs(4610) <= not (a xor b);
    layer1_outputs(4611) <= not b;
    layer1_outputs(4612) <= not b or a;
    layer1_outputs(4613) <= a and not b;
    layer1_outputs(4614) <= a or b;
    layer1_outputs(4615) <= not a;
    layer1_outputs(4616) <= a or b;
    layer1_outputs(4617) <= not (a or b);
    layer1_outputs(4618) <= not b;
    layer1_outputs(4619) <= not (a or b);
    layer1_outputs(4620) <= a and not b;
    layer1_outputs(4621) <= not b;
    layer1_outputs(4622) <= 1'b0;
    layer1_outputs(4623) <= not a or b;
    layer1_outputs(4624) <= not (a xor b);
    layer1_outputs(4625) <= b;
    layer1_outputs(4626) <= a;
    layer1_outputs(4627) <= not a;
    layer1_outputs(4628) <= a or b;
    layer1_outputs(4629) <= not b or a;
    layer1_outputs(4630) <= not a;
    layer1_outputs(4631) <= a;
    layer1_outputs(4632) <= b;
    layer1_outputs(4633) <= b;
    layer1_outputs(4634) <= not b;
    layer1_outputs(4635) <= not (a or b);
    layer1_outputs(4636) <= b;
    layer1_outputs(4637) <= not (a or b);
    layer1_outputs(4638) <= not a or b;
    layer1_outputs(4639) <= not (a or b);
    layer1_outputs(4640) <= b;
    layer1_outputs(4641) <= a and b;
    layer1_outputs(4642) <= not a or b;
    layer1_outputs(4643) <= a;
    layer1_outputs(4644) <= not (a xor b);
    layer1_outputs(4645) <= a or b;
    layer1_outputs(4646) <= 1'b1;
    layer1_outputs(4647) <= a;
    layer1_outputs(4648) <= a and not b;
    layer1_outputs(4649) <= a xor b;
    layer1_outputs(4650) <= a or b;
    layer1_outputs(4651) <= not a or b;
    layer1_outputs(4652) <= not (a and b);
    layer1_outputs(4653) <= not (a and b);
    layer1_outputs(4654) <= not (a xor b);
    layer1_outputs(4655) <= not b or a;
    layer1_outputs(4656) <= a or b;
    layer1_outputs(4657) <= a xor b;
    layer1_outputs(4658) <= not a;
    layer1_outputs(4659) <= not a or b;
    layer1_outputs(4660) <= not b;
    layer1_outputs(4661) <= a or b;
    layer1_outputs(4662) <= not (a or b);
    layer1_outputs(4663) <= not b or a;
    layer1_outputs(4664) <= a xor b;
    layer1_outputs(4665) <= a and not b;
    layer1_outputs(4666) <= not (a and b);
    layer1_outputs(4667) <= not a or b;
    layer1_outputs(4668) <= not a;
    layer1_outputs(4669) <= not b;
    layer1_outputs(4670) <= b;
    layer1_outputs(4671) <= a or b;
    layer1_outputs(4672) <= not (a and b);
    layer1_outputs(4673) <= b and not a;
    layer1_outputs(4674) <= a and b;
    layer1_outputs(4675) <= not a;
    layer1_outputs(4676) <= not a;
    layer1_outputs(4677) <= not a or b;
    layer1_outputs(4678) <= not a;
    layer1_outputs(4679) <= not b or a;
    layer1_outputs(4680) <= not a;
    layer1_outputs(4681) <= a or b;
    layer1_outputs(4682) <= b and not a;
    layer1_outputs(4683) <= 1'b0;
    layer1_outputs(4684) <= not (a or b);
    layer1_outputs(4685) <= not b or a;
    layer1_outputs(4686) <= not a;
    layer1_outputs(4687) <= a;
    layer1_outputs(4688) <= not a;
    layer1_outputs(4689) <= not b or a;
    layer1_outputs(4690) <= a;
    layer1_outputs(4691) <= not (a and b);
    layer1_outputs(4692) <= a xor b;
    layer1_outputs(4693) <= not a;
    layer1_outputs(4694) <= b;
    layer1_outputs(4695) <= a and not b;
    layer1_outputs(4696) <= not (a or b);
    layer1_outputs(4697) <= not (a xor b);
    layer1_outputs(4698) <= not (a and b);
    layer1_outputs(4699) <= 1'b1;
    layer1_outputs(4700) <= a;
    layer1_outputs(4701) <= not (a and b);
    layer1_outputs(4702) <= a and not b;
    layer1_outputs(4703) <= not b or a;
    layer1_outputs(4704) <= not (a xor b);
    layer1_outputs(4705) <= not b or a;
    layer1_outputs(4706) <= a or b;
    layer1_outputs(4707) <= not b;
    layer1_outputs(4708) <= a xor b;
    layer1_outputs(4709) <= a and b;
    layer1_outputs(4710) <= a and b;
    layer1_outputs(4711) <= not (a xor b);
    layer1_outputs(4712) <= not b;
    layer1_outputs(4713) <= not b or a;
    layer1_outputs(4714) <= not b or a;
    layer1_outputs(4715) <= not a;
    layer1_outputs(4716) <= a or b;
    layer1_outputs(4717) <= not (a xor b);
    layer1_outputs(4718) <= a and not b;
    layer1_outputs(4719) <= b;
    layer1_outputs(4720) <= 1'b0;
    layer1_outputs(4721) <= not (a or b);
    layer1_outputs(4722) <= a xor b;
    layer1_outputs(4723) <= a and b;
    layer1_outputs(4724) <= b;
    layer1_outputs(4725) <= b and not a;
    layer1_outputs(4726) <= a and b;
    layer1_outputs(4727) <= b and not a;
    layer1_outputs(4728) <= not a or b;
    layer1_outputs(4729) <= b;
    layer1_outputs(4730) <= not (a or b);
    layer1_outputs(4731) <= not a;
    layer1_outputs(4732) <= b and not a;
    layer1_outputs(4733) <= not b or a;
    layer1_outputs(4734) <= not b;
    layer1_outputs(4735) <= not (a or b);
    layer1_outputs(4736) <= not b;
    layer1_outputs(4737) <= a and not b;
    layer1_outputs(4738) <= not (a and b);
    layer1_outputs(4739) <= not a;
    layer1_outputs(4740) <= b;
    layer1_outputs(4741) <= not b or a;
    layer1_outputs(4742) <= not b;
    layer1_outputs(4743) <= a and b;
    layer1_outputs(4744) <= a;
    layer1_outputs(4745) <= a and not b;
    layer1_outputs(4746) <= not (a and b);
    layer1_outputs(4747) <= b and not a;
    layer1_outputs(4748) <= b and not a;
    layer1_outputs(4749) <= not b or a;
    layer1_outputs(4750) <= not b;
    layer1_outputs(4751) <= a;
    layer1_outputs(4752) <= not b;
    layer1_outputs(4753) <= a and b;
    layer1_outputs(4754) <= b;
    layer1_outputs(4755) <= a;
    layer1_outputs(4756) <= not (a and b);
    layer1_outputs(4757) <= b;
    layer1_outputs(4758) <= not (a and b);
    layer1_outputs(4759) <= not a or b;
    layer1_outputs(4760) <= a xor b;
    layer1_outputs(4761) <= a;
    layer1_outputs(4762) <= b;
    layer1_outputs(4763) <= a and not b;
    layer1_outputs(4764) <= a;
    layer1_outputs(4765) <= not b;
    layer1_outputs(4766) <= a;
    layer1_outputs(4767) <= not b or a;
    layer1_outputs(4768) <= not (a xor b);
    layer1_outputs(4769) <= not a;
    layer1_outputs(4770) <= a and b;
    layer1_outputs(4771) <= not (a or b);
    layer1_outputs(4772) <= not (a xor b);
    layer1_outputs(4773) <= not a;
    layer1_outputs(4774) <= not a;
    layer1_outputs(4775) <= not (a xor b);
    layer1_outputs(4776) <= a and b;
    layer1_outputs(4777) <= not (a or b);
    layer1_outputs(4778) <= not b or a;
    layer1_outputs(4779) <= a or b;
    layer1_outputs(4780) <= a or b;
    layer1_outputs(4781) <= not (a and b);
    layer1_outputs(4782) <= not (a xor b);
    layer1_outputs(4783) <= a or b;
    layer1_outputs(4784) <= a or b;
    layer1_outputs(4785) <= a xor b;
    layer1_outputs(4786) <= not a;
    layer1_outputs(4787) <= a;
    layer1_outputs(4788) <= b and not a;
    layer1_outputs(4789) <= a;
    layer1_outputs(4790) <= not a;
    layer1_outputs(4791) <= not (a xor b);
    layer1_outputs(4792) <= not b or a;
    layer1_outputs(4793) <= a and b;
    layer1_outputs(4794) <= a and not b;
    layer1_outputs(4795) <= not (a or b);
    layer1_outputs(4796) <= not b or a;
    layer1_outputs(4797) <= not a;
    layer1_outputs(4798) <= not b;
    layer1_outputs(4799) <= not a;
    layer1_outputs(4800) <= not (a xor b);
    layer1_outputs(4801) <= not a;
    layer1_outputs(4802) <= not (a xor b);
    layer1_outputs(4803) <= not b;
    layer1_outputs(4804) <= not (a or b);
    layer1_outputs(4805) <= b;
    layer1_outputs(4806) <= b;
    layer1_outputs(4807) <= a and not b;
    layer1_outputs(4808) <= not (a xor b);
    layer1_outputs(4809) <= a xor b;
    layer1_outputs(4810) <= b and not a;
    layer1_outputs(4811) <= not a;
    layer1_outputs(4812) <= not b;
    layer1_outputs(4813) <= not (a xor b);
    layer1_outputs(4814) <= a xor b;
    layer1_outputs(4815) <= not b;
    layer1_outputs(4816) <= b;
    layer1_outputs(4817) <= not b;
    layer1_outputs(4818) <= a and b;
    layer1_outputs(4819) <= a;
    layer1_outputs(4820) <= not b or a;
    layer1_outputs(4821) <= not a or b;
    layer1_outputs(4822) <= a or b;
    layer1_outputs(4823) <= not (a and b);
    layer1_outputs(4824) <= b;
    layer1_outputs(4825) <= not b or a;
    layer1_outputs(4826) <= not b;
    layer1_outputs(4827) <= a or b;
    layer1_outputs(4828) <= not b or a;
    layer1_outputs(4829) <= a and not b;
    layer1_outputs(4830) <= a and b;
    layer1_outputs(4831) <= not (a xor b);
    layer1_outputs(4832) <= not (a and b);
    layer1_outputs(4833) <= not a;
    layer1_outputs(4834) <= a xor b;
    layer1_outputs(4835) <= not (a or b);
    layer1_outputs(4836) <= b and not a;
    layer1_outputs(4837) <= not (a or b);
    layer1_outputs(4838) <= not b or a;
    layer1_outputs(4839) <= not b;
    layer1_outputs(4840) <= not a;
    layer1_outputs(4841) <= not (a or b);
    layer1_outputs(4842) <= b and not a;
    layer1_outputs(4843) <= not a;
    layer1_outputs(4844) <= not a;
    layer1_outputs(4845) <= b and not a;
    layer1_outputs(4846) <= not (a or b);
    layer1_outputs(4847) <= not b;
    layer1_outputs(4848) <= a and not b;
    layer1_outputs(4849) <= not (a xor b);
    layer1_outputs(4850) <= not (a or b);
    layer1_outputs(4851) <= a and b;
    layer1_outputs(4852) <= b;
    layer1_outputs(4853) <= not b;
    layer1_outputs(4854) <= not b;
    layer1_outputs(4855) <= a xor b;
    layer1_outputs(4856) <= not (a or b);
    layer1_outputs(4857) <= not b or a;
    layer1_outputs(4858) <= not b;
    layer1_outputs(4859) <= not (a or b);
    layer1_outputs(4860) <= a or b;
    layer1_outputs(4861) <= a;
    layer1_outputs(4862) <= not a or b;
    layer1_outputs(4863) <= a xor b;
    layer1_outputs(4864) <= a or b;
    layer1_outputs(4865) <= a;
    layer1_outputs(4866) <= not (a or b);
    layer1_outputs(4867) <= a xor b;
    layer1_outputs(4868) <= a and b;
    layer1_outputs(4869) <= not b;
    layer1_outputs(4870) <= a xor b;
    layer1_outputs(4871) <= not b;
    layer1_outputs(4872) <= not (a xor b);
    layer1_outputs(4873) <= not (a xor b);
    layer1_outputs(4874) <= not a;
    layer1_outputs(4875) <= 1'b0;
    layer1_outputs(4876) <= not (a and b);
    layer1_outputs(4877) <= not (a and b);
    layer1_outputs(4878) <= b and not a;
    layer1_outputs(4879) <= not b or a;
    layer1_outputs(4880) <= not b or a;
    layer1_outputs(4881) <= b;
    layer1_outputs(4882) <= not b;
    layer1_outputs(4883) <= not b;
    layer1_outputs(4884) <= not b;
    layer1_outputs(4885) <= a xor b;
    layer1_outputs(4886) <= not a or b;
    layer1_outputs(4887) <= not a;
    layer1_outputs(4888) <= b;
    layer1_outputs(4889) <= not (a xor b);
    layer1_outputs(4890) <= not b or a;
    layer1_outputs(4891) <= a and b;
    layer1_outputs(4892) <= b and not a;
    layer1_outputs(4893) <= not (a and b);
    layer1_outputs(4894) <= a and b;
    layer1_outputs(4895) <= a or b;
    layer1_outputs(4896) <= a or b;
    layer1_outputs(4897) <= b;
    layer1_outputs(4898) <= a xor b;
    layer1_outputs(4899) <= not (a or b);
    layer1_outputs(4900) <= b;
    layer1_outputs(4901) <= not b;
    layer1_outputs(4902) <= b;
    layer1_outputs(4903) <= a xor b;
    layer1_outputs(4904) <= a and not b;
    layer1_outputs(4905) <= not b or a;
    layer1_outputs(4906) <= a or b;
    layer1_outputs(4907) <= a and b;
    layer1_outputs(4908) <= a xor b;
    layer1_outputs(4909) <= not a;
    layer1_outputs(4910) <= a;
    layer1_outputs(4911) <= not (a and b);
    layer1_outputs(4912) <= not a;
    layer1_outputs(4913) <= not (a or b);
    layer1_outputs(4914) <= a;
    layer1_outputs(4915) <= a and not b;
    layer1_outputs(4916) <= a or b;
    layer1_outputs(4917) <= b;
    layer1_outputs(4918) <= b and not a;
    layer1_outputs(4919) <= 1'b1;
    layer1_outputs(4920) <= a and not b;
    layer1_outputs(4921) <= not a;
    layer1_outputs(4922) <= b and not a;
    layer1_outputs(4923) <= not a;
    layer1_outputs(4924) <= not b or a;
    layer1_outputs(4925) <= b;
    layer1_outputs(4926) <= a;
    layer1_outputs(4927) <= not (a or b);
    layer1_outputs(4928) <= a or b;
    layer1_outputs(4929) <= not a;
    layer1_outputs(4930) <= a and b;
    layer1_outputs(4931) <= a or b;
    layer1_outputs(4932) <= a;
    layer1_outputs(4933) <= a;
    layer1_outputs(4934) <= b;
    layer1_outputs(4935) <= not (a xor b);
    layer1_outputs(4936) <= a and not b;
    layer1_outputs(4937) <= a xor b;
    layer1_outputs(4938) <= b;
    layer1_outputs(4939) <= a or b;
    layer1_outputs(4940) <= not (a and b);
    layer1_outputs(4941) <= not (a and b);
    layer1_outputs(4942) <= not (a or b);
    layer1_outputs(4943) <= not b;
    layer1_outputs(4944) <= a xor b;
    layer1_outputs(4945) <= a;
    layer1_outputs(4946) <= b;
    layer1_outputs(4947) <= not a;
    layer1_outputs(4948) <= b;
    layer1_outputs(4949) <= a and b;
    layer1_outputs(4950) <= not (a or b);
    layer1_outputs(4951) <= not (a xor b);
    layer1_outputs(4952) <= not (a or b);
    layer1_outputs(4953) <= a xor b;
    layer1_outputs(4954) <= a and b;
    layer1_outputs(4955) <= not b or a;
    layer1_outputs(4956) <= not b;
    layer1_outputs(4957) <= b;
    layer1_outputs(4958) <= not a;
    layer1_outputs(4959) <= b;
    layer1_outputs(4960) <= a;
    layer1_outputs(4961) <= not (a or b);
    layer1_outputs(4962) <= not a or b;
    layer1_outputs(4963) <= not b;
    layer1_outputs(4964) <= a and not b;
    layer1_outputs(4965) <= not (a or b);
    layer1_outputs(4966) <= not b;
    layer1_outputs(4967) <= b and not a;
    layer1_outputs(4968) <= not (a or b);
    layer1_outputs(4969) <= not (a xor b);
    layer1_outputs(4970) <= a or b;
    layer1_outputs(4971) <= not (a or b);
    layer1_outputs(4972) <= not (a xor b);
    layer1_outputs(4973) <= b;
    layer1_outputs(4974) <= a and b;
    layer1_outputs(4975) <= a xor b;
    layer1_outputs(4976) <= b and not a;
    layer1_outputs(4977) <= not b;
    layer1_outputs(4978) <= not b;
    layer1_outputs(4979) <= not (a and b);
    layer1_outputs(4980) <= a;
    layer1_outputs(4981) <= a and b;
    layer1_outputs(4982) <= a;
    layer1_outputs(4983) <= a or b;
    layer1_outputs(4984) <= a xor b;
    layer1_outputs(4985) <= not b or a;
    layer1_outputs(4986) <= a or b;
    layer1_outputs(4987) <= not b;
    layer1_outputs(4988) <= a and not b;
    layer1_outputs(4989) <= a and b;
    layer1_outputs(4990) <= not (a and b);
    layer1_outputs(4991) <= not a or b;
    layer1_outputs(4992) <= b and not a;
    layer1_outputs(4993) <= not b;
    layer1_outputs(4994) <= b;
    layer1_outputs(4995) <= not a;
    layer1_outputs(4996) <= b and not a;
    layer1_outputs(4997) <= not b or a;
    layer1_outputs(4998) <= not b;
    layer1_outputs(4999) <= a and b;
    layer1_outputs(5000) <= a and b;
    layer1_outputs(5001) <= not b;
    layer1_outputs(5002) <= not (a xor b);
    layer1_outputs(5003) <= a and not b;
    layer1_outputs(5004) <= not a or b;
    layer1_outputs(5005) <= b;
    layer1_outputs(5006) <= 1'b1;
    layer1_outputs(5007) <= not (a xor b);
    layer1_outputs(5008) <= not (a or b);
    layer1_outputs(5009) <= a or b;
    layer1_outputs(5010) <= a xor b;
    layer1_outputs(5011) <= not (a or b);
    layer1_outputs(5012) <= not a;
    layer1_outputs(5013) <= a and b;
    layer1_outputs(5014) <= not (a and b);
    layer1_outputs(5015) <= not (a and b);
    layer1_outputs(5016) <= a;
    layer1_outputs(5017) <= a;
    layer1_outputs(5018) <= b and not a;
    layer1_outputs(5019) <= not b or a;
    layer1_outputs(5020) <= not (a xor b);
    layer1_outputs(5021) <= not (a and b);
    layer1_outputs(5022) <= not (a and b);
    layer1_outputs(5023) <= not (a xor b);
    layer1_outputs(5024) <= not b or a;
    layer1_outputs(5025) <= not b or a;
    layer1_outputs(5026) <= b;
    layer1_outputs(5027) <= a and b;
    layer1_outputs(5028) <= not b;
    layer1_outputs(5029) <= not (a xor b);
    layer1_outputs(5030) <= a and not b;
    layer1_outputs(5031) <= not b or a;
    layer1_outputs(5032) <= a xor b;
    layer1_outputs(5033) <= not (a or b);
    layer1_outputs(5034) <= not b;
    layer1_outputs(5035) <= not a or b;
    layer1_outputs(5036) <= a or b;
    layer1_outputs(5037) <= not a or b;
    layer1_outputs(5038) <= not b;
    layer1_outputs(5039) <= not (a and b);
    layer1_outputs(5040) <= not (a xor b);
    layer1_outputs(5041) <= b and not a;
    layer1_outputs(5042) <= a xor b;
    layer1_outputs(5043) <= not b;
    layer1_outputs(5044) <= not a or b;
    layer1_outputs(5045) <= a or b;
    layer1_outputs(5046) <= not a;
    layer1_outputs(5047) <= not a;
    layer1_outputs(5048) <= a and b;
    layer1_outputs(5049) <= a or b;
    layer1_outputs(5050) <= 1'b0;
    layer1_outputs(5051) <= not a;
    layer1_outputs(5052) <= b;
    layer1_outputs(5053) <= not b or a;
    layer1_outputs(5054) <= not (a and b);
    layer1_outputs(5055) <= not (a or b);
    layer1_outputs(5056) <= not b;
    layer1_outputs(5057) <= not a;
    layer1_outputs(5058) <= not a;
    layer1_outputs(5059) <= a;
    layer1_outputs(5060) <= a and b;
    layer1_outputs(5061) <= b;
    layer1_outputs(5062) <= not a or b;
    layer1_outputs(5063) <= not (a or b);
    layer1_outputs(5064) <= 1'b1;
    layer1_outputs(5065) <= not a;
    layer1_outputs(5066) <= a and not b;
    layer1_outputs(5067) <= not b;
    layer1_outputs(5068) <= not b or a;
    layer1_outputs(5069) <= not a or b;
    layer1_outputs(5070) <= a;
    layer1_outputs(5071) <= not (a and b);
    layer1_outputs(5072) <= b and not a;
    layer1_outputs(5073) <= a and b;
    layer1_outputs(5074) <= not a or b;
    layer1_outputs(5075) <= not b;
    layer1_outputs(5076) <= not b or a;
    layer1_outputs(5077) <= not a;
    layer1_outputs(5078) <= not a;
    layer1_outputs(5079) <= b;
    layer1_outputs(5080) <= not b or a;
    layer1_outputs(5081) <= a xor b;
    layer1_outputs(5082) <= not a;
    layer1_outputs(5083) <= not (a and b);
    layer1_outputs(5084) <= not (a and b);
    layer1_outputs(5085) <= a and b;
    layer1_outputs(5086) <= not a or b;
    layer1_outputs(5087) <= not b;
    layer1_outputs(5088) <= a;
    layer1_outputs(5089) <= a xor b;
    layer1_outputs(5090) <= not b or a;
    layer1_outputs(5091) <= not (a and b);
    layer1_outputs(5092) <= b and not a;
    layer1_outputs(5093) <= a or b;
    layer1_outputs(5094) <= b;
    layer1_outputs(5095) <= not (a or b);
    layer1_outputs(5096) <= b;
    layer1_outputs(5097) <= not (a or b);
    layer1_outputs(5098) <= not (a xor b);
    layer1_outputs(5099) <= not (a xor b);
    layer1_outputs(5100) <= not a;
    layer1_outputs(5101) <= not (a xor b);
    layer1_outputs(5102) <= not b;
    layer1_outputs(5103) <= b and not a;
    layer1_outputs(5104) <= not a or b;
    layer1_outputs(5105) <= not b;
    layer1_outputs(5106) <= 1'b1;
    layer1_outputs(5107) <= a;
    layer1_outputs(5108) <= not a;
    layer1_outputs(5109) <= a;
    layer1_outputs(5110) <= a and not b;
    layer1_outputs(5111) <= not b;
    layer1_outputs(5112) <= a;
    layer1_outputs(5113) <= not (a or b);
    layer1_outputs(5114) <= b;
    layer1_outputs(5115) <= not b or a;
    layer1_outputs(5116) <= a or b;
    layer1_outputs(5117) <= not (a xor b);
    layer1_outputs(5118) <= a;
    layer1_outputs(5119) <= a or b;
    layer2_outputs(0) <= not (a and b);
    layer2_outputs(1) <= not (a xor b);
    layer2_outputs(2) <= a and not b;
    layer2_outputs(3) <= a and not b;
    layer2_outputs(4) <= not a or b;
    layer2_outputs(5) <= not (a and b);
    layer2_outputs(6) <= 1'b0;
    layer2_outputs(7) <= a and b;
    layer2_outputs(8) <= not a;
    layer2_outputs(9) <= not a;
    layer2_outputs(10) <= a;
    layer2_outputs(11) <= a;
    layer2_outputs(12) <= not (a and b);
    layer2_outputs(13) <= b;
    layer2_outputs(14) <= b;
    layer2_outputs(15) <= not (a xor b);
    layer2_outputs(16) <= not (a and b);
    layer2_outputs(17) <= a;
    layer2_outputs(18) <= a and not b;
    layer2_outputs(19) <= 1'b1;
    layer2_outputs(20) <= a xor b;
    layer2_outputs(21) <= not (a or b);
    layer2_outputs(22) <= a and b;
    layer2_outputs(23) <= not b;
    layer2_outputs(24) <= a xor b;
    layer2_outputs(25) <= a and not b;
    layer2_outputs(26) <= not a or b;
    layer2_outputs(27) <= a;
    layer2_outputs(28) <= not (a or b);
    layer2_outputs(29) <= a;
    layer2_outputs(30) <= not b;
    layer2_outputs(31) <= not b;
    layer2_outputs(32) <= a;
    layer2_outputs(33) <= not a or b;
    layer2_outputs(34) <= not (a and b);
    layer2_outputs(35) <= not a or b;
    layer2_outputs(36) <= not b;
    layer2_outputs(37) <= a or b;
    layer2_outputs(38) <= b and not a;
    layer2_outputs(39) <= not (a and b);
    layer2_outputs(40) <= b;
    layer2_outputs(41) <= a or b;
    layer2_outputs(42) <= a;
    layer2_outputs(43) <= 1'b0;
    layer2_outputs(44) <= not a;
    layer2_outputs(45) <= b;
    layer2_outputs(46) <= a xor b;
    layer2_outputs(47) <= a;
    layer2_outputs(48) <= a and not b;
    layer2_outputs(49) <= not b or a;
    layer2_outputs(50) <= not (a or b);
    layer2_outputs(51) <= not a or b;
    layer2_outputs(52) <= b;
    layer2_outputs(53) <= a or b;
    layer2_outputs(54) <= a and not b;
    layer2_outputs(55) <= not (a and b);
    layer2_outputs(56) <= a;
    layer2_outputs(57) <= not a;
    layer2_outputs(58) <= not b;
    layer2_outputs(59) <= not (a or b);
    layer2_outputs(60) <= a or b;
    layer2_outputs(61) <= not a;
    layer2_outputs(62) <= b;
    layer2_outputs(63) <= not (a and b);
    layer2_outputs(64) <= not (a xor b);
    layer2_outputs(65) <= a and not b;
    layer2_outputs(66) <= not b;
    layer2_outputs(67) <= not (a or b);
    layer2_outputs(68) <= b;
    layer2_outputs(69) <= a;
    layer2_outputs(70) <= a xor b;
    layer2_outputs(71) <= a xor b;
    layer2_outputs(72) <= a;
    layer2_outputs(73) <= not b;
    layer2_outputs(74) <= not (a or b);
    layer2_outputs(75) <= not a;
    layer2_outputs(76) <= b and not a;
    layer2_outputs(77) <= a;
    layer2_outputs(78) <= not (a and b);
    layer2_outputs(79) <= a xor b;
    layer2_outputs(80) <= a or b;
    layer2_outputs(81) <= not b or a;
    layer2_outputs(82) <= b and not a;
    layer2_outputs(83) <= b;
    layer2_outputs(84) <= not (a and b);
    layer2_outputs(85) <= a and not b;
    layer2_outputs(86) <= a and not b;
    layer2_outputs(87) <= not a;
    layer2_outputs(88) <= b;
    layer2_outputs(89) <= not b;
    layer2_outputs(90) <= a and b;
    layer2_outputs(91) <= a and not b;
    layer2_outputs(92) <= a and b;
    layer2_outputs(93) <= a;
    layer2_outputs(94) <= not (a or b);
    layer2_outputs(95) <= not a or b;
    layer2_outputs(96) <= not a or b;
    layer2_outputs(97) <= not b or a;
    layer2_outputs(98) <= a xor b;
    layer2_outputs(99) <= a;
    layer2_outputs(100) <= not b;
    layer2_outputs(101) <= a and b;
    layer2_outputs(102) <= a and not b;
    layer2_outputs(103) <= not a;
    layer2_outputs(104) <= a xor b;
    layer2_outputs(105) <= not b;
    layer2_outputs(106) <= not b;
    layer2_outputs(107) <= not a;
    layer2_outputs(108) <= a or b;
    layer2_outputs(109) <= not b or a;
    layer2_outputs(110) <= not b or a;
    layer2_outputs(111) <= not (a xor b);
    layer2_outputs(112) <= not a or b;
    layer2_outputs(113) <= a;
    layer2_outputs(114) <= not (a xor b);
    layer2_outputs(115) <= a;
    layer2_outputs(116) <= a or b;
    layer2_outputs(117) <= a and not b;
    layer2_outputs(118) <= not b;
    layer2_outputs(119) <= b and not a;
    layer2_outputs(120) <= a and b;
    layer2_outputs(121) <= not (a and b);
    layer2_outputs(122) <= not b or a;
    layer2_outputs(123) <= a;
    layer2_outputs(124) <= not (a and b);
    layer2_outputs(125) <= not b;
    layer2_outputs(126) <= not (a and b);
    layer2_outputs(127) <= not (a or b);
    layer2_outputs(128) <= a or b;
    layer2_outputs(129) <= b;
    layer2_outputs(130) <= not (a xor b);
    layer2_outputs(131) <= not (a xor b);
    layer2_outputs(132) <= not (a or b);
    layer2_outputs(133) <= b;
    layer2_outputs(134) <= not (a and b);
    layer2_outputs(135) <= a;
    layer2_outputs(136) <= a and not b;
    layer2_outputs(137) <= a;
    layer2_outputs(138) <= not (a or b);
    layer2_outputs(139) <= a and not b;
    layer2_outputs(140) <= not b;
    layer2_outputs(141) <= not a or b;
    layer2_outputs(142) <= a;
    layer2_outputs(143) <= not a or b;
    layer2_outputs(144) <= b and not a;
    layer2_outputs(145) <= not (a xor b);
    layer2_outputs(146) <= a;
    layer2_outputs(147) <= not a or b;
    layer2_outputs(148) <= a xor b;
    layer2_outputs(149) <= a or b;
    layer2_outputs(150) <= not a;
    layer2_outputs(151) <= not (a and b);
    layer2_outputs(152) <= a xor b;
    layer2_outputs(153) <= not b or a;
    layer2_outputs(154) <= not b;
    layer2_outputs(155) <= b;
    layer2_outputs(156) <= a and b;
    layer2_outputs(157) <= a;
    layer2_outputs(158) <= a and b;
    layer2_outputs(159) <= a and not b;
    layer2_outputs(160) <= not a;
    layer2_outputs(161) <= b;
    layer2_outputs(162) <= not b;
    layer2_outputs(163) <= a or b;
    layer2_outputs(164) <= b;
    layer2_outputs(165) <= not (a and b);
    layer2_outputs(166) <= b and not a;
    layer2_outputs(167) <= not b or a;
    layer2_outputs(168) <= a or b;
    layer2_outputs(169) <= b and not a;
    layer2_outputs(170) <= not b or a;
    layer2_outputs(171) <= not a;
    layer2_outputs(172) <= not (a and b);
    layer2_outputs(173) <= not (a xor b);
    layer2_outputs(174) <= a and not b;
    layer2_outputs(175) <= not (a and b);
    layer2_outputs(176) <= a xor b;
    layer2_outputs(177) <= not b;
    layer2_outputs(178) <= b and not a;
    layer2_outputs(179) <= a xor b;
    layer2_outputs(180) <= b;
    layer2_outputs(181) <= not a;
    layer2_outputs(182) <= a;
    layer2_outputs(183) <= not b;
    layer2_outputs(184) <= a;
    layer2_outputs(185) <= a or b;
    layer2_outputs(186) <= not a;
    layer2_outputs(187) <= not a;
    layer2_outputs(188) <= b and not a;
    layer2_outputs(189) <= a and b;
    layer2_outputs(190) <= not (a or b);
    layer2_outputs(191) <= not b or a;
    layer2_outputs(192) <= b and not a;
    layer2_outputs(193) <= b and not a;
    layer2_outputs(194) <= a and b;
    layer2_outputs(195) <= not (a xor b);
    layer2_outputs(196) <= not (a or b);
    layer2_outputs(197) <= a and not b;
    layer2_outputs(198) <= a or b;
    layer2_outputs(199) <= a and b;
    layer2_outputs(200) <= b;
    layer2_outputs(201) <= not (a and b);
    layer2_outputs(202) <= b and not a;
    layer2_outputs(203) <= a;
    layer2_outputs(204) <= b and not a;
    layer2_outputs(205) <= not a or b;
    layer2_outputs(206) <= not (a and b);
    layer2_outputs(207) <= not a;
    layer2_outputs(208) <= not a;
    layer2_outputs(209) <= b and not a;
    layer2_outputs(210) <= a;
    layer2_outputs(211) <= a or b;
    layer2_outputs(212) <= b;
    layer2_outputs(213) <= not a or b;
    layer2_outputs(214) <= not b or a;
    layer2_outputs(215) <= a and not b;
    layer2_outputs(216) <= b;
    layer2_outputs(217) <= not b or a;
    layer2_outputs(218) <= a and b;
    layer2_outputs(219) <= not (a or b);
    layer2_outputs(220) <= not b;
    layer2_outputs(221) <= a and not b;
    layer2_outputs(222) <= b and not a;
    layer2_outputs(223) <= a or b;
    layer2_outputs(224) <= a and not b;
    layer2_outputs(225) <= a and b;
    layer2_outputs(226) <= not a;
    layer2_outputs(227) <= a or b;
    layer2_outputs(228) <= b;
    layer2_outputs(229) <= not (a and b);
    layer2_outputs(230) <= not (a xor b);
    layer2_outputs(231) <= b and not a;
    layer2_outputs(232) <= not a;
    layer2_outputs(233) <= not a or b;
    layer2_outputs(234) <= not (a or b);
    layer2_outputs(235) <= a xor b;
    layer2_outputs(236) <= 1'b0;
    layer2_outputs(237) <= not (a and b);
    layer2_outputs(238) <= not a or b;
    layer2_outputs(239) <= a xor b;
    layer2_outputs(240) <= b and not a;
    layer2_outputs(241) <= a and b;
    layer2_outputs(242) <= a;
    layer2_outputs(243) <= a;
    layer2_outputs(244) <= a or b;
    layer2_outputs(245) <= not a;
    layer2_outputs(246) <= a;
    layer2_outputs(247) <= a;
    layer2_outputs(248) <= b;
    layer2_outputs(249) <= not (a or b);
    layer2_outputs(250) <= a;
    layer2_outputs(251) <= not (a xor b);
    layer2_outputs(252) <= a;
    layer2_outputs(253) <= a xor b;
    layer2_outputs(254) <= a;
    layer2_outputs(255) <= not (a and b);
    layer2_outputs(256) <= b;
    layer2_outputs(257) <= not (a and b);
    layer2_outputs(258) <= not (a xor b);
    layer2_outputs(259) <= a xor b;
    layer2_outputs(260) <= a and not b;
    layer2_outputs(261) <= not b or a;
    layer2_outputs(262) <= 1'b1;
    layer2_outputs(263) <= not a;
    layer2_outputs(264) <= a;
    layer2_outputs(265) <= a or b;
    layer2_outputs(266) <= a and not b;
    layer2_outputs(267) <= not b;
    layer2_outputs(268) <= not a;
    layer2_outputs(269) <= b;
    layer2_outputs(270) <= not (a or b);
    layer2_outputs(271) <= b and not a;
    layer2_outputs(272) <= not b;
    layer2_outputs(273) <= not (a or b);
    layer2_outputs(274) <= a and b;
    layer2_outputs(275) <= not b or a;
    layer2_outputs(276) <= a xor b;
    layer2_outputs(277) <= a;
    layer2_outputs(278) <= not a;
    layer2_outputs(279) <= not a or b;
    layer2_outputs(280) <= a;
    layer2_outputs(281) <= b;
    layer2_outputs(282) <= not b;
    layer2_outputs(283) <= not (a xor b);
    layer2_outputs(284) <= not a or b;
    layer2_outputs(285) <= not a;
    layer2_outputs(286) <= not b;
    layer2_outputs(287) <= a;
    layer2_outputs(288) <= a xor b;
    layer2_outputs(289) <= a;
    layer2_outputs(290) <= not b;
    layer2_outputs(291) <= not b;
    layer2_outputs(292) <= a or b;
    layer2_outputs(293) <= not a or b;
    layer2_outputs(294) <= not a or b;
    layer2_outputs(295) <= a;
    layer2_outputs(296) <= a and b;
    layer2_outputs(297) <= not a or b;
    layer2_outputs(298) <= not b or a;
    layer2_outputs(299) <= not b;
    layer2_outputs(300) <= a or b;
    layer2_outputs(301) <= not b;
    layer2_outputs(302) <= a;
    layer2_outputs(303) <= b;
    layer2_outputs(304) <= b;
    layer2_outputs(305) <= a and not b;
    layer2_outputs(306) <= not (a or b);
    layer2_outputs(307) <= not b;
    layer2_outputs(308) <= not a;
    layer2_outputs(309) <= not (a and b);
    layer2_outputs(310) <= b and not a;
    layer2_outputs(311) <= not b or a;
    layer2_outputs(312) <= not b or a;
    layer2_outputs(313) <= b;
    layer2_outputs(314) <= not (a xor b);
    layer2_outputs(315) <= a and b;
    layer2_outputs(316) <= not (a or b);
    layer2_outputs(317) <= b;
    layer2_outputs(318) <= not b or a;
    layer2_outputs(319) <= b and not a;
    layer2_outputs(320) <= a or b;
    layer2_outputs(321) <= not (a and b);
    layer2_outputs(322) <= a;
    layer2_outputs(323) <= not (a xor b);
    layer2_outputs(324) <= not b;
    layer2_outputs(325) <= b;
    layer2_outputs(326) <= a and not b;
    layer2_outputs(327) <= a;
    layer2_outputs(328) <= not (a or b);
    layer2_outputs(329) <= a;
    layer2_outputs(330) <= not (a and b);
    layer2_outputs(331) <= b;
    layer2_outputs(332) <= not a;
    layer2_outputs(333) <= b;
    layer2_outputs(334) <= a and not b;
    layer2_outputs(335) <= b;
    layer2_outputs(336) <= not (a xor b);
    layer2_outputs(337) <= b;
    layer2_outputs(338) <= a and b;
    layer2_outputs(339) <= not a;
    layer2_outputs(340) <= a and not b;
    layer2_outputs(341) <= not a or b;
    layer2_outputs(342) <= not a;
    layer2_outputs(343) <= a;
    layer2_outputs(344) <= a and not b;
    layer2_outputs(345) <= not (a and b);
    layer2_outputs(346) <= not b;
    layer2_outputs(347) <= not b;
    layer2_outputs(348) <= not b;
    layer2_outputs(349) <= a or b;
    layer2_outputs(350) <= a and not b;
    layer2_outputs(351) <= a;
    layer2_outputs(352) <= not a;
    layer2_outputs(353) <= a or b;
    layer2_outputs(354) <= a;
    layer2_outputs(355) <= not a or b;
    layer2_outputs(356) <= not (a and b);
    layer2_outputs(357) <= not (a and b);
    layer2_outputs(358) <= b and not a;
    layer2_outputs(359) <= b;
    layer2_outputs(360) <= not (a or b);
    layer2_outputs(361) <= b and not a;
    layer2_outputs(362) <= a or b;
    layer2_outputs(363) <= not a;
    layer2_outputs(364) <= b;
    layer2_outputs(365) <= not b;
    layer2_outputs(366) <= not a;
    layer2_outputs(367) <= not (a xor b);
    layer2_outputs(368) <= a;
    layer2_outputs(369) <= a and not b;
    layer2_outputs(370) <= a and b;
    layer2_outputs(371) <= not (a xor b);
    layer2_outputs(372) <= b and not a;
    layer2_outputs(373) <= not (a or b);
    layer2_outputs(374) <= b;
    layer2_outputs(375) <= not (a or b);
    layer2_outputs(376) <= a;
    layer2_outputs(377) <= b and not a;
    layer2_outputs(378) <= a xor b;
    layer2_outputs(379) <= a;
    layer2_outputs(380) <= not (a and b);
    layer2_outputs(381) <= a;
    layer2_outputs(382) <= a;
    layer2_outputs(383) <= a and not b;
    layer2_outputs(384) <= a or b;
    layer2_outputs(385) <= a;
    layer2_outputs(386) <= a and b;
    layer2_outputs(387) <= b and not a;
    layer2_outputs(388) <= not (a and b);
    layer2_outputs(389) <= a;
    layer2_outputs(390) <= not a;
    layer2_outputs(391) <= not a or b;
    layer2_outputs(392) <= b and not a;
    layer2_outputs(393) <= not b;
    layer2_outputs(394) <= b;
    layer2_outputs(395) <= a and b;
    layer2_outputs(396) <= not (a or b);
    layer2_outputs(397) <= b;
    layer2_outputs(398) <= not (a and b);
    layer2_outputs(399) <= a;
    layer2_outputs(400) <= not a;
    layer2_outputs(401) <= b and not a;
    layer2_outputs(402) <= not a or b;
    layer2_outputs(403) <= not (a xor b);
    layer2_outputs(404) <= a or b;
    layer2_outputs(405) <= b;
    layer2_outputs(406) <= a and not b;
    layer2_outputs(407) <= not b;
    layer2_outputs(408) <= a or b;
    layer2_outputs(409) <= a;
    layer2_outputs(410) <= not b;
    layer2_outputs(411) <= not b;
    layer2_outputs(412) <= not a or b;
    layer2_outputs(413) <= not (a or b);
    layer2_outputs(414) <= a or b;
    layer2_outputs(415) <= not (a xor b);
    layer2_outputs(416) <= not (a and b);
    layer2_outputs(417) <= a xor b;
    layer2_outputs(418) <= not a;
    layer2_outputs(419) <= a xor b;
    layer2_outputs(420) <= not a;
    layer2_outputs(421) <= not b;
    layer2_outputs(422) <= b;
    layer2_outputs(423) <= not a;
    layer2_outputs(424) <= not a;
    layer2_outputs(425) <= a;
    layer2_outputs(426) <= not a or b;
    layer2_outputs(427) <= not b;
    layer2_outputs(428) <= b;
    layer2_outputs(429) <= not (a or b);
    layer2_outputs(430) <= a xor b;
    layer2_outputs(431) <= a and b;
    layer2_outputs(432) <= not a;
    layer2_outputs(433) <= not b;
    layer2_outputs(434) <= not b;
    layer2_outputs(435) <= not (a or b);
    layer2_outputs(436) <= not (a xor b);
    layer2_outputs(437) <= not b;
    layer2_outputs(438) <= not b or a;
    layer2_outputs(439) <= a and not b;
    layer2_outputs(440) <= b and not a;
    layer2_outputs(441) <= b;
    layer2_outputs(442) <= a and b;
    layer2_outputs(443) <= a;
    layer2_outputs(444) <= not (a or b);
    layer2_outputs(445) <= a and b;
    layer2_outputs(446) <= not a;
    layer2_outputs(447) <= not (a xor b);
    layer2_outputs(448) <= b;
    layer2_outputs(449) <= not a;
    layer2_outputs(450) <= not a or b;
    layer2_outputs(451) <= b and not a;
    layer2_outputs(452) <= a and b;
    layer2_outputs(453) <= not a or b;
    layer2_outputs(454) <= a;
    layer2_outputs(455) <= not (a and b);
    layer2_outputs(456) <= a and not b;
    layer2_outputs(457) <= not (a xor b);
    layer2_outputs(458) <= not (a or b);
    layer2_outputs(459) <= b and not a;
    layer2_outputs(460) <= a or b;
    layer2_outputs(461) <= b;
    layer2_outputs(462) <= b and not a;
    layer2_outputs(463) <= b and not a;
    layer2_outputs(464) <= a;
    layer2_outputs(465) <= a xor b;
    layer2_outputs(466) <= a or b;
    layer2_outputs(467) <= not (a and b);
    layer2_outputs(468) <= not b;
    layer2_outputs(469) <= a and not b;
    layer2_outputs(470) <= a and b;
    layer2_outputs(471) <= not a or b;
    layer2_outputs(472) <= a and b;
    layer2_outputs(473) <= b;
    layer2_outputs(474) <= a xor b;
    layer2_outputs(475) <= not b or a;
    layer2_outputs(476) <= a;
    layer2_outputs(477) <= a or b;
    layer2_outputs(478) <= a and b;
    layer2_outputs(479) <= a and b;
    layer2_outputs(480) <= not (a xor b);
    layer2_outputs(481) <= not (a and b);
    layer2_outputs(482) <= a;
    layer2_outputs(483) <= not b or a;
    layer2_outputs(484) <= not b or a;
    layer2_outputs(485) <= a and not b;
    layer2_outputs(486) <= b;
    layer2_outputs(487) <= not b;
    layer2_outputs(488) <= b;
    layer2_outputs(489) <= not b;
    layer2_outputs(490) <= a or b;
    layer2_outputs(491) <= b and not a;
    layer2_outputs(492) <= not b or a;
    layer2_outputs(493) <= not (a xor b);
    layer2_outputs(494) <= a and not b;
    layer2_outputs(495) <= not a;
    layer2_outputs(496) <= not b;
    layer2_outputs(497) <= not (a or b);
    layer2_outputs(498) <= not b;
    layer2_outputs(499) <= not (a and b);
    layer2_outputs(500) <= a xor b;
    layer2_outputs(501) <= not b or a;
    layer2_outputs(502) <= a;
    layer2_outputs(503) <= not a or b;
    layer2_outputs(504) <= a and not b;
    layer2_outputs(505) <= a xor b;
    layer2_outputs(506) <= not (a or b);
    layer2_outputs(507) <= a and not b;
    layer2_outputs(508) <= a xor b;
    layer2_outputs(509) <= not (a xor b);
    layer2_outputs(510) <= not a;
    layer2_outputs(511) <= not (a or b);
    layer2_outputs(512) <= not (a or b);
    layer2_outputs(513) <= a and b;
    layer2_outputs(514) <= not (a or b);
    layer2_outputs(515) <= not (a and b);
    layer2_outputs(516) <= not a;
    layer2_outputs(517) <= a;
    layer2_outputs(518) <= b;
    layer2_outputs(519) <= a;
    layer2_outputs(520) <= not a or b;
    layer2_outputs(521) <= a or b;
    layer2_outputs(522) <= not (a or b);
    layer2_outputs(523) <= not a or b;
    layer2_outputs(524) <= a xor b;
    layer2_outputs(525) <= not a or b;
    layer2_outputs(526) <= a and b;
    layer2_outputs(527) <= not (a and b);
    layer2_outputs(528) <= b and not a;
    layer2_outputs(529) <= not (a and b);
    layer2_outputs(530) <= a;
    layer2_outputs(531) <= a xor b;
    layer2_outputs(532) <= not a;
    layer2_outputs(533) <= a;
    layer2_outputs(534) <= not (a and b);
    layer2_outputs(535) <= not b or a;
    layer2_outputs(536) <= a and not b;
    layer2_outputs(537) <= a;
    layer2_outputs(538) <= b;
    layer2_outputs(539) <= 1'b1;
    layer2_outputs(540) <= b and not a;
    layer2_outputs(541) <= not (a or b);
    layer2_outputs(542) <= not a;
    layer2_outputs(543) <= not (a xor b);
    layer2_outputs(544) <= not b;
    layer2_outputs(545) <= a and b;
    layer2_outputs(546) <= a xor b;
    layer2_outputs(547) <= 1'b1;
    layer2_outputs(548) <= not (a and b);
    layer2_outputs(549) <= not b or a;
    layer2_outputs(550) <= a;
    layer2_outputs(551) <= a or b;
    layer2_outputs(552) <= not (a xor b);
    layer2_outputs(553) <= a xor b;
    layer2_outputs(554) <= not (a or b);
    layer2_outputs(555) <= not (a and b);
    layer2_outputs(556) <= a and not b;
    layer2_outputs(557) <= b and not a;
    layer2_outputs(558) <= a and not b;
    layer2_outputs(559) <= a xor b;
    layer2_outputs(560) <= a and b;
    layer2_outputs(561) <= not b;
    layer2_outputs(562) <= not b;
    layer2_outputs(563) <= not (a or b);
    layer2_outputs(564) <= not b;
    layer2_outputs(565) <= a or b;
    layer2_outputs(566) <= b;
    layer2_outputs(567) <= not (a and b);
    layer2_outputs(568) <= a;
    layer2_outputs(569) <= not b;
    layer2_outputs(570) <= not a or b;
    layer2_outputs(571) <= not a;
    layer2_outputs(572) <= b;
    layer2_outputs(573) <= a and b;
    layer2_outputs(574) <= a;
    layer2_outputs(575) <= a or b;
    layer2_outputs(576) <= not (a and b);
    layer2_outputs(577) <= a or b;
    layer2_outputs(578) <= a or b;
    layer2_outputs(579) <= not b;
    layer2_outputs(580) <= not b;
    layer2_outputs(581) <= not b;
    layer2_outputs(582) <= b;
    layer2_outputs(583) <= not (a or b);
    layer2_outputs(584) <= a;
    layer2_outputs(585) <= not (a and b);
    layer2_outputs(586) <= not a;
    layer2_outputs(587) <= b;
    layer2_outputs(588) <= a and b;
    layer2_outputs(589) <= a and not b;
    layer2_outputs(590) <= not b;
    layer2_outputs(591) <= a and not b;
    layer2_outputs(592) <= a;
    layer2_outputs(593) <= not a;
    layer2_outputs(594) <= a and b;
    layer2_outputs(595) <= b and not a;
    layer2_outputs(596) <= a;
    layer2_outputs(597) <= not a;
    layer2_outputs(598) <= a or b;
    layer2_outputs(599) <= a or b;
    layer2_outputs(600) <= not (a xor b);
    layer2_outputs(601) <= a or b;
    layer2_outputs(602) <= b;
    layer2_outputs(603) <= not b;
    layer2_outputs(604) <= not a;
    layer2_outputs(605) <= not a;
    layer2_outputs(606) <= b;
    layer2_outputs(607) <= a;
    layer2_outputs(608) <= not b or a;
    layer2_outputs(609) <= a;
    layer2_outputs(610) <= not a or b;
    layer2_outputs(611) <= not (a xor b);
    layer2_outputs(612) <= a and not b;
    layer2_outputs(613) <= not a or b;
    layer2_outputs(614) <= not a;
    layer2_outputs(615) <= b and not a;
    layer2_outputs(616) <= not a or b;
    layer2_outputs(617) <= not (a xor b);
    layer2_outputs(618) <= not (a or b);
    layer2_outputs(619) <= a;
    layer2_outputs(620) <= not b;
    layer2_outputs(621) <= a;
    layer2_outputs(622) <= not a or b;
    layer2_outputs(623) <= a;
    layer2_outputs(624) <= not a;
    layer2_outputs(625) <= a or b;
    layer2_outputs(626) <= b and not a;
    layer2_outputs(627) <= a;
    layer2_outputs(628) <= a xor b;
    layer2_outputs(629) <= a and not b;
    layer2_outputs(630) <= not a or b;
    layer2_outputs(631) <= b;
    layer2_outputs(632) <= not (a and b);
    layer2_outputs(633) <= a;
    layer2_outputs(634) <= a and not b;
    layer2_outputs(635) <= a and b;
    layer2_outputs(636) <= not (a or b);
    layer2_outputs(637) <= a;
    layer2_outputs(638) <= not (a or b);
    layer2_outputs(639) <= not (a and b);
    layer2_outputs(640) <= not (a or b);
    layer2_outputs(641) <= b and not a;
    layer2_outputs(642) <= a xor b;
    layer2_outputs(643) <= not a;
    layer2_outputs(644) <= not b;
    layer2_outputs(645) <= not (a or b);
    layer2_outputs(646) <= b;
    layer2_outputs(647) <= 1'b0;
    layer2_outputs(648) <= a;
    layer2_outputs(649) <= not (a xor b);
    layer2_outputs(650) <= a or b;
    layer2_outputs(651) <= a and b;
    layer2_outputs(652) <= not a or b;
    layer2_outputs(653) <= not b;
    layer2_outputs(654) <= not (a xor b);
    layer2_outputs(655) <= b and not a;
    layer2_outputs(656) <= b;
    layer2_outputs(657) <= a and not b;
    layer2_outputs(658) <= a or b;
    layer2_outputs(659) <= not (a xor b);
    layer2_outputs(660) <= b;
    layer2_outputs(661) <= b;
    layer2_outputs(662) <= a and not b;
    layer2_outputs(663) <= a and not b;
    layer2_outputs(664) <= 1'b1;
    layer2_outputs(665) <= a;
    layer2_outputs(666) <= a and not b;
    layer2_outputs(667) <= not (a or b);
    layer2_outputs(668) <= a and b;
    layer2_outputs(669) <= not (a xor b);
    layer2_outputs(670) <= a and b;
    layer2_outputs(671) <= b and not a;
    layer2_outputs(672) <= a;
    layer2_outputs(673) <= not b;
    layer2_outputs(674) <= b;
    layer2_outputs(675) <= not (a and b);
    layer2_outputs(676) <= not b;
    layer2_outputs(677) <= not (a and b);
    layer2_outputs(678) <= not a;
    layer2_outputs(679) <= not (a and b);
    layer2_outputs(680) <= b;
    layer2_outputs(681) <= a and not b;
    layer2_outputs(682) <= not b;
    layer2_outputs(683) <= not a or b;
    layer2_outputs(684) <= not (a or b);
    layer2_outputs(685) <= a;
    layer2_outputs(686) <= b;
    layer2_outputs(687) <= a or b;
    layer2_outputs(688) <= b;
    layer2_outputs(689) <= b;
    layer2_outputs(690) <= not (a and b);
    layer2_outputs(691) <= not b or a;
    layer2_outputs(692) <= not a;
    layer2_outputs(693) <= not (a and b);
    layer2_outputs(694) <= b;
    layer2_outputs(695) <= not b;
    layer2_outputs(696) <= not b or a;
    layer2_outputs(697) <= a and not b;
    layer2_outputs(698) <= not b;
    layer2_outputs(699) <= a xor b;
    layer2_outputs(700) <= a and b;
    layer2_outputs(701) <= not b or a;
    layer2_outputs(702) <= a and b;
    layer2_outputs(703) <= a;
    layer2_outputs(704) <= not b;
    layer2_outputs(705) <= a and not b;
    layer2_outputs(706) <= not (a or b);
    layer2_outputs(707) <= a and not b;
    layer2_outputs(708) <= a and b;
    layer2_outputs(709) <= not a;
    layer2_outputs(710) <= a;
    layer2_outputs(711) <= 1'b1;
    layer2_outputs(712) <= a xor b;
    layer2_outputs(713) <= not b or a;
    layer2_outputs(714) <= b and not a;
    layer2_outputs(715) <= a and b;
    layer2_outputs(716) <= not b or a;
    layer2_outputs(717) <= a;
    layer2_outputs(718) <= a and b;
    layer2_outputs(719) <= not (a and b);
    layer2_outputs(720) <= not b;
    layer2_outputs(721) <= not b;
    layer2_outputs(722) <= not b or a;
    layer2_outputs(723) <= b;
    layer2_outputs(724) <= not a;
    layer2_outputs(725) <= a and not b;
    layer2_outputs(726) <= a or b;
    layer2_outputs(727) <= a;
    layer2_outputs(728) <= a xor b;
    layer2_outputs(729) <= not a;
    layer2_outputs(730) <= not a or b;
    layer2_outputs(731) <= not b or a;
    layer2_outputs(732) <= a;
    layer2_outputs(733) <= b;
    layer2_outputs(734) <= not a or b;
    layer2_outputs(735) <= not b;
    layer2_outputs(736) <= not a;
    layer2_outputs(737) <= a and b;
    layer2_outputs(738) <= a and not b;
    layer2_outputs(739) <= a or b;
    layer2_outputs(740) <= a xor b;
    layer2_outputs(741) <= not (a xor b);
    layer2_outputs(742) <= not b;
    layer2_outputs(743) <= a and not b;
    layer2_outputs(744) <= not b;
    layer2_outputs(745) <= not a or b;
    layer2_outputs(746) <= b and not a;
    layer2_outputs(747) <= not b;
    layer2_outputs(748) <= not a;
    layer2_outputs(749) <= a and not b;
    layer2_outputs(750) <= a xor b;
    layer2_outputs(751) <= b;
    layer2_outputs(752) <= a xor b;
    layer2_outputs(753) <= not (a and b);
    layer2_outputs(754) <= not (a or b);
    layer2_outputs(755) <= a or b;
    layer2_outputs(756) <= a and b;
    layer2_outputs(757) <= not b;
    layer2_outputs(758) <= b and not a;
    layer2_outputs(759) <= a or b;
    layer2_outputs(760) <= not (a xor b);
    layer2_outputs(761) <= 1'b0;
    layer2_outputs(762) <= b and not a;
    layer2_outputs(763) <= a and b;
    layer2_outputs(764) <= not a or b;
    layer2_outputs(765) <= b and not a;
    layer2_outputs(766) <= not b;
    layer2_outputs(767) <= a;
    layer2_outputs(768) <= not b or a;
    layer2_outputs(769) <= b;
    layer2_outputs(770) <= b;
    layer2_outputs(771) <= not b;
    layer2_outputs(772) <= not b or a;
    layer2_outputs(773) <= not a;
    layer2_outputs(774) <= not (a and b);
    layer2_outputs(775) <= b;
    layer2_outputs(776) <= a;
    layer2_outputs(777) <= not a;
    layer2_outputs(778) <= a and b;
    layer2_outputs(779) <= not (a xor b);
    layer2_outputs(780) <= not b;
    layer2_outputs(781) <= a and not b;
    layer2_outputs(782) <= not (a or b);
    layer2_outputs(783) <= a xor b;
    layer2_outputs(784) <= not a or b;
    layer2_outputs(785) <= not (a or b);
    layer2_outputs(786) <= not a;
    layer2_outputs(787) <= not (a xor b);
    layer2_outputs(788) <= 1'b0;
    layer2_outputs(789) <= a;
    layer2_outputs(790) <= b;
    layer2_outputs(791) <= b;
    layer2_outputs(792) <= a;
    layer2_outputs(793) <= a and b;
    layer2_outputs(794) <= a or b;
    layer2_outputs(795) <= not b or a;
    layer2_outputs(796) <= not (a or b);
    layer2_outputs(797) <= not b;
    layer2_outputs(798) <= a xor b;
    layer2_outputs(799) <= not b;
    layer2_outputs(800) <= not (a xor b);
    layer2_outputs(801) <= a and b;
    layer2_outputs(802) <= not (a or b);
    layer2_outputs(803) <= not b;
    layer2_outputs(804) <= not (a and b);
    layer2_outputs(805) <= not b or a;
    layer2_outputs(806) <= not a;
    layer2_outputs(807) <= a and b;
    layer2_outputs(808) <= not (a and b);
    layer2_outputs(809) <= a and b;
    layer2_outputs(810) <= not (a xor b);
    layer2_outputs(811) <= not b;
    layer2_outputs(812) <= a and not b;
    layer2_outputs(813) <= a xor b;
    layer2_outputs(814) <= b;
    layer2_outputs(815) <= a xor b;
    layer2_outputs(816) <= a and not b;
    layer2_outputs(817) <= not b;
    layer2_outputs(818) <= b;
    layer2_outputs(819) <= b;
    layer2_outputs(820) <= not b;
    layer2_outputs(821) <= not b or a;
    layer2_outputs(822) <= not (a and b);
    layer2_outputs(823) <= a xor b;
    layer2_outputs(824) <= b;
    layer2_outputs(825) <= b;
    layer2_outputs(826) <= not (a and b);
    layer2_outputs(827) <= not a;
    layer2_outputs(828) <= not b;
    layer2_outputs(829) <= a and not b;
    layer2_outputs(830) <= not (a or b);
    layer2_outputs(831) <= not (a and b);
    layer2_outputs(832) <= not (a and b);
    layer2_outputs(833) <= a and b;
    layer2_outputs(834) <= not a or b;
    layer2_outputs(835) <= not b;
    layer2_outputs(836) <= a xor b;
    layer2_outputs(837) <= not (a or b);
    layer2_outputs(838) <= not b or a;
    layer2_outputs(839) <= a and b;
    layer2_outputs(840) <= b;
    layer2_outputs(841) <= a;
    layer2_outputs(842) <= a xor b;
    layer2_outputs(843) <= a or b;
    layer2_outputs(844) <= not a or b;
    layer2_outputs(845) <= a or b;
    layer2_outputs(846) <= not a;
    layer2_outputs(847) <= b;
    layer2_outputs(848) <= a;
    layer2_outputs(849) <= not b;
    layer2_outputs(850) <= not (a xor b);
    layer2_outputs(851) <= not (a xor b);
    layer2_outputs(852) <= not a or b;
    layer2_outputs(853) <= not a or b;
    layer2_outputs(854) <= b and not a;
    layer2_outputs(855) <= a and b;
    layer2_outputs(856) <= not b or a;
    layer2_outputs(857) <= not (a and b);
    layer2_outputs(858) <= not (a xor b);
    layer2_outputs(859) <= a;
    layer2_outputs(860) <= not b;
    layer2_outputs(861) <= a;
    layer2_outputs(862) <= not a;
    layer2_outputs(863) <= not (a xor b);
    layer2_outputs(864) <= a or b;
    layer2_outputs(865) <= not b or a;
    layer2_outputs(866) <= b;
    layer2_outputs(867) <= not (a or b);
    layer2_outputs(868) <= a and b;
    layer2_outputs(869) <= b and not a;
    layer2_outputs(870) <= not a or b;
    layer2_outputs(871) <= not a;
    layer2_outputs(872) <= not (a or b);
    layer2_outputs(873) <= not a;
    layer2_outputs(874) <= not a;
    layer2_outputs(875) <= a;
    layer2_outputs(876) <= not a;
    layer2_outputs(877) <= b and not a;
    layer2_outputs(878) <= not (a xor b);
    layer2_outputs(879) <= not b;
    layer2_outputs(880) <= a;
    layer2_outputs(881) <= a and b;
    layer2_outputs(882) <= a;
    layer2_outputs(883) <= a and b;
    layer2_outputs(884) <= not (a or b);
    layer2_outputs(885) <= a and not b;
    layer2_outputs(886) <= not b or a;
    layer2_outputs(887) <= b and not a;
    layer2_outputs(888) <= not (a or b);
    layer2_outputs(889) <= a and b;
    layer2_outputs(890) <= a and b;
    layer2_outputs(891) <= a and b;
    layer2_outputs(892) <= a;
    layer2_outputs(893) <= b;
    layer2_outputs(894) <= not (a xor b);
    layer2_outputs(895) <= not a;
    layer2_outputs(896) <= not (a and b);
    layer2_outputs(897) <= not a or b;
    layer2_outputs(898) <= b and not a;
    layer2_outputs(899) <= not a;
    layer2_outputs(900) <= not b;
    layer2_outputs(901) <= not b or a;
    layer2_outputs(902) <= not (a or b);
    layer2_outputs(903) <= a and b;
    layer2_outputs(904) <= not b;
    layer2_outputs(905) <= b and not a;
    layer2_outputs(906) <= a xor b;
    layer2_outputs(907) <= b;
    layer2_outputs(908) <= a or b;
    layer2_outputs(909) <= a and b;
    layer2_outputs(910) <= a xor b;
    layer2_outputs(911) <= not a;
    layer2_outputs(912) <= not b;
    layer2_outputs(913) <= not (a xor b);
    layer2_outputs(914) <= a and not b;
    layer2_outputs(915) <= not b;
    layer2_outputs(916) <= a;
    layer2_outputs(917) <= b;
    layer2_outputs(918) <= not (a xor b);
    layer2_outputs(919) <= a;
    layer2_outputs(920) <= a or b;
    layer2_outputs(921) <= a or b;
    layer2_outputs(922) <= b and not a;
    layer2_outputs(923) <= a;
    layer2_outputs(924) <= b;
    layer2_outputs(925) <= not (a and b);
    layer2_outputs(926) <= not (a or b);
    layer2_outputs(927) <= a and b;
    layer2_outputs(928) <= b;
    layer2_outputs(929) <= not b or a;
    layer2_outputs(930) <= not a;
    layer2_outputs(931) <= not (a or b);
    layer2_outputs(932) <= not a;
    layer2_outputs(933) <= not a or b;
    layer2_outputs(934) <= not (a and b);
    layer2_outputs(935) <= a and not b;
    layer2_outputs(936) <= not b;
    layer2_outputs(937) <= a and b;
    layer2_outputs(938) <= b and not a;
    layer2_outputs(939) <= not a;
    layer2_outputs(940) <= a;
    layer2_outputs(941) <= b;
    layer2_outputs(942) <= not a;
    layer2_outputs(943) <= not b;
    layer2_outputs(944) <= a;
    layer2_outputs(945) <= b;
    layer2_outputs(946) <= a and not b;
    layer2_outputs(947) <= not (a and b);
    layer2_outputs(948) <= not b;
    layer2_outputs(949) <= b and not a;
    layer2_outputs(950) <= a xor b;
    layer2_outputs(951) <= a and b;
    layer2_outputs(952) <= a xor b;
    layer2_outputs(953) <= a and not b;
    layer2_outputs(954) <= not a;
    layer2_outputs(955) <= a or b;
    layer2_outputs(956) <= b and not a;
    layer2_outputs(957) <= not b;
    layer2_outputs(958) <= b and not a;
    layer2_outputs(959) <= not a;
    layer2_outputs(960) <= not b;
    layer2_outputs(961) <= b;
    layer2_outputs(962) <= a;
    layer2_outputs(963) <= not (a and b);
    layer2_outputs(964) <= a or b;
    layer2_outputs(965) <= b;
    layer2_outputs(966) <= not (a xor b);
    layer2_outputs(967) <= not (a and b);
    layer2_outputs(968) <= not (a xor b);
    layer2_outputs(969) <= not (a and b);
    layer2_outputs(970) <= not (a xor b);
    layer2_outputs(971) <= b and not a;
    layer2_outputs(972) <= a;
    layer2_outputs(973) <= a xor b;
    layer2_outputs(974) <= a and b;
    layer2_outputs(975) <= a xor b;
    layer2_outputs(976) <= a and not b;
    layer2_outputs(977) <= not b;
    layer2_outputs(978) <= a or b;
    layer2_outputs(979) <= b;
    layer2_outputs(980) <= not (a or b);
    layer2_outputs(981) <= not a or b;
    layer2_outputs(982) <= not a;
    layer2_outputs(983) <= a;
    layer2_outputs(984) <= a and not b;
    layer2_outputs(985) <= a xor b;
    layer2_outputs(986) <= a xor b;
    layer2_outputs(987) <= a and not b;
    layer2_outputs(988) <= not b or a;
    layer2_outputs(989) <= not (a xor b);
    layer2_outputs(990) <= a;
    layer2_outputs(991) <= not a;
    layer2_outputs(992) <= not (a xor b);
    layer2_outputs(993) <= not a;
    layer2_outputs(994) <= a;
    layer2_outputs(995) <= not (a or b);
    layer2_outputs(996) <= not a;
    layer2_outputs(997) <= not b or a;
    layer2_outputs(998) <= not a;
    layer2_outputs(999) <= a;
    layer2_outputs(1000) <= b;
    layer2_outputs(1001) <= not a;
    layer2_outputs(1002) <= not a;
    layer2_outputs(1003) <= a xor b;
    layer2_outputs(1004) <= 1'b1;
    layer2_outputs(1005) <= b;
    layer2_outputs(1006) <= a;
    layer2_outputs(1007) <= not (a or b);
    layer2_outputs(1008) <= a xor b;
    layer2_outputs(1009) <= a;
    layer2_outputs(1010) <= not b or a;
    layer2_outputs(1011) <= not (a and b);
    layer2_outputs(1012) <= b and not a;
    layer2_outputs(1013) <= not (a or b);
    layer2_outputs(1014) <= not (a xor b);
    layer2_outputs(1015) <= a;
    layer2_outputs(1016) <= not b or a;
    layer2_outputs(1017) <= a;
    layer2_outputs(1018) <= a or b;
    layer2_outputs(1019) <= a and not b;
    layer2_outputs(1020) <= a;
    layer2_outputs(1021) <= a xor b;
    layer2_outputs(1022) <= not a;
    layer2_outputs(1023) <= a and b;
    layer2_outputs(1024) <= not b;
    layer2_outputs(1025) <= a and b;
    layer2_outputs(1026) <= b;
    layer2_outputs(1027) <= not b;
    layer2_outputs(1028) <= a xor b;
    layer2_outputs(1029) <= b;
    layer2_outputs(1030) <= a;
    layer2_outputs(1031) <= not b or a;
    layer2_outputs(1032) <= not (a and b);
    layer2_outputs(1033) <= b;
    layer2_outputs(1034) <= not b or a;
    layer2_outputs(1035) <= not b;
    layer2_outputs(1036) <= a xor b;
    layer2_outputs(1037) <= a or b;
    layer2_outputs(1038) <= not (a and b);
    layer2_outputs(1039) <= not (a and b);
    layer2_outputs(1040) <= b;
    layer2_outputs(1041) <= b and not a;
    layer2_outputs(1042) <= a;
    layer2_outputs(1043) <= a;
    layer2_outputs(1044) <= a;
    layer2_outputs(1045) <= not (a and b);
    layer2_outputs(1046) <= not a;
    layer2_outputs(1047) <= not b;
    layer2_outputs(1048) <= not (a and b);
    layer2_outputs(1049) <= not b or a;
    layer2_outputs(1050) <= not a;
    layer2_outputs(1051) <= not a or b;
    layer2_outputs(1052) <= b;
    layer2_outputs(1053) <= not a or b;
    layer2_outputs(1054) <= not (a xor b);
    layer2_outputs(1055) <= a;
    layer2_outputs(1056) <= not b;
    layer2_outputs(1057) <= a xor b;
    layer2_outputs(1058) <= a and not b;
    layer2_outputs(1059) <= not b;
    layer2_outputs(1060) <= a or b;
    layer2_outputs(1061) <= a xor b;
    layer2_outputs(1062) <= 1'b1;
    layer2_outputs(1063) <= a and b;
    layer2_outputs(1064) <= a;
    layer2_outputs(1065) <= not (a xor b);
    layer2_outputs(1066) <= b;
    layer2_outputs(1067) <= not b or a;
    layer2_outputs(1068) <= not b;
    layer2_outputs(1069) <= a;
    layer2_outputs(1070) <= b and not a;
    layer2_outputs(1071) <= not a or b;
    layer2_outputs(1072) <= a xor b;
    layer2_outputs(1073) <= not b;
    layer2_outputs(1074) <= a;
    layer2_outputs(1075) <= not a or b;
    layer2_outputs(1076) <= not b;
    layer2_outputs(1077) <= b;
    layer2_outputs(1078) <= not b or a;
    layer2_outputs(1079) <= not a or b;
    layer2_outputs(1080) <= a and b;
    layer2_outputs(1081) <= a xor b;
    layer2_outputs(1082) <= not b or a;
    layer2_outputs(1083) <= not b or a;
    layer2_outputs(1084) <= not a;
    layer2_outputs(1085) <= not b or a;
    layer2_outputs(1086) <= b and not a;
    layer2_outputs(1087) <= not (a or b);
    layer2_outputs(1088) <= a;
    layer2_outputs(1089) <= a;
    layer2_outputs(1090) <= b;
    layer2_outputs(1091) <= a and b;
    layer2_outputs(1092) <= not (a xor b);
    layer2_outputs(1093) <= not b or a;
    layer2_outputs(1094) <= a or b;
    layer2_outputs(1095) <= a xor b;
    layer2_outputs(1096) <= b;
    layer2_outputs(1097) <= not a;
    layer2_outputs(1098) <= a or b;
    layer2_outputs(1099) <= not b;
    layer2_outputs(1100) <= not a or b;
    layer2_outputs(1101) <= a;
    layer2_outputs(1102) <= 1'b0;
    layer2_outputs(1103) <= a;
    layer2_outputs(1104) <= b;
    layer2_outputs(1105) <= b;
    layer2_outputs(1106) <= not a;
    layer2_outputs(1107) <= a;
    layer2_outputs(1108) <= not (a or b);
    layer2_outputs(1109) <= not b;
    layer2_outputs(1110) <= a and b;
    layer2_outputs(1111) <= b;
    layer2_outputs(1112) <= a or b;
    layer2_outputs(1113) <= b;
    layer2_outputs(1114) <= a and b;
    layer2_outputs(1115) <= a;
    layer2_outputs(1116) <= a and b;
    layer2_outputs(1117) <= not (a xor b);
    layer2_outputs(1118) <= b;
    layer2_outputs(1119) <= a and not b;
    layer2_outputs(1120) <= 1'b1;
    layer2_outputs(1121) <= b and not a;
    layer2_outputs(1122) <= a or b;
    layer2_outputs(1123) <= b;
    layer2_outputs(1124) <= not (a and b);
    layer2_outputs(1125) <= a or b;
    layer2_outputs(1126) <= a or b;
    layer2_outputs(1127) <= not a;
    layer2_outputs(1128) <= not a;
    layer2_outputs(1129) <= a and not b;
    layer2_outputs(1130) <= not a or b;
    layer2_outputs(1131) <= not b;
    layer2_outputs(1132) <= b;
    layer2_outputs(1133) <= b;
    layer2_outputs(1134) <= b;
    layer2_outputs(1135) <= b and not a;
    layer2_outputs(1136) <= not a or b;
    layer2_outputs(1137) <= not (a xor b);
    layer2_outputs(1138) <= b and not a;
    layer2_outputs(1139) <= not (a or b);
    layer2_outputs(1140) <= a and b;
    layer2_outputs(1141) <= a;
    layer2_outputs(1142) <= a and b;
    layer2_outputs(1143) <= b;
    layer2_outputs(1144) <= not b;
    layer2_outputs(1145) <= not (a xor b);
    layer2_outputs(1146) <= a and b;
    layer2_outputs(1147) <= a xor b;
    layer2_outputs(1148) <= a and b;
    layer2_outputs(1149) <= a and not b;
    layer2_outputs(1150) <= not a;
    layer2_outputs(1151) <= not b;
    layer2_outputs(1152) <= not b or a;
    layer2_outputs(1153) <= b;
    layer2_outputs(1154) <= b;
    layer2_outputs(1155) <= b and not a;
    layer2_outputs(1156) <= not a;
    layer2_outputs(1157) <= not (a and b);
    layer2_outputs(1158) <= not (a and b);
    layer2_outputs(1159) <= a;
    layer2_outputs(1160) <= a and not b;
    layer2_outputs(1161) <= not (a xor b);
    layer2_outputs(1162) <= a xor b;
    layer2_outputs(1163) <= not (a and b);
    layer2_outputs(1164) <= not b;
    layer2_outputs(1165) <= not b or a;
    layer2_outputs(1166) <= not (a and b);
    layer2_outputs(1167) <= not b;
    layer2_outputs(1168) <= a or b;
    layer2_outputs(1169) <= not (a or b);
    layer2_outputs(1170) <= b;
    layer2_outputs(1171) <= not (a and b);
    layer2_outputs(1172) <= 1'b1;
    layer2_outputs(1173) <= b and not a;
    layer2_outputs(1174) <= not b or a;
    layer2_outputs(1175) <= not a;
    layer2_outputs(1176) <= not b or a;
    layer2_outputs(1177) <= a or b;
    layer2_outputs(1178) <= a;
    layer2_outputs(1179) <= b;
    layer2_outputs(1180) <= not (a or b);
    layer2_outputs(1181) <= not (a or b);
    layer2_outputs(1182) <= not (a or b);
    layer2_outputs(1183) <= not b;
    layer2_outputs(1184) <= a or b;
    layer2_outputs(1185) <= b;
    layer2_outputs(1186) <= b;
    layer2_outputs(1187) <= not (a xor b);
    layer2_outputs(1188) <= not (a xor b);
    layer2_outputs(1189) <= b and not a;
    layer2_outputs(1190) <= not b;
    layer2_outputs(1191) <= a and b;
    layer2_outputs(1192) <= not (a or b);
    layer2_outputs(1193) <= not (a xor b);
    layer2_outputs(1194) <= a;
    layer2_outputs(1195) <= not a or b;
    layer2_outputs(1196) <= not (a and b);
    layer2_outputs(1197) <= not a;
    layer2_outputs(1198) <= b;
    layer2_outputs(1199) <= not b;
    layer2_outputs(1200) <= a xor b;
    layer2_outputs(1201) <= b and not a;
    layer2_outputs(1202) <= not a;
    layer2_outputs(1203) <= a;
    layer2_outputs(1204) <= not (a xor b);
    layer2_outputs(1205) <= a and b;
    layer2_outputs(1206) <= b;
    layer2_outputs(1207) <= b;
    layer2_outputs(1208) <= not (a or b);
    layer2_outputs(1209) <= a and b;
    layer2_outputs(1210) <= not b;
    layer2_outputs(1211) <= not a or b;
    layer2_outputs(1212) <= b;
    layer2_outputs(1213) <= not a or b;
    layer2_outputs(1214) <= b and not a;
    layer2_outputs(1215) <= not a or b;
    layer2_outputs(1216) <= not (a and b);
    layer2_outputs(1217) <= 1'b0;
    layer2_outputs(1218) <= not (a xor b);
    layer2_outputs(1219) <= not a or b;
    layer2_outputs(1220) <= a or b;
    layer2_outputs(1221) <= not (a or b);
    layer2_outputs(1222) <= not (a xor b);
    layer2_outputs(1223) <= a and not b;
    layer2_outputs(1224) <= a;
    layer2_outputs(1225) <= b;
    layer2_outputs(1226) <= a and not b;
    layer2_outputs(1227) <= not (a or b);
    layer2_outputs(1228) <= not a or b;
    layer2_outputs(1229) <= not a or b;
    layer2_outputs(1230) <= not (a or b);
    layer2_outputs(1231) <= a or b;
    layer2_outputs(1232) <= a and not b;
    layer2_outputs(1233) <= not (a and b);
    layer2_outputs(1234) <= not (a xor b);
    layer2_outputs(1235) <= 1'b1;
    layer2_outputs(1236) <= a;
    layer2_outputs(1237) <= a;
    layer2_outputs(1238) <= not b;
    layer2_outputs(1239) <= b and not a;
    layer2_outputs(1240) <= not (a or b);
    layer2_outputs(1241) <= a;
    layer2_outputs(1242) <= a and b;
    layer2_outputs(1243) <= a xor b;
    layer2_outputs(1244) <= not (a or b);
    layer2_outputs(1245) <= a or b;
    layer2_outputs(1246) <= not (a xor b);
    layer2_outputs(1247) <= not a;
    layer2_outputs(1248) <= a and b;
    layer2_outputs(1249) <= b;
    layer2_outputs(1250) <= b and not a;
    layer2_outputs(1251) <= not (a xor b);
    layer2_outputs(1252) <= not a;
    layer2_outputs(1253) <= a and not b;
    layer2_outputs(1254) <= b;
    layer2_outputs(1255) <= not (a xor b);
    layer2_outputs(1256) <= a xor b;
    layer2_outputs(1257) <= a;
    layer2_outputs(1258) <= b and not a;
    layer2_outputs(1259) <= a or b;
    layer2_outputs(1260) <= not a or b;
    layer2_outputs(1261) <= not a;
    layer2_outputs(1262) <= not (a xor b);
    layer2_outputs(1263) <= b;
    layer2_outputs(1264) <= not a or b;
    layer2_outputs(1265) <= a;
    layer2_outputs(1266) <= a;
    layer2_outputs(1267) <= a and b;
    layer2_outputs(1268) <= a and not b;
    layer2_outputs(1269) <= not (a and b);
    layer2_outputs(1270) <= not a or b;
    layer2_outputs(1271) <= a and not b;
    layer2_outputs(1272) <= a;
    layer2_outputs(1273) <= not b;
    layer2_outputs(1274) <= not b;
    layer2_outputs(1275) <= not (a and b);
    layer2_outputs(1276) <= a;
    layer2_outputs(1277) <= a or b;
    layer2_outputs(1278) <= not a;
    layer2_outputs(1279) <= not b;
    layer2_outputs(1280) <= not b;
    layer2_outputs(1281) <= a xor b;
    layer2_outputs(1282) <= a and not b;
    layer2_outputs(1283) <= b;
    layer2_outputs(1284) <= a xor b;
    layer2_outputs(1285) <= a and b;
    layer2_outputs(1286) <= a xor b;
    layer2_outputs(1287) <= not (a xor b);
    layer2_outputs(1288) <= a;
    layer2_outputs(1289) <= b and not a;
    layer2_outputs(1290) <= not b;
    layer2_outputs(1291) <= a or b;
    layer2_outputs(1292) <= a or b;
    layer2_outputs(1293) <= not a;
    layer2_outputs(1294) <= a or b;
    layer2_outputs(1295) <= a and not b;
    layer2_outputs(1296) <= not a or b;
    layer2_outputs(1297) <= b and not a;
    layer2_outputs(1298) <= not a;
    layer2_outputs(1299) <= a or b;
    layer2_outputs(1300) <= not b;
    layer2_outputs(1301) <= not (a xor b);
    layer2_outputs(1302) <= not (a xor b);
    layer2_outputs(1303) <= a and b;
    layer2_outputs(1304) <= not b;
    layer2_outputs(1305) <= not (a or b);
    layer2_outputs(1306) <= not a;
    layer2_outputs(1307) <= a and not b;
    layer2_outputs(1308) <= a and not b;
    layer2_outputs(1309) <= a and b;
    layer2_outputs(1310) <= not (a xor b);
    layer2_outputs(1311) <= a;
    layer2_outputs(1312) <= a;
    layer2_outputs(1313) <= not (a or b);
    layer2_outputs(1314) <= b;
    layer2_outputs(1315) <= not a or b;
    layer2_outputs(1316) <= b;
    layer2_outputs(1317) <= not a;
    layer2_outputs(1318) <= not b;
    layer2_outputs(1319) <= b;
    layer2_outputs(1320) <= not a or b;
    layer2_outputs(1321) <= not (a or b);
    layer2_outputs(1322) <= a or b;
    layer2_outputs(1323) <= a xor b;
    layer2_outputs(1324) <= a or b;
    layer2_outputs(1325) <= 1'b1;
    layer2_outputs(1326) <= not (a xor b);
    layer2_outputs(1327) <= a and b;
    layer2_outputs(1328) <= not b or a;
    layer2_outputs(1329) <= not (a xor b);
    layer2_outputs(1330) <= a and not b;
    layer2_outputs(1331) <= a;
    layer2_outputs(1332) <= a and not b;
    layer2_outputs(1333) <= b and not a;
    layer2_outputs(1334) <= a xor b;
    layer2_outputs(1335) <= not b;
    layer2_outputs(1336) <= not (a and b);
    layer2_outputs(1337) <= not (a xor b);
    layer2_outputs(1338) <= not (a xor b);
    layer2_outputs(1339) <= not b;
    layer2_outputs(1340) <= not a or b;
    layer2_outputs(1341) <= not (a and b);
    layer2_outputs(1342) <= a or b;
    layer2_outputs(1343) <= a;
    layer2_outputs(1344) <= b and not a;
    layer2_outputs(1345) <= not (a or b);
    layer2_outputs(1346) <= not a;
    layer2_outputs(1347) <= not a or b;
    layer2_outputs(1348) <= not a or b;
    layer2_outputs(1349) <= a or b;
    layer2_outputs(1350) <= not b;
    layer2_outputs(1351) <= not (a and b);
    layer2_outputs(1352) <= b;
    layer2_outputs(1353) <= not (a xor b);
    layer2_outputs(1354) <= a or b;
    layer2_outputs(1355) <= not (a or b);
    layer2_outputs(1356) <= not a;
    layer2_outputs(1357) <= not b;
    layer2_outputs(1358) <= not b or a;
    layer2_outputs(1359) <= not (a and b);
    layer2_outputs(1360) <= b and not a;
    layer2_outputs(1361) <= not (a or b);
    layer2_outputs(1362) <= a;
    layer2_outputs(1363) <= not a or b;
    layer2_outputs(1364) <= not a;
    layer2_outputs(1365) <= not (a xor b);
    layer2_outputs(1366) <= not (a xor b);
    layer2_outputs(1367) <= a and b;
    layer2_outputs(1368) <= not b;
    layer2_outputs(1369) <= a xor b;
    layer2_outputs(1370) <= a or b;
    layer2_outputs(1371) <= not a or b;
    layer2_outputs(1372) <= a and not b;
    layer2_outputs(1373) <= not b or a;
    layer2_outputs(1374) <= not (a xor b);
    layer2_outputs(1375) <= b;
    layer2_outputs(1376) <= not (a and b);
    layer2_outputs(1377) <= not (a and b);
    layer2_outputs(1378) <= not (a and b);
    layer2_outputs(1379) <= b;
    layer2_outputs(1380) <= not a;
    layer2_outputs(1381) <= not b;
    layer2_outputs(1382) <= a xor b;
    layer2_outputs(1383) <= a and not b;
    layer2_outputs(1384) <= not (a and b);
    layer2_outputs(1385) <= a and not b;
    layer2_outputs(1386) <= not b or a;
    layer2_outputs(1387) <= not (a xor b);
    layer2_outputs(1388) <= b;
    layer2_outputs(1389) <= not b or a;
    layer2_outputs(1390) <= not b or a;
    layer2_outputs(1391) <= not b or a;
    layer2_outputs(1392) <= a or b;
    layer2_outputs(1393) <= a;
    layer2_outputs(1394) <= a and not b;
    layer2_outputs(1395) <= not (a and b);
    layer2_outputs(1396) <= a xor b;
    layer2_outputs(1397) <= b and not a;
    layer2_outputs(1398) <= not b;
    layer2_outputs(1399) <= a xor b;
    layer2_outputs(1400) <= not b or a;
    layer2_outputs(1401) <= not b;
    layer2_outputs(1402) <= not (a or b);
    layer2_outputs(1403) <= not b;
    layer2_outputs(1404) <= not (a and b);
    layer2_outputs(1405) <= a xor b;
    layer2_outputs(1406) <= a and b;
    layer2_outputs(1407) <= 1'b1;
    layer2_outputs(1408) <= not a;
    layer2_outputs(1409) <= a;
    layer2_outputs(1410) <= not b or a;
    layer2_outputs(1411) <= b and not a;
    layer2_outputs(1412) <= a and not b;
    layer2_outputs(1413) <= not b or a;
    layer2_outputs(1414) <= b and not a;
    layer2_outputs(1415) <= not (a or b);
    layer2_outputs(1416) <= a and not b;
    layer2_outputs(1417) <= not (a and b);
    layer2_outputs(1418) <= not b or a;
    layer2_outputs(1419) <= a and not b;
    layer2_outputs(1420) <= b;
    layer2_outputs(1421) <= not a or b;
    layer2_outputs(1422) <= a xor b;
    layer2_outputs(1423) <= not (a and b);
    layer2_outputs(1424) <= not (a or b);
    layer2_outputs(1425) <= not (a xor b);
    layer2_outputs(1426) <= b;
    layer2_outputs(1427) <= a xor b;
    layer2_outputs(1428) <= not (a and b);
    layer2_outputs(1429) <= not (a and b);
    layer2_outputs(1430) <= a xor b;
    layer2_outputs(1431) <= not (a or b);
    layer2_outputs(1432) <= a;
    layer2_outputs(1433) <= a;
    layer2_outputs(1434) <= a or b;
    layer2_outputs(1435) <= a or b;
    layer2_outputs(1436) <= not (a or b);
    layer2_outputs(1437) <= not a;
    layer2_outputs(1438) <= not (a or b);
    layer2_outputs(1439) <= not b;
    layer2_outputs(1440) <= not (a xor b);
    layer2_outputs(1441) <= a;
    layer2_outputs(1442) <= not a;
    layer2_outputs(1443) <= not a;
    layer2_outputs(1444) <= a;
    layer2_outputs(1445) <= not a;
    layer2_outputs(1446) <= not b;
    layer2_outputs(1447) <= not b or a;
    layer2_outputs(1448) <= a or b;
    layer2_outputs(1449) <= not a;
    layer2_outputs(1450) <= a xor b;
    layer2_outputs(1451) <= not (a or b);
    layer2_outputs(1452) <= not a;
    layer2_outputs(1453) <= not (a or b);
    layer2_outputs(1454) <= a;
    layer2_outputs(1455) <= not b;
    layer2_outputs(1456) <= a or b;
    layer2_outputs(1457) <= not (a xor b);
    layer2_outputs(1458) <= a;
    layer2_outputs(1459) <= not b or a;
    layer2_outputs(1460) <= not a;
    layer2_outputs(1461) <= not (a xor b);
    layer2_outputs(1462) <= a;
    layer2_outputs(1463) <= b;
    layer2_outputs(1464) <= not (a xor b);
    layer2_outputs(1465) <= not (a and b);
    layer2_outputs(1466) <= a xor b;
    layer2_outputs(1467) <= a;
    layer2_outputs(1468) <= not a or b;
    layer2_outputs(1469) <= a xor b;
    layer2_outputs(1470) <= b;
    layer2_outputs(1471) <= not a or b;
    layer2_outputs(1472) <= not b or a;
    layer2_outputs(1473) <= not (a and b);
    layer2_outputs(1474) <= a or b;
    layer2_outputs(1475) <= not b or a;
    layer2_outputs(1476) <= a or b;
    layer2_outputs(1477) <= a;
    layer2_outputs(1478) <= not a;
    layer2_outputs(1479) <= not b or a;
    layer2_outputs(1480) <= a;
    layer2_outputs(1481) <= b and not a;
    layer2_outputs(1482) <= not (a or b);
    layer2_outputs(1483) <= a xor b;
    layer2_outputs(1484) <= a xor b;
    layer2_outputs(1485) <= not (a and b);
    layer2_outputs(1486) <= a and not b;
    layer2_outputs(1487) <= a;
    layer2_outputs(1488) <= a xor b;
    layer2_outputs(1489) <= a and b;
    layer2_outputs(1490) <= not a or b;
    layer2_outputs(1491) <= not a or b;
    layer2_outputs(1492) <= a and not b;
    layer2_outputs(1493) <= a xor b;
    layer2_outputs(1494) <= a;
    layer2_outputs(1495) <= a and not b;
    layer2_outputs(1496) <= not (a xor b);
    layer2_outputs(1497) <= not (a and b);
    layer2_outputs(1498) <= not a;
    layer2_outputs(1499) <= not a;
    layer2_outputs(1500) <= b;
    layer2_outputs(1501) <= a;
    layer2_outputs(1502) <= not a;
    layer2_outputs(1503) <= not (a xor b);
    layer2_outputs(1504) <= not b;
    layer2_outputs(1505) <= a xor b;
    layer2_outputs(1506) <= not (a and b);
    layer2_outputs(1507) <= not a or b;
    layer2_outputs(1508) <= a xor b;
    layer2_outputs(1509) <= a and not b;
    layer2_outputs(1510) <= not (a and b);
    layer2_outputs(1511) <= not (a and b);
    layer2_outputs(1512) <= a or b;
    layer2_outputs(1513) <= not a;
    layer2_outputs(1514) <= not a;
    layer2_outputs(1515) <= a or b;
    layer2_outputs(1516) <= not a;
    layer2_outputs(1517) <= a xor b;
    layer2_outputs(1518) <= not a or b;
    layer2_outputs(1519) <= b;
    layer2_outputs(1520) <= not b;
    layer2_outputs(1521) <= not (a xor b);
    layer2_outputs(1522) <= not b;
    layer2_outputs(1523) <= b;
    layer2_outputs(1524) <= not b;
    layer2_outputs(1525) <= b and not a;
    layer2_outputs(1526) <= not (a xor b);
    layer2_outputs(1527) <= not b;
    layer2_outputs(1528) <= not a;
    layer2_outputs(1529) <= a xor b;
    layer2_outputs(1530) <= not (a or b);
    layer2_outputs(1531) <= not b;
    layer2_outputs(1532) <= not (a xor b);
    layer2_outputs(1533) <= not (a or b);
    layer2_outputs(1534) <= a or b;
    layer2_outputs(1535) <= not b;
    layer2_outputs(1536) <= not a;
    layer2_outputs(1537) <= not b or a;
    layer2_outputs(1538) <= not a;
    layer2_outputs(1539) <= not b or a;
    layer2_outputs(1540) <= not (a and b);
    layer2_outputs(1541) <= a and b;
    layer2_outputs(1542) <= not b;
    layer2_outputs(1543) <= b;
    layer2_outputs(1544) <= not (a and b);
    layer2_outputs(1545) <= not (a and b);
    layer2_outputs(1546) <= not (a xor b);
    layer2_outputs(1547) <= not b;
    layer2_outputs(1548) <= not a;
    layer2_outputs(1549) <= not (a xor b);
    layer2_outputs(1550) <= not a or b;
    layer2_outputs(1551) <= not a;
    layer2_outputs(1552) <= b;
    layer2_outputs(1553) <= not b;
    layer2_outputs(1554) <= not (a xor b);
    layer2_outputs(1555) <= b and not a;
    layer2_outputs(1556) <= not a or b;
    layer2_outputs(1557) <= a or b;
    layer2_outputs(1558) <= not a;
    layer2_outputs(1559) <= b and not a;
    layer2_outputs(1560) <= b;
    layer2_outputs(1561) <= b and not a;
    layer2_outputs(1562) <= not b;
    layer2_outputs(1563) <= not b or a;
    layer2_outputs(1564) <= not a;
    layer2_outputs(1565) <= a;
    layer2_outputs(1566) <= not b or a;
    layer2_outputs(1567) <= a and not b;
    layer2_outputs(1568) <= a;
    layer2_outputs(1569) <= a and not b;
    layer2_outputs(1570) <= not b or a;
    layer2_outputs(1571) <= a;
    layer2_outputs(1572) <= a xor b;
    layer2_outputs(1573) <= a xor b;
    layer2_outputs(1574) <= not (a or b);
    layer2_outputs(1575) <= a or b;
    layer2_outputs(1576) <= a or b;
    layer2_outputs(1577) <= not a;
    layer2_outputs(1578) <= 1'b0;
    layer2_outputs(1579) <= 1'b1;
    layer2_outputs(1580) <= not b or a;
    layer2_outputs(1581) <= not a or b;
    layer2_outputs(1582) <= a and b;
    layer2_outputs(1583) <= not a or b;
    layer2_outputs(1584) <= not a;
    layer2_outputs(1585) <= a;
    layer2_outputs(1586) <= a;
    layer2_outputs(1587) <= not (a xor b);
    layer2_outputs(1588) <= not b;
    layer2_outputs(1589) <= a xor b;
    layer2_outputs(1590) <= b;
    layer2_outputs(1591) <= not b;
    layer2_outputs(1592) <= b;
    layer2_outputs(1593) <= a;
    layer2_outputs(1594) <= b;
    layer2_outputs(1595) <= b and not a;
    layer2_outputs(1596) <= not (a or b);
    layer2_outputs(1597) <= not a;
    layer2_outputs(1598) <= not a or b;
    layer2_outputs(1599) <= a and b;
    layer2_outputs(1600) <= not (a or b);
    layer2_outputs(1601) <= a and not b;
    layer2_outputs(1602) <= not a;
    layer2_outputs(1603) <= not (a and b);
    layer2_outputs(1604) <= a and not b;
    layer2_outputs(1605) <= a;
    layer2_outputs(1606) <= a and not b;
    layer2_outputs(1607) <= not (a and b);
    layer2_outputs(1608) <= a;
    layer2_outputs(1609) <= b;
    layer2_outputs(1610) <= b;
    layer2_outputs(1611) <= not b;
    layer2_outputs(1612) <= b and not a;
    layer2_outputs(1613) <= not a or b;
    layer2_outputs(1614) <= a and not b;
    layer2_outputs(1615) <= not a;
    layer2_outputs(1616) <= not (a and b);
    layer2_outputs(1617) <= not a;
    layer2_outputs(1618) <= a or b;
    layer2_outputs(1619) <= a and b;
    layer2_outputs(1620) <= not (a and b);
    layer2_outputs(1621) <= not a or b;
    layer2_outputs(1622) <= a or b;
    layer2_outputs(1623) <= a or b;
    layer2_outputs(1624) <= b;
    layer2_outputs(1625) <= not b;
    layer2_outputs(1626) <= b and not a;
    layer2_outputs(1627) <= a xor b;
    layer2_outputs(1628) <= not (a and b);
    layer2_outputs(1629) <= not a;
    layer2_outputs(1630) <= a and not b;
    layer2_outputs(1631) <= not b;
    layer2_outputs(1632) <= not a or b;
    layer2_outputs(1633) <= not (a or b);
    layer2_outputs(1634) <= not a;
    layer2_outputs(1635) <= not b;
    layer2_outputs(1636) <= b;
    layer2_outputs(1637) <= not a;
    layer2_outputs(1638) <= a and not b;
    layer2_outputs(1639) <= not a or b;
    layer2_outputs(1640) <= not a;
    layer2_outputs(1641) <= b;
    layer2_outputs(1642) <= a;
    layer2_outputs(1643) <= a or b;
    layer2_outputs(1644) <= b;
    layer2_outputs(1645) <= not (a or b);
    layer2_outputs(1646) <= not (a xor b);
    layer2_outputs(1647) <= not b;
    layer2_outputs(1648) <= not (a or b);
    layer2_outputs(1649) <= a and b;
    layer2_outputs(1650) <= not b or a;
    layer2_outputs(1651) <= not a or b;
    layer2_outputs(1652) <= not (a and b);
    layer2_outputs(1653) <= a and b;
    layer2_outputs(1654) <= not a;
    layer2_outputs(1655) <= not b;
    layer2_outputs(1656) <= not b or a;
    layer2_outputs(1657) <= b;
    layer2_outputs(1658) <= a and not b;
    layer2_outputs(1659) <= not (a xor b);
    layer2_outputs(1660) <= not b or a;
    layer2_outputs(1661) <= not a;
    layer2_outputs(1662) <= not (a or b);
    layer2_outputs(1663) <= a xor b;
    layer2_outputs(1664) <= not a or b;
    layer2_outputs(1665) <= b;
    layer2_outputs(1666) <= not a;
    layer2_outputs(1667) <= not a;
    layer2_outputs(1668) <= a xor b;
    layer2_outputs(1669) <= a;
    layer2_outputs(1670) <= a xor b;
    layer2_outputs(1671) <= not (a or b);
    layer2_outputs(1672) <= not (a and b);
    layer2_outputs(1673) <= not b or a;
    layer2_outputs(1674) <= not b or a;
    layer2_outputs(1675) <= a and not b;
    layer2_outputs(1676) <= not b;
    layer2_outputs(1677) <= not a;
    layer2_outputs(1678) <= a;
    layer2_outputs(1679) <= a and b;
    layer2_outputs(1680) <= not (a or b);
    layer2_outputs(1681) <= b;
    layer2_outputs(1682) <= a or b;
    layer2_outputs(1683) <= a and not b;
    layer2_outputs(1684) <= not (a or b);
    layer2_outputs(1685) <= b;
    layer2_outputs(1686) <= not b or a;
    layer2_outputs(1687) <= b and not a;
    layer2_outputs(1688) <= b and not a;
    layer2_outputs(1689) <= not a or b;
    layer2_outputs(1690) <= not a;
    layer2_outputs(1691) <= a xor b;
    layer2_outputs(1692) <= b and not a;
    layer2_outputs(1693) <= a xor b;
    layer2_outputs(1694) <= a;
    layer2_outputs(1695) <= not (a xor b);
    layer2_outputs(1696) <= not (a xor b);
    layer2_outputs(1697) <= a and not b;
    layer2_outputs(1698) <= not a or b;
    layer2_outputs(1699) <= a xor b;
    layer2_outputs(1700) <= a;
    layer2_outputs(1701) <= a or b;
    layer2_outputs(1702) <= a or b;
    layer2_outputs(1703) <= b;
    layer2_outputs(1704) <= 1'b0;
    layer2_outputs(1705) <= not (a xor b);
    layer2_outputs(1706) <= a or b;
    layer2_outputs(1707) <= not (a and b);
    layer2_outputs(1708) <= not b or a;
    layer2_outputs(1709) <= not a;
    layer2_outputs(1710) <= a;
    layer2_outputs(1711) <= not a or b;
    layer2_outputs(1712) <= b;
    layer2_outputs(1713) <= not a;
    layer2_outputs(1714) <= not (a and b);
    layer2_outputs(1715) <= not a or b;
    layer2_outputs(1716) <= not a or b;
    layer2_outputs(1717) <= a and b;
    layer2_outputs(1718) <= b;
    layer2_outputs(1719) <= not (a and b);
    layer2_outputs(1720) <= a and b;
    layer2_outputs(1721) <= b;
    layer2_outputs(1722) <= a;
    layer2_outputs(1723) <= not (a and b);
    layer2_outputs(1724) <= not a;
    layer2_outputs(1725) <= a xor b;
    layer2_outputs(1726) <= not b;
    layer2_outputs(1727) <= a and not b;
    layer2_outputs(1728) <= not b;
    layer2_outputs(1729) <= not b;
    layer2_outputs(1730) <= not (a and b);
    layer2_outputs(1731) <= not (a or b);
    layer2_outputs(1732) <= a and b;
    layer2_outputs(1733) <= a and b;
    layer2_outputs(1734) <= not a;
    layer2_outputs(1735) <= b;
    layer2_outputs(1736) <= a and b;
    layer2_outputs(1737) <= not b;
    layer2_outputs(1738) <= not (a and b);
    layer2_outputs(1739) <= not b or a;
    layer2_outputs(1740) <= not b or a;
    layer2_outputs(1741) <= a or b;
    layer2_outputs(1742) <= not (a or b);
    layer2_outputs(1743) <= not (a and b);
    layer2_outputs(1744) <= not (a xor b);
    layer2_outputs(1745) <= a;
    layer2_outputs(1746) <= a;
    layer2_outputs(1747) <= not (a and b);
    layer2_outputs(1748) <= not b or a;
    layer2_outputs(1749) <= not (a and b);
    layer2_outputs(1750) <= a;
    layer2_outputs(1751) <= a;
    layer2_outputs(1752) <= a and not b;
    layer2_outputs(1753) <= not (a xor b);
    layer2_outputs(1754) <= not a;
    layer2_outputs(1755) <= not a or b;
    layer2_outputs(1756) <= not a;
    layer2_outputs(1757) <= a;
    layer2_outputs(1758) <= b;
    layer2_outputs(1759) <= a or b;
    layer2_outputs(1760) <= not a;
    layer2_outputs(1761) <= not (a and b);
    layer2_outputs(1762) <= b and not a;
    layer2_outputs(1763) <= a and b;
    layer2_outputs(1764) <= a and b;
    layer2_outputs(1765) <= a xor b;
    layer2_outputs(1766) <= b and not a;
    layer2_outputs(1767) <= a;
    layer2_outputs(1768) <= a xor b;
    layer2_outputs(1769) <= b;
    layer2_outputs(1770) <= b and not a;
    layer2_outputs(1771) <= b;
    layer2_outputs(1772) <= b;
    layer2_outputs(1773) <= a;
    layer2_outputs(1774) <= a and not b;
    layer2_outputs(1775) <= not a or b;
    layer2_outputs(1776) <= a and not b;
    layer2_outputs(1777) <= not a;
    layer2_outputs(1778) <= a or b;
    layer2_outputs(1779) <= a and b;
    layer2_outputs(1780) <= not b or a;
    layer2_outputs(1781) <= b;
    layer2_outputs(1782) <= not b;
    layer2_outputs(1783) <= not (a and b);
    layer2_outputs(1784) <= not (a or b);
    layer2_outputs(1785) <= not a;
    layer2_outputs(1786) <= not (a xor b);
    layer2_outputs(1787) <= a xor b;
    layer2_outputs(1788) <= not b or a;
    layer2_outputs(1789) <= not b or a;
    layer2_outputs(1790) <= not a or b;
    layer2_outputs(1791) <= not a;
    layer2_outputs(1792) <= a;
    layer2_outputs(1793) <= b;
    layer2_outputs(1794) <= a and b;
    layer2_outputs(1795) <= a or b;
    layer2_outputs(1796) <= not a;
    layer2_outputs(1797) <= not b;
    layer2_outputs(1798) <= a or b;
    layer2_outputs(1799) <= not a;
    layer2_outputs(1800) <= b;
    layer2_outputs(1801) <= not (a xor b);
    layer2_outputs(1802) <= a and b;
    layer2_outputs(1803) <= not (a xor b);
    layer2_outputs(1804) <= a xor b;
    layer2_outputs(1805) <= not (a or b);
    layer2_outputs(1806) <= not a or b;
    layer2_outputs(1807) <= not a or b;
    layer2_outputs(1808) <= a xor b;
    layer2_outputs(1809) <= b;
    layer2_outputs(1810) <= not b;
    layer2_outputs(1811) <= not a or b;
    layer2_outputs(1812) <= a xor b;
    layer2_outputs(1813) <= a;
    layer2_outputs(1814) <= a or b;
    layer2_outputs(1815) <= b;
    layer2_outputs(1816) <= a;
    layer2_outputs(1817) <= not b or a;
    layer2_outputs(1818) <= a and not b;
    layer2_outputs(1819) <= not b;
    layer2_outputs(1820) <= not b or a;
    layer2_outputs(1821) <= b;
    layer2_outputs(1822) <= not b or a;
    layer2_outputs(1823) <= not (a or b);
    layer2_outputs(1824) <= not a or b;
    layer2_outputs(1825) <= b and not a;
    layer2_outputs(1826) <= b and not a;
    layer2_outputs(1827) <= a and b;
    layer2_outputs(1828) <= b;
    layer2_outputs(1829) <= a or b;
    layer2_outputs(1830) <= not a;
    layer2_outputs(1831) <= a;
    layer2_outputs(1832) <= a;
    layer2_outputs(1833) <= not a or b;
    layer2_outputs(1834) <= a;
    layer2_outputs(1835) <= not a;
    layer2_outputs(1836) <= not (a xor b);
    layer2_outputs(1837) <= not b;
    layer2_outputs(1838) <= not a;
    layer2_outputs(1839) <= not b;
    layer2_outputs(1840) <= b;
    layer2_outputs(1841) <= a or b;
    layer2_outputs(1842) <= a;
    layer2_outputs(1843) <= a;
    layer2_outputs(1844) <= not (a and b);
    layer2_outputs(1845) <= b;
    layer2_outputs(1846) <= a and not b;
    layer2_outputs(1847) <= a and b;
    layer2_outputs(1848) <= not b or a;
    layer2_outputs(1849) <= not (a and b);
    layer2_outputs(1850) <= a;
    layer2_outputs(1851) <= a;
    layer2_outputs(1852) <= a or b;
    layer2_outputs(1853) <= a or b;
    layer2_outputs(1854) <= not a or b;
    layer2_outputs(1855) <= b and not a;
    layer2_outputs(1856) <= b;
    layer2_outputs(1857) <= not b or a;
    layer2_outputs(1858) <= b and not a;
    layer2_outputs(1859) <= a and b;
    layer2_outputs(1860) <= not b;
    layer2_outputs(1861) <= b;
    layer2_outputs(1862) <= not b or a;
    layer2_outputs(1863) <= a or b;
    layer2_outputs(1864) <= not (a xor b);
    layer2_outputs(1865) <= not (a and b);
    layer2_outputs(1866) <= not a or b;
    layer2_outputs(1867) <= not b;
    layer2_outputs(1868) <= a;
    layer2_outputs(1869) <= a;
    layer2_outputs(1870) <= a or b;
    layer2_outputs(1871) <= a and not b;
    layer2_outputs(1872) <= not a or b;
    layer2_outputs(1873) <= b and not a;
    layer2_outputs(1874) <= not (a or b);
    layer2_outputs(1875) <= not b;
    layer2_outputs(1876) <= b;
    layer2_outputs(1877) <= 1'b0;
    layer2_outputs(1878) <= not b;
    layer2_outputs(1879) <= a;
    layer2_outputs(1880) <= not a or b;
    layer2_outputs(1881) <= not a;
    layer2_outputs(1882) <= a and not b;
    layer2_outputs(1883) <= a and not b;
    layer2_outputs(1884) <= not a or b;
    layer2_outputs(1885) <= a xor b;
    layer2_outputs(1886) <= not (a xor b);
    layer2_outputs(1887) <= not b;
    layer2_outputs(1888) <= a;
    layer2_outputs(1889) <= not b or a;
    layer2_outputs(1890) <= b;
    layer2_outputs(1891) <= a or b;
    layer2_outputs(1892) <= a;
    layer2_outputs(1893) <= a xor b;
    layer2_outputs(1894) <= not b or a;
    layer2_outputs(1895) <= a;
    layer2_outputs(1896) <= not b;
    layer2_outputs(1897) <= not a;
    layer2_outputs(1898) <= not (a or b);
    layer2_outputs(1899) <= not b;
    layer2_outputs(1900) <= a xor b;
    layer2_outputs(1901) <= not a;
    layer2_outputs(1902) <= a or b;
    layer2_outputs(1903) <= not a;
    layer2_outputs(1904) <= not a or b;
    layer2_outputs(1905) <= not (a and b);
    layer2_outputs(1906) <= a or b;
    layer2_outputs(1907) <= not (a xor b);
    layer2_outputs(1908) <= 1'b0;
    layer2_outputs(1909) <= not (a or b);
    layer2_outputs(1910) <= not (a and b);
    layer2_outputs(1911) <= a and not b;
    layer2_outputs(1912) <= b and not a;
    layer2_outputs(1913) <= not a;
    layer2_outputs(1914) <= not b;
    layer2_outputs(1915) <= not b;
    layer2_outputs(1916) <= b;
    layer2_outputs(1917) <= not b;
    layer2_outputs(1918) <= a and b;
    layer2_outputs(1919) <= a and not b;
    layer2_outputs(1920) <= not a or b;
    layer2_outputs(1921) <= not (a xor b);
    layer2_outputs(1922) <= a;
    layer2_outputs(1923) <= b;
    layer2_outputs(1924) <= b and not a;
    layer2_outputs(1925) <= a and not b;
    layer2_outputs(1926) <= b;
    layer2_outputs(1927) <= not (a xor b);
    layer2_outputs(1928) <= not b;
    layer2_outputs(1929) <= a;
    layer2_outputs(1930) <= a;
    layer2_outputs(1931) <= not (a and b);
    layer2_outputs(1932) <= b and not a;
    layer2_outputs(1933) <= b;
    layer2_outputs(1934) <= a and b;
    layer2_outputs(1935) <= not (a or b);
    layer2_outputs(1936) <= b;
    layer2_outputs(1937) <= a or b;
    layer2_outputs(1938) <= b;
    layer2_outputs(1939) <= b;
    layer2_outputs(1940) <= not b or a;
    layer2_outputs(1941) <= a;
    layer2_outputs(1942) <= not b or a;
    layer2_outputs(1943) <= a or b;
    layer2_outputs(1944) <= a;
    layer2_outputs(1945) <= not b or a;
    layer2_outputs(1946) <= a;
    layer2_outputs(1947) <= a xor b;
    layer2_outputs(1948) <= not a or b;
    layer2_outputs(1949) <= not (a or b);
    layer2_outputs(1950) <= not b;
    layer2_outputs(1951) <= a and not b;
    layer2_outputs(1952) <= a;
    layer2_outputs(1953) <= not b or a;
    layer2_outputs(1954) <= b;
    layer2_outputs(1955) <= a;
    layer2_outputs(1956) <= a and not b;
    layer2_outputs(1957) <= not b or a;
    layer2_outputs(1958) <= not b or a;
    layer2_outputs(1959) <= not a;
    layer2_outputs(1960) <= not a;
    layer2_outputs(1961) <= not a;
    layer2_outputs(1962) <= a xor b;
    layer2_outputs(1963) <= a or b;
    layer2_outputs(1964) <= b;
    layer2_outputs(1965) <= not (a or b);
    layer2_outputs(1966) <= a or b;
    layer2_outputs(1967) <= a and not b;
    layer2_outputs(1968) <= b and not a;
    layer2_outputs(1969) <= a and not b;
    layer2_outputs(1970) <= not (a xor b);
    layer2_outputs(1971) <= not a;
    layer2_outputs(1972) <= a xor b;
    layer2_outputs(1973) <= a and b;
    layer2_outputs(1974) <= b;
    layer2_outputs(1975) <= a xor b;
    layer2_outputs(1976) <= not a;
    layer2_outputs(1977) <= not a;
    layer2_outputs(1978) <= b;
    layer2_outputs(1979) <= a and b;
    layer2_outputs(1980) <= a xor b;
    layer2_outputs(1981) <= a;
    layer2_outputs(1982) <= not a;
    layer2_outputs(1983) <= a and b;
    layer2_outputs(1984) <= not (a xor b);
    layer2_outputs(1985) <= b and not a;
    layer2_outputs(1986) <= b;
    layer2_outputs(1987) <= not b or a;
    layer2_outputs(1988) <= not (a and b);
    layer2_outputs(1989) <= 1'b1;
    layer2_outputs(1990) <= not (a xor b);
    layer2_outputs(1991) <= b;
    layer2_outputs(1992) <= a;
    layer2_outputs(1993) <= not a or b;
    layer2_outputs(1994) <= not (a or b);
    layer2_outputs(1995) <= b and not a;
    layer2_outputs(1996) <= a and b;
    layer2_outputs(1997) <= not b;
    layer2_outputs(1998) <= not a;
    layer2_outputs(1999) <= not b;
    layer2_outputs(2000) <= not a or b;
    layer2_outputs(2001) <= not a or b;
    layer2_outputs(2002) <= 1'b1;
    layer2_outputs(2003) <= a xor b;
    layer2_outputs(2004) <= a or b;
    layer2_outputs(2005) <= not b;
    layer2_outputs(2006) <= a and not b;
    layer2_outputs(2007) <= not a;
    layer2_outputs(2008) <= not b;
    layer2_outputs(2009) <= not (a and b);
    layer2_outputs(2010) <= a and not b;
    layer2_outputs(2011) <= not a or b;
    layer2_outputs(2012) <= not (a xor b);
    layer2_outputs(2013) <= a;
    layer2_outputs(2014) <= not a;
    layer2_outputs(2015) <= b and not a;
    layer2_outputs(2016) <= a xor b;
    layer2_outputs(2017) <= not (a or b);
    layer2_outputs(2018) <= a xor b;
    layer2_outputs(2019) <= not a or b;
    layer2_outputs(2020) <= not (a xor b);
    layer2_outputs(2021) <= not b;
    layer2_outputs(2022) <= not a;
    layer2_outputs(2023) <= not a or b;
    layer2_outputs(2024) <= a;
    layer2_outputs(2025) <= a xor b;
    layer2_outputs(2026) <= not b or a;
    layer2_outputs(2027) <= not a;
    layer2_outputs(2028) <= a and b;
    layer2_outputs(2029) <= not b;
    layer2_outputs(2030) <= not (a and b);
    layer2_outputs(2031) <= not a or b;
    layer2_outputs(2032) <= not (a xor b);
    layer2_outputs(2033) <= b;
    layer2_outputs(2034) <= not b;
    layer2_outputs(2035) <= not a;
    layer2_outputs(2036) <= not (a xor b);
    layer2_outputs(2037) <= a or b;
    layer2_outputs(2038) <= not a;
    layer2_outputs(2039) <= not (a or b);
    layer2_outputs(2040) <= a;
    layer2_outputs(2041) <= not b;
    layer2_outputs(2042) <= not b;
    layer2_outputs(2043) <= a and b;
    layer2_outputs(2044) <= not a;
    layer2_outputs(2045) <= a;
    layer2_outputs(2046) <= not b;
    layer2_outputs(2047) <= b;
    layer2_outputs(2048) <= not a;
    layer2_outputs(2049) <= a;
    layer2_outputs(2050) <= not (a or b);
    layer2_outputs(2051) <= 1'b0;
    layer2_outputs(2052) <= not a;
    layer2_outputs(2053) <= a and not b;
    layer2_outputs(2054) <= a and not b;
    layer2_outputs(2055) <= not (a xor b);
    layer2_outputs(2056) <= a xor b;
    layer2_outputs(2057) <= not (a and b);
    layer2_outputs(2058) <= not b;
    layer2_outputs(2059) <= not b or a;
    layer2_outputs(2060) <= not a;
    layer2_outputs(2061) <= not (a and b);
    layer2_outputs(2062) <= a and b;
    layer2_outputs(2063) <= b;
    layer2_outputs(2064) <= not (a and b);
    layer2_outputs(2065) <= b;
    layer2_outputs(2066) <= not (a xor b);
    layer2_outputs(2067) <= a and b;
    layer2_outputs(2068) <= a and b;
    layer2_outputs(2069) <= a and b;
    layer2_outputs(2070) <= a or b;
    layer2_outputs(2071) <= b and not a;
    layer2_outputs(2072) <= not (a and b);
    layer2_outputs(2073) <= b and not a;
    layer2_outputs(2074) <= a;
    layer2_outputs(2075) <= b;
    layer2_outputs(2076) <= b and not a;
    layer2_outputs(2077) <= not (a xor b);
    layer2_outputs(2078) <= a;
    layer2_outputs(2079) <= not a or b;
    layer2_outputs(2080) <= a xor b;
    layer2_outputs(2081) <= not a or b;
    layer2_outputs(2082) <= not (a or b);
    layer2_outputs(2083) <= not (a and b);
    layer2_outputs(2084) <= b;
    layer2_outputs(2085) <= b;
    layer2_outputs(2086) <= a;
    layer2_outputs(2087) <= not a;
    layer2_outputs(2088) <= not b;
    layer2_outputs(2089) <= a and b;
    layer2_outputs(2090) <= not (a and b);
    layer2_outputs(2091) <= a xor b;
    layer2_outputs(2092) <= not (a xor b);
    layer2_outputs(2093) <= not b or a;
    layer2_outputs(2094) <= a and not b;
    layer2_outputs(2095) <= not b;
    layer2_outputs(2096) <= a and not b;
    layer2_outputs(2097) <= not (a or b);
    layer2_outputs(2098) <= a and not b;
    layer2_outputs(2099) <= a and b;
    layer2_outputs(2100) <= a xor b;
    layer2_outputs(2101) <= not b or a;
    layer2_outputs(2102) <= not a or b;
    layer2_outputs(2103) <= not (a or b);
    layer2_outputs(2104) <= a;
    layer2_outputs(2105) <= a and b;
    layer2_outputs(2106) <= not (a xor b);
    layer2_outputs(2107) <= a and not b;
    layer2_outputs(2108) <= b;
    layer2_outputs(2109) <= b;
    layer2_outputs(2110) <= not a;
    layer2_outputs(2111) <= a or b;
    layer2_outputs(2112) <= a or b;
    layer2_outputs(2113) <= not b;
    layer2_outputs(2114) <= b;
    layer2_outputs(2115) <= not a;
    layer2_outputs(2116) <= a and b;
    layer2_outputs(2117) <= a and not b;
    layer2_outputs(2118) <= not (a xor b);
    layer2_outputs(2119) <= a;
    layer2_outputs(2120) <= 1'b1;
    layer2_outputs(2121) <= a xor b;
    layer2_outputs(2122) <= a and b;
    layer2_outputs(2123) <= not (a or b);
    layer2_outputs(2124) <= not a or b;
    layer2_outputs(2125) <= a xor b;
    layer2_outputs(2126) <= a;
    layer2_outputs(2127) <= not (a or b);
    layer2_outputs(2128) <= not (a or b);
    layer2_outputs(2129) <= not b;
    layer2_outputs(2130) <= not (a and b);
    layer2_outputs(2131) <= a and not b;
    layer2_outputs(2132) <= b;
    layer2_outputs(2133) <= a xor b;
    layer2_outputs(2134) <= a;
    layer2_outputs(2135) <= not (a or b);
    layer2_outputs(2136) <= a and b;
    layer2_outputs(2137) <= not b;
    layer2_outputs(2138) <= not a;
    layer2_outputs(2139) <= not b or a;
    layer2_outputs(2140) <= b;
    layer2_outputs(2141) <= not a or b;
    layer2_outputs(2142) <= a and b;
    layer2_outputs(2143) <= not b;
    layer2_outputs(2144) <= not (a or b);
    layer2_outputs(2145) <= a and not b;
    layer2_outputs(2146) <= a and b;
    layer2_outputs(2147) <= a;
    layer2_outputs(2148) <= a xor b;
    layer2_outputs(2149) <= not (a or b);
    layer2_outputs(2150) <= not a or b;
    layer2_outputs(2151) <= not a;
    layer2_outputs(2152) <= a;
    layer2_outputs(2153) <= a or b;
    layer2_outputs(2154) <= not a;
    layer2_outputs(2155) <= a and b;
    layer2_outputs(2156) <= a;
    layer2_outputs(2157) <= not a;
    layer2_outputs(2158) <= a xor b;
    layer2_outputs(2159) <= not a;
    layer2_outputs(2160) <= a or b;
    layer2_outputs(2161) <= 1'b1;
    layer2_outputs(2162) <= a and not b;
    layer2_outputs(2163) <= a or b;
    layer2_outputs(2164) <= not a;
    layer2_outputs(2165) <= not b or a;
    layer2_outputs(2166) <= a or b;
    layer2_outputs(2167) <= a and not b;
    layer2_outputs(2168) <= a and b;
    layer2_outputs(2169) <= not (a and b);
    layer2_outputs(2170) <= not b or a;
    layer2_outputs(2171) <= 1'b1;
    layer2_outputs(2172) <= not b or a;
    layer2_outputs(2173) <= a and b;
    layer2_outputs(2174) <= a;
    layer2_outputs(2175) <= not a or b;
    layer2_outputs(2176) <= b;
    layer2_outputs(2177) <= a and b;
    layer2_outputs(2178) <= a;
    layer2_outputs(2179) <= a and not b;
    layer2_outputs(2180) <= a or b;
    layer2_outputs(2181) <= a and b;
    layer2_outputs(2182) <= b and not a;
    layer2_outputs(2183) <= not (a or b);
    layer2_outputs(2184) <= a and b;
    layer2_outputs(2185) <= a xor b;
    layer2_outputs(2186) <= not b;
    layer2_outputs(2187) <= a;
    layer2_outputs(2188) <= not a;
    layer2_outputs(2189) <= a;
    layer2_outputs(2190) <= not a;
    layer2_outputs(2191) <= not b or a;
    layer2_outputs(2192) <= 1'b1;
    layer2_outputs(2193) <= a and not b;
    layer2_outputs(2194) <= not a;
    layer2_outputs(2195) <= not a;
    layer2_outputs(2196) <= not (a and b);
    layer2_outputs(2197) <= not b;
    layer2_outputs(2198) <= not (a and b);
    layer2_outputs(2199) <= not (a and b);
    layer2_outputs(2200) <= b;
    layer2_outputs(2201) <= a and b;
    layer2_outputs(2202) <= not b or a;
    layer2_outputs(2203) <= b and not a;
    layer2_outputs(2204) <= not (a or b);
    layer2_outputs(2205) <= not a;
    layer2_outputs(2206) <= a;
    layer2_outputs(2207) <= not a;
    layer2_outputs(2208) <= not (a or b);
    layer2_outputs(2209) <= a xor b;
    layer2_outputs(2210) <= not a;
    layer2_outputs(2211) <= not (a and b);
    layer2_outputs(2212) <= a or b;
    layer2_outputs(2213) <= not (a xor b);
    layer2_outputs(2214) <= a and not b;
    layer2_outputs(2215) <= a xor b;
    layer2_outputs(2216) <= a and b;
    layer2_outputs(2217) <= not b;
    layer2_outputs(2218) <= b and not a;
    layer2_outputs(2219) <= b and not a;
    layer2_outputs(2220) <= not a or b;
    layer2_outputs(2221) <= a;
    layer2_outputs(2222) <= b;
    layer2_outputs(2223) <= not b;
    layer2_outputs(2224) <= not b or a;
    layer2_outputs(2225) <= not (a or b);
    layer2_outputs(2226) <= b;
    layer2_outputs(2227) <= not (a and b);
    layer2_outputs(2228) <= not b;
    layer2_outputs(2229) <= a xor b;
    layer2_outputs(2230) <= a and not b;
    layer2_outputs(2231) <= not a;
    layer2_outputs(2232) <= a and b;
    layer2_outputs(2233) <= not a;
    layer2_outputs(2234) <= 1'b1;
    layer2_outputs(2235) <= b and not a;
    layer2_outputs(2236) <= b and not a;
    layer2_outputs(2237) <= a and b;
    layer2_outputs(2238) <= not (a or b);
    layer2_outputs(2239) <= not a;
    layer2_outputs(2240) <= not b;
    layer2_outputs(2241) <= a and not b;
    layer2_outputs(2242) <= a or b;
    layer2_outputs(2243) <= not b;
    layer2_outputs(2244) <= not (a xor b);
    layer2_outputs(2245) <= b;
    layer2_outputs(2246) <= b;
    layer2_outputs(2247) <= a;
    layer2_outputs(2248) <= a or b;
    layer2_outputs(2249) <= 1'b1;
    layer2_outputs(2250) <= a and not b;
    layer2_outputs(2251) <= not (a xor b);
    layer2_outputs(2252) <= a xor b;
    layer2_outputs(2253) <= a or b;
    layer2_outputs(2254) <= not a;
    layer2_outputs(2255) <= not (a or b);
    layer2_outputs(2256) <= not a;
    layer2_outputs(2257) <= not a or b;
    layer2_outputs(2258) <= not (a xor b);
    layer2_outputs(2259) <= a and b;
    layer2_outputs(2260) <= a xor b;
    layer2_outputs(2261) <= not a;
    layer2_outputs(2262) <= not a or b;
    layer2_outputs(2263) <= a xor b;
    layer2_outputs(2264) <= a;
    layer2_outputs(2265) <= not a or b;
    layer2_outputs(2266) <= a and not b;
    layer2_outputs(2267) <= a;
    layer2_outputs(2268) <= a xor b;
    layer2_outputs(2269) <= a;
    layer2_outputs(2270) <= a xor b;
    layer2_outputs(2271) <= not b;
    layer2_outputs(2272) <= a and not b;
    layer2_outputs(2273) <= not a;
    layer2_outputs(2274) <= not (a or b);
    layer2_outputs(2275) <= a or b;
    layer2_outputs(2276) <= not b;
    layer2_outputs(2277) <= a;
    layer2_outputs(2278) <= b;
    layer2_outputs(2279) <= not (a xor b);
    layer2_outputs(2280) <= b and not a;
    layer2_outputs(2281) <= not (a or b);
    layer2_outputs(2282) <= b and not a;
    layer2_outputs(2283) <= not (a or b);
    layer2_outputs(2284) <= a;
    layer2_outputs(2285) <= a and b;
    layer2_outputs(2286) <= not (a or b);
    layer2_outputs(2287) <= a and b;
    layer2_outputs(2288) <= not (a and b);
    layer2_outputs(2289) <= a and b;
    layer2_outputs(2290) <= b;
    layer2_outputs(2291) <= b;
    layer2_outputs(2292) <= not a or b;
    layer2_outputs(2293) <= a or b;
    layer2_outputs(2294) <= not (a or b);
    layer2_outputs(2295) <= not (a or b);
    layer2_outputs(2296) <= a and not b;
    layer2_outputs(2297) <= not (a and b);
    layer2_outputs(2298) <= not b;
    layer2_outputs(2299) <= a;
    layer2_outputs(2300) <= b;
    layer2_outputs(2301) <= a or b;
    layer2_outputs(2302) <= not (a xor b);
    layer2_outputs(2303) <= b and not a;
    layer2_outputs(2304) <= not a or b;
    layer2_outputs(2305) <= not (a and b);
    layer2_outputs(2306) <= b and not a;
    layer2_outputs(2307) <= b and not a;
    layer2_outputs(2308) <= not a;
    layer2_outputs(2309) <= a and not b;
    layer2_outputs(2310) <= b;
    layer2_outputs(2311) <= a;
    layer2_outputs(2312) <= b and not a;
    layer2_outputs(2313) <= a;
    layer2_outputs(2314) <= b and not a;
    layer2_outputs(2315) <= b and not a;
    layer2_outputs(2316) <= not (a or b);
    layer2_outputs(2317) <= not a;
    layer2_outputs(2318) <= a and b;
    layer2_outputs(2319) <= a or b;
    layer2_outputs(2320) <= not (a and b);
    layer2_outputs(2321) <= not b;
    layer2_outputs(2322) <= b;
    layer2_outputs(2323) <= not b;
    layer2_outputs(2324) <= not b or a;
    layer2_outputs(2325) <= a or b;
    layer2_outputs(2326) <= a;
    layer2_outputs(2327) <= not (a and b);
    layer2_outputs(2328) <= not b;
    layer2_outputs(2329) <= not a;
    layer2_outputs(2330) <= not b or a;
    layer2_outputs(2331) <= a and b;
    layer2_outputs(2332) <= b;
    layer2_outputs(2333) <= b and not a;
    layer2_outputs(2334) <= not (a xor b);
    layer2_outputs(2335) <= not (a or b);
    layer2_outputs(2336) <= a;
    layer2_outputs(2337) <= not b;
    layer2_outputs(2338) <= a or b;
    layer2_outputs(2339) <= not (a and b);
    layer2_outputs(2340) <= not b;
    layer2_outputs(2341) <= not (a xor b);
    layer2_outputs(2342) <= a xor b;
    layer2_outputs(2343) <= b;
    layer2_outputs(2344) <= b;
    layer2_outputs(2345) <= not (a or b);
    layer2_outputs(2346) <= a and b;
    layer2_outputs(2347) <= not a;
    layer2_outputs(2348) <= a and b;
    layer2_outputs(2349) <= not b;
    layer2_outputs(2350) <= not b or a;
    layer2_outputs(2351) <= not b;
    layer2_outputs(2352) <= not b;
    layer2_outputs(2353) <= a and not b;
    layer2_outputs(2354) <= a and not b;
    layer2_outputs(2355) <= a;
    layer2_outputs(2356) <= not (a or b);
    layer2_outputs(2357) <= b;
    layer2_outputs(2358) <= b and not a;
    layer2_outputs(2359) <= not (a or b);
    layer2_outputs(2360) <= not a;
    layer2_outputs(2361) <= a and b;
    layer2_outputs(2362) <= not a;
    layer2_outputs(2363) <= not b or a;
    layer2_outputs(2364) <= not a;
    layer2_outputs(2365) <= b and not a;
    layer2_outputs(2366) <= not (a and b);
    layer2_outputs(2367) <= not b or a;
    layer2_outputs(2368) <= not (a and b);
    layer2_outputs(2369) <= a;
    layer2_outputs(2370) <= not b;
    layer2_outputs(2371) <= a and not b;
    layer2_outputs(2372) <= not a or b;
    layer2_outputs(2373) <= not (a and b);
    layer2_outputs(2374) <= b and not a;
    layer2_outputs(2375) <= b;
    layer2_outputs(2376) <= b and not a;
    layer2_outputs(2377) <= not b or a;
    layer2_outputs(2378) <= not b;
    layer2_outputs(2379) <= a;
    layer2_outputs(2380) <= not (a xor b);
    layer2_outputs(2381) <= b;
    layer2_outputs(2382) <= not (a xor b);
    layer2_outputs(2383) <= not b or a;
    layer2_outputs(2384) <= not (a or b);
    layer2_outputs(2385) <= a and not b;
    layer2_outputs(2386) <= not a;
    layer2_outputs(2387) <= a and b;
    layer2_outputs(2388) <= not b or a;
    layer2_outputs(2389) <= not b;
    layer2_outputs(2390) <= a or b;
    layer2_outputs(2391) <= not b or a;
    layer2_outputs(2392) <= a or b;
    layer2_outputs(2393) <= b;
    layer2_outputs(2394) <= b and not a;
    layer2_outputs(2395) <= a and not b;
    layer2_outputs(2396) <= not (a and b);
    layer2_outputs(2397) <= a xor b;
    layer2_outputs(2398) <= a and not b;
    layer2_outputs(2399) <= not b;
    layer2_outputs(2400) <= a and b;
    layer2_outputs(2401) <= a;
    layer2_outputs(2402) <= a and b;
    layer2_outputs(2403) <= a and not b;
    layer2_outputs(2404) <= b;
    layer2_outputs(2405) <= b and not a;
    layer2_outputs(2406) <= not a;
    layer2_outputs(2407) <= not (a and b);
    layer2_outputs(2408) <= b and not a;
    layer2_outputs(2409) <= not b;
    layer2_outputs(2410) <= a;
    layer2_outputs(2411) <= a and not b;
    layer2_outputs(2412) <= b;
    layer2_outputs(2413) <= not b;
    layer2_outputs(2414) <= not a;
    layer2_outputs(2415) <= not (a or b);
    layer2_outputs(2416) <= not b;
    layer2_outputs(2417) <= a;
    layer2_outputs(2418) <= a and not b;
    layer2_outputs(2419) <= a and not b;
    layer2_outputs(2420) <= 1'b0;
    layer2_outputs(2421) <= not (a and b);
    layer2_outputs(2422) <= a xor b;
    layer2_outputs(2423) <= a or b;
    layer2_outputs(2424) <= a and b;
    layer2_outputs(2425) <= b;
    layer2_outputs(2426) <= b;
    layer2_outputs(2427) <= b and not a;
    layer2_outputs(2428) <= b;
    layer2_outputs(2429) <= a and not b;
    layer2_outputs(2430) <= a;
    layer2_outputs(2431) <= not a;
    layer2_outputs(2432) <= a and b;
    layer2_outputs(2433) <= not b or a;
    layer2_outputs(2434) <= not (a or b);
    layer2_outputs(2435) <= not a;
    layer2_outputs(2436) <= not a;
    layer2_outputs(2437) <= not b;
    layer2_outputs(2438) <= not (a xor b);
    layer2_outputs(2439) <= a or b;
    layer2_outputs(2440) <= not (a xor b);
    layer2_outputs(2441) <= a and b;
    layer2_outputs(2442) <= not a;
    layer2_outputs(2443) <= a and not b;
    layer2_outputs(2444) <= not a or b;
    layer2_outputs(2445) <= b;
    layer2_outputs(2446) <= 1'b1;
    layer2_outputs(2447) <= not b or a;
    layer2_outputs(2448) <= a xor b;
    layer2_outputs(2449) <= 1'b1;
    layer2_outputs(2450) <= b;
    layer2_outputs(2451) <= not (a and b);
    layer2_outputs(2452) <= a;
    layer2_outputs(2453) <= not (a xor b);
    layer2_outputs(2454) <= not b or a;
    layer2_outputs(2455) <= not b;
    layer2_outputs(2456) <= not (a and b);
    layer2_outputs(2457) <= a;
    layer2_outputs(2458) <= a;
    layer2_outputs(2459) <= a;
    layer2_outputs(2460) <= not a or b;
    layer2_outputs(2461) <= not b;
    layer2_outputs(2462) <= not a;
    layer2_outputs(2463) <= not b or a;
    layer2_outputs(2464) <= not (a and b);
    layer2_outputs(2465) <= b;
    layer2_outputs(2466) <= a;
    layer2_outputs(2467) <= a xor b;
    layer2_outputs(2468) <= a xor b;
    layer2_outputs(2469) <= a xor b;
    layer2_outputs(2470) <= not (a and b);
    layer2_outputs(2471) <= not a or b;
    layer2_outputs(2472) <= b and not a;
    layer2_outputs(2473) <= a;
    layer2_outputs(2474) <= not (a xor b);
    layer2_outputs(2475) <= not a;
    layer2_outputs(2476) <= not (a or b);
    layer2_outputs(2477) <= b;
    layer2_outputs(2478) <= a xor b;
    layer2_outputs(2479) <= not a;
    layer2_outputs(2480) <= a or b;
    layer2_outputs(2481) <= b;
    layer2_outputs(2482) <= not b;
    layer2_outputs(2483) <= not a;
    layer2_outputs(2484) <= not (a or b);
    layer2_outputs(2485) <= a and not b;
    layer2_outputs(2486) <= b;
    layer2_outputs(2487) <= a;
    layer2_outputs(2488) <= a;
    layer2_outputs(2489) <= a and not b;
    layer2_outputs(2490) <= a;
    layer2_outputs(2491) <= not b or a;
    layer2_outputs(2492) <= a xor b;
    layer2_outputs(2493) <= a;
    layer2_outputs(2494) <= b and not a;
    layer2_outputs(2495) <= not b;
    layer2_outputs(2496) <= not a;
    layer2_outputs(2497) <= a or b;
    layer2_outputs(2498) <= not a;
    layer2_outputs(2499) <= b and not a;
    layer2_outputs(2500) <= a;
    layer2_outputs(2501) <= not a;
    layer2_outputs(2502) <= b;
    layer2_outputs(2503) <= b;
    layer2_outputs(2504) <= not a or b;
    layer2_outputs(2505) <= a;
    layer2_outputs(2506) <= not b;
    layer2_outputs(2507) <= a and not b;
    layer2_outputs(2508) <= not a or b;
    layer2_outputs(2509) <= a xor b;
    layer2_outputs(2510) <= not b or a;
    layer2_outputs(2511) <= not a;
    layer2_outputs(2512) <= not a;
    layer2_outputs(2513) <= not a or b;
    layer2_outputs(2514) <= b;
    layer2_outputs(2515) <= not (a and b);
    layer2_outputs(2516) <= not b or a;
    layer2_outputs(2517) <= a;
    layer2_outputs(2518) <= b;
    layer2_outputs(2519) <= not (a and b);
    layer2_outputs(2520) <= not a or b;
    layer2_outputs(2521) <= not a;
    layer2_outputs(2522) <= not a or b;
    layer2_outputs(2523) <= not (a or b);
    layer2_outputs(2524) <= not b;
    layer2_outputs(2525) <= not a or b;
    layer2_outputs(2526) <= a and b;
    layer2_outputs(2527) <= b;
    layer2_outputs(2528) <= a or b;
    layer2_outputs(2529) <= a and not b;
    layer2_outputs(2530) <= not a or b;
    layer2_outputs(2531) <= b and not a;
    layer2_outputs(2532) <= not (a and b);
    layer2_outputs(2533) <= a and b;
    layer2_outputs(2534) <= not b;
    layer2_outputs(2535) <= not a;
    layer2_outputs(2536) <= b;
    layer2_outputs(2537) <= a;
    layer2_outputs(2538) <= not a or b;
    layer2_outputs(2539) <= a and b;
    layer2_outputs(2540) <= not b;
    layer2_outputs(2541) <= b;
    layer2_outputs(2542) <= a;
    layer2_outputs(2543) <= a and not b;
    layer2_outputs(2544) <= not a or b;
    layer2_outputs(2545) <= a and not b;
    layer2_outputs(2546) <= a and not b;
    layer2_outputs(2547) <= a;
    layer2_outputs(2548) <= b;
    layer2_outputs(2549) <= b and not a;
    layer2_outputs(2550) <= a and b;
    layer2_outputs(2551) <= a or b;
    layer2_outputs(2552) <= b and not a;
    layer2_outputs(2553) <= not a or b;
    layer2_outputs(2554) <= not (a xor b);
    layer2_outputs(2555) <= a or b;
    layer2_outputs(2556) <= a;
    layer2_outputs(2557) <= b;
    layer2_outputs(2558) <= not a;
    layer2_outputs(2559) <= a;
    layer2_outputs(2560) <= not a or b;
    layer2_outputs(2561) <= not b;
    layer2_outputs(2562) <= a or b;
    layer2_outputs(2563) <= not a or b;
    layer2_outputs(2564) <= a or b;
    layer2_outputs(2565) <= not a or b;
    layer2_outputs(2566) <= b and not a;
    layer2_outputs(2567) <= not (a or b);
    layer2_outputs(2568) <= a or b;
    layer2_outputs(2569) <= a and not b;
    layer2_outputs(2570) <= 1'b0;
    layer2_outputs(2571) <= not (a and b);
    layer2_outputs(2572) <= not a;
    layer2_outputs(2573) <= b;
    layer2_outputs(2574) <= not (a or b);
    layer2_outputs(2575) <= not (a xor b);
    layer2_outputs(2576) <= a or b;
    layer2_outputs(2577) <= not b or a;
    layer2_outputs(2578) <= a or b;
    layer2_outputs(2579) <= not (a xor b);
    layer2_outputs(2580) <= a or b;
    layer2_outputs(2581) <= b and not a;
    layer2_outputs(2582) <= not (a xor b);
    layer2_outputs(2583) <= not b;
    layer2_outputs(2584) <= a;
    layer2_outputs(2585) <= not (a or b);
    layer2_outputs(2586) <= not (a and b);
    layer2_outputs(2587) <= not a;
    layer2_outputs(2588) <= a and b;
    layer2_outputs(2589) <= not a;
    layer2_outputs(2590) <= a or b;
    layer2_outputs(2591) <= not a or b;
    layer2_outputs(2592) <= 1'b0;
    layer2_outputs(2593) <= not b or a;
    layer2_outputs(2594) <= not (a xor b);
    layer2_outputs(2595) <= not (a xor b);
    layer2_outputs(2596) <= a;
    layer2_outputs(2597) <= a xor b;
    layer2_outputs(2598) <= not a;
    layer2_outputs(2599) <= a or b;
    layer2_outputs(2600) <= not a;
    layer2_outputs(2601) <= a and b;
    layer2_outputs(2602) <= a;
    layer2_outputs(2603) <= not a;
    layer2_outputs(2604) <= 1'b0;
    layer2_outputs(2605) <= a and not b;
    layer2_outputs(2606) <= b;
    layer2_outputs(2607) <= a or b;
    layer2_outputs(2608) <= not b or a;
    layer2_outputs(2609) <= not a;
    layer2_outputs(2610) <= b;
    layer2_outputs(2611) <= not a;
    layer2_outputs(2612) <= not (a xor b);
    layer2_outputs(2613) <= not b or a;
    layer2_outputs(2614) <= b and not a;
    layer2_outputs(2615) <= not b;
    layer2_outputs(2616) <= not b;
    layer2_outputs(2617) <= a xor b;
    layer2_outputs(2618) <= b;
    layer2_outputs(2619) <= not (a or b);
    layer2_outputs(2620) <= a or b;
    layer2_outputs(2621) <= not (a or b);
    layer2_outputs(2622) <= b and not a;
    layer2_outputs(2623) <= not (a or b);
    layer2_outputs(2624) <= not (a xor b);
    layer2_outputs(2625) <= a and b;
    layer2_outputs(2626) <= not a or b;
    layer2_outputs(2627) <= b;
    layer2_outputs(2628) <= not a;
    layer2_outputs(2629) <= a xor b;
    layer2_outputs(2630) <= not (a xor b);
    layer2_outputs(2631) <= not (a and b);
    layer2_outputs(2632) <= not b or a;
    layer2_outputs(2633) <= not a;
    layer2_outputs(2634) <= a xor b;
    layer2_outputs(2635) <= a and b;
    layer2_outputs(2636) <= a and not b;
    layer2_outputs(2637) <= a;
    layer2_outputs(2638) <= not (a xor b);
    layer2_outputs(2639) <= a or b;
    layer2_outputs(2640) <= not a or b;
    layer2_outputs(2641) <= a and not b;
    layer2_outputs(2642) <= a and not b;
    layer2_outputs(2643) <= not a or b;
    layer2_outputs(2644) <= a and not b;
    layer2_outputs(2645) <= not (a xor b);
    layer2_outputs(2646) <= a;
    layer2_outputs(2647) <= not (a xor b);
    layer2_outputs(2648) <= not a;
    layer2_outputs(2649) <= b;
    layer2_outputs(2650) <= not a;
    layer2_outputs(2651) <= not (a and b);
    layer2_outputs(2652) <= not (a or b);
    layer2_outputs(2653) <= not a or b;
    layer2_outputs(2654) <= not b;
    layer2_outputs(2655) <= not b;
    layer2_outputs(2656) <= not b or a;
    layer2_outputs(2657) <= a and not b;
    layer2_outputs(2658) <= a and not b;
    layer2_outputs(2659) <= a;
    layer2_outputs(2660) <= not a;
    layer2_outputs(2661) <= not (a xor b);
    layer2_outputs(2662) <= not a;
    layer2_outputs(2663) <= not (a or b);
    layer2_outputs(2664) <= a;
    layer2_outputs(2665) <= b;
    layer2_outputs(2666) <= a;
    layer2_outputs(2667) <= not a;
    layer2_outputs(2668) <= not a;
    layer2_outputs(2669) <= a or b;
    layer2_outputs(2670) <= not a;
    layer2_outputs(2671) <= a;
    layer2_outputs(2672) <= not a;
    layer2_outputs(2673) <= not (a and b);
    layer2_outputs(2674) <= not a or b;
    layer2_outputs(2675) <= not (a or b);
    layer2_outputs(2676) <= not b or a;
    layer2_outputs(2677) <= not b;
    layer2_outputs(2678) <= a and b;
    layer2_outputs(2679) <= not a or b;
    layer2_outputs(2680) <= b and not a;
    layer2_outputs(2681) <= b;
    layer2_outputs(2682) <= not a;
    layer2_outputs(2683) <= not a;
    layer2_outputs(2684) <= not (a and b);
    layer2_outputs(2685) <= a or b;
    layer2_outputs(2686) <= a and not b;
    layer2_outputs(2687) <= not a;
    layer2_outputs(2688) <= 1'b1;
    layer2_outputs(2689) <= not (a xor b);
    layer2_outputs(2690) <= 1'b0;
    layer2_outputs(2691) <= a;
    layer2_outputs(2692) <= not a or b;
    layer2_outputs(2693) <= not (a or b);
    layer2_outputs(2694) <= a;
    layer2_outputs(2695) <= b;
    layer2_outputs(2696) <= a and not b;
    layer2_outputs(2697) <= b and not a;
    layer2_outputs(2698) <= not (a xor b);
    layer2_outputs(2699) <= b;
    layer2_outputs(2700) <= b and not a;
    layer2_outputs(2701) <= b and not a;
    layer2_outputs(2702) <= not b;
    layer2_outputs(2703) <= not a;
    layer2_outputs(2704) <= b and not a;
    layer2_outputs(2705) <= b;
    layer2_outputs(2706) <= not a;
    layer2_outputs(2707) <= b;
    layer2_outputs(2708) <= a xor b;
    layer2_outputs(2709) <= not (a and b);
    layer2_outputs(2710) <= a and not b;
    layer2_outputs(2711) <= b and not a;
    layer2_outputs(2712) <= b and not a;
    layer2_outputs(2713) <= a or b;
    layer2_outputs(2714) <= not (a and b);
    layer2_outputs(2715) <= a and not b;
    layer2_outputs(2716) <= a and not b;
    layer2_outputs(2717) <= a or b;
    layer2_outputs(2718) <= not a or b;
    layer2_outputs(2719) <= a xor b;
    layer2_outputs(2720) <= a;
    layer2_outputs(2721) <= a xor b;
    layer2_outputs(2722) <= not a;
    layer2_outputs(2723) <= not a or b;
    layer2_outputs(2724) <= not a or b;
    layer2_outputs(2725) <= not (a and b);
    layer2_outputs(2726) <= a and b;
    layer2_outputs(2727) <= not a;
    layer2_outputs(2728) <= a;
    layer2_outputs(2729) <= b and not a;
    layer2_outputs(2730) <= b and not a;
    layer2_outputs(2731) <= a;
    layer2_outputs(2732) <= not a;
    layer2_outputs(2733) <= not (a and b);
    layer2_outputs(2734) <= not b;
    layer2_outputs(2735) <= a or b;
    layer2_outputs(2736) <= b and not a;
    layer2_outputs(2737) <= a or b;
    layer2_outputs(2738) <= not a or b;
    layer2_outputs(2739) <= b;
    layer2_outputs(2740) <= not a;
    layer2_outputs(2741) <= not (a xor b);
    layer2_outputs(2742) <= not b or a;
    layer2_outputs(2743) <= a;
    layer2_outputs(2744) <= not (a or b);
    layer2_outputs(2745) <= a or b;
    layer2_outputs(2746) <= a xor b;
    layer2_outputs(2747) <= a and not b;
    layer2_outputs(2748) <= not b;
    layer2_outputs(2749) <= not b or a;
    layer2_outputs(2750) <= a and not b;
    layer2_outputs(2751) <= not (a xor b);
    layer2_outputs(2752) <= not b or a;
    layer2_outputs(2753) <= not a;
    layer2_outputs(2754) <= not a;
    layer2_outputs(2755) <= not a or b;
    layer2_outputs(2756) <= b;
    layer2_outputs(2757) <= not (a or b);
    layer2_outputs(2758) <= a and b;
    layer2_outputs(2759) <= not a or b;
    layer2_outputs(2760) <= b;
    layer2_outputs(2761) <= a xor b;
    layer2_outputs(2762) <= a;
    layer2_outputs(2763) <= a xor b;
    layer2_outputs(2764) <= a xor b;
    layer2_outputs(2765) <= not a;
    layer2_outputs(2766) <= b;
    layer2_outputs(2767) <= not b;
    layer2_outputs(2768) <= not b;
    layer2_outputs(2769) <= not (a xor b);
    layer2_outputs(2770) <= b;
    layer2_outputs(2771) <= not (a xor b);
    layer2_outputs(2772) <= a or b;
    layer2_outputs(2773) <= b and not a;
    layer2_outputs(2774) <= b;
    layer2_outputs(2775) <= a;
    layer2_outputs(2776) <= a or b;
    layer2_outputs(2777) <= a and not b;
    layer2_outputs(2778) <= not b;
    layer2_outputs(2779) <= not (a xor b);
    layer2_outputs(2780) <= a xor b;
    layer2_outputs(2781) <= b;
    layer2_outputs(2782) <= a xor b;
    layer2_outputs(2783) <= a and b;
    layer2_outputs(2784) <= a;
    layer2_outputs(2785) <= b;
    layer2_outputs(2786) <= a or b;
    layer2_outputs(2787) <= b;
    layer2_outputs(2788) <= a and not b;
    layer2_outputs(2789) <= b;
    layer2_outputs(2790) <= a xor b;
    layer2_outputs(2791) <= not a or b;
    layer2_outputs(2792) <= b and not a;
    layer2_outputs(2793) <= b and not a;
    layer2_outputs(2794) <= not (a and b);
    layer2_outputs(2795) <= a and b;
    layer2_outputs(2796) <= not a or b;
    layer2_outputs(2797) <= a xor b;
    layer2_outputs(2798) <= not a or b;
    layer2_outputs(2799) <= a or b;
    layer2_outputs(2800) <= not b;
    layer2_outputs(2801) <= not (a xor b);
    layer2_outputs(2802) <= b;
    layer2_outputs(2803) <= not a;
    layer2_outputs(2804) <= not (a xor b);
    layer2_outputs(2805) <= not b;
    layer2_outputs(2806) <= not a;
    layer2_outputs(2807) <= not (a or b);
    layer2_outputs(2808) <= a;
    layer2_outputs(2809) <= not b or a;
    layer2_outputs(2810) <= a xor b;
    layer2_outputs(2811) <= a;
    layer2_outputs(2812) <= not b;
    layer2_outputs(2813) <= not (a and b);
    layer2_outputs(2814) <= not (a or b);
    layer2_outputs(2815) <= a and not b;
    layer2_outputs(2816) <= a;
    layer2_outputs(2817) <= a;
    layer2_outputs(2818) <= a and b;
    layer2_outputs(2819) <= b;
    layer2_outputs(2820) <= not b or a;
    layer2_outputs(2821) <= not (a xor b);
    layer2_outputs(2822) <= not (a and b);
    layer2_outputs(2823) <= a xor b;
    layer2_outputs(2824) <= not (a and b);
    layer2_outputs(2825) <= not (a or b);
    layer2_outputs(2826) <= not a;
    layer2_outputs(2827) <= not (a or b);
    layer2_outputs(2828) <= not (a and b);
    layer2_outputs(2829) <= not a;
    layer2_outputs(2830) <= not a;
    layer2_outputs(2831) <= not b or a;
    layer2_outputs(2832) <= not b;
    layer2_outputs(2833) <= a or b;
    layer2_outputs(2834) <= not a;
    layer2_outputs(2835) <= b;
    layer2_outputs(2836) <= a or b;
    layer2_outputs(2837) <= a xor b;
    layer2_outputs(2838) <= not b or a;
    layer2_outputs(2839) <= 1'b0;
    layer2_outputs(2840) <= not a;
    layer2_outputs(2841) <= a;
    layer2_outputs(2842) <= not a;
    layer2_outputs(2843) <= a and not b;
    layer2_outputs(2844) <= b;
    layer2_outputs(2845) <= not a;
    layer2_outputs(2846) <= not b;
    layer2_outputs(2847) <= not (a or b);
    layer2_outputs(2848) <= a xor b;
    layer2_outputs(2849) <= not (a xor b);
    layer2_outputs(2850) <= b;
    layer2_outputs(2851) <= b;
    layer2_outputs(2852) <= b;
    layer2_outputs(2853) <= a;
    layer2_outputs(2854) <= not (a and b);
    layer2_outputs(2855) <= b;
    layer2_outputs(2856) <= not b;
    layer2_outputs(2857) <= not (a xor b);
    layer2_outputs(2858) <= not b;
    layer2_outputs(2859) <= b;
    layer2_outputs(2860) <= b and not a;
    layer2_outputs(2861) <= a or b;
    layer2_outputs(2862) <= b and not a;
    layer2_outputs(2863) <= not (a and b);
    layer2_outputs(2864) <= not b;
    layer2_outputs(2865) <= not a or b;
    layer2_outputs(2866) <= not b;
    layer2_outputs(2867) <= not b or a;
    layer2_outputs(2868) <= not (a xor b);
    layer2_outputs(2869) <= a or b;
    layer2_outputs(2870) <= not (a or b);
    layer2_outputs(2871) <= not b;
    layer2_outputs(2872) <= b;
    layer2_outputs(2873) <= a or b;
    layer2_outputs(2874) <= not (a xor b);
    layer2_outputs(2875) <= 1'b0;
    layer2_outputs(2876) <= a and b;
    layer2_outputs(2877) <= not (a or b);
    layer2_outputs(2878) <= not a;
    layer2_outputs(2879) <= not b;
    layer2_outputs(2880) <= not (a and b);
    layer2_outputs(2881) <= not a;
    layer2_outputs(2882) <= a or b;
    layer2_outputs(2883) <= not b;
    layer2_outputs(2884) <= a and b;
    layer2_outputs(2885) <= a;
    layer2_outputs(2886) <= a and b;
    layer2_outputs(2887) <= a;
    layer2_outputs(2888) <= a and b;
    layer2_outputs(2889) <= not (a xor b);
    layer2_outputs(2890) <= not a or b;
    layer2_outputs(2891) <= not (a xor b);
    layer2_outputs(2892) <= b;
    layer2_outputs(2893) <= not (a and b);
    layer2_outputs(2894) <= not b;
    layer2_outputs(2895) <= b;
    layer2_outputs(2896) <= a;
    layer2_outputs(2897) <= b;
    layer2_outputs(2898) <= not (a and b);
    layer2_outputs(2899) <= not a;
    layer2_outputs(2900) <= a and not b;
    layer2_outputs(2901) <= a and not b;
    layer2_outputs(2902) <= not (a xor b);
    layer2_outputs(2903) <= b;
    layer2_outputs(2904) <= a and b;
    layer2_outputs(2905) <= a or b;
    layer2_outputs(2906) <= a;
    layer2_outputs(2907) <= a or b;
    layer2_outputs(2908) <= not a;
    layer2_outputs(2909) <= a and b;
    layer2_outputs(2910) <= not a;
    layer2_outputs(2911) <= not b or a;
    layer2_outputs(2912) <= not b or a;
    layer2_outputs(2913) <= not b;
    layer2_outputs(2914) <= not (a and b);
    layer2_outputs(2915) <= a;
    layer2_outputs(2916) <= not b;
    layer2_outputs(2917) <= b;
    layer2_outputs(2918) <= not a or b;
    layer2_outputs(2919) <= b and not a;
    layer2_outputs(2920) <= not b;
    layer2_outputs(2921) <= not b;
    layer2_outputs(2922) <= b;
    layer2_outputs(2923) <= not b;
    layer2_outputs(2924) <= not b;
    layer2_outputs(2925) <= b;
    layer2_outputs(2926) <= b;
    layer2_outputs(2927) <= not b;
    layer2_outputs(2928) <= not b;
    layer2_outputs(2929) <= a xor b;
    layer2_outputs(2930) <= a and b;
    layer2_outputs(2931) <= not b;
    layer2_outputs(2932) <= not b or a;
    layer2_outputs(2933) <= not (a xor b);
    layer2_outputs(2934) <= not (a or b);
    layer2_outputs(2935) <= a and not b;
    layer2_outputs(2936) <= not a;
    layer2_outputs(2937) <= a and not b;
    layer2_outputs(2938) <= not b;
    layer2_outputs(2939) <= a xor b;
    layer2_outputs(2940) <= not b;
    layer2_outputs(2941) <= a or b;
    layer2_outputs(2942) <= a or b;
    layer2_outputs(2943) <= a and not b;
    layer2_outputs(2944) <= not a;
    layer2_outputs(2945) <= a and not b;
    layer2_outputs(2946) <= not (a xor b);
    layer2_outputs(2947) <= a and not b;
    layer2_outputs(2948) <= b;
    layer2_outputs(2949) <= b;
    layer2_outputs(2950) <= not (a xor b);
    layer2_outputs(2951) <= a and not b;
    layer2_outputs(2952) <= not a;
    layer2_outputs(2953) <= a and not b;
    layer2_outputs(2954) <= not b or a;
    layer2_outputs(2955) <= b and not a;
    layer2_outputs(2956) <= a;
    layer2_outputs(2957) <= a and b;
    layer2_outputs(2958) <= not (a xor b);
    layer2_outputs(2959) <= not (a xor b);
    layer2_outputs(2960) <= not b or a;
    layer2_outputs(2961) <= not b;
    layer2_outputs(2962) <= not a;
    layer2_outputs(2963) <= 1'b1;
    layer2_outputs(2964) <= b and not a;
    layer2_outputs(2965) <= a or b;
    layer2_outputs(2966) <= a;
    layer2_outputs(2967) <= not b;
    layer2_outputs(2968) <= a and b;
    layer2_outputs(2969) <= a and b;
    layer2_outputs(2970) <= a xor b;
    layer2_outputs(2971) <= b;
    layer2_outputs(2972) <= a and b;
    layer2_outputs(2973) <= 1'b0;
    layer2_outputs(2974) <= not a;
    layer2_outputs(2975) <= a;
    layer2_outputs(2976) <= not b or a;
    layer2_outputs(2977) <= not a;
    layer2_outputs(2978) <= not b or a;
    layer2_outputs(2979) <= b;
    layer2_outputs(2980) <= not b or a;
    layer2_outputs(2981) <= b;
    layer2_outputs(2982) <= b and not a;
    layer2_outputs(2983) <= b and not a;
    layer2_outputs(2984) <= a and b;
    layer2_outputs(2985) <= not b or a;
    layer2_outputs(2986) <= b;
    layer2_outputs(2987) <= b;
    layer2_outputs(2988) <= a and not b;
    layer2_outputs(2989) <= b;
    layer2_outputs(2990) <= a;
    layer2_outputs(2991) <= not (a xor b);
    layer2_outputs(2992) <= a;
    layer2_outputs(2993) <= not b;
    layer2_outputs(2994) <= b;
    layer2_outputs(2995) <= not b;
    layer2_outputs(2996) <= not b or a;
    layer2_outputs(2997) <= not (a xor b);
    layer2_outputs(2998) <= not b or a;
    layer2_outputs(2999) <= not a;
    layer2_outputs(3000) <= b;
    layer2_outputs(3001) <= a and b;
    layer2_outputs(3002) <= not (a or b);
    layer2_outputs(3003) <= b;
    layer2_outputs(3004) <= not (a and b);
    layer2_outputs(3005) <= not (a or b);
    layer2_outputs(3006) <= a and not b;
    layer2_outputs(3007) <= not (a and b);
    layer2_outputs(3008) <= a;
    layer2_outputs(3009) <= a or b;
    layer2_outputs(3010) <= not b or a;
    layer2_outputs(3011) <= b;
    layer2_outputs(3012) <= not b;
    layer2_outputs(3013) <= a xor b;
    layer2_outputs(3014) <= not b;
    layer2_outputs(3015) <= a;
    layer2_outputs(3016) <= a;
    layer2_outputs(3017) <= a and b;
    layer2_outputs(3018) <= not (a xor b);
    layer2_outputs(3019) <= not a;
    layer2_outputs(3020) <= not a;
    layer2_outputs(3021) <= not a;
    layer2_outputs(3022) <= not a;
    layer2_outputs(3023) <= not b;
    layer2_outputs(3024) <= a and b;
    layer2_outputs(3025) <= not b or a;
    layer2_outputs(3026) <= not a;
    layer2_outputs(3027) <= 1'b0;
    layer2_outputs(3028) <= not (a or b);
    layer2_outputs(3029) <= a or b;
    layer2_outputs(3030) <= b;
    layer2_outputs(3031) <= not (a or b);
    layer2_outputs(3032) <= not (a and b);
    layer2_outputs(3033) <= not (a xor b);
    layer2_outputs(3034) <= not (a or b);
    layer2_outputs(3035) <= a;
    layer2_outputs(3036) <= not (a or b);
    layer2_outputs(3037) <= a and b;
    layer2_outputs(3038) <= a;
    layer2_outputs(3039) <= a and not b;
    layer2_outputs(3040) <= b;
    layer2_outputs(3041) <= a and not b;
    layer2_outputs(3042) <= a and b;
    layer2_outputs(3043) <= a xor b;
    layer2_outputs(3044) <= not (a xor b);
    layer2_outputs(3045) <= a xor b;
    layer2_outputs(3046) <= not a;
    layer2_outputs(3047) <= not b;
    layer2_outputs(3048) <= not (a xor b);
    layer2_outputs(3049) <= a;
    layer2_outputs(3050) <= b;
    layer2_outputs(3051) <= not b;
    layer2_outputs(3052) <= not a or b;
    layer2_outputs(3053) <= b;
    layer2_outputs(3054) <= a and not b;
    layer2_outputs(3055) <= not a or b;
    layer2_outputs(3056) <= a;
    layer2_outputs(3057) <= a xor b;
    layer2_outputs(3058) <= b;
    layer2_outputs(3059) <= not b;
    layer2_outputs(3060) <= not b;
    layer2_outputs(3061) <= a and not b;
    layer2_outputs(3062) <= a and b;
    layer2_outputs(3063) <= b and not a;
    layer2_outputs(3064) <= not (a or b);
    layer2_outputs(3065) <= not b;
    layer2_outputs(3066) <= b;
    layer2_outputs(3067) <= b;
    layer2_outputs(3068) <= a xor b;
    layer2_outputs(3069) <= a;
    layer2_outputs(3070) <= not a;
    layer2_outputs(3071) <= a xor b;
    layer2_outputs(3072) <= not a or b;
    layer2_outputs(3073) <= a and not b;
    layer2_outputs(3074) <= not b;
    layer2_outputs(3075) <= b;
    layer2_outputs(3076) <= not b or a;
    layer2_outputs(3077) <= a and not b;
    layer2_outputs(3078) <= not b or a;
    layer2_outputs(3079) <= a;
    layer2_outputs(3080) <= a xor b;
    layer2_outputs(3081) <= a or b;
    layer2_outputs(3082) <= a and not b;
    layer2_outputs(3083) <= not b;
    layer2_outputs(3084) <= a;
    layer2_outputs(3085) <= a and b;
    layer2_outputs(3086) <= b;
    layer2_outputs(3087) <= not a;
    layer2_outputs(3088) <= a or b;
    layer2_outputs(3089) <= not b;
    layer2_outputs(3090) <= b;
    layer2_outputs(3091) <= b and not a;
    layer2_outputs(3092) <= not a;
    layer2_outputs(3093) <= a and not b;
    layer2_outputs(3094) <= not a or b;
    layer2_outputs(3095) <= a and not b;
    layer2_outputs(3096) <= not a;
    layer2_outputs(3097) <= not (a and b);
    layer2_outputs(3098) <= a xor b;
    layer2_outputs(3099) <= not a;
    layer2_outputs(3100) <= a and not b;
    layer2_outputs(3101) <= not b or a;
    layer2_outputs(3102) <= b;
    layer2_outputs(3103) <= a and b;
    layer2_outputs(3104) <= not (a or b);
    layer2_outputs(3105) <= not a;
    layer2_outputs(3106) <= b and not a;
    layer2_outputs(3107) <= a xor b;
    layer2_outputs(3108) <= a and b;
    layer2_outputs(3109) <= not a or b;
    layer2_outputs(3110) <= a;
    layer2_outputs(3111) <= not b;
    layer2_outputs(3112) <= b;
    layer2_outputs(3113) <= b;
    layer2_outputs(3114) <= not (a and b);
    layer2_outputs(3115) <= a;
    layer2_outputs(3116) <= not (a and b);
    layer2_outputs(3117) <= a xor b;
    layer2_outputs(3118) <= a;
    layer2_outputs(3119) <= a and b;
    layer2_outputs(3120) <= not (a or b);
    layer2_outputs(3121) <= a and b;
    layer2_outputs(3122) <= a xor b;
    layer2_outputs(3123) <= b;
    layer2_outputs(3124) <= a;
    layer2_outputs(3125) <= not (a xor b);
    layer2_outputs(3126) <= a;
    layer2_outputs(3127) <= b;
    layer2_outputs(3128) <= not b or a;
    layer2_outputs(3129) <= not (a or b);
    layer2_outputs(3130) <= not b;
    layer2_outputs(3131) <= not b;
    layer2_outputs(3132) <= a;
    layer2_outputs(3133) <= a;
    layer2_outputs(3134) <= a;
    layer2_outputs(3135) <= b;
    layer2_outputs(3136) <= not a;
    layer2_outputs(3137) <= 1'b1;
    layer2_outputs(3138) <= not b;
    layer2_outputs(3139) <= b and not a;
    layer2_outputs(3140) <= a;
    layer2_outputs(3141) <= not (a or b);
    layer2_outputs(3142) <= a xor b;
    layer2_outputs(3143) <= 1'b0;
    layer2_outputs(3144) <= not b or a;
    layer2_outputs(3145) <= not b;
    layer2_outputs(3146) <= a and not b;
    layer2_outputs(3147) <= a;
    layer2_outputs(3148) <= not b;
    layer2_outputs(3149) <= not (a or b);
    layer2_outputs(3150) <= not a;
    layer2_outputs(3151) <= not b;
    layer2_outputs(3152) <= not (a and b);
    layer2_outputs(3153) <= b;
    layer2_outputs(3154) <= not (a xor b);
    layer2_outputs(3155) <= not (a or b);
    layer2_outputs(3156) <= not (a or b);
    layer2_outputs(3157) <= not b;
    layer2_outputs(3158) <= a xor b;
    layer2_outputs(3159) <= not b or a;
    layer2_outputs(3160) <= not b;
    layer2_outputs(3161) <= a xor b;
    layer2_outputs(3162) <= not (a xor b);
    layer2_outputs(3163) <= not (a or b);
    layer2_outputs(3164) <= not a;
    layer2_outputs(3165) <= not a;
    layer2_outputs(3166) <= not (a or b);
    layer2_outputs(3167) <= not b or a;
    layer2_outputs(3168) <= a xor b;
    layer2_outputs(3169) <= a;
    layer2_outputs(3170) <= b;
    layer2_outputs(3171) <= a;
    layer2_outputs(3172) <= b;
    layer2_outputs(3173) <= not b;
    layer2_outputs(3174) <= a and not b;
    layer2_outputs(3175) <= b and not a;
    layer2_outputs(3176) <= a or b;
    layer2_outputs(3177) <= a xor b;
    layer2_outputs(3178) <= not a;
    layer2_outputs(3179) <= b;
    layer2_outputs(3180) <= b;
    layer2_outputs(3181) <= a and not b;
    layer2_outputs(3182) <= b and not a;
    layer2_outputs(3183) <= a;
    layer2_outputs(3184) <= b;
    layer2_outputs(3185) <= b;
    layer2_outputs(3186) <= not b or a;
    layer2_outputs(3187) <= not b or a;
    layer2_outputs(3188) <= not a;
    layer2_outputs(3189) <= not (a and b);
    layer2_outputs(3190) <= a and b;
    layer2_outputs(3191) <= 1'b1;
    layer2_outputs(3192) <= not b;
    layer2_outputs(3193) <= not (a xor b);
    layer2_outputs(3194) <= not (a and b);
    layer2_outputs(3195) <= not (a or b);
    layer2_outputs(3196) <= not b;
    layer2_outputs(3197) <= b;
    layer2_outputs(3198) <= a;
    layer2_outputs(3199) <= not b;
    layer2_outputs(3200) <= a;
    layer2_outputs(3201) <= b;
    layer2_outputs(3202) <= b and not a;
    layer2_outputs(3203) <= a xor b;
    layer2_outputs(3204) <= not a or b;
    layer2_outputs(3205) <= a;
    layer2_outputs(3206) <= a and not b;
    layer2_outputs(3207) <= b;
    layer2_outputs(3208) <= not b;
    layer2_outputs(3209) <= a;
    layer2_outputs(3210) <= a or b;
    layer2_outputs(3211) <= not a or b;
    layer2_outputs(3212) <= a;
    layer2_outputs(3213) <= not (a and b);
    layer2_outputs(3214) <= a and b;
    layer2_outputs(3215) <= a and not b;
    layer2_outputs(3216) <= a;
    layer2_outputs(3217) <= a;
    layer2_outputs(3218) <= a and not b;
    layer2_outputs(3219) <= not b;
    layer2_outputs(3220) <= b and not a;
    layer2_outputs(3221) <= a or b;
    layer2_outputs(3222) <= a and b;
    layer2_outputs(3223) <= not (a xor b);
    layer2_outputs(3224) <= a xor b;
    layer2_outputs(3225) <= not (a and b);
    layer2_outputs(3226) <= 1'b0;
    layer2_outputs(3227) <= b;
    layer2_outputs(3228) <= not a;
    layer2_outputs(3229) <= b;
    layer2_outputs(3230) <= not b or a;
    layer2_outputs(3231) <= not a or b;
    layer2_outputs(3232) <= not (a or b);
    layer2_outputs(3233) <= not b or a;
    layer2_outputs(3234) <= a;
    layer2_outputs(3235) <= not a or b;
    layer2_outputs(3236) <= not (a and b);
    layer2_outputs(3237) <= a xor b;
    layer2_outputs(3238) <= a;
    layer2_outputs(3239) <= not a or b;
    layer2_outputs(3240) <= not a or b;
    layer2_outputs(3241) <= not a or b;
    layer2_outputs(3242) <= not a;
    layer2_outputs(3243) <= not b;
    layer2_outputs(3244) <= not (a and b);
    layer2_outputs(3245) <= a;
    layer2_outputs(3246) <= not (a or b);
    layer2_outputs(3247) <= not (a or b);
    layer2_outputs(3248) <= not (a or b);
    layer2_outputs(3249) <= a;
    layer2_outputs(3250) <= a;
    layer2_outputs(3251) <= a;
    layer2_outputs(3252) <= not a;
    layer2_outputs(3253) <= not b;
    layer2_outputs(3254) <= not a;
    layer2_outputs(3255) <= not (a and b);
    layer2_outputs(3256) <= a and not b;
    layer2_outputs(3257) <= a or b;
    layer2_outputs(3258) <= a and b;
    layer2_outputs(3259) <= not a;
    layer2_outputs(3260) <= a;
    layer2_outputs(3261) <= not a or b;
    layer2_outputs(3262) <= a or b;
    layer2_outputs(3263) <= not (a or b);
    layer2_outputs(3264) <= not (a xor b);
    layer2_outputs(3265) <= not (a xor b);
    layer2_outputs(3266) <= not b;
    layer2_outputs(3267) <= not b;
    layer2_outputs(3268) <= not b or a;
    layer2_outputs(3269) <= not b;
    layer2_outputs(3270) <= b and not a;
    layer2_outputs(3271) <= a or b;
    layer2_outputs(3272) <= a;
    layer2_outputs(3273) <= a;
    layer2_outputs(3274) <= a;
    layer2_outputs(3275) <= a and b;
    layer2_outputs(3276) <= not b;
    layer2_outputs(3277) <= not b or a;
    layer2_outputs(3278) <= not a;
    layer2_outputs(3279) <= a;
    layer2_outputs(3280) <= not b;
    layer2_outputs(3281) <= not (a xor b);
    layer2_outputs(3282) <= a;
    layer2_outputs(3283) <= not a;
    layer2_outputs(3284) <= a or b;
    layer2_outputs(3285) <= 1'b0;
    layer2_outputs(3286) <= not a;
    layer2_outputs(3287) <= not b;
    layer2_outputs(3288) <= b;
    layer2_outputs(3289) <= not a or b;
    layer2_outputs(3290) <= a and not b;
    layer2_outputs(3291) <= a xor b;
    layer2_outputs(3292) <= not (a or b);
    layer2_outputs(3293) <= not b;
    layer2_outputs(3294) <= a and not b;
    layer2_outputs(3295) <= 1'b0;
    layer2_outputs(3296) <= a and not b;
    layer2_outputs(3297) <= not a;
    layer2_outputs(3298) <= not a;
    layer2_outputs(3299) <= not (a xor b);
    layer2_outputs(3300) <= not (a and b);
    layer2_outputs(3301) <= a and b;
    layer2_outputs(3302) <= not b or a;
    layer2_outputs(3303) <= not (a and b);
    layer2_outputs(3304) <= not b;
    layer2_outputs(3305) <= a or b;
    layer2_outputs(3306) <= not a or b;
    layer2_outputs(3307) <= a or b;
    layer2_outputs(3308) <= b and not a;
    layer2_outputs(3309) <= not a or b;
    layer2_outputs(3310) <= a or b;
    layer2_outputs(3311) <= not (a or b);
    layer2_outputs(3312) <= a;
    layer2_outputs(3313) <= not a;
    layer2_outputs(3314) <= not (a xor b);
    layer2_outputs(3315) <= not (a and b);
    layer2_outputs(3316) <= a;
    layer2_outputs(3317) <= not a;
    layer2_outputs(3318) <= a xor b;
    layer2_outputs(3319) <= a and not b;
    layer2_outputs(3320) <= not b or a;
    layer2_outputs(3321) <= not a;
    layer2_outputs(3322) <= a or b;
    layer2_outputs(3323) <= not a;
    layer2_outputs(3324) <= not b or a;
    layer2_outputs(3325) <= a and not b;
    layer2_outputs(3326) <= b;
    layer2_outputs(3327) <= not (a or b);
    layer2_outputs(3328) <= not a;
    layer2_outputs(3329) <= a xor b;
    layer2_outputs(3330) <= not a or b;
    layer2_outputs(3331) <= a and b;
    layer2_outputs(3332) <= a and not b;
    layer2_outputs(3333) <= not a or b;
    layer2_outputs(3334) <= not b or a;
    layer2_outputs(3335) <= a and not b;
    layer2_outputs(3336) <= a xor b;
    layer2_outputs(3337) <= b and not a;
    layer2_outputs(3338) <= not a;
    layer2_outputs(3339) <= not (a xor b);
    layer2_outputs(3340) <= not (a and b);
    layer2_outputs(3341) <= a;
    layer2_outputs(3342) <= a;
    layer2_outputs(3343) <= b;
    layer2_outputs(3344) <= b;
    layer2_outputs(3345) <= not (a and b);
    layer2_outputs(3346) <= not a or b;
    layer2_outputs(3347) <= a xor b;
    layer2_outputs(3348) <= a and b;
    layer2_outputs(3349) <= not a;
    layer2_outputs(3350) <= a or b;
    layer2_outputs(3351) <= a;
    layer2_outputs(3352) <= a and not b;
    layer2_outputs(3353) <= not b or a;
    layer2_outputs(3354) <= a or b;
    layer2_outputs(3355) <= a and b;
    layer2_outputs(3356) <= not a;
    layer2_outputs(3357) <= a and not b;
    layer2_outputs(3358) <= a and not b;
    layer2_outputs(3359) <= b;
    layer2_outputs(3360) <= a and b;
    layer2_outputs(3361) <= not a;
    layer2_outputs(3362) <= a xor b;
    layer2_outputs(3363) <= a or b;
    layer2_outputs(3364) <= not a or b;
    layer2_outputs(3365) <= not a;
    layer2_outputs(3366) <= not b;
    layer2_outputs(3367) <= not (a and b);
    layer2_outputs(3368) <= not b or a;
    layer2_outputs(3369) <= not a or b;
    layer2_outputs(3370) <= b;
    layer2_outputs(3371) <= a;
    layer2_outputs(3372) <= not b;
    layer2_outputs(3373) <= b and not a;
    layer2_outputs(3374) <= b and not a;
    layer2_outputs(3375) <= a;
    layer2_outputs(3376) <= b;
    layer2_outputs(3377) <= a;
    layer2_outputs(3378) <= b;
    layer2_outputs(3379) <= not a;
    layer2_outputs(3380) <= a xor b;
    layer2_outputs(3381) <= not b;
    layer2_outputs(3382) <= a;
    layer2_outputs(3383) <= a or b;
    layer2_outputs(3384) <= not b;
    layer2_outputs(3385) <= b;
    layer2_outputs(3386) <= a xor b;
    layer2_outputs(3387) <= not (a and b);
    layer2_outputs(3388) <= not (a xor b);
    layer2_outputs(3389) <= b;
    layer2_outputs(3390) <= a;
    layer2_outputs(3391) <= not (a xor b);
    layer2_outputs(3392) <= a and b;
    layer2_outputs(3393) <= a or b;
    layer2_outputs(3394) <= not (a and b);
    layer2_outputs(3395) <= a and b;
    layer2_outputs(3396) <= a or b;
    layer2_outputs(3397) <= a and b;
    layer2_outputs(3398) <= b and not a;
    layer2_outputs(3399) <= not a or b;
    layer2_outputs(3400) <= not b;
    layer2_outputs(3401) <= a and b;
    layer2_outputs(3402) <= b;
    layer2_outputs(3403) <= not a;
    layer2_outputs(3404) <= a;
    layer2_outputs(3405) <= b and not a;
    layer2_outputs(3406) <= not a or b;
    layer2_outputs(3407) <= not b or a;
    layer2_outputs(3408) <= a xor b;
    layer2_outputs(3409) <= a and not b;
    layer2_outputs(3410) <= a;
    layer2_outputs(3411) <= not b or a;
    layer2_outputs(3412) <= not a or b;
    layer2_outputs(3413) <= not b or a;
    layer2_outputs(3414) <= not (a and b);
    layer2_outputs(3415) <= not a;
    layer2_outputs(3416) <= b;
    layer2_outputs(3417) <= not b or a;
    layer2_outputs(3418) <= a and not b;
    layer2_outputs(3419) <= a and b;
    layer2_outputs(3420) <= a xor b;
    layer2_outputs(3421) <= a xor b;
    layer2_outputs(3422) <= a or b;
    layer2_outputs(3423) <= a and not b;
    layer2_outputs(3424) <= a and not b;
    layer2_outputs(3425) <= a or b;
    layer2_outputs(3426) <= not b or a;
    layer2_outputs(3427) <= not a;
    layer2_outputs(3428) <= a xor b;
    layer2_outputs(3429) <= not (a and b);
    layer2_outputs(3430) <= b;
    layer2_outputs(3431) <= not (a and b);
    layer2_outputs(3432) <= not (a and b);
    layer2_outputs(3433) <= not (a and b);
    layer2_outputs(3434) <= a and b;
    layer2_outputs(3435) <= a xor b;
    layer2_outputs(3436) <= b;
    layer2_outputs(3437) <= not b or a;
    layer2_outputs(3438) <= not a or b;
    layer2_outputs(3439) <= a and not b;
    layer2_outputs(3440) <= a and not b;
    layer2_outputs(3441) <= not (a xor b);
    layer2_outputs(3442) <= a;
    layer2_outputs(3443) <= not a;
    layer2_outputs(3444) <= not b;
    layer2_outputs(3445) <= not b or a;
    layer2_outputs(3446) <= not (a xor b);
    layer2_outputs(3447) <= a;
    layer2_outputs(3448) <= not a or b;
    layer2_outputs(3449) <= b;
    layer2_outputs(3450) <= not b or a;
    layer2_outputs(3451) <= b;
    layer2_outputs(3452) <= a or b;
    layer2_outputs(3453) <= not b;
    layer2_outputs(3454) <= b;
    layer2_outputs(3455) <= b;
    layer2_outputs(3456) <= b;
    layer2_outputs(3457) <= b and not a;
    layer2_outputs(3458) <= not a or b;
    layer2_outputs(3459) <= a;
    layer2_outputs(3460) <= not a or b;
    layer2_outputs(3461) <= b;
    layer2_outputs(3462) <= not (a xor b);
    layer2_outputs(3463) <= 1'b0;
    layer2_outputs(3464) <= not a;
    layer2_outputs(3465) <= b and not a;
    layer2_outputs(3466) <= not (a or b);
    layer2_outputs(3467) <= a and not b;
    layer2_outputs(3468) <= a;
    layer2_outputs(3469) <= a and not b;
    layer2_outputs(3470) <= b;
    layer2_outputs(3471) <= not b or a;
    layer2_outputs(3472) <= a or b;
    layer2_outputs(3473) <= 1'b1;
    layer2_outputs(3474) <= not a;
    layer2_outputs(3475) <= not b;
    layer2_outputs(3476) <= not a or b;
    layer2_outputs(3477) <= not a or b;
    layer2_outputs(3478) <= a or b;
    layer2_outputs(3479) <= not a or b;
    layer2_outputs(3480) <= not a;
    layer2_outputs(3481) <= a and not b;
    layer2_outputs(3482) <= b and not a;
    layer2_outputs(3483) <= not (a and b);
    layer2_outputs(3484) <= not b;
    layer2_outputs(3485) <= not (a or b);
    layer2_outputs(3486) <= not a;
    layer2_outputs(3487) <= not (a or b);
    layer2_outputs(3488) <= a xor b;
    layer2_outputs(3489) <= not b;
    layer2_outputs(3490) <= not a;
    layer2_outputs(3491) <= not (a xor b);
    layer2_outputs(3492) <= not (a or b);
    layer2_outputs(3493) <= b;
    layer2_outputs(3494) <= not a or b;
    layer2_outputs(3495) <= a;
    layer2_outputs(3496) <= not (a or b);
    layer2_outputs(3497) <= b and not a;
    layer2_outputs(3498) <= a or b;
    layer2_outputs(3499) <= b;
    layer2_outputs(3500) <= a or b;
    layer2_outputs(3501) <= not b;
    layer2_outputs(3502) <= a and b;
    layer2_outputs(3503) <= not (a xor b);
    layer2_outputs(3504) <= not (a or b);
    layer2_outputs(3505) <= not (a or b);
    layer2_outputs(3506) <= not (a and b);
    layer2_outputs(3507) <= not a;
    layer2_outputs(3508) <= not a or b;
    layer2_outputs(3509) <= a and b;
    layer2_outputs(3510) <= not a;
    layer2_outputs(3511) <= not b;
    layer2_outputs(3512) <= a;
    layer2_outputs(3513) <= a xor b;
    layer2_outputs(3514) <= b and not a;
    layer2_outputs(3515) <= not b;
    layer2_outputs(3516) <= not b or a;
    layer2_outputs(3517) <= b and not a;
    layer2_outputs(3518) <= not (a and b);
    layer2_outputs(3519) <= a;
    layer2_outputs(3520) <= not (a and b);
    layer2_outputs(3521) <= a and not b;
    layer2_outputs(3522) <= b;
    layer2_outputs(3523) <= a and b;
    layer2_outputs(3524) <= b;
    layer2_outputs(3525) <= not a;
    layer2_outputs(3526) <= not a;
    layer2_outputs(3527) <= not b or a;
    layer2_outputs(3528) <= b;
    layer2_outputs(3529) <= not (a or b);
    layer2_outputs(3530) <= not b;
    layer2_outputs(3531) <= not (a and b);
    layer2_outputs(3532) <= not (a xor b);
    layer2_outputs(3533) <= b;
    layer2_outputs(3534) <= a;
    layer2_outputs(3535) <= not b;
    layer2_outputs(3536) <= b;
    layer2_outputs(3537) <= not a or b;
    layer2_outputs(3538) <= b and not a;
    layer2_outputs(3539) <= not (a xor b);
    layer2_outputs(3540) <= b;
    layer2_outputs(3541) <= not b or a;
    layer2_outputs(3542) <= a;
    layer2_outputs(3543) <= not b or a;
    layer2_outputs(3544) <= not b;
    layer2_outputs(3545) <= b;
    layer2_outputs(3546) <= a and b;
    layer2_outputs(3547) <= a;
    layer2_outputs(3548) <= a and b;
    layer2_outputs(3549) <= a;
    layer2_outputs(3550) <= a;
    layer2_outputs(3551) <= not a or b;
    layer2_outputs(3552) <= a and not b;
    layer2_outputs(3553) <= b;
    layer2_outputs(3554) <= a xor b;
    layer2_outputs(3555) <= a or b;
    layer2_outputs(3556) <= not a or b;
    layer2_outputs(3557) <= a and b;
    layer2_outputs(3558) <= not b or a;
    layer2_outputs(3559) <= a and b;
    layer2_outputs(3560) <= b;
    layer2_outputs(3561) <= a;
    layer2_outputs(3562) <= a or b;
    layer2_outputs(3563) <= a or b;
    layer2_outputs(3564) <= not (a or b);
    layer2_outputs(3565) <= not b or a;
    layer2_outputs(3566) <= a or b;
    layer2_outputs(3567) <= not (a or b);
    layer2_outputs(3568) <= not (a xor b);
    layer2_outputs(3569) <= a or b;
    layer2_outputs(3570) <= b and not a;
    layer2_outputs(3571) <= not b or a;
    layer2_outputs(3572) <= a or b;
    layer2_outputs(3573) <= not (a xor b);
    layer2_outputs(3574) <= a and not b;
    layer2_outputs(3575) <= b;
    layer2_outputs(3576) <= not b or a;
    layer2_outputs(3577) <= b and not a;
    layer2_outputs(3578) <= b and not a;
    layer2_outputs(3579) <= not a or b;
    layer2_outputs(3580) <= b;
    layer2_outputs(3581) <= a and b;
    layer2_outputs(3582) <= b;
    layer2_outputs(3583) <= a or b;
    layer2_outputs(3584) <= b;
    layer2_outputs(3585) <= b and not a;
    layer2_outputs(3586) <= b and not a;
    layer2_outputs(3587) <= not a;
    layer2_outputs(3588) <= a or b;
    layer2_outputs(3589) <= not a or b;
    layer2_outputs(3590) <= a or b;
    layer2_outputs(3591) <= not (a xor b);
    layer2_outputs(3592) <= a;
    layer2_outputs(3593) <= not b or a;
    layer2_outputs(3594) <= not (a or b);
    layer2_outputs(3595) <= a xor b;
    layer2_outputs(3596) <= not b or a;
    layer2_outputs(3597) <= not a;
    layer2_outputs(3598) <= not (a and b);
    layer2_outputs(3599) <= not a or b;
    layer2_outputs(3600) <= not (a and b);
    layer2_outputs(3601) <= a and not b;
    layer2_outputs(3602) <= b and not a;
    layer2_outputs(3603) <= not (a or b);
    layer2_outputs(3604) <= a and b;
    layer2_outputs(3605) <= a;
    layer2_outputs(3606) <= a;
    layer2_outputs(3607) <= b;
    layer2_outputs(3608) <= a and b;
    layer2_outputs(3609) <= not b or a;
    layer2_outputs(3610) <= not b or a;
    layer2_outputs(3611) <= not (a and b);
    layer2_outputs(3612) <= b and not a;
    layer2_outputs(3613) <= not b or a;
    layer2_outputs(3614) <= not (a and b);
    layer2_outputs(3615) <= not a or b;
    layer2_outputs(3616) <= a;
    layer2_outputs(3617) <= not (a xor b);
    layer2_outputs(3618) <= not a;
    layer2_outputs(3619) <= not (a xor b);
    layer2_outputs(3620) <= not (a or b);
    layer2_outputs(3621) <= not a;
    layer2_outputs(3622) <= b and not a;
    layer2_outputs(3623) <= a;
    layer2_outputs(3624) <= a xor b;
    layer2_outputs(3625) <= not (a or b);
    layer2_outputs(3626) <= not a or b;
    layer2_outputs(3627) <= not a;
    layer2_outputs(3628) <= not b;
    layer2_outputs(3629) <= not (a or b);
    layer2_outputs(3630) <= a and not b;
    layer2_outputs(3631) <= not b;
    layer2_outputs(3632) <= a;
    layer2_outputs(3633) <= not (a and b);
    layer2_outputs(3634) <= not b;
    layer2_outputs(3635) <= b and not a;
    layer2_outputs(3636) <= not b;
    layer2_outputs(3637) <= not (a xor b);
    layer2_outputs(3638) <= not b;
    layer2_outputs(3639) <= not (a or b);
    layer2_outputs(3640) <= not a;
    layer2_outputs(3641) <= b;
    layer2_outputs(3642) <= not (a or b);
    layer2_outputs(3643) <= not b;
    layer2_outputs(3644) <= not (a or b);
    layer2_outputs(3645) <= not a or b;
    layer2_outputs(3646) <= not b;
    layer2_outputs(3647) <= not b or a;
    layer2_outputs(3648) <= not a;
    layer2_outputs(3649) <= not a or b;
    layer2_outputs(3650) <= b;
    layer2_outputs(3651) <= b;
    layer2_outputs(3652) <= not (a and b);
    layer2_outputs(3653) <= a or b;
    layer2_outputs(3654) <= not a or b;
    layer2_outputs(3655) <= not (a or b);
    layer2_outputs(3656) <= a;
    layer2_outputs(3657) <= 1'b1;
    layer2_outputs(3658) <= not (a or b);
    layer2_outputs(3659) <= b and not a;
    layer2_outputs(3660) <= not b;
    layer2_outputs(3661) <= not b;
    layer2_outputs(3662) <= a or b;
    layer2_outputs(3663) <= not (a xor b);
    layer2_outputs(3664) <= b;
    layer2_outputs(3665) <= a;
    layer2_outputs(3666) <= not (a or b);
    layer2_outputs(3667) <= not (a or b);
    layer2_outputs(3668) <= not (a xor b);
    layer2_outputs(3669) <= b;
    layer2_outputs(3670) <= a and not b;
    layer2_outputs(3671) <= a;
    layer2_outputs(3672) <= not a;
    layer2_outputs(3673) <= not (a and b);
    layer2_outputs(3674) <= not (a and b);
    layer2_outputs(3675) <= a and not b;
    layer2_outputs(3676) <= not (a or b);
    layer2_outputs(3677) <= a xor b;
    layer2_outputs(3678) <= not b or a;
    layer2_outputs(3679) <= a;
    layer2_outputs(3680) <= a or b;
    layer2_outputs(3681) <= b;
    layer2_outputs(3682) <= a and b;
    layer2_outputs(3683) <= a and b;
    layer2_outputs(3684) <= a xor b;
    layer2_outputs(3685) <= not (a or b);
    layer2_outputs(3686) <= not a;
    layer2_outputs(3687) <= not b;
    layer2_outputs(3688) <= not b or a;
    layer2_outputs(3689) <= a or b;
    layer2_outputs(3690) <= not (a or b);
    layer2_outputs(3691) <= not a;
    layer2_outputs(3692) <= not (a or b);
    layer2_outputs(3693) <= not (a and b);
    layer2_outputs(3694) <= b;
    layer2_outputs(3695) <= not b;
    layer2_outputs(3696) <= not b or a;
    layer2_outputs(3697) <= a;
    layer2_outputs(3698) <= a and not b;
    layer2_outputs(3699) <= a and b;
    layer2_outputs(3700) <= a or b;
    layer2_outputs(3701) <= not b or a;
    layer2_outputs(3702) <= not b;
    layer2_outputs(3703) <= not (a and b);
    layer2_outputs(3704) <= not (a xor b);
    layer2_outputs(3705) <= not b or a;
    layer2_outputs(3706) <= not (a or b);
    layer2_outputs(3707) <= not (a and b);
    layer2_outputs(3708) <= a xor b;
    layer2_outputs(3709) <= b;
    layer2_outputs(3710) <= not a;
    layer2_outputs(3711) <= a and not b;
    layer2_outputs(3712) <= b;
    layer2_outputs(3713) <= a;
    layer2_outputs(3714) <= not (a or b);
    layer2_outputs(3715) <= b;
    layer2_outputs(3716) <= not (a and b);
    layer2_outputs(3717) <= not (a or b);
    layer2_outputs(3718) <= not a;
    layer2_outputs(3719) <= not a or b;
    layer2_outputs(3720) <= a;
    layer2_outputs(3721) <= a xor b;
    layer2_outputs(3722) <= not (a and b);
    layer2_outputs(3723) <= a xor b;
    layer2_outputs(3724) <= a and not b;
    layer2_outputs(3725) <= not (a or b);
    layer2_outputs(3726) <= not (a and b);
    layer2_outputs(3727) <= not (a and b);
    layer2_outputs(3728) <= not a;
    layer2_outputs(3729) <= a;
    layer2_outputs(3730) <= not b or a;
    layer2_outputs(3731) <= not (a or b);
    layer2_outputs(3732) <= not b or a;
    layer2_outputs(3733) <= a or b;
    layer2_outputs(3734) <= a xor b;
    layer2_outputs(3735) <= b and not a;
    layer2_outputs(3736) <= not (a xor b);
    layer2_outputs(3737) <= not b;
    layer2_outputs(3738) <= b and not a;
    layer2_outputs(3739) <= a and b;
    layer2_outputs(3740) <= b;
    layer2_outputs(3741) <= not a;
    layer2_outputs(3742) <= a;
    layer2_outputs(3743) <= not (a and b);
    layer2_outputs(3744) <= not (a xor b);
    layer2_outputs(3745) <= not a;
    layer2_outputs(3746) <= not a;
    layer2_outputs(3747) <= b;
    layer2_outputs(3748) <= not b or a;
    layer2_outputs(3749) <= not (a xor b);
    layer2_outputs(3750) <= not (a xor b);
    layer2_outputs(3751) <= b and not a;
    layer2_outputs(3752) <= not b or a;
    layer2_outputs(3753) <= a;
    layer2_outputs(3754) <= not a;
    layer2_outputs(3755) <= b and not a;
    layer2_outputs(3756) <= a and b;
    layer2_outputs(3757) <= not (a or b);
    layer2_outputs(3758) <= not b or a;
    layer2_outputs(3759) <= not (a xor b);
    layer2_outputs(3760) <= b and not a;
    layer2_outputs(3761) <= not (a xor b);
    layer2_outputs(3762) <= b;
    layer2_outputs(3763) <= not (a or b);
    layer2_outputs(3764) <= not b or a;
    layer2_outputs(3765) <= a xor b;
    layer2_outputs(3766) <= not a;
    layer2_outputs(3767) <= not (a and b);
    layer2_outputs(3768) <= not (a or b);
    layer2_outputs(3769) <= b;
    layer2_outputs(3770) <= not b;
    layer2_outputs(3771) <= not a;
    layer2_outputs(3772) <= not a or b;
    layer2_outputs(3773) <= not (a or b);
    layer2_outputs(3774) <= not (a or b);
    layer2_outputs(3775) <= a xor b;
    layer2_outputs(3776) <= not a;
    layer2_outputs(3777) <= not a;
    layer2_outputs(3778) <= b and not a;
    layer2_outputs(3779) <= not b;
    layer2_outputs(3780) <= b;
    layer2_outputs(3781) <= not a;
    layer2_outputs(3782) <= not (a or b);
    layer2_outputs(3783) <= not (a xor b);
    layer2_outputs(3784) <= not a;
    layer2_outputs(3785) <= not b or a;
    layer2_outputs(3786) <= b;
    layer2_outputs(3787) <= not a;
    layer2_outputs(3788) <= 1'b0;
    layer2_outputs(3789) <= not (a or b);
    layer2_outputs(3790) <= not b or a;
    layer2_outputs(3791) <= a and not b;
    layer2_outputs(3792) <= not (a or b);
    layer2_outputs(3793) <= not a or b;
    layer2_outputs(3794) <= a and b;
    layer2_outputs(3795) <= not (a or b);
    layer2_outputs(3796) <= b and not a;
    layer2_outputs(3797) <= a and b;
    layer2_outputs(3798) <= not b;
    layer2_outputs(3799) <= a xor b;
    layer2_outputs(3800) <= a;
    layer2_outputs(3801) <= a;
    layer2_outputs(3802) <= a;
    layer2_outputs(3803) <= a xor b;
    layer2_outputs(3804) <= not a;
    layer2_outputs(3805) <= 1'b0;
    layer2_outputs(3806) <= a;
    layer2_outputs(3807) <= a;
    layer2_outputs(3808) <= not (a or b);
    layer2_outputs(3809) <= not b;
    layer2_outputs(3810) <= a xor b;
    layer2_outputs(3811) <= not a or b;
    layer2_outputs(3812) <= a;
    layer2_outputs(3813) <= not (a and b);
    layer2_outputs(3814) <= not (a or b);
    layer2_outputs(3815) <= b and not a;
    layer2_outputs(3816) <= a or b;
    layer2_outputs(3817) <= not a;
    layer2_outputs(3818) <= b;
    layer2_outputs(3819) <= not b or a;
    layer2_outputs(3820) <= not b;
    layer2_outputs(3821) <= not b;
    layer2_outputs(3822) <= not a;
    layer2_outputs(3823) <= a or b;
    layer2_outputs(3824) <= not b or a;
    layer2_outputs(3825) <= a and b;
    layer2_outputs(3826) <= not a or b;
    layer2_outputs(3827) <= a xor b;
    layer2_outputs(3828) <= a and not b;
    layer2_outputs(3829) <= a and not b;
    layer2_outputs(3830) <= not a;
    layer2_outputs(3831) <= not (a xor b);
    layer2_outputs(3832) <= a;
    layer2_outputs(3833) <= a;
    layer2_outputs(3834) <= a;
    layer2_outputs(3835) <= not b;
    layer2_outputs(3836) <= not a;
    layer2_outputs(3837) <= a and b;
    layer2_outputs(3838) <= a and b;
    layer2_outputs(3839) <= a;
    layer2_outputs(3840) <= not (a or b);
    layer2_outputs(3841) <= not a;
    layer2_outputs(3842) <= a xor b;
    layer2_outputs(3843) <= a and not b;
    layer2_outputs(3844) <= not a;
    layer2_outputs(3845) <= a and not b;
    layer2_outputs(3846) <= not (a and b);
    layer2_outputs(3847) <= a xor b;
    layer2_outputs(3848) <= a;
    layer2_outputs(3849) <= a and not b;
    layer2_outputs(3850) <= a or b;
    layer2_outputs(3851) <= not b or a;
    layer2_outputs(3852) <= b;
    layer2_outputs(3853) <= b;
    layer2_outputs(3854) <= not (a and b);
    layer2_outputs(3855) <= a and not b;
    layer2_outputs(3856) <= not a or b;
    layer2_outputs(3857) <= a and b;
    layer2_outputs(3858) <= a and not b;
    layer2_outputs(3859) <= not a;
    layer2_outputs(3860) <= not (a and b);
    layer2_outputs(3861) <= a or b;
    layer2_outputs(3862) <= not (a or b);
    layer2_outputs(3863) <= b;
    layer2_outputs(3864) <= not b;
    layer2_outputs(3865) <= a;
    layer2_outputs(3866) <= not a;
    layer2_outputs(3867) <= a xor b;
    layer2_outputs(3868) <= b;
    layer2_outputs(3869) <= not a or b;
    layer2_outputs(3870) <= not b or a;
    layer2_outputs(3871) <= not (a and b);
    layer2_outputs(3872) <= not a or b;
    layer2_outputs(3873) <= b;
    layer2_outputs(3874) <= a and b;
    layer2_outputs(3875) <= not b;
    layer2_outputs(3876) <= not a;
    layer2_outputs(3877) <= not (a or b);
    layer2_outputs(3878) <= a or b;
    layer2_outputs(3879) <= not (a and b);
    layer2_outputs(3880) <= not b or a;
    layer2_outputs(3881) <= not b or a;
    layer2_outputs(3882) <= b and not a;
    layer2_outputs(3883) <= not (a or b);
    layer2_outputs(3884) <= not a;
    layer2_outputs(3885) <= a or b;
    layer2_outputs(3886) <= not b;
    layer2_outputs(3887) <= a xor b;
    layer2_outputs(3888) <= not b or a;
    layer2_outputs(3889) <= b;
    layer2_outputs(3890) <= not b or a;
    layer2_outputs(3891) <= b;
    layer2_outputs(3892) <= b;
    layer2_outputs(3893) <= not a;
    layer2_outputs(3894) <= not b;
    layer2_outputs(3895) <= b and not a;
    layer2_outputs(3896) <= b;
    layer2_outputs(3897) <= not b;
    layer2_outputs(3898) <= not (a xor b);
    layer2_outputs(3899) <= not a;
    layer2_outputs(3900) <= not b or a;
    layer2_outputs(3901) <= not (a or b);
    layer2_outputs(3902) <= not (a and b);
    layer2_outputs(3903) <= not b;
    layer2_outputs(3904) <= not b;
    layer2_outputs(3905) <= a or b;
    layer2_outputs(3906) <= a;
    layer2_outputs(3907) <= a and b;
    layer2_outputs(3908) <= not (a or b);
    layer2_outputs(3909) <= a;
    layer2_outputs(3910) <= not b;
    layer2_outputs(3911) <= not b or a;
    layer2_outputs(3912) <= b and not a;
    layer2_outputs(3913) <= not a or b;
    layer2_outputs(3914) <= not a or b;
    layer2_outputs(3915) <= b;
    layer2_outputs(3916) <= not (a and b);
    layer2_outputs(3917) <= b;
    layer2_outputs(3918) <= a;
    layer2_outputs(3919) <= a and not b;
    layer2_outputs(3920) <= b;
    layer2_outputs(3921) <= a;
    layer2_outputs(3922) <= a or b;
    layer2_outputs(3923) <= not a or b;
    layer2_outputs(3924) <= a;
    layer2_outputs(3925) <= a;
    layer2_outputs(3926) <= a;
    layer2_outputs(3927) <= not a;
    layer2_outputs(3928) <= not (a xor b);
    layer2_outputs(3929) <= not (a or b);
    layer2_outputs(3930) <= a;
    layer2_outputs(3931) <= b;
    layer2_outputs(3932) <= b;
    layer2_outputs(3933) <= a xor b;
    layer2_outputs(3934) <= b;
    layer2_outputs(3935) <= b and not a;
    layer2_outputs(3936) <= b;
    layer2_outputs(3937) <= not a;
    layer2_outputs(3938) <= b and not a;
    layer2_outputs(3939) <= b;
    layer2_outputs(3940) <= not a;
    layer2_outputs(3941) <= not (a and b);
    layer2_outputs(3942) <= b;
    layer2_outputs(3943) <= b;
    layer2_outputs(3944) <= a and b;
    layer2_outputs(3945) <= not a;
    layer2_outputs(3946) <= not (a or b);
    layer2_outputs(3947) <= a;
    layer2_outputs(3948) <= b;
    layer2_outputs(3949) <= not b;
    layer2_outputs(3950) <= a;
    layer2_outputs(3951) <= not b;
    layer2_outputs(3952) <= not (a xor b);
    layer2_outputs(3953) <= not b;
    layer2_outputs(3954) <= b;
    layer2_outputs(3955) <= not a or b;
    layer2_outputs(3956) <= not a;
    layer2_outputs(3957) <= a and not b;
    layer2_outputs(3958) <= a and b;
    layer2_outputs(3959) <= 1'b0;
    layer2_outputs(3960) <= a and not b;
    layer2_outputs(3961) <= not a or b;
    layer2_outputs(3962) <= a or b;
    layer2_outputs(3963) <= a or b;
    layer2_outputs(3964) <= not a;
    layer2_outputs(3965) <= a or b;
    layer2_outputs(3966) <= not b;
    layer2_outputs(3967) <= not (a and b);
    layer2_outputs(3968) <= b;
    layer2_outputs(3969) <= not a;
    layer2_outputs(3970) <= not (a xor b);
    layer2_outputs(3971) <= not b or a;
    layer2_outputs(3972) <= not (a or b);
    layer2_outputs(3973) <= a;
    layer2_outputs(3974) <= not (a and b);
    layer2_outputs(3975) <= not (a xor b);
    layer2_outputs(3976) <= not b or a;
    layer2_outputs(3977) <= a or b;
    layer2_outputs(3978) <= not (a xor b);
    layer2_outputs(3979) <= not a or b;
    layer2_outputs(3980) <= not a;
    layer2_outputs(3981) <= a and b;
    layer2_outputs(3982) <= not b or a;
    layer2_outputs(3983) <= 1'b1;
    layer2_outputs(3984) <= not a;
    layer2_outputs(3985) <= a xor b;
    layer2_outputs(3986) <= not b or a;
    layer2_outputs(3987) <= not (a xor b);
    layer2_outputs(3988) <= a xor b;
    layer2_outputs(3989) <= b and not a;
    layer2_outputs(3990) <= not a;
    layer2_outputs(3991) <= a;
    layer2_outputs(3992) <= not (a xor b);
    layer2_outputs(3993) <= b and not a;
    layer2_outputs(3994) <= a and not b;
    layer2_outputs(3995) <= not b;
    layer2_outputs(3996) <= b;
    layer2_outputs(3997) <= a or b;
    layer2_outputs(3998) <= b;
    layer2_outputs(3999) <= not a or b;
    layer2_outputs(4000) <= b;
    layer2_outputs(4001) <= a or b;
    layer2_outputs(4002) <= not a or b;
    layer2_outputs(4003) <= not a or b;
    layer2_outputs(4004) <= b and not a;
    layer2_outputs(4005) <= a or b;
    layer2_outputs(4006) <= not a or b;
    layer2_outputs(4007) <= a and not b;
    layer2_outputs(4008) <= b;
    layer2_outputs(4009) <= a xor b;
    layer2_outputs(4010) <= not (a and b);
    layer2_outputs(4011) <= not a;
    layer2_outputs(4012) <= not b or a;
    layer2_outputs(4013) <= not (a and b);
    layer2_outputs(4014) <= a or b;
    layer2_outputs(4015) <= b;
    layer2_outputs(4016) <= not (a xor b);
    layer2_outputs(4017) <= a;
    layer2_outputs(4018) <= a;
    layer2_outputs(4019) <= a and not b;
    layer2_outputs(4020) <= b;
    layer2_outputs(4021) <= a and not b;
    layer2_outputs(4022) <= not b;
    layer2_outputs(4023) <= not b or a;
    layer2_outputs(4024) <= not (a xor b);
    layer2_outputs(4025) <= not b;
    layer2_outputs(4026) <= a or b;
    layer2_outputs(4027) <= not b or a;
    layer2_outputs(4028) <= b;
    layer2_outputs(4029) <= not b;
    layer2_outputs(4030) <= a and not b;
    layer2_outputs(4031) <= not (a or b);
    layer2_outputs(4032) <= b;
    layer2_outputs(4033) <= not b;
    layer2_outputs(4034) <= not a;
    layer2_outputs(4035) <= a;
    layer2_outputs(4036) <= a and not b;
    layer2_outputs(4037) <= not a or b;
    layer2_outputs(4038) <= 1'b0;
    layer2_outputs(4039) <= b and not a;
    layer2_outputs(4040) <= a;
    layer2_outputs(4041) <= a and not b;
    layer2_outputs(4042) <= not a or b;
    layer2_outputs(4043) <= not b or a;
    layer2_outputs(4044) <= not a;
    layer2_outputs(4045) <= not b;
    layer2_outputs(4046) <= b and not a;
    layer2_outputs(4047) <= not (a and b);
    layer2_outputs(4048) <= a xor b;
    layer2_outputs(4049) <= not (a and b);
    layer2_outputs(4050) <= not (a xor b);
    layer2_outputs(4051) <= not (a or b);
    layer2_outputs(4052) <= a and not b;
    layer2_outputs(4053) <= not b or a;
    layer2_outputs(4054) <= a;
    layer2_outputs(4055) <= not b or a;
    layer2_outputs(4056) <= b;
    layer2_outputs(4057) <= a;
    layer2_outputs(4058) <= not (a and b);
    layer2_outputs(4059) <= not a;
    layer2_outputs(4060) <= not (a or b);
    layer2_outputs(4061) <= b;
    layer2_outputs(4062) <= b;
    layer2_outputs(4063) <= not a;
    layer2_outputs(4064) <= a and b;
    layer2_outputs(4065) <= not a or b;
    layer2_outputs(4066) <= not b;
    layer2_outputs(4067) <= b;
    layer2_outputs(4068) <= a and b;
    layer2_outputs(4069) <= a and not b;
    layer2_outputs(4070) <= a and b;
    layer2_outputs(4071) <= b and not a;
    layer2_outputs(4072) <= not a;
    layer2_outputs(4073) <= not b;
    layer2_outputs(4074) <= not a or b;
    layer2_outputs(4075) <= not b;
    layer2_outputs(4076) <= not a;
    layer2_outputs(4077) <= a or b;
    layer2_outputs(4078) <= b;
    layer2_outputs(4079) <= not b or a;
    layer2_outputs(4080) <= a;
    layer2_outputs(4081) <= a xor b;
    layer2_outputs(4082) <= a;
    layer2_outputs(4083) <= a and not b;
    layer2_outputs(4084) <= b and not a;
    layer2_outputs(4085) <= not a;
    layer2_outputs(4086) <= a or b;
    layer2_outputs(4087) <= 1'b0;
    layer2_outputs(4088) <= a;
    layer2_outputs(4089) <= a or b;
    layer2_outputs(4090) <= not (a and b);
    layer2_outputs(4091) <= b and not a;
    layer2_outputs(4092) <= b;
    layer2_outputs(4093) <= a and not b;
    layer2_outputs(4094) <= b;
    layer2_outputs(4095) <= b and not a;
    layer2_outputs(4096) <= not (a and b);
    layer2_outputs(4097) <= not a;
    layer2_outputs(4098) <= not (a and b);
    layer2_outputs(4099) <= not (a and b);
    layer2_outputs(4100) <= a;
    layer2_outputs(4101) <= a and not b;
    layer2_outputs(4102) <= not a;
    layer2_outputs(4103) <= not a or b;
    layer2_outputs(4104) <= not (a and b);
    layer2_outputs(4105) <= a and not b;
    layer2_outputs(4106) <= a;
    layer2_outputs(4107) <= not (a and b);
    layer2_outputs(4108) <= b and not a;
    layer2_outputs(4109) <= not (a and b);
    layer2_outputs(4110) <= not (a and b);
    layer2_outputs(4111) <= 1'b1;
    layer2_outputs(4112) <= b and not a;
    layer2_outputs(4113) <= not a or b;
    layer2_outputs(4114) <= not (a and b);
    layer2_outputs(4115) <= not (a or b);
    layer2_outputs(4116) <= not (a or b);
    layer2_outputs(4117) <= not (a xor b);
    layer2_outputs(4118) <= a and b;
    layer2_outputs(4119) <= not b;
    layer2_outputs(4120) <= not a;
    layer2_outputs(4121) <= a;
    layer2_outputs(4122) <= b and not a;
    layer2_outputs(4123) <= a and not b;
    layer2_outputs(4124) <= not (a and b);
    layer2_outputs(4125) <= not a;
    layer2_outputs(4126) <= b;
    layer2_outputs(4127) <= a and b;
    layer2_outputs(4128) <= not (a xor b);
    layer2_outputs(4129) <= a;
    layer2_outputs(4130) <= b;
    layer2_outputs(4131) <= b;
    layer2_outputs(4132) <= b;
    layer2_outputs(4133) <= a or b;
    layer2_outputs(4134) <= a;
    layer2_outputs(4135) <= not (a xor b);
    layer2_outputs(4136) <= a and b;
    layer2_outputs(4137) <= b;
    layer2_outputs(4138) <= b and not a;
    layer2_outputs(4139) <= b;
    layer2_outputs(4140) <= a and b;
    layer2_outputs(4141) <= not a;
    layer2_outputs(4142) <= not b;
    layer2_outputs(4143) <= a;
    layer2_outputs(4144) <= a and b;
    layer2_outputs(4145) <= not b;
    layer2_outputs(4146) <= a and not b;
    layer2_outputs(4147) <= a;
    layer2_outputs(4148) <= not (a and b);
    layer2_outputs(4149) <= not (a or b);
    layer2_outputs(4150) <= a or b;
    layer2_outputs(4151) <= not (a and b);
    layer2_outputs(4152) <= a and not b;
    layer2_outputs(4153) <= not (a and b);
    layer2_outputs(4154) <= not (a and b);
    layer2_outputs(4155) <= b and not a;
    layer2_outputs(4156) <= a;
    layer2_outputs(4157) <= not a;
    layer2_outputs(4158) <= not (a or b);
    layer2_outputs(4159) <= b;
    layer2_outputs(4160) <= b and not a;
    layer2_outputs(4161) <= b and not a;
    layer2_outputs(4162) <= not b;
    layer2_outputs(4163) <= a xor b;
    layer2_outputs(4164) <= a and not b;
    layer2_outputs(4165) <= a or b;
    layer2_outputs(4166) <= a;
    layer2_outputs(4167) <= not (a xor b);
    layer2_outputs(4168) <= b and not a;
    layer2_outputs(4169) <= b;
    layer2_outputs(4170) <= not (a or b);
    layer2_outputs(4171) <= b and not a;
    layer2_outputs(4172) <= a;
    layer2_outputs(4173) <= not a or b;
    layer2_outputs(4174) <= not (a or b);
    layer2_outputs(4175) <= a or b;
    layer2_outputs(4176) <= not a;
    layer2_outputs(4177) <= b and not a;
    layer2_outputs(4178) <= a and not b;
    layer2_outputs(4179) <= a or b;
    layer2_outputs(4180) <= not (a and b);
    layer2_outputs(4181) <= a and b;
    layer2_outputs(4182) <= not b;
    layer2_outputs(4183) <= b;
    layer2_outputs(4184) <= a xor b;
    layer2_outputs(4185) <= not b;
    layer2_outputs(4186) <= a;
    layer2_outputs(4187) <= not (a and b);
    layer2_outputs(4188) <= not (a and b);
    layer2_outputs(4189) <= not (a and b);
    layer2_outputs(4190) <= not (a and b);
    layer2_outputs(4191) <= not b;
    layer2_outputs(4192) <= not (a or b);
    layer2_outputs(4193) <= not a;
    layer2_outputs(4194) <= b;
    layer2_outputs(4195) <= b;
    layer2_outputs(4196) <= not a;
    layer2_outputs(4197) <= a xor b;
    layer2_outputs(4198) <= not b;
    layer2_outputs(4199) <= a and b;
    layer2_outputs(4200) <= not (a and b);
    layer2_outputs(4201) <= not b or a;
    layer2_outputs(4202) <= 1'b0;
    layer2_outputs(4203) <= a and b;
    layer2_outputs(4204) <= not b or a;
    layer2_outputs(4205) <= not (a xor b);
    layer2_outputs(4206) <= a or b;
    layer2_outputs(4207) <= not (a or b);
    layer2_outputs(4208) <= not (a and b);
    layer2_outputs(4209) <= not (a xor b);
    layer2_outputs(4210) <= b and not a;
    layer2_outputs(4211) <= not (a or b);
    layer2_outputs(4212) <= not b;
    layer2_outputs(4213) <= a and b;
    layer2_outputs(4214) <= not (a or b);
    layer2_outputs(4215) <= b;
    layer2_outputs(4216) <= not b;
    layer2_outputs(4217) <= a and b;
    layer2_outputs(4218) <= not a;
    layer2_outputs(4219) <= b;
    layer2_outputs(4220) <= b;
    layer2_outputs(4221) <= not b;
    layer2_outputs(4222) <= b and not a;
    layer2_outputs(4223) <= b;
    layer2_outputs(4224) <= not b or a;
    layer2_outputs(4225) <= a and not b;
    layer2_outputs(4226) <= a;
    layer2_outputs(4227) <= not a or b;
    layer2_outputs(4228) <= not (a xor b);
    layer2_outputs(4229) <= b and not a;
    layer2_outputs(4230) <= not a;
    layer2_outputs(4231) <= not a or b;
    layer2_outputs(4232) <= b;
    layer2_outputs(4233) <= a xor b;
    layer2_outputs(4234) <= b;
    layer2_outputs(4235) <= a;
    layer2_outputs(4236) <= not a or b;
    layer2_outputs(4237) <= not a;
    layer2_outputs(4238) <= not a or b;
    layer2_outputs(4239) <= not (a or b);
    layer2_outputs(4240) <= not a;
    layer2_outputs(4241) <= a and not b;
    layer2_outputs(4242) <= b and not a;
    layer2_outputs(4243) <= a;
    layer2_outputs(4244) <= b;
    layer2_outputs(4245) <= not (a xor b);
    layer2_outputs(4246) <= not (a or b);
    layer2_outputs(4247) <= not (a and b);
    layer2_outputs(4248) <= not (a or b);
    layer2_outputs(4249) <= a and b;
    layer2_outputs(4250) <= not a;
    layer2_outputs(4251) <= not (a xor b);
    layer2_outputs(4252) <= a;
    layer2_outputs(4253) <= a and not b;
    layer2_outputs(4254) <= b;
    layer2_outputs(4255) <= not a;
    layer2_outputs(4256) <= not (a and b);
    layer2_outputs(4257) <= 1'b1;
    layer2_outputs(4258) <= a;
    layer2_outputs(4259) <= a xor b;
    layer2_outputs(4260) <= b;
    layer2_outputs(4261) <= b and not a;
    layer2_outputs(4262) <= not a or b;
    layer2_outputs(4263) <= not (a xor b);
    layer2_outputs(4264) <= a and b;
    layer2_outputs(4265) <= a;
    layer2_outputs(4266) <= a xor b;
    layer2_outputs(4267) <= not (a and b);
    layer2_outputs(4268) <= not a;
    layer2_outputs(4269) <= not b;
    layer2_outputs(4270) <= a;
    layer2_outputs(4271) <= not a;
    layer2_outputs(4272) <= b and not a;
    layer2_outputs(4273) <= a and b;
    layer2_outputs(4274) <= a xor b;
    layer2_outputs(4275) <= b;
    layer2_outputs(4276) <= a or b;
    layer2_outputs(4277) <= a and not b;
    layer2_outputs(4278) <= not b or a;
    layer2_outputs(4279) <= a and b;
    layer2_outputs(4280) <= not b;
    layer2_outputs(4281) <= a or b;
    layer2_outputs(4282) <= a;
    layer2_outputs(4283) <= b;
    layer2_outputs(4284) <= not a or b;
    layer2_outputs(4285) <= not (a and b);
    layer2_outputs(4286) <= not (a xor b);
    layer2_outputs(4287) <= a;
    layer2_outputs(4288) <= not (a and b);
    layer2_outputs(4289) <= not a or b;
    layer2_outputs(4290) <= not b;
    layer2_outputs(4291) <= b and not a;
    layer2_outputs(4292) <= 1'b1;
    layer2_outputs(4293) <= not a or b;
    layer2_outputs(4294) <= b and not a;
    layer2_outputs(4295) <= not b;
    layer2_outputs(4296) <= not (a or b);
    layer2_outputs(4297) <= a and b;
    layer2_outputs(4298) <= a and b;
    layer2_outputs(4299) <= a and not b;
    layer2_outputs(4300) <= not b or a;
    layer2_outputs(4301) <= not (a xor b);
    layer2_outputs(4302) <= not (a and b);
    layer2_outputs(4303) <= a and b;
    layer2_outputs(4304) <= not b or a;
    layer2_outputs(4305) <= not a;
    layer2_outputs(4306) <= not b;
    layer2_outputs(4307) <= not a;
    layer2_outputs(4308) <= a;
    layer2_outputs(4309) <= not (a xor b);
    layer2_outputs(4310) <= not (a and b);
    layer2_outputs(4311) <= a;
    layer2_outputs(4312) <= a;
    layer2_outputs(4313) <= 1'b0;
    layer2_outputs(4314) <= a and b;
    layer2_outputs(4315) <= a or b;
    layer2_outputs(4316) <= b;
    layer2_outputs(4317) <= not b;
    layer2_outputs(4318) <= a and not b;
    layer2_outputs(4319) <= a or b;
    layer2_outputs(4320) <= not (a or b);
    layer2_outputs(4321) <= not a or b;
    layer2_outputs(4322) <= a and b;
    layer2_outputs(4323) <= a;
    layer2_outputs(4324) <= not b or a;
    layer2_outputs(4325) <= not (a or b);
    layer2_outputs(4326) <= b and not a;
    layer2_outputs(4327) <= not b or a;
    layer2_outputs(4328) <= not (a or b);
    layer2_outputs(4329) <= not a;
    layer2_outputs(4330) <= not (a xor b);
    layer2_outputs(4331) <= b;
    layer2_outputs(4332) <= a and b;
    layer2_outputs(4333) <= not b;
    layer2_outputs(4334) <= not (a xor b);
    layer2_outputs(4335) <= not (a and b);
    layer2_outputs(4336) <= a or b;
    layer2_outputs(4337) <= a and not b;
    layer2_outputs(4338) <= not a or b;
    layer2_outputs(4339) <= not (a or b);
    layer2_outputs(4340) <= not b;
    layer2_outputs(4341) <= b;
    layer2_outputs(4342) <= a;
    layer2_outputs(4343) <= a xor b;
    layer2_outputs(4344) <= a and not b;
    layer2_outputs(4345) <= a or b;
    layer2_outputs(4346) <= not a;
    layer2_outputs(4347) <= not (a xor b);
    layer2_outputs(4348) <= not b or a;
    layer2_outputs(4349) <= 1'b1;
    layer2_outputs(4350) <= b and not a;
    layer2_outputs(4351) <= not b or a;
    layer2_outputs(4352) <= a;
    layer2_outputs(4353) <= not b or a;
    layer2_outputs(4354) <= a;
    layer2_outputs(4355) <= not b or a;
    layer2_outputs(4356) <= not b;
    layer2_outputs(4357) <= not b;
    layer2_outputs(4358) <= a;
    layer2_outputs(4359) <= not (a or b);
    layer2_outputs(4360) <= a and not b;
    layer2_outputs(4361) <= not (a or b);
    layer2_outputs(4362) <= not a or b;
    layer2_outputs(4363) <= a;
    layer2_outputs(4364) <= not a or b;
    layer2_outputs(4365) <= b and not a;
    layer2_outputs(4366) <= not a;
    layer2_outputs(4367) <= not (a xor b);
    layer2_outputs(4368) <= not (a and b);
    layer2_outputs(4369) <= a xor b;
    layer2_outputs(4370) <= not (a or b);
    layer2_outputs(4371) <= b and not a;
    layer2_outputs(4372) <= not b;
    layer2_outputs(4373) <= not (a xor b);
    layer2_outputs(4374) <= not b or a;
    layer2_outputs(4375) <= b;
    layer2_outputs(4376) <= a;
    layer2_outputs(4377) <= not b;
    layer2_outputs(4378) <= not (a or b);
    layer2_outputs(4379) <= b;
    layer2_outputs(4380) <= a and not b;
    layer2_outputs(4381) <= a;
    layer2_outputs(4382) <= a;
    layer2_outputs(4383) <= b;
    layer2_outputs(4384) <= a and b;
    layer2_outputs(4385) <= 1'b0;
    layer2_outputs(4386) <= b;
    layer2_outputs(4387) <= a and not b;
    layer2_outputs(4388) <= a and not b;
    layer2_outputs(4389) <= not (a xor b);
    layer2_outputs(4390) <= not b;
    layer2_outputs(4391) <= not a;
    layer2_outputs(4392) <= not b;
    layer2_outputs(4393) <= a;
    layer2_outputs(4394) <= not b or a;
    layer2_outputs(4395) <= not (a xor b);
    layer2_outputs(4396) <= not a or b;
    layer2_outputs(4397) <= not (a xor b);
    layer2_outputs(4398) <= not a;
    layer2_outputs(4399) <= not (a or b);
    layer2_outputs(4400) <= not a or b;
    layer2_outputs(4401) <= not (a or b);
    layer2_outputs(4402) <= b and not a;
    layer2_outputs(4403) <= not a;
    layer2_outputs(4404) <= not a or b;
    layer2_outputs(4405) <= not (a and b);
    layer2_outputs(4406) <= a and not b;
    layer2_outputs(4407) <= not a;
    layer2_outputs(4408) <= not a;
    layer2_outputs(4409) <= b;
    layer2_outputs(4410) <= b and not a;
    layer2_outputs(4411) <= not b or a;
    layer2_outputs(4412) <= not a;
    layer2_outputs(4413) <= not a;
    layer2_outputs(4414) <= not (a or b);
    layer2_outputs(4415) <= not b;
    layer2_outputs(4416) <= a and b;
    layer2_outputs(4417) <= 1'b0;
    layer2_outputs(4418) <= b;
    layer2_outputs(4419) <= b and not a;
    layer2_outputs(4420) <= not a;
    layer2_outputs(4421) <= b;
    layer2_outputs(4422) <= 1'b1;
    layer2_outputs(4423) <= not (a xor b);
    layer2_outputs(4424) <= a or b;
    layer2_outputs(4425) <= a xor b;
    layer2_outputs(4426) <= not (a or b);
    layer2_outputs(4427) <= not (a and b);
    layer2_outputs(4428) <= not b;
    layer2_outputs(4429) <= a and not b;
    layer2_outputs(4430) <= not (a and b);
    layer2_outputs(4431) <= a or b;
    layer2_outputs(4432) <= not (a and b);
    layer2_outputs(4433) <= b and not a;
    layer2_outputs(4434) <= not b or a;
    layer2_outputs(4435) <= b;
    layer2_outputs(4436) <= not b;
    layer2_outputs(4437) <= a and b;
    layer2_outputs(4438) <= not a or b;
    layer2_outputs(4439) <= not a;
    layer2_outputs(4440) <= not (a xor b);
    layer2_outputs(4441) <= b;
    layer2_outputs(4442) <= a and not b;
    layer2_outputs(4443) <= not b;
    layer2_outputs(4444) <= a xor b;
    layer2_outputs(4445) <= not (a or b);
    layer2_outputs(4446) <= not (a and b);
    layer2_outputs(4447) <= not (a and b);
    layer2_outputs(4448) <= not (a or b);
    layer2_outputs(4449) <= not (a xor b);
    layer2_outputs(4450) <= a or b;
    layer2_outputs(4451) <= not b;
    layer2_outputs(4452) <= a and b;
    layer2_outputs(4453) <= not a;
    layer2_outputs(4454) <= not b;
    layer2_outputs(4455) <= not (a and b);
    layer2_outputs(4456) <= not a;
    layer2_outputs(4457) <= not (a xor b);
    layer2_outputs(4458) <= not (a or b);
    layer2_outputs(4459) <= not b;
    layer2_outputs(4460) <= not b;
    layer2_outputs(4461) <= not b or a;
    layer2_outputs(4462) <= b;
    layer2_outputs(4463) <= a and b;
    layer2_outputs(4464) <= not (a xor b);
    layer2_outputs(4465) <= not (a xor b);
    layer2_outputs(4466) <= 1'b0;
    layer2_outputs(4467) <= b;
    layer2_outputs(4468) <= a and b;
    layer2_outputs(4469) <= not (a and b);
    layer2_outputs(4470) <= b;
    layer2_outputs(4471) <= not (a and b);
    layer2_outputs(4472) <= a;
    layer2_outputs(4473) <= b and not a;
    layer2_outputs(4474) <= not b;
    layer2_outputs(4475) <= b;
    layer2_outputs(4476) <= not (a xor b);
    layer2_outputs(4477) <= not b or a;
    layer2_outputs(4478) <= not (a and b);
    layer2_outputs(4479) <= not a;
    layer2_outputs(4480) <= b and not a;
    layer2_outputs(4481) <= b and not a;
    layer2_outputs(4482) <= b and not a;
    layer2_outputs(4483) <= not (a or b);
    layer2_outputs(4484) <= b and not a;
    layer2_outputs(4485) <= a and b;
    layer2_outputs(4486) <= not (a and b);
    layer2_outputs(4487) <= not a or b;
    layer2_outputs(4488) <= not (a xor b);
    layer2_outputs(4489) <= 1'b1;
    layer2_outputs(4490) <= b and not a;
    layer2_outputs(4491) <= not (a xor b);
    layer2_outputs(4492) <= not b or a;
    layer2_outputs(4493) <= not (a or b);
    layer2_outputs(4494) <= a and not b;
    layer2_outputs(4495) <= a or b;
    layer2_outputs(4496) <= a and b;
    layer2_outputs(4497) <= b and not a;
    layer2_outputs(4498) <= a xor b;
    layer2_outputs(4499) <= not b or a;
    layer2_outputs(4500) <= a and b;
    layer2_outputs(4501) <= not b;
    layer2_outputs(4502) <= not a;
    layer2_outputs(4503) <= not b or a;
    layer2_outputs(4504) <= a xor b;
    layer2_outputs(4505) <= not a or b;
    layer2_outputs(4506) <= a and b;
    layer2_outputs(4507) <= a xor b;
    layer2_outputs(4508) <= a;
    layer2_outputs(4509) <= not (a and b);
    layer2_outputs(4510) <= a;
    layer2_outputs(4511) <= a and b;
    layer2_outputs(4512) <= a and not b;
    layer2_outputs(4513) <= not b;
    layer2_outputs(4514) <= not a;
    layer2_outputs(4515) <= a;
    layer2_outputs(4516) <= not b;
    layer2_outputs(4517) <= not a;
    layer2_outputs(4518) <= not b;
    layer2_outputs(4519) <= b;
    layer2_outputs(4520) <= not a or b;
    layer2_outputs(4521) <= not b or a;
    layer2_outputs(4522) <= a and b;
    layer2_outputs(4523) <= not b;
    layer2_outputs(4524) <= not a;
    layer2_outputs(4525) <= not b;
    layer2_outputs(4526) <= a;
    layer2_outputs(4527) <= not a or b;
    layer2_outputs(4528) <= not b;
    layer2_outputs(4529) <= a xor b;
    layer2_outputs(4530) <= not b;
    layer2_outputs(4531) <= not a or b;
    layer2_outputs(4532) <= a and b;
    layer2_outputs(4533) <= not a;
    layer2_outputs(4534) <= not (a xor b);
    layer2_outputs(4535) <= not a;
    layer2_outputs(4536) <= a and not b;
    layer2_outputs(4537) <= a and b;
    layer2_outputs(4538) <= not b;
    layer2_outputs(4539) <= not (a and b);
    layer2_outputs(4540) <= a xor b;
    layer2_outputs(4541) <= not (a or b);
    layer2_outputs(4542) <= b and not a;
    layer2_outputs(4543) <= a;
    layer2_outputs(4544) <= not (a xor b);
    layer2_outputs(4545) <= not b or a;
    layer2_outputs(4546) <= not b;
    layer2_outputs(4547) <= not (a xor b);
    layer2_outputs(4548) <= b and not a;
    layer2_outputs(4549) <= not (a xor b);
    layer2_outputs(4550) <= a;
    layer2_outputs(4551) <= not b or a;
    layer2_outputs(4552) <= a xor b;
    layer2_outputs(4553) <= b;
    layer2_outputs(4554) <= not b or a;
    layer2_outputs(4555) <= a xor b;
    layer2_outputs(4556) <= not (a and b);
    layer2_outputs(4557) <= not a;
    layer2_outputs(4558) <= not (a or b);
    layer2_outputs(4559) <= a and not b;
    layer2_outputs(4560) <= not (a and b);
    layer2_outputs(4561) <= not b or a;
    layer2_outputs(4562) <= b;
    layer2_outputs(4563) <= a and not b;
    layer2_outputs(4564) <= a and not b;
    layer2_outputs(4565) <= b and not a;
    layer2_outputs(4566) <= not b;
    layer2_outputs(4567) <= not b or a;
    layer2_outputs(4568) <= b;
    layer2_outputs(4569) <= not b;
    layer2_outputs(4570) <= a;
    layer2_outputs(4571) <= not a;
    layer2_outputs(4572) <= not (a xor b);
    layer2_outputs(4573) <= a;
    layer2_outputs(4574) <= a and not b;
    layer2_outputs(4575) <= not b;
    layer2_outputs(4576) <= not a;
    layer2_outputs(4577) <= not b;
    layer2_outputs(4578) <= a xor b;
    layer2_outputs(4579) <= not a or b;
    layer2_outputs(4580) <= a xor b;
    layer2_outputs(4581) <= a xor b;
    layer2_outputs(4582) <= a xor b;
    layer2_outputs(4583) <= not b;
    layer2_outputs(4584) <= a;
    layer2_outputs(4585) <= not a or b;
    layer2_outputs(4586) <= not (a or b);
    layer2_outputs(4587) <= not b;
    layer2_outputs(4588) <= b;
    layer2_outputs(4589) <= not b or a;
    layer2_outputs(4590) <= a xor b;
    layer2_outputs(4591) <= a and b;
    layer2_outputs(4592) <= a or b;
    layer2_outputs(4593) <= not b or a;
    layer2_outputs(4594) <= not (a xor b);
    layer2_outputs(4595) <= a xor b;
    layer2_outputs(4596) <= b;
    layer2_outputs(4597) <= a;
    layer2_outputs(4598) <= a xor b;
    layer2_outputs(4599) <= not a or b;
    layer2_outputs(4600) <= a and b;
    layer2_outputs(4601) <= a;
    layer2_outputs(4602) <= not a or b;
    layer2_outputs(4603) <= not b or a;
    layer2_outputs(4604) <= not (a or b);
    layer2_outputs(4605) <= a and b;
    layer2_outputs(4606) <= a and not b;
    layer2_outputs(4607) <= not (a xor b);
    layer2_outputs(4608) <= a;
    layer2_outputs(4609) <= b;
    layer2_outputs(4610) <= a and b;
    layer2_outputs(4611) <= not (a or b);
    layer2_outputs(4612) <= not b or a;
    layer2_outputs(4613) <= not (a or b);
    layer2_outputs(4614) <= not b;
    layer2_outputs(4615) <= a;
    layer2_outputs(4616) <= a and not b;
    layer2_outputs(4617) <= b and not a;
    layer2_outputs(4618) <= not (a and b);
    layer2_outputs(4619) <= a and b;
    layer2_outputs(4620) <= not (a xor b);
    layer2_outputs(4621) <= not (a and b);
    layer2_outputs(4622) <= not b;
    layer2_outputs(4623) <= not a;
    layer2_outputs(4624) <= not (a and b);
    layer2_outputs(4625) <= a;
    layer2_outputs(4626) <= a or b;
    layer2_outputs(4627) <= a and b;
    layer2_outputs(4628) <= a;
    layer2_outputs(4629) <= not b or a;
    layer2_outputs(4630) <= a and not b;
    layer2_outputs(4631) <= not (a and b);
    layer2_outputs(4632) <= not (a xor b);
    layer2_outputs(4633) <= not a;
    layer2_outputs(4634) <= a and not b;
    layer2_outputs(4635) <= not a or b;
    layer2_outputs(4636) <= not (a xor b);
    layer2_outputs(4637) <= not a;
    layer2_outputs(4638) <= a and b;
    layer2_outputs(4639) <= a xor b;
    layer2_outputs(4640) <= not b;
    layer2_outputs(4641) <= a or b;
    layer2_outputs(4642) <= a and b;
    layer2_outputs(4643) <= a xor b;
    layer2_outputs(4644) <= not (a xor b);
    layer2_outputs(4645) <= a and b;
    layer2_outputs(4646) <= not (a or b);
    layer2_outputs(4647) <= not (a or b);
    layer2_outputs(4648) <= a and b;
    layer2_outputs(4649) <= not b or a;
    layer2_outputs(4650) <= a and b;
    layer2_outputs(4651) <= b;
    layer2_outputs(4652) <= not a or b;
    layer2_outputs(4653) <= a xor b;
    layer2_outputs(4654) <= a xor b;
    layer2_outputs(4655) <= not a or b;
    layer2_outputs(4656) <= not a;
    layer2_outputs(4657) <= b;
    layer2_outputs(4658) <= a xor b;
    layer2_outputs(4659) <= a and not b;
    layer2_outputs(4660) <= b;
    layer2_outputs(4661) <= not (a xor b);
    layer2_outputs(4662) <= not b;
    layer2_outputs(4663) <= a;
    layer2_outputs(4664) <= a or b;
    layer2_outputs(4665) <= b and not a;
    layer2_outputs(4666) <= a or b;
    layer2_outputs(4667) <= a xor b;
    layer2_outputs(4668) <= b;
    layer2_outputs(4669) <= a or b;
    layer2_outputs(4670) <= a and not b;
    layer2_outputs(4671) <= not a;
    layer2_outputs(4672) <= not a;
    layer2_outputs(4673) <= a;
    layer2_outputs(4674) <= not a;
    layer2_outputs(4675) <= not (a or b);
    layer2_outputs(4676) <= not b;
    layer2_outputs(4677) <= a;
    layer2_outputs(4678) <= not (a and b);
    layer2_outputs(4679) <= a or b;
    layer2_outputs(4680) <= not a;
    layer2_outputs(4681) <= not (a xor b);
    layer2_outputs(4682) <= not a;
    layer2_outputs(4683) <= a or b;
    layer2_outputs(4684) <= not a;
    layer2_outputs(4685) <= a xor b;
    layer2_outputs(4686) <= not (a and b);
    layer2_outputs(4687) <= not b;
    layer2_outputs(4688) <= not b or a;
    layer2_outputs(4689) <= b and not a;
    layer2_outputs(4690) <= b;
    layer2_outputs(4691) <= not (a or b);
    layer2_outputs(4692) <= not (a or b);
    layer2_outputs(4693) <= a xor b;
    layer2_outputs(4694) <= a and not b;
    layer2_outputs(4695) <= not a or b;
    layer2_outputs(4696) <= a and not b;
    layer2_outputs(4697) <= a xor b;
    layer2_outputs(4698) <= a;
    layer2_outputs(4699) <= a and b;
    layer2_outputs(4700) <= b and not a;
    layer2_outputs(4701) <= not a;
    layer2_outputs(4702) <= not b or a;
    layer2_outputs(4703) <= not (a and b);
    layer2_outputs(4704) <= b and not a;
    layer2_outputs(4705) <= a;
    layer2_outputs(4706) <= a;
    layer2_outputs(4707) <= b;
    layer2_outputs(4708) <= a and b;
    layer2_outputs(4709) <= not (a or b);
    layer2_outputs(4710) <= b and not a;
    layer2_outputs(4711) <= not (a and b);
    layer2_outputs(4712) <= a or b;
    layer2_outputs(4713) <= not (a or b);
    layer2_outputs(4714) <= a xor b;
    layer2_outputs(4715) <= a xor b;
    layer2_outputs(4716) <= a and not b;
    layer2_outputs(4717) <= not b or a;
    layer2_outputs(4718) <= not (a xor b);
    layer2_outputs(4719) <= not (a or b);
    layer2_outputs(4720) <= a xor b;
    layer2_outputs(4721) <= not a or b;
    layer2_outputs(4722) <= a or b;
    layer2_outputs(4723) <= not b;
    layer2_outputs(4724) <= not (a xor b);
    layer2_outputs(4725) <= b;
    layer2_outputs(4726) <= a and not b;
    layer2_outputs(4727) <= a and b;
    layer2_outputs(4728) <= b;
    layer2_outputs(4729) <= a and b;
    layer2_outputs(4730) <= b;
    layer2_outputs(4731) <= a xor b;
    layer2_outputs(4732) <= a or b;
    layer2_outputs(4733) <= a and b;
    layer2_outputs(4734) <= not (a or b);
    layer2_outputs(4735) <= a;
    layer2_outputs(4736) <= b;
    layer2_outputs(4737) <= not b or a;
    layer2_outputs(4738) <= not b or a;
    layer2_outputs(4739) <= not b;
    layer2_outputs(4740) <= b;
    layer2_outputs(4741) <= not a;
    layer2_outputs(4742) <= not (a or b);
    layer2_outputs(4743) <= a;
    layer2_outputs(4744) <= a and b;
    layer2_outputs(4745) <= not b or a;
    layer2_outputs(4746) <= b;
    layer2_outputs(4747) <= b;
    layer2_outputs(4748) <= b and not a;
    layer2_outputs(4749) <= a xor b;
    layer2_outputs(4750) <= not (a and b);
    layer2_outputs(4751) <= b;
    layer2_outputs(4752) <= not b;
    layer2_outputs(4753) <= a and not b;
    layer2_outputs(4754) <= a xor b;
    layer2_outputs(4755) <= b and not a;
    layer2_outputs(4756) <= a or b;
    layer2_outputs(4757) <= not (a and b);
    layer2_outputs(4758) <= not (a or b);
    layer2_outputs(4759) <= 1'b1;
    layer2_outputs(4760) <= not a or b;
    layer2_outputs(4761) <= a and b;
    layer2_outputs(4762) <= not (a and b);
    layer2_outputs(4763) <= a and not b;
    layer2_outputs(4764) <= not b;
    layer2_outputs(4765) <= not (a xor b);
    layer2_outputs(4766) <= not b or a;
    layer2_outputs(4767) <= b and not a;
    layer2_outputs(4768) <= not b;
    layer2_outputs(4769) <= a;
    layer2_outputs(4770) <= not b;
    layer2_outputs(4771) <= not a;
    layer2_outputs(4772) <= a xor b;
    layer2_outputs(4773) <= not (a and b);
    layer2_outputs(4774) <= a xor b;
    layer2_outputs(4775) <= b and not a;
    layer2_outputs(4776) <= not b;
    layer2_outputs(4777) <= b and not a;
    layer2_outputs(4778) <= not b;
    layer2_outputs(4779) <= not b or a;
    layer2_outputs(4780) <= not a or b;
    layer2_outputs(4781) <= not b or a;
    layer2_outputs(4782) <= not b;
    layer2_outputs(4783) <= not b or a;
    layer2_outputs(4784) <= not (a xor b);
    layer2_outputs(4785) <= b and not a;
    layer2_outputs(4786) <= a;
    layer2_outputs(4787) <= b;
    layer2_outputs(4788) <= 1'b0;
    layer2_outputs(4789) <= not (a or b);
    layer2_outputs(4790) <= not a or b;
    layer2_outputs(4791) <= not (a or b);
    layer2_outputs(4792) <= a xor b;
    layer2_outputs(4793) <= b and not a;
    layer2_outputs(4794) <= not (a and b);
    layer2_outputs(4795) <= not b;
    layer2_outputs(4796) <= not (a and b);
    layer2_outputs(4797) <= not (a xor b);
    layer2_outputs(4798) <= not b;
    layer2_outputs(4799) <= a;
    layer2_outputs(4800) <= not (a or b);
    layer2_outputs(4801) <= not b;
    layer2_outputs(4802) <= not (a and b);
    layer2_outputs(4803) <= b and not a;
    layer2_outputs(4804) <= not (a or b);
    layer2_outputs(4805) <= b;
    layer2_outputs(4806) <= a and not b;
    layer2_outputs(4807) <= b;
    layer2_outputs(4808) <= a;
    layer2_outputs(4809) <= b;
    layer2_outputs(4810) <= a;
    layer2_outputs(4811) <= b;
    layer2_outputs(4812) <= a and b;
    layer2_outputs(4813) <= not a;
    layer2_outputs(4814) <= a;
    layer2_outputs(4815) <= not a;
    layer2_outputs(4816) <= not (a xor b);
    layer2_outputs(4817) <= not a or b;
    layer2_outputs(4818) <= not a;
    layer2_outputs(4819) <= not b;
    layer2_outputs(4820) <= a or b;
    layer2_outputs(4821) <= not a or b;
    layer2_outputs(4822) <= not b;
    layer2_outputs(4823) <= not a or b;
    layer2_outputs(4824) <= not a;
    layer2_outputs(4825) <= not a;
    layer2_outputs(4826) <= not a;
    layer2_outputs(4827) <= not (a xor b);
    layer2_outputs(4828) <= not b;
    layer2_outputs(4829) <= not b or a;
    layer2_outputs(4830) <= not a;
    layer2_outputs(4831) <= not (a or b);
    layer2_outputs(4832) <= not (a and b);
    layer2_outputs(4833) <= a xor b;
    layer2_outputs(4834) <= not b or a;
    layer2_outputs(4835) <= b;
    layer2_outputs(4836) <= a or b;
    layer2_outputs(4837) <= b and not a;
    layer2_outputs(4838) <= 1'b0;
    layer2_outputs(4839) <= not b;
    layer2_outputs(4840) <= a and b;
    layer2_outputs(4841) <= a and not b;
    layer2_outputs(4842) <= a xor b;
    layer2_outputs(4843) <= a and not b;
    layer2_outputs(4844) <= b;
    layer2_outputs(4845) <= a and not b;
    layer2_outputs(4846) <= a and b;
    layer2_outputs(4847) <= not (a xor b);
    layer2_outputs(4848) <= b and not a;
    layer2_outputs(4849) <= a and not b;
    layer2_outputs(4850) <= b;
    layer2_outputs(4851) <= not b;
    layer2_outputs(4852) <= a or b;
    layer2_outputs(4853) <= a;
    layer2_outputs(4854) <= not (a xor b);
    layer2_outputs(4855) <= not (a or b);
    layer2_outputs(4856) <= not b;
    layer2_outputs(4857) <= a or b;
    layer2_outputs(4858) <= b and not a;
    layer2_outputs(4859) <= b;
    layer2_outputs(4860) <= not b or a;
    layer2_outputs(4861) <= not a;
    layer2_outputs(4862) <= a;
    layer2_outputs(4863) <= a and not b;
    layer2_outputs(4864) <= not a;
    layer2_outputs(4865) <= b and not a;
    layer2_outputs(4866) <= a;
    layer2_outputs(4867) <= a;
    layer2_outputs(4868) <= a or b;
    layer2_outputs(4869) <= a;
    layer2_outputs(4870) <= a;
    layer2_outputs(4871) <= not a;
    layer2_outputs(4872) <= not (a and b);
    layer2_outputs(4873) <= not (a or b);
    layer2_outputs(4874) <= a and b;
    layer2_outputs(4875) <= not a or b;
    layer2_outputs(4876) <= not b;
    layer2_outputs(4877) <= not (a xor b);
    layer2_outputs(4878) <= not a or b;
    layer2_outputs(4879) <= a;
    layer2_outputs(4880) <= a;
    layer2_outputs(4881) <= a;
    layer2_outputs(4882) <= a and not b;
    layer2_outputs(4883) <= not (a or b);
    layer2_outputs(4884) <= not a;
    layer2_outputs(4885) <= a;
    layer2_outputs(4886) <= a and not b;
    layer2_outputs(4887) <= not b;
    layer2_outputs(4888) <= a and not b;
    layer2_outputs(4889) <= not a;
    layer2_outputs(4890) <= not (a or b);
    layer2_outputs(4891) <= a and b;
    layer2_outputs(4892) <= a or b;
    layer2_outputs(4893) <= not b;
    layer2_outputs(4894) <= b and not a;
    layer2_outputs(4895) <= 1'b0;
    layer2_outputs(4896) <= not b;
    layer2_outputs(4897) <= a and b;
    layer2_outputs(4898) <= not b or a;
    layer2_outputs(4899) <= a xor b;
    layer2_outputs(4900) <= a or b;
    layer2_outputs(4901) <= 1'b1;
    layer2_outputs(4902) <= a xor b;
    layer2_outputs(4903) <= not (a xor b);
    layer2_outputs(4904) <= a;
    layer2_outputs(4905) <= a and b;
    layer2_outputs(4906) <= not b or a;
    layer2_outputs(4907) <= a or b;
    layer2_outputs(4908) <= not (a xor b);
    layer2_outputs(4909) <= b;
    layer2_outputs(4910) <= a;
    layer2_outputs(4911) <= a xor b;
    layer2_outputs(4912) <= not (a and b);
    layer2_outputs(4913) <= not b or a;
    layer2_outputs(4914) <= b;
    layer2_outputs(4915) <= not b or a;
    layer2_outputs(4916) <= not (a xor b);
    layer2_outputs(4917) <= not a;
    layer2_outputs(4918) <= not (a or b);
    layer2_outputs(4919) <= not a;
    layer2_outputs(4920) <= b;
    layer2_outputs(4921) <= b;
    layer2_outputs(4922) <= not (a and b);
    layer2_outputs(4923) <= not (a or b);
    layer2_outputs(4924) <= not a or b;
    layer2_outputs(4925) <= b;
    layer2_outputs(4926) <= 1'b1;
    layer2_outputs(4927) <= a;
    layer2_outputs(4928) <= a xor b;
    layer2_outputs(4929) <= not (a xor b);
    layer2_outputs(4930) <= not b;
    layer2_outputs(4931) <= a and b;
    layer2_outputs(4932) <= a and not b;
    layer2_outputs(4933) <= b and not a;
    layer2_outputs(4934) <= not (a and b);
    layer2_outputs(4935) <= not a or b;
    layer2_outputs(4936) <= b;
    layer2_outputs(4937) <= not (a or b);
    layer2_outputs(4938) <= not (a xor b);
    layer2_outputs(4939) <= not a or b;
    layer2_outputs(4940) <= not b or a;
    layer2_outputs(4941) <= not a;
    layer2_outputs(4942) <= a;
    layer2_outputs(4943) <= a or b;
    layer2_outputs(4944) <= 1'b1;
    layer2_outputs(4945) <= a and not b;
    layer2_outputs(4946) <= a and not b;
    layer2_outputs(4947) <= a and b;
    layer2_outputs(4948) <= not (a xor b);
    layer2_outputs(4949) <= a and not b;
    layer2_outputs(4950) <= a or b;
    layer2_outputs(4951) <= b;
    layer2_outputs(4952) <= a xor b;
    layer2_outputs(4953) <= not (a xor b);
    layer2_outputs(4954) <= b and not a;
    layer2_outputs(4955) <= b and not a;
    layer2_outputs(4956) <= not (a xor b);
    layer2_outputs(4957) <= not a;
    layer2_outputs(4958) <= not a or b;
    layer2_outputs(4959) <= a and not b;
    layer2_outputs(4960) <= a and not b;
    layer2_outputs(4961) <= not a or b;
    layer2_outputs(4962) <= a and not b;
    layer2_outputs(4963) <= a or b;
    layer2_outputs(4964) <= not a;
    layer2_outputs(4965) <= b;
    layer2_outputs(4966) <= not b or a;
    layer2_outputs(4967) <= a and b;
    layer2_outputs(4968) <= not b;
    layer2_outputs(4969) <= a;
    layer2_outputs(4970) <= not b or a;
    layer2_outputs(4971) <= a xor b;
    layer2_outputs(4972) <= not a or b;
    layer2_outputs(4973) <= not a or b;
    layer2_outputs(4974) <= b;
    layer2_outputs(4975) <= a and b;
    layer2_outputs(4976) <= a or b;
    layer2_outputs(4977) <= a;
    layer2_outputs(4978) <= b and not a;
    layer2_outputs(4979) <= b and not a;
    layer2_outputs(4980) <= not a;
    layer2_outputs(4981) <= not a;
    layer2_outputs(4982) <= a xor b;
    layer2_outputs(4983) <= b;
    layer2_outputs(4984) <= a and b;
    layer2_outputs(4985) <= not b or a;
    layer2_outputs(4986) <= b;
    layer2_outputs(4987) <= not (a and b);
    layer2_outputs(4988) <= not (a and b);
    layer2_outputs(4989) <= a xor b;
    layer2_outputs(4990) <= b;
    layer2_outputs(4991) <= not b or a;
    layer2_outputs(4992) <= not a or b;
    layer2_outputs(4993) <= not a;
    layer2_outputs(4994) <= not b;
    layer2_outputs(4995) <= a and not b;
    layer2_outputs(4996) <= a;
    layer2_outputs(4997) <= not (a and b);
    layer2_outputs(4998) <= a or b;
    layer2_outputs(4999) <= not (a and b);
    layer2_outputs(5000) <= a or b;
    layer2_outputs(5001) <= b and not a;
    layer2_outputs(5002) <= not (a or b);
    layer2_outputs(5003) <= not b;
    layer2_outputs(5004) <= a xor b;
    layer2_outputs(5005) <= a xor b;
    layer2_outputs(5006) <= a and not b;
    layer2_outputs(5007) <= not b;
    layer2_outputs(5008) <= not a;
    layer2_outputs(5009) <= not (a or b);
    layer2_outputs(5010) <= a xor b;
    layer2_outputs(5011) <= not b or a;
    layer2_outputs(5012) <= not b;
    layer2_outputs(5013) <= b and not a;
    layer2_outputs(5014) <= not a;
    layer2_outputs(5015) <= not b;
    layer2_outputs(5016) <= a and b;
    layer2_outputs(5017) <= not a or b;
    layer2_outputs(5018) <= a and b;
    layer2_outputs(5019) <= a;
    layer2_outputs(5020) <= not (a or b);
    layer2_outputs(5021) <= not b;
    layer2_outputs(5022) <= a xor b;
    layer2_outputs(5023) <= not a or b;
    layer2_outputs(5024) <= b;
    layer2_outputs(5025) <= a;
    layer2_outputs(5026) <= not b or a;
    layer2_outputs(5027) <= not a or b;
    layer2_outputs(5028) <= a and not b;
    layer2_outputs(5029) <= not a;
    layer2_outputs(5030) <= b and not a;
    layer2_outputs(5031) <= not (a and b);
    layer2_outputs(5032) <= not (a or b);
    layer2_outputs(5033) <= not (a or b);
    layer2_outputs(5034) <= not (a or b);
    layer2_outputs(5035) <= not b;
    layer2_outputs(5036) <= not b;
    layer2_outputs(5037) <= a;
    layer2_outputs(5038) <= a;
    layer2_outputs(5039) <= a and not b;
    layer2_outputs(5040) <= a xor b;
    layer2_outputs(5041) <= b and not a;
    layer2_outputs(5042) <= not (a xor b);
    layer2_outputs(5043) <= b;
    layer2_outputs(5044) <= not a or b;
    layer2_outputs(5045) <= b;
    layer2_outputs(5046) <= b;
    layer2_outputs(5047) <= not (a and b);
    layer2_outputs(5048) <= not a or b;
    layer2_outputs(5049) <= not (a xor b);
    layer2_outputs(5050) <= b;
    layer2_outputs(5051) <= a and not b;
    layer2_outputs(5052) <= not (a and b);
    layer2_outputs(5053) <= a;
    layer2_outputs(5054) <= not (a and b);
    layer2_outputs(5055) <= not (a or b);
    layer2_outputs(5056) <= not (a xor b);
    layer2_outputs(5057) <= a and not b;
    layer2_outputs(5058) <= not a or b;
    layer2_outputs(5059) <= a xor b;
    layer2_outputs(5060) <= a and b;
    layer2_outputs(5061) <= not b;
    layer2_outputs(5062) <= a xor b;
    layer2_outputs(5063) <= not a or b;
    layer2_outputs(5064) <= 1'b0;
    layer2_outputs(5065) <= a and not b;
    layer2_outputs(5066) <= not a;
    layer2_outputs(5067) <= not a;
    layer2_outputs(5068) <= a;
    layer2_outputs(5069) <= not b;
    layer2_outputs(5070) <= not b;
    layer2_outputs(5071) <= not b;
    layer2_outputs(5072) <= not a;
    layer2_outputs(5073) <= a or b;
    layer2_outputs(5074) <= not a or b;
    layer2_outputs(5075) <= a and b;
    layer2_outputs(5076) <= a and not b;
    layer2_outputs(5077) <= a xor b;
    layer2_outputs(5078) <= not (a xor b);
    layer2_outputs(5079) <= a and not b;
    layer2_outputs(5080) <= a;
    layer2_outputs(5081) <= not (a or b);
    layer2_outputs(5082) <= a and not b;
    layer2_outputs(5083) <= not (a and b);
    layer2_outputs(5084) <= not b or a;
    layer2_outputs(5085) <= not (a xor b);
    layer2_outputs(5086) <= a xor b;
    layer2_outputs(5087) <= not b or a;
    layer2_outputs(5088) <= not a;
    layer2_outputs(5089) <= b and not a;
    layer2_outputs(5090) <= not a or b;
    layer2_outputs(5091) <= b;
    layer2_outputs(5092) <= b;
    layer2_outputs(5093) <= a;
    layer2_outputs(5094) <= not a or b;
    layer2_outputs(5095) <= not (a or b);
    layer2_outputs(5096) <= not (a or b);
    layer2_outputs(5097) <= not b;
    layer2_outputs(5098) <= a;
    layer2_outputs(5099) <= b and not a;
    layer2_outputs(5100) <= a and not b;
    layer2_outputs(5101) <= not (a xor b);
    layer2_outputs(5102) <= a and not b;
    layer2_outputs(5103) <= not b or a;
    layer2_outputs(5104) <= a xor b;
    layer2_outputs(5105) <= b;
    layer2_outputs(5106) <= b;
    layer2_outputs(5107) <= a and not b;
    layer2_outputs(5108) <= not (a xor b);
    layer2_outputs(5109) <= a xor b;
    layer2_outputs(5110) <= a;
    layer2_outputs(5111) <= not a or b;
    layer2_outputs(5112) <= not (a or b);
    layer2_outputs(5113) <= not a;
    layer2_outputs(5114) <= not (a or b);
    layer2_outputs(5115) <= not a or b;
    layer2_outputs(5116) <= a;
    layer2_outputs(5117) <= not a;
    layer2_outputs(5118) <= a and b;
    layer2_outputs(5119) <= 1'b1;
    outputs(0) <= not (a or b);
    outputs(1) <= a and not b;
    outputs(2) <= a and b;
    outputs(3) <= b;
    outputs(4) <= not b;
    outputs(5) <= a xor b;
    outputs(6) <= not (a or b);
    outputs(7) <= not (a and b);
    outputs(8) <= not b or a;
    outputs(9) <= a xor b;
    outputs(10) <= a;
    outputs(11) <= b;
    outputs(12) <= a and b;
    outputs(13) <= a xor b;
    outputs(14) <= b and not a;
    outputs(15) <= not b;
    outputs(16) <= b and not a;
    outputs(17) <= not a;
    outputs(18) <= b;
    outputs(19) <= not b;
    outputs(20) <= not (a xor b);
    outputs(21) <= a and not b;
    outputs(22) <= b;
    outputs(23) <= a;
    outputs(24) <= a xor b;
    outputs(25) <= a;
    outputs(26) <= a and b;
    outputs(27) <= a and not b;
    outputs(28) <= b;
    outputs(29) <= a and not b;
    outputs(30) <= not b or a;
    outputs(31) <= not b;
    outputs(32) <= not b;
    outputs(33) <= b and not a;
    outputs(34) <= a or b;
    outputs(35) <= a;
    outputs(36) <= not a;
    outputs(37) <= not b;
    outputs(38) <= not b;
    outputs(39) <= a;
    outputs(40) <= a;
    outputs(41) <= not b or a;
    outputs(42) <= b;
    outputs(43) <= not b;
    outputs(44) <= a and not b;
    outputs(45) <= b;
    outputs(46) <= b;
    outputs(47) <= not b or a;
    outputs(48) <= a and b;
    outputs(49) <= not b;
    outputs(50) <= b;
    outputs(51) <= a;
    outputs(52) <= a;
    outputs(53) <= a;
    outputs(54) <= a and not b;
    outputs(55) <= a and not b;
    outputs(56) <= not b or a;
    outputs(57) <= a and b;
    outputs(58) <= not (a xor b);
    outputs(59) <= a and b;
    outputs(60) <= not (a and b);
    outputs(61) <= a;
    outputs(62) <= a;
    outputs(63) <= not (a xor b);
    outputs(64) <= a;
    outputs(65) <= not (a xor b);
    outputs(66) <= not (a or b);
    outputs(67) <= not a;
    outputs(68) <= not b or a;
    outputs(69) <= b and not a;
    outputs(70) <= not b;
    outputs(71) <= a;
    outputs(72) <= a and b;
    outputs(73) <= not a or b;
    outputs(74) <= not a;
    outputs(75) <= a;
    outputs(76) <= a and b;
    outputs(77) <= not b;
    outputs(78) <= a;
    outputs(79) <= not (a xor b);
    outputs(80) <= a;
    outputs(81) <= not a;
    outputs(82) <= not b;
    outputs(83) <= a xor b;
    outputs(84) <= a and not b;
    outputs(85) <= a xor b;
    outputs(86) <= not b;
    outputs(87) <= not a;
    outputs(88) <= a and not b;
    outputs(89) <= not a;
    outputs(90) <= a;
    outputs(91) <= b;
    outputs(92) <= not (a and b);
    outputs(93) <= a;
    outputs(94) <= a and b;
    outputs(95) <= b;
    outputs(96) <= b;
    outputs(97) <= not (a xor b);
    outputs(98) <= b and not a;
    outputs(99) <= a;
    outputs(100) <= a xor b;
    outputs(101) <= a xor b;
    outputs(102) <= not a or b;
    outputs(103) <= not b;
    outputs(104) <= b and not a;
    outputs(105) <= b;
    outputs(106) <= a;
    outputs(107) <= not a;
    outputs(108) <= not (a and b);
    outputs(109) <= not a;
    outputs(110) <= a and b;
    outputs(111) <= b;
    outputs(112) <= not (a and b);
    outputs(113) <= a xor b;
    outputs(114) <= a;
    outputs(115) <= a;
    outputs(116) <= a or b;
    outputs(117) <= not b;
    outputs(118) <= not b or a;
    outputs(119) <= not b or a;
    outputs(120) <= b;
    outputs(121) <= b;
    outputs(122) <= not b;
    outputs(123) <= b and not a;
    outputs(124) <= not (a xor b);
    outputs(125) <= a;
    outputs(126) <= not a;
    outputs(127) <= b;
    outputs(128) <= not a or b;
    outputs(129) <= a;
    outputs(130) <= a xor b;
    outputs(131) <= not b or a;
    outputs(132) <= not a;
    outputs(133) <= b;
    outputs(134) <= not a;
    outputs(135) <= a xor b;
    outputs(136) <= a;
    outputs(137) <= not a;
    outputs(138) <= not b or a;
    outputs(139) <= not a;
    outputs(140) <= b;
    outputs(141) <= a and not b;
    outputs(142) <= b;
    outputs(143) <= not a or b;
    outputs(144) <= not a;
    outputs(145) <= b;
    outputs(146) <= b;
    outputs(147) <= not a;
    outputs(148) <= b;
    outputs(149) <= not (a xor b);
    outputs(150) <= not (a or b);
    outputs(151) <= not b;
    outputs(152) <= a and b;
    outputs(153) <= a;
    outputs(154) <= not b;
    outputs(155) <= not (a or b);
    outputs(156) <= not b;
    outputs(157) <= a and b;
    outputs(158) <= not a;
    outputs(159) <= a;
    outputs(160) <= not a;
    outputs(161) <= a and b;
    outputs(162) <= b and not a;
    outputs(163) <= a;
    outputs(164) <= b;
    outputs(165) <= not a;
    outputs(166) <= not a;
    outputs(167) <= not (a or b);
    outputs(168) <= a and b;
    outputs(169) <= b;
    outputs(170) <= not a;
    outputs(171) <= a xor b;
    outputs(172) <= not (a or b);
    outputs(173) <= b;
    outputs(174) <= not b or a;
    outputs(175) <= not (a xor b);
    outputs(176) <= not a;
    outputs(177) <= a and b;
    outputs(178) <= a xor b;
    outputs(179) <= not (a xor b);
    outputs(180) <= not (a xor b);
    outputs(181) <= b;
    outputs(182) <= a and b;
    outputs(183) <= a and b;
    outputs(184) <= not (a or b);
    outputs(185) <= a;
    outputs(186) <= not a or b;
    outputs(187) <= b and not a;
    outputs(188) <= a;
    outputs(189) <= a and not b;
    outputs(190) <= not (a xor b);
    outputs(191) <= a and b;
    outputs(192) <= a and b;
    outputs(193) <= not (a xor b);
    outputs(194) <= a xor b;
    outputs(195) <= not (a xor b);
    outputs(196) <= b;
    outputs(197) <= b and not a;
    outputs(198) <= a and b;
    outputs(199) <= not a or b;
    outputs(200) <= not a;
    outputs(201) <= a and not b;
    outputs(202) <= b;
    outputs(203) <= a xor b;
    outputs(204) <= a xor b;
    outputs(205) <= not a or b;
    outputs(206) <= b;
    outputs(207) <= b;
    outputs(208) <= a and b;
    outputs(209) <= not (a xor b);
    outputs(210) <= b;
    outputs(211) <= a xor b;
    outputs(212) <= not b;
    outputs(213) <= not a;
    outputs(214) <= a and not b;
    outputs(215) <= not a;
    outputs(216) <= not (a or b);
    outputs(217) <= b;
    outputs(218) <= a;
    outputs(219) <= a and not b;
    outputs(220) <= not (a or b);
    outputs(221) <= not (a and b);
    outputs(222) <= not (a or b);
    outputs(223) <= not a;
    outputs(224) <= not (a and b);
    outputs(225) <= not (a or b);
    outputs(226) <= not (a or b);
    outputs(227) <= a and b;
    outputs(228) <= a;
    outputs(229) <= b;
    outputs(230) <= b;
    outputs(231) <= a and not b;
    outputs(232) <= not b;
    outputs(233) <= a and b;
    outputs(234) <= a and b;
    outputs(235) <= b;
    outputs(236) <= a and b;
    outputs(237) <= not b;
    outputs(238) <= not (a xor b);
    outputs(239) <= b;
    outputs(240) <= not a;
    outputs(241) <= not a;
    outputs(242) <= not b;
    outputs(243) <= a and b;
    outputs(244) <= a and b;
    outputs(245) <= not (a and b);
    outputs(246) <= not a;
    outputs(247) <= a and b;
    outputs(248) <= not a or b;
    outputs(249) <= not (a or b);
    outputs(250) <= not (a and b);
    outputs(251) <= not (a xor b);
    outputs(252) <= b and not a;
    outputs(253) <= a xor b;
    outputs(254) <= b;
    outputs(255) <= not b;
    outputs(256) <= a and b;
    outputs(257) <= a and b;
    outputs(258) <= b and not a;
    outputs(259) <= a;
    outputs(260) <= not (a or b);
    outputs(261) <= not a or b;
    outputs(262) <= not b;
    outputs(263) <= a;
    outputs(264) <= not b;
    outputs(265) <= a xor b;
    outputs(266) <= not a;
    outputs(267) <= not b or a;
    outputs(268) <= b;
    outputs(269) <= not a or b;
    outputs(270) <= not (a or b);
    outputs(271) <= not a;
    outputs(272) <= not a;
    outputs(273) <= not b;
    outputs(274) <= a xor b;
    outputs(275) <= a;
    outputs(276) <= not b;
    outputs(277) <= a and b;
    outputs(278) <= b;
    outputs(279) <= not a;
    outputs(280) <= not b;
    outputs(281) <= not b;
    outputs(282) <= not b;
    outputs(283) <= not b;
    outputs(284) <= not (a or b);
    outputs(285) <= not a;
    outputs(286) <= not (a xor b);
    outputs(287) <= a and not b;
    outputs(288) <= not a;
    outputs(289) <= b;
    outputs(290) <= not b;
    outputs(291) <= a or b;
    outputs(292) <= a;
    outputs(293) <= b;
    outputs(294) <= not a or b;
    outputs(295) <= not a;
    outputs(296) <= b and not a;
    outputs(297) <= not a;
    outputs(298) <= not (a or b);
    outputs(299) <= a;
    outputs(300) <= a xor b;
    outputs(301) <= not b;
    outputs(302) <= b;
    outputs(303) <= a and not b;
    outputs(304) <= a;
    outputs(305) <= a;
    outputs(306) <= not b;
    outputs(307) <= a;
    outputs(308) <= a and b;
    outputs(309) <= not a;
    outputs(310) <= b;
    outputs(311) <= not b;
    outputs(312) <= b;
    outputs(313) <= not (a and b);
    outputs(314) <= a;
    outputs(315) <= not b or a;
    outputs(316) <= a xor b;
    outputs(317) <= not (a and b);
    outputs(318) <= a and b;
    outputs(319) <= a xor b;
    outputs(320) <= a xor b;
    outputs(321) <= a and not b;
    outputs(322) <= not a;
    outputs(323) <= a;
    outputs(324) <= not b;
    outputs(325) <= not b or a;
    outputs(326) <= not (a and b);
    outputs(327) <= not (a and b);
    outputs(328) <= b and not a;
    outputs(329) <= a;
    outputs(330) <= not a or b;
    outputs(331) <= not (a or b);
    outputs(332) <= b;
    outputs(333) <= b;
    outputs(334) <= a and not b;
    outputs(335) <= not a;
    outputs(336) <= not b;
    outputs(337) <= not b or a;
    outputs(338) <= b and not a;
    outputs(339) <= a;
    outputs(340) <= not a;
    outputs(341) <= not (a and b);
    outputs(342) <= not b;
    outputs(343) <= a xor b;
    outputs(344) <= not b;
    outputs(345) <= not (a xor b);
    outputs(346) <= not a or b;
    outputs(347) <= not b;
    outputs(348) <= not (a xor b);
    outputs(349) <= not b;
    outputs(350) <= a and b;
    outputs(351) <= b;
    outputs(352) <= a or b;
    outputs(353) <= a and not b;
    outputs(354) <= a xor b;
    outputs(355) <= a;
    outputs(356) <= not a;
    outputs(357) <= a and not b;
    outputs(358) <= b;
    outputs(359) <= a xor b;
    outputs(360) <= not b;
    outputs(361) <= b;
    outputs(362) <= b;
    outputs(363) <= a;
    outputs(364) <= not b;
    outputs(365) <= not b;
    outputs(366) <= not a;
    outputs(367) <= b and not a;
    outputs(368) <= a or b;
    outputs(369) <= not a;
    outputs(370) <= a;
    outputs(371) <= a or b;
    outputs(372) <= not (a xor b);
    outputs(373) <= a;
    outputs(374) <= not a;
    outputs(375) <= b;
    outputs(376) <= not b;
    outputs(377) <= b;
    outputs(378) <= a;
    outputs(379) <= a and b;
    outputs(380) <= not a;
    outputs(381) <= a and not b;
    outputs(382) <= b;
    outputs(383) <= a;
    outputs(384) <= a xor b;
    outputs(385) <= not (a and b);
    outputs(386) <= not a;
    outputs(387) <= a;
    outputs(388) <= a and not b;
    outputs(389) <= a;
    outputs(390) <= a and b;
    outputs(391) <= not a;
    outputs(392) <= not a;
    outputs(393) <= not a;
    outputs(394) <= a;
    outputs(395) <= not b;
    outputs(396) <= b;
    outputs(397) <= not b;
    outputs(398) <= not b;
    outputs(399) <= a xor b;
    outputs(400) <= a;
    outputs(401) <= a;
    outputs(402) <= not (a xor b);
    outputs(403) <= not (a and b);
    outputs(404) <= not b;
    outputs(405) <= a xor b;
    outputs(406) <= not (a or b);
    outputs(407) <= not (a xor b);
    outputs(408) <= not b;
    outputs(409) <= not a;
    outputs(410) <= not a;
    outputs(411) <= not a;
    outputs(412) <= not b;
    outputs(413) <= not (a or b);
    outputs(414) <= a and not b;
    outputs(415) <= b;
    outputs(416) <= not b;
    outputs(417) <= not (a xor b);
    outputs(418) <= b;
    outputs(419) <= not b;
    outputs(420) <= not a;
    outputs(421) <= not b;
    outputs(422) <= not b;
    outputs(423) <= not b;
    outputs(424) <= a;
    outputs(425) <= a and b;
    outputs(426) <= not b;
    outputs(427) <= b;
    outputs(428) <= b and not a;
    outputs(429) <= a xor b;
    outputs(430) <= a or b;
    outputs(431) <= a;
    outputs(432) <= not b;
    outputs(433) <= a and b;
    outputs(434) <= not b;
    outputs(435) <= not a;
    outputs(436) <= not b;
    outputs(437) <= not b;
    outputs(438) <= a and not b;
    outputs(439) <= not a;
    outputs(440) <= not a;
    outputs(441) <= not b or a;
    outputs(442) <= a;
    outputs(443) <= b and not a;
    outputs(444) <= not a;
    outputs(445) <= not (a xor b);
    outputs(446) <= b;
    outputs(447) <= a xor b;
    outputs(448) <= not a;
    outputs(449) <= a;
    outputs(450) <= b;
    outputs(451) <= not a;
    outputs(452) <= a xor b;
    outputs(453) <= a and not b;
    outputs(454) <= not a;
    outputs(455) <= not b;
    outputs(456) <= a and not b;
    outputs(457) <= not b;
    outputs(458) <= not a;
    outputs(459) <= a xor b;
    outputs(460) <= a xor b;
    outputs(461) <= not a or b;
    outputs(462) <= a;
    outputs(463) <= not a;
    outputs(464) <= a and b;
    outputs(465) <= not b;
    outputs(466) <= b;
    outputs(467) <= not (a or b);
    outputs(468) <= a xor b;
    outputs(469) <= not b;
    outputs(470) <= not a;
    outputs(471) <= a;
    outputs(472) <= not (a or b);
    outputs(473) <= not a;
    outputs(474) <= b and not a;
    outputs(475) <= a xor b;
    outputs(476) <= not a;
    outputs(477) <= a or b;
    outputs(478) <= not b or a;
    outputs(479) <= not a or b;
    outputs(480) <= not (a or b);
    outputs(481) <= b;
    outputs(482) <= a or b;
    outputs(483) <= a and b;
    outputs(484) <= not b;
    outputs(485) <= not a;
    outputs(486) <= a;
    outputs(487) <= not a or b;
    outputs(488) <= not a or b;
    outputs(489) <= b and not a;
    outputs(490) <= b;
    outputs(491) <= not b;
    outputs(492) <= b;
    outputs(493) <= not a;
    outputs(494) <= a xor b;
    outputs(495) <= b;
    outputs(496) <= a;
    outputs(497) <= a;
    outputs(498) <= b and not a;
    outputs(499) <= not b;
    outputs(500) <= a and not b;
    outputs(501) <= not a;
    outputs(502) <= not b or a;
    outputs(503) <= not a;
    outputs(504) <= not b;
    outputs(505) <= a xor b;
    outputs(506) <= a;
    outputs(507) <= a xor b;
    outputs(508) <= not (a xor b);
    outputs(509) <= not b;
    outputs(510) <= a;
    outputs(511) <= not (a or b);
    outputs(512) <= b;
    outputs(513) <= b;
    outputs(514) <= not a;
    outputs(515) <= not (a or b);
    outputs(516) <= a xor b;
    outputs(517) <= a and b;
    outputs(518) <= a and not b;
    outputs(519) <= a and not b;
    outputs(520) <= not (a or b);
    outputs(521) <= a and b;
    outputs(522) <= a;
    outputs(523) <= not a;
    outputs(524) <= not (a or b);
    outputs(525) <= a and not b;
    outputs(526) <= not (a or b);
    outputs(527) <= b and not a;
    outputs(528) <= not b;
    outputs(529) <= a xor b;
    outputs(530) <= a and not b;
    outputs(531) <= not (a or b);
    outputs(532) <= not (a or b);
    outputs(533) <= not (a or b);
    outputs(534) <= a xor b;
    outputs(535) <= not (a or b);
    outputs(536) <= not (a or b);
    outputs(537) <= b and not a;
    outputs(538) <= not (a or b);
    outputs(539) <= a;
    outputs(540) <= a xor b;
    outputs(541) <= b;
    outputs(542) <= not a;
    outputs(543) <= b;
    outputs(544) <= not (a or b);
    outputs(545) <= a and b;
    outputs(546) <= not (a xor b);
    outputs(547) <= b;
    outputs(548) <= not a;
    outputs(549) <= b and not a;
    outputs(550) <= a and b;
    outputs(551) <= not (a or b);
    outputs(552) <= a and b;
    outputs(553) <= a and b;
    outputs(554) <= not a;
    outputs(555) <= a;
    outputs(556) <= not a;
    outputs(557) <= b and not a;
    outputs(558) <= not b;
    outputs(559) <= a;
    outputs(560) <= a;
    outputs(561) <= b and not a;
    outputs(562) <= b and not a;
    outputs(563) <= a and b;
    outputs(564) <= a xor b;
    outputs(565) <= not b;
    outputs(566) <= a and b;
    outputs(567) <= not (a or b);
    outputs(568) <= not (a or b);
    outputs(569) <= b and not a;
    outputs(570) <= not (a or b);
    outputs(571) <= 1'b0;
    outputs(572) <= b and not a;
    outputs(573) <= not (a or b);
    outputs(574) <= not b;
    outputs(575) <= not (a or b);
    outputs(576) <= b and not a;
    outputs(577) <= a and not b;
    outputs(578) <= b and not a;
    outputs(579) <= b and not a;
    outputs(580) <= a and b;
    outputs(581) <= a and b;
    outputs(582) <= a and not b;
    outputs(583) <= a;
    outputs(584) <= b;
    outputs(585) <= b and not a;
    outputs(586) <= a;
    outputs(587) <= a and not b;
    outputs(588) <= b and not a;
    outputs(589) <= a and b;
    outputs(590) <= b and not a;
    outputs(591) <= a xor b;
    outputs(592) <= a and not b;
    outputs(593) <= b and not a;
    outputs(594) <= not b;
    outputs(595) <= a and not b;
    outputs(596) <= a and b;
    outputs(597) <= not (a xor b);
    outputs(598) <= a and b;
    outputs(599) <= not (a or b);
    outputs(600) <= a and b;
    outputs(601) <= not (a or b);
    outputs(602) <= a and b;
    outputs(603) <= not b;
    outputs(604) <= a and not b;
    outputs(605) <= not b;
    outputs(606) <= a and not b;
    outputs(607) <= b and not a;
    outputs(608) <= b and not a;
    outputs(609) <= a and not b;
    outputs(610) <= a;
    outputs(611) <= a and b;
    outputs(612) <= not (a or b);
    outputs(613) <= a and not b;
    outputs(614) <= not (a or b);
    outputs(615) <= a and b;
    outputs(616) <= b and not a;
    outputs(617) <= a and not b;
    outputs(618) <= a and b;
    outputs(619) <= not (a xor b);
    outputs(620) <= b and not a;
    outputs(621) <= a and b;
    outputs(622) <= not (a or b);
    outputs(623) <= not (a or b);
    outputs(624) <= a and not b;
    outputs(625) <= a and not b;
    outputs(626) <= b and not a;
    outputs(627) <= not a;
    outputs(628) <= a and b;
    outputs(629) <= a and b;
    outputs(630) <= a xor b;
    outputs(631) <= a and b;
    outputs(632) <= a;
    outputs(633) <= a and b;
    outputs(634) <= a;
    outputs(635) <= b and not a;
    outputs(636) <= not (a xor b);
    outputs(637) <= a and b;
    outputs(638) <= a;
    outputs(639) <= a and b;
    outputs(640) <= a and not b;
    outputs(641) <= not b;
    outputs(642) <= a and not b;
    outputs(643) <= not (a xor b);
    outputs(644) <= a;
    outputs(645) <= a and not b;
    outputs(646) <= not (a xor b);
    outputs(647) <= b and not a;
    outputs(648) <= a and not b;
    outputs(649) <= b and not a;
    outputs(650) <= a;
    outputs(651) <= not (a xor b);
    outputs(652) <= b;
    outputs(653) <= not (a xor b);
    outputs(654) <= a and not b;
    outputs(655) <= not (a or b);
    outputs(656) <= a xor b;
    outputs(657) <= a or b;
    outputs(658) <= a and not b;
    outputs(659) <= not (a or b);
    outputs(660) <= not (a or b);
    outputs(661) <= not (a or b);
    outputs(662) <= b;
    outputs(663) <= b;
    outputs(664) <= not a;
    outputs(665) <= not (a or b);
    outputs(666) <= a and b;
    outputs(667) <= a and b;
    outputs(668) <= not b;
    outputs(669) <= a xor b;
    outputs(670) <= not b or a;
    outputs(671) <= a and not b;
    outputs(672) <= b and not a;
    outputs(673) <= not a;
    outputs(674) <= a and b;
    outputs(675) <= a and b;
    outputs(676) <= not b;
    outputs(677) <= a and not b;
    outputs(678) <= not a;
    outputs(679) <= not b;
    outputs(680) <= not b;
    outputs(681) <= a xor b;
    outputs(682) <= not (a or b);
    outputs(683) <= b;
    outputs(684) <= a xor b;
    outputs(685) <= a and not b;
    outputs(686) <= not (a or b);
    outputs(687) <= a and b;
    outputs(688) <= a and b;
    outputs(689) <= not b;
    outputs(690) <= not (a or b);
    outputs(691) <= not (a xor b);
    outputs(692) <= not (a or b);
    outputs(693) <= a and not b;
    outputs(694) <= a and b;
    outputs(695) <= a and b;
    outputs(696) <= a and not b;
    outputs(697) <= not b;
    outputs(698) <= a and b;
    outputs(699) <= not a;
    outputs(700) <= not (a xor b);
    outputs(701) <= a and b;
    outputs(702) <= not a;
    outputs(703) <= a;
    outputs(704) <= b and not a;
    outputs(705) <= a and not b;
    outputs(706) <= not b;
    outputs(707) <= not (a or b);
    outputs(708) <= not b;
    outputs(709) <= b and not a;
    outputs(710) <= not (a or b);
    outputs(711) <= not (a or b);
    outputs(712) <= a and b;
    outputs(713) <= b and not a;
    outputs(714) <= b and not a;
    outputs(715) <= not b;
    outputs(716) <= 1'b0;
    outputs(717) <= b;
    outputs(718) <= 1'b0;
    outputs(719) <= not (a or b);
    outputs(720) <= b;
    outputs(721) <= not (a or b);
    outputs(722) <= b and not a;
    outputs(723) <= not b or a;
    outputs(724) <= b and not a;
    outputs(725) <= not b;
    outputs(726) <= not (a xor b);
    outputs(727) <= not a;
    outputs(728) <= b and not a;
    outputs(729) <= not (a xor b);
    outputs(730) <= not a;
    outputs(731) <= a and not b;
    outputs(732) <= b and not a;
    outputs(733) <= a and b;
    outputs(734) <= b;
    outputs(735) <= not (a xor b);
    outputs(736) <= a and not b;
    outputs(737) <= b and not a;
    outputs(738) <= b and not a;
    outputs(739) <= not (a or b);
    outputs(740) <= a and not b;
    outputs(741) <= not (a xor b);
    outputs(742) <= not a;
    outputs(743) <= a and not b;
    outputs(744) <= not b;
    outputs(745) <= a xor b;
    outputs(746) <= a and not b;
    outputs(747) <= a and not b;
    outputs(748) <= not (a and b);
    outputs(749) <= not a;
    outputs(750) <= not a or b;
    outputs(751) <= not (a xor b);
    outputs(752) <= not (a or b);
    outputs(753) <= b;
    outputs(754) <= a and b;
    outputs(755) <= a and not b;
    outputs(756) <= a xor b;
    outputs(757) <= not b;
    outputs(758) <= b;
    outputs(759) <= not (a or b);
    outputs(760) <= 1'b0;
    outputs(761) <= not (a xor b);
    outputs(762) <= a and not b;
    outputs(763) <= not (a xor b);
    outputs(764) <= not (a or b);
    outputs(765) <= b and not a;
    outputs(766) <= a xor b;
    outputs(767) <= a and not b;
    outputs(768) <= a and not b;
    outputs(769) <= a and not b;
    outputs(770) <= a;
    outputs(771) <= a and b;
    outputs(772) <= a;
    outputs(773) <= b and not a;
    outputs(774) <= a and not b;
    outputs(775) <= not (a or b);
    outputs(776) <= not (a xor b);
    outputs(777) <= b and not a;
    outputs(778) <= not b;
    outputs(779) <= not (a or b);
    outputs(780) <= b;
    outputs(781) <= b and not a;
    outputs(782) <= b;
    outputs(783) <= a and b;
    outputs(784) <= not (a xor b);
    outputs(785) <= not a;
    outputs(786) <= b;
    outputs(787) <= a and b;
    outputs(788) <= not (a xor b);
    outputs(789) <= not (a or b);
    outputs(790) <= not (a or b);
    outputs(791) <= b and not a;
    outputs(792) <= b and not a;
    outputs(793) <= b and not a;
    outputs(794) <= a and not b;
    outputs(795) <= a and b;
    outputs(796) <= b;
    outputs(797) <= a and b;
    outputs(798) <= a and not b;
    outputs(799) <= b;
    outputs(800) <= not a;
    outputs(801) <= b and not a;
    outputs(802) <= a and not b;
    outputs(803) <= not (a xor b);
    outputs(804) <= not a;
    outputs(805) <= a and b;
    outputs(806) <= not (a or b);
    outputs(807) <= not b;
    outputs(808) <= a xor b;
    outputs(809) <= not (a or b);
    outputs(810) <= not (a xor b);
    outputs(811) <= b and not a;
    outputs(812) <= not a;
    outputs(813) <= a;
    outputs(814) <= b and not a;
    outputs(815) <= not (a or b);
    outputs(816) <= a and b;
    outputs(817) <= a xor b;
    outputs(818) <= a and not b;
    outputs(819) <= a;
    outputs(820) <= b;
    outputs(821) <= a;
    outputs(822) <= a and not b;
    outputs(823) <= a xor b;
    outputs(824) <= b and not a;
    outputs(825) <= a;
    outputs(826) <= a and not b;
    outputs(827) <= a and b;
    outputs(828) <= not (a or b);
    outputs(829) <= b;
    outputs(830) <= b and not a;
    outputs(831) <= not (a or b);
    outputs(832) <= not a;
    outputs(833) <= a xor b;
    outputs(834) <= a xor b;
    outputs(835) <= not (a xor b);
    outputs(836) <= a and b;
    outputs(837) <= a;
    outputs(838) <= a xor b;
    outputs(839) <= b;
    outputs(840) <= not (a or b);
    outputs(841) <= b;
    outputs(842) <= a and not b;
    outputs(843) <= not b;
    outputs(844) <= not b;
    outputs(845) <= a and b;
    outputs(846) <= a and not b;
    outputs(847) <= a and not b;
    outputs(848) <= b and not a;
    outputs(849) <= b and not a;
    outputs(850) <= a and not b;
    outputs(851) <= a and not b;
    outputs(852) <= not (a xor b);
    outputs(853) <= b and not a;
    outputs(854) <= b and not a;
    outputs(855) <= a;
    outputs(856) <= a and not b;
    outputs(857) <= a and b;
    outputs(858) <= b and not a;
    outputs(859) <= not (a or b);
    outputs(860) <= not a;
    outputs(861) <= a xor b;
    outputs(862) <= a and b;
    outputs(863) <= not (a or b);
    outputs(864) <= b;
    outputs(865) <= a xor b;
    outputs(866) <= b and not a;
    outputs(867) <= b and not a;
    outputs(868) <= not (a xor b);
    outputs(869) <= a;
    outputs(870) <= not b;
    outputs(871) <= a xor b;
    outputs(872) <= b and not a;
    outputs(873) <= b and not a;
    outputs(874) <= not b;
    outputs(875) <= not (a or b);
    outputs(876) <= not (a or b);
    outputs(877) <= not (a or b);
    outputs(878) <= a;
    outputs(879) <= a;
    outputs(880) <= a;
    outputs(881) <= a and not b;
    outputs(882) <= b;
    outputs(883) <= a and not b;
    outputs(884) <= not a;
    outputs(885) <= not (a or b);
    outputs(886) <= a or b;
    outputs(887) <= not (a or b);
    outputs(888) <= not b;
    outputs(889) <= not (a and b);
    outputs(890) <= b and not a;
    outputs(891) <= a;
    outputs(892) <= not (a or b);
    outputs(893) <= not (a or b);
    outputs(894) <= b;
    outputs(895) <= not (a or b);
    outputs(896) <= b;
    outputs(897) <= a and b;
    outputs(898) <= b and not a;
    outputs(899) <= not b;
    outputs(900) <= a and b;
    outputs(901) <= not (a or b);
    outputs(902) <= a and b;
    outputs(903) <= b and not a;
    outputs(904) <= a;
    outputs(905) <= a;
    outputs(906) <= a and b;
    outputs(907) <= not (a or b);
    outputs(908) <= a xor b;
    outputs(909) <= a and b;
    outputs(910) <= a and b;
    outputs(911) <= a and not b;
    outputs(912) <= not a or b;
    outputs(913) <= a and not b;
    outputs(914) <= b;
    outputs(915) <= not (a or b);
    outputs(916) <= a and b;
    outputs(917) <= a;
    outputs(918) <= b and not a;
    outputs(919) <= b and not a;
    outputs(920) <= not b;
    outputs(921) <= a and not b;
    outputs(922) <= a and not b;
    outputs(923) <= a and not b;
    outputs(924) <= a;
    outputs(925) <= not (a xor b);
    outputs(926) <= not a;
    outputs(927) <= a and not b;
    outputs(928) <= a and b;
    outputs(929) <= a and b;
    outputs(930) <= b;
    outputs(931) <= not (a xor b);
    outputs(932) <= b and not a;
    outputs(933) <= a and b;
    outputs(934) <= not (a or b);
    outputs(935) <= a or b;
    outputs(936) <= a and b;
    outputs(937) <= a and b;
    outputs(938) <= a and b;
    outputs(939) <= not a;
    outputs(940) <= a and b;
    outputs(941) <= b and not a;
    outputs(942) <= a and not b;
    outputs(943) <= b;
    outputs(944) <= b;
    outputs(945) <= a and b;
    outputs(946) <= a and b;
    outputs(947) <= not (a or b);
    outputs(948) <= not (a or b);
    outputs(949) <= a and not b;
    outputs(950) <= not a;
    outputs(951) <= b and not a;
    outputs(952) <= not (a xor b);
    outputs(953) <= a xor b;
    outputs(954) <= not (a xor b);
    outputs(955) <= not (a or b);
    outputs(956) <= a;
    outputs(957) <= not b;
    outputs(958) <= a and b;
    outputs(959) <= a and b;
    outputs(960) <= b and not a;
    outputs(961) <= a xor b;
    outputs(962) <= b;
    outputs(963) <= 1'b0;
    outputs(964) <= a and b;
    outputs(965) <= not (a or b);
    outputs(966) <= b and not a;
    outputs(967) <= a and b;
    outputs(968) <= b and not a;
    outputs(969) <= not (a xor b);
    outputs(970) <= b and not a;
    outputs(971) <= not a;
    outputs(972) <= a and not b;
    outputs(973) <= a;
    outputs(974) <= b and not a;
    outputs(975) <= a xor b;
    outputs(976) <= a and b;
    outputs(977) <= b and not a;
    outputs(978) <= a;
    outputs(979) <= a xor b;
    outputs(980) <= not b;
    outputs(981) <= a and b;
    outputs(982) <= a and b;
    outputs(983) <= not a;
    outputs(984) <= not a;
    outputs(985) <= a and not b;
    outputs(986) <= a and not b;
    outputs(987) <= b and not a;
    outputs(988) <= a xor b;
    outputs(989) <= a and b;
    outputs(990) <= not b;
    outputs(991) <= b and not a;
    outputs(992) <= a xor b;
    outputs(993) <= b and not a;
    outputs(994) <= not (a or b);
    outputs(995) <= not (a or b);
    outputs(996) <= a and not b;
    outputs(997) <= a xor b;
    outputs(998) <= a;
    outputs(999) <= not b;
    outputs(1000) <= not (a xor b);
    outputs(1001) <= a and b;
    outputs(1002) <= b;
    outputs(1003) <= not (a or b);
    outputs(1004) <= a and b;
    outputs(1005) <= not (a xor b);
    outputs(1006) <= not b;
    outputs(1007) <= a and not b;
    outputs(1008) <= not (a or b);
    outputs(1009) <= b and not a;
    outputs(1010) <= not b;
    outputs(1011) <= b;
    outputs(1012) <= a and b;
    outputs(1013) <= b and not a;
    outputs(1014) <= b and not a;
    outputs(1015) <= not (a or b);
    outputs(1016) <= a and not b;
    outputs(1017) <= not (a xor b);
    outputs(1018) <= not (a or b);
    outputs(1019) <= a and b;
    outputs(1020) <= b and not a;
    outputs(1021) <= a;
    outputs(1022) <= b and not a;
    outputs(1023) <= a;
    outputs(1024) <= not (a xor b);
    outputs(1025) <= a and b;
    outputs(1026) <= not (a xor b);
    outputs(1027) <= b;
    outputs(1028) <= not b;
    outputs(1029) <= a and b;
    outputs(1030) <= b;
    outputs(1031) <= not (a xor b);
    outputs(1032) <= a;
    outputs(1033) <= b;
    outputs(1034) <= a or b;
    outputs(1035) <= a and b;
    outputs(1036) <= b;
    outputs(1037) <= not a;
    outputs(1038) <= a;
    outputs(1039) <= b;
    outputs(1040) <= a or b;
    outputs(1041) <= not (a or b);
    outputs(1042) <= a or b;
    outputs(1043) <= a and not b;
    outputs(1044) <= a;
    outputs(1045) <= not b or a;
    outputs(1046) <= not a;
    outputs(1047) <= not a;
    outputs(1048) <= a and b;
    outputs(1049) <= b;
    outputs(1050) <= a and not b;
    outputs(1051) <= not (a and b);
    outputs(1052) <= a;
    outputs(1053) <= not (a and b);
    outputs(1054) <= a and b;
    outputs(1055) <= not (a and b);
    outputs(1056) <= a or b;
    outputs(1057) <= not a;
    outputs(1058) <= not a or b;
    outputs(1059) <= a xor b;
    outputs(1060) <= not a or b;
    outputs(1061) <= b;
    outputs(1062) <= b;
    outputs(1063) <= b;
    outputs(1064) <= not b or a;
    outputs(1065) <= a;
    outputs(1066) <= not (a and b);
    outputs(1067) <= not (a xor b);
    outputs(1068) <= a xor b;
    outputs(1069) <= not a or b;
    outputs(1070) <= b;
    outputs(1071) <= not (a or b);
    outputs(1072) <= not b;
    outputs(1073) <= a or b;
    outputs(1074) <= not b;
    outputs(1075) <= a;
    outputs(1076) <= not b;
    outputs(1077) <= a xor b;
    outputs(1078) <= a or b;
    outputs(1079) <= not b;
    outputs(1080) <= a;
    outputs(1081) <= b;
    outputs(1082) <= b and not a;
    outputs(1083) <= a;
    outputs(1084) <= not (a xor b);
    outputs(1085) <= a;
    outputs(1086) <= a and b;
    outputs(1087) <= not b;
    outputs(1088) <= not (a and b);
    outputs(1089) <= not a;
    outputs(1090) <= not (a or b);
    outputs(1091) <= not (a and b);
    outputs(1092) <= not a;
    outputs(1093) <= a and not b;
    outputs(1094) <= a xor b;
    outputs(1095) <= not b;
    outputs(1096) <= not (a and b);
    outputs(1097) <= b;
    outputs(1098) <= not b;
    outputs(1099) <= a and not b;
    outputs(1100) <= not a or b;
    outputs(1101) <= b;
    outputs(1102) <= not (a and b);
    outputs(1103) <= not a or b;
    outputs(1104) <= a;
    outputs(1105) <= a and b;
    outputs(1106) <= not (a or b);
    outputs(1107) <= not a;
    outputs(1108) <= not (a or b);
    outputs(1109) <= a and not b;
    outputs(1110) <= not a or b;
    outputs(1111) <= a or b;
    outputs(1112) <= b;
    outputs(1113) <= not a or b;
    outputs(1114) <= not (a and b);
    outputs(1115) <= not a;
    outputs(1116) <= a;
    outputs(1117) <= a or b;
    outputs(1118) <= a and not b;
    outputs(1119) <= b;
    outputs(1120) <= b;
    outputs(1121) <= a;
    outputs(1122) <= a;
    outputs(1123) <= a xor b;
    outputs(1124) <= not a;
    outputs(1125) <= a and b;
    outputs(1126) <= a and b;
    outputs(1127) <= b;
    outputs(1128) <= a and not b;
    outputs(1129) <= a or b;
    outputs(1130) <= not a;
    outputs(1131) <= not (a and b);
    outputs(1132) <= b;
    outputs(1133) <= a;
    outputs(1134) <= a xor b;
    outputs(1135) <= a xor b;
    outputs(1136) <= b;
    outputs(1137) <= b;
    outputs(1138) <= not b or a;
    outputs(1139) <= not (a and b);
    outputs(1140) <= not (a xor b);
    outputs(1141) <= not a;
    outputs(1142) <= not b or a;
    outputs(1143) <= b;
    outputs(1144) <= not a;
    outputs(1145) <= not b;
    outputs(1146) <= a and not b;
    outputs(1147) <= b;
    outputs(1148) <= not (a and b);
    outputs(1149) <= b;
    outputs(1150) <= not (a and b);
    outputs(1151) <= a;
    outputs(1152) <= not (a or b);
    outputs(1153) <= not (a or b);
    outputs(1154) <= a;
    outputs(1155) <= not b;
    outputs(1156) <= a and not b;
    outputs(1157) <= b;
    outputs(1158) <= b;
    outputs(1159) <= a xor b;
    outputs(1160) <= b;
    outputs(1161) <= not (a or b);
    outputs(1162) <= not (a xor b);
    outputs(1163) <= a;
    outputs(1164) <= not (a and b);
    outputs(1165) <= b;
    outputs(1166) <= not (a or b);
    outputs(1167) <= b;
    outputs(1168) <= a and b;
    outputs(1169) <= b;
    outputs(1170) <= b;
    outputs(1171) <= a and not b;
    outputs(1172) <= not (a xor b);
    outputs(1173) <= not (a and b);
    outputs(1174) <= not (a xor b);
    outputs(1175) <= a;
    outputs(1176) <= not (a xor b);
    outputs(1177) <= a xor b;
    outputs(1178) <= not (a or b);
    outputs(1179) <= not a;
    outputs(1180) <= not (a xor b);
    outputs(1181) <= not b;
    outputs(1182) <= not a;
    outputs(1183) <= b;
    outputs(1184) <= not a or b;
    outputs(1185) <= a and b;
    outputs(1186) <= b and not a;
    outputs(1187) <= not b;
    outputs(1188) <= not b or a;
    outputs(1189) <= not b;
    outputs(1190) <= not (a xor b);
    outputs(1191) <= not a;
    outputs(1192) <= a xor b;
    outputs(1193) <= not a;
    outputs(1194) <= not b;
    outputs(1195) <= b;
    outputs(1196) <= a xor b;
    outputs(1197) <= a or b;
    outputs(1198) <= not b;
    outputs(1199) <= b;
    outputs(1200) <= not b;
    outputs(1201) <= not b;
    outputs(1202) <= a and not b;
    outputs(1203) <= a;
    outputs(1204) <= a;
    outputs(1205) <= not b or a;
    outputs(1206) <= b;
    outputs(1207) <= not a or b;
    outputs(1208) <= not a;
    outputs(1209) <= a;
    outputs(1210) <= not b;
    outputs(1211) <= not b;
    outputs(1212) <= not b or a;
    outputs(1213) <= a and not b;
    outputs(1214) <= not (a xor b);
    outputs(1215) <= not a;
    outputs(1216) <= not a or b;
    outputs(1217) <= not b;
    outputs(1218) <= not b or a;
    outputs(1219) <= a or b;
    outputs(1220) <= not (a and b);
    outputs(1221) <= a xor b;
    outputs(1222) <= not a or b;
    outputs(1223) <= not b or a;
    outputs(1224) <= not (a or b);
    outputs(1225) <= not b;
    outputs(1226) <= not b;
    outputs(1227) <= b;
    outputs(1228) <= a or b;
    outputs(1229) <= a;
    outputs(1230) <= a xor b;
    outputs(1231) <= a;
    outputs(1232) <= not (a and b);
    outputs(1233) <= not (a or b);
    outputs(1234) <= not b or a;
    outputs(1235) <= a xor b;
    outputs(1236) <= a or b;
    outputs(1237) <= not b;
    outputs(1238) <= not (a or b);
    outputs(1239) <= not (a xor b);
    outputs(1240) <= not a;
    outputs(1241) <= not (a xor b);
    outputs(1242) <= a;
    outputs(1243) <= not b or a;
    outputs(1244) <= not b;
    outputs(1245) <= not (a or b);
    outputs(1246) <= not b;
    outputs(1247) <= a xor b;
    outputs(1248) <= not a or b;
    outputs(1249) <= a;
    outputs(1250) <= b;
    outputs(1251) <= a xor b;
    outputs(1252) <= b and not a;
    outputs(1253) <= not (a or b);
    outputs(1254) <= b;
    outputs(1255) <= not a or b;
    outputs(1256) <= a and b;
    outputs(1257) <= not a;
    outputs(1258) <= a xor b;
    outputs(1259) <= not b or a;
    outputs(1260) <= not (a xor b);
    outputs(1261) <= a;
    outputs(1262) <= b;
    outputs(1263) <= not (a xor b);
    outputs(1264) <= not a or b;
    outputs(1265) <= a and b;
    outputs(1266) <= not a or b;
    outputs(1267) <= not (a xor b);
    outputs(1268) <= a and not b;
    outputs(1269) <= not a;
    outputs(1270) <= not b;
    outputs(1271) <= a or b;
    outputs(1272) <= not (a or b);
    outputs(1273) <= not b;
    outputs(1274) <= b;
    outputs(1275) <= a;
    outputs(1276) <= b;
    outputs(1277) <= not (a or b);
    outputs(1278) <= b and not a;
    outputs(1279) <= not b;
    outputs(1280) <= not (a or b);
    outputs(1281) <= not a or b;
    outputs(1282) <= not b or a;
    outputs(1283) <= a;
    outputs(1284) <= b;
    outputs(1285) <= not b;
    outputs(1286) <= not a;
    outputs(1287) <= not b;
    outputs(1288) <= not a;
    outputs(1289) <= not a;
    outputs(1290) <= not (a xor b);
    outputs(1291) <= not b;
    outputs(1292) <= not a;
    outputs(1293) <= a and b;
    outputs(1294) <= b;
    outputs(1295) <= not (a xor b);
    outputs(1296) <= a;
    outputs(1297) <= not a;
    outputs(1298) <= not (a xor b);
    outputs(1299) <= a;
    outputs(1300) <= not b;
    outputs(1301) <= b;
    outputs(1302) <= a or b;
    outputs(1303) <= not a;
    outputs(1304) <= b;
    outputs(1305) <= b;
    outputs(1306) <= not a;
    outputs(1307) <= not a;
    outputs(1308) <= not a;
    outputs(1309) <= b and not a;
    outputs(1310) <= a or b;
    outputs(1311) <= b;
    outputs(1312) <= not b;
    outputs(1313) <= b;
    outputs(1314) <= b and not a;
    outputs(1315) <= not b;
    outputs(1316) <= not a;
    outputs(1317) <= not b;
    outputs(1318) <= a xor b;
    outputs(1319) <= b;
    outputs(1320) <= a and not b;
    outputs(1321) <= a xor b;
    outputs(1322) <= b;
    outputs(1323) <= not (a and b);
    outputs(1324) <= a;
    outputs(1325) <= a;
    outputs(1326) <= a;
    outputs(1327) <= a and not b;
    outputs(1328) <= not a;
    outputs(1329) <= not (a xor b);
    outputs(1330) <= not (a xor b);
    outputs(1331) <= not a;
    outputs(1332) <= not (a and b);
    outputs(1333) <= not b;
    outputs(1334) <= not b;
    outputs(1335) <= a xor b;
    outputs(1336) <= not b;
    outputs(1337) <= b;
    outputs(1338) <= not (a and b);
    outputs(1339) <= not (a or b);
    outputs(1340) <= a or b;
    outputs(1341) <= a or b;
    outputs(1342) <= a;
    outputs(1343) <= not (a xor b);
    outputs(1344) <= a and b;
    outputs(1345) <= not b or a;
    outputs(1346) <= a or b;
    outputs(1347) <= not b;
    outputs(1348) <= not (a xor b);
    outputs(1349) <= b;
    outputs(1350) <= not a or b;
    outputs(1351) <= a;
    outputs(1352) <= a or b;
    outputs(1353) <= a and b;
    outputs(1354) <= not (a or b);
    outputs(1355) <= a;
    outputs(1356) <= not b;
    outputs(1357) <= a;
    outputs(1358) <= b;
    outputs(1359) <= b;
    outputs(1360) <= a or b;
    outputs(1361) <= a and b;
    outputs(1362) <= not b;
    outputs(1363) <= not a;
    outputs(1364) <= not b;
    outputs(1365) <= not b;
    outputs(1366) <= not b or a;
    outputs(1367) <= b;
    outputs(1368) <= not a;
    outputs(1369) <= not b;
    outputs(1370) <= not (a and b);
    outputs(1371) <= a;
    outputs(1372) <= a and not b;
    outputs(1373) <= not a or b;
    outputs(1374) <= a;
    outputs(1375) <= not a;
    outputs(1376) <= not a or b;
    outputs(1377) <= a xor b;
    outputs(1378) <= not b or a;
    outputs(1379) <= b and not a;
    outputs(1380) <= a or b;
    outputs(1381) <= b;
    outputs(1382) <= not a or b;
    outputs(1383) <= not a or b;
    outputs(1384) <= a xor b;
    outputs(1385) <= b and not a;
    outputs(1386) <= a or b;
    outputs(1387) <= a and b;
    outputs(1388) <= not (a xor b);
    outputs(1389) <= a;
    outputs(1390) <= not b;
    outputs(1391) <= a and b;
    outputs(1392) <= not a;
    outputs(1393) <= a xor b;
    outputs(1394) <= not (a xor b);
    outputs(1395) <= a;
    outputs(1396) <= not a;
    outputs(1397) <= not (a xor b);
    outputs(1398) <= a and b;
    outputs(1399) <= not b;
    outputs(1400) <= a;
    outputs(1401) <= not (a xor b);
    outputs(1402) <= not b;
    outputs(1403) <= a or b;
    outputs(1404) <= not a;
    outputs(1405) <= not a;
    outputs(1406) <= a and b;
    outputs(1407) <= a;
    outputs(1408) <= b;
    outputs(1409) <= not a;
    outputs(1410) <= not b;
    outputs(1411) <= not b;
    outputs(1412) <= not b;
    outputs(1413) <= b and not a;
    outputs(1414) <= not (a and b);
    outputs(1415) <= not (a xor b);
    outputs(1416) <= not (a or b);
    outputs(1417) <= not a;
    outputs(1418) <= a and not b;
    outputs(1419) <= not b;
    outputs(1420) <= b and not a;
    outputs(1421) <= a;
    outputs(1422) <= a or b;
    outputs(1423) <= a;
    outputs(1424) <= not a;
    outputs(1425) <= b and not a;
    outputs(1426) <= not b or a;
    outputs(1427) <= a;
    outputs(1428) <= not b;
    outputs(1429) <= not (a xor b);
    outputs(1430) <= b;
    outputs(1431) <= not b;
    outputs(1432) <= not a;
    outputs(1433) <= a and not b;
    outputs(1434) <= a;
    outputs(1435) <= not (a or b);
    outputs(1436) <= not b;
    outputs(1437) <= a;
    outputs(1438) <= not a or b;
    outputs(1439) <= not (a or b);
    outputs(1440) <= b and not a;
    outputs(1441) <= b;
    outputs(1442) <= a and not b;
    outputs(1443) <= a xor b;
    outputs(1444) <= not b;
    outputs(1445) <= not b or a;
    outputs(1446) <= not a;
    outputs(1447) <= b;
    outputs(1448) <= a;
    outputs(1449) <= not (a or b);
    outputs(1450) <= not (a xor b);
    outputs(1451) <= b;
    outputs(1452) <= not b;
    outputs(1453) <= not b;
    outputs(1454) <= b;
    outputs(1455) <= not a or b;
    outputs(1456) <= not a or b;
    outputs(1457) <= b;
    outputs(1458) <= not (a xor b);
    outputs(1459) <= b;
    outputs(1460) <= not b;
    outputs(1461) <= not a;
    outputs(1462) <= a;
    outputs(1463) <= a;
    outputs(1464) <= a and b;
    outputs(1465) <= not a or b;
    outputs(1466) <= b and not a;
    outputs(1467) <= a;
    outputs(1468) <= not (a and b);
    outputs(1469) <= not b;
    outputs(1470) <= a;
    outputs(1471) <= a;
    outputs(1472) <= a xor b;
    outputs(1473) <= a and b;
    outputs(1474) <= a and b;
    outputs(1475) <= a;
    outputs(1476) <= not b;
    outputs(1477) <= a and not b;
    outputs(1478) <= not a;
    outputs(1479) <= not a;
    outputs(1480) <= not a;
    outputs(1481) <= not (a xor b);
    outputs(1482) <= not b or a;
    outputs(1483) <= not a;
    outputs(1484) <= not (a and b);
    outputs(1485) <= not b or a;
    outputs(1486) <= b and not a;
    outputs(1487) <= not b or a;
    outputs(1488) <= not a;
    outputs(1489) <= a xor b;
    outputs(1490) <= b;
    outputs(1491) <= not b or a;
    outputs(1492) <= not a;
    outputs(1493) <= not (a or b);
    outputs(1494) <= a and not b;
    outputs(1495) <= a and b;
    outputs(1496) <= a xor b;
    outputs(1497) <= not a;
    outputs(1498) <= b and not a;
    outputs(1499) <= not a or b;
    outputs(1500) <= not a;
    outputs(1501) <= a xor b;
    outputs(1502) <= b;
    outputs(1503) <= not b;
    outputs(1504) <= not a;
    outputs(1505) <= not (a or b);
    outputs(1506) <= a and b;
    outputs(1507) <= not b;
    outputs(1508) <= b;
    outputs(1509) <= a and not b;
    outputs(1510) <= not a;
    outputs(1511) <= a;
    outputs(1512) <= a and b;
    outputs(1513) <= b and not a;
    outputs(1514) <= a and b;
    outputs(1515) <= b;
    outputs(1516) <= b and not a;
    outputs(1517) <= b;
    outputs(1518) <= not (a and b);
    outputs(1519) <= a;
    outputs(1520) <= not (a xor b);
    outputs(1521) <= b;
    outputs(1522) <= not a or b;
    outputs(1523) <= not (a xor b);
    outputs(1524) <= not b;
    outputs(1525) <= not b;
    outputs(1526) <= not a;
    outputs(1527) <= not a;
    outputs(1528) <= not a;
    outputs(1529) <= not a;
    outputs(1530) <= a;
    outputs(1531) <= a;
    outputs(1532) <= not a;
    outputs(1533) <= a and not b;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= b;
    outputs(1536) <= not (a xor b);
    outputs(1537) <= not (a xor b);
    outputs(1538) <= not b or a;
    outputs(1539) <= a;
    outputs(1540) <= a and b;
    outputs(1541) <= b;
    outputs(1542) <= not b;
    outputs(1543) <= b;
    outputs(1544) <= b;
    outputs(1545) <= a;
    outputs(1546) <= not (a and b);
    outputs(1547) <= not a or b;
    outputs(1548) <= a;
    outputs(1549) <= a xor b;
    outputs(1550) <= not a or b;
    outputs(1551) <= a xor b;
    outputs(1552) <= b;
    outputs(1553) <= b;
    outputs(1554) <= a xor b;
    outputs(1555) <= not (a or b);
    outputs(1556) <= a;
    outputs(1557) <= not (a xor b);
    outputs(1558) <= a;
    outputs(1559) <= not a;
    outputs(1560) <= not a;
    outputs(1561) <= not a;
    outputs(1562) <= b;
    outputs(1563) <= not (a xor b);
    outputs(1564) <= a or b;
    outputs(1565) <= not b;
    outputs(1566) <= not b or a;
    outputs(1567) <= b;
    outputs(1568) <= b and not a;
    outputs(1569) <= not (a or b);
    outputs(1570) <= not b;
    outputs(1571) <= a;
    outputs(1572) <= a and not b;
    outputs(1573) <= not a;
    outputs(1574) <= not a or b;
    outputs(1575) <= a and b;
    outputs(1576) <= not a;
    outputs(1577) <= b;
    outputs(1578) <= a and b;
    outputs(1579) <= not a;
    outputs(1580) <= not b;
    outputs(1581) <= not a;
    outputs(1582) <= a;
    outputs(1583) <= not (a xor b);
    outputs(1584) <= not a;
    outputs(1585) <= a;
    outputs(1586) <= not a;
    outputs(1587) <= not a;
    outputs(1588) <= not a;
    outputs(1589) <= not b;
    outputs(1590) <= not b or a;
    outputs(1591) <= not a or b;
    outputs(1592) <= not (a xor b);
    outputs(1593) <= not (a xor b);
    outputs(1594) <= a and not b;
    outputs(1595) <= not (a and b);
    outputs(1596) <= not a or b;
    outputs(1597) <= b and not a;
    outputs(1598) <= a and not b;
    outputs(1599) <= 1'b0;
    outputs(1600) <= b and not a;
    outputs(1601) <= not b;
    outputs(1602) <= not b;
    outputs(1603) <= not b;
    outputs(1604) <= not b;
    outputs(1605) <= not a;
    outputs(1606) <= a;
    outputs(1607) <= a;
    outputs(1608) <= a or b;
    outputs(1609) <= a or b;
    outputs(1610) <= not (a xor b);
    outputs(1611) <= not (a or b);
    outputs(1612) <= not b;
    outputs(1613) <= not a;
    outputs(1614) <= a and not b;
    outputs(1615) <= not a;
    outputs(1616) <= not (a or b);
    outputs(1617) <= not b;
    outputs(1618) <= a and b;
    outputs(1619) <= a and b;
    outputs(1620) <= a xor b;
    outputs(1621) <= a xor b;
    outputs(1622) <= b;
    outputs(1623) <= a and b;
    outputs(1624) <= b;
    outputs(1625) <= not (a xor b);
    outputs(1626) <= a xor b;
    outputs(1627) <= a and b;
    outputs(1628) <= b and not a;
    outputs(1629) <= a;
    outputs(1630) <= a;
    outputs(1631) <= not (a or b);
    outputs(1632) <= b;
    outputs(1633) <= a and b;
    outputs(1634) <= b and not a;
    outputs(1635) <= b and not a;
    outputs(1636) <= not a or b;
    outputs(1637) <= a xor b;
    outputs(1638) <= a;
    outputs(1639) <= a;
    outputs(1640) <= not (a or b);
    outputs(1641) <= not (a xor b);
    outputs(1642) <= b and not a;
    outputs(1643) <= a;
    outputs(1644) <= not a or b;
    outputs(1645) <= b;
    outputs(1646) <= not b;
    outputs(1647) <= b;
    outputs(1648) <= not b;
    outputs(1649) <= not (a or b);
    outputs(1650) <= a;
    outputs(1651) <= a and not b;
    outputs(1652) <= not (a xor b);
    outputs(1653) <= b;
    outputs(1654) <= not a or b;
    outputs(1655) <= a and b;
    outputs(1656) <= not b;
    outputs(1657) <= b;
    outputs(1658) <= b;
    outputs(1659) <= a xor b;
    outputs(1660) <= not b;
    outputs(1661) <= a xor b;
    outputs(1662) <= not (a or b);
    outputs(1663) <= b and not a;
    outputs(1664) <= not (a xor b);
    outputs(1665) <= not (a xor b);
    outputs(1666) <= not a;
    outputs(1667) <= not (a and b);
    outputs(1668) <= not a;
    outputs(1669) <= not a;
    outputs(1670) <= not b;
    outputs(1671) <= a and b;
    outputs(1672) <= not a;
    outputs(1673) <= a;
    outputs(1674) <= a or b;
    outputs(1675) <= a or b;
    outputs(1676) <= b and not a;
    outputs(1677) <= b;
    outputs(1678) <= not b;
    outputs(1679) <= not b or a;
    outputs(1680) <= not a or b;
    outputs(1681) <= a;
    outputs(1682) <= not (a xor b);
    outputs(1683) <= not b;
    outputs(1684) <= not b;
    outputs(1685) <= a;
    outputs(1686) <= a and b;
    outputs(1687) <= a;
    outputs(1688) <= not b;
    outputs(1689) <= not b;
    outputs(1690) <= not (a xor b);
    outputs(1691) <= not (a xor b);
    outputs(1692) <= a xor b;
    outputs(1693) <= not b;
    outputs(1694) <= not (a or b);
    outputs(1695) <= not (a and b);
    outputs(1696) <= a xor b;
    outputs(1697) <= a or b;
    outputs(1698) <= b;
    outputs(1699) <= a or b;
    outputs(1700) <= not b;
    outputs(1701) <= b and not a;
    outputs(1702) <= not (a xor b);
    outputs(1703) <= not (a or b);
    outputs(1704) <= a;
    outputs(1705) <= not (a and b);
    outputs(1706) <= not (a or b);
    outputs(1707) <= not a;
    outputs(1708) <= not a;
    outputs(1709) <= not a or b;
    outputs(1710) <= a xor b;
    outputs(1711) <= b and not a;
    outputs(1712) <= a xor b;
    outputs(1713) <= a and not b;
    outputs(1714) <= not b;
    outputs(1715) <= a xor b;
    outputs(1716) <= not b or a;
    outputs(1717) <= not (a and b);
    outputs(1718) <= not a;
    outputs(1719) <= not (a or b);
    outputs(1720) <= a;
    outputs(1721) <= b;
    outputs(1722) <= a;
    outputs(1723) <= not b;
    outputs(1724) <= a and not b;
    outputs(1725) <= not b;
    outputs(1726) <= a or b;
    outputs(1727) <= a and b;
    outputs(1728) <= a and not b;
    outputs(1729) <= b;
    outputs(1730) <= not b;
    outputs(1731) <= b and not a;
    outputs(1732) <= not a or b;
    outputs(1733) <= b;
    outputs(1734) <= not b;
    outputs(1735) <= not b;
    outputs(1736) <= b;
    outputs(1737) <= not b;
    outputs(1738) <= not b;
    outputs(1739) <= a;
    outputs(1740) <= b and not a;
    outputs(1741) <= a xor b;
    outputs(1742) <= not (a xor b);
    outputs(1743) <= not (a or b);
    outputs(1744) <= not a;
    outputs(1745) <= not b or a;
    outputs(1746) <= a xor b;
    outputs(1747) <= not b;
    outputs(1748) <= not b;
    outputs(1749) <= a or b;
    outputs(1750) <= not b;
    outputs(1751) <= not b;
    outputs(1752) <= a;
    outputs(1753) <= b and not a;
    outputs(1754) <= not (a xor b);
    outputs(1755) <= a;
    outputs(1756) <= not (a or b);
    outputs(1757) <= a xor b;
    outputs(1758) <= not (a or b);
    outputs(1759) <= a and not b;
    outputs(1760) <= not a or b;
    outputs(1761) <= b;
    outputs(1762) <= not b;
    outputs(1763) <= a or b;
    outputs(1764) <= not b;
    outputs(1765) <= not (a or b);
    outputs(1766) <= a;
    outputs(1767) <= not (a and b);
    outputs(1768) <= not b or a;
    outputs(1769) <= a and not b;
    outputs(1770) <= a or b;
    outputs(1771) <= a;
    outputs(1772) <= not (a xor b);
    outputs(1773) <= not b or a;
    outputs(1774) <= not b;
    outputs(1775) <= b and not a;
    outputs(1776) <= a and not b;
    outputs(1777) <= not b;
    outputs(1778) <= a xor b;
    outputs(1779) <= not a;
    outputs(1780) <= a;
    outputs(1781) <= not a;
    outputs(1782) <= b and not a;
    outputs(1783) <= a xor b;
    outputs(1784) <= b and not a;
    outputs(1785) <= not a or b;
    outputs(1786) <= not b;
    outputs(1787) <= a or b;
    outputs(1788) <= not a;
    outputs(1789) <= not (a xor b);
    outputs(1790) <= a and not b;
    outputs(1791) <= not (a or b);
    outputs(1792) <= b;
    outputs(1793) <= b and not a;
    outputs(1794) <= a;
    outputs(1795) <= a and b;
    outputs(1796) <= not b;
    outputs(1797) <= a and not b;
    outputs(1798) <= not b;
    outputs(1799) <= a and b;
    outputs(1800) <= not b;
    outputs(1801) <= not a;
    outputs(1802) <= not (a xor b);
    outputs(1803) <= b;
    outputs(1804) <= b and not a;
    outputs(1805) <= a;
    outputs(1806) <= not b;
    outputs(1807) <= not a;
    outputs(1808) <= not a;
    outputs(1809) <= a or b;
    outputs(1810) <= a or b;
    outputs(1811) <= not a or b;
    outputs(1812) <= not b;
    outputs(1813) <= not a;
    outputs(1814) <= not (a or b);
    outputs(1815) <= not (a or b);
    outputs(1816) <= a and not b;
    outputs(1817) <= a;
    outputs(1818) <= not a;
    outputs(1819) <= b and not a;
    outputs(1820) <= not (a or b);
    outputs(1821) <= not a;
    outputs(1822) <= a xor b;
    outputs(1823) <= a;
    outputs(1824) <= not a;
    outputs(1825) <= b;
    outputs(1826) <= not (a xor b);
    outputs(1827) <= a xor b;
    outputs(1828) <= not b;
    outputs(1829) <= a or b;
    outputs(1830) <= not a;
    outputs(1831) <= a xor b;
    outputs(1832) <= not a;
    outputs(1833) <= not (a or b);
    outputs(1834) <= a xor b;
    outputs(1835) <= not (a xor b);
    outputs(1836) <= b;
    outputs(1837) <= not (a and b);
    outputs(1838) <= a;
    outputs(1839) <= a or b;
    outputs(1840) <= not b;
    outputs(1841) <= not b or a;
    outputs(1842) <= a;
    outputs(1843) <= a and not b;
    outputs(1844) <= not a;
    outputs(1845) <= not b;
    outputs(1846) <= b and not a;
    outputs(1847) <= not (a or b);
    outputs(1848) <= b;
    outputs(1849) <= not b;
    outputs(1850) <= a and b;
    outputs(1851) <= not b or a;
    outputs(1852) <= not (a xor b);
    outputs(1853) <= not b;
    outputs(1854) <= not a;
    outputs(1855) <= not (a or b);
    outputs(1856) <= a xor b;
    outputs(1857) <= not b;
    outputs(1858) <= a and not b;
    outputs(1859) <= a;
    outputs(1860) <= not (a xor b);
    outputs(1861) <= not b or a;
    outputs(1862) <= not b;
    outputs(1863) <= not b;
    outputs(1864) <= not a or b;
    outputs(1865) <= a;
    outputs(1866) <= a and b;
    outputs(1867) <= a and b;
    outputs(1868) <= not b;
    outputs(1869) <= not (a xor b);
    outputs(1870) <= a and b;
    outputs(1871) <= not (a or b);
    outputs(1872) <= a xor b;
    outputs(1873) <= not b;
    outputs(1874) <= a and not b;
    outputs(1875) <= b;
    outputs(1876) <= a;
    outputs(1877) <= b;
    outputs(1878) <= a and not b;
    outputs(1879) <= not a;
    outputs(1880) <= a and not b;
    outputs(1881) <= not a;
    outputs(1882) <= not (a xor b);
    outputs(1883) <= not b;
    outputs(1884) <= a and b;
    outputs(1885) <= not b;
    outputs(1886) <= a xor b;
    outputs(1887) <= b;
    outputs(1888) <= a xor b;
    outputs(1889) <= not (a xor b);
    outputs(1890) <= a and b;
    outputs(1891) <= b;
    outputs(1892) <= b;
    outputs(1893) <= not b;
    outputs(1894) <= b and not a;
    outputs(1895) <= not (a or b);
    outputs(1896) <= b and not a;
    outputs(1897) <= a;
    outputs(1898) <= a or b;
    outputs(1899) <= not a;
    outputs(1900) <= b;
    outputs(1901) <= a;
    outputs(1902) <= not b;
    outputs(1903) <= a and b;
    outputs(1904) <= b and not a;
    outputs(1905) <= a and not b;
    outputs(1906) <= a or b;
    outputs(1907) <= a xor b;
    outputs(1908) <= b;
    outputs(1909) <= not a;
    outputs(1910) <= not b or a;
    outputs(1911) <= b;
    outputs(1912) <= not b;
    outputs(1913) <= not a;
    outputs(1914) <= a and b;
    outputs(1915) <= a;
    outputs(1916) <= b and not a;
    outputs(1917) <= not a or b;
    outputs(1918) <= not a;
    outputs(1919) <= b and not a;
    outputs(1920) <= a xor b;
    outputs(1921) <= not (a and b);
    outputs(1922) <= a;
    outputs(1923) <= a;
    outputs(1924) <= a and not b;
    outputs(1925) <= not (a or b);
    outputs(1926) <= a xor b;
    outputs(1927) <= not a or b;
    outputs(1928) <= not b;
    outputs(1929) <= b and not a;
    outputs(1930) <= not b;
    outputs(1931) <= b and not a;
    outputs(1932) <= a xor b;
    outputs(1933) <= a or b;
    outputs(1934) <= b and not a;
    outputs(1935) <= b;
    outputs(1936) <= not (a or b);
    outputs(1937) <= not (a or b);
    outputs(1938) <= a;
    outputs(1939) <= not a;
    outputs(1940) <= not b;
    outputs(1941) <= a and b;
    outputs(1942) <= not a or b;
    outputs(1943) <= not (a xor b);
    outputs(1944) <= a and b;
    outputs(1945) <= not b;
    outputs(1946) <= a;
    outputs(1947) <= b;
    outputs(1948) <= b;
    outputs(1949) <= not b or a;
    outputs(1950) <= not (a and b);
    outputs(1951) <= not a;
    outputs(1952) <= not (a or b);
    outputs(1953) <= b;
    outputs(1954) <= a;
    outputs(1955) <= b;
    outputs(1956) <= not a;
    outputs(1957) <= not b;
    outputs(1958) <= b;
    outputs(1959) <= b;
    outputs(1960) <= not a;
    outputs(1961) <= a xor b;
    outputs(1962) <= a and b;
    outputs(1963) <= b;
    outputs(1964) <= not (a or b);
    outputs(1965) <= not b;
    outputs(1966) <= b;
    outputs(1967) <= a and b;
    outputs(1968) <= b and not a;
    outputs(1969) <= b;
    outputs(1970) <= b;
    outputs(1971) <= not b;
    outputs(1972) <= not a or b;
    outputs(1973) <= a;
    outputs(1974) <= not b;
    outputs(1975) <= a;
    outputs(1976) <= a;
    outputs(1977) <= not a or b;
    outputs(1978) <= a xor b;
    outputs(1979) <= not a;
    outputs(1980) <= not (a xor b);
    outputs(1981) <= a;
    outputs(1982) <= a and not b;
    outputs(1983) <= a and b;
    outputs(1984) <= a and not b;
    outputs(1985) <= a xor b;
    outputs(1986) <= not (a and b);
    outputs(1987) <= not b or a;
    outputs(1988) <= b;
    outputs(1989) <= not b;
    outputs(1990) <= a xor b;
    outputs(1991) <= not (a or b);
    outputs(1992) <= b;
    outputs(1993) <= not b;
    outputs(1994) <= not a;
    outputs(1995) <= a or b;
    outputs(1996) <= b and not a;
    outputs(1997) <= a;
    outputs(1998) <= not (a xor b);
    outputs(1999) <= b and not a;
    outputs(2000) <= a and b;
    outputs(2001) <= a and not b;
    outputs(2002) <= a and b;
    outputs(2003) <= a and not b;
    outputs(2004) <= not (a xor b);
    outputs(2005) <= not (a xor b);
    outputs(2006) <= b;
    outputs(2007) <= not (a or b);
    outputs(2008) <= a and not b;
    outputs(2009) <= not b;
    outputs(2010) <= b and not a;
    outputs(2011) <= b and not a;
    outputs(2012) <= b;
    outputs(2013) <= b;
    outputs(2014) <= b and not a;
    outputs(2015) <= not (a and b);
    outputs(2016) <= a xor b;
    outputs(2017) <= not a;
    outputs(2018) <= b;
    outputs(2019) <= a and not b;
    outputs(2020) <= a and not b;
    outputs(2021) <= not a or b;
    outputs(2022) <= b and not a;
    outputs(2023) <= not b;
    outputs(2024) <= a;
    outputs(2025) <= not (a xor b);
    outputs(2026) <= a and not b;
    outputs(2027) <= not (a xor b);
    outputs(2028) <= a and not b;
    outputs(2029) <= a and b;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= a;
    outputs(2032) <= b;
    outputs(2033) <= a;
    outputs(2034) <= b;
    outputs(2035) <= b;
    outputs(2036) <= not a;
    outputs(2037) <= a and not b;
    outputs(2038) <= b;
    outputs(2039) <= not b or a;
    outputs(2040) <= b and not a;
    outputs(2041) <= not b;
    outputs(2042) <= not a;
    outputs(2043) <= a xor b;
    outputs(2044) <= a xor b;
    outputs(2045) <= not b;
    outputs(2046) <= b and not a;
    outputs(2047) <= a and b;
    outputs(2048) <= a and b;
    outputs(2049) <= a and not b;
    outputs(2050) <= not a;
    outputs(2051) <= b;
    outputs(2052) <= not a;
    outputs(2053) <= not b or a;
    outputs(2054) <= not a;
    outputs(2055) <= a and not b;
    outputs(2056) <= a and not b;
    outputs(2057) <= a and not b;
    outputs(2058) <= b;
    outputs(2059) <= b;
    outputs(2060) <= a and not b;
    outputs(2061) <= a;
    outputs(2062) <= a;
    outputs(2063) <= b;
    outputs(2064) <= b and not a;
    outputs(2065) <= b;
    outputs(2066) <= not (a or b);
    outputs(2067) <= b;
    outputs(2068) <= not (a xor b);
    outputs(2069) <= a;
    outputs(2070) <= a and b;
    outputs(2071) <= a;
    outputs(2072) <= not b;
    outputs(2073) <= not a;
    outputs(2074) <= not (a and b);
    outputs(2075) <= a and b;
    outputs(2076) <= not (a and b);
    outputs(2077) <= b and not a;
    outputs(2078) <= b;
    outputs(2079) <= a and not b;
    outputs(2080) <= not (a xor b);
    outputs(2081) <= a xor b;
    outputs(2082) <= a and b;
    outputs(2083) <= not b;
    outputs(2084) <= a and b;
    outputs(2085) <= a and not b;
    outputs(2086) <= b and not a;
    outputs(2087) <= a and b;
    outputs(2088) <= not b;
    outputs(2089) <= not a;
    outputs(2090) <= not b or a;
    outputs(2091) <= b and not a;
    outputs(2092) <= b;
    outputs(2093) <= a and not b;
    outputs(2094) <= a and b;
    outputs(2095) <= a and b;
    outputs(2096) <= a and not b;
    outputs(2097) <= not a;
    outputs(2098) <= not b;
    outputs(2099) <= b;
    outputs(2100) <= b and not a;
    outputs(2101) <= not (a xor b);
    outputs(2102) <= a and not b;
    outputs(2103) <= b;
    outputs(2104) <= not a;
    outputs(2105) <= not a;
    outputs(2106) <= b and not a;
    outputs(2107) <= a xor b;
    outputs(2108) <= b and not a;
    outputs(2109) <= not b;
    outputs(2110) <= not (a and b);
    outputs(2111) <= b;
    outputs(2112) <= b;
    outputs(2113) <= b and not a;
    outputs(2114) <= not (a xor b);
    outputs(2115) <= b and not a;
    outputs(2116) <= not (a and b);
    outputs(2117) <= a;
    outputs(2118) <= b;
    outputs(2119) <= a;
    outputs(2120) <= not (a and b);
    outputs(2121) <= b and not a;
    outputs(2122) <= a and not b;
    outputs(2123) <= a xor b;
    outputs(2124) <= not b;
    outputs(2125) <= a;
    outputs(2126) <= not (a or b);
    outputs(2127) <= a and b;
    outputs(2128) <= b;
    outputs(2129) <= b;
    outputs(2130) <= not b;
    outputs(2131) <= not a;
    outputs(2132) <= b and not a;
    outputs(2133) <= not a or b;
    outputs(2134) <= not b;
    outputs(2135) <= b;
    outputs(2136) <= a xor b;
    outputs(2137) <= a;
    outputs(2138) <= not b;
    outputs(2139) <= b and not a;
    outputs(2140) <= not b;
    outputs(2141) <= b;
    outputs(2142) <= a and b;
    outputs(2143) <= not a;
    outputs(2144) <= b and not a;
    outputs(2145) <= not a;
    outputs(2146) <= a and not b;
    outputs(2147) <= a xor b;
    outputs(2148) <= a and b;
    outputs(2149) <= a;
    outputs(2150) <= a xor b;
    outputs(2151) <= a;
    outputs(2152) <= not (a or b);
    outputs(2153) <= a;
    outputs(2154) <= not (a or b);
    outputs(2155) <= not a;
    outputs(2156) <= a;
    outputs(2157) <= a;
    outputs(2158) <= a and b;
    outputs(2159) <= a and b;
    outputs(2160) <= a and b;
    outputs(2161) <= a;
    outputs(2162) <= a and not b;
    outputs(2163) <= not b;
    outputs(2164) <= a xor b;
    outputs(2165) <= a and b;
    outputs(2166) <= a and not b;
    outputs(2167) <= not (a or b);
    outputs(2168) <= b;
    outputs(2169) <= not (a or b);
    outputs(2170) <= a;
    outputs(2171) <= a;
    outputs(2172) <= not (a or b);
    outputs(2173) <= a;
    outputs(2174) <= not a;
    outputs(2175) <= not b;
    outputs(2176) <= not a;
    outputs(2177) <= a xor b;
    outputs(2178) <= a and not b;
    outputs(2179) <= b;
    outputs(2180) <= b;
    outputs(2181) <= a and b;
    outputs(2182) <= a and not b;
    outputs(2183) <= a;
    outputs(2184) <= a;
    outputs(2185) <= a and b;
    outputs(2186) <= a;
    outputs(2187) <= not a;
    outputs(2188) <= not a;
    outputs(2189) <= a and not b;
    outputs(2190) <= a and b;
    outputs(2191) <= a xor b;
    outputs(2192) <= a and b;
    outputs(2193) <= b;
    outputs(2194) <= not (a or b);
    outputs(2195) <= a and b;
    outputs(2196) <= a;
    outputs(2197) <= b and not a;
    outputs(2198) <= a;
    outputs(2199) <= b and not a;
    outputs(2200) <= b;
    outputs(2201) <= b and not a;
    outputs(2202) <= b and not a;
    outputs(2203) <= a;
    outputs(2204) <= b;
    outputs(2205) <= a or b;
    outputs(2206) <= b and not a;
    outputs(2207) <= not a;
    outputs(2208) <= not a;
    outputs(2209) <= not a;
    outputs(2210) <= not (a or b);
    outputs(2211) <= a and not b;
    outputs(2212) <= a and b;
    outputs(2213) <= a;
    outputs(2214) <= b and not a;
    outputs(2215) <= not a;
    outputs(2216) <= b and not a;
    outputs(2217) <= b;
    outputs(2218) <= not b;
    outputs(2219) <= b and not a;
    outputs(2220) <= not (a xor b);
    outputs(2221) <= b and not a;
    outputs(2222) <= b;
    outputs(2223) <= not a;
    outputs(2224) <= a xor b;
    outputs(2225) <= b;
    outputs(2226) <= not (a xor b);
    outputs(2227) <= not b;
    outputs(2228) <= b;
    outputs(2229) <= not a;
    outputs(2230) <= a and b;
    outputs(2231) <= a xor b;
    outputs(2232) <= a and b;
    outputs(2233) <= a or b;
    outputs(2234) <= not a;
    outputs(2235) <= b and not a;
    outputs(2236) <= not b;
    outputs(2237) <= not (a or b);
    outputs(2238) <= b;
    outputs(2239) <= a;
    outputs(2240) <= not (a xor b);
    outputs(2241) <= a;
    outputs(2242) <= not a or b;
    outputs(2243) <= not b;
    outputs(2244) <= a and b;
    outputs(2245) <= b and not a;
    outputs(2246) <= b;
    outputs(2247) <= a or b;
    outputs(2248) <= not (a and b);
    outputs(2249) <= not b;
    outputs(2250) <= a;
    outputs(2251) <= not a;
    outputs(2252) <= not a;
    outputs(2253) <= a and not b;
    outputs(2254) <= b;
    outputs(2255) <= a xor b;
    outputs(2256) <= not a;
    outputs(2257) <= a;
    outputs(2258) <= b;
    outputs(2259) <= a and not b;
    outputs(2260) <= not b;
    outputs(2261) <= a;
    outputs(2262) <= not a;
    outputs(2263) <= not a;
    outputs(2264) <= a and not b;
    outputs(2265) <= a and not b;
    outputs(2266) <= b and not a;
    outputs(2267) <= not a;
    outputs(2268) <= a;
    outputs(2269) <= a and not b;
    outputs(2270) <= not (a or b);
    outputs(2271) <= not a;
    outputs(2272) <= not a;
    outputs(2273) <= not a;
    outputs(2274) <= a xor b;
    outputs(2275) <= b;
    outputs(2276) <= not (a and b);
    outputs(2277) <= b;
    outputs(2278) <= not a;
    outputs(2279) <= not (a or b);
    outputs(2280) <= not b;
    outputs(2281) <= a xor b;
    outputs(2282) <= not (a xor b);
    outputs(2283) <= a and b;
    outputs(2284) <= b;
    outputs(2285) <= a;
    outputs(2286) <= b and not a;
    outputs(2287) <= not b or a;
    outputs(2288) <= a;
    outputs(2289) <= not b or a;
    outputs(2290) <= not a;
    outputs(2291) <= not b;
    outputs(2292) <= not (a xor b);
    outputs(2293) <= a and b;
    outputs(2294) <= not b;
    outputs(2295) <= not a or b;
    outputs(2296) <= a;
    outputs(2297) <= not (a or b);
    outputs(2298) <= a xor b;
    outputs(2299) <= not a or b;
    outputs(2300) <= a or b;
    outputs(2301) <= a;
    outputs(2302) <= b;
    outputs(2303) <= a and b;
    outputs(2304) <= not b;
    outputs(2305) <= not b;
    outputs(2306) <= a xor b;
    outputs(2307) <= a;
    outputs(2308) <= a and not b;
    outputs(2309) <= b;
    outputs(2310) <= not a or b;
    outputs(2311) <= not b;
    outputs(2312) <= b;
    outputs(2313) <= a and b;
    outputs(2314) <= a and not b;
    outputs(2315) <= not a;
    outputs(2316) <= a;
    outputs(2317) <= a and not b;
    outputs(2318) <= not (a xor b);
    outputs(2319) <= a;
    outputs(2320) <= not (a xor b);
    outputs(2321) <= a and b;
    outputs(2322) <= not (a xor b);
    outputs(2323) <= a;
    outputs(2324) <= a and b;
    outputs(2325) <= a xor b;
    outputs(2326) <= a xor b;
    outputs(2327) <= a;
    outputs(2328) <= not (a or b);
    outputs(2329) <= b;
    outputs(2330) <= not b;
    outputs(2331) <= not a;
    outputs(2332) <= not a;
    outputs(2333) <= b;
    outputs(2334) <= a and not b;
    outputs(2335) <= a and b;
    outputs(2336) <= not (a xor b);
    outputs(2337) <= not (a and b);
    outputs(2338) <= not (a or b);
    outputs(2339) <= b and not a;
    outputs(2340) <= a and b;
    outputs(2341) <= not b or a;
    outputs(2342) <= a and b;
    outputs(2343) <= a;
    outputs(2344) <= not (a xor b);
    outputs(2345) <= a and b;
    outputs(2346) <= b;
    outputs(2347) <= not (a xor b);
    outputs(2348) <= a and b;
    outputs(2349) <= a xor b;
    outputs(2350) <= not (a xor b);
    outputs(2351) <= a and b;
    outputs(2352) <= not a;
    outputs(2353) <= not a;
    outputs(2354) <= not (a xor b);
    outputs(2355) <= a and b;
    outputs(2356) <= a and not b;
    outputs(2357) <= not b;
    outputs(2358) <= a;
    outputs(2359) <= not b or a;
    outputs(2360) <= b;
    outputs(2361) <= a xor b;
    outputs(2362) <= a;
    outputs(2363) <= b;
    outputs(2364) <= not b;
    outputs(2365) <= a;
    outputs(2366) <= not b;
    outputs(2367) <= not a;
    outputs(2368) <= not (a or b);
    outputs(2369) <= not b;
    outputs(2370) <= b;
    outputs(2371) <= a and b;
    outputs(2372) <= not (a and b);
    outputs(2373) <= not b;
    outputs(2374) <= a xor b;
    outputs(2375) <= not b;
    outputs(2376) <= b and not a;
    outputs(2377) <= b and not a;
    outputs(2378) <= a and not b;
    outputs(2379) <= b;
    outputs(2380) <= b and not a;
    outputs(2381) <= not a;
    outputs(2382) <= a;
    outputs(2383) <= a and not b;
    outputs(2384) <= a and b;
    outputs(2385) <= not (a or b);
    outputs(2386) <= a and not b;
    outputs(2387) <= a;
    outputs(2388) <= not (a or b);
    outputs(2389) <= not a;
    outputs(2390) <= not (a and b);
    outputs(2391) <= a and b;
    outputs(2392) <= not a;
    outputs(2393) <= not (a or b);
    outputs(2394) <= a and b;
    outputs(2395) <= not a;
    outputs(2396) <= not (a xor b);
    outputs(2397) <= b and not a;
    outputs(2398) <= a and b;
    outputs(2399) <= b;
    outputs(2400) <= not a or b;
    outputs(2401) <= not a;
    outputs(2402) <= not b;
    outputs(2403) <= a and not b;
    outputs(2404) <= a;
    outputs(2405) <= not (a or b);
    outputs(2406) <= not a;
    outputs(2407) <= not (a xor b);
    outputs(2408) <= a and b;
    outputs(2409) <= not (a or b);
    outputs(2410) <= not (a xor b);
    outputs(2411) <= a xor b;
    outputs(2412) <= not (a or b);
    outputs(2413) <= a and b;
    outputs(2414) <= a and not b;
    outputs(2415) <= a;
    outputs(2416) <= not (a or b);
    outputs(2417) <= not (a or b);
    outputs(2418) <= a;
    outputs(2419) <= not b;
    outputs(2420) <= not a;
    outputs(2421) <= a or b;
    outputs(2422) <= a;
    outputs(2423) <= a and not b;
    outputs(2424) <= b;
    outputs(2425) <= not b;
    outputs(2426) <= a and not b;
    outputs(2427) <= not b;
    outputs(2428) <= a or b;
    outputs(2429) <= b and not a;
    outputs(2430) <= not (a or b);
    outputs(2431) <= a;
    outputs(2432) <= not a;
    outputs(2433) <= a and b;
    outputs(2434) <= a;
    outputs(2435) <= not (a or b);
    outputs(2436) <= a and not b;
    outputs(2437) <= not (a and b);
    outputs(2438) <= a;
    outputs(2439) <= a;
    outputs(2440) <= a and not b;
    outputs(2441) <= a and not b;
    outputs(2442) <= a;
    outputs(2443) <= a;
    outputs(2444) <= b and not a;
    outputs(2445) <= a;
    outputs(2446) <= b and not a;
    outputs(2447) <= b;
    outputs(2448) <= b and not a;
    outputs(2449) <= not b or a;
    outputs(2450) <= not (a or b);
    outputs(2451) <= not a;
    outputs(2452) <= a or b;
    outputs(2453) <= not (a xor b);
    outputs(2454) <= not (a xor b);
    outputs(2455) <= a and not b;
    outputs(2456) <= not a or b;
    outputs(2457) <= a xor b;
    outputs(2458) <= a and not b;
    outputs(2459) <= b;
    outputs(2460) <= not (a or b);
    outputs(2461) <= a;
    outputs(2462) <= not (a or b);
    outputs(2463) <= not (a xor b);
    outputs(2464) <= not b;
    outputs(2465) <= not b;
    outputs(2466) <= a and b;
    outputs(2467) <= a;
    outputs(2468) <= a xor b;
    outputs(2469) <= b and not a;
    outputs(2470) <= b;
    outputs(2471) <= not a;
    outputs(2472) <= b;
    outputs(2473) <= a;
    outputs(2474) <= not (a or b);
    outputs(2475) <= a;
    outputs(2476) <= not (a and b);
    outputs(2477) <= b and not a;
    outputs(2478) <= not a;
    outputs(2479) <= a and b;
    outputs(2480) <= not (a xor b);
    outputs(2481) <= a xor b;
    outputs(2482) <= a and b;
    outputs(2483) <= b and not a;
    outputs(2484) <= not (a and b);
    outputs(2485) <= b;
    outputs(2486) <= not (a xor b);
    outputs(2487) <= a and b;
    outputs(2488) <= a and b;
    outputs(2489) <= a and b;
    outputs(2490) <= a and not b;
    outputs(2491) <= not b;
    outputs(2492) <= a;
    outputs(2493) <= b and not a;
    outputs(2494) <= b;
    outputs(2495) <= not (a or b);
    outputs(2496) <= not a;
    outputs(2497) <= a xor b;
    outputs(2498) <= a xor b;
    outputs(2499) <= not (a xor b);
    outputs(2500) <= a and not b;
    outputs(2501) <= a;
    outputs(2502) <= not (a or b);
    outputs(2503) <= a;
    outputs(2504) <= a and not b;
    outputs(2505) <= a and b;
    outputs(2506) <= a and b;
    outputs(2507) <= a and b;
    outputs(2508) <= not a or b;
    outputs(2509) <= not (a xor b);
    outputs(2510) <= not b;
    outputs(2511) <= not b;
    outputs(2512) <= a and not b;
    outputs(2513) <= a;
    outputs(2514) <= a and not b;
    outputs(2515) <= a xor b;
    outputs(2516) <= not a or b;
    outputs(2517) <= a;
    outputs(2518) <= a and not b;
    outputs(2519) <= a and not b;
    outputs(2520) <= not a;
    outputs(2521) <= a and b;
    outputs(2522) <= not a;
    outputs(2523) <= b;
    outputs(2524) <= a and not b;
    outputs(2525) <= not b or a;
    outputs(2526) <= a xor b;
    outputs(2527) <= a xor b;
    outputs(2528) <= a;
    outputs(2529) <= not (a or b);
    outputs(2530) <= a xor b;
    outputs(2531) <= b and not a;
    outputs(2532) <= b;
    outputs(2533) <= b;
    outputs(2534) <= a;
    outputs(2535) <= not (a or b);
    outputs(2536) <= a and b;
    outputs(2537) <= a and b;
    outputs(2538) <= a and not b;
    outputs(2539) <= a xor b;
    outputs(2540) <= a;
    outputs(2541) <= a;
    outputs(2542) <= not b or a;
    outputs(2543) <= a;
    outputs(2544) <= a and b;
    outputs(2545) <= not (a or b);
    outputs(2546) <= a or b;
    outputs(2547) <= not (a xor b);
    outputs(2548) <= a xor b;
    outputs(2549) <= a xor b;
    outputs(2550) <= not a;
    outputs(2551) <= a xor b;
    outputs(2552) <= a xor b;
    outputs(2553) <= a;
    outputs(2554) <= not a;
    outputs(2555) <= not (a or b);
    outputs(2556) <= a or b;
    outputs(2557) <= b and not a;
    outputs(2558) <= not (a or b);
    outputs(2559) <= a;
    outputs(2560) <= b;
    outputs(2561) <= not b;
    outputs(2562) <= not b or a;
    outputs(2563) <= a and not b;
    outputs(2564) <= not (a and b);
    outputs(2565) <= not b;
    outputs(2566) <= a or b;
    outputs(2567) <= a and b;
    outputs(2568) <= not a;
    outputs(2569) <= a xor b;
    outputs(2570) <= not a;
    outputs(2571) <= a and b;
    outputs(2572) <= not (a or b);
    outputs(2573) <= a xor b;
    outputs(2574) <= b;
    outputs(2575) <= b;
    outputs(2576) <= a xor b;
    outputs(2577) <= a and b;
    outputs(2578) <= not (a and b);
    outputs(2579) <= not (a xor b);
    outputs(2580) <= not a;
    outputs(2581) <= b;
    outputs(2582) <= a and b;
    outputs(2583) <= not b;
    outputs(2584) <= a and b;
    outputs(2585) <= not (a and b);
    outputs(2586) <= a xor b;
    outputs(2587) <= not (a or b);
    outputs(2588) <= a and not b;
    outputs(2589) <= not (a xor b);
    outputs(2590) <= not b;
    outputs(2591) <= not (a and b);
    outputs(2592) <= not b;
    outputs(2593) <= not b;
    outputs(2594) <= a xor b;
    outputs(2595) <= a and not b;
    outputs(2596) <= not b;
    outputs(2597) <= not (a xor b);
    outputs(2598) <= not (a xor b);
    outputs(2599) <= a xor b;
    outputs(2600) <= b;
    outputs(2601) <= not (a xor b);
    outputs(2602) <= a and b;
    outputs(2603) <= a xor b;
    outputs(2604) <= a;
    outputs(2605) <= a or b;
    outputs(2606) <= not a or b;
    outputs(2607) <= a or b;
    outputs(2608) <= not (a xor b);
    outputs(2609) <= not b;
    outputs(2610) <= not (a and b);
    outputs(2611) <= a and not b;
    outputs(2612) <= a and b;
    outputs(2613) <= not (a xor b);
    outputs(2614) <= not (a or b);
    outputs(2615) <= not b;
    outputs(2616) <= not b;
    outputs(2617) <= not (a xor b);
    outputs(2618) <= not b;
    outputs(2619) <= a xor b;
    outputs(2620) <= not (a xor b);
    outputs(2621) <= a and b;
    outputs(2622) <= b and not a;
    outputs(2623) <= not (a xor b);
    outputs(2624) <= not a;
    outputs(2625) <= not b;
    outputs(2626) <= not b;
    outputs(2627) <= a and not b;
    outputs(2628) <= b;
    outputs(2629) <= a xor b;
    outputs(2630) <= a;
    outputs(2631) <= not (a xor b);
    outputs(2632) <= b;
    outputs(2633) <= a;
    outputs(2634) <= a xor b;
    outputs(2635) <= not a;
    outputs(2636) <= b;
    outputs(2637) <= b and not a;
    outputs(2638) <= not a;
    outputs(2639) <= a;
    outputs(2640) <= not b or a;
    outputs(2641) <= b and not a;
    outputs(2642) <= a or b;
    outputs(2643) <= a and b;
    outputs(2644) <= not b;
    outputs(2645) <= not (a xor b);
    outputs(2646) <= a;
    outputs(2647) <= a xor b;
    outputs(2648) <= not a or b;
    outputs(2649) <= not (a xor b);
    outputs(2650) <= a and not b;
    outputs(2651) <= a and not b;
    outputs(2652) <= not b;
    outputs(2653) <= not b or a;
    outputs(2654) <= not (a xor b);
    outputs(2655) <= b and not a;
    outputs(2656) <= not (a or b);
    outputs(2657) <= b and not a;
    outputs(2658) <= a xor b;
    outputs(2659) <= not a;
    outputs(2660) <= not (a xor b);
    outputs(2661) <= b;
    outputs(2662) <= a and not b;
    outputs(2663) <= not a;
    outputs(2664) <= a xor b;
    outputs(2665) <= a and not b;
    outputs(2666) <= a;
    outputs(2667) <= not (a xor b);
    outputs(2668) <= not a or b;
    outputs(2669) <= a;
    outputs(2670) <= a;
    outputs(2671) <= a xor b;
    outputs(2672) <= not (a xor b);
    outputs(2673) <= a and not b;
    outputs(2674) <= not (a or b);
    outputs(2675) <= not b;
    outputs(2676) <= b and not a;
    outputs(2677) <= not a;
    outputs(2678) <= not (a or b);
    outputs(2679) <= b;
    outputs(2680) <= a and not b;
    outputs(2681) <= a;
    outputs(2682) <= not b or a;
    outputs(2683) <= a or b;
    outputs(2684) <= not a;
    outputs(2685) <= b;
    outputs(2686) <= not (a or b);
    outputs(2687) <= a and b;
    outputs(2688) <= a xor b;
    outputs(2689) <= a xor b;
    outputs(2690) <= a and b;
    outputs(2691) <= b;
    outputs(2692) <= not b or a;
    outputs(2693) <= a xor b;
    outputs(2694) <= a;
    outputs(2695) <= not a;
    outputs(2696) <= a and b;
    outputs(2697) <= b;
    outputs(2698) <= a and not b;
    outputs(2699) <= a;
    outputs(2700) <= b and not a;
    outputs(2701) <= a;
    outputs(2702) <= a or b;
    outputs(2703) <= a xor b;
    outputs(2704) <= not b;
    outputs(2705) <= a;
    outputs(2706) <= a or b;
    outputs(2707) <= not a;
    outputs(2708) <= not b;
    outputs(2709) <= not a or b;
    outputs(2710) <= a xor b;
    outputs(2711) <= a and not b;
    outputs(2712) <= a xor b;
    outputs(2713) <= not a;
    outputs(2714) <= not b;
    outputs(2715) <= not b;
    outputs(2716) <= b;
    outputs(2717) <= a and not b;
    outputs(2718) <= not a;
    outputs(2719) <= a and b;
    outputs(2720) <= a;
    outputs(2721) <= a xor b;
    outputs(2722) <= not (a or b);
    outputs(2723) <= not (a xor b);
    outputs(2724) <= not a;
    outputs(2725) <= a;
    outputs(2726) <= b and not a;
    outputs(2727) <= a and not b;
    outputs(2728) <= a xor b;
    outputs(2729) <= not (a and b);
    outputs(2730) <= not b;
    outputs(2731) <= a xor b;
    outputs(2732) <= a and not b;
    outputs(2733) <= a and not b;
    outputs(2734) <= b;
    outputs(2735) <= not a;
    outputs(2736) <= a;
    outputs(2737) <= not (a or b);
    outputs(2738) <= a and b;
    outputs(2739) <= b;
    outputs(2740) <= b and not a;
    outputs(2741) <= b and not a;
    outputs(2742) <= a;
    outputs(2743) <= not (a xor b);
    outputs(2744) <= not (a xor b);
    outputs(2745) <= not a;
    outputs(2746) <= b and not a;
    outputs(2747) <= not b;
    outputs(2748) <= b and not a;
    outputs(2749) <= not b;
    outputs(2750) <= a;
    outputs(2751) <= a;
    outputs(2752) <= not b;
    outputs(2753) <= a xor b;
    outputs(2754) <= a xor b;
    outputs(2755) <= not a;
    outputs(2756) <= not b or a;
    outputs(2757) <= not a;
    outputs(2758) <= b;
    outputs(2759) <= b;
    outputs(2760) <= a;
    outputs(2761) <= not b;
    outputs(2762) <= not b or a;
    outputs(2763) <= a or b;
    outputs(2764) <= a xor b;
    outputs(2765) <= not b;
    outputs(2766) <= a;
    outputs(2767) <= not (a or b);
    outputs(2768) <= a;
    outputs(2769) <= not (a and b);
    outputs(2770) <= b;
    outputs(2771) <= a and b;
    outputs(2772) <= not a;
    outputs(2773) <= a;
    outputs(2774) <= a xor b;
    outputs(2775) <= not (a xor b);
    outputs(2776) <= b and not a;
    outputs(2777) <= not b or a;
    outputs(2778) <= a and not b;
    outputs(2779) <= b;
    outputs(2780) <= not a or b;
    outputs(2781) <= b and not a;
    outputs(2782) <= a and not b;
    outputs(2783) <= a or b;
    outputs(2784) <= not (a xor b);
    outputs(2785) <= b and not a;
    outputs(2786) <= not a;
    outputs(2787) <= a xor b;
    outputs(2788) <= not b;
    outputs(2789) <= b and not a;
    outputs(2790) <= not (a and b);
    outputs(2791) <= a xor b;
    outputs(2792) <= a xor b;
    outputs(2793) <= not (a xor b);
    outputs(2794) <= not b or a;
    outputs(2795) <= not b;
    outputs(2796) <= not (a or b);
    outputs(2797) <= a;
    outputs(2798) <= not a;
    outputs(2799) <= b;
    outputs(2800) <= not a;
    outputs(2801) <= not a or b;
    outputs(2802) <= not a;
    outputs(2803) <= not a;
    outputs(2804) <= a or b;
    outputs(2805) <= not a or b;
    outputs(2806) <= not b;
    outputs(2807) <= b;
    outputs(2808) <= a and b;
    outputs(2809) <= a;
    outputs(2810) <= b and not a;
    outputs(2811) <= not (a or b);
    outputs(2812) <= a xor b;
    outputs(2813) <= a xor b;
    outputs(2814) <= a;
    outputs(2815) <= not a;
    outputs(2816) <= a xor b;
    outputs(2817) <= a;
    outputs(2818) <= not (a or b);
    outputs(2819) <= b;
    outputs(2820) <= a and b;
    outputs(2821) <= not b;
    outputs(2822) <= a and not b;
    outputs(2823) <= not b;
    outputs(2824) <= a and not b;
    outputs(2825) <= not (a xor b);
    outputs(2826) <= not a;
    outputs(2827) <= a and not b;
    outputs(2828) <= not b;
    outputs(2829) <= not b;
    outputs(2830) <= not (a xor b);
    outputs(2831) <= a xor b;
    outputs(2832) <= a and b;
    outputs(2833) <= not (a xor b);
    outputs(2834) <= not b;
    outputs(2835) <= b;
    outputs(2836) <= a;
    outputs(2837) <= a xor b;
    outputs(2838) <= not (a or b);
    outputs(2839) <= not (a xor b);
    outputs(2840) <= a;
    outputs(2841) <= not a;
    outputs(2842) <= not a or b;
    outputs(2843) <= not a;
    outputs(2844) <= a xor b;
    outputs(2845) <= not a;
    outputs(2846) <= b and not a;
    outputs(2847) <= not b;
    outputs(2848) <= a;
    outputs(2849) <= a and b;
    outputs(2850) <= a or b;
    outputs(2851) <= not a;
    outputs(2852) <= a or b;
    outputs(2853) <= not (a xor b);
    outputs(2854) <= a xor b;
    outputs(2855) <= b;
    outputs(2856) <= not (a xor b);
    outputs(2857) <= not a or b;
    outputs(2858) <= a;
    outputs(2859) <= a xor b;
    outputs(2860) <= b;
    outputs(2861) <= b;
    outputs(2862) <= a xor b;
    outputs(2863) <= a and b;
    outputs(2864) <= not a;
    outputs(2865) <= b and not a;
    outputs(2866) <= a xor b;
    outputs(2867) <= a and b;
    outputs(2868) <= not (a xor b);
    outputs(2869) <= not (a or b);
    outputs(2870) <= b and not a;
    outputs(2871) <= a xor b;
    outputs(2872) <= not a;
    outputs(2873) <= not (a or b);
    outputs(2874) <= a xor b;
    outputs(2875) <= a or b;
    outputs(2876) <= a or b;
    outputs(2877) <= a xor b;
    outputs(2878) <= a and not b;
    outputs(2879) <= not a or b;
    outputs(2880) <= a or b;
    outputs(2881) <= a xor b;
    outputs(2882) <= not (a xor b);
    outputs(2883) <= a;
    outputs(2884) <= not (a and b);
    outputs(2885) <= not b or a;
    outputs(2886) <= not b or a;
    outputs(2887) <= a;
    outputs(2888) <= a;
    outputs(2889) <= a and b;
    outputs(2890) <= a xor b;
    outputs(2891) <= not a;
    outputs(2892) <= not a or b;
    outputs(2893) <= b;
    outputs(2894) <= not (a xor b);
    outputs(2895) <= not b or a;
    outputs(2896) <= not a;
    outputs(2897) <= a and not b;
    outputs(2898) <= a;
    outputs(2899) <= not (a or b);
    outputs(2900) <= not a;
    outputs(2901) <= a xor b;
    outputs(2902) <= not b;
    outputs(2903) <= a and not b;
    outputs(2904) <= a or b;
    outputs(2905) <= not (a or b);
    outputs(2906) <= a or b;
    outputs(2907) <= not (a xor b);
    outputs(2908) <= a;
    outputs(2909) <= b;
    outputs(2910) <= a xor b;
    outputs(2911) <= not a;
    outputs(2912) <= a and b;
    outputs(2913) <= a and b;
    outputs(2914) <= not (a and b);
    outputs(2915) <= not a;
    outputs(2916) <= a xor b;
    outputs(2917) <= not (a xor b);
    outputs(2918) <= not b;
    outputs(2919) <= not (a or b);
    outputs(2920) <= b;
    outputs(2921) <= not a;
    outputs(2922) <= a xor b;
    outputs(2923) <= a xor b;
    outputs(2924) <= a xor b;
    outputs(2925) <= a xor b;
    outputs(2926) <= not a;
    outputs(2927) <= a xor b;
    outputs(2928) <= not (a xor b);
    outputs(2929) <= not b;
    outputs(2930) <= a and not b;
    outputs(2931) <= a and not b;
    outputs(2932) <= a;
    outputs(2933) <= a xor b;
    outputs(2934) <= not (a xor b);
    outputs(2935) <= not a or b;
    outputs(2936) <= a xor b;
    outputs(2937) <= not a;
    outputs(2938) <= a xor b;
    outputs(2939) <= a xor b;
    outputs(2940) <= a xor b;
    outputs(2941) <= a;
    outputs(2942) <= not (a xor b);
    outputs(2943) <= not a;
    outputs(2944) <= not b;
    outputs(2945) <= not (a xor b);
    outputs(2946) <= a xor b;
    outputs(2947) <= not b;
    outputs(2948) <= not (a and b);
    outputs(2949) <= a;
    outputs(2950) <= not a;
    outputs(2951) <= not b;
    outputs(2952) <= b;
    outputs(2953) <= b;
    outputs(2954) <= not (a xor b);
    outputs(2955) <= a and b;
    outputs(2956) <= not a or b;
    outputs(2957) <= b;
    outputs(2958) <= a and not b;
    outputs(2959) <= not (a xor b);
    outputs(2960) <= not (a or b);
    outputs(2961) <= a;
    outputs(2962) <= not a;
    outputs(2963) <= b and not a;
    outputs(2964) <= not b;
    outputs(2965) <= b;
    outputs(2966) <= a;
    outputs(2967) <= a;
    outputs(2968) <= not a;
    outputs(2969) <= not a;
    outputs(2970) <= b and not a;
    outputs(2971) <= a;
    outputs(2972) <= not a;
    outputs(2973) <= a and not b;
    outputs(2974) <= a and not b;
    outputs(2975) <= not a or b;
    outputs(2976) <= not b;
    outputs(2977) <= b;
    outputs(2978) <= a or b;
    outputs(2979) <= a and b;
    outputs(2980) <= b;
    outputs(2981) <= b and not a;
    outputs(2982) <= a xor b;
    outputs(2983) <= not b;
    outputs(2984) <= not (a xor b);
    outputs(2985) <= not (a xor b);
    outputs(2986) <= not (a or b);
    outputs(2987) <= not b;
    outputs(2988) <= not (a xor b);
    outputs(2989) <= a and not b;
    outputs(2990) <= a or b;
    outputs(2991) <= a and not b;
    outputs(2992) <= a xor b;
    outputs(2993) <= a or b;
    outputs(2994) <= b;
    outputs(2995) <= not b;
    outputs(2996) <= a xor b;
    outputs(2997) <= a and not b;
    outputs(2998) <= a and not b;
    outputs(2999) <= a;
    outputs(3000) <= not a;
    outputs(3001) <= a and not b;
    outputs(3002) <= a and b;
    outputs(3003) <= not a;
    outputs(3004) <= not b;
    outputs(3005) <= not b or a;
    outputs(3006) <= b;
    outputs(3007) <= b and not a;
    outputs(3008) <= not a or b;
    outputs(3009) <= not a;
    outputs(3010) <= b and not a;
    outputs(3011) <= not a;
    outputs(3012) <= a and not b;
    outputs(3013) <= not (a xor b);
    outputs(3014) <= b;
    outputs(3015) <= not (a or b);
    outputs(3016) <= not a or b;
    outputs(3017) <= a xor b;
    outputs(3018) <= a and b;
    outputs(3019) <= not a;
    outputs(3020) <= a;
    outputs(3021) <= a and not b;
    outputs(3022) <= not (a xor b);
    outputs(3023) <= not (a xor b);
    outputs(3024) <= a and not b;
    outputs(3025) <= not (a or b);
    outputs(3026) <= b;
    outputs(3027) <= b;
    outputs(3028) <= b;
    outputs(3029) <= not b or a;
    outputs(3030) <= not b;
    outputs(3031) <= not (a and b);
    outputs(3032) <= not (a xor b);
    outputs(3033) <= not a;
    outputs(3034) <= not (a xor b);
    outputs(3035) <= not b;
    outputs(3036) <= a xor b;
    outputs(3037) <= b;
    outputs(3038) <= a or b;
    outputs(3039) <= not b;
    outputs(3040) <= not b or a;
    outputs(3041) <= a and b;
    outputs(3042) <= not b;
    outputs(3043) <= not (a xor b);
    outputs(3044) <= not (a xor b);
    outputs(3045) <= not (a or b);
    outputs(3046) <= not a or b;
    outputs(3047) <= b;
    outputs(3048) <= a xor b;
    outputs(3049) <= a and b;
    outputs(3050) <= a xor b;
    outputs(3051) <= a xor b;
    outputs(3052) <= not b;
    outputs(3053) <= a xor b;
    outputs(3054) <= a xor b;
    outputs(3055) <= b and not a;
    outputs(3056) <= a and b;
    outputs(3057) <= not a or b;
    outputs(3058) <= not b;
    outputs(3059) <= a;
    outputs(3060) <= not b;
    outputs(3061) <= not (a xor b);
    outputs(3062) <= b;
    outputs(3063) <= not b;
    outputs(3064) <= b and not a;
    outputs(3065) <= a;
    outputs(3066) <= not a;
    outputs(3067) <= not a;
    outputs(3068) <= a;
    outputs(3069) <= not (a or b);
    outputs(3070) <= b;
    outputs(3071) <= not b;
    outputs(3072) <= not b;
    outputs(3073) <= a and b;
    outputs(3074) <= b;
    outputs(3075) <= a and b;
    outputs(3076) <= a and b;
    outputs(3077) <= not (a or b);
    outputs(3078) <= a;
    outputs(3079) <= a;
    outputs(3080) <= b;
    outputs(3081) <= not a;
    outputs(3082) <= b;
    outputs(3083) <= not a;
    outputs(3084) <= not (a xor b);
    outputs(3085) <= b;
    outputs(3086) <= b and not a;
    outputs(3087) <= a;
    outputs(3088) <= not a or b;
    outputs(3089) <= not (a or b);
    outputs(3090) <= not b;
    outputs(3091) <= a or b;
    outputs(3092) <= a xor b;
    outputs(3093) <= not a;
    outputs(3094) <= b;
    outputs(3095) <= b;
    outputs(3096) <= a xor b;
    outputs(3097) <= not (a xor b);
    outputs(3098) <= not a;
    outputs(3099) <= b;
    outputs(3100) <= a;
    outputs(3101) <= not b;
    outputs(3102) <= b and not a;
    outputs(3103) <= a;
    outputs(3104) <= not a;
    outputs(3105) <= not a;
    outputs(3106) <= a and not b;
    outputs(3107) <= not b;
    outputs(3108) <= not (a or b);
    outputs(3109) <= not b;
    outputs(3110) <= not a;
    outputs(3111) <= a and b;
    outputs(3112) <= a;
    outputs(3113) <= b and not a;
    outputs(3114) <= a;
    outputs(3115) <= a xor b;
    outputs(3116) <= not b;
    outputs(3117) <= b;
    outputs(3118) <= not b;
    outputs(3119) <= a or b;
    outputs(3120) <= b;
    outputs(3121) <= not a;
    outputs(3122) <= a;
    outputs(3123) <= not (a xor b);
    outputs(3124) <= not a;
    outputs(3125) <= not b;
    outputs(3126) <= a and b;
    outputs(3127) <= a and not b;
    outputs(3128) <= not (a xor b);
    outputs(3129) <= a;
    outputs(3130) <= not b;
    outputs(3131) <= not b or a;
    outputs(3132) <= b and not a;
    outputs(3133) <= not a;
    outputs(3134) <= not a;
    outputs(3135) <= a or b;
    outputs(3136) <= a xor b;
    outputs(3137) <= b;
    outputs(3138) <= not b;
    outputs(3139) <= a;
    outputs(3140) <= not a;
    outputs(3141) <= not b;
    outputs(3142) <= not a;
    outputs(3143) <= not (a or b);
    outputs(3144) <= not b;
    outputs(3145) <= not a;
    outputs(3146) <= not a;
    outputs(3147) <= a;
    outputs(3148) <= not (a xor b);
    outputs(3149) <= not a;
    outputs(3150) <= b and not a;
    outputs(3151) <= a and b;
    outputs(3152) <= b and not a;
    outputs(3153) <= a xor b;
    outputs(3154) <= not (a or b);
    outputs(3155) <= not a;
    outputs(3156) <= not a;
    outputs(3157) <= not b;
    outputs(3158) <= not (a or b);
    outputs(3159) <= a;
    outputs(3160) <= a;
    outputs(3161) <= not b;
    outputs(3162) <= not (a xor b);
    outputs(3163) <= not b;
    outputs(3164) <= b and not a;
    outputs(3165) <= a xor b;
    outputs(3166) <= b;
    outputs(3167) <= not a;
    outputs(3168) <= not a;
    outputs(3169) <= a and not b;
    outputs(3170) <= not a or b;
    outputs(3171) <= not a;
    outputs(3172) <= a or b;
    outputs(3173) <= a and b;
    outputs(3174) <= not b;
    outputs(3175) <= not a or b;
    outputs(3176) <= a or b;
    outputs(3177) <= not b;
    outputs(3178) <= a;
    outputs(3179) <= b and not a;
    outputs(3180) <= not b;
    outputs(3181) <= a and b;
    outputs(3182) <= b;
    outputs(3183) <= a and b;
    outputs(3184) <= not (a or b);
    outputs(3185) <= a and b;
    outputs(3186) <= a;
    outputs(3187) <= b;
    outputs(3188) <= a and not b;
    outputs(3189) <= not a;
    outputs(3190) <= not b;
    outputs(3191) <= not b or a;
    outputs(3192) <= not a;
    outputs(3193) <= not b;
    outputs(3194) <= a;
    outputs(3195) <= not (a xor b);
    outputs(3196) <= a and not b;
    outputs(3197) <= not b;
    outputs(3198) <= not a;
    outputs(3199) <= b;
    outputs(3200) <= b and not a;
    outputs(3201) <= not (a or b);
    outputs(3202) <= not b;
    outputs(3203) <= b and not a;
    outputs(3204) <= not (a xor b);
    outputs(3205) <= not b or a;
    outputs(3206) <= not (a or b);
    outputs(3207) <= a and b;
    outputs(3208) <= a and not b;
    outputs(3209) <= b;
    outputs(3210) <= b;
    outputs(3211) <= a;
    outputs(3212) <= a;
    outputs(3213) <= not a;
    outputs(3214) <= not (a or b);
    outputs(3215) <= not b;
    outputs(3216) <= b and not a;
    outputs(3217) <= b;
    outputs(3218) <= not a;
    outputs(3219) <= b;
    outputs(3220) <= b;
    outputs(3221) <= b and not a;
    outputs(3222) <= a or b;
    outputs(3223) <= not a;
    outputs(3224) <= not b or a;
    outputs(3225) <= not b;
    outputs(3226) <= a and not b;
    outputs(3227) <= a xor b;
    outputs(3228) <= a;
    outputs(3229) <= a and b;
    outputs(3230) <= not b or a;
    outputs(3231) <= a;
    outputs(3232) <= not a;
    outputs(3233) <= a and not b;
    outputs(3234) <= not b;
    outputs(3235) <= not (a xor b);
    outputs(3236) <= b;
    outputs(3237) <= not b;
    outputs(3238) <= a and b;
    outputs(3239) <= a and b;
    outputs(3240) <= a;
    outputs(3241) <= not (a xor b);
    outputs(3242) <= b;
    outputs(3243) <= not b or a;
    outputs(3244) <= not (a and b);
    outputs(3245) <= a;
    outputs(3246) <= a and b;
    outputs(3247) <= a;
    outputs(3248) <= a xor b;
    outputs(3249) <= a and not b;
    outputs(3250) <= a and b;
    outputs(3251) <= not (a or b);
    outputs(3252) <= a;
    outputs(3253) <= not b or a;
    outputs(3254) <= not b;
    outputs(3255) <= b and not a;
    outputs(3256) <= not a;
    outputs(3257) <= not b;
    outputs(3258) <= a;
    outputs(3259) <= b;
    outputs(3260) <= not a;
    outputs(3261) <= a and not b;
    outputs(3262) <= a;
    outputs(3263) <= a;
    outputs(3264) <= not b;
    outputs(3265) <= b;
    outputs(3266) <= not b;
    outputs(3267) <= b;
    outputs(3268) <= a;
    outputs(3269) <= a;
    outputs(3270) <= not (a or b);
    outputs(3271) <= b;
    outputs(3272) <= not a;
    outputs(3273) <= a;
    outputs(3274) <= not (a xor b);
    outputs(3275) <= b;
    outputs(3276) <= not a;
    outputs(3277) <= b;
    outputs(3278) <= a and not b;
    outputs(3279) <= a;
    outputs(3280) <= not (a and b);
    outputs(3281) <= not a;
    outputs(3282) <= b;
    outputs(3283) <= b and not a;
    outputs(3284) <= not a;
    outputs(3285) <= not (a or b);
    outputs(3286) <= a and b;
    outputs(3287) <= a and not b;
    outputs(3288) <= not b;
    outputs(3289) <= not a or b;
    outputs(3290) <= a and b;
    outputs(3291) <= not b;
    outputs(3292) <= not b;
    outputs(3293) <= not b;
    outputs(3294) <= a and not b;
    outputs(3295) <= a;
    outputs(3296) <= a and not b;
    outputs(3297) <= not b;
    outputs(3298) <= not a;
    outputs(3299) <= a and b;
    outputs(3300) <= not (a or b);
    outputs(3301) <= not b;
    outputs(3302) <= not (a and b);
    outputs(3303) <= b;
    outputs(3304) <= b;
    outputs(3305) <= not a;
    outputs(3306) <= b;
    outputs(3307) <= not (a or b);
    outputs(3308) <= a;
    outputs(3309) <= b and not a;
    outputs(3310) <= b and not a;
    outputs(3311) <= b;
    outputs(3312) <= b;
    outputs(3313) <= not a;
    outputs(3314) <= b and not a;
    outputs(3315) <= a;
    outputs(3316) <= a;
    outputs(3317) <= a;
    outputs(3318) <= a;
    outputs(3319) <= a and not b;
    outputs(3320) <= b and not a;
    outputs(3321) <= a or b;
    outputs(3322) <= a;
    outputs(3323) <= b and not a;
    outputs(3324) <= b and not a;
    outputs(3325) <= not (a or b);
    outputs(3326) <= not b or a;
    outputs(3327) <= a xor b;
    outputs(3328) <= not (a or b);
    outputs(3329) <= a or b;
    outputs(3330) <= b;
    outputs(3331) <= a;
    outputs(3332) <= not (a or b);
    outputs(3333) <= a and not b;
    outputs(3334) <= a;
    outputs(3335) <= a xor b;
    outputs(3336) <= not b;
    outputs(3337) <= not (a xor b);
    outputs(3338) <= b;
    outputs(3339) <= a xor b;
    outputs(3340) <= b;
    outputs(3341) <= a and not b;
    outputs(3342) <= not a;
    outputs(3343) <= not a or b;
    outputs(3344) <= not (a xor b);
    outputs(3345) <= not a;
    outputs(3346) <= b;
    outputs(3347) <= a;
    outputs(3348) <= not b;
    outputs(3349) <= a and not b;
    outputs(3350) <= a or b;
    outputs(3351) <= a and b;
    outputs(3352) <= not a;
    outputs(3353) <= not a or b;
    outputs(3354) <= not a;
    outputs(3355) <= b;
    outputs(3356) <= not (a or b);
    outputs(3357) <= not b or a;
    outputs(3358) <= a and b;
    outputs(3359) <= a and b;
    outputs(3360) <= b and not a;
    outputs(3361) <= a and b;
    outputs(3362) <= a and not b;
    outputs(3363) <= not (a and b);
    outputs(3364) <= a;
    outputs(3365) <= a or b;
    outputs(3366) <= a;
    outputs(3367) <= a;
    outputs(3368) <= a xor b;
    outputs(3369) <= a and not b;
    outputs(3370) <= a;
    outputs(3371) <= not (a xor b);
    outputs(3372) <= not a;
    outputs(3373) <= not b;
    outputs(3374) <= a;
    outputs(3375) <= b;
    outputs(3376) <= a xor b;
    outputs(3377) <= not a;
    outputs(3378) <= not b;
    outputs(3379) <= a;
    outputs(3380) <= a;
    outputs(3381) <= a or b;
    outputs(3382) <= a;
    outputs(3383) <= not b;
    outputs(3384) <= not b;
    outputs(3385) <= b;
    outputs(3386) <= not (a or b);
    outputs(3387) <= a or b;
    outputs(3388) <= not (a or b);
    outputs(3389) <= not b;
    outputs(3390) <= not a;
    outputs(3391) <= b;
    outputs(3392) <= not b;
    outputs(3393) <= not b;
    outputs(3394) <= a xor b;
    outputs(3395) <= a;
    outputs(3396) <= a xor b;
    outputs(3397) <= not b;
    outputs(3398) <= a;
    outputs(3399) <= not a;
    outputs(3400) <= not b or a;
    outputs(3401) <= a and not b;
    outputs(3402) <= a;
    outputs(3403) <= a and b;
    outputs(3404) <= b;
    outputs(3405) <= b;
    outputs(3406) <= not b;
    outputs(3407) <= not (a xor b);
    outputs(3408) <= not b or a;
    outputs(3409) <= not (a or b);
    outputs(3410) <= not a;
    outputs(3411) <= not a;
    outputs(3412) <= not (a or b);
    outputs(3413) <= not b;
    outputs(3414) <= not (a or b);
    outputs(3415) <= b;
    outputs(3416) <= b;
    outputs(3417) <= not b;
    outputs(3418) <= a;
    outputs(3419) <= b;
    outputs(3420) <= not b;
    outputs(3421) <= b;
    outputs(3422) <= a or b;
    outputs(3423) <= b;
    outputs(3424) <= not (a or b);
    outputs(3425) <= a and not b;
    outputs(3426) <= not (a or b);
    outputs(3427) <= b;
    outputs(3428) <= a xor b;
    outputs(3429) <= not b or a;
    outputs(3430) <= not a;
    outputs(3431) <= a;
    outputs(3432) <= a and not b;
    outputs(3433) <= a xor b;
    outputs(3434) <= a;
    outputs(3435) <= not (a or b);
    outputs(3436) <= not (a or b);
    outputs(3437) <= not (a xor b);
    outputs(3438) <= b;
    outputs(3439) <= a xor b;
    outputs(3440) <= not a or b;
    outputs(3441) <= a and not b;
    outputs(3442) <= a and not b;
    outputs(3443) <= b;
    outputs(3444) <= b;
    outputs(3445) <= b;
    outputs(3446) <= a;
    outputs(3447) <= a xor b;
    outputs(3448) <= b and not a;
    outputs(3449) <= not (a or b);
    outputs(3450) <= not (a xor b);
    outputs(3451) <= not (a xor b);
    outputs(3452) <= a and not b;
    outputs(3453) <= not b or a;
    outputs(3454) <= not (a xor b);
    outputs(3455) <= not (a xor b);
    outputs(3456) <= b;
    outputs(3457) <= a and b;
    outputs(3458) <= not (a and b);
    outputs(3459) <= a or b;
    outputs(3460) <= a xor b;
    outputs(3461) <= a xor b;
    outputs(3462) <= not (a or b);
    outputs(3463) <= b;
    outputs(3464) <= a and not b;
    outputs(3465) <= a and b;
    outputs(3466) <= not (a or b);
    outputs(3467) <= not (a or b);
    outputs(3468) <= a and b;
    outputs(3469) <= a;
    outputs(3470) <= not b;
    outputs(3471) <= not a;
    outputs(3472) <= not (a and b);
    outputs(3473) <= a and not b;
    outputs(3474) <= not a or b;
    outputs(3475) <= a and b;
    outputs(3476) <= not a;
    outputs(3477) <= not b;
    outputs(3478) <= not b;
    outputs(3479) <= not (a and b);
    outputs(3480) <= a and not b;
    outputs(3481) <= not a;
    outputs(3482) <= not (a or b);
    outputs(3483) <= b and not a;
    outputs(3484) <= a and not b;
    outputs(3485) <= not a;
    outputs(3486) <= not (a or b);
    outputs(3487) <= a and not b;
    outputs(3488) <= a;
    outputs(3489) <= not a or b;
    outputs(3490) <= b;
    outputs(3491) <= b and not a;
    outputs(3492) <= a;
    outputs(3493) <= not (a and b);
    outputs(3494) <= not (a or b);
    outputs(3495) <= not a;
    outputs(3496) <= not a;
    outputs(3497) <= not a or b;
    outputs(3498) <= not b;
    outputs(3499) <= not (a or b);
    outputs(3500) <= a;
    outputs(3501) <= a and b;
    outputs(3502) <= b and not a;
    outputs(3503) <= not a or b;
    outputs(3504) <= b;
    outputs(3505) <= b and not a;
    outputs(3506) <= not (a or b);
    outputs(3507) <= not b;
    outputs(3508) <= not b;
    outputs(3509) <= not (a xor b);
    outputs(3510) <= b and not a;
    outputs(3511) <= a;
    outputs(3512) <= a and not b;
    outputs(3513) <= not a;
    outputs(3514) <= not (a and b);
    outputs(3515) <= a and b;
    outputs(3516) <= not (a and b);
    outputs(3517) <= not b;
    outputs(3518) <= not a;
    outputs(3519) <= a and b;
    outputs(3520) <= b;
    outputs(3521) <= not (a or b);
    outputs(3522) <= b;
    outputs(3523) <= not b;
    outputs(3524) <= b;
    outputs(3525) <= a;
    outputs(3526) <= not (a xor b);
    outputs(3527) <= a;
    outputs(3528) <= b and not a;
    outputs(3529) <= not a;
    outputs(3530) <= b;
    outputs(3531) <= not (a or b);
    outputs(3532) <= not b;
    outputs(3533) <= not b or a;
    outputs(3534) <= b and not a;
    outputs(3535) <= not b;
    outputs(3536) <= not (a or b);
    outputs(3537) <= a;
    outputs(3538) <= b;
    outputs(3539) <= b;
    outputs(3540) <= a;
    outputs(3541) <= not b;
    outputs(3542) <= not a;
    outputs(3543) <= not b or a;
    outputs(3544) <= a;
    outputs(3545) <= a xor b;
    outputs(3546) <= b;
    outputs(3547) <= a xor b;
    outputs(3548) <= not a or b;
    outputs(3549) <= a or b;
    outputs(3550) <= not a;
    outputs(3551) <= b and not a;
    outputs(3552) <= not (a or b);
    outputs(3553) <= not a;
    outputs(3554) <= a and not b;
    outputs(3555) <= b;
    outputs(3556) <= b;
    outputs(3557) <= a and b;
    outputs(3558) <= not b or a;
    outputs(3559) <= a;
    outputs(3560) <= b;
    outputs(3561) <= not (a or b);
    outputs(3562) <= not a;
    outputs(3563) <= not (a xor b);
    outputs(3564) <= not b;
    outputs(3565) <= a and not b;
    outputs(3566) <= not (a or b);
    outputs(3567) <= a;
    outputs(3568) <= not a;
    outputs(3569) <= not a;
    outputs(3570) <= not (a or b);
    outputs(3571) <= not a;
    outputs(3572) <= a and b;
    outputs(3573) <= not (a xor b);
    outputs(3574) <= b;
    outputs(3575) <= b and not a;
    outputs(3576) <= b;
    outputs(3577) <= b and not a;
    outputs(3578) <= a and b;
    outputs(3579) <= a and not b;
    outputs(3580) <= a and b;
    outputs(3581) <= not b;
    outputs(3582) <= a and not b;
    outputs(3583) <= a and b;
    outputs(3584) <= a xor b;
    outputs(3585) <= b and not a;
    outputs(3586) <= not a;
    outputs(3587) <= b;
    outputs(3588) <= a;
    outputs(3589) <= a and b;
    outputs(3590) <= a and not b;
    outputs(3591) <= not a;
    outputs(3592) <= a or b;
    outputs(3593) <= a and not b;
    outputs(3594) <= b and not a;
    outputs(3595) <= b;
    outputs(3596) <= a and b;
    outputs(3597) <= b;
    outputs(3598) <= not (a or b);
    outputs(3599) <= b and not a;
    outputs(3600) <= not (a or b);
    outputs(3601) <= not (a or b);
    outputs(3602) <= a xor b;
    outputs(3603) <= not (a xor b);
    outputs(3604) <= a xor b;
    outputs(3605) <= a and not b;
    outputs(3606) <= not a;
    outputs(3607) <= b;
    outputs(3608) <= not b;
    outputs(3609) <= a and b;
    outputs(3610) <= not (a or b);
    outputs(3611) <= not b or a;
    outputs(3612) <= a and b;
    outputs(3613) <= a and b;
    outputs(3614) <= a or b;
    outputs(3615) <= not b;
    outputs(3616) <= a and not b;
    outputs(3617) <= b;
    outputs(3618) <= b and not a;
    outputs(3619) <= not b;
    outputs(3620) <= not a;
    outputs(3621) <= not b;
    outputs(3622) <= a and not b;
    outputs(3623) <= not (a or b);
    outputs(3624) <= b and not a;
    outputs(3625) <= not (a xor b);
    outputs(3626) <= a and b;
    outputs(3627) <= not (a or b);
    outputs(3628) <= a and b;
    outputs(3629) <= a;
    outputs(3630) <= a;
    outputs(3631) <= a xor b;
    outputs(3632) <= a xor b;
    outputs(3633) <= a xor b;
    outputs(3634) <= not a;
    outputs(3635) <= a and b;
    outputs(3636) <= b and not a;
    outputs(3637) <= not b or a;
    outputs(3638) <= not a;
    outputs(3639) <= b and not a;
    outputs(3640) <= b;
    outputs(3641) <= not b;
    outputs(3642) <= a;
    outputs(3643) <= a;
    outputs(3644) <= b and not a;
    outputs(3645) <= not a;
    outputs(3646) <= a and not b;
    outputs(3647) <= a or b;
    outputs(3648) <= a and b;
    outputs(3649) <= not a;
    outputs(3650) <= not b;
    outputs(3651) <= a and not b;
    outputs(3652) <= a and b;
    outputs(3653) <= not a or b;
    outputs(3654) <= not (a xor b);
    outputs(3655) <= a;
    outputs(3656) <= not a;
    outputs(3657) <= not (a xor b);
    outputs(3658) <= not a or b;
    outputs(3659) <= a and not b;
    outputs(3660) <= a and b;
    outputs(3661) <= a;
    outputs(3662) <= a;
    outputs(3663) <= a and b;
    outputs(3664) <= a or b;
    outputs(3665) <= a;
    outputs(3666) <= b and not a;
    outputs(3667) <= a and b;
    outputs(3668) <= a;
    outputs(3669) <= not b or a;
    outputs(3670) <= not a or b;
    outputs(3671) <= not a;
    outputs(3672) <= a xor b;
    outputs(3673) <= not b;
    outputs(3674) <= a xor b;
    outputs(3675) <= b and not a;
    outputs(3676) <= b and not a;
    outputs(3677) <= not a;
    outputs(3678) <= not b;
    outputs(3679) <= a or b;
    outputs(3680) <= not a;
    outputs(3681) <= not a;
    outputs(3682) <= not (a or b);
    outputs(3683) <= not b;
    outputs(3684) <= a;
    outputs(3685) <= a;
    outputs(3686) <= a xor b;
    outputs(3687) <= b;
    outputs(3688) <= not (a or b);
    outputs(3689) <= a and b;
    outputs(3690) <= b and not a;
    outputs(3691) <= a and b;
    outputs(3692) <= b and not a;
    outputs(3693) <= b;
    outputs(3694) <= a and not b;
    outputs(3695) <= b;
    outputs(3696) <= not a or b;
    outputs(3697) <= a xor b;
    outputs(3698) <= a and b;
    outputs(3699) <= not (a or b);
    outputs(3700) <= not b or a;
    outputs(3701) <= not b;
    outputs(3702) <= a and not b;
    outputs(3703) <= a and b;
    outputs(3704) <= not (a xor b);
    outputs(3705) <= a and b;
    outputs(3706) <= a and b;
    outputs(3707) <= not b;
    outputs(3708) <= not (a xor b);
    outputs(3709) <= not (a or b);
    outputs(3710) <= not (a xor b);
    outputs(3711) <= b;
    outputs(3712) <= not a;
    outputs(3713) <= not (a or b);
    outputs(3714) <= a and b;
    outputs(3715) <= a and not b;
    outputs(3716) <= a;
    outputs(3717) <= not (a or b);
    outputs(3718) <= not (a or b);
    outputs(3719) <= not b;
    outputs(3720) <= a and not b;
    outputs(3721) <= a xor b;
    outputs(3722) <= a and not b;
    outputs(3723) <= a xor b;
    outputs(3724) <= a and not b;
    outputs(3725) <= not (a or b);
    outputs(3726) <= a;
    outputs(3727) <= b;
    outputs(3728) <= not a or b;
    outputs(3729) <= a and not b;
    outputs(3730) <= not (a or b);
    outputs(3731) <= not (a and b);
    outputs(3732) <= not (a and b);
    outputs(3733) <= a or b;
    outputs(3734) <= not (a or b);
    outputs(3735) <= a xor b;
    outputs(3736) <= not b;
    outputs(3737) <= not (a and b);
    outputs(3738) <= not (a and b);
    outputs(3739) <= a and b;
    outputs(3740) <= a;
    outputs(3741) <= not (a xor b);
    outputs(3742) <= b;
    outputs(3743) <= b and not a;
    outputs(3744) <= not (a or b);
    outputs(3745) <= a and b;
    outputs(3746) <= not b;
    outputs(3747) <= a and not b;
    outputs(3748) <= b and not a;
    outputs(3749) <= not b or a;
    outputs(3750) <= not b;
    outputs(3751) <= not (a or b);
    outputs(3752) <= b and not a;
    outputs(3753) <= a xor b;
    outputs(3754) <= not a;
    outputs(3755) <= b;
    outputs(3756) <= a and b;
    outputs(3757) <= not (a or b);
    outputs(3758) <= a and b;
    outputs(3759) <= not (a xor b);
    outputs(3760) <= not a;
    outputs(3761) <= not a;
    outputs(3762) <= b and not a;
    outputs(3763) <= not (a xor b);
    outputs(3764) <= b;
    outputs(3765) <= not b;
    outputs(3766) <= a;
    outputs(3767) <= not (a or b);
    outputs(3768) <= not (a and b);
    outputs(3769) <= not b;
    outputs(3770) <= b;
    outputs(3771) <= a and b;
    outputs(3772) <= a and not b;
    outputs(3773) <= not a;
    outputs(3774) <= b and not a;
    outputs(3775) <= not a;
    outputs(3776) <= not a;
    outputs(3777) <= a and b;
    outputs(3778) <= not (a xor b);
    outputs(3779) <= not (a or b);
    outputs(3780) <= b and not a;
    outputs(3781) <= not b;
    outputs(3782) <= not (a or b);
    outputs(3783) <= not (a or b);
    outputs(3784) <= b;
    outputs(3785) <= b and not a;
    outputs(3786) <= b and not a;
    outputs(3787) <= not a;
    outputs(3788) <= not (a xor b);
    outputs(3789) <= a xor b;
    outputs(3790) <= b;
    outputs(3791) <= not a or b;
    outputs(3792) <= not a;
    outputs(3793) <= a and not b;
    outputs(3794) <= not b;
    outputs(3795) <= b;
    outputs(3796) <= a xor b;
    outputs(3797) <= not a;
    outputs(3798) <= b and not a;
    outputs(3799) <= b;
    outputs(3800) <= b;
    outputs(3801) <= a xor b;
    outputs(3802) <= b;
    outputs(3803) <= not a or b;
    outputs(3804) <= not a;
    outputs(3805) <= a or b;
    outputs(3806) <= not a;
    outputs(3807) <= not b;
    outputs(3808) <= a;
    outputs(3809) <= b;
    outputs(3810) <= b;
    outputs(3811) <= not a;
    outputs(3812) <= not a;
    outputs(3813) <= a and b;
    outputs(3814) <= not (a or b);
    outputs(3815) <= not a;
    outputs(3816) <= not (a or b);
    outputs(3817) <= not a;
    outputs(3818) <= a;
    outputs(3819) <= a;
    outputs(3820) <= not b;
    outputs(3821) <= not (a or b);
    outputs(3822) <= b and not a;
    outputs(3823) <= not (a and b);
    outputs(3824) <= a and b;
    outputs(3825) <= not (a or b);
    outputs(3826) <= not (a xor b);
    outputs(3827) <= a and not b;
    outputs(3828) <= not b;
    outputs(3829) <= b;
    outputs(3830) <= not (a xor b);
    outputs(3831) <= not a;
    outputs(3832) <= b and not a;
    outputs(3833) <= a;
    outputs(3834) <= a;
    outputs(3835) <= a and not b;
    outputs(3836) <= a and not b;
    outputs(3837) <= a and not b;
    outputs(3838) <= a and b;
    outputs(3839) <= a and b;
    outputs(3840) <= b and not a;
    outputs(3841) <= b;
    outputs(3842) <= not (a and b);
    outputs(3843) <= not (a or b);
    outputs(3844) <= a or b;
    outputs(3845) <= b;
    outputs(3846) <= a xor b;
    outputs(3847) <= not a;
    outputs(3848) <= not b;
    outputs(3849) <= not b;
    outputs(3850) <= not b;
    outputs(3851) <= b and not a;
    outputs(3852) <= a;
    outputs(3853) <= a xor b;
    outputs(3854) <= not a;
    outputs(3855) <= not a;
    outputs(3856) <= not a;
    outputs(3857) <= a and b;
    outputs(3858) <= a and not b;
    outputs(3859) <= not (a or b);
    outputs(3860) <= b;
    outputs(3861) <= not (a or b);
    outputs(3862) <= a and not b;
    outputs(3863) <= b;
    outputs(3864) <= a;
    outputs(3865) <= a and not b;
    outputs(3866) <= b;
    outputs(3867) <= a;
    outputs(3868) <= b and not a;
    outputs(3869) <= not (a and b);
    outputs(3870) <= b;
    outputs(3871) <= not a;
    outputs(3872) <= not (a xor b);
    outputs(3873) <= b;
    outputs(3874) <= not (a or b);
    outputs(3875) <= not b or a;
    outputs(3876) <= a;
    outputs(3877) <= a and not b;
    outputs(3878) <= not a;
    outputs(3879) <= not b;
    outputs(3880) <= not b;
    outputs(3881) <= not (a and b);
    outputs(3882) <= a and b;
    outputs(3883) <= not (a xor b);
    outputs(3884) <= not a;
    outputs(3885) <= not a;
    outputs(3886) <= b;
    outputs(3887) <= not b or a;
    outputs(3888) <= a and b;
    outputs(3889) <= not (a or b);
    outputs(3890) <= a;
    outputs(3891) <= a and b;
    outputs(3892) <= a and b;
    outputs(3893) <= not b;
    outputs(3894) <= b;
    outputs(3895) <= not (a or b);
    outputs(3896) <= b;
    outputs(3897) <= not (a or b);
    outputs(3898) <= not (a or b);
    outputs(3899) <= not (a or b);
    outputs(3900) <= not b;
    outputs(3901) <= not (a and b);
    outputs(3902) <= not (a or b);
    outputs(3903) <= a;
    outputs(3904) <= a and not b;
    outputs(3905) <= a;
    outputs(3906) <= not (a xor b);
    outputs(3907) <= b;
    outputs(3908) <= b and not a;
    outputs(3909) <= a and b;
    outputs(3910) <= a;
    outputs(3911) <= b;
    outputs(3912) <= a or b;
    outputs(3913) <= b and not a;
    outputs(3914) <= a;
    outputs(3915) <= not a or b;
    outputs(3916) <= not (a or b);
    outputs(3917) <= not a;
    outputs(3918) <= not (a or b);
    outputs(3919) <= not a;
    outputs(3920) <= not (a or b);
    outputs(3921) <= b;
    outputs(3922) <= not b;
    outputs(3923) <= a and not b;
    outputs(3924) <= not b or a;
    outputs(3925) <= a and not b;
    outputs(3926) <= a and b;
    outputs(3927) <= not b or a;
    outputs(3928) <= not (a or b);
    outputs(3929) <= not a;
    outputs(3930) <= b;
    outputs(3931) <= not a;
    outputs(3932) <= a;
    outputs(3933) <= a and not b;
    outputs(3934) <= b and not a;
    outputs(3935) <= a;
    outputs(3936) <= b;
    outputs(3937) <= not (a xor b);
    outputs(3938) <= a and b;
    outputs(3939) <= a or b;
    outputs(3940) <= b;
    outputs(3941) <= a and b;
    outputs(3942) <= b;
    outputs(3943) <= b;
    outputs(3944) <= not (a or b);
    outputs(3945) <= not (a xor b);
    outputs(3946) <= b and not a;
    outputs(3947) <= a xor b;
    outputs(3948) <= not b;
    outputs(3949) <= not b or a;
    outputs(3950) <= a;
    outputs(3951) <= not (a xor b);
    outputs(3952) <= a and b;
    outputs(3953) <= b and not a;
    outputs(3954) <= not (a or b);
    outputs(3955) <= a;
    outputs(3956) <= b and not a;
    outputs(3957) <= a and not b;
    outputs(3958) <= not a;
    outputs(3959) <= b;
    outputs(3960) <= a;
    outputs(3961) <= not (a or b);
    outputs(3962) <= not b;
    outputs(3963) <= not a;
    outputs(3964) <= b;
    outputs(3965) <= not a;
    outputs(3966) <= a;
    outputs(3967) <= not b;
    outputs(3968) <= a and not b;
    outputs(3969) <= a and b;
    outputs(3970) <= not b;
    outputs(3971) <= b and not a;
    outputs(3972) <= not (a or b);
    outputs(3973) <= b;
    outputs(3974) <= b and not a;
    outputs(3975) <= not b;
    outputs(3976) <= not a;
    outputs(3977) <= b;
    outputs(3978) <= b;
    outputs(3979) <= a and not b;
    outputs(3980) <= b and not a;
    outputs(3981) <= not a or b;
    outputs(3982) <= a or b;
    outputs(3983) <= not (a or b);
    outputs(3984) <= not b;
    outputs(3985) <= a;
    outputs(3986) <= b;
    outputs(3987) <= a and not b;
    outputs(3988) <= not (a or b);
    outputs(3989) <= b;
    outputs(3990) <= a;
    outputs(3991) <= not a;
    outputs(3992) <= a and b;
    outputs(3993) <= b and not a;
    outputs(3994) <= not b;
    outputs(3995) <= b;
    outputs(3996) <= not a;
    outputs(3997) <= not a;
    outputs(3998) <= b;
    outputs(3999) <= a;
    outputs(4000) <= not a or b;
    outputs(4001) <= not b or a;
    outputs(4002) <= not (a or b);
    outputs(4003) <= a and not b;
    outputs(4004) <= not a;
    outputs(4005) <= not (a or b);
    outputs(4006) <= a and b;
    outputs(4007) <= not a;
    outputs(4008) <= b and not a;
    outputs(4009) <= b and not a;
    outputs(4010) <= b and not a;
    outputs(4011) <= not b;
    outputs(4012) <= not (a or b);
    outputs(4013) <= not a;
    outputs(4014) <= not b;
    outputs(4015) <= not a;
    outputs(4016) <= not b;
    outputs(4017) <= a;
    outputs(4018) <= a;
    outputs(4019) <= a and b;
    outputs(4020) <= a and not b;
    outputs(4021) <= a and not b;
    outputs(4022) <= not b or a;
    outputs(4023) <= not a or b;
    outputs(4024) <= not b;
    outputs(4025) <= a and b;
    outputs(4026) <= b and not a;
    outputs(4027) <= b;
    outputs(4028) <= not a;
    outputs(4029) <= a;
    outputs(4030) <= not b or a;
    outputs(4031) <= a;
    outputs(4032) <= b;
    outputs(4033) <= a;
    outputs(4034) <= a and not b;
    outputs(4035) <= b;
    outputs(4036) <= not (a xor b);
    outputs(4037) <= b;
    outputs(4038) <= a and b;
    outputs(4039) <= not b;
    outputs(4040) <= a;
    outputs(4041) <= not b;
    outputs(4042) <= b and not a;
    outputs(4043) <= b and not a;
    outputs(4044) <= not b;
    outputs(4045) <= not (a or b);
    outputs(4046) <= a xor b;
    outputs(4047) <= a;
    outputs(4048) <= a and b;
    outputs(4049) <= not (a and b);
    outputs(4050) <= a;
    outputs(4051) <= not (a or b);
    outputs(4052) <= a;
    outputs(4053) <= b and not a;
    outputs(4054) <= a;
    outputs(4055) <= a;
    outputs(4056) <= not (a or b);
    outputs(4057) <= not a;
    outputs(4058) <= not b;
    outputs(4059) <= a and b;
    outputs(4060) <= not b;
    outputs(4061) <= b and not a;
    outputs(4062) <= not b;
    outputs(4063) <= a and b;
    outputs(4064) <= a;
    outputs(4065) <= b and not a;
    outputs(4066) <= not b;
    outputs(4067) <= b;
    outputs(4068) <= a;
    outputs(4069) <= b;
    outputs(4070) <= not b;
    outputs(4071) <= a and not b;
    outputs(4072) <= a and b;
    outputs(4073) <= b and not a;
    outputs(4074) <= b;
    outputs(4075) <= b and not a;
    outputs(4076) <= not b;
    outputs(4077) <= not a or b;
    outputs(4078) <= not b or a;
    outputs(4079) <= not (a xor b);
    outputs(4080) <= not b or a;
    outputs(4081) <= a;
    outputs(4082) <= not (a xor b);
    outputs(4083) <= not (a or b);
    outputs(4084) <= b;
    outputs(4085) <= b and not a;
    outputs(4086) <= b and not a;
    outputs(4087) <= a xor b;
    outputs(4088) <= not a;
    outputs(4089) <= a;
    outputs(4090) <= a;
    outputs(4091) <= a and b;
    outputs(4092) <= a;
    outputs(4093) <= not a;
    outputs(4094) <= a;
    outputs(4095) <= a and b;
    outputs(4096) <= a or b;
    outputs(4097) <= a;
    outputs(4098) <= a;
    outputs(4099) <= not b or a;
    outputs(4100) <= a or b;
    outputs(4101) <= not a or b;
    outputs(4102) <= a;
    outputs(4103) <= not b;
    outputs(4104) <= a;
    outputs(4105) <= a;
    outputs(4106) <= not b;
    outputs(4107) <= not b;
    outputs(4108) <= not b or a;
    outputs(4109) <= a;
    outputs(4110) <= b;
    outputs(4111) <= not (a or b);
    outputs(4112) <= not (a or b);
    outputs(4113) <= a xor b;
    outputs(4114) <= not a;
    outputs(4115) <= not (a xor b);
    outputs(4116) <= a or b;
    outputs(4117) <= not (a xor b);
    outputs(4118) <= a and not b;
    outputs(4119) <= b;
    outputs(4120) <= a xor b;
    outputs(4121) <= a xor b;
    outputs(4122) <= not b or a;
    outputs(4123) <= a and not b;
    outputs(4124) <= b;
    outputs(4125) <= b and not a;
    outputs(4126) <= not a;
    outputs(4127) <= not b;
    outputs(4128) <= a xor b;
    outputs(4129) <= a and not b;
    outputs(4130) <= a xor b;
    outputs(4131) <= not a;
    outputs(4132) <= a or b;
    outputs(4133) <= not b;
    outputs(4134) <= not a or b;
    outputs(4135) <= a xor b;
    outputs(4136) <= not b;
    outputs(4137) <= a xor b;
    outputs(4138) <= a;
    outputs(4139) <= a or b;
    outputs(4140) <= a and b;
    outputs(4141) <= a xor b;
    outputs(4142) <= not a;
    outputs(4143) <= not b;
    outputs(4144) <= a and not b;
    outputs(4145) <= not b or a;
    outputs(4146) <= a;
    outputs(4147) <= a;
    outputs(4148) <= b;
    outputs(4149) <= not b;
    outputs(4150) <= not b;
    outputs(4151) <= a;
    outputs(4152) <= a or b;
    outputs(4153) <= a;
    outputs(4154) <= b;
    outputs(4155) <= not (a and b);
    outputs(4156) <= a and not b;
    outputs(4157) <= b;
    outputs(4158) <= not b;
    outputs(4159) <= a;
    outputs(4160) <= not a;
    outputs(4161) <= a and not b;
    outputs(4162) <= b;
    outputs(4163) <= not b or a;
    outputs(4164) <= not a;
    outputs(4165) <= not (a xor b);
    outputs(4166) <= not (a xor b);
    outputs(4167) <= not (a and b);
    outputs(4168) <= a xor b;
    outputs(4169) <= not b;
    outputs(4170) <= a;
    outputs(4171) <= a;
    outputs(4172) <= b;
    outputs(4173) <= a and not b;
    outputs(4174) <= not (a xor b);
    outputs(4175) <= not (a or b);
    outputs(4176) <= a;
    outputs(4177) <= a xor b;
    outputs(4178) <= a;
    outputs(4179) <= not a;
    outputs(4180) <= a and not b;
    outputs(4181) <= b;
    outputs(4182) <= b and not a;
    outputs(4183) <= not (a or b);
    outputs(4184) <= not a or b;
    outputs(4185) <= a xor b;
    outputs(4186) <= a or b;
    outputs(4187) <= not b;
    outputs(4188) <= a and b;
    outputs(4189) <= b;
    outputs(4190) <= a and not b;
    outputs(4191) <= a;
    outputs(4192) <= not (a xor b);
    outputs(4193) <= b and not a;
    outputs(4194) <= not b or a;
    outputs(4195) <= a xor b;
    outputs(4196) <= a;
    outputs(4197) <= not (a xor b);
    outputs(4198) <= a and not b;
    outputs(4199) <= a and not b;
    outputs(4200) <= b;
    outputs(4201) <= a and not b;
    outputs(4202) <= not (a xor b);
    outputs(4203) <= not (a or b);
    outputs(4204) <= not a;
    outputs(4205) <= a or b;
    outputs(4206) <= not (a or b);
    outputs(4207) <= not a;
    outputs(4208) <= not a;
    outputs(4209) <= not b or a;
    outputs(4210) <= not a or b;
    outputs(4211) <= b;
    outputs(4212) <= not a;
    outputs(4213) <= not a;
    outputs(4214) <= not a;
    outputs(4215) <= b;
    outputs(4216) <= a or b;
    outputs(4217) <= a or b;
    outputs(4218) <= b and not a;
    outputs(4219) <= b;
    outputs(4220) <= not (a and b);
    outputs(4221) <= b;
    outputs(4222) <= a and not b;
    outputs(4223) <= not (a xor b);
    outputs(4224) <= b;
    outputs(4225) <= a;
    outputs(4226) <= a and b;
    outputs(4227) <= a and not b;
    outputs(4228) <= not b or a;
    outputs(4229) <= a and b;
    outputs(4230) <= not (a xor b);
    outputs(4231) <= not a or b;
    outputs(4232) <= b;
    outputs(4233) <= b;
    outputs(4234) <= not (a xor b);
    outputs(4235) <= a and b;
    outputs(4236) <= not a;
    outputs(4237) <= a;
    outputs(4238) <= a;
    outputs(4239) <= b;
    outputs(4240) <= a or b;
    outputs(4241) <= not (a and b);
    outputs(4242) <= not b;
    outputs(4243) <= a and not b;
    outputs(4244) <= a and b;
    outputs(4245) <= a;
    outputs(4246) <= a;
    outputs(4247) <= not b;
    outputs(4248) <= not b or a;
    outputs(4249) <= a xor b;
    outputs(4250) <= not b;
    outputs(4251) <= a xor b;
    outputs(4252) <= a xor b;
    outputs(4253) <= not (a xor b);
    outputs(4254) <= not (a and b);
    outputs(4255) <= not b or a;
    outputs(4256) <= a or b;
    outputs(4257) <= a;
    outputs(4258) <= not a;
    outputs(4259) <= b;
    outputs(4260) <= not (a and b);
    outputs(4261) <= b and not a;
    outputs(4262) <= a and b;
    outputs(4263) <= not (a or b);
    outputs(4264) <= a xor b;
    outputs(4265) <= not b;
    outputs(4266) <= a;
    outputs(4267) <= b;
    outputs(4268) <= b;
    outputs(4269) <= not b or a;
    outputs(4270) <= not a;
    outputs(4271) <= not (a xor b);
    outputs(4272) <= not a;
    outputs(4273) <= a;
    outputs(4274) <= a or b;
    outputs(4275) <= a xor b;
    outputs(4276) <= b;
    outputs(4277) <= not b or a;
    outputs(4278) <= not a;
    outputs(4279) <= a xor b;
    outputs(4280) <= a xor b;
    outputs(4281) <= b;
    outputs(4282) <= not (a and b);
    outputs(4283) <= a and b;
    outputs(4284) <= not a or b;
    outputs(4285) <= a and not b;
    outputs(4286) <= not (a or b);
    outputs(4287) <= not (a xor b);
    outputs(4288) <= b and not a;
    outputs(4289) <= a and b;
    outputs(4290) <= not (a xor b);
    outputs(4291) <= a;
    outputs(4292) <= b;
    outputs(4293) <= a xor b;
    outputs(4294) <= a;
    outputs(4295) <= not b or a;
    outputs(4296) <= b;
    outputs(4297) <= not a;
    outputs(4298) <= not a;
    outputs(4299) <= b;
    outputs(4300) <= not b or a;
    outputs(4301) <= a;
    outputs(4302) <= b;
    outputs(4303) <= not b;
    outputs(4304) <= a;
    outputs(4305) <= a or b;
    outputs(4306) <= a xor b;
    outputs(4307) <= not a;
    outputs(4308) <= b;
    outputs(4309) <= not b;
    outputs(4310) <= not a;
    outputs(4311) <= not b;
    outputs(4312) <= not b;
    outputs(4313) <= not a or b;
    outputs(4314) <= b;
    outputs(4315) <= not a;
    outputs(4316) <= a or b;
    outputs(4317) <= not a;
    outputs(4318) <= not a;
    outputs(4319) <= not b;
    outputs(4320) <= not (a and b);
    outputs(4321) <= b and not a;
    outputs(4322) <= a xor b;
    outputs(4323) <= a xor b;
    outputs(4324) <= a and b;
    outputs(4325) <= b and not a;
    outputs(4326) <= a xor b;
    outputs(4327) <= b;
    outputs(4328) <= a xor b;
    outputs(4329) <= a;
    outputs(4330) <= a xor b;
    outputs(4331) <= a and b;
    outputs(4332) <= b;
    outputs(4333) <= not (a xor b);
    outputs(4334) <= not b;
    outputs(4335) <= not a;
    outputs(4336) <= not (a or b);
    outputs(4337) <= not (a or b);
    outputs(4338) <= not b;
    outputs(4339) <= not a;
    outputs(4340) <= not (a or b);
    outputs(4341) <= not (a xor b);
    outputs(4342) <= b;
    outputs(4343) <= not a or b;
    outputs(4344) <= not (a xor b);
    outputs(4345) <= b;
    outputs(4346) <= not (a or b);
    outputs(4347) <= a and b;
    outputs(4348) <= a or b;
    outputs(4349) <= a or b;
    outputs(4350) <= b;
    outputs(4351) <= a;
    outputs(4352) <= not a or b;
    outputs(4353) <= not b;
    outputs(4354) <= a xor b;
    outputs(4355) <= not b;
    outputs(4356) <= not (a or b);
    outputs(4357) <= a and not b;
    outputs(4358) <= b and not a;
    outputs(4359) <= not a;
    outputs(4360) <= not (a and b);
    outputs(4361) <= not a;
    outputs(4362) <= b;
    outputs(4363) <= a;
    outputs(4364) <= b;
    outputs(4365) <= not a;
    outputs(4366) <= not (a xor b);
    outputs(4367) <= b;
    outputs(4368) <= b and not a;
    outputs(4369) <= not a;
    outputs(4370) <= b;
    outputs(4371) <= a or b;
    outputs(4372) <= a and b;
    outputs(4373) <= a;
    outputs(4374) <= a;
    outputs(4375) <= b;
    outputs(4376) <= not a;
    outputs(4377) <= not a or b;
    outputs(4378) <= a xor b;
    outputs(4379) <= not (a xor b);
    outputs(4380) <= not (a xor b);
    outputs(4381) <= not a;
    outputs(4382) <= not a or b;
    outputs(4383) <= a xor b;
    outputs(4384) <= not (a or b);
    outputs(4385) <= a and b;
    outputs(4386) <= a and not b;
    outputs(4387) <= b;
    outputs(4388) <= not a;
    outputs(4389) <= a;
    outputs(4390) <= a;
    outputs(4391) <= a and not b;
    outputs(4392) <= not b or a;
    outputs(4393) <= a and b;
    outputs(4394) <= b;
    outputs(4395) <= a;
    outputs(4396) <= not (a xor b);
    outputs(4397) <= not (a xor b);
    outputs(4398) <= not a or b;
    outputs(4399) <= not a;
    outputs(4400) <= a and b;
    outputs(4401) <= not a;
    outputs(4402) <= not (a and b);
    outputs(4403) <= not b or a;
    outputs(4404) <= not b;
    outputs(4405) <= not (a and b);
    outputs(4406) <= b;
    outputs(4407) <= a;
    outputs(4408) <= not b;
    outputs(4409) <= a;
    outputs(4410) <= a xor b;
    outputs(4411) <= a xor b;
    outputs(4412) <= a xor b;
    outputs(4413) <= b and not a;
    outputs(4414) <= a and b;
    outputs(4415) <= not b or a;
    outputs(4416) <= b and not a;
    outputs(4417) <= not a;
    outputs(4418) <= b;
    outputs(4419) <= b;
    outputs(4420) <= not a or b;
    outputs(4421) <= not a;
    outputs(4422) <= not a or b;
    outputs(4423) <= a and b;
    outputs(4424) <= not (a and b);
    outputs(4425) <= a;
    outputs(4426) <= a and not b;
    outputs(4427) <= a xor b;
    outputs(4428) <= not b or a;
    outputs(4429) <= not (a and b);
    outputs(4430) <= not b;
    outputs(4431) <= not b or a;
    outputs(4432) <= not a;
    outputs(4433) <= not (a and b);
    outputs(4434) <= not a or b;
    outputs(4435) <= not b;
    outputs(4436) <= a xor b;
    outputs(4437) <= a;
    outputs(4438) <= not b;
    outputs(4439) <= b;
    outputs(4440) <= a xor b;
    outputs(4441) <= not b;
    outputs(4442) <= a xor b;
    outputs(4443) <= not a or b;
    outputs(4444) <= not (a xor b);
    outputs(4445) <= b;
    outputs(4446) <= not (a xor b);
    outputs(4447) <= not (a xor b);
    outputs(4448) <= not b;
    outputs(4449) <= b;
    outputs(4450) <= not a or b;
    outputs(4451) <= not a;
    outputs(4452) <= a or b;
    outputs(4453) <= b and not a;
    outputs(4454) <= a xor b;
    outputs(4455) <= not a;
    outputs(4456) <= a and not b;
    outputs(4457) <= a xor b;
    outputs(4458) <= not a;
    outputs(4459) <= b;
    outputs(4460) <= b;
    outputs(4461) <= not b;
    outputs(4462) <= not a;
    outputs(4463) <= a or b;
    outputs(4464) <= not b;
    outputs(4465) <= a;
    outputs(4466) <= a and b;
    outputs(4467) <= a;
    outputs(4468) <= not a;
    outputs(4469) <= not b;
    outputs(4470) <= a and b;
    outputs(4471) <= a;
    outputs(4472) <= not a;
    outputs(4473) <= not a;
    outputs(4474) <= not a;
    outputs(4475) <= not (a xor b);
    outputs(4476) <= b;
    outputs(4477) <= not (a or b);
    outputs(4478) <= a and not b;
    outputs(4479) <= not (a or b);
    outputs(4480) <= not a;
    outputs(4481) <= not (a or b);
    outputs(4482) <= b and not a;
    outputs(4483) <= a xor b;
    outputs(4484) <= not b;
    outputs(4485) <= not (a xor b);
    outputs(4486) <= not a or b;
    outputs(4487) <= b;
    outputs(4488) <= not b or a;
    outputs(4489) <= b;
    outputs(4490) <= b and not a;
    outputs(4491) <= a;
    outputs(4492) <= not (a xor b);
    outputs(4493) <= b and not a;
    outputs(4494) <= b and not a;
    outputs(4495) <= b and not a;
    outputs(4496) <= not a;
    outputs(4497) <= a or b;
    outputs(4498) <= not a;
    outputs(4499) <= a or b;
    outputs(4500) <= not b;
    outputs(4501) <= not a;
    outputs(4502) <= a;
    outputs(4503) <= not (a or b);
    outputs(4504) <= not b;
    outputs(4505) <= a;
    outputs(4506) <= not (a or b);
    outputs(4507) <= not b;
    outputs(4508) <= b;
    outputs(4509) <= not (a xor b);
    outputs(4510) <= a xor b;
    outputs(4511) <= b;
    outputs(4512) <= not (a and b);
    outputs(4513) <= a or b;
    outputs(4514) <= not (a xor b);
    outputs(4515) <= a;
    outputs(4516) <= not a or b;
    outputs(4517) <= not (a xor b);
    outputs(4518) <= a xor b;
    outputs(4519) <= not a or b;
    outputs(4520) <= a and not b;
    outputs(4521) <= b;
    outputs(4522) <= b;
    outputs(4523) <= not (a xor b);
    outputs(4524) <= not a;
    outputs(4525) <= not a or b;
    outputs(4526) <= not b;
    outputs(4527) <= not (a and b);
    outputs(4528) <= a;
    outputs(4529) <= b;
    outputs(4530) <= not b;
    outputs(4531) <= b;
    outputs(4532) <= a;
    outputs(4533) <= not a;
    outputs(4534) <= not b;
    outputs(4535) <= a and not b;
    outputs(4536) <= not a;
    outputs(4537) <= a;
    outputs(4538) <= not (a and b);
    outputs(4539) <= not (a xor b);
    outputs(4540) <= not (a xor b);
    outputs(4541) <= not a or b;
    outputs(4542) <= a and b;
    outputs(4543) <= not b;
    outputs(4544) <= not a;
    outputs(4545) <= b;
    outputs(4546) <= not b;
    outputs(4547) <= b;
    outputs(4548) <= a or b;
    outputs(4549) <= a;
    outputs(4550) <= b;
    outputs(4551) <= b;
    outputs(4552) <= a;
    outputs(4553) <= a;
    outputs(4554) <= a or b;
    outputs(4555) <= b and not a;
    outputs(4556) <= not (a or b);
    outputs(4557) <= a;
    outputs(4558) <= a;
    outputs(4559) <= a and not b;
    outputs(4560) <= not b;
    outputs(4561) <= b;
    outputs(4562) <= b and not a;
    outputs(4563) <= a xor b;
    outputs(4564) <= a xor b;
    outputs(4565) <= not (a and b);
    outputs(4566) <= a and not b;
    outputs(4567) <= not (a xor b);
    outputs(4568) <= not (a xor b);
    outputs(4569) <= b;
    outputs(4570) <= b;
    outputs(4571) <= a and b;
    outputs(4572) <= not (a xor b);
    outputs(4573) <= not (a xor b);
    outputs(4574) <= not (a or b);
    outputs(4575) <= a;
    outputs(4576) <= a and b;
    outputs(4577) <= b and not a;
    outputs(4578) <= not (a or b);
    outputs(4579) <= b and not a;
    outputs(4580) <= a xor b;
    outputs(4581) <= a xor b;
    outputs(4582) <= not (a and b);
    outputs(4583) <= not (a and b);
    outputs(4584) <= not (a xor b);
    outputs(4585) <= not b or a;
    outputs(4586) <= not b;
    outputs(4587) <= b and not a;
    outputs(4588) <= not a;
    outputs(4589) <= b;
    outputs(4590) <= b;
    outputs(4591) <= not b;
    outputs(4592) <= not b;
    outputs(4593) <= b;
    outputs(4594) <= not b;
    outputs(4595) <= a;
    outputs(4596) <= not a;
    outputs(4597) <= not b;
    outputs(4598) <= a;
    outputs(4599) <= not (a or b);
    outputs(4600) <= a;
    outputs(4601) <= not (a or b);
    outputs(4602) <= not (a xor b);
    outputs(4603) <= a;
    outputs(4604) <= a;
    outputs(4605) <= not b or a;
    outputs(4606) <= a;
    outputs(4607) <= a xor b;
    outputs(4608) <= a;
    outputs(4609) <= b and not a;
    outputs(4610) <= not b;
    outputs(4611) <= a xor b;
    outputs(4612) <= not (a or b);
    outputs(4613) <= a or b;
    outputs(4614) <= b;
    outputs(4615) <= not b;
    outputs(4616) <= a xor b;
    outputs(4617) <= not (a or b);
    outputs(4618) <= not (a xor b);
    outputs(4619) <= not (a xor b);
    outputs(4620) <= not (a xor b);
    outputs(4621) <= not a;
    outputs(4622) <= not (a xor b);
    outputs(4623) <= a and not b;
    outputs(4624) <= a and not b;
    outputs(4625) <= a and not b;
    outputs(4626) <= not (a xor b);
    outputs(4627) <= b and not a;
    outputs(4628) <= not (a and b);
    outputs(4629) <= a;
    outputs(4630) <= not a;
    outputs(4631) <= b and not a;
    outputs(4632) <= not (a xor b);
    outputs(4633) <= not (a or b);
    outputs(4634) <= b;
    outputs(4635) <= not (a xor b);
    outputs(4636) <= not a or b;
    outputs(4637) <= not a;
    outputs(4638) <= b;
    outputs(4639) <= b;
    outputs(4640) <= b;
    outputs(4641) <= not a;
    outputs(4642) <= a xor b;
    outputs(4643) <= a;
    outputs(4644) <= a;
    outputs(4645) <= a and not b;
    outputs(4646) <= a or b;
    outputs(4647) <= not a or b;
    outputs(4648) <= not (a or b);
    outputs(4649) <= not b;
    outputs(4650) <= not b or a;
    outputs(4651) <= a and b;
    outputs(4652) <= a and b;
    outputs(4653) <= b and not a;
    outputs(4654) <= not a;
    outputs(4655) <= a and not b;
    outputs(4656) <= not a or b;
    outputs(4657) <= a and not b;
    outputs(4658) <= a and not b;
    outputs(4659) <= a and not b;
    outputs(4660) <= a;
    outputs(4661) <= not (a xor b);
    outputs(4662) <= not (a xor b);
    outputs(4663) <= not (a or b);
    outputs(4664) <= not a;
    outputs(4665) <= not b;
    outputs(4666) <= not a or b;
    outputs(4667) <= not a;
    outputs(4668) <= a;
    outputs(4669) <= not b or a;
    outputs(4670) <= b;
    outputs(4671) <= a and b;
    outputs(4672) <= not (a or b);
    outputs(4673) <= b and not a;
    outputs(4674) <= a;
    outputs(4675) <= b and not a;
    outputs(4676) <= not (a and b);
    outputs(4677) <= not (a xor b);
    outputs(4678) <= a and b;
    outputs(4679) <= a xor b;
    outputs(4680) <= not (a or b);
    outputs(4681) <= not (a xor b);
    outputs(4682) <= a and not b;
    outputs(4683) <= b;
    outputs(4684) <= not (a xor b);
    outputs(4685) <= a;
    outputs(4686) <= b and not a;
    outputs(4687) <= not a;
    outputs(4688) <= b and not a;
    outputs(4689) <= b;
    outputs(4690) <= a xor b;
    outputs(4691) <= not b;
    outputs(4692) <= a and not b;
    outputs(4693) <= a;
    outputs(4694) <= b;
    outputs(4695) <= b;
    outputs(4696) <= not b or a;
    outputs(4697) <= not a;
    outputs(4698) <= not (a or b);
    outputs(4699) <= not (a or b);
    outputs(4700) <= not b;
    outputs(4701) <= b;
    outputs(4702) <= a;
    outputs(4703) <= a;
    outputs(4704) <= a xor b;
    outputs(4705) <= not (a xor b);
    outputs(4706) <= not (a or b);
    outputs(4707) <= not b;
    outputs(4708) <= a and not b;
    outputs(4709) <= a and b;
    outputs(4710) <= not a;
    outputs(4711) <= not (a xor b);
    outputs(4712) <= b;
    outputs(4713) <= a or b;
    outputs(4714) <= a xor b;
    outputs(4715) <= not a;
    outputs(4716) <= a and not b;
    outputs(4717) <= a and b;
    outputs(4718) <= not a;
    outputs(4719) <= b and not a;
    outputs(4720) <= a;
    outputs(4721) <= b;
    outputs(4722) <= b and not a;
    outputs(4723) <= a xor b;
    outputs(4724) <= a xor b;
    outputs(4725) <= a xor b;
    outputs(4726) <= a xor b;
    outputs(4727) <= not (a or b);
    outputs(4728) <= not b;
    outputs(4729) <= not (a or b);
    outputs(4730) <= not a;
    outputs(4731) <= a;
    outputs(4732) <= not (a or b);
    outputs(4733) <= not a;
    outputs(4734) <= not (a or b);
    outputs(4735) <= b and not a;
    outputs(4736) <= not b;
    outputs(4737) <= a and b;
    outputs(4738) <= not (a or b);
    outputs(4739) <= b and not a;
    outputs(4740) <= a and b;
    outputs(4741) <= b and not a;
    outputs(4742) <= not (a xor b);
    outputs(4743) <= a xor b;
    outputs(4744) <= not b;
    outputs(4745) <= a xor b;
    outputs(4746) <= b and not a;
    outputs(4747) <= not (a xor b);
    outputs(4748) <= a xor b;
    outputs(4749) <= not (a xor b);
    outputs(4750) <= a;
    outputs(4751) <= b and not a;
    outputs(4752) <= not (a or b);
    outputs(4753) <= a;
    outputs(4754) <= a and not b;
    outputs(4755) <= a xor b;
    outputs(4756) <= b;
    outputs(4757) <= b;
    outputs(4758) <= b;
    outputs(4759) <= not b;
    outputs(4760) <= a and not b;
    outputs(4761) <= a or b;
    outputs(4762) <= b;
    outputs(4763) <= a;
    outputs(4764) <= a xor b;
    outputs(4765) <= not (a or b);
    outputs(4766) <= not a;
    outputs(4767) <= b and not a;
    outputs(4768) <= not b;
    outputs(4769) <= not b;
    outputs(4770) <= a xor b;
    outputs(4771) <= not b;
    outputs(4772) <= not (a or b);
    outputs(4773) <= not (a and b);
    outputs(4774) <= not (a xor b);
    outputs(4775) <= a;
    outputs(4776) <= a and b;
    outputs(4777) <= not (a xor b);
    outputs(4778) <= a and not b;
    outputs(4779) <= not b or a;
    outputs(4780) <= a;
    outputs(4781) <= not (a xor b);
    outputs(4782) <= a xor b;
    outputs(4783) <= not b or a;
    outputs(4784) <= not (a xor b);
    outputs(4785) <= not a;
    outputs(4786) <= b;
    outputs(4787) <= not (a xor b);
    outputs(4788) <= b;
    outputs(4789) <= not a;
    outputs(4790) <= not (a xor b);
    outputs(4791) <= b;
    outputs(4792) <= not a or b;
    outputs(4793) <= a;
    outputs(4794) <= not (a xor b);
    outputs(4795) <= a and not b;
    outputs(4796) <= a xor b;
    outputs(4797) <= b;
    outputs(4798) <= b;
    outputs(4799) <= b;
    outputs(4800) <= not (a xor b);
    outputs(4801) <= a and b;
    outputs(4802) <= a xor b;
    outputs(4803) <= not (a or b);
    outputs(4804) <= a and not b;
    outputs(4805) <= a xor b;
    outputs(4806) <= not a;
    outputs(4807) <= not (a or b);
    outputs(4808) <= not a;
    outputs(4809) <= b and not a;
    outputs(4810) <= not (a xor b);
    outputs(4811) <= not b;
    outputs(4812) <= b;
    outputs(4813) <= a;
    outputs(4814) <= not a or b;
    outputs(4815) <= not a;
    outputs(4816) <= b;
    outputs(4817) <= b and not a;
    outputs(4818) <= a and b;
    outputs(4819) <= not (a or b);
    outputs(4820) <= a or b;
    outputs(4821) <= b;
    outputs(4822) <= not (a or b);
    outputs(4823) <= not a;
    outputs(4824) <= a;
    outputs(4825) <= a;
    outputs(4826) <= b and not a;
    outputs(4827) <= b;
    outputs(4828) <= not a;
    outputs(4829) <= not (a xor b);
    outputs(4830) <= a and not b;
    outputs(4831) <= a and b;
    outputs(4832) <= not (a xor b);
    outputs(4833) <= not b;
    outputs(4834) <= not (a xor b);
    outputs(4835) <= not b or a;
    outputs(4836) <= not b;
    outputs(4837) <= a xor b;
    outputs(4838) <= b;
    outputs(4839) <= not b;
    outputs(4840) <= not (a xor b);
    outputs(4841) <= a xor b;
    outputs(4842) <= a and not b;
    outputs(4843) <= a;
    outputs(4844) <= a and b;
    outputs(4845) <= a and not b;
    outputs(4846) <= a;
    outputs(4847) <= b;
    outputs(4848) <= a and b;
    outputs(4849) <= not a;
    outputs(4850) <= not (a or b);
    outputs(4851) <= not a;
    outputs(4852) <= a and not b;
    outputs(4853) <= b;
    outputs(4854) <= not (a xor b);
    outputs(4855) <= a and not b;
    outputs(4856) <= a or b;
    outputs(4857) <= a and not b;
    outputs(4858) <= b and not a;
    outputs(4859) <= a and b;
    outputs(4860) <= b;
    outputs(4861) <= b and not a;
    outputs(4862) <= a;
    outputs(4863) <= not b or a;
    outputs(4864) <= b and not a;
    outputs(4865) <= not (a or b);
    outputs(4866) <= b;
    outputs(4867) <= b;
    outputs(4868) <= not (a or b);
    outputs(4869) <= a;
    outputs(4870) <= a and not b;
    outputs(4871) <= not (a or b);
    outputs(4872) <= not a;
    outputs(4873) <= a and not b;
    outputs(4874) <= not b;
    outputs(4875) <= a;
    outputs(4876) <= not b;
    outputs(4877) <= a xor b;
    outputs(4878) <= not b;
    outputs(4879) <= not a;
    outputs(4880) <= not b or a;
    outputs(4881) <= b;
    outputs(4882) <= a and not b;
    outputs(4883) <= a or b;
    outputs(4884) <= not a;
    outputs(4885) <= not b;
    outputs(4886) <= b and not a;
    outputs(4887) <= a and not b;
    outputs(4888) <= not b;
    outputs(4889) <= not b;
    outputs(4890) <= not (a or b);
    outputs(4891) <= not (a or b);
    outputs(4892) <= a xor b;
    outputs(4893) <= not b;
    outputs(4894) <= not b or a;
    outputs(4895) <= a or b;
    outputs(4896) <= not (a and b);
    outputs(4897) <= not (a xor b);
    outputs(4898) <= not (a or b);
    outputs(4899) <= a and b;
    outputs(4900) <= a;
    outputs(4901) <= a or b;
    outputs(4902) <= a and not b;
    outputs(4903) <= a xor b;
    outputs(4904) <= not (a and b);
    outputs(4905) <= b and not a;
    outputs(4906) <= not a;
    outputs(4907) <= a xor b;
    outputs(4908) <= b;
    outputs(4909) <= a or b;
    outputs(4910) <= not a or b;
    outputs(4911) <= a and not b;
    outputs(4912) <= a and not b;
    outputs(4913) <= a and not b;
    outputs(4914) <= a;
    outputs(4915) <= b and not a;
    outputs(4916) <= a xor b;
    outputs(4917) <= not a;
    outputs(4918) <= a;
    outputs(4919) <= b;
    outputs(4920) <= not b;
    outputs(4921) <= a;
    outputs(4922) <= b;
    outputs(4923) <= a and b;
    outputs(4924) <= not b or a;
    outputs(4925) <= a and not b;
    outputs(4926) <= a xor b;
    outputs(4927) <= a and b;
    outputs(4928) <= a and b;
    outputs(4929) <= not (a or b);
    outputs(4930) <= not (a xor b);
    outputs(4931) <= not b;
    outputs(4932) <= not b;
    outputs(4933) <= not (a xor b);
    outputs(4934) <= b and not a;
    outputs(4935) <= b and not a;
    outputs(4936) <= a and b;
    outputs(4937) <= not (a or b);
    outputs(4938) <= not a;
    outputs(4939) <= a xor b;
    outputs(4940) <= not b;
    outputs(4941) <= not a or b;
    outputs(4942) <= not (a xor b);
    outputs(4943) <= a and b;
    outputs(4944) <= a and b;
    outputs(4945) <= b;
    outputs(4946) <= not (a or b);
    outputs(4947) <= a and not b;
    outputs(4948) <= b and not a;
    outputs(4949) <= not a;
    outputs(4950) <= a xor b;
    outputs(4951) <= not a;
    outputs(4952) <= not (a xor b);
    outputs(4953) <= b;
    outputs(4954) <= a and not b;
    outputs(4955) <= b;
    outputs(4956) <= a xor b;
    outputs(4957) <= b;
    outputs(4958) <= not (a xor b);
    outputs(4959) <= a xor b;
    outputs(4960) <= a and not b;
    outputs(4961) <= a and not b;
    outputs(4962) <= not (a or b);
    outputs(4963) <= a and not b;
    outputs(4964) <= b and not a;
    outputs(4965) <= a;
    outputs(4966) <= a xor b;
    outputs(4967) <= a and not b;
    outputs(4968) <= a xor b;
    outputs(4969) <= not (a xor b);
    outputs(4970) <= a;
    outputs(4971) <= a xor b;
    outputs(4972) <= b and not a;
    outputs(4973) <= not (a xor b);
    outputs(4974) <= not b;
    outputs(4975) <= not a;
    outputs(4976) <= a;
    outputs(4977) <= a and not b;
    outputs(4978) <= a or b;
    outputs(4979) <= not b;
    outputs(4980) <= a;
    outputs(4981) <= b and not a;
    outputs(4982) <= a and b;
    outputs(4983) <= a and not b;
    outputs(4984) <= a or b;
    outputs(4985) <= b and not a;
    outputs(4986) <= a;
    outputs(4987) <= b;
    outputs(4988) <= b and not a;
    outputs(4989) <= not (a xor b);
    outputs(4990) <= not b;
    outputs(4991) <= a xor b;
    outputs(4992) <= b and not a;
    outputs(4993) <= a xor b;
    outputs(4994) <= b and not a;
    outputs(4995) <= a and b;
    outputs(4996) <= a xor b;
    outputs(4997) <= not (a and b);
    outputs(4998) <= b;
    outputs(4999) <= a;
    outputs(5000) <= not a or b;
    outputs(5001) <= a and not b;
    outputs(5002) <= b and not a;
    outputs(5003) <= b;
    outputs(5004) <= not (a xor b);
    outputs(5005) <= not b;
    outputs(5006) <= b;
    outputs(5007) <= not (a or b);
    outputs(5008) <= a and b;
    outputs(5009) <= a;
    outputs(5010) <= b;
    outputs(5011) <= not b;
    outputs(5012) <= b;
    outputs(5013) <= a xor b;
    outputs(5014) <= a and not b;
    outputs(5015) <= not (a xor b);
    outputs(5016) <= a and b;
    outputs(5017) <= not b;
    outputs(5018) <= not (a or b);
    outputs(5019) <= a and b;
    outputs(5020) <= a and b;
    outputs(5021) <= not b;
    outputs(5022) <= not (a or b);
    outputs(5023) <= not (a xor b);
    outputs(5024) <= a and not b;
    outputs(5025) <= a xor b;
    outputs(5026) <= a xor b;
    outputs(5027) <= not b;
    outputs(5028) <= b and not a;
    outputs(5029) <= not b;
    outputs(5030) <= b;
    outputs(5031) <= not (a or b);
    outputs(5032) <= not (a xor b);
    outputs(5033) <= not b;
    outputs(5034) <= a and not b;
    outputs(5035) <= a;
    outputs(5036) <= a xor b;
    outputs(5037) <= b;
    outputs(5038) <= not b;
    outputs(5039) <= not (a or b);
    outputs(5040) <= not b;
    outputs(5041) <= a and not b;
    outputs(5042) <= a xor b;
    outputs(5043) <= not a;
    outputs(5044) <= not b;
    outputs(5045) <= b;
    outputs(5046) <= not b;
    outputs(5047) <= a and not b;
    outputs(5048) <= not b;
    outputs(5049) <= a and not b;
    outputs(5050) <= b and not a;
    outputs(5051) <= not a;
    outputs(5052) <= not (a xor b);
    outputs(5053) <= not a or b;
    outputs(5054) <= a;
    outputs(5055) <= not (a and b);
    outputs(5056) <= not b;
    outputs(5057) <= not b;
    outputs(5058) <= a;
    outputs(5059) <= not (a or b);
    outputs(5060) <= a and not b;
    outputs(5061) <= not (a or b);
    outputs(5062) <= b and not a;
    outputs(5063) <= not a or b;
    outputs(5064) <= a;
    outputs(5065) <= a;
    outputs(5066) <= a xor b;
    outputs(5067) <= a xor b;
    outputs(5068) <= not a;
    outputs(5069) <= a;
    outputs(5070) <= not b;
    outputs(5071) <= not b;
    outputs(5072) <= not (a xor b);
    outputs(5073) <= not (a or b);
    outputs(5074) <= a;
    outputs(5075) <= a;
    outputs(5076) <= a and b;
    outputs(5077) <= a xor b;
    outputs(5078) <= a or b;
    outputs(5079) <= not b;
    outputs(5080) <= not a;
    outputs(5081) <= a and not b;
    outputs(5082) <= b and not a;
    outputs(5083) <= not b;
    outputs(5084) <= a;
    outputs(5085) <= not a or b;
    outputs(5086) <= b and not a;
    outputs(5087) <= b and not a;
    outputs(5088) <= a;
    outputs(5089) <= a;
    outputs(5090) <= b;
    outputs(5091) <= a and not b;
    outputs(5092) <= not (a xor b);
    outputs(5093) <= not b;
    outputs(5094) <= a and b;
    outputs(5095) <= b;
    outputs(5096) <= not (a or b);
    outputs(5097) <= b;
    outputs(5098) <= b and not a;
    outputs(5099) <= a;
    outputs(5100) <= not a;
    outputs(5101) <= not b or a;
    outputs(5102) <= not a or b;
    outputs(5103) <= b and not a;
    outputs(5104) <= a;
    outputs(5105) <= not a;
    outputs(5106) <= a and b;
    outputs(5107) <= not b;
    outputs(5108) <= not (a or b);
    outputs(5109) <= a;
    outputs(5110) <= not a or b;
    outputs(5111) <= not b;
    outputs(5112) <= b;
    outputs(5113) <= a and not b;
    outputs(5114) <= not (a xor b);
    outputs(5115) <= not (a xor b);
    outputs(5116) <= not a;
    outputs(5117) <= not (a or b);
    outputs(5118) <= not b;
    outputs(5119) <= not (a or b);
end Behavioral;
